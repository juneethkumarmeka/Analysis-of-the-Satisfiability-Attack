module basic_5000_50000_5000_5_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nand U0 (N_0,In_2819,In_1434);
xor U1 (N_1,In_4767,In_880);
nand U2 (N_2,In_3822,In_3728);
and U3 (N_3,In_3398,In_4773);
xnor U4 (N_4,In_4855,In_23);
xor U5 (N_5,In_73,In_405);
nand U6 (N_6,In_29,In_2909);
or U7 (N_7,In_1593,In_887);
nor U8 (N_8,In_4113,In_1576);
and U9 (N_9,In_4971,In_3482);
nand U10 (N_10,In_4228,In_1038);
xnor U11 (N_11,In_245,In_3365);
xnor U12 (N_12,In_1879,In_515);
nand U13 (N_13,In_3669,In_651);
nor U14 (N_14,In_674,In_507);
nand U15 (N_15,In_766,In_2446);
xor U16 (N_16,In_1603,In_3154);
or U17 (N_17,In_1435,In_3668);
nand U18 (N_18,In_1983,In_2539);
and U19 (N_19,In_4571,In_2675);
nor U20 (N_20,In_3520,In_2850);
xnor U21 (N_21,In_3255,In_4827);
and U22 (N_22,In_1343,In_4628);
nor U23 (N_23,In_2105,In_2740);
xnor U24 (N_24,In_2842,In_4487);
or U25 (N_25,In_4106,In_3132);
nor U26 (N_26,In_1242,In_4050);
xnor U27 (N_27,In_3581,In_2001);
or U28 (N_28,In_2508,In_3713);
xor U29 (N_29,In_4423,In_1499);
and U30 (N_30,In_217,In_2219);
nand U31 (N_31,In_1536,In_792);
nor U32 (N_32,In_2989,In_3552);
nand U33 (N_33,In_1075,In_1243);
xor U34 (N_34,In_2235,In_1862);
nand U35 (N_35,In_1590,In_3051);
or U36 (N_36,In_3362,In_3468);
xnor U37 (N_37,In_1975,In_2527);
nor U38 (N_38,In_2249,In_3896);
or U39 (N_39,In_3428,In_122);
xnor U40 (N_40,In_3211,In_2595);
or U41 (N_41,In_51,In_3408);
or U42 (N_42,In_4616,In_2845);
xor U43 (N_43,In_829,In_2283);
and U44 (N_44,In_192,In_4021);
nor U45 (N_45,In_4730,In_2182);
xor U46 (N_46,In_1269,In_3329);
nand U47 (N_47,In_2829,In_585);
nor U48 (N_48,In_1699,In_1552);
xor U49 (N_49,In_4499,In_2672);
nand U50 (N_50,In_4999,In_1107);
xnor U51 (N_51,In_4706,In_2493);
and U52 (N_52,In_4359,In_270);
or U53 (N_53,In_4196,In_3129);
nand U54 (N_54,In_438,In_2003);
and U55 (N_55,In_4932,In_35);
nor U56 (N_56,In_693,In_1199);
xor U57 (N_57,In_2149,In_3455);
xnor U58 (N_58,In_1511,In_3002);
or U59 (N_59,In_3740,In_599);
nand U60 (N_60,In_3662,In_1755);
nor U61 (N_61,In_3445,In_1870);
nand U62 (N_62,In_2621,In_2);
nor U63 (N_63,In_2005,In_2949);
nand U64 (N_64,In_4047,In_571);
or U65 (N_65,In_4335,In_1047);
and U66 (N_66,In_4379,In_162);
xor U67 (N_67,In_38,In_3845);
or U68 (N_68,In_1407,In_732);
xor U69 (N_69,In_4116,In_4655);
nor U70 (N_70,In_4131,In_1144);
xnor U71 (N_71,In_3157,In_2831);
and U72 (N_72,In_1664,In_4143);
xnor U73 (N_73,In_2253,In_2677);
xnor U74 (N_74,In_2919,In_4702);
nand U75 (N_75,In_784,In_2967);
nand U76 (N_76,In_3328,In_740);
xor U77 (N_77,In_1646,In_2368);
nor U78 (N_78,In_2222,In_2168);
nor U79 (N_79,In_2029,In_2280);
nand U80 (N_80,In_2440,In_1145);
and U81 (N_81,In_2987,In_2132);
xnor U82 (N_82,In_3017,In_2087);
and U83 (N_83,In_4604,In_452);
nand U84 (N_84,In_4358,In_3931);
xnor U85 (N_85,In_4124,In_128);
nor U86 (N_86,In_2646,In_2101);
and U87 (N_87,In_4251,In_3401);
or U88 (N_88,In_812,In_2510);
xnor U89 (N_89,In_2973,In_746);
and U90 (N_90,In_3557,In_2543);
xor U91 (N_91,In_3433,In_44);
or U92 (N_92,In_4274,In_606);
xor U93 (N_93,In_2802,In_3969);
nand U94 (N_94,In_269,In_4919);
nand U95 (N_95,In_2433,In_4204);
nor U96 (N_96,In_4667,In_3603);
xor U97 (N_97,In_1017,In_2504);
xnor U98 (N_98,In_431,In_1829);
nor U99 (N_99,In_1609,In_3864);
nand U100 (N_100,In_512,In_479);
xor U101 (N_101,In_3039,In_605);
nand U102 (N_102,In_4085,In_4651);
nor U103 (N_103,In_2277,In_3608);
nor U104 (N_104,In_2955,In_1373);
nor U105 (N_105,In_226,In_2801);
xnor U106 (N_106,In_1201,In_1185);
nor U107 (N_107,In_232,In_2478);
nor U108 (N_108,In_439,In_3184);
and U109 (N_109,In_2158,In_345);
or U110 (N_110,In_809,In_4237);
or U111 (N_111,In_4502,In_3617);
nor U112 (N_112,In_3403,In_621);
nor U113 (N_113,In_1789,In_1337);
nor U114 (N_114,In_4843,In_1284);
or U115 (N_115,In_3963,In_1495);
nor U116 (N_116,In_3402,In_4012);
or U117 (N_117,In_2995,In_1830);
xnor U118 (N_118,In_109,In_1375);
or U119 (N_119,In_3673,In_4275);
nor U120 (N_120,In_475,In_3676);
nand U121 (N_121,In_3835,In_4447);
and U122 (N_122,In_3061,In_4213);
xor U123 (N_123,In_2361,In_1167);
nor U124 (N_124,In_1106,In_1541);
xor U125 (N_125,In_542,In_2847);
or U126 (N_126,In_158,In_3330);
or U127 (N_127,In_4852,In_319);
nor U128 (N_128,In_4534,In_3000);
nor U129 (N_129,In_2913,In_2922);
nand U130 (N_130,In_2934,In_4581);
nand U131 (N_131,In_2771,In_3201);
or U132 (N_132,In_731,In_1124);
xnor U133 (N_133,In_259,In_1503);
nor U134 (N_134,In_4829,In_4067);
nor U135 (N_135,In_851,In_3353);
and U136 (N_136,In_4775,In_4090);
or U137 (N_137,In_4300,In_4934);
nor U138 (N_138,In_4301,In_642);
nor U139 (N_139,In_2221,In_4678);
and U140 (N_140,In_3757,In_2367);
nor U141 (N_141,In_2747,In_4974);
nor U142 (N_142,In_87,In_1923);
xor U143 (N_143,In_4191,In_3674);
or U144 (N_144,In_1631,In_3786);
nand U145 (N_145,In_957,In_85);
nor U146 (N_146,In_785,In_3653);
nor U147 (N_147,In_1449,In_2920);
nor U148 (N_148,In_3092,In_627);
nor U149 (N_149,In_3553,In_4685);
and U150 (N_150,In_1611,In_2820);
or U151 (N_151,In_64,In_2560);
xnor U152 (N_152,In_2971,In_2661);
and U153 (N_153,In_3773,In_3332);
nand U154 (N_154,In_2898,In_2507);
and U155 (N_155,In_1594,In_407);
nor U156 (N_156,In_2725,In_3677);
nor U157 (N_157,In_1143,In_3271);
and U158 (N_158,In_3776,In_2320);
or U159 (N_159,In_3506,In_3731);
nor U160 (N_160,In_4327,In_4283);
nor U161 (N_161,In_22,In_4178);
and U162 (N_162,In_1384,In_1223);
nand U163 (N_163,In_3885,In_1648);
nand U164 (N_164,In_2393,In_1818);
or U165 (N_165,In_4620,In_497);
nor U166 (N_166,In_1527,In_853);
or U167 (N_167,In_3366,In_3256);
nor U168 (N_168,In_3264,In_2274);
or U169 (N_169,In_4378,In_4916);
nand U170 (N_170,In_4698,In_2805);
and U171 (N_171,In_1355,In_3796);
and U172 (N_172,In_4060,In_4874);
xor U173 (N_173,In_2714,In_3452);
xor U174 (N_174,In_959,In_3216);
xnor U175 (N_175,In_883,In_3208);
nand U176 (N_176,In_1005,In_1799);
nand U177 (N_177,In_1994,In_2051);
nand U178 (N_178,In_4026,In_3381);
or U179 (N_179,In_4809,In_4710);
nand U180 (N_180,In_534,In_1558);
nand U181 (N_181,In_3373,In_3869);
xor U182 (N_182,In_4167,In_4933);
xnor U183 (N_183,In_796,In_3344);
or U184 (N_184,In_327,In_91);
nor U185 (N_185,In_969,In_838);
and U186 (N_186,In_1087,In_2759);
xor U187 (N_187,In_547,In_2389);
xnor U188 (N_188,In_4192,In_645);
xor U189 (N_189,In_981,In_1441);
nor U190 (N_190,In_3269,In_2064);
nor U191 (N_191,In_100,In_1131);
or U192 (N_192,In_2216,In_978);
nor U193 (N_193,In_2945,In_3592);
or U194 (N_194,In_2080,In_4878);
nor U195 (N_195,In_2142,In_4492);
or U196 (N_196,In_460,In_1346);
nor U197 (N_197,In_3546,In_2653);
xnor U198 (N_198,In_3912,In_1625);
or U199 (N_199,In_1857,In_1283);
xnor U200 (N_200,In_963,In_4430);
and U201 (N_201,In_4304,In_1200);
nand U202 (N_202,In_708,In_4324);
xor U203 (N_203,In_4579,In_419);
nand U204 (N_204,In_1379,In_1888);
nor U205 (N_205,In_4170,In_3347);
nand U206 (N_206,In_4136,In_230);
nor U207 (N_207,In_3315,In_4253);
and U208 (N_208,In_488,In_3792);
xor U209 (N_209,In_1127,In_3503);
or U210 (N_210,In_3620,In_4076);
nand U211 (N_211,In_2438,In_4294);
xor U212 (N_212,In_4794,In_4724);
and U213 (N_213,In_1986,In_404);
nor U214 (N_214,In_758,In_1657);
nand U215 (N_215,In_3739,In_2376);
nor U216 (N_216,In_678,In_4466);
or U217 (N_217,In_2115,In_4104);
and U218 (N_218,In_1610,In_924);
and U219 (N_219,In_2822,In_1917);
xnor U220 (N_220,In_46,In_1619);
or U221 (N_221,In_3294,In_4406);
nand U222 (N_222,In_3029,In_1866);
or U223 (N_223,In_1703,In_3938);
nand U224 (N_224,In_3656,In_3508);
nand U225 (N_225,In_2727,In_3724);
nand U226 (N_226,In_4397,In_2636);
nand U227 (N_227,In_4473,In_209);
and U228 (N_228,In_4326,In_2745);
and U229 (N_229,In_1754,In_1961);
and U230 (N_230,In_4547,In_4210);
or U231 (N_231,In_1976,In_494);
xor U232 (N_232,In_3016,In_2015);
or U233 (N_233,In_4478,In_3479);
xor U234 (N_234,In_3429,In_1523);
or U235 (N_235,In_2194,In_4781);
and U236 (N_236,In_114,In_2624);
and U237 (N_237,In_1876,In_2057);
or U238 (N_238,In_1007,In_2983);
nand U239 (N_239,In_890,In_2673);
and U240 (N_240,In_2021,In_359);
nand U241 (N_241,In_381,In_4558);
and U242 (N_242,In_4778,In_1216);
or U243 (N_243,In_4911,In_3743);
nand U244 (N_244,In_2710,In_1544);
nor U245 (N_245,In_2642,In_2263);
nor U246 (N_246,In_4238,In_3231);
and U247 (N_247,In_15,In_1908);
or U248 (N_248,In_3512,In_4688);
nand U249 (N_249,In_2326,In_1710);
xnor U250 (N_250,In_4647,In_176);
and U251 (N_251,In_3040,In_17);
nor U252 (N_252,In_2887,In_3317);
nor U253 (N_253,In_2649,In_4004);
nor U254 (N_254,In_2900,In_3139);
nor U255 (N_255,In_3660,In_194);
nand U256 (N_256,In_2117,In_397);
nand U257 (N_257,In_4519,In_1898);
or U258 (N_258,In_1309,In_2704);
xnor U259 (N_259,In_4316,In_4930);
xnor U260 (N_260,In_2840,In_3680);
and U261 (N_261,In_2996,In_1171);
nand U262 (N_262,In_1068,In_3838);
xnor U263 (N_263,In_3371,In_2223);
nor U264 (N_264,In_3910,In_2529);
xnor U265 (N_265,In_828,In_4340);
nand U266 (N_266,In_1993,In_2733);
nor U267 (N_267,In_1341,In_4446);
xor U268 (N_268,In_4037,In_1746);
and U269 (N_269,In_968,In_1484);
and U270 (N_270,In_1275,In_221);
and U271 (N_271,In_3,In_3424);
nand U272 (N_272,In_4491,In_4783);
or U273 (N_273,In_843,In_4469);
xnor U274 (N_274,In_4239,In_4858);
nor U275 (N_275,In_3204,In_997);
or U276 (N_276,In_4943,In_2520);
and U277 (N_277,In_1860,In_63);
nand U278 (N_278,In_2668,In_1585);
or U279 (N_279,In_4675,In_273);
nor U280 (N_280,In_491,In_244);
nand U281 (N_281,In_4895,In_6);
nand U282 (N_282,In_2450,In_1874);
or U283 (N_283,In_47,In_313);
and U284 (N_284,In_3238,In_1924);
and U285 (N_285,In_1996,In_1489);
nand U286 (N_286,In_3149,In_2550);
nand U287 (N_287,In_4583,In_3405);
nor U288 (N_288,In_1230,In_1388);
xnor U289 (N_289,In_4811,In_3960);
and U290 (N_290,In_1638,In_2036);
xnor U291 (N_291,In_2776,In_2917);
or U292 (N_292,In_2127,In_954);
or U293 (N_293,In_2839,In_3984);
and U294 (N_294,In_303,In_2106);
xor U295 (N_295,In_1026,In_522);
nand U296 (N_296,In_4684,In_4433);
xnor U297 (N_297,In_3529,In_735);
nor U298 (N_298,In_2757,In_805);
nor U299 (N_299,In_1372,In_3339);
and U300 (N_300,In_4789,In_3666);
nor U301 (N_301,In_3397,In_3919);
nand U302 (N_302,In_2939,In_1479);
nor U303 (N_303,In_24,In_4475);
nor U304 (N_304,In_2028,In_2122);
nand U305 (N_305,In_3823,In_1922);
nand U306 (N_306,In_349,In_2738);
nand U307 (N_307,In_2120,In_388);
xnor U308 (N_308,In_3011,In_4841);
or U309 (N_309,In_4642,In_323);
and U310 (N_310,In_976,In_1316);
or U311 (N_311,In_590,In_932);
nor U312 (N_312,In_1121,In_1166);
nor U313 (N_313,In_1240,In_4453);
xor U314 (N_314,In_1405,In_2655);
or U315 (N_315,In_2144,In_3357);
nand U316 (N_316,In_369,In_2734);
and U317 (N_317,In_117,In_2578);
xor U318 (N_318,In_4205,In_3214);
xnor U319 (N_319,In_416,In_3057);
xnor U320 (N_320,In_712,In_3809);
or U321 (N_321,In_3649,In_4312);
xnor U322 (N_322,In_1367,In_3251);
nand U323 (N_323,In_4471,In_2399);
and U324 (N_324,In_912,In_3215);
nand U325 (N_325,In_3037,In_223);
nor U326 (N_326,In_1488,In_4859);
or U327 (N_327,In_265,In_4649);
nand U328 (N_328,In_3393,In_3941);
nor U329 (N_329,In_188,In_1728);
and U330 (N_330,In_4162,In_1000);
or U331 (N_331,In_2644,In_4603);
nand U332 (N_332,In_3582,In_1324);
and U333 (N_333,In_164,In_1120);
nor U334 (N_334,In_3987,In_1759);
xor U335 (N_335,In_4554,In_3693);
or U336 (N_336,In_206,In_43);
or U337 (N_337,In_3654,In_1852);
and U338 (N_338,In_3642,In_837);
nor U339 (N_339,In_2855,In_425);
xnor U340 (N_340,In_500,In_482);
nor U341 (N_341,In_3052,In_2824);
and U342 (N_342,In_478,In_2960);
nand U343 (N_343,In_3534,In_710);
nand U344 (N_344,In_1482,In_560);
nor U345 (N_345,In_533,In_242);
and U346 (N_346,In_926,In_2910);
xnor U347 (N_347,In_1767,In_4606);
xor U348 (N_348,In_2310,In_596);
nor U349 (N_349,In_4721,In_1285);
and U350 (N_350,In_3527,In_2515);
or U351 (N_351,In_4753,In_1861);
xnor U352 (N_352,In_1859,In_734);
nand U353 (N_353,In_871,In_3417);
nor U354 (N_354,In_2085,In_211);
or U355 (N_355,In_2071,In_846);
nand U356 (N_356,In_282,In_1605);
and U357 (N_357,In_2506,In_2108);
xnor U358 (N_358,In_2359,In_324);
or U359 (N_359,In_3537,In_527);
nand U360 (N_360,In_3391,In_4262);
or U361 (N_361,In_4184,In_2075);
or U362 (N_362,In_4850,In_4736);
nand U363 (N_363,In_518,In_611);
xnor U364 (N_364,In_1249,In_3262);
nand U365 (N_365,In_2549,In_4008);
nand U366 (N_366,In_103,In_4907);
nand U367 (N_367,In_703,In_2882);
xor U368 (N_368,In_2525,In_1785);
nand U369 (N_369,In_318,In_4799);
nand U370 (N_370,In_2709,In_1615);
and U371 (N_371,In_640,In_4381);
nand U372 (N_372,In_1915,In_930);
nor U373 (N_373,In_2395,In_827);
or U374 (N_374,In_4777,In_3406);
nor U375 (N_375,In_3273,In_3156);
nand U376 (N_376,In_2240,In_748);
and U377 (N_377,In_2712,In_3022);
and U378 (N_378,In_240,In_810);
or U379 (N_379,In_689,In_2289);
or U380 (N_380,In_506,In_1190);
xnor U381 (N_381,In_3863,In_53);
and U382 (N_382,In_1140,In_4278);
or U383 (N_383,In_3672,In_695);
or U384 (N_384,In_4595,In_4297);
xnor U385 (N_385,In_262,In_935);
or U386 (N_386,In_4810,In_2041);
nor U387 (N_387,In_4966,In_1307);
nor U388 (N_388,In_95,In_3470);
or U389 (N_389,In_2279,In_3291);
nand U390 (N_390,In_4230,In_1639);
and U391 (N_391,In_423,In_3049);
nor U392 (N_392,In_4816,In_3980);
nand U393 (N_393,In_2159,In_4861);
nand U394 (N_394,In_4769,In_3112);
or U395 (N_395,In_1538,In_4224);
nand U396 (N_396,In_4339,In_3952);
nand U397 (N_397,In_1053,In_2889);
or U398 (N_398,In_3663,In_4483);
xor U399 (N_399,In_3778,In_3521);
nor U400 (N_400,In_408,In_1058);
nor U401 (N_401,In_4498,In_3278);
nor U402 (N_402,In_1687,In_2927);
and U403 (N_403,In_891,In_4069);
xnor U404 (N_404,In_3986,In_905);
xnor U405 (N_405,In_1039,In_2301);
xor U406 (N_406,In_2626,In_3383);
nor U407 (N_407,In_3093,In_331);
nor U408 (N_408,In_4972,In_34);
xor U409 (N_409,In_1587,In_3538);
and U410 (N_410,In_3545,In_1278);
nor U411 (N_411,In_698,In_3684);
xor U412 (N_412,In_402,In_3193);
nor U413 (N_413,In_4015,In_4893);
or U414 (N_414,In_2435,In_1276);
and U415 (N_415,In_4140,In_4656);
or U416 (N_416,In_4477,In_683);
nand U417 (N_417,In_4699,In_2942);
xnor U418 (N_418,In_2979,In_1747);
xnor U419 (N_419,In_2488,In_2573);
or U420 (N_420,In_2706,In_3004);
nand U421 (N_421,In_1690,In_1947);
nor U422 (N_422,In_2137,In_1310);
xnor U423 (N_423,In_2705,In_1842);
nand U424 (N_424,In_4520,In_3075);
nor U425 (N_425,In_275,In_304);
xnor U426 (N_426,In_3060,In_3694);
and U427 (N_427,In_3095,In_2016);
or U428 (N_428,In_2147,In_1914);
xor U429 (N_429,In_2189,In_3058);
and U430 (N_430,In_4095,In_675);
and U431 (N_431,In_4209,In_4577);
or U432 (N_432,In_2095,In_581);
nor U433 (N_433,In_4399,In_412);
nand U434 (N_434,In_1694,In_3179);
nor U435 (N_435,In_3631,In_915);
nor U436 (N_436,In_4942,In_4059);
and U437 (N_437,In_815,In_2566);
and U438 (N_438,In_1850,In_156);
or U439 (N_439,In_4232,In_1073);
nor U440 (N_440,In_3070,In_1612);
nor U441 (N_441,In_2449,In_544);
and U442 (N_442,In_3504,In_2766);
nor U443 (N_443,In_3472,In_4121);
nand U444 (N_444,In_4017,In_4034);
nand U445 (N_445,In_4006,In_1526);
nor U446 (N_446,In_636,In_2724);
nor U447 (N_447,In_297,In_2412);
nor U448 (N_448,In_2584,In_3804);
nand U449 (N_449,In_3426,In_4005);
and U450 (N_450,In_60,In_662);
and U451 (N_451,In_2143,In_634);
xnor U452 (N_452,In_4996,In_3150);
xor U453 (N_453,In_2492,In_802);
and U454 (N_454,In_3114,In_3410);
nor U455 (N_455,In_2201,In_3542);
nor U456 (N_456,In_4757,In_2225);
and U457 (N_457,In_3247,In_1882);
xor U458 (N_458,In_2294,In_551);
xor U459 (N_459,In_2414,In_1682);
nor U460 (N_460,In_4389,In_1551);
or U461 (N_461,In_548,In_559);
xor U462 (N_462,In_2031,In_2116);
nor U463 (N_463,In_308,In_1164);
or U464 (N_464,In_3828,In_3050);
nor U465 (N_465,In_4640,In_4485);
nand U466 (N_466,In_4556,In_806);
nor U467 (N_467,In_789,In_3942);
and U468 (N_468,In_437,In_937);
or U469 (N_469,In_3103,In_3888);
nor U470 (N_470,In_3842,In_3734);
nand U471 (N_471,In_2073,In_4803);
nand U472 (N_472,In_2247,In_2683);
and U473 (N_473,In_2770,In_1035);
or U474 (N_474,In_4635,In_2717);
or U475 (N_475,In_3242,In_2811);
or U476 (N_476,In_649,In_1505);
nor U477 (N_477,In_260,In_2443);
or U478 (N_478,In_3925,In_4780);
nor U479 (N_479,In_1466,In_3737);
nor U480 (N_480,In_3024,In_487);
nand U481 (N_481,In_676,In_4716);
nand U482 (N_482,In_4202,In_4719);
or U483 (N_483,In_1598,In_3812);
nor U484 (N_484,In_3361,In_1467);
or U485 (N_485,In_1776,In_3342);
nor U486 (N_486,In_2832,In_2447);
or U487 (N_487,In_1084,In_236);
nor U488 (N_488,In_1832,In_196);
or U489 (N_489,In_1030,In_3687);
or U490 (N_490,In_3783,In_4686);
xor U491 (N_491,In_4515,In_4646);
xor U492 (N_492,In_1041,In_2089);
nand U493 (N_493,In_3732,In_893);
nor U494 (N_494,In_3126,In_1351);
xor U495 (N_495,In_4882,In_45);
or U496 (N_496,In_2070,In_3300);
nor U497 (N_497,In_4985,In_2030);
nand U498 (N_498,In_562,In_3892);
or U499 (N_499,In_3413,In_2444);
nor U500 (N_500,In_1938,In_4681);
nand U501 (N_501,In_1032,In_2735);
xor U502 (N_502,In_2422,In_1439);
nand U503 (N_503,In_3003,In_3277);
or U504 (N_504,In_102,In_1504);
xnor U505 (N_505,In_1192,In_4052);
nor U506 (N_506,In_4369,In_1327);
and U507 (N_507,In_1116,In_2690);
or U508 (N_508,In_4514,In_3736);
and U509 (N_509,In_724,In_1863);
or U510 (N_510,In_3370,In_4174);
xor U511 (N_511,In_2613,In_2769);
or U512 (N_512,In_4820,In_2176);
nand U513 (N_513,In_4695,In_1067);
and U514 (N_514,In_3906,In_3511);
and U515 (N_515,In_4391,In_2755);
nand U516 (N_516,In_4043,In_4914);
nand U517 (N_517,In_3140,In_3021);
or U518 (N_518,In_1298,In_1193);
nand U519 (N_519,In_2135,In_2916);
and U520 (N_520,In_4877,In_1608);
nor U521 (N_521,In_4036,In_1114);
or U522 (N_522,In_1008,In_577);
or U523 (N_523,In_4525,In_2869);
nor U524 (N_524,In_3257,In_1119);
nor U525 (N_525,In_2808,In_2431);
or U526 (N_526,In_1793,In_739);
and U527 (N_527,In_1214,In_2401);
nor U528 (N_528,In_3120,In_2929);
nor U529 (N_529,In_797,In_2411);
or U530 (N_530,In_1202,In_4917);
xor U531 (N_531,In_3167,In_76);
and U532 (N_532,In_2061,In_33);
or U533 (N_533,In_2055,In_4445);
and U534 (N_534,In_4467,In_207);
nand U535 (N_535,In_844,In_3715);
or U536 (N_536,In_3355,In_4308);
xor U537 (N_537,In_637,In_1456);
nand U538 (N_538,In_4458,In_3974);
or U539 (N_539,In_4127,In_4311);
and U540 (N_540,In_2591,In_2930);
nand U541 (N_541,In_3905,In_4051);
and U542 (N_542,In_3624,In_384);
and U543 (N_543,In_1903,In_1797);
and U544 (N_544,In_3703,In_1021);
nor U545 (N_545,In_2352,In_2325);
xor U546 (N_546,In_4845,In_1258);
xor U547 (N_547,In_664,In_4956);
nor U548 (N_548,In_867,In_3042);
nor U549 (N_549,In_2139,In_2564);
and U550 (N_550,In_266,In_3758);
or U551 (N_551,In_903,In_252);
nand U552 (N_552,In_3182,In_3130);
or U553 (N_553,In_410,In_3733);
or U554 (N_554,In_775,In_2637);
or U555 (N_555,In_4885,In_171);
nor U556 (N_556,In_2157,In_955);
nor U557 (N_557,In_1779,In_1497);
nand U558 (N_558,In_1618,In_4030);
and U559 (N_559,In_3164,In_4997);
xnor U560 (N_560,In_1623,In_1239);
or U561 (N_561,In_4918,In_2551);
nor U562 (N_562,In_2275,In_1233);
or U563 (N_563,In_4134,In_2963);
xnor U564 (N_564,In_639,In_2282);
nand U565 (N_565,In_1656,In_4976);
xor U566 (N_566,In_4559,In_4098);
xnor U567 (N_567,In_1622,In_3948);
xnor U568 (N_568,In_4435,In_2475);
nand U569 (N_569,In_4263,In_1386);
xnor U570 (N_570,In_4153,In_3558);
or U571 (N_571,In_1323,In_718);
xnor U572 (N_572,In_1264,In_3720);
or U573 (N_573,In_1142,In_3759);
and U574 (N_574,In_1052,In_1913);
or U575 (N_575,In_119,In_579);
nand U576 (N_576,In_646,In_1393);
nand U577 (N_577,In_3258,In_4225);
xnor U578 (N_578,In_3889,In_1224);
nand U579 (N_579,In_3437,In_286);
nor U580 (N_580,In_233,In_4876);
xor U581 (N_581,In_2397,In_2448);
nor U582 (N_582,In_3138,In_4835);
nor U583 (N_583,In_4227,In_2849);
nand U584 (N_584,In_1380,In_174);
nand U585 (N_585,In_3566,In_2437);
and U586 (N_586,In_4284,In_1387);
nand U587 (N_587,In_4982,In_3219);
or U588 (N_588,In_1952,In_2796);
xnor U589 (N_589,In_1838,In_4958);
and U590 (N_590,In_3585,In_771);
and U591 (N_591,In_1071,In_2104);
nand U592 (N_592,In_1568,In_690);
xor U593 (N_593,In_1620,In_3601);
nor U594 (N_594,In_4819,In_4531);
or U595 (N_595,In_750,In_4745);
and U596 (N_596,In_4725,In_1153);
and U597 (N_597,In_4122,In_2490);
or U598 (N_598,In_1334,In_2729);
or U599 (N_599,In_3600,In_264);
and U600 (N_600,In_4668,In_4544);
nand U601 (N_601,In_3902,In_4693);
and U602 (N_602,In_833,In_4529);
and U603 (N_603,In_2313,In_630);
nand U604 (N_604,In_3465,In_1256);
xnor U605 (N_605,In_2467,In_3555);
xnor U606 (N_606,In_2946,In_2332);
nor U607 (N_607,In_208,In_1222);
or U608 (N_608,In_1586,In_3327);
xor U609 (N_609,In_1179,In_4844);
and U610 (N_610,In_1501,In_4049);
or U611 (N_611,In_991,In_4959);
or U612 (N_612,In_3469,In_1529);
or U613 (N_613,In_904,In_906);
or U614 (N_614,In_2163,In_428);
nand U615 (N_615,In_3806,In_864);
nor U616 (N_616,In_1229,In_3685);
or U617 (N_617,In_2602,In_4382);
or U618 (N_618,In_271,In_1381);
and U619 (N_619,In_4086,In_2944);
xor U620 (N_620,In_456,In_629);
and U621 (N_621,In_272,In_1263);
nand U622 (N_622,In_4594,In_714);
and U623 (N_623,In_182,In_25);
and U624 (N_624,In_1766,In_650);
and U625 (N_625,In_4815,In_2582);
nor U626 (N_626,In_2121,In_4875);
nand U627 (N_627,In_2146,In_2689);
nor U628 (N_628,In_2185,In_2477);
xor U629 (N_629,In_4223,In_795);
or U630 (N_630,In_424,In_2096);
and U631 (N_631,In_1281,In_4530);
or U632 (N_632,In_553,In_1802);
or U633 (N_633,In_2482,In_3270);
or U634 (N_634,In_1013,In_2879);
nand U635 (N_635,In_4244,In_2992);
nand U636 (N_636,In_4631,In_3868);
or U637 (N_637,In_2009,In_3874);
or U638 (N_638,In_3241,In_3858);
nand U639 (N_639,In_4618,In_4909);
nand U640 (N_640,In_4100,In_3547);
xor U641 (N_641,In_2744,In_4797);
xnor U642 (N_642,In_2321,In_1930);
nor U643 (N_643,In_1732,In_2686);
nor U644 (N_644,In_1083,In_3459);
and U645 (N_645,In_4459,In_3185);
nand U646 (N_646,In_4790,In_290);
xnor U647 (N_647,In_1663,In_2786);
nor U648 (N_648,In_3186,In_3374);
and U649 (N_649,In_779,In_909);
or U650 (N_650,In_3949,In_3671);
and U651 (N_651,In_2303,In_4401);
or U652 (N_652,In_4347,In_2540);
nor U653 (N_653,In_112,In_1494);
and U654 (N_654,In_2086,In_199);
xor U655 (N_655,In_1556,In_3338);
nor U656 (N_656,In_4497,In_1630);
and U657 (N_657,In_1718,In_4089);
or U658 (N_658,In_2347,In_4680);
xor U659 (N_659,In_3813,In_2342);
xnor U660 (N_660,In_4383,In_2198);
nand U661 (N_661,In_298,In_3882);
nand U662 (N_662,In_2737,In_247);
nor U663 (N_663,In_3460,In_4000);
nor U664 (N_664,In_3354,In_4836);
or U665 (N_665,In_1251,In_354);
xor U666 (N_666,In_1542,In_4241);
or U667 (N_667,In_1806,In_3305);
and U668 (N_668,In_150,In_896);
nor U669 (N_669,In_330,In_1642);
and U670 (N_670,In_429,In_3036);
or U671 (N_671,In_3852,In_2823);
and U672 (N_672,In_1016,In_1474);
nor U673 (N_673,In_3043,In_3735);
or U674 (N_674,In_3807,In_3427);
and U675 (N_675,In_1864,In_4532);
nor U676 (N_676,In_3533,In_1665);
nor U677 (N_677,In_1183,In_2950);
xor U678 (N_678,In_691,In_868);
or U679 (N_679,In_3001,In_3924);
xor U680 (N_680,In_3222,In_1725);
nor U681 (N_681,In_3711,In_141);
and U682 (N_682,In_2885,In_210);
nor U683 (N_683,In_198,In_2726);
and U684 (N_684,In_4325,In_2896);
xnor U685 (N_685,In_1085,In_1217);
nand U686 (N_686,In_2456,In_1231);
and U687 (N_687,In_900,In_1234);
xnor U688 (N_688,In_4354,In_523);
or U689 (N_689,In_1211,In_1040);
and U690 (N_690,In_3627,In_3097);
or U691 (N_691,In_1936,In_254);
and U692 (N_692,In_4615,In_441);
nand U693 (N_693,In_2698,In_4772);
nor U694 (N_694,In_2844,In_1460);
or U695 (N_695,In_4733,In_2948);
or U696 (N_696,In_2410,In_1535);
xor U697 (N_697,In_4570,In_42);
and U698 (N_698,In_4994,In_409);
or U699 (N_699,In_2299,In_4768);
nor U700 (N_700,In_2363,In_3814);
or U701 (N_701,In_958,In_3825);
and U702 (N_702,In_4279,In_3643);
or U703 (N_703,In_3692,In_2846);
and U704 (N_704,In_1825,In_1260);
nor U705 (N_705,In_1816,In_4711);
xnor U706 (N_706,In_931,In_3081);
nor U707 (N_707,In_1571,In_1347);
and U708 (N_708,In_4526,In_519);
nand U709 (N_709,In_757,In_3977);
nand U710 (N_710,In_4443,In_427);
nand U711 (N_711,In_3400,In_3509);
xnor U712 (N_712,In_3619,In_3719);
nand U713 (N_713,In_3280,In_2674);
and U714 (N_714,In_555,In_759);
or U715 (N_715,In_2575,In_325);
xnor U716 (N_716,In_847,In_2093);
or U717 (N_717,In_4181,In_1098);
or U718 (N_718,In_3577,In_4897);
xor U719 (N_719,In_2666,In_3175);
nor U720 (N_720,In_2298,In_1189);
nor U721 (N_721,In_705,In_791);
or U722 (N_722,In_3861,In_1636);
and U723 (N_723,In_965,In_3321);
nor U724 (N_724,In_3744,In_3569);
xor U725 (N_725,In_878,In_202);
or U726 (N_726,In_1076,In_3876);
nor U727 (N_727,In_4587,In_1833);
nor U728 (N_728,In_1778,In_3700);
nor U729 (N_729,In_3352,In_663);
nor U730 (N_730,In_2351,In_3444);
or U731 (N_731,In_1440,In_688);
nor U732 (N_732,In_3657,In_2118);
nand U733 (N_733,In_1969,In_4137);
nor U734 (N_734,In_4713,In_3260);
xnor U735 (N_735,In_3223,In_480);
or U736 (N_736,In_653,In_2069);
and U737 (N_737,In_1382,In_2935);
and U738 (N_738,In_4744,In_4660);
nand U739 (N_739,In_4057,In_537);
nor U740 (N_740,In_461,In_396);
nor U741 (N_741,In_1985,In_3490);
or U742 (N_742,In_61,In_3995);
nor U743 (N_743,In_1563,In_132);
nand U744 (N_744,In_800,In_2544);
nor U745 (N_745,In_3855,In_398);
or U746 (N_746,In_2416,In_1509);
nand U747 (N_747,In_1186,In_3730);
nor U748 (N_748,In_4367,In_4);
nor U749 (N_749,In_1396,In_933);
or U750 (N_750,In_4629,In_1321);
xor U751 (N_751,In_4662,In_3483);
or U752 (N_752,In_4922,In_4417);
xnor U753 (N_753,In_2977,In_3904);
or U754 (N_754,In_3964,In_3009);
nor U755 (N_755,In_3388,In_1515);
xor U756 (N_756,In_4866,In_2033);
or U757 (N_757,In_4824,In_1868);
or U758 (N_758,In_951,In_3419);
nand U759 (N_759,In_2962,In_4872);
and U760 (N_760,In_3319,In_4490);
and U761 (N_761,In_3623,In_3944);
nand U762 (N_762,In_1899,In_1130);
xnor U763 (N_763,In_1492,In_4019);
and U764 (N_764,In_1721,In_2237);
xor U765 (N_765,In_477,In_2398);
xor U766 (N_766,In_922,In_643);
and U767 (N_767,In_2568,In_3937);
or U768 (N_768,In_3268,In_104);
nand U769 (N_769,In_717,In_4593);
and U770 (N_770,In_2523,In_4042);
xor U771 (N_771,In_4002,In_1853);
nand U772 (N_772,In_2090,In_4343);
nor U773 (N_773,In_2818,In_1477);
xnor U774 (N_774,In_595,In_1742);
nand U775 (N_775,In_1156,In_1319);
nor U776 (N_776,In_4752,In_447);
nand U777 (N_777,In_4787,In_1463);
xnor U778 (N_778,In_287,In_4538);
nand U779 (N_779,In_2167,In_4418);
nand U780 (N_780,In_4194,In_2660);
nor U781 (N_781,In_4853,In_1419);
or U782 (N_782,In_3131,In_2841);
or U783 (N_783,In_2323,In_58);
nand U784 (N_784,In_4273,In_2794);
nand U785 (N_785,In_3360,In_3747);
or U786 (N_786,In_1237,In_1118);
xor U787 (N_787,In_2091,In_3900);
and U788 (N_788,In_4120,In_552);
or U789 (N_789,In_2893,In_4240);
nand U790 (N_790,In_2630,In_2337);
nand U791 (N_791,In_4512,In_3116);
nor U792 (N_792,In_2304,In_869);
xnor U793 (N_793,In_75,In_2888);
nor U794 (N_794,In_2570,In_4001);
xor U795 (N_795,In_4611,In_3782);
xnor U796 (N_796,In_2954,In_4357);
nor U797 (N_797,In_4868,In_3083);
nand U798 (N_798,In_2494,In_2063);
xnor U799 (N_799,In_3237,In_2335);
xor U800 (N_800,In_3899,In_4365);
nor U801 (N_801,In_3539,In_1342);
and U802 (N_802,In_1940,In_390);
xor U803 (N_803,In_2899,In_1951);
or U804 (N_804,In_4689,In_2843);
nor U805 (N_805,In_813,In_2262);
nand U806 (N_806,In_3541,In_3486);
nand U807 (N_807,In_3891,In_2557);
nand U808 (N_808,In_2251,In_4831);
nor U809 (N_809,In_1159,In_159);
or U810 (N_810,In_4812,In_1430);
or U811 (N_811,In_1077,In_3591);
or U812 (N_812,In_770,In_3117);
and U813 (N_813,In_3466,In_4915);
nand U814 (N_814,In_4926,In_2233);
nand U815 (N_815,In_2152,In_3707);
or U816 (N_816,In_768,In_3917);
nor U817 (N_817,In_1412,In_357);
nor U818 (N_818,In_4975,In_4896);
nor U819 (N_819,In_3972,In_754);
nor U820 (N_820,In_875,In_1562);
or U821 (N_821,In_3895,In_3229);
or U822 (N_822,In_2370,In_120);
and U823 (N_823,In_2651,In_155);
and U824 (N_824,In_4407,In_1160);
nor U825 (N_825,In_2453,In_1939);
or U826 (N_826,In_366,In_3761);
nor U827 (N_827,In_660,In_2736);
nand U828 (N_828,In_633,In_2338);
nand U829 (N_829,In_3072,In_2124);
nor U830 (N_830,In_1426,In_444);
or U831 (N_831,In_4676,In_1854);
nand U832 (N_832,In_2994,In_3228);
or U833 (N_833,In_1023,In_3918);
or U834 (N_834,In_1932,In_1398);
and U835 (N_835,In_3375,In_1927);
xor U836 (N_836,In_2519,In_2150);
or U837 (N_837,In_463,In_2076);
xnor U838 (N_838,In_2228,In_873);
xnor U839 (N_839,In_1086,In_2719);
nand U840 (N_840,In_4715,In_701);
nand U841 (N_841,In_3059,In_4048);
xnor U842 (N_842,In_2513,In_3302);
xnor U843 (N_843,In_3146,In_4509);
nor U844 (N_844,In_4535,In_2319);
and U845 (N_845,In_3598,In_3499);
nor U846 (N_846,In_1152,In_4682);
nor U847 (N_847,In_4395,In_2783);
and U848 (N_848,In_11,In_255);
or U849 (N_849,In_626,In_3540);
xor U850 (N_850,In_2538,In_3833);
or U851 (N_851,In_2534,In_1294);
xor U852 (N_852,In_4427,In_1312);
and U853 (N_853,In_2765,In_1545);
and U854 (N_854,In_2810,In_2531);
or U855 (N_855,In_3652,In_4132);
nor U856 (N_856,In_738,In_3205);
and U857 (N_857,In_2866,In_2532);
nand U858 (N_858,In_854,In_1684);
nor U859 (N_859,In_744,In_4518);
nor U860 (N_860,In_4252,In_2825);
nor U861 (N_861,In_2514,In_1433);
xnor U862 (N_862,In_899,In_1676);
xnor U863 (N_863,In_4890,In_1769);
xnor U864 (N_864,In_2480,In_2789);
nor U865 (N_865,In_1018,In_2205);
xor U866 (N_866,In_2779,In_4652);
nand U867 (N_867,In_2608,In_4077);
nand U868 (N_868,In_2877,In_2700);
or U869 (N_869,In_445,In_1647);
xor U870 (N_870,In_4879,In_4666);
nand U871 (N_871,In_360,In_2053);
or U872 (N_872,In_1573,In_3580);
or U873 (N_873,In_3023,In_3463);
or U874 (N_874,In_406,In_4857);
and U875 (N_875,In_2606,In_1700);
nor U876 (N_876,In_4923,In_941);
or U877 (N_877,In_529,In_4981);
and U878 (N_878,In_2555,In_4368);
xnor U879 (N_879,In_496,In_2391);
or U880 (N_880,In_1090,In_3610);
xnor U881 (N_881,In_614,In_2092);
nand U882 (N_882,In_814,In_3638);
nor U883 (N_883,In_4426,In_2894);
and U884 (N_884,In_3526,In_707);
nor U885 (N_885,In_3614,In_4450);
or U886 (N_886,In_4889,In_3837);
xor U887 (N_887,In_4763,In_4505);
or U888 (N_888,In_4776,In_3471);
or U889 (N_889,In_820,In_4270);
nor U890 (N_890,In_3956,In_1417);
and U891 (N_891,In_3632,In_2803);
nor U892 (N_892,In_752,In_2165);
or U893 (N_893,In_2835,In_1350);
nand U894 (N_894,In_1128,In_4648);
and U895 (N_895,In_1954,In_3501);
or U896 (N_896,In_4066,In_490);
nand U897 (N_897,In_3041,In_4639);
or U898 (N_898,In_3474,In_1287);
or U899 (N_899,In_589,In_1964);
nor U900 (N_900,In_3159,In_3839);
nor U901 (N_901,In_1437,In_3076);
and U902 (N_902,In_1057,In_1680);
or U903 (N_903,In_4336,In_2267);
and U904 (N_904,In_3789,In_3055);
or U905 (N_905,In_4287,In_2966);
nor U906 (N_906,In_1228,In_375);
nor U907 (N_907,In_4031,In_2334);
or U908 (N_908,In_3045,In_3560);
and U909 (N_909,In_2815,In_1454);
nand U910 (N_910,In_3594,In_892);
and U911 (N_911,In_3725,In_1675);
or U912 (N_912,In_2305,In_2388);
nand U913 (N_913,In_20,In_3698);
xnor U914 (N_914,In_4175,In_4949);
nor U915 (N_915,In_4792,In_2836);
or U916 (N_916,In_2854,In_3416);
and U917 (N_917,In_1313,In_2629);
or U918 (N_918,In_2306,In_1652);
nand U919 (N_919,In_446,In_219);
or U920 (N_920,In_835,In_4672);
or U921 (N_921,In_2042,In_684);
nand U922 (N_922,In_2580,In_1774);
nor U923 (N_923,In_4508,In_3505);
or U924 (N_924,In_4552,In_4727);
or U925 (N_925,In_2119,In_2614);
nor U926 (N_926,In_2430,In_2486);
and U927 (N_927,In_1897,In_1154);
and U928 (N_928,In_3082,In_2943);
nor U929 (N_929,In_1752,In_459);
xnor U930 (N_930,In_2207,In_4834);
and U931 (N_931,In_1604,In_3768);
xor U932 (N_932,In_3218,In_615);
xor U933 (N_933,In_1227,In_294);
xnor U934 (N_934,In_616,In_720);
nand U935 (N_935,In_4659,In_952);
nand U936 (N_936,In_2290,In_3818);
and U937 (N_937,In_3575,In_3981);
and U938 (N_938,In_1919,In_1056);
nand U939 (N_939,In_1795,In_3312);
and U940 (N_940,In_2360,In_934);
or U941 (N_941,In_3854,In_652);
or U942 (N_942,In_2278,In_3843);
nand U943 (N_943,In_3411,In_3187);
and U944 (N_944,In_1002,In_2239);
nand U945 (N_945,In_1674,In_2040);
and U946 (N_946,In_530,In_2522);
nand U947 (N_947,In_913,In_78);
xor U948 (N_948,In_4404,In_4814);
and U949 (N_949,In_4454,In_2407);
or U950 (N_950,In_2068,In_1750);
or U951 (N_951,In_391,In_4561);
and U952 (N_952,In_501,In_881);
xnor U953 (N_953,In_56,In_1796);
or U954 (N_954,In_3073,In_2990);
and U955 (N_955,In_4786,In_1901);
nand U956 (N_956,In_2988,In_1362);
nand U957 (N_957,In_3295,In_3609);
or U958 (N_958,In_4771,In_4259);
xnor U959 (N_959,In_1480,In_670);
xor U960 (N_960,In_755,In_4242);
and U961 (N_961,In_1301,In_4276);
xor U962 (N_962,In_3670,In_1650);
nand U963 (N_963,In_2880,In_1060);
xnor U964 (N_964,In_4795,In_2517);
or U965 (N_965,In_3844,In_2937);
or U966 (N_966,In_4176,In_3532);
and U967 (N_967,In_679,In_2723);
xnor U968 (N_968,In_96,In_727);
nand U969 (N_969,In_1979,In_3990);
or U970 (N_970,In_1079,In_1314);
nand U971 (N_971,In_1413,In_1708);
nor U972 (N_972,In_4883,In_3785);
nor U973 (N_973,In_4542,In_4206);
nand U974 (N_974,In_3683,In_2358);
or U975 (N_975,In_2795,In_2924);
nand U976 (N_976,In_1633,In_3507);
nand U977 (N_977,In_130,In_2697);
nor U978 (N_978,In_3212,In_715);
nand U979 (N_979,In_2362,In_1521);
nor U980 (N_980,In_3929,In_983);
or U981 (N_981,In_3233,In_3962);
or U982 (N_982,In_2019,In_295);
xor U983 (N_983,In_1918,In_1760);
or U984 (N_984,In_1432,In_2138);
or U985 (N_985,In_101,In_4322);
or U986 (N_986,In_13,In_1025);
nor U987 (N_987,In_914,In_1696);
or U988 (N_988,In_961,In_4375);
xor U989 (N_989,In_4020,In_2383);
and U990 (N_990,In_1065,In_285);
and U991 (N_991,In_498,In_3128);
or U992 (N_992,In_3717,In_635);
xnor U993 (N_993,In_2126,In_510);
and U994 (N_994,In_4439,In_2623);
xor U995 (N_995,In_2638,In_106);
xor U996 (N_996,In_1855,In_203);
xor U997 (N_997,In_2161,In_2348);
and U998 (N_998,In_4084,In_235);
nand U999 (N_999,In_3596,In_4481);
xnor U1000 (N_1000,In_2038,In_2763);
nor U1001 (N_1001,In_772,In_977);
and U1002 (N_1002,In_2314,In_3920);
nand U1003 (N_1003,In_316,In_4608);
or U1004 (N_1004,In_2276,In_3456);
nand U1005 (N_1005,In_3226,In_1400);
nor U1006 (N_1006,In_4523,In_4886);
xnor U1007 (N_1007,In_3637,In_923);
and U1008 (N_1008,In_1686,In_939);
nor U1009 (N_1009,In_3510,In_3166);
xnor U1010 (N_1010,In_2141,In_747);
or U1011 (N_1011,In_1582,In_2350);
nor U1012 (N_1012,In_3395,In_2639);
nand U1013 (N_1013,In_2413,In_173);
or U1014 (N_1014,In_741,In_3811);
nor U1015 (N_1015,In_2432,In_3326);
and U1016 (N_1016,In_257,In_4160);
xnor U1017 (N_1017,In_1896,In_218);
nand U1018 (N_1018,In_602,In_4770);
nor U1019 (N_1019,In_989,In_1024);
or U1020 (N_1020,In_1575,In_4575);
or U1021 (N_1021,In_1010,In_4363);
xor U1022 (N_1022,In_4182,In_2300);
and U1023 (N_1023,In_3853,In_4964);
nand U1024 (N_1024,In_593,In_1787);
and U1025 (N_1025,In_3597,In_32);
nor U1026 (N_1026,In_4256,In_385);
nand U1027 (N_1027,In_1539,In_492);
and U1028 (N_1028,In_3898,In_4609);
and U1029 (N_1029,In_4746,In_4723);
nand U1030 (N_1030,In_3290,In_3763);
and U1031 (N_1031,In_2858,In_2609);
xor U1032 (N_1032,In_1997,In_2574);
nand U1033 (N_1033,In_309,In_4574);
nand U1034 (N_1034,In_3880,In_3945);
and U1035 (N_1035,In_1788,In_2680);
xor U1036 (N_1036,In_763,In_2203);
or U1037 (N_1037,In_4612,In_4250);
nor U1038 (N_1038,In_3611,In_2292);
or U1039 (N_1039,In_568,In_945);
nor U1040 (N_1040,In_54,In_2535);
xor U1041 (N_1041,In_572,In_4690);
nand U1042 (N_1042,In_3372,In_4740);
or U1043 (N_1043,In_2423,In_3475);
or U1044 (N_1044,In_2978,In_3239);
or U1045 (N_1045,In_819,In_697);
nor U1046 (N_1046,In_3458,In_4557);
nand U1047 (N_1047,In_2114,In_4314);
or U1048 (N_1048,In_4751,In_414);
and U1049 (N_1049,In_1906,In_4856);
nor U1050 (N_1050,In_565,In_4386);
nand U1051 (N_1051,In_2242,In_4480);
nor U1052 (N_1052,In_1916,In_2654);
nor U1053 (N_1053,In_3448,In_1366);
and U1054 (N_1054,In_2039,In_1672);
and U1055 (N_1055,In_4419,In_279);
xnor U1056 (N_1056,In_471,In_4333);
nor U1057 (N_1057,In_3699,In_2394);
nand U1058 (N_1058,In_4431,In_870);
and U1059 (N_1059,In_1332,In_3993);
nand U1060 (N_1060,In_4078,In_1296);
or U1061 (N_1061,In_803,In_576);
nand U1062 (N_1062,In_1322,In_3245);
xnor U1063 (N_1063,In_2627,In_2466);
or U1064 (N_1064,In_1557,In_246);
nor U1065 (N_1065,In_3836,In_2346);
nand U1066 (N_1066,In_3544,In_3359);
nor U1067 (N_1067,In_1990,In_3587);
or U1068 (N_1068,In_1377,In_778);
nand U1069 (N_1069,In_144,In_4105);
xor U1070 (N_1070,In_3109,In_1485);
and U1071 (N_1071,In_3752,In_1317);
nor U1072 (N_1072,In_4189,In_4755);
or U1073 (N_1073,In_4438,In_2722);
nor U1074 (N_1074,In_4849,In_394);
or U1075 (N_1075,In_3650,In_3859);
xnor U1076 (N_1076,In_2485,In_3172);
or U1077 (N_1077,In_600,In_2718);
xnor U1078 (N_1078,In_3646,In_4578);
and U1079 (N_1079,In_3679,In_2890);
nor U1080 (N_1080,In_558,In_4567);
nor U1081 (N_1081,In_3841,In_2390);
nand U1082 (N_1082,In_804,In_816);
nor U1083 (N_1083,In_2703,In_3171);
nand U1084 (N_1084,In_4208,In_2622);
nand U1085 (N_1085,In_764,In_1662);
xnor U1086 (N_1086,In_489,In_1009);
nor U1087 (N_1087,In_1911,In_625);
or U1088 (N_1088,In_4373,In_3062);
or U1089 (N_1089,In_2230,In_426);
xnor U1090 (N_1090,In_3764,In_1999);
or U1091 (N_1091,In_307,In_4484);
and U1092 (N_1092,In_733,In_8);
nor U1093 (N_1093,In_1629,In_648);
xnor U1094 (N_1094,In_2865,In_1707);
xor U1095 (N_1095,In_2218,In_3350);
xor U1096 (N_1096,In_1653,In_3018);
nor U1097 (N_1097,In_4924,In_2008);
xor U1098 (N_1098,In_1740,In_3137);
and U1099 (N_1099,In_987,In_4296);
and U1100 (N_1100,In_1184,In_2011);
nand U1101 (N_1101,In_320,In_1592);
or U1102 (N_1102,In_885,In_2234);
nand U1103 (N_1103,In_4318,In_2160);
nand U1104 (N_1104,In_526,In_3894);
nand U1105 (N_1105,In_4035,In_4510);
xor U1106 (N_1106,In_908,In_3173);
nand U1107 (N_1107,In_4521,In_2311);
nor U1108 (N_1108,In_3727,In_52);
nand U1109 (N_1109,In_2017,In_3570);
and U1110 (N_1110,In_258,In_3152);
and U1111 (N_1111,In_3316,In_2957);
or U1112 (N_1112,In_2258,In_2199);
or U1113 (N_1113,In_4904,In_280);
xnor U1114 (N_1114,In_2341,In_1570);
nand U1115 (N_1115,In_1453,In_186);
xnor U1116 (N_1116,In_1113,In_3498);
xnor U1117 (N_1117,In_1522,In_3054);
or U1118 (N_1118,In_4180,In_2871);
nand U1119 (N_1119,In_1869,In_2007);
or U1120 (N_1120,In_709,In_3513);
nand U1121 (N_1121,In_299,In_1884);
and U1122 (N_1122,In_1977,In_877);
nand U1123 (N_1123,In_3314,In_187);
and U1124 (N_1124,In_4323,In_1715);
xnor U1125 (N_1125,In_3142,In_4097);
nor U1126 (N_1126,In_730,In_3613);
nor U1127 (N_1127,In_1749,In_2154);
or U1128 (N_1128,In_767,In_2500);
xnor U1129 (N_1129,In_1963,In_588);
or U1130 (N_1130,In_3840,In_895);
or U1131 (N_1131,In_879,In_4110);
nand U1132 (N_1132,In_3133,In_2928);
nor U1133 (N_1133,In_3621,In_2463);
or U1134 (N_1134,In_3034,In_2281);
and U1135 (N_1135,In_3968,In_1391);
nand U1136 (N_1136,In_1326,In_3769);
nor U1137 (N_1137,In_4854,In_1805);
or U1138 (N_1138,In_2800,In_4320);
or U1139 (N_1139,In_3829,In_140);
nor U1140 (N_1140,In_1673,In_1014);
and U1141 (N_1141,In_1397,In_4601);
nand U1142 (N_1142,In_1514,In_3252);
nor U1143 (N_1143,In_3379,In_692);
nand U1144 (N_1144,In_2864,In_4806);
xnor U1145 (N_1145,In_1800,In_4372);
nand U1146 (N_1146,In_2895,In_1092);
and U1147 (N_1147,In_2254,In_4957);
or U1148 (N_1148,In_3303,In_1681);
xnor U1149 (N_1149,In_1271,In_204);
nor U1150 (N_1150,In_2066,In_4258);
nor U1151 (N_1151,In_3078,In_3386);
and U1152 (N_1152,In_2378,In_3584);
and U1153 (N_1153,In_3380,In_66);
xor U1154 (N_1154,In_545,In_4585);
or U1155 (N_1155,In_1401,In_1841);
xnor U1156 (N_1156,In_3485,In_3141);
nand U1157 (N_1157,In_3629,In_2669);
xor U1158 (N_1158,In_4597,In_3203);
or U1159 (N_1159,In_3702,In_966);
and U1160 (N_1160,In_2285,In_1103);
nor U1161 (N_1161,In_3068,In_1945);
or U1162 (N_1162,In_4272,In_1757);
nor U1163 (N_1163,In_3382,In_2183);
nor U1164 (N_1164,In_1409,In_3940);
or U1165 (N_1165,In_1006,In_2860);
xnor U1166 (N_1166,In_532,In_1404);
nor U1167 (N_1167,In_469,In_2442);
nor U1168 (N_1168,In_2461,In_1157);
xnor U1169 (N_1169,In_4010,In_3760);
and U1170 (N_1170,In_4541,In_1578);
nand U1171 (N_1171,In_2856,In_2904);
xnor U1172 (N_1172,In_1383,In_2065);
and U1173 (N_1173,In_1900,In_3543);
or U1174 (N_1174,In_1845,In_2405);
xnor U1175 (N_1175,In_1645,In_1768);
xor U1176 (N_1176,In_143,In_1814);
xor U1177 (N_1177,In_2472,In_1502);
xnor U1178 (N_1178,In_574,In_2330);
and U1179 (N_1179,In_4592,In_988);
or U1180 (N_1180,In_3442,In_267);
and U1181 (N_1181,In_3430,In_4925);
nor U1182 (N_1182,In_2054,In_2084);
or U1183 (N_1183,In_4154,In_1719);
and U1184 (N_1184,In_3518,In_2861);
or U1185 (N_1185,In_2693,In_546);
nand U1186 (N_1186,In_4633,In_4440);
nand U1187 (N_1187,In_1764,In_2400);
and U1188 (N_1188,In_773,In_3562);
nor U1189 (N_1189,In_3243,In_2170);
nor U1190 (N_1190,In_4229,In_3850);
xnor U1191 (N_1191,In_3748,In_4900);
nor U1192 (N_1192,In_107,In_364);
nor U1193 (N_1193,In_2384,In_1093);
xnor U1194 (N_1194,In_4489,In_2664);
and U1195 (N_1195,In_2470,In_372);
and U1196 (N_1196,In_2248,In_3235);
or U1197 (N_1197,In_4696,In_2951);
nand U1198 (N_1198,In_4793,In_4298);
nand U1199 (N_1199,In_2473,In_2993);
or U1200 (N_1200,In_3493,In_2002);
nor U1201 (N_1201,In_3877,In_4188);
and U1202 (N_1202,In_3209,In_465);
xor U1203 (N_1203,In_4669,In_4146);
and U1204 (N_1204,In_4482,In_1880);
or U1205 (N_1205,In_237,In_4762);
nor U1206 (N_1206,In_4249,In_4046);
nor U1207 (N_1207,In_1780,In_1363);
and U1208 (N_1208,In_2312,In_3119);
xnor U1209 (N_1209,In_3590,In_3425);
nand U1210 (N_1210,In_3871,In_921);
xnor U1211 (N_1211,In_4053,In_1253);
or U1212 (N_1212,In_4576,In_1105);
xnor U1213 (N_1213,In_165,In_4337);
xor U1214 (N_1214,In_2062,In_4898);
nand U1215 (N_1215,In_4560,In_3358);
xor U1216 (N_1216,In_4704,In_4550);
nor U1217 (N_1217,In_4555,In_476);
and U1218 (N_1218,In_2503,In_2569);
nand U1219 (N_1219,In_998,In_3599);
nand U1220 (N_1220,In_587,In_97);
and U1221 (N_1221,In_2788,In_536);
and U1222 (N_1222,In_3101,In_4705);
nor U1223 (N_1223,In_3421,In_2266);
nor U1224 (N_1224,In_2601,In_2556);
nand U1225 (N_1225,In_3578,In_1967);
nor U1226 (N_1226,In_3928,In_1288);
nand U1227 (N_1227,In_1360,In_597);
nand U1228 (N_1228,In_4070,In_3234);
or U1229 (N_1229,In_4364,In_3766);
or U1230 (N_1230,In_2874,In_4112);
and U1231 (N_1231,In_4351,In_1691);
or U1232 (N_1232,In_2761,In_1837);
or U1233 (N_1233,In_2356,In_3875);
nand U1234 (N_1234,In_3378,In_849);
nand U1235 (N_1235,In_4269,In_1427);
xnor U1236 (N_1236,In_170,In_1942);
nand U1237 (N_1237,In_288,In_860);
xnor U1238 (N_1238,In_2502,In_2536);
nand U1239 (N_1239,In_694,In_3111);
nor U1240 (N_1240,In_1266,In_4860);
xor U1241 (N_1241,In_3834,In_3932);
nand U1242 (N_1242,In_2187,In_2392);
and U1243 (N_1243,In_26,In_2938);
or U1244 (N_1244,In_1628,In_3751);
and U1245 (N_1245,In_3635,In_3461);
or U1246 (N_1246,In_711,In_862);
xor U1247 (N_1247,In_4353,In_3020);
and U1248 (N_1248,In_2581,In_1839);
nand U1249 (N_1249,In_3701,In_3343);
nor U1250 (N_1250,In_2169,In_146);
or U1251 (N_1251,In_3821,In_2576);
xor U1252 (N_1252,In_4183,In_2817);
or U1253 (N_1253,In_4062,In_3158);
nand U1254 (N_1254,In_2565,In_704);
and U1255 (N_1255,In_3308,In_2439);
nor U1256 (N_1256,In_293,In_4673);
nand U1257 (N_1257,In_2286,In_4217);
nand U1258 (N_1258,In_3202,In_350);
xor U1259 (N_1259,In_4384,In_1210);
xor U1260 (N_1260,In_4295,In_1390);
nor U1261 (N_1261,In_1102,In_1820);
nand U1262 (N_1262,In_322,In_2308);
nand U1263 (N_1263,In_1835,In_4345);
nand U1264 (N_1264,In_4980,In_3640);
nor U1265 (N_1265,In_1235,In_1150);
nand U1266 (N_1266,In_4081,In_84);
nor U1267 (N_1267,In_4758,In_4147);
or U1268 (N_1268,In_3363,In_2307);
and U1269 (N_1269,In_3102,In_1299);
and U1270 (N_1270,In_4064,In_3696);
or U1271 (N_1271,In_160,In_1094);
xor U1272 (N_1272,In_3678,In_4671);
nor U1273 (N_1273,In_4707,In_2553);
nor U1274 (N_1274,In_3484,In_2881);
xnor U1275 (N_1275,In_2462,In_4501);
xor U1276 (N_1276,In_3695,In_1272);
or U1277 (N_1277,In_984,In_4334);
nor U1278 (N_1278,In_4186,In_4494);
xnor U1279 (N_1279,In_610,In_1689);
nor U1280 (N_1280,In_2837,In_3819);
nand U1281 (N_1281,In_4679,In_2175);
or U1282 (N_1282,In_3901,In_2296);
or U1283 (N_1283,In_4516,In_3340);
and U1284 (N_1284,In_1478,In_2941);
xor U1285 (N_1285,In_3301,In_3495);
nor U1286 (N_1286,In_4220,In_2798);
nor U1287 (N_1287,In_88,In_315);
or U1288 (N_1288,In_1490,In_666);
xor U1289 (N_1289,In_3477,In_19);
nand U1290 (N_1290,In_4377,In_1225);
or U1291 (N_1291,In_80,In_3946);
nand U1292 (N_1292,In_3106,In_21);
xor U1293 (N_1293,In_2188,In_2526);
and U1294 (N_1294,In_4356,In_1935);
or U1295 (N_1295,In_1506,In_938);
nor U1296 (N_1296,In_355,In_3516);
or U1297 (N_1297,In_3749,In_3069);
xor U1298 (N_1298,In_421,In_910);
nor U1299 (N_1299,In_3467,In_4114);
or U1300 (N_1300,In_1207,In_786);
nor U1301 (N_1301,In_145,In_1727);
nand U1302 (N_1302,In_3080,In_2468);
nand U1303 (N_1303,In_1865,In_4978);
and U1304 (N_1304,In_243,In_762);
xor U1305 (N_1305,In_2210,In_2489);
or U1306 (N_1306,In_278,In_2915);
nor U1307 (N_1307,In_3121,In_3276);
xnor U1308 (N_1308,In_4195,In_4870);
or U1309 (N_1309,In_4350,In_3489);
or U1310 (N_1310,In_1753,In_4717);
and U1311 (N_1311,In_4749,In_2227);
and U1312 (N_1312,In_2246,In_4396);
nand U1313 (N_1313,In_1019,In_1265);
nor U1314 (N_1314,In_1187,In_3548);
nand U1315 (N_1315,In_1297,In_4332);
or U1316 (N_1316,In_918,In_1465);
or U1317 (N_1317,In_499,In_399);
nor U1318 (N_1318,In_2046,In_185);
and U1319 (N_1319,In_256,In_2056);
xnor U1320 (N_1320,In_4436,In_979);
or U1321 (N_1321,In_940,In_612);
nor U1322 (N_1322,In_2780,In_486);
nand U1323 (N_1323,In_4761,In_3178);
and U1324 (N_1324,In_2931,In_4692);
nor U1325 (N_1325,In_4474,In_1425);
nand U1326 (N_1326,In_4961,In_1469);
and U1327 (N_1327,In_2200,In_4388);
nor U1328 (N_1328,In_2959,In_2982);
nor U1329 (N_1329,In_344,In_3124);
xor U1330 (N_1330,In_4729,In_3473);
xor U1331 (N_1331,In_1070,In_592);
nor U1332 (N_1332,In_866,In_363);
and U1333 (N_1333,In_1175,In_4425);
or U1334 (N_1334,In_3263,In_2914);
and U1335 (N_1335,In_333,In_3309);
and U1336 (N_1336,In_3957,In_946);
nor U1337 (N_1337,In_2428,In_4569);
and U1338 (N_1338,In_3324,In_2804);
or U1339 (N_1339,In_2701,In_3688);
and U1340 (N_1340,In_4080,In_3005);
or U1341 (N_1341,In_2749,In_3457);
and U1342 (N_1342,In_2912,In_3230);
nand U1343 (N_1343,In_4977,In_1572);
and U1344 (N_1344,In_2752,In_4236);
nand U1345 (N_1345,In_2172,In_1974);
nand U1346 (N_1346,In_3922,In_3376);
xnor U1347 (N_1347,In_2474,In_668);
and U1348 (N_1348,In_2471,In_3012);
nor U1349 (N_1349,In_4955,In_2074);
or U1350 (N_1350,In_3714,In_4969);
nand U1351 (N_1351,In_2424,In_1720);
nor U1352 (N_1352,In_1912,In_3293);
xor U1353 (N_1353,In_2481,In_4808);
xor U1354 (N_1354,In_2548,In_1537);
or U1355 (N_1355,In_2562,In_1751);
xor U1356 (N_1356,In_3887,In_4448);
nand U1357 (N_1357,In_2873,In_2640);
xor U1358 (N_1358,In_4619,In_1443);
or U1359 (N_1359,In_3195,In_4623);
or U1360 (N_1360,In_3721,In_671);
nor U1361 (N_1361,In_2434,In_1931);
and U1362 (N_1362,In_2643,In_4644);
nor U1363 (N_1363,In_3921,In_2317);
and U1364 (N_1364,In_716,In_964);
and U1365 (N_1365,In_3476,In_2908);
and U1366 (N_1366,In_1772,In_2103);
or U1367 (N_1367,In_4622,In_2848);
or U1368 (N_1368,In_3847,In_1370);
nand U1369 (N_1369,In_2784,In_2657);
or U1370 (N_1370,In_3762,In_1277);
nand U1371 (N_1371,In_4231,In_4421);
and U1372 (N_1372,In_1221,In_1667);
and U1373 (N_1373,In_539,In_3893);
or U1374 (N_1374,In_4963,In_1134);
xnor U1375 (N_1375,In_3144,In_1236);
nand U1376 (N_1376,In_2379,In_889);
and U1377 (N_1377,In_111,In_69);
nor U1378 (N_1378,In_224,In_831);
nand U1379 (N_1379,In_2484,In_2821);
and U1380 (N_1380,In_177,In_4290);
nor U1381 (N_1381,In_3681,In_4912);
or U1382 (N_1382,In_1928,In_706);
nand U1383 (N_1383,In_4677,In_2940);
nor U1384 (N_1384,In_1588,In_1632);
nand U1385 (N_1385,In_3390,In_4234);
xor U1386 (N_1386,In_3729,In_3565);
or U1387 (N_1387,In_3971,In_72);
or U1388 (N_1388,In_2099,In_4764);
and U1389 (N_1389,In_4214,In_2357);
xnor U1390 (N_1390,In_4553,In_3053);
and U1391 (N_1391,In_4145,In_2812);
nor U1392 (N_1392,In_3192,In_4522);
or U1393 (N_1393,In_4476,In_2128);
nand U1394 (N_1394,In_1411,In_1205);
and U1395 (N_1395,In_1257,In_3035);
and U1396 (N_1396,In_442,In_973);
xor U1397 (N_1397,In_1881,In_4144);
or U1398 (N_1398,In_1828,In_1600);
and U1399 (N_1399,In_2293,In_4944);
xor U1400 (N_1400,In_4061,In_886);
or U1401 (N_1401,In_2711,In_4130);
xor U1402 (N_1402,In_253,In_2260);
and U1403 (N_1403,In_2171,In_3517);
nor U1404 (N_1404,In_1878,In_808);
or U1405 (N_1405,In_1937,In_1671);
and U1406 (N_1406,In_4187,In_3780);
and U1407 (N_1407,In_3071,In_1597);
or U1408 (N_1408,In_4307,In_4286);
nand U1409 (N_1409,In_1822,In_1181);
and U1410 (N_1410,In_1616,In_4936);
and U1411 (N_1411,In_2110,In_1464);
xor U1412 (N_1412,In_3056,In_3753);
nor U1413 (N_1413,In_212,In_2530);
or U1414 (N_1414,In_677,In_49);
and U1415 (N_1415,In_3846,In_4281);
nor U1416 (N_1416,In_3622,In_3439);
or U1417 (N_1417,In_2464,In_4779);
and U1418 (N_1418,In_1135,In_517);
or U1419 (N_1419,In_2684,In_3225);
or U1420 (N_1420,In_3088,In_274);
and U1421 (N_1421,In_1735,In_4099);
xnor U1422 (N_1422,In_848,In_3890);
xnor U1423 (N_1423,In_4257,In_464);
nand U1424 (N_1424,In_4164,In_3407);
and U1425 (N_1425,In_3127,In_4756);
xnor U1426 (N_1426,In_2026,In_4948);
nand U1427 (N_1427,In_3399,In_3438);
nand U1428 (N_1428,In_3155,In_1950);
nand U1429 (N_1429,In_3014,In_4759);
or U1430 (N_1430,In_2628,In_1);
nand U1431 (N_1431,In_591,In_1339);
and U1432 (N_1432,In_722,In_570);
or U1433 (N_1433,In_685,In_2707);
nor U1434 (N_1434,In_4434,In_1001);
and U1435 (N_1435,In_1232,In_3207);
nor U1436 (N_1436,In_2694,In_852);
nor U1437 (N_1437,In_845,In_205);
nor U1438 (N_1438,In_2833,In_3086);
or U1439 (N_1439,In_3108,In_1943);
or U1440 (N_1440,In_2353,In_1902);
nand U1441 (N_1441,In_1042,In_1758);
and U1442 (N_1442,In_3651,In_3983);
xnor U1443 (N_1443,In_2072,In_3689);
and U1444 (N_1444,In_4995,In_3915);
or U1445 (N_1445,In_4796,In_2932);
nand U1446 (N_1446,In_1238,In_3047);
or U1447 (N_1447,In_4039,In_3177);
or U1448 (N_1448,In_3094,In_4023);
and U1449 (N_1449,In_2758,In_3169);
xor U1450 (N_1450,In_4989,In_4954);
and U1451 (N_1451,In_1722,In_200);
xor U1452 (N_1452,In_2354,In_4701);
nand U1453 (N_1453,In_509,In_2241);
and U1454 (N_1454,In_1978,In_346);
xor U1455 (N_1455,In_2329,In_1748);
nor U1456 (N_1456,In_2713,In_1762);
nor U1457 (N_1457,In_1871,In_1846);
xnor U1458 (N_1458,In_3716,In_1770);
xnor U1459 (N_1459,In_2597,In_2559);
nor U1460 (N_1460,In_502,In_3008);
and U1461 (N_1461,In_2615,In_2374);
nand U1462 (N_1462,In_3310,In_4533);
or U1463 (N_1463,In_335,In_2238);
and U1464 (N_1464,In_3265,In_123);
nor U1465 (N_1465,In_4346,In_4869);
xnor U1466 (N_1466,In_4201,In_1765);
xnor U1467 (N_1467,In_4331,In_4650);
xnor U1468 (N_1468,In_4468,In_1126);
xnor U1469 (N_1469,In_2583,In_3183);
nand U1470 (N_1470,In_1462,In_2315);
xor U1471 (N_1471,In_948,In_2605);
nand U1472 (N_1472,In_4101,In_1338);
or U1473 (N_1473,In_1471,In_4193);
or U1474 (N_1474,In_4414,In_1962);
nor U1475 (N_1475,In_139,In_4694);
or U1476 (N_1476,In_3423,In_2123);
nor U1477 (N_1477,In_3973,In_1640);
xnor U1478 (N_1478,In_865,In_857);
and U1479 (N_1479,In_3464,In_134);
and U1480 (N_1480,In_3827,In_2676);
nor U1481 (N_1481,In_3927,In_2231);
or U1482 (N_1482,In_721,In_2742);
nand U1483 (N_1483,In_3860,In_2807);
xnor U1484 (N_1484,In_3573,In_1966);
and U1485 (N_1485,In_453,In_4968);
nand U1486 (N_1486,In_4032,In_3115);
nand U1487 (N_1487,In_4341,In_2647);
nand U1488 (N_1488,In_3404,In_628);
and U1489 (N_1489,In_2476,In_2318);
nor U1490 (N_1490,In_3451,In_4545);
nand U1491 (N_1491,In_178,In_1066);
nor U1492 (N_1492,In_220,In_1984);
nor U1493 (N_1493,In_3639,In_2933);
xor U1494 (N_1494,In_2018,In_2633);
or U1495 (N_1495,In_4513,In_1305);
xnor U1496 (N_1496,In_92,In_753);
and U1497 (N_1497,In_3522,In_531);
nor U1498 (N_1498,In_4962,In_2772);
and U1499 (N_1499,In_3285,In_1055);
and U1500 (N_1500,In_3318,In_481);
xnor U1501 (N_1501,In_1784,In_3961);
or U1502 (N_1502,In_2077,In_1944);
or U1503 (N_1503,In_4865,In_189);
nor U1504 (N_1504,In_1843,In_1108);
or U1505 (N_1505,In_4785,In_2487);
nand U1506 (N_1506,In_378,In_1244);
or U1507 (N_1507,In_2452,In_2999);
xnor U1508 (N_1508,In_667,In_2863);
nor U1509 (N_1509,In_4215,In_1550);
nor U1510 (N_1510,In_1410,In_3634);
and U1511 (N_1511,In_4568,In_1431);
nand U1512 (N_1512,In_1096,In_1450);
nand U1513 (N_1513,In_4267,In_190);
and U1514 (N_1514,In_2322,In_4862);
xnor U1515 (N_1515,In_3805,In_657);
nor U1516 (N_1516,In_2785,In_1020);
xnor U1517 (N_1517,In_1325,In_2229);
xnor U1518 (N_1518,In_3389,In_4842);
nor U1519 (N_1519,In_3198,In_4543);
xnor U1520 (N_1520,In_700,In_1534);
or U1521 (N_1521,In_1161,In_4500);
xnor U1522 (N_1522,In_3777,In_1340);
nand U1523 (N_1523,In_4641,In_4221);
nor U1524 (N_1524,In_3817,In_647);
xor U1525 (N_1525,In_4653,In_4741);
nor U1526 (N_1526,In_4607,In_4451);
nor U1527 (N_1527,In_263,In_3190);
nor U1528 (N_1528,In_2111,In_289);
nor U1529 (N_1529,In_1798,In_470);
nor U1530 (N_1530,In_1731,In_168);
or U1531 (N_1531,In_4864,In_2255);
and U1532 (N_1532,In_4441,In_1734);
xnor U1533 (N_1533,In_4235,In_659);
nand U1534 (N_1534,In_2417,In_2050);
or U1535 (N_1535,In_1643,In_3435);
xnor U1536 (N_1536,In_4822,In_2671);
nor U1537 (N_1537,In_2585,In_3325);
xor U1538 (N_1538,In_215,In_2155);
xor U1539 (N_1539,In_3462,In_4349);
and U1540 (N_1540,In_2451,In_4456);
nand U1541 (N_1541,In_2035,In_3706);
nand U1542 (N_1542,In_4461,In_1306);
xor U1543 (N_1543,In_4998,In_115);
xnor U1544 (N_1544,In_1834,In_1851);
and U1545 (N_1545,In_338,In_4362);
nand U1546 (N_1546,In_3862,In_1209);
xnor U1547 (N_1547,In_291,In_2925);
or U1548 (N_1548,In_4617,In_3337);
xnor U1549 (N_1549,In_3636,In_4302);
nor U1550 (N_1550,In_1555,In_4946);
xnor U1551 (N_1551,In_4091,In_573);
or U1552 (N_1552,In_1483,In_440);
and U1553 (N_1553,In_3125,In_118);
nand U1554 (N_1554,In_3955,In_4605);
nor U1555 (N_1555,In_2047,In_807);
nand U1556 (N_1556,In_3648,In_4200);
nand U1557 (N_1557,In_4185,In_3336);
and U1558 (N_1558,In_1037,In_3994);
and U1559 (N_1559,In_1973,In_373);
and U1560 (N_1560,In_93,In_888);
and U1561 (N_1561,In_3497,In_3134);
nor U1562 (N_1562,In_1971,In_3206);
nor U1563 (N_1563,In_4292,In_3959);
nor U1564 (N_1564,In_1213,In_2685);
nor U1565 (N_1565,In_3153,In_1813);
or U1566 (N_1566,In_2645,In_57);
xor U1567 (N_1567,In_1138,In_702);
nand U1568 (N_1568,In_3992,In_2662);
xor U1569 (N_1569,In_4415,In_466);
nand U1570 (N_1570,In_2387,In_3718);
or U1571 (N_1571,In_1254,In_2214);
nand U1572 (N_1572,In_4927,In_3298);
or U1573 (N_1573,In_4190,In_1446);
nor U1574 (N_1574,In_4737,In_897);
and U1575 (N_1575,In_3136,In_2331);
nand U1576 (N_1576,In_569,In_898);
xor U1577 (N_1577,In_3593,In_4412);
nor U1578 (N_1578,In_3723,In_1359);
and U1579 (N_1579,In_367,In_936);
nor U1580 (N_1580,In_4657,In_1315);
xnor U1581 (N_1581,In_1335,In_3063);
and U1582 (N_1582,In_4452,In_2936);
nor U1583 (N_1583,In_4562,In_3267);
xnor U1584 (N_1584,In_336,In_1406);
xnor U1585 (N_1585,In_1626,In_4088);
or U1586 (N_1586,In_834,In_1507);
nor U1587 (N_1587,In_4838,In_1267);
nor U1588 (N_1588,In_2083,In_3873);
xor U1589 (N_1589,In_1566,In_4179);
or U1590 (N_1590,In_4586,In_3213);
nor U1591 (N_1591,In_342,In_3191);
nor U1592 (N_1592,In_3857,In_4665);
or U1593 (N_1593,In_3549,In_4709);
and U1594 (N_1594,In_4040,In_2025);
nor U1595 (N_1595,In_4058,In_2097);
nor U1596 (N_1596,In_4163,In_167);
nor U1597 (N_1597,In_2516,In_3978);
nand U1598 (N_1598,In_863,In_2590);
and U1599 (N_1599,In_2754,In_927);
and U1600 (N_1600,In_2838,In_2542);
xor U1601 (N_1601,In_2730,In_435);
xor U1602 (N_1602,In_2746,In_2587);
or U1603 (N_1603,In_1516,In_2380);
and U1604 (N_1604,In_321,In_3525);
nand U1605 (N_1605,In_2156,In_2921);
or U1606 (N_1606,In_3176,In_4245);
and U1607 (N_1607,In_3210,In_822);
and U1608 (N_1608,In_1596,In_1088);
and U1609 (N_1609,In_1402,In_3775);
and U1610 (N_1610,In_2012,In_175);
nand U1611 (N_1611,In_4169,In_1577);
or U1612 (N_1612,In_1203,In_1109);
or U1613 (N_1613,In_3253,In_1015);
and U1614 (N_1614,In_1651,In_227);
nor U1615 (N_1615,In_1965,In_4572);
nand U1616 (N_1616,In_1713,In_411);
nand U1617 (N_1617,In_3965,In_4506);
xnor U1618 (N_1618,In_4825,In_129);
or U1619 (N_1619,In_598,In_4888);
and U1620 (N_1620,In_3304,In_1821);
nor U1621 (N_1621,In_2596,In_4207);
or U1622 (N_1622,In_2611,In_131);
xor U1623 (N_1623,In_4159,In_1290);
nor U1624 (N_1624,In_197,In_1533);
nand U1625 (N_1625,In_4507,In_4991);
nor U1626 (N_1626,In_2455,In_340);
nand U1627 (N_1627,In_516,In_283);
or U1628 (N_1628,In_81,In_3284);
and U1629 (N_1629,In_1886,In_3934);
nand U1630 (N_1630,In_4449,In_1292);
nand U1631 (N_1631,In_1698,In_1929);
nor U1632 (N_1632,In_3563,In_4712);
xnor U1633 (N_1633,In_3881,In_3331);
and U1634 (N_1634,In_1840,In_1925);
nand U1635 (N_1635,In_541,In_184);
xnor U1636 (N_1636,In_3148,In_4992);
and U1637 (N_1637,In_4370,In_1374);
nor U1638 (N_1638,In_2419,In_1448);
or U1639 (N_1639,In_4488,In_2220);
xor U1640 (N_1640,In_1972,In_1693);
or U1641 (N_1641,In_296,In_521);
and U1642 (N_1642,In_4599,In_4271);
and U1643 (N_1643,In_4022,In_2426);
and U1644 (N_1644,In_3019,In_1304);
or U1645 (N_1645,In_2375,In_4645);
or U1646 (N_1646,In_1195,In_3431);
and U1647 (N_1647,In_4720,In_4625);
nor U1648 (N_1648,In_1248,In_2616);
nor U1649 (N_1649,In_3027,In_2554);
nand U1650 (N_1650,In_665,In_2178);
nor U1651 (N_1651,In_1268,In_3283);
or U1652 (N_1652,In_1579,In_457);
nor U1653 (N_1653,In_2720,In_2589);
and U1654 (N_1654,In_4798,In_2679);
xor U1655 (N_1655,In_567,In_2760);
and U1656 (N_1656,In_71,In_4222);
nor U1657 (N_1657,In_36,In_2148);
nand U1658 (N_1658,In_2045,In_7);
or U1659 (N_1659,In_4462,In_986);
nor U1660 (N_1660,In_3615,In_2663);
nor U1661 (N_1661,In_990,In_1513);
nand U1662 (N_1662,In_1122,In_2134);
xor U1663 (N_1663,In_1602,In_1981);
nor U1664 (N_1664,In_2681,In_2791);
and U1665 (N_1665,In_1530,In_4083);
or U1666 (N_1666,In_2546,In_3930);
or U1667 (N_1667,In_2268,In_1649);
nor U1668 (N_1668,In_505,In_4282);
nand U1669 (N_1669,In_4118,In_4661);
xnor U1670 (N_1670,In_1781,In_2420);
nor U1671 (N_1671,In_1811,In_248);
or U1672 (N_1672,In_1168,In_916);
xnor U1673 (N_1673,In_1354,In_1554);
xnor U1674 (N_1674,In_3686,In_2906);
and U1675 (N_1675,In_3307,In_2558);
nand U1676 (N_1676,In_3606,In_3625);
and U1677 (N_1677,In_1204,In_2792);
nand U1678 (N_1678,In_3259,In_4385);
or U1679 (N_1679,In_1311,In_2793);
nand U1680 (N_1680,In_2491,In_1560);
xnor U1681 (N_1681,In_4987,In_2059);
or U1682 (N_1682,In_3595,In_1392);
and U1683 (N_1683,In_4638,In_2166);
and U1684 (N_1684,In_4960,In_3346);
nand U1685 (N_1685,In_4800,In_3951);
xor U1686 (N_1686,In_4027,In_4670);
xor U1687 (N_1687,In_1921,In_4582);
or U1688 (N_1688,In_826,In_4138);
nand U1689 (N_1689,In_3616,In_90);
xnor U1690 (N_1690,In_3165,In_3659);
xor U1691 (N_1691,In_1246,In_2658);
nand U1692 (N_1692,In_780,In_840);
and U1693 (N_1693,In_1920,In_950);
nor U1694 (N_1694,In_2799,In_3989);
or U1695 (N_1695,In_3281,In_1669);
or U1696 (N_1696,In_1110,In_1889);
and U1697 (N_1697,In_4315,In_277);
xnor U1698 (N_1698,In_4371,In_1461);
or U1699 (N_1699,In_4539,In_3820);
or U1700 (N_1700,In_4028,In_3084);
nand U1701 (N_1701,In_1280,In_3030);
nand U1702 (N_1702,In_607,In_1659);
xnor U1703 (N_1703,In_169,In_4158);
nand U1704 (N_1704,In_3641,In_3559);
nand U1705 (N_1705,In_310,In_2859);
xnor U1706 (N_1706,In_2291,In_996);
and U1707 (N_1707,In_1395,In_538);
xor U1708 (N_1708,In_1827,In_1949);
or U1709 (N_1709,In_2577,In_314);
nand U1710 (N_1710,In_234,In_3536);
nand U1711 (N_1711,In_2923,In_1046);
nor U1712 (N_1712,In_3936,In_4846);
nor U1713 (N_1713,In_696,In_3897);
and U1714 (N_1714,In_2511,In_2970);
nor U1715 (N_1715,In_3756,In_2956);
nand U1716 (N_1716,In_2883,In_2814);
and U1717 (N_1717,In_3333,In_4108);
nand U1718 (N_1718,In_1584,In_400);
or U1719 (N_1719,In_2878,In_4129);
or U1720 (N_1720,In_4906,In_1357);
or U1721 (N_1721,In_222,In_872);
nor U1722 (N_1722,In_580,In_4760);
xor U1723 (N_1723,In_2250,In_55);
nor U1724 (N_1724,In_4168,In_911);
nor U1725 (N_1725,In_3664,In_74);
xnor U1726 (N_1726,In_4965,In_2193);
nor U1727 (N_1727,In_4056,In_1137);
nor U1728 (N_1728,In_3392,In_798);
or U1729 (N_1729,In_4621,In_1546);
or U1730 (N_1730,In_1162,In_4938);
nand U1731 (N_1731,In_362,In_4931);
xor U1732 (N_1732,In_4899,In_1293);
nand U1733 (N_1733,In_1050,In_4735);
or U1734 (N_1734,In_1775,In_2129);
nor U1735 (N_1735,In_2813,In_1599);
or U1736 (N_1736,In_2381,In_3135);
and U1737 (N_1737,In_2081,In_586);
and U1738 (N_1738,In_2648,In_1136);
xor U1739 (N_1739,In_1803,In_1415);
nor U1740 (N_1740,In_682,In_3576);
nor U1741 (N_1741,In_2911,In_1291);
xor U1742 (N_1742,In_3879,In_681);
nor U1743 (N_1743,In_4079,In_1583);
xor U1744 (N_1744,In_654,In_448);
nand U1745 (N_1745,In_371,In_2715);
nand U1746 (N_1746,In_4708,In_1716);
nand U1747 (N_1747,In_4288,In_4177);
nor U1748 (N_1748,In_947,In_514);
nand U1749 (N_1749,In_472,In_4387);
and U1750 (N_1750,In_1371,In_756);
nand U1751 (N_1751,In_655,In_4003);
nand U1752 (N_1752,In_417,In_3865);
nand U1753 (N_1753,In_1424,In_4065);
nand U1754 (N_1754,In_1022,In_2197);
nand U1755 (N_1755,In_1635,In_3272);
and U1756 (N_1756,In_2037,In_450);
nor U1757 (N_1757,In_1910,In_1422);
nand U1758 (N_1758,In_3754,In_907);
xnor U1759 (N_1759,In_3519,In_769);
nor U1760 (N_1760,In_1352,In_4598);
nor U1761 (N_1761,In_1688,In_2588);
nand U1762 (N_1762,In_962,In_1957);
xnor U1763 (N_1763,In_4947,In_2078);
nor U1764 (N_1764,In_4254,In_1414);
or U1765 (N_1765,In_2634,In_1428);
and U1766 (N_1766,In_2191,In_638);
nand U1767 (N_1767,In_149,In_1970);
or U1768 (N_1768,In_980,In_2004);
and U1769 (N_1769,In_28,In_4929);
or U1770 (N_1770,In_1420,In_4390);
or U1771 (N_1771,In_765,In_2625);
xor U1772 (N_1772,In_1569,In_3954);
xor U1773 (N_1773,In_4361,In_1790);
nor U1774 (N_1774,In_1353,In_4374);
or U1775 (N_1775,In_4941,In_4742);
nand U1776 (N_1776,In_949,In_4952);
and U1777 (N_1777,In_1512,In_4527);
and U1778 (N_1778,In_1982,In_3583);
nand U1779 (N_1779,In_3574,In_4155);
nor U1780 (N_1780,In_4219,In_2459);
and U1781 (N_1781,In_3147,In_401);
nor U1782 (N_1782,In_4464,In_4117);
or U1783 (N_1783,In_2696,In_94);
nor U1784 (N_1784,In_2868,In_4123);
nor U1785 (N_1785,In_4634,In_2790);
and U1786 (N_1786,In_462,In_48);
nand U1787 (N_1787,In_1436,In_1011);
or U1788 (N_1788,In_2533,In_1487);
nand U1789 (N_1789,In_4953,In_2382);
and U1790 (N_1790,In_1333,In_1666);
xnor U1791 (N_1791,In_1361,In_3123);
nand U1792 (N_1792,In_1080,In_3443);
xnor U1793 (N_1793,In_1451,In_603);
nand U1794 (N_1794,In_1445,In_154);
nor U1795 (N_1795,In_4610,In_2010);
or U1796 (N_1796,In_1791,In_4355);
and U1797 (N_1797,In_3447,In_443);
xnor U1798 (N_1798,In_261,In_3033);
nor U1799 (N_1799,In_3907,In_3633);
xor U1800 (N_1800,In_1737,In_543);
nor U1801 (N_1801,In_37,In_618);
nand U1802 (N_1802,In_2708,In_4013);
or U1803 (N_1803,In_4428,In_1062);
nor U1804 (N_1804,In_2991,In_774);
nand U1805 (N_1805,In_89,In_1282);
xnor U1806 (N_1806,In_971,In_2682);
nor U1807 (N_1807,In_2665,In_1517);
nor U1808 (N_1808,In_613,In_1658);
nor U1809 (N_1809,In_524,In_4055);
nand U1810 (N_1810,In_4600,In_1644);
or U1811 (N_1811,In_4074,In_328);
nand U1812 (N_1812,In_1524,In_1500);
nor U1813 (N_1813,In_3933,In_2603);
and U1814 (N_1814,In_4319,In_2857);
xor U1815 (N_1815,In_2586,In_1063);
xnor U1816 (N_1816,In_1170,In_3903);
xor U1817 (N_1817,In_1815,In_306);
nand U1818 (N_1818,In_3998,In_4291);
xnor U1819 (N_1819,In_2402,In_2345);
xor U1820 (N_1820,In_1677,In_392);
nor U1821 (N_1821,In_1763,In_3908);
or U1822 (N_1822,In_1197,In_4054);
xnor U1823 (N_1823,In_728,In_902);
nor U1824 (N_1824,In_2567,In_1418);
or U1825 (N_1825,In_3551,In_193);
or U1826 (N_1826,In_4405,In_1989);
xnor U1827 (N_1827,In_2501,In_919);
and U1828 (N_1828,In_3494,In_2961);
nand U1829 (N_1829,In_4403,In_4891);
xnor U1830 (N_1830,In_2349,In_760);
and U1831 (N_1831,In_3420,In_3364);
and U1832 (N_1832,In_4937,In_1172);
xnor U1833 (N_1833,In_583,In_2958);
and U1834 (N_1834,In_1378,In_4901);
and U1835 (N_1835,In_956,In_3815);
xor U1836 (N_1836,In_3966,In_3113);
and U1837 (N_1837,In_2528,In_1476);
or U1838 (N_1838,In_1621,In_2297);
nor U1839 (N_1839,In_4967,In_3644);
and U1840 (N_1840,In_673,In_4135);
nand U1841 (N_1841,In_1255,In_994);
xor U1842 (N_1842,In_1043,In_1877);
or U1843 (N_1843,In_3145,In_2179);
nor U1844 (N_1844,In_687,In_658);
nand U1845 (N_1845,In_3567,In_3032);
nor U1846 (N_1846,In_467,In_454);
and U1847 (N_1847,In_2140,In_894);
xnor U1848 (N_1848,In_1960,In_858);
or U1849 (N_1849,In_1348,In_4627);
or U1850 (N_1850,In_138,In_2901);
and U1851 (N_1851,In_3396,In_2340);
or U1852 (N_1852,In_3500,In_3647);
xor U1853 (N_1853,In_393,In_944);
nand U1854 (N_1854,In_18,In_2130);
nand U1855 (N_1855,In_967,In_127);
nor U1856 (N_1856,In_4903,In_3496);
nand U1857 (N_1857,In_3248,In_249);
or U1858 (N_1858,In_2385,In_4309);
or U1859 (N_1859,In_1247,In_2721);
or U1860 (N_1860,In_4394,In_3531);
or U1861 (N_1861,In_3450,In_2620);
xnor U1862 (N_1862,In_4216,In_2469);
and U1863 (N_1863,In_1457,In_4038);
xor U1864 (N_1864,In_3923,In_2607);
nand U1865 (N_1865,In_3588,In_3436);
and U1866 (N_1866,In_181,In_1756);
nor U1867 (N_1867,In_2259,In_3174);
and U1868 (N_1868,In_2741,In_2495);
xor U1869 (N_1869,In_719,In_3161);
or U1870 (N_1870,In_1100,In_3770);
and U1871 (N_1871,In_2743,In_379);
nand U1872 (N_1872,In_3289,In_4243);
or U1873 (N_1873,In_4344,In_4264);
xor U1874 (N_1874,In_1385,In_3975);
nor U1875 (N_1875,In_1824,In_50);
xnor U1876 (N_1876,In_4636,In_1259);
xor U1877 (N_1877,In_929,In_2244);
nand U1878 (N_1878,In_3950,In_3096);
or U1879 (N_1879,In_2750,In_2125);
or U1880 (N_1880,In_3279,In_302);
and U1881 (N_1881,In_433,In_2667);
nor U1882 (N_1882,In_3067,In_1303);
and U1883 (N_1883,In_326,In_1177);
xor U1884 (N_1884,In_334,In_561);
nand U1885 (N_1885,In_737,In_2827);
or U1886 (N_1886,In_4092,In_1262);
xor U1887 (N_1887,In_3851,In_2269);
and U1888 (N_1888,In_4303,In_1289);
nor U1889 (N_1889,In_1792,In_3038);
xnor U1890 (N_1890,In_1704,In_4432);
or U1891 (N_1891,In_4801,In_2828);
or U1892 (N_1892,In_2236,In_2107);
and U1893 (N_1893,In_2316,In_2131);
and U1894 (N_1894,In_14,In_3572);
nand U1895 (N_1895,In_1543,In_2404);
nand U1896 (N_1896,In_2202,In_449);
xnor U1897 (N_1897,In_1613,In_59);
and U1898 (N_1898,In_2782,In_3709);
and U1899 (N_1899,In_1783,In_1111);
or U1900 (N_1900,In_4463,In_2650);
and U1901 (N_1901,In_1995,In_1712);
xor U1902 (N_1902,In_113,In_751);
and U1903 (N_1903,In_1250,In_1029);
nand U1904 (N_1904,In_3976,In_4986);
nand U1905 (N_1905,In_1723,In_917);
and U1906 (N_1906,In_1549,In_1394);
nor U1907 (N_1907,In_2457,In_4111);
nand U1908 (N_1908,In_3856,In_3089);
or U1909 (N_1909,In_4524,In_1992);
nor U1910 (N_1910,In_1998,In_1045);
xnor U1911 (N_1911,In_1028,In_2212);
or U1912 (N_1912,In_358,In_1245);
xor U1913 (N_1913,In_4493,In_1955);
or U1914 (N_1914,In_4536,In_337);
xnor U1915 (N_1915,In_4277,In_2907);
nor U1916 (N_1916,In_4268,In_4951);
nor U1917 (N_1917,In_3795,In_1178);
nor U1918 (N_1918,In_554,In_3988);
and U1919 (N_1919,In_484,In_2232);
and U1920 (N_1920,In_1308,In_4528);
nand U1921 (N_1921,In_1336,In_4071);
xor U1922 (N_1922,In_3297,In_4218);
or U1923 (N_1923,In_3369,In_3514);
or U1924 (N_1924,In_3335,In_3712);
or U1925 (N_1925,In_284,In_942);
or U1926 (N_1926,In_329,In_10);
xor U1927 (N_1927,In_656,In_1637);
nor U1928 (N_1928,In_4171,In_2870);
nor U1929 (N_1929,In_3535,In_790);
or U1930 (N_1930,In_2524,In_2067);
xor U1931 (N_1931,In_3013,In_4211);
xor U1932 (N_1932,In_2604,In_4830);
nand U1933 (N_1933,In_2243,In_1726);
nor U1934 (N_1934,In_1678,In_3798);
and U1935 (N_1935,In_1496,In_3217);
or U1936 (N_1936,In_1141,In_4016);
or U1937 (N_1937,In_4289,In_2164);
xnor U1938 (N_1938,In_2034,In_2369);
and U1939 (N_1939,In_2006,In_4596);
nor U1940 (N_1940,In_4950,In_3384);
nand U1941 (N_1941,In_1660,In_4643);
and U1942 (N_1942,In_251,In_3848);
or U1943 (N_1943,In_4007,In_4663);
and U1944 (N_1944,In_4157,In_4107);
nand U1945 (N_1945,In_3612,In_1933);
nor U1946 (N_1946,In_3991,In_725);
and U1947 (N_1947,In_745,In_4894);
nand U1948 (N_1948,In_4697,In_1438);
nor U1949 (N_1949,In_528,In_901);
nand U1950 (N_1950,In_455,In_3970);
nand U1951 (N_1951,In_4376,In_2151);
or U1952 (N_1952,In_4410,In_4400);
nand U1953 (N_1953,In_4804,In_3044);
or U1954 (N_1954,In_4265,In_2834);
nor U1955 (N_1955,In_2762,In_1867);
xor U1956 (N_1956,In_1614,In_4075);
nand U1957 (N_1957,In_356,In_3618);
xnor U1958 (N_1958,In_116,In_1104);
nor U1959 (N_1959,In_799,In_2965);
nor U1960 (N_1960,In_4072,In_4818);
or U1961 (N_1961,In_3322,In_4993);
or U1962 (N_1962,In_485,In_1510);
nand U1963 (N_1963,In_3007,In_2406);
nor U1964 (N_1964,In_2213,In_157);
nor U1965 (N_1965,In_874,In_1894);
or U1966 (N_1966,In_1941,In_1082);
xor U1967 (N_1967,In_3196,In_3412);
nand U1968 (N_1968,In_1810,In_241);
or U1969 (N_1969,In_12,In_3568);
xnor U1970 (N_1970,In_3046,In_1627);
nor U1971 (N_1971,In_1069,In_2652);
nor U1972 (N_1972,In_1697,In_793);
nor U1973 (N_1973,In_2610,In_3449);
xnor U1974 (N_1974,In_920,In_3530);
nor U1975 (N_1975,In_4813,In_4094);
nand U1976 (N_1976,In_4728,In_2479);
and U1977 (N_1977,In_2986,In_3334);
xor U1978 (N_1978,In_312,In_4429);
or U1979 (N_1979,In_1520,In_1486);
nand U1980 (N_1980,In_861,In_2545);
nand U1981 (N_1981,In_4602,In_3799);
and U1982 (N_1982,In_2695,In_213);
nor U1983 (N_1983,In_2518,In_1856);
nand U1984 (N_1984,In_3299,In_4102);
nand U1985 (N_1985,In_1051,In_575);
or U1986 (N_1986,In_4044,In_1953);
nor U1987 (N_1987,In_4731,In_1059);
or U1988 (N_1988,In_4691,In_3550);
or U1989 (N_1989,In_2458,In_2903);
xnor U1990 (N_1990,In_992,In_4940);
xor U1991 (N_1991,In_3292,In_1559);
and U1992 (N_1992,In_1429,In_4306);
or U1993 (N_1993,In_3107,In_1709);
nand U1994 (N_1994,In_4470,In_2371);
nor U1995 (N_1995,In_4173,In_4782);
or U1996 (N_1996,In_4125,In_1831);
xor U1997 (N_1997,In_2756,In_1892);
nand U1998 (N_1998,In_823,In_2816);
nor U1999 (N_1999,In_1389,In_970);
nor U2000 (N_2000,In_1695,In_3491);
nand U2001 (N_2001,In_601,In_4115);
or U2002 (N_2002,In_3105,In_2496);
and U2003 (N_2003,In_4626,In_4873);
nand U2004 (N_2004,In_3926,In_4139);
or U2005 (N_2005,In_557,In_2599);
xnor U2006 (N_2006,In_2265,In_1286);
nor U2007 (N_2007,In_2436,In_2287);
nor U2008 (N_2008,In_2328,In_4979);
or U2009 (N_2009,In_1679,In_3074);
and U2010 (N_2010,In_3943,In_2396);
or U2011 (N_2011,In_3556,In_3010);
xnor U2012 (N_2012,In_353,In_1146);
and U2013 (N_2013,In_3348,In_3767);
nor U2014 (N_2014,In_3810,In_1318);
xnor U2015 (N_2015,In_582,In_40);
or U2016 (N_2016,In_2013,In_311);
nor U2017 (N_2017,In_3118,In_4247);
nand U2018 (N_2018,In_1714,In_3691);
or U2019 (N_2019,In_2418,In_2113);
nor U2020 (N_2020,In_4398,In_2632);
xnor U2021 (N_2021,In_859,In_1155);
nand U2022 (N_2022,In_3661,In_2806);
nor U2023 (N_2023,In_4465,In_3958);
nand U2024 (N_2024,In_3771,In_3528);
and U2025 (N_2025,In_4613,In_999);
nand U2026 (N_2026,In_2499,In_943);
nand U2027 (N_2027,In_31,In_3800);
and U2028 (N_2028,In_781,In_1455);
xor U2029 (N_2029,In_4411,In_1356);
and U2030 (N_2030,In_3502,In_1115);
xnor U2031 (N_2031,In_1905,In_4166);
nand U2032 (N_2032,In_4313,In_1498);
xnor U2033 (N_2033,In_1804,In_3866);
and U2034 (N_2034,In_504,In_1872);
nor U2035 (N_2035,In_3478,In_2184);
xor U2036 (N_2036,In_374,In_3122);
xor U2037 (N_2037,In_830,In_1564);
xnor U2038 (N_2038,In_982,In_395);
and U2039 (N_2039,In_4045,In_1773);
or U2040 (N_2040,In_850,In_3085);
nor U2041 (N_2041,In_1591,In_876);
nor U2042 (N_2042,In_79,In_609);
nand U2043 (N_2043,In_508,In_458);
nor U2044 (N_2044,In_3523,In_3026);
or U2045 (N_2045,In_3066,In_2136);
or U2046 (N_2046,In_3488,In_4774);
or U2047 (N_2047,In_228,In_1345);
nand U2048 (N_2048,In_387,In_4141);
nor U2049 (N_2049,In_1875,In_3607);
or U2050 (N_2050,In_617,In_339);
and U2051 (N_2051,In_3181,In_0);
nand U2052 (N_2052,In_3481,In_3999);
xor U2053 (N_2053,In_3221,In_2905);
nor U2054 (N_2054,In_292,In_1148);
or U2055 (N_2055,In_817,In_4517);
nand U2056 (N_2056,In_1885,In_644);
nor U2057 (N_2057,In_1692,In_2691);
and U2058 (N_2058,In_4537,In_1574);
nor U2059 (N_2059,In_2688,In_2377);
nor U2060 (N_2060,In_403,In_1473);
and U2061 (N_2061,In_2133,In_1072);
nand U2062 (N_2062,In_1081,In_1421);
or U2063 (N_2063,In_4765,In_434);
and U2064 (N_2064,In_67,In_4203);
or U2065 (N_2065,In_191,In_2014);
or U2066 (N_2066,In_1470,In_2044);
xor U2067 (N_2067,In_3979,In_535);
and U2068 (N_2068,In_2302,In_2186);
and U2069 (N_2069,In_928,In_3254);
and U2070 (N_2070,In_4226,In_1270);
and U2071 (N_2071,In_4832,In_1274);
and U2072 (N_2072,In_2256,In_4212);
or U2073 (N_2073,In_2415,In_608);
xor U2074 (N_2074,In_4805,In_3630);
or U2075 (N_2075,In_1226,In_2592);
or U2076 (N_2076,In_1654,In_2670);
and U2077 (N_2077,In_2355,In_4748);
xor U2078 (N_2078,In_2975,In_3602);
nand U2079 (N_2079,In_3367,In_1091);
or U2080 (N_2080,In_619,In_3345);
nor U2081 (N_2081,In_1241,In_4352);
and U2082 (N_2082,In_2716,In_3831);
xor U2083 (N_2083,In_1123,In_3099);
nor U2084 (N_2084,In_2261,In_3816);
nand U2085 (N_2085,In_83,In_352);
and U2086 (N_2086,In_4348,In_3996);
nand U2087 (N_2087,In_3710,In_16);
and U2088 (N_2088,In_126,In_1891);
xnor U2089 (N_2089,In_1782,In_2195);
and U2090 (N_2090,In_2173,In_2656);
or U2091 (N_2091,In_3100,In_2969);
nor U2092 (N_2092,In_2022,In_124);
and U2093 (N_2093,In_1685,In_4718);
or U2094 (N_2094,In_3787,In_4821);
xor U2095 (N_2095,In_3913,In_495);
xnor U2096 (N_2096,In_4549,In_1528);
xor U2097 (N_2097,In_1220,In_594);
xor U2098 (N_2098,In_3170,In_1493);
nand U2099 (N_2099,In_3454,In_1273);
xor U2100 (N_2100,In_2692,In_70);
nand U2101 (N_2101,In_332,In_3826);
nor U2102 (N_2102,In_300,In_3738);
or U2103 (N_2103,In_180,In_4109);
xnor U2104 (N_2104,In_4637,In_4285);
or U2105 (N_2105,In_3160,In_4366);
nor U2106 (N_2106,In_882,In_2020);
xnor U2107 (N_2107,In_4299,In_1794);
nor U2108 (N_2108,In_3194,In_2048);
nor U2109 (N_2109,In_1349,In_3015);
and U2110 (N_2110,In_2732,In_4928);
nor U2111 (N_2111,In_3189,In_4973);
and U2112 (N_2112,In_4902,In_4563);
xnor U2113 (N_2113,In_305,In_1595);
and U2114 (N_2114,In_1004,In_1655);
and U2115 (N_2115,In_1182,In_2976);
xor U2116 (N_2116,In_4380,In_3794);
nand U2117 (N_2117,In_4068,In_1472);
nand U2118 (N_2118,In_2429,In_1525);
or U2119 (N_2119,In_3480,In_4880);
nor U2120 (N_2120,In_3524,In_525);
nand U2121 (N_2121,In_1904,In_3313);
or U2122 (N_2122,In_238,In_2579);
nand U2123 (N_2123,In_1117,In_4851);
xnor U2124 (N_2124,In_4409,In_4413);
xnor U2125 (N_2125,In_474,In_4041);
nor U2126 (N_2126,In_4165,In_4328);
or U2127 (N_2127,In_4664,In_2181);
nor U2128 (N_2128,In_2678,In_3275);
and U2129 (N_2129,In_2563,In_3872);
and U2130 (N_2130,In_2498,In_3722);
xor U2131 (N_2131,In_4082,In_1219);
and U2132 (N_2132,In_4833,In_3997);
nand U2133 (N_2133,In_818,In_2600);
nand U2134 (N_2134,In_1331,In_1733);
or U2135 (N_2135,In_3274,In_855);
or U2136 (N_2136,In_4881,In_3655);
xnor U2137 (N_2137,In_137,In_3064);
or U2138 (N_2138,In_1634,In_4073);
nor U2139 (N_2139,In_317,In_723);
xor U2140 (N_2140,In_975,In_1031);
xnor U2141 (N_2141,In_3849,In_4126);
or U2142 (N_2142,In_27,In_2774);
or U2143 (N_2143,In_3048,In_3163);
nor U2144 (N_2144,In_3824,In_3168);
nor U2145 (N_2145,In_4632,In_4255);
and U2146 (N_2146,In_3006,In_2373);
nor U2147 (N_2147,In_2024,In_2631);
or U2148 (N_2148,In_1948,In_2748);
nor U2149 (N_2149,In_1956,In_842);
nand U2150 (N_2150,In_584,In_4884);
nor U2151 (N_2151,In_4921,In_604);
and U2152 (N_2152,In_4472,In_4444);
nor U2153 (N_2153,In_4261,In_3765);
or U2154 (N_2154,In_1959,In_549);
and U2155 (N_2155,In_3162,In_4743);
nor U2156 (N_2156,In_4033,In_672);
nand U2157 (N_2157,In_2571,In_2270);
xor U2158 (N_2158,In_3091,In_151);
or U2159 (N_2159,In_3571,In_2781);
nor U2160 (N_2160,In_2867,In_1958);
and U2161 (N_2161,In_1358,In_216);
xor U2162 (N_2162,In_1099,In_1849);
nor U2163 (N_2163,In_4908,In_972);
and U2164 (N_2164,In_2365,In_2058);
nor U2165 (N_2165,In_4310,In_4393);
xor U2166 (N_2166,In_4791,In_4246);
nand U2167 (N_2167,In_2753,In_250);
xor U2168 (N_2168,In_1208,In_787);
nand U2169 (N_2169,In_418,In_1369);
or U2170 (N_2170,In_2425,In_4984);
xor U2171 (N_2171,In_2088,In_4504);
nor U2172 (N_2172,In_2211,In_2273);
nand U2173 (N_2173,In_4700,In_2180);
and U2174 (N_2174,In_430,In_383);
xnor U2175 (N_2175,In_1194,In_4103);
or U2176 (N_2176,In_3665,In_3418);
xnor U2177 (N_2177,In_451,In_1364);
nand U2178 (N_2178,In_2023,In_3422);
nor U2179 (N_2179,In_3250,In_3886);
nand U2180 (N_2180,In_3409,In_4087);
and U2181 (N_2181,In_4546,In_3605);
nor U2182 (N_2182,In_1300,In_836);
xnor U2183 (N_2183,In_2947,In_1302);
or U2184 (N_2184,In_2079,In_4420);
nor U2185 (N_2185,In_2739,In_4148);
or U2186 (N_2186,In_4564,In_1893);
nand U2187 (N_2187,In_3434,In_4591);
nor U2188 (N_2188,In_1054,In_1808);
and U2189 (N_2189,In_2968,In_3939);
nand U2190 (N_2190,In_794,In_3199);
or U2191 (N_2191,In_1909,In_1561);
nand U2192 (N_2192,In_1196,In_3180);
or U2193 (N_2193,In_4548,In_1547);
or U2194 (N_2194,In_1617,In_4674);
nor U2195 (N_2195,In_3286,In_2364);
nor U2196 (N_2196,In_3441,In_3697);
and U2197 (N_2197,In_413,In_2728);
xor U2198 (N_2198,In_4848,In_4014);
nand U2199 (N_2199,In_2505,In_3784);
nand U2200 (N_2200,In_2409,In_281);
and U2201 (N_2201,In_1452,In_1218);
nand U2202 (N_2202,In_3788,In_1416);
and U2203 (N_2203,In_4739,In_77);
and U2204 (N_2204,In_566,In_2918);
and U2205 (N_2205,In_3914,In_2981);
xnor U2206 (N_2206,In_166,In_121);
or U2207 (N_2207,In_4573,In_3883);
nand U2208 (N_2208,In_2974,In_179);
and U2209 (N_2209,In_3028,In_1089);
nor U2210 (N_2210,In_3446,In_1606);
xnor U2211 (N_2211,In_3197,In_1033);
and U2212 (N_2212,In_3791,In_2257);
nand U2213 (N_2213,In_4063,In_468);
nand U2214 (N_2214,In_3726,In_1163);
nand U2215 (N_2215,In_2052,In_4867);
xor U2216 (N_2216,In_1661,In_1565);
and U2217 (N_2217,In_4766,In_3236);
nor U2218 (N_2218,In_2100,In_3296);
and U2219 (N_2219,In_1847,In_389);
xnor U2220 (N_2220,In_3878,In_3755);
and U2221 (N_2221,In_4172,In_2372);
and U2222 (N_2222,In_2635,In_1328);
and U2223 (N_2223,In_3453,In_239);
xnor U2224 (N_2224,In_4887,In_1095);
nand U2225 (N_2225,In_1481,In_2797);
and U2226 (N_2226,In_4750,In_4495);
or U2227 (N_2227,In_578,In_761);
nand U2228 (N_2228,In_4714,In_620);
nor U2229 (N_2229,In_147,In_2196);
xor U2230 (N_2230,In_3143,In_3935);
nor U2231 (N_2231,In_3645,In_1097);
or U2232 (N_2232,In_3779,In_1459);
and U2233 (N_2233,In_4486,In_623);
and U2234 (N_2234,In_3947,In_2288);
nor U2235 (N_2235,In_1812,In_4442);
xor U2236 (N_2236,In_1706,In_201);
nor U2237 (N_2237,In_1176,In_483);
nand U2238 (N_2238,In_3377,In_4988);
nand U2239 (N_2239,In_2998,In_420);
and U2240 (N_2240,In_1807,In_4260);
nor U2241 (N_2241,In_841,In_2109);
xnor U2242 (N_2242,In_2082,In_268);
xor U2243 (N_2243,In_3306,In_3414);
and U2244 (N_2244,In_2972,In_825);
nor U2245 (N_2245,In_2454,In_3065);
and U2246 (N_2246,In_370,In_3200);
nor U2247 (N_2247,In_4329,In_108);
nand U2248 (N_2248,In_4233,In_3745);
and U2249 (N_2249,In_3110,In_2997);
xor U2250 (N_2250,In_4455,In_1151);
or U2251 (N_2251,In_195,In_4457);
nor U2252 (N_2252,In_2593,In_3626);
and U2253 (N_2253,In_98,In_2598);
xor U2254 (N_2254,In_540,In_3867);
and U2255 (N_2255,In_4837,In_1252);
nand U2256 (N_2256,In_1705,In_3916);
and U2257 (N_2257,In_9,In_2787);
nand U2258 (N_2258,In_3704,In_1771);
or U2259 (N_2259,In_1887,In_4338);
nand U2260 (N_2260,In_4863,In_3220);
or U2261 (N_2261,In_4913,In_351);
nor U2262 (N_2262,In_556,In_1074);
and U2263 (N_2263,In_382,In_1329);
or U2264 (N_2264,In_1589,In_782);
nor U2265 (N_2265,In_3356,In_3909);
nor U2266 (N_2266,In_1701,In_3774);
xor U2267 (N_2267,In_343,In_4839);
or U2268 (N_2268,In_1112,In_2209);
or U2269 (N_2269,In_225,In_729);
and U2270 (N_2270,In_3227,In_2309);
xor U2271 (N_2271,In_4784,In_4321);
or U2272 (N_2272,In_1738,In_2641);
xnor U2273 (N_2273,In_3090,In_801);
or U2274 (N_2274,In_3232,In_163);
xnor U2275 (N_2275,In_4029,In_564);
and U2276 (N_2276,In_1149,In_550);
or U2277 (N_2277,In_1736,In_1848);
nand U2278 (N_2278,In_3772,In_1061);
nand U2279 (N_2279,In_1344,In_4133);
nand U2280 (N_2280,In_3087,In_153);
and U2281 (N_2281,In_4920,In_41);
xor U2282 (N_2282,In_1475,In_3079);
nand U2283 (N_2283,In_2336,In_2826);
or U2284 (N_2284,In_2853,In_4248);
and U2285 (N_2285,In_2547,In_4156);
nor U2286 (N_2286,In_3667,In_2094);
nor U2287 (N_2287,In_1934,In_1553);
xor U2288 (N_2288,In_148,In_4479);
and U2289 (N_2289,In_1012,In_2208);
or U2290 (N_2290,In_3440,In_661);
or U2291 (N_2291,In_4018,In_2112);
or U2292 (N_2292,In_3492,In_2060);
xnor U2293 (N_2293,In_3104,In_1548);
nand U2294 (N_2294,In_669,In_993);
or U2295 (N_2295,In_4150,In_432);
xor U2296 (N_2296,In_4511,In_3288);
nor U2297 (N_2297,In_3741,In_86);
nand U2298 (N_2298,In_1741,In_2731);
xor U2299 (N_2299,In_4460,In_4817);
and U2300 (N_2300,In_1580,In_503);
or U2301 (N_2301,In_1641,In_1044);
nor U2302 (N_2302,In_110,In_4565);
nand U2303 (N_2303,In_65,In_4738);
or U2304 (N_2304,In_30,In_4722);
nor U2305 (N_2305,In_2174,In_3808);
nand U2306 (N_2306,In_1817,In_2295);
nand U2307 (N_2307,In_2980,In_2775);
xor U2308 (N_2308,In_2102,In_4754);
xor U2309 (N_2309,In_301,In_4437);
xnor U2310 (N_2310,In_68,In_3801);
nand U2311 (N_2311,In_1174,In_347);
or U2312 (N_2312,In_985,In_1926);
and U2313 (N_2313,In_4703,In_925);
nor U2314 (N_2314,In_4939,In_4011);
or U2315 (N_2315,In_386,In_4024);
nor U2316 (N_2316,In_2619,In_3224);
and U2317 (N_2317,In_2098,In_1786);
or U2318 (N_2318,In_2897,In_1873);
nand U2319 (N_2319,In_2043,In_3188);
or U2320 (N_2320,In_3793,In_422);
nand U2321 (N_2321,In_348,In_3031);
and U2322 (N_2322,In_4732,In_105);
nand U2323 (N_2323,In_4614,In_4747);
nand U2324 (N_2324,In_4589,In_632);
or U2325 (N_2325,In_1048,In_4726);
nor U2326 (N_2326,In_3589,In_4630);
nor U2327 (N_2327,In_2561,In_1724);
and U2328 (N_2328,In_4151,In_3341);
xor U2329 (N_2329,In_2572,In_3351);
and U2330 (N_2330,In_1777,In_4734);
or U2331 (N_2331,In_777,In_2027);
nor U2332 (N_2332,In_1717,In_473);
nor U2333 (N_2333,In_2190,In_1188);
and U2334 (N_2334,In_365,In_4990);
nand U2335 (N_2335,In_4624,In_3675);
nor U2336 (N_2336,In_2177,In_856);
nand U2337 (N_2337,In_960,In_4360);
or U2338 (N_2338,In_1365,In_2891);
xor U2339 (N_2339,In_2875,In_4422);
and U2340 (N_2340,In_3790,In_1125);
and U2341 (N_2341,In_2751,In_2541);
or U2342 (N_2342,In_3282,In_4847);
and U2343 (N_2343,In_1320,In_3870);
xor U2344 (N_2344,In_1468,In_1968);
nand U2345 (N_2345,In_3705,In_4142);
nor U2346 (N_2346,In_2773,In_736);
nand U2347 (N_2347,In_3246,In_4910);
and U2348 (N_2348,In_1895,In_2460);
and U2349 (N_2349,In_3385,In_622);
nor U2350 (N_2350,In_1532,In_3586);
xnor U2351 (N_2351,In_2465,In_3750);
xor U2352 (N_2352,In_1823,In_136);
xor U2353 (N_2353,In_4096,In_3415);
and U2354 (N_2354,In_624,In_1729);
nand U2355 (N_2355,In_686,In_1034);
nor U2356 (N_2356,In_2252,In_2699);
nand U2357 (N_2357,In_4119,In_1027);
or U2358 (N_2358,In_743,In_2594);
nor U2359 (N_2359,In_3323,In_4198);
and U2360 (N_2360,In_1399,In_1991);
and U2361 (N_2361,In_4823,In_1624);
and U2362 (N_2362,In_4392,In_214);
or U2363 (N_2363,In_2902,In_231);
nand U2364 (N_2364,In_2884,In_4161);
or U2365 (N_2365,In_1519,In_4197);
nor U2366 (N_2366,In_4342,In_776);
nor U2367 (N_2367,In_1826,In_3287);
nand U2368 (N_2368,In_3554,In_631);
xnor U2369 (N_2369,In_161,In_2952);
nand U2370 (N_2370,In_641,In_4402);
nand U2371 (N_2371,In_3487,In_2876);
or U2372 (N_2372,In_1147,In_1683);
or U2373 (N_2373,In_1458,In_2224);
or U2374 (N_2374,In_1601,In_1198);
or U2375 (N_2375,In_4025,In_3311);
nand U2376 (N_2376,In_2445,In_1444);
and U2377 (N_2377,In_436,In_3781);
xor U2378 (N_2378,In_1447,In_3368);
nand U2379 (N_2379,In_4580,In_1295);
and U2380 (N_2380,In_4828,In_1423);
and U2381 (N_2381,In_2217,In_133);
xnor U2382 (N_2382,In_2284,In_3604);
nand U2383 (N_2383,In_4687,In_1212);
nand U2384 (N_2384,In_3832,In_4093);
or U2385 (N_2385,In_39,In_4330);
and U2386 (N_2386,In_4199,In_2145);
nor U2387 (N_2387,In_1064,In_2272);
xnor U2388 (N_2388,In_2618,In_1049);
and U2389 (N_2389,In_2851,In_1101);
nor U2390 (N_2390,In_4566,In_2000);
xnor U2391 (N_2391,In_2333,In_824);
and U2392 (N_2392,In_1836,In_4503);
nand U2393 (N_2393,In_4280,In_2497);
or U2394 (N_2394,In_1215,In_1988);
or U2395 (N_2395,In_3098,In_62);
and U2396 (N_2396,In_2521,In_4658);
or U2397 (N_2397,In_2777,In_3742);
and U2398 (N_2398,In_2344,In_1946);
or U2399 (N_2399,In_4945,In_3244);
nor U2400 (N_2400,In_4807,In_953);
nor U2401 (N_2401,In_2206,In_3432);
nand U2402 (N_2402,In_2245,In_4408);
nand U2403 (N_2403,In_2386,In_783);
nor U2404 (N_2404,In_368,In_2702);
xor U2405 (N_2405,In_3025,In_513);
nor U2406 (N_2406,In_4871,In_3746);
and U2407 (N_2407,In_1711,In_4424);
xnor U2408 (N_2408,In_276,In_3579);
and U2409 (N_2409,In_742,In_99);
nor U2410 (N_2410,In_229,In_3561);
and U2411 (N_2411,In_3682,In_4683);
nor U2412 (N_2412,In_1844,In_2767);
nor U2413 (N_2413,In_2617,In_995);
xor U2414 (N_2414,In_2862,In_1206);
nor U2415 (N_2415,In_4551,In_2427);
xnor U2416 (N_2416,In_1607,In_1567);
or U2417 (N_2417,In_680,In_125);
nor U2418 (N_2418,In_3985,In_2032);
and U2419 (N_2419,In_511,In_2964);
nor U2420 (N_2420,In_1801,In_1702);
nand U2421 (N_2421,In_1261,In_2886);
nor U2422 (N_2422,In_4128,In_1518);
nand U2423 (N_2423,In_82,In_4416);
nand U2424 (N_2424,In_2659,In_361);
or U2425 (N_2425,In_3151,In_2809);
nor U2426 (N_2426,In_2830,In_4788);
xnor U2427 (N_2427,In_713,In_3077);
xnor U2428 (N_2428,In_4496,In_1907);
or U2429 (N_2429,In_520,In_4266);
nand U2430 (N_2430,In_4540,In_135);
xor U2431 (N_2431,In_1139,In_4935);
nor U2432 (N_2432,In_3690,In_1376);
nand U2433 (N_2433,In_2892,In_2343);
nand U2434 (N_2434,In_4305,In_2687);
or U2435 (N_2435,In_2984,In_1890);
nor U2436 (N_2436,In_4590,In_2324);
or U2437 (N_2437,In_2537,In_2483);
or U2438 (N_2438,In_3658,In_3628);
or U2439 (N_2439,In_341,In_1987);
or U2440 (N_2440,In_183,In_974);
nand U2441 (N_2441,In_2192,In_376);
or U2442 (N_2442,In_1883,In_2408);
xor U2443 (N_2443,In_1442,In_1819);
xnor U2444 (N_2444,In_4983,In_2339);
and U2445 (N_2445,In_2872,In_1670);
nand U2446 (N_2446,In_4293,In_4826);
or U2447 (N_2447,In_4802,In_1858);
xnor U2448 (N_2448,In_1491,In_3708);
nor U2449 (N_2449,In_1368,In_3564);
nand U2450 (N_2450,In_3953,In_726);
nor U2451 (N_2451,In_5,In_2768);
nor U2452 (N_2452,In_2509,In_3802);
nor U2453 (N_2453,In_4009,In_832);
nand U2454 (N_2454,In_1745,In_811);
xor U2455 (N_2455,In_2612,In_4840);
xnor U2456 (N_2456,In_2153,In_2162);
nor U2457 (N_2457,In_1133,In_3394);
or U2458 (N_2458,In_3320,In_2421);
xor U2459 (N_2459,In_1330,In_1132);
nor U2460 (N_2460,In_2226,In_1668);
or U2461 (N_2461,In_2852,In_3797);
and U2462 (N_2462,In_1743,In_2204);
and U2463 (N_2463,In_2215,In_3884);
xnor U2464 (N_2464,In_2985,In_2264);
and U2465 (N_2465,In_1403,In_3387);
nand U2466 (N_2466,In_1003,In_1531);
nand U2467 (N_2467,In_749,In_4905);
nor U2468 (N_2468,In_2271,In_3515);
nand U2469 (N_2469,In_3982,In_4588);
nor U2470 (N_2470,In_1980,In_1581);
nand U2471 (N_2471,In_1078,In_4970);
and U2472 (N_2472,In_884,In_3349);
and U2473 (N_2473,In_3249,In_380);
and U2474 (N_2474,In_2926,In_2552);
or U2475 (N_2475,In_2403,In_4892);
xnor U2476 (N_2476,In_821,In_1173);
nand U2477 (N_2477,In_2441,In_1540);
nand U2478 (N_2478,In_2327,In_1279);
and U2479 (N_2479,In_1180,In_2764);
and U2480 (N_2480,In_1739,In_377);
xnor U2481 (N_2481,In_2778,In_4584);
nand U2482 (N_2482,In_493,In_3261);
nand U2483 (N_2483,In_1508,In_1730);
and U2484 (N_2484,In_3240,In_1191);
nor U2485 (N_2485,In_699,In_2953);
or U2486 (N_2486,In_1744,In_4152);
or U2487 (N_2487,In_1165,In_839);
or U2488 (N_2488,In_2512,In_172);
and U2489 (N_2489,In_4317,In_4149);
xnor U2490 (N_2490,In_1809,In_415);
or U2491 (N_2491,In_152,In_3911);
xor U2492 (N_2492,In_1158,In_3803);
nor U2493 (N_2493,In_142,In_3967);
nand U2494 (N_2494,In_1169,In_3266);
nor U2495 (N_2495,In_4654,In_1408);
nor U2496 (N_2496,In_788,In_563);
xnor U2497 (N_2497,In_2049,In_3830);
and U2498 (N_2498,In_2366,In_1129);
or U2499 (N_2499,In_1036,In_1761);
and U2500 (N_2500,In_2852,In_2663);
xor U2501 (N_2501,In_1323,In_552);
xor U2502 (N_2502,In_3979,In_3942);
or U2503 (N_2503,In_2070,In_685);
nor U2504 (N_2504,In_3246,In_2556);
nor U2505 (N_2505,In_3834,In_2747);
nand U2506 (N_2506,In_1773,In_939);
nor U2507 (N_2507,In_4550,In_2457);
or U2508 (N_2508,In_1904,In_4667);
xnor U2509 (N_2509,In_3420,In_1475);
or U2510 (N_2510,In_3418,In_1415);
nor U2511 (N_2511,In_3784,In_1868);
nand U2512 (N_2512,In_4393,In_2946);
nand U2513 (N_2513,In_681,In_3296);
and U2514 (N_2514,In_4228,In_3927);
nand U2515 (N_2515,In_418,In_875);
nand U2516 (N_2516,In_4545,In_795);
and U2517 (N_2517,In_4626,In_4133);
xnor U2518 (N_2518,In_1713,In_408);
xnor U2519 (N_2519,In_1226,In_646);
nor U2520 (N_2520,In_2328,In_4721);
nor U2521 (N_2521,In_4101,In_1905);
xor U2522 (N_2522,In_784,In_2257);
xnor U2523 (N_2523,In_620,In_278);
nand U2524 (N_2524,In_4369,In_1536);
nand U2525 (N_2525,In_1868,In_505);
nor U2526 (N_2526,In_1905,In_2898);
nor U2527 (N_2527,In_371,In_2949);
nand U2528 (N_2528,In_2546,In_691);
nand U2529 (N_2529,In_57,In_2636);
or U2530 (N_2530,In_137,In_1526);
nor U2531 (N_2531,In_2701,In_381);
nand U2532 (N_2532,In_1660,In_2765);
or U2533 (N_2533,In_1261,In_1893);
nor U2534 (N_2534,In_1247,In_1181);
and U2535 (N_2535,In_440,In_680);
or U2536 (N_2536,In_2845,In_3107);
and U2537 (N_2537,In_4776,In_1137);
nor U2538 (N_2538,In_2413,In_4459);
or U2539 (N_2539,In_3772,In_4819);
xor U2540 (N_2540,In_816,In_391);
nor U2541 (N_2541,In_929,In_2802);
xnor U2542 (N_2542,In_237,In_113);
and U2543 (N_2543,In_3733,In_4517);
or U2544 (N_2544,In_3374,In_312);
and U2545 (N_2545,In_1453,In_3278);
and U2546 (N_2546,In_3952,In_3542);
or U2547 (N_2547,In_597,In_3093);
nor U2548 (N_2548,In_865,In_3287);
nand U2549 (N_2549,In_516,In_3765);
and U2550 (N_2550,In_487,In_2015);
and U2551 (N_2551,In_4978,In_4800);
and U2552 (N_2552,In_310,In_1456);
nor U2553 (N_2553,In_459,In_2798);
and U2554 (N_2554,In_4353,In_1448);
nor U2555 (N_2555,In_4490,In_3092);
nand U2556 (N_2556,In_4286,In_3884);
nand U2557 (N_2557,In_3036,In_438);
xor U2558 (N_2558,In_2047,In_2756);
nor U2559 (N_2559,In_1724,In_517);
xnor U2560 (N_2560,In_1130,In_3402);
nor U2561 (N_2561,In_3254,In_4856);
nor U2562 (N_2562,In_3611,In_2670);
nor U2563 (N_2563,In_908,In_4312);
nor U2564 (N_2564,In_3687,In_2726);
or U2565 (N_2565,In_4730,In_1063);
xnor U2566 (N_2566,In_3097,In_4018);
nand U2567 (N_2567,In_4554,In_3610);
xnor U2568 (N_2568,In_1858,In_2406);
or U2569 (N_2569,In_780,In_3870);
nor U2570 (N_2570,In_1470,In_2132);
xor U2571 (N_2571,In_4977,In_3036);
or U2572 (N_2572,In_19,In_3443);
or U2573 (N_2573,In_3018,In_3318);
xor U2574 (N_2574,In_3217,In_3049);
or U2575 (N_2575,In_4809,In_4240);
nand U2576 (N_2576,In_159,In_3455);
xor U2577 (N_2577,In_507,In_1527);
nor U2578 (N_2578,In_2398,In_4163);
and U2579 (N_2579,In_3372,In_4160);
and U2580 (N_2580,In_3770,In_137);
or U2581 (N_2581,In_1084,In_2633);
and U2582 (N_2582,In_556,In_4004);
and U2583 (N_2583,In_276,In_1633);
xor U2584 (N_2584,In_975,In_1244);
or U2585 (N_2585,In_1460,In_4405);
nor U2586 (N_2586,In_3658,In_3058);
xnor U2587 (N_2587,In_729,In_3654);
xnor U2588 (N_2588,In_3474,In_1111);
nand U2589 (N_2589,In_4320,In_3502);
nor U2590 (N_2590,In_3192,In_587);
nand U2591 (N_2591,In_1698,In_4531);
nand U2592 (N_2592,In_2519,In_353);
or U2593 (N_2593,In_3156,In_247);
xnor U2594 (N_2594,In_546,In_1823);
or U2595 (N_2595,In_4927,In_590);
nand U2596 (N_2596,In_1090,In_4714);
xnor U2597 (N_2597,In_3015,In_1051);
and U2598 (N_2598,In_4296,In_4555);
or U2599 (N_2599,In_4369,In_2295);
nand U2600 (N_2600,In_3949,In_908);
or U2601 (N_2601,In_1453,In_4576);
nand U2602 (N_2602,In_975,In_3025);
xnor U2603 (N_2603,In_3611,In_4235);
xor U2604 (N_2604,In_2558,In_425);
nand U2605 (N_2605,In_2521,In_683);
or U2606 (N_2606,In_2881,In_1022);
or U2607 (N_2607,In_1213,In_4174);
nor U2608 (N_2608,In_1599,In_2686);
or U2609 (N_2609,In_1195,In_4701);
nand U2610 (N_2610,In_2373,In_2931);
and U2611 (N_2611,In_2257,In_2985);
or U2612 (N_2612,In_87,In_536);
xnor U2613 (N_2613,In_2072,In_1381);
nor U2614 (N_2614,In_4551,In_4501);
nand U2615 (N_2615,In_3935,In_3749);
and U2616 (N_2616,In_603,In_4587);
or U2617 (N_2617,In_2186,In_3219);
and U2618 (N_2618,In_2450,In_4902);
nor U2619 (N_2619,In_403,In_4911);
and U2620 (N_2620,In_1162,In_3631);
and U2621 (N_2621,In_1402,In_1651);
nor U2622 (N_2622,In_411,In_2054);
xor U2623 (N_2623,In_4865,In_4149);
or U2624 (N_2624,In_1347,In_401);
or U2625 (N_2625,In_644,In_2333);
nor U2626 (N_2626,In_2220,In_4690);
xor U2627 (N_2627,In_2789,In_3428);
nand U2628 (N_2628,In_476,In_479);
and U2629 (N_2629,In_2343,In_3815);
and U2630 (N_2630,In_837,In_1544);
and U2631 (N_2631,In_4271,In_3623);
nor U2632 (N_2632,In_4503,In_911);
nand U2633 (N_2633,In_4926,In_1568);
xor U2634 (N_2634,In_659,In_2939);
nor U2635 (N_2635,In_2901,In_3080);
xnor U2636 (N_2636,In_2332,In_3716);
nor U2637 (N_2637,In_1834,In_812);
nor U2638 (N_2638,In_2952,In_2830);
or U2639 (N_2639,In_1677,In_4592);
and U2640 (N_2640,In_952,In_1369);
or U2641 (N_2641,In_1417,In_1845);
xnor U2642 (N_2642,In_4422,In_1271);
and U2643 (N_2643,In_4861,In_5);
nor U2644 (N_2644,In_2644,In_822);
or U2645 (N_2645,In_3235,In_1886);
nand U2646 (N_2646,In_2002,In_2643);
nor U2647 (N_2647,In_2333,In_133);
xnor U2648 (N_2648,In_547,In_4740);
nand U2649 (N_2649,In_4746,In_470);
and U2650 (N_2650,In_4216,In_3430);
nand U2651 (N_2651,In_3074,In_1222);
nand U2652 (N_2652,In_1129,In_2380);
nor U2653 (N_2653,In_1114,In_3769);
nand U2654 (N_2654,In_4724,In_2139);
and U2655 (N_2655,In_172,In_4816);
nor U2656 (N_2656,In_1618,In_4750);
nor U2657 (N_2657,In_161,In_669);
xor U2658 (N_2658,In_2879,In_3994);
nor U2659 (N_2659,In_3895,In_2242);
nand U2660 (N_2660,In_4351,In_4836);
or U2661 (N_2661,In_638,In_403);
nand U2662 (N_2662,In_357,In_1671);
and U2663 (N_2663,In_4626,In_366);
nand U2664 (N_2664,In_3915,In_139);
or U2665 (N_2665,In_4844,In_532);
nor U2666 (N_2666,In_4751,In_4133);
or U2667 (N_2667,In_3464,In_4227);
or U2668 (N_2668,In_2495,In_4948);
or U2669 (N_2669,In_493,In_3379);
nor U2670 (N_2670,In_2858,In_1225);
nor U2671 (N_2671,In_3430,In_2274);
nand U2672 (N_2672,In_2733,In_2889);
and U2673 (N_2673,In_2044,In_2943);
nor U2674 (N_2674,In_2093,In_915);
nor U2675 (N_2675,In_4068,In_426);
nand U2676 (N_2676,In_3414,In_745);
nor U2677 (N_2677,In_633,In_4156);
or U2678 (N_2678,In_3289,In_3605);
nand U2679 (N_2679,In_3442,In_1395);
nand U2680 (N_2680,In_2960,In_1269);
and U2681 (N_2681,In_4611,In_3525);
and U2682 (N_2682,In_1719,In_556);
and U2683 (N_2683,In_248,In_630);
or U2684 (N_2684,In_3569,In_4802);
or U2685 (N_2685,In_1496,In_2190);
and U2686 (N_2686,In_2010,In_591);
and U2687 (N_2687,In_1163,In_1785);
or U2688 (N_2688,In_1179,In_293);
or U2689 (N_2689,In_1879,In_1573);
nand U2690 (N_2690,In_4858,In_3696);
nand U2691 (N_2691,In_2974,In_1119);
nand U2692 (N_2692,In_342,In_4782);
nand U2693 (N_2693,In_904,In_2373);
or U2694 (N_2694,In_2170,In_1640);
nand U2695 (N_2695,In_4447,In_2006);
or U2696 (N_2696,In_1468,In_2817);
nand U2697 (N_2697,In_4355,In_811);
nor U2698 (N_2698,In_603,In_759);
and U2699 (N_2699,In_197,In_13);
xnor U2700 (N_2700,In_342,In_4490);
nand U2701 (N_2701,In_1449,In_1603);
nor U2702 (N_2702,In_871,In_1035);
nand U2703 (N_2703,In_4954,In_1574);
nand U2704 (N_2704,In_2789,In_4830);
and U2705 (N_2705,In_2202,In_1486);
and U2706 (N_2706,In_3099,In_3313);
xor U2707 (N_2707,In_1335,In_3103);
and U2708 (N_2708,In_1539,In_2319);
nand U2709 (N_2709,In_4917,In_3086);
nor U2710 (N_2710,In_2364,In_4121);
nor U2711 (N_2711,In_1214,In_626);
and U2712 (N_2712,In_3682,In_2535);
and U2713 (N_2713,In_1462,In_3946);
and U2714 (N_2714,In_2339,In_1220);
or U2715 (N_2715,In_2953,In_1742);
nand U2716 (N_2716,In_1558,In_1368);
and U2717 (N_2717,In_102,In_939);
nand U2718 (N_2718,In_1378,In_906);
and U2719 (N_2719,In_4275,In_3199);
nor U2720 (N_2720,In_3445,In_3757);
nor U2721 (N_2721,In_2819,In_2925);
xnor U2722 (N_2722,In_546,In_2003);
or U2723 (N_2723,In_3276,In_243);
xor U2724 (N_2724,In_1703,In_1155);
nand U2725 (N_2725,In_3456,In_4747);
nor U2726 (N_2726,In_633,In_4108);
xnor U2727 (N_2727,In_4443,In_439);
and U2728 (N_2728,In_1757,In_2077);
and U2729 (N_2729,In_831,In_1905);
or U2730 (N_2730,In_4212,In_2051);
nor U2731 (N_2731,In_1945,In_2633);
or U2732 (N_2732,In_73,In_935);
nand U2733 (N_2733,In_4831,In_4184);
nand U2734 (N_2734,In_4111,In_1991);
and U2735 (N_2735,In_2378,In_329);
xnor U2736 (N_2736,In_3045,In_3715);
and U2737 (N_2737,In_1226,In_1427);
nor U2738 (N_2738,In_3237,In_1654);
or U2739 (N_2739,In_717,In_4881);
xnor U2740 (N_2740,In_103,In_1395);
nor U2741 (N_2741,In_4959,In_2361);
xnor U2742 (N_2742,In_740,In_4339);
and U2743 (N_2743,In_3780,In_274);
or U2744 (N_2744,In_1626,In_2267);
and U2745 (N_2745,In_3066,In_149);
and U2746 (N_2746,In_4946,In_3192);
nand U2747 (N_2747,In_1724,In_2443);
and U2748 (N_2748,In_807,In_3655);
and U2749 (N_2749,In_1164,In_3938);
and U2750 (N_2750,In_3401,In_2692);
nor U2751 (N_2751,In_3222,In_178);
or U2752 (N_2752,In_4164,In_4251);
and U2753 (N_2753,In_1343,In_4126);
nor U2754 (N_2754,In_3054,In_3155);
nand U2755 (N_2755,In_544,In_2802);
nand U2756 (N_2756,In_1552,In_3864);
or U2757 (N_2757,In_2599,In_4414);
nand U2758 (N_2758,In_2738,In_1358);
or U2759 (N_2759,In_3868,In_2156);
xnor U2760 (N_2760,In_4343,In_2788);
or U2761 (N_2761,In_3931,In_4963);
or U2762 (N_2762,In_406,In_653);
xor U2763 (N_2763,In_4108,In_3558);
xor U2764 (N_2764,In_4539,In_4176);
or U2765 (N_2765,In_2890,In_1463);
nor U2766 (N_2766,In_2752,In_2480);
and U2767 (N_2767,In_397,In_3216);
or U2768 (N_2768,In_2011,In_2351);
xor U2769 (N_2769,In_2519,In_3951);
nor U2770 (N_2770,In_2296,In_4541);
nand U2771 (N_2771,In_734,In_1747);
and U2772 (N_2772,In_3965,In_4776);
xor U2773 (N_2773,In_624,In_3196);
or U2774 (N_2774,In_944,In_3607);
nand U2775 (N_2775,In_445,In_625);
and U2776 (N_2776,In_508,In_627);
or U2777 (N_2777,In_3812,In_4420);
and U2778 (N_2778,In_1427,In_4672);
or U2779 (N_2779,In_2380,In_681);
or U2780 (N_2780,In_3504,In_803);
and U2781 (N_2781,In_3782,In_2072);
nand U2782 (N_2782,In_3523,In_2323);
nand U2783 (N_2783,In_179,In_4481);
nand U2784 (N_2784,In_1873,In_3631);
or U2785 (N_2785,In_2320,In_1776);
or U2786 (N_2786,In_738,In_1663);
or U2787 (N_2787,In_4455,In_4123);
nor U2788 (N_2788,In_4884,In_3208);
nor U2789 (N_2789,In_14,In_4432);
and U2790 (N_2790,In_4369,In_2961);
or U2791 (N_2791,In_1292,In_4778);
and U2792 (N_2792,In_2275,In_3399);
and U2793 (N_2793,In_1007,In_510);
or U2794 (N_2794,In_4629,In_4245);
or U2795 (N_2795,In_2107,In_4233);
nor U2796 (N_2796,In_4269,In_1381);
and U2797 (N_2797,In_4505,In_4299);
nor U2798 (N_2798,In_4248,In_4595);
nor U2799 (N_2799,In_1425,In_3266);
or U2800 (N_2800,In_3373,In_4719);
or U2801 (N_2801,In_3069,In_2562);
nand U2802 (N_2802,In_250,In_4312);
or U2803 (N_2803,In_1919,In_1810);
nand U2804 (N_2804,In_2695,In_4272);
nand U2805 (N_2805,In_1750,In_2331);
and U2806 (N_2806,In_198,In_545);
or U2807 (N_2807,In_584,In_4273);
xnor U2808 (N_2808,In_3586,In_2192);
xor U2809 (N_2809,In_2748,In_2622);
xnor U2810 (N_2810,In_1861,In_3546);
nand U2811 (N_2811,In_1686,In_1667);
nor U2812 (N_2812,In_1707,In_3520);
and U2813 (N_2813,In_3086,In_635);
nand U2814 (N_2814,In_1968,In_4130);
xnor U2815 (N_2815,In_546,In_4527);
and U2816 (N_2816,In_977,In_970);
or U2817 (N_2817,In_4068,In_326);
nor U2818 (N_2818,In_169,In_2523);
and U2819 (N_2819,In_1225,In_3066);
or U2820 (N_2820,In_3918,In_4956);
nor U2821 (N_2821,In_3913,In_1409);
and U2822 (N_2822,In_3571,In_1548);
or U2823 (N_2823,In_2511,In_631);
nor U2824 (N_2824,In_3621,In_2183);
and U2825 (N_2825,In_2753,In_3605);
and U2826 (N_2826,In_2463,In_4960);
xor U2827 (N_2827,In_101,In_1601);
or U2828 (N_2828,In_400,In_1604);
or U2829 (N_2829,In_1750,In_893);
and U2830 (N_2830,In_4391,In_3342);
xor U2831 (N_2831,In_1214,In_2793);
and U2832 (N_2832,In_3474,In_156);
nand U2833 (N_2833,In_2944,In_4406);
or U2834 (N_2834,In_212,In_610);
nor U2835 (N_2835,In_26,In_1680);
nand U2836 (N_2836,In_2866,In_708);
nand U2837 (N_2837,In_3359,In_4129);
nor U2838 (N_2838,In_705,In_1591);
and U2839 (N_2839,In_1101,In_3017);
nand U2840 (N_2840,In_905,In_2188);
and U2841 (N_2841,In_3343,In_4129);
xnor U2842 (N_2842,In_1482,In_260);
nand U2843 (N_2843,In_4049,In_3386);
nor U2844 (N_2844,In_4091,In_2772);
nor U2845 (N_2845,In_4192,In_2617);
or U2846 (N_2846,In_3327,In_4799);
nor U2847 (N_2847,In_598,In_1197);
and U2848 (N_2848,In_4597,In_312);
or U2849 (N_2849,In_3415,In_2081);
nor U2850 (N_2850,In_4597,In_3783);
nand U2851 (N_2851,In_2922,In_2054);
nand U2852 (N_2852,In_1349,In_3782);
and U2853 (N_2853,In_2830,In_2918);
nand U2854 (N_2854,In_4985,In_2188);
or U2855 (N_2855,In_76,In_3874);
nor U2856 (N_2856,In_1620,In_1281);
or U2857 (N_2857,In_3358,In_1869);
nand U2858 (N_2858,In_3152,In_3926);
or U2859 (N_2859,In_863,In_1190);
nand U2860 (N_2860,In_3560,In_1361);
nand U2861 (N_2861,In_3786,In_1638);
nand U2862 (N_2862,In_640,In_535);
nor U2863 (N_2863,In_2126,In_4599);
xnor U2864 (N_2864,In_350,In_1043);
or U2865 (N_2865,In_1966,In_4425);
nor U2866 (N_2866,In_4091,In_2034);
or U2867 (N_2867,In_1517,In_4329);
or U2868 (N_2868,In_1138,In_4160);
or U2869 (N_2869,In_2005,In_598);
xnor U2870 (N_2870,In_3066,In_2351);
or U2871 (N_2871,In_922,In_2032);
nand U2872 (N_2872,In_4694,In_779);
xor U2873 (N_2873,In_137,In_302);
or U2874 (N_2874,In_3115,In_640);
xor U2875 (N_2875,In_1634,In_3171);
and U2876 (N_2876,In_2400,In_4039);
and U2877 (N_2877,In_3073,In_806);
or U2878 (N_2878,In_1251,In_209);
nand U2879 (N_2879,In_2461,In_2121);
xor U2880 (N_2880,In_1346,In_3319);
nor U2881 (N_2881,In_2928,In_1019);
or U2882 (N_2882,In_274,In_4673);
and U2883 (N_2883,In_270,In_2715);
xnor U2884 (N_2884,In_2312,In_3185);
nand U2885 (N_2885,In_4820,In_1057);
nand U2886 (N_2886,In_980,In_787);
xor U2887 (N_2887,In_754,In_1455);
nor U2888 (N_2888,In_1184,In_2530);
nand U2889 (N_2889,In_127,In_3259);
nand U2890 (N_2890,In_2307,In_4913);
or U2891 (N_2891,In_1109,In_3837);
and U2892 (N_2892,In_2811,In_1276);
xor U2893 (N_2893,In_4276,In_1152);
and U2894 (N_2894,In_4705,In_2592);
or U2895 (N_2895,In_3673,In_2662);
nor U2896 (N_2896,In_3767,In_962);
nand U2897 (N_2897,In_4590,In_1809);
nor U2898 (N_2898,In_4308,In_3697);
or U2899 (N_2899,In_3592,In_3122);
and U2900 (N_2900,In_814,In_1612);
and U2901 (N_2901,In_2233,In_4295);
xor U2902 (N_2902,In_4052,In_212);
xnor U2903 (N_2903,In_3763,In_2315);
nand U2904 (N_2904,In_437,In_2629);
nand U2905 (N_2905,In_3545,In_1114);
xor U2906 (N_2906,In_1253,In_4177);
xnor U2907 (N_2907,In_4844,In_3087);
or U2908 (N_2908,In_482,In_2788);
xnor U2909 (N_2909,In_1488,In_2184);
nand U2910 (N_2910,In_2619,In_3409);
nor U2911 (N_2911,In_4926,In_3963);
and U2912 (N_2912,In_1419,In_4296);
and U2913 (N_2913,In_2312,In_1898);
or U2914 (N_2914,In_2883,In_3513);
and U2915 (N_2915,In_4875,In_1239);
or U2916 (N_2916,In_3034,In_2007);
nor U2917 (N_2917,In_1980,In_1066);
and U2918 (N_2918,In_1573,In_528);
nor U2919 (N_2919,In_3549,In_1112);
and U2920 (N_2920,In_2861,In_4832);
xnor U2921 (N_2921,In_2729,In_124);
nor U2922 (N_2922,In_3667,In_143);
nor U2923 (N_2923,In_278,In_1142);
xnor U2924 (N_2924,In_862,In_4466);
or U2925 (N_2925,In_1304,In_1052);
or U2926 (N_2926,In_2161,In_3304);
nand U2927 (N_2927,In_3423,In_524);
xor U2928 (N_2928,In_4212,In_1017);
or U2929 (N_2929,In_2141,In_43);
nand U2930 (N_2930,In_3436,In_318);
or U2931 (N_2931,In_4030,In_1933);
or U2932 (N_2932,In_3622,In_3711);
nor U2933 (N_2933,In_2170,In_505);
or U2934 (N_2934,In_1471,In_3538);
nand U2935 (N_2935,In_3769,In_561);
nand U2936 (N_2936,In_75,In_2721);
and U2937 (N_2937,In_4968,In_3219);
nor U2938 (N_2938,In_4736,In_977);
nor U2939 (N_2939,In_3313,In_3454);
nand U2940 (N_2940,In_3535,In_58);
nor U2941 (N_2941,In_537,In_4507);
nand U2942 (N_2942,In_235,In_2164);
or U2943 (N_2943,In_4042,In_2842);
nor U2944 (N_2944,In_4774,In_2656);
nor U2945 (N_2945,In_2483,In_4510);
nor U2946 (N_2946,In_3275,In_522);
and U2947 (N_2947,In_326,In_3434);
and U2948 (N_2948,In_4901,In_2949);
nand U2949 (N_2949,In_4218,In_2325);
or U2950 (N_2950,In_2,In_4707);
nand U2951 (N_2951,In_1077,In_4533);
xor U2952 (N_2952,In_2696,In_438);
nor U2953 (N_2953,In_1567,In_4011);
nor U2954 (N_2954,In_366,In_1401);
xor U2955 (N_2955,In_1808,In_2087);
and U2956 (N_2956,In_2402,In_690);
nand U2957 (N_2957,In_4809,In_1629);
and U2958 (N_2958,In_3431,In_3404);
nor U2959 (N_2959,In_640,In_4244);
or U2960 (N_2960,In_1880,In_2950);
and U2961 (N_2961,In_387,In_2343);
xnor U2962 (N_2962,In_3359,In_4047);
or U2963 (N_2963,In_2567,In_2765);
and U2964 (N_2964,In_3789,In_2955);
nor U2965 (N_2965,In_3695,In_4167);
or U2966 (N_2966,In_1879,In_4231);
or U2967 (N_2967,In_2989,In_87);
xnor U2968 (N_2968,In_2440,In_760);
nand U2969 (N_2969,In_4436,In_1949);
xor U2970 (N_2970,In_2001,In_4768);
nor U2971 (N_2971,In_2324,In_1306);
nand U2972 (N_2972,In_688,In_4425);
nand U2973 (N_2973,In_2365,In_3252);
nand U2974 (N_2974,In_811,In_1237);
nor U2975 (N_2975,In_383,In_2274);
and U2976 (N_2976,In_1383,In_1423);
and U2977 (N_2977,In_2119,In_2046);
or U2978 (N_2978,In_4039,In_2476);
and U2979 (N_2979,In_4304,In_4441);
or U2980 (N_2980,In_4522,In_4730);
and U2981 (N_2981,In_1272,In_117);
or U2982 (N_2982,In_3148,In_4706);
and U2983 (N_2983,In_2462,In_1858);
and U2984 (N_2984,In_1824,In_981);
nor U2985 (N_2985,In_4297,In_4778);
or U2986 (N_2986,In_560,In_3946);
nor U2987 (N_2987,In_797,In_2207);
nor U2988 (N_2988,In_709,In_1233);
xnor U2989 (N_2989,In_581,In_2610);
and U2990 (N_2990,In_1620,In_1894);
and U2991 (N_2991,In_2048,In_4304);
xnor U2992 (N_2992,In_35,In_4795);
and U2993 (N_2993,In_1333,In_1218);
and U2994 (N_2994,In_3908,In_2687);
or U2995 (N_2995,In_3952,In_1984);
xor U2996 (N_2996,In_625,In_1494);
nor U2997 (N_2997,In_420,In_938);
xor U2998 (N_2998,In_3308,In_1737);
and U2999 (N_2999,In_4213,In_1584);
xnor U3000 (N_3000,In_4765,In_1219);
nand U3001 (N_3001,In_2198,In_545);
xor U3002 (N_3002,In_3879,In_2435);
and U3003 (N_3003,In_2542,In_304);
nor U3004 (N_3004,In_2717,In_2723);
xor U3005 (N_3005,In_1083,In_1383);
nand U3006 (N_3006,In_1005,In_4723);
and U3007 (N_3007,In_4180,In_4124);
xnor U3008 (N_3008,In_264,In_600);
nor U3009 (N_3009,In_3147,In_4044);
or U3010 (N_3010,In_1497,In_2021);
nor U3011 (N_3011,In_1232,In_291);
or U3012 (N_3012,In_725,In_4907);
nand U3013 (N_3013,In_2346,In_1798);
or U3014 (N_3014,In_4331,In_3196);
nand U3015 (N_3015,In_2112,In_3582);
or U3016 (N_3016,In_3057,In_4377);
nand U3017 (N_3017,In_2045,In_4519);
or U3018 (N_3018,In_3727,In_681);
and U3019 (N_3019,In_3231,In_2496);
and U3020 (N_3020,In_831,In_1023);
or U3021 (N_3021,In_550,In_1426);
nand U3022 (N_3022,In_1605,In_508);
nor U3023 (N_3023,In_202,In_499);
and U3024 (N_3024,In_57,In_2649);
or U3025 (N_3025,In_620,In_2627);
or U3026 (N_3026,In_4589,In_253);
nor U3027 (N_3027,In_1090,In_2136);
and U3028 (N_3028,In_4073,In_2366);
nor U3029 (N_3029,In_40,In_4816);
xor U3030 (N_3030,In_3431,In_568);
xnor U3031 (N_3031,In_243,In_163);
nand U3032 (N_3032,In_1327,In_1690);
or U3033 (N_3033,In_1972,In_1502);
nor U3034 (N_3034,In_1185,In_1741);
or U3035 (N_3035,In_158,In_1231);
nor U3036 (N_3036,In_3144,In_3725);
xnor U3037 (N_3037,In_893,In_3703);
xor U3038 (N_3038,In_1028,In_571);
or U3039 (N_3039,In_298,In_2078);
and U3040 (N_3040,In_3884,In_4986);
xor U3041 (N_3041,In_4910,In_1265);
nand U3042 (N_3042,In_1060,In_1072);
or U3043 (N_3043,In_1974,In_253);
xor U3044 (N_3044,In_1498,In_16);
and U3045 (N_3045,In_1578,In_3208);
and U3046 (N_3046,In_2111,In_1284);
nand U3047 (N_3047,In_117,In_1561);
or U3048 (N_3048,In_2114,In_4067);
or U3049 (N_3049,In_1091,In_167);
or U3050 (N_3050,In_416,In_1745);
nor U3051 (N_3051,In_2694,In_3658);
and U3052 (N_3052,In_3387,In_1751);
nor U3053 (N_3053,In_1166,In_759);
nor U3054 (N_3054,In_4519,In_3342);
xor U3055 (N_3055,In_769,In_2752);
or U3056 (N_3056,In_3337,In_4116);
xor U3057 (N_3057,In_3895,In_2592);
nor U3058 (N_3058,In_310,In_714);
or U3059 (N_3059,In_4687,In_1634);
or U3060 (N_3060,In_4103,In_693);
or U3061 (N_3061,In_415,In_4861);
nand U3062 (N_3062,In_4434,In_789);
nor U3063 (N_3063,In_4408,In_2338);
nand U3064 (N_3064,In_2096,In_3766);
nor U3065 (N_3065,In_869,In_4570);
nand U3066 (N_3066,In_4994,In_745);
nand U3067 (N_3067,In_4860,In_3459);
and U3068 (N_3068,In_2580,In_1047);
nor U3069 (N_3069,In_3099,In_4331);
nor U3070 (N_3070,In_229,In_3748);
or U3071 (N_3071,In_2619,In_1225);
or U3072 (N_3072,In_3991,In_106);
and U3073 (N_3073,In_4578,In_4407);
or U3074 (N_3074,In_2339,In_2926);
nor U3075 (N_3075,In_4997,In_3457);
nand U3076 (N_3076,In_684,In_4760);
or U3077 (N_3077,In_3095,In_3140);
xnor U3078 (N_3078,In_3672,In_673);
nor U3079 (N_3079,In_2487,In_1055);
and U3080 (N_3080,In_4500,In_4847);
nor U3081 (N_3081,In_3559,In_2303);
xnor U3082 (N_3082,In_3689,In_1058);
or U3083 (N_3083,In_3032,In_1758);
and U3084 (N_3084,In_3209,In_2710);
nand U3085 (N_3085,In_4183,In_3459);
or U3086 (N_3086,In_1723,In_1939);
xnor U3087 (N_3087,In_1297,In_3078);
and U3088 (N_3088,In_4039,In_504);
and U3089 (N_3089,In_2183,In_603);
nor U3090 (N_3090,In_2992,In_81);
xor U3091 (N_3091,In_3884,In_852);
nor U3092 (N_3092,In_1388,In_2154);
or U3093 (N_3093,In_2006,In_421);
and U3094 (N_3094,In_1165,In_2945);
and U3095 (N_3095,In_1456,In_3879);
or U3096 (N_3096,In_703,In_443);
and U3097 (N_3097,In_1595,In_2912);
nor U3098 (N_3098,In_3933,In_3870);
xnor U3099 (N_3099,In_2430,In_1205);
nor U3100 (N_3100,In_1533,In_1030);
nand U3101 (N_3101,In_52,In_709);
and U3102 (N_3102,In_2824,In_537);
and U3103 (N_3103,In_4852,In_676);
nor U3104 (N_3104,In_3528,In_624);
nor U3105 (N_3105,In_651,In_1580);
nand U3106 (N_3106,In_3685,In_1231);
xor U3107 (N_3107,In_875,In_4720);
or U3108 (N_3108,In_4283,In_2238);
nor U3109 (N_3109,In_1929,In_2424);
or U3110 (N_3110,In_1719,In_2872);
or U3111 (N_3111,In_139,In_1387);
nor U3112 (N_3112,In_26,In_3553);
and U3113 (N_3113,In_2715,In_329);
or U3114 (N_3114,In_2910,In_4693);
xor U3115 (N_3115,In_1097,In_4692);
nand U3116 (N_3116,In_715,In_4777);
nand U3117 (N_3117,In_3451,In_1423);
nor U3118 (N_3118,In_4325,In_4767);
nand U3119 (N_3119,In_4905,In_1099);
nor U3120 (N_3120,In_691,In_1239);
nor U3121 (N_3121,In_1616,In_111);
nor U3122 (N_3122,In_4149,In_248);
and U3123 (N_3123,In_2607,In_3003);
xnor U3124 (N_3124,In_2269,In_1912);
nand U3125 (N_3125,In_3325,In_2957);
nand U3126 (N_3126,In_1359,In_1279);
nor U3127 (N_3127,In_4680,In_49);
or U3128 (N_3128,In_2574,In_2439);
and U3129 (N_3129,In_2319,In_697);
and U3130 (N_3130,In_4949,In_4098);
xor U3131 (N_3131,In_883,In_1171);
nor U3132 (N_3132,In_3500,In_4615);
nand U3133 (N_3133,In_1639,In_3460);
nand U3134 (N_3134,In_4623,In_1447);
xor U3135 (N_3135,In_1316,In_3107);
xnor U3136 (N_3136,In_3504,In_2848);
or U3137 (N_3137,In_1754,In_3108);
xor U3138 (N_3138,In_1838,In_285);
and U3139 (N_3139,In_3681,In_4210);
and U3140 (N_3140,In_2756,In_352);
nand U3141 (N_3141,In_2965,In_1846);
nor U3142 (N_3142,In_1570,In_1616);
and U3143 (N_3143,In_252,In_575);
xor U3144 (N_3144,In_555,In_2121);
nand U3145 (N_3145,In_960,In_877);
nor U3146 (N_3146,In_1352,In_181);
xnor U3147 (N_3147,In_1960,In_1096);
nand U3148 (N_3148,In_3877,In_4517);
xnor U3149 (N_3149,In_1630,In_1865);
nor U3150 (N_3150,In_2284,In_3075);
and U3151 (N_3151,In_4507,In_2066);
and U3152 (N_3152,In_4124,In_1914);
xor U3153 (N_3153,In_3416,In_588);
nor U3154 (N_3154,In_4034,In_3469);
or U3155 (N_3155,In_722,In_4756);
or U3156 (N_3156,In_3941,In_871);
and U3157 (N_3157,In_1689,In_3940);
and U3158 (N_3158,In_908,In_2267);
or U3159 (N_3159,In_2640,In_615);
or U3160 (N_3160,In_1685,In_3214);
and U3161 (N_3161,In_28,In_3393);
and U3162 (N_3162,In_3203,In_1437);
and U3163 (N_3163,In_4830,In_1440);
nand U3164 (N_3164,In_4857,In_2867);
xor U3165 (N_3165,In_4886,In_2543);
nand U3166 (N_3166,In_540,In_1644);
and U3167 (N_3167,In_3728,In_4783);
xnor U3168 (N_3168,In_3924,In_1986);
nand U3169 (N_3169,In_2629,In_4798);
nand U3170 (N_3170,In_2064,In_1598);
nor U3171 (N_3171,In_2726,In_1492);
or U3172 (N_3172,In_1909,In_4185);
nor U3173 (N_3173,In_4266,In_2209);
xnor U3174 (N_3174,In_4721,In_4572);
xnor U3175 (N_3175,In_3714,In_1750);
and U3176 (N_3176,In_3551,In_135);
or U3177 (N_3177,In_2333,In_1246);
xor U3178 (N_3178,In_272,In_4862);
nand U3179 (N_3179,In_150,In_2766);
or U3180 (N_3180,In_2470,In_3526);
nor U3181 (N_3181,In_4414,In_1627);
and U3182 (N_3182,In_3631,In_4823);
nand U3183 (N_3183,In_3249,In_4156);
and U3184 (N_3184,In_4940,In_327);
nor U3185 (N_3185,In_1059,In_3454);
and U3186 (N_3186,In_2317,In_389);
nand U3187 (N_3187,In_1027,In_2889);
nand U3188 (N_3188,In_3881,In_1837);
or U3189 (N_3189,In_4297,In_4308);
nand U3190 (N_3190,In_825,In_1635);
or U3191 (N_3191,In_2092,In_461);
xor U3192 (N_3192,In_2678,In_3057);
or U3193 (N_3193,In_1821,In_2369);
and U3194 (N_3194,In_374,In_4474);
or U3195 (N_3195,In_2984,In_152);
and U3196 (N_3196,In_2232,In_2421);
nand U3197 (N_3197,In_4357,In_667);
and U3198 (N_3198,In_1728,In_2654);
xnor U3199 (N_3199,In_2189,In_3091);
and U3200 (N_3200,In_2148,In_3956);
or U3201 (N_3201,In_841,In_3989);
xor U3202 (N_3202,In_2363,In_4204);
or U3203 (N_3203,In_4985,In_1379);
nor U3204 (N_3204,In_1854,In_958);
or U3205 (N_3205,In_2443,In_2154);
nand U3206 (N_3206,In_3283,In_180);
nor U3207 (N_3207,In_2119,In_4051);
and U3208 (N_3208,In_4336,In_3038);
nor U3209 (N_3209,In_3902,In_2583);
and U3210 (N_3210,In_2234,In_898);
nand U3211 (N_3211,In_68,In_4957);
or U3212 (N_3212,In_3193,In_4973);
nand U3213 (N_3213,In_4345,In_4379);
nand U3214 (N_3214,In_1374,In_1066);
and U3215 (N_3215,In_2416,In_4755);
and U3216 (N_3216,In_3863,In_4756);
nor U3217 (N_3217,In_2732,In_3356);
xnor U3218 (N_3218,In_1917,In_1934);
or U3219 (N_3219,In_2545,In_1493);
and U3220 (N_3220,In_4196,In_2785);
nor U3221 (N_3221,In_3408,In_2069);
nor U3222 (N_3222,In_3724,In_1527);
nand U3223 (N_3223,In_1466,In_2196);
nand U3224 (N_3224,In_2140,In_3832);
nor U3225 (N_3225,In_1861,In_2442);
xor U3226 (N_3226,In_2395,In_4816);
xnor U3227 (N_3227,In_4596,In_3428);
nor U3228 (N_3228,In_825,In_2395);
nor U3229 (N_3229,In_1847,In_2135);
or U3230 (N_3230,In_3463,In_3369);
and U3231 (N_3231,In_1410,In_4785);
xor U3232 (N_3232,In_1830,In_4479);
and U3233 (N_3233,In_3452,In_291);
and U3234 (N_3234,In_3719,In_1021);
or U3235 (N_3235,In_4737,In_1595);
and U3236 (N_3236,In_3764,In_2472);
and U3237 (N_3237,In_3719,In_4521);
or U3238 (N_3238,In_168,In_337);
nor U3239 (N_3239,In_773,In_2335);
xnor U3240 (N_3240,In_359,In_3257);
and U3241 (N_3241,In_1225,In_275);
nor U3242 (N_3242,In_1354,In_1265);
nand U3243 (N_3243,In_3528,In_168);
or U3244 (N_3244,In_3017,In_3347);
xor U3245 (N_3245,In_1058,In_1406);
or U3246 (N_3246,In_4190,In_3789);
xnor U3247 (N_3247,In_4259,In_4609);
xnor U3248 (N_3248,In_1087,In_4440);
nand U3249 (N_3249,In_1302,In_3320);
and U3250 (N_3250,In_2485,In_973);
nand U3251 (N_3251,In_420,In_4216);
and U3252 (N_3252,In_791,In_4356);
nand U3253 (N_3253,In_3855,In_1026);
nor U3254 (N_3254,In_1195,In_3752);
xnor U3255 (N_3255,In_1133,In_2391);
and U3256 (N_3256,In_444,In_1975);
xor U3257 (N_3257,In_3276,In_411);
nand U3258 (N_3258,In_3424,In_413);
xnor U3259 (N_3259,In_322,In_325);
nand U3260 (N_3260,In_1470,In_1981);
nor U3261 (N_3261,In_1871,In_2266);
and U3262 (N_3262,In_3864,In_430);
nand U3263 (N_3263,In_3821,In_1218);
nand U3264 (N_3264,In_3932,In_1563);
and U3265 (N_3265,In_897,In_1313);
nor U3266 (N_3266,In_1517,In_2100);
nand U3267 (N_3267,In_1706,In_2415);
nor U3268 (N_3268,In_4027,In_3029);
or U3269 (N_3269,In_1651,In_3288);
nand U3270 (N_3270,In_3627,In_4600);
nand U3271 (N_3271,In_2302,In_4422);
nor U3272 (N_3272,In_1059,In_4040);
or U3273 (N_3273,In_3972,In_2272);
nand U3274 (N_3274,In_4376,In_1571);
nand U3275 (N_3275,In_2027,In_1978);
nor U3276 (N_3276,In_3951,In_2097);
or U3277 (N_3277,In_920,In_4476);
nand U3278 (N_3278,In_290,In_3608);
nor U3279 (N_3279,In_2739,In_982);
nor U3280 (N_3280,In_4553,In_2918);
nand U3281 (N_3281,In_3788,In_2658);
xnor U3282 (N_3282,In_4468,In_443);
and U3283 (N_3283,In_2750,In_2664);
nand U3284 (N_3284,In_4802,In_3623);
and U3285 (N_3285,In_4273,In_4637);
nor U3286 (N_3286,In_2049,In_27);
and U3287 (N_3287,In_1455,In_4249);
and U3288 (N_3288,In_3289,In_478);
and U3289 (N_3289,In_227,In_4221);
nor U3290 (N_3290,In_2319,In_385);
nand U3291 (N_3291,In_4997,In_3197);
nand U3292 (N_3292,In_601,In_3030);
nor U3293 (N_3293,In_3018,In_2320);
xor U3294 (N_3294,In_472,In_4444);
and U3295 (N_3295,In_636,In_1607);
nor U3296 (N_3296,In_1813,In_976);
or U3297 (N_3297,In_3766,In_4276);
or U3298 (N_3298,In_1494,In_297);
and U3299 (N_3299,In_2578,In_377);
nand U3300 (N_3300,In_3402,In_1836);
and U3301 (N_3301,In_3281,In_717);
nor U3302 (N_3302,In_169,In_4798);
nand U3303 (N_3303,In_4490,In_3875);
nor U3304 (N_3304,In_3287,In_3800);
or U3305 (N_3305,In_34,In_1719);
nor U3306 (N_3306,In_1514,In_4864);
or U3307 (N_3307,In_3960,In_658);
or U3308 (N_3308,In_4226,In_1649);
xor U3309 (N_3309,In_3738,In_1194);
nand U3310 (N_3310,In_3317,In_4517);
or U3311 (N_3311,In_255,In_4452);
and U3312 (N_3312,In_1337,In_3208);
nand U3313 (N_3313,In_1109,In_4030);
nand U3314 (N_3314,In_3465,In_2996);
nor U3315 (N_3315,In_186,In_33);
nand U3316 (N_3316,In_3969,In_570);
nand U3317 (N_3317,In_1875,In_3158);
and U3318 (N_3318,In_235,In_2000);
and U3319 (N_3319,In_2227,In_4536);
or U3320 (N_3320,In_2660,In_2280);
nor U3321 (N_3321,In_3340,In_208);
or U3322 (N_3322,In_2825,In_2637);
or U3323 (N_3323,In_4172,In_1976);
and U3324 (N_3324,In_988,In_4890);
and U3325 (N_3325,In_3920,In_4451);
nand U3326 (N_3326,In_1136,In_1298);
or U3327 (N_3327,In_4424,In_1232);
nor U3328 (N_3328,In_1591,In_1584);
xnor U3329 (N_3329,In_3668,In_4085);
and U3330 (N_3330,In_2311,In_601);
nor U3331 (N_3331,In_968,In_3020);
xor U3332 (N_3332,In_797,In_4609);
and U3333 (N_3333,In_2253,In_2895);
or U3334 (N_3334,In_1981,In_2342);
xor U3335 (N_3335,In_2700,In_1452);
xor U3336 (N_3336,In_1314,In_4813);
or U3337 (N_3337,In_4031,In_1758);
xor U3338 (N_3338,In_4250,In_1232);
or U3339 (N_3339,In_4709,In_2388);
nand U3340 (N_3340,In_4021,In_4013);
or U3341 (N_3341,In_2862,In_3729);
nand U3342 (N_3342,In_1984,In_4807);
nand U3343 (N_3343,In_3841,In_1661);
nand U3344 (N_3344,In_2561,In_801);
nand U3345 (N_3345,In_2699,In_1036);
xor U3346 (N_3346,In_3386,In_3484);
nor U3347 (N_3347,In_1609,In_230);
or U3348 (N_3348,In_485,In_3453);
xnor U3349 (N_3349,In_3108,In_4604);
nand U3350 (N_3350,In_3649,In_4158);
nor U3351 (N_3351,In_975,In_203);
and U3352 (N_3352,In_1472,In_363);
or U3353 (N_3353,In_766,In_909);
or U3354 (N_3354,In_1578,In_3928);
nor U3355 (N_3355,In_984,In_380);
xor U3356 (N_3356,In_3595,In_3629);
nor U3357 (N_3357,In_1625,In_3581);
or U3358 (N_3358,In_4262,In_4899);
and U3359 (N_3359,In_3832,In_699);
nand U3360 (N_3360,In_3292,In_4651);
nor U3361 (N_3361,In_4443,In_2591);
and U3362 (N_3362,In_3788,In_1327);
nor U3363 (N_3363,In_706,In_3398);
xor U3364 (N_3364,In_1352,In_4406);
xor U3365 (N_3365,In_4602,In_151);
or U3366 (N_3366,In_4765,In_3752);
or U3367 (N_3367,In_2780,In_1395);
or U3368 (N_3368,In_3028,In_1397);
nor U3369 (N_3369,In_3761,In_2512);
or U3370 (N_3370,In_2243,In_1434);
nand U3371 (N_3371,In_3236,In_3504);
nand U3372 (N_3372,In_3003,In_679);
nand U3373 (N_3373,In_350,In_2244);
and U3374 (N_3374,In_3860,In_3601);
nand U3375 (N_3375,In_1061,In_1350);
xnor U3376 (N_3376,In_3417,In_894);
and U3377 (N_3377,In_1275,In_362);
xor U3378 (N_3378,In_1254,In_472);
or U3379 (N_3379,In_96,In_4034);
or U3380 (N_3380,In_635,In_559);
nor U3381 (N_3381,In_784,In_2217);
nand U3382 (N_3382,In_4210,In_2315);
xor U3383 (N_3383,In_1527,In_2145);
nand U3384 (N_3384,In_1012,In_2105);
or U3385 (N_3385,In_2766,In_1706);
or U3386 (N_3386,In_3177,In_1083);
and U3387 (N_3387,In_2224,In_953);
and U3388 (N_3388,In_3377,In_371);
or U3389 (N_3389,In_1876,In_4833);
nand U3390 (N_3390,In_2919,In_2454);
nand U3391 (N_3391,In_507,In_1310);
or U3392 (N_3392,In_125,In_691);
or U3393 (N_3393,In_4917,In_4687);
and U3394 (N_3394,In_4060,In_857);
nand U3395 (N_3395,In_223,In_4381);
nand U3396 (N_3396,In_925,In_1749);
xor U3397 (N_3397,In_568,In_4490);
and U3398 (N_3398,In_1483,In_2157);
or U3399 (N_3399,In_4916,In_4486);
nand U3400 (N_3400,In_1065,In_1498);
nor U3401 (N_3401,In_1203,In_3650);
or U3402 (N_3402,In_4238,In_4484);
xnor U3403 (N_3403,In_4407,In_2727);
xor U3404 (N_3404,In_2945,In_3897);
or U3405 (N_3405,In_2519,In_257);
nand U3406 (N_3406,In_4101,In_1325);
and U3407 (N_3407,In_692,In_1451);
nand U3408 (N_3408,In_4663,In_4785);
xor U3409 (N_3409,In_3650,In_686);
nor U3410 (N_3410,In_776,In_3542);
or U3411 (N_3411,In_484,In_2589);
or U3412 (N_3412,In_3512,In_2809);
nor U3413 (N_3413,In_970,In_2266);
nor U3414 (N_3414,In_3129,In_3407);
nand U3415 (N_3415,In_4046,In_4977);
nor U3416 (N_3416,In_4067,In_4964);
and U3417 (N_3417,In_1753,In_1374);
xnor U3418 (N_3418,In_541,In_1834);
nor U3419 (N_3419,In_504,In_1619);
nor U3420 (N_3420,In_1760,In_4540);
nand U3421 (N_3421,In_1454,In_2515);
nand U3422 (N_3422,In_164,In_4206);
nor U3423 (N_3423,In_4825,In_2857);
xnor U3424 (N_3424,In_3207,In_2133);
nand U3425 (N_3425,In_4681,In_3883);
or U3426 (N_3426,In_987,In_2796);
or U3427 (N_3427,In_729,In_4898);
xor U3428 (N_3428,In_2321,In_3973);
and U3429 (N_3429,In_4525,In_221);
or U3430 (N_3430,In_4534,In_491);
or U3431 (N_3431,In_743,In_2709);
nand U3432 (N_3432,In_3394,In_2179);
or U3433 (N_3433,In_3416,In_4429);
and U3434 (N_3434,In_1852,In_4725);
and U3435 (N_3435,In_4266,In_1022);
nor U3436 (N_3436,In_3747,In_1261);
and U3437 (N_3437,In_2003,In_3148);
nand U3438 (N_3438,In_2671,In_4376);
and U3439 (N_3439,In_4606,In_1892);
xor U3440 (N_3440,In_2566,In_1927);
and U3441 (N_3441,In_3901,In_4831);
xnor U3442 (N_3442,In_2018,In_1858);
and U3443 (N_3443,In_2253,In_917);
or U3444 (N_3444,In_529,In_2846);
nor U3445 (N_3445,In_1384,In_4739);
or U3446 (N_3446,In_559,In_3112);
nor U3447 (N_3447,In_3498,In_1132);
or U3448 (N_3448,In_1482,In_2435);
xnor U3449 (N_3449,In_3179,In_251);
or U3450 (N_3450,In_4665,In_2089);
xnor U3451 (N_3451,In_4998,In_391);
xor U3452 (N_3452,In_609,In_4242);
nand U3453 (N_3453,In_2969,In_1538);
and U3454 (N_3454,In_1380,In_4710);
and U3455 (N_3455,In_3626,In_1302);
xnor U3456 (N_3456,In_3224,In_2021);
and U3457 (N_3457,In_2150,In_4669);
or U3458 (N_3458,In_3452,In_2361);
or U3459 (N_3459,In_3695,In_224);
and U3460 (N_3460,In_3023,In_4626);
nand U3461 (N_3461,In_232,In_2460);
nor U3462 (N_3462,In_4750,In_4342);
nand U3463 (N_3463,In_2240,In_711);
xnor U3464 (N_3464,In_2427,In_4825);
nor U3465 (N_3465,In_3969,In_4349);
nand U3466 (N_3466,In_2515,In_4006);
and U3467 (N_3467,In_3834,In_3234);
or U3468 (N_3468,In_757,In_4664);
xnor U3469 (N_3469,In_316,In_3207);
xnor U3470 (N_3470,In_2715,In_1169);
nand U3471 (N_3471,In_4704,In_4167);
and U3472 (N_3472,In_996,In_230);
and U3473 (N_3473,In_2280,In_1063);
nand U3474 (N_3474,In_2580,In_1797);
or U3475 (N_3475,In_2889,In_1813);
xnor U3476 (N_3476,In_932,In_1916);
nor U3477 (N_3477,In_4479,In_523);
nor U3478 (N_3478,In_4937,In_1845);
nand U3479 (N_3479,In_1177,In_1240);
nand U3480 (N_3480,In_1793,In_3099);
or U3481 (N_3481,In_2886,In_241);
and U3482 (N_3482,In_1080,In_62);
or U3483 (N_3483,In_2274,In_105);
nand U3484 (N_3484,In_90,In_4135);
xor U3485 (N_3485,In_2860,In_1694);
xnor U3486 (N_3486,In_1756,In_1895);
nor U3487 (N_3487,In_2295,In_3364);
nor U3488 (N_3488,In_1799,In_3804);
and U3489 (N_3489,In_636,In_4549);
nand U3490 (N_3490,In_218,In_996);
xnor U3491 (N_3491,In_491,In_1599);
and U3492 (N_3492,In_1485,In_120);
nand U3493 (N_3493,In_2862,In_1611);
and U3494 (N_3494,In_4075,In_2423);
xnor U3495 (N_3495,In_2096,In_2140);
nor U3496 (N_3496,In_4596,In_751);
or U3497 (N_3497,In_1340,In_875);
xnor U3498 (N_3498,In_3630,In_784);
or U3499 (N_3499,In_904,In_4941);
nand U3500 (N_3500,In_1969,In_1195);
and U3501 (N_3501,In_420,In_1295);
nor U3502 (N_3502,In_1744,In_1677);
and U3503 (N_3503,In_3478,In_3871);
or U3504 (N_3504,In_843,In_39);
nand U3505 (N_3505,In_3233,In_2266);
nand U3506 (N_3506,In_2779,In_3608);
nand U3507 (N_3507,In_3644,In_4994);
or U3508 (N_3508,In_2253,In_2278);
nor U3509 (N_3509,In_2673,In_4832);
nor U3510 (N_3510,In_442,In_3007);
or U3511 (N_3511,In_1742,In_2012);
nor U3512 (N_3512,In_962,In_2354);
nand U3513 (N_3513,In_2963,In_889);
nand U3514 (N_3514,In_108,In_1538);
and U3515 (N_3515,In_2840,In_4934);
nand U3516 (N_3516,In_2060,In_3652);
and U3517 (N_3517,In_2268,In_2136);
nor U3518 (N_3518,In_1604,In_2032);
xor U3519 (N_3519,In_1035,In_4333);
nor U3520 (N_3520,In_277,In_3863);
nand U3521 (N_3521,In_3821,In_2193);
and U3522 (N_3522,In_3653,In_3447);
nand U3523 (N_3523,In_2267,In_3686);
nand U3524 (N_3524,In_959,In_955);
or U3525 (N_3525,In_3443,In_2257);
nand U3526 (N_3526,In_3323,In_481);
nand U3527 (N_3527,In_2424,In_433);
nor U3528 (N_3528,In_2701,In_4645);
or U3529 (N_3529,In_4587,In_1303);
nand U3530 (N_3530,In_4244,In_4923);
or U3531 (N_3531,In_2139,In_2614);
xnor U3532 (N_3532,In_3800,In_958);
xnor U3533 (N_3533,In_4222,In_2519);
or U3534 (N_3534,In_2522,In_4719);
nor U3535 (N_3535,In_1451,In_4778);
or U3536 (N_3536,In_2929,In_3716);
nor U3537 (N_3537,In_4176,In_2529);
and U3538 (N_3538,In_3496,In_2239);
nor U3539 (N_3539,In_2726,In_3877);
and U3540 (N_3540,In_3520,In_2418);
and U3541 (N_3541,In_4388,In_3670);
nand U3542 (N_3542,In_1298,In_2737);
or U3543 (N_3543,In_638,In_2711);
or U3544 (N_3544,In_322,In_2810);
xnor U3545 (N_3545,In_4712,In_3976);
nor U3546 (N_3546,In_2369,In_2428);
xnor U3547 (N_3547,In_1348,In_4439);
nor U3548 (N_3548,In_1707,In_4310);
nand U3549 (N_3549,In_1529,In_1824);
or U3550 (N_3550,In_333,In_4107);
or U3551 (N_3551,In_4359,In_2361);
or U3552 (N_3552,In_1752,In_4413);
xnor U3553 (N_3553,In_1407,In_4123);
xnor U3554 (N_3554,In_3580,In_1983);
or U3555 (N_3555,In_4610,In_1324);
or U3556 (N_3556,In_3210,In_3586);
or U3557 (N_3557,In_4202,In_77);
and U3558 (N_3558,In_1015,In_142);
nor U3559 (N_3559,In_1986,In_3995);
or U3560 (N_3560,In_146,In_4469);
or U3561 (N_3561,In_4129,In_878);
or U3562 (N_3562,In_2540,In_3904);
and U3563 (N_3563,In_2959,In_823);
nand U3564 (N_3564,In_220,In_3448);
xnor U3565 (N_3565,In_2052,In_35);
nor U3566 (N_3566,In_2874,In_2525);
and U3567 (N_3567,In_4305,In_4238);
nor U3568 (N_3568,In_648,In_920);
nor U3569 (N_3569,In_65,In_4560);
and U3570 (N_3570,In_1300,In_806);
xor U3571 (N_3571,In_3289,In_4646);
nor U3572 (N_3572,In_4960,In_2408);
and U3573 (N_3573,In_1279,In_772);
nand U3574 (N_3574,In_2486,In_3851);
or U3575 (N_3575,In_1409,In_1518);
or U3576 (N_3576,In_3097,In_1331);
nor U3577 (N_3577,In_4926,In_1896);
nand U3578 (N_3578,In_1392,In_4587);
nand U3579 (N_3579,In_2111,In_3792);
and U3580 (N_3580,In_4547,In_4805);
nand U3581 (N_3581,In_103,In_897);
or U3582 (N_3582,In_338,In_522);
xnor U3583 (N_3583,In_1501,In_713);
or U3584 (N_3584,In_3628,In_3108);
or U3585 (N_3585,In_4732,In_1440);
and U3586 (N_3586,In_1221,In_4789);
and U3587 (N_3587,In_2603,In_4272);
nor U3588 (N_3588,In_3891,In_2003);
or U3589 (N_3589,In_1305,In_4779);
and U3590 (N_3590,In_1345,In_3594);
or U3591 (N_3591,In_2752,In_3786);
xnor U3592 (N_3592,In_2411,In_1376);
nand U3593 (N_3593,In_4820,In_4718);
nand U3594 (N_3594,In_1479,In_3356);
and U3595 (N_3595,In_4869,In_1239);
nand U3596 (N_3596,In_3378,In_1346);
nor U3597 (N_3597,In_4038,In_1584);
or U3598 (N_3598,In_1101,In_2877);
nor U3599 (N_3599,In_3213,In_3727);
or U3600 (N_3600,In_2898,In_34);
xnor U3601 (N_3601,In_1894,In_628);
xnor U3602 (N_3602,In_3440,In_2885);
xnor U3603 (N_3603,In_2447,In_4092);
nand U3604 (N_3604,In_3210,In_4454);
nor U3605 (N_3605,In_963,In_901);
and U3606 (N_3606,In_3793,In_2781);
nand U3607 (N_3607,In_1020,In_1190);
or U3608 (N_3608,In_380,In_4990);
xor U3609 (N_3609,In_3882,In_933);
nor U3610 (N_3610,In_41,In_3985);
or U3611 (N_3611,In_1990,In_3275);
and U3612 (N_3612,In_569,In_1194);
nor U3613 (N_3613,In_4699,In_3185);
nand U3614 (N_3614,In_138,In_2553);
or U3615 (N_3615,In_3049,In_4946);
or U3616 (N_3616,In_3880,In_1428);
nand U3617 (N_3617,In_2597,In_4750);
or U3618 (N_3618,In_4971,In_1081);
or U3619 (N_3619,In_2530,In_368);
nand U3620 (N_3620,In_2843,In_1462);
nand U3621 (N_3621,In_2188,In_629);
xnor U3622 (N_3622,In_4193,In_1290);
nand U3623 (N_3623,In_3063,In_127);
xor U3624 (N_3624,In_3102,In_4055);
or U3625 (N_3625,In_457,In_1221);
xnor U3626 (N_3626,In_4677,In_4379);
and U3627 (N_3627,In_493,In_4958);
or U3628 (N_3628,In_4292,In_2736);
nand U3629 (N_3629,In_3309,In_2876);
nand U3630 (N_3630,In_3757,In_3628);
nand U3631 (N_3631,In_1011,In_295);
nor U3632 (N_3632,In_2501,In_6);
and U3633 (N_3633,In_3669,In_577);
and U3634 (N_3634,In_1762,In_2510);
and U3635 (N_3635,In_156,In_3861);
xnor U3636 (N_3636,In_3983,In_2218);
xnor U3637 (N_3637,In_802,In_3882);
nor U3638 (N_3638,In_1066,In_1767);
and U3639 (N_3639,In_466,In_828);
nor U3640 (N_3640,In_2181,In_3858);
xor U3641 (N_3641,In_2587,In_3169);
nand U3642 (N_3642,In_3024,In_332);
nand U3643 (N_3643,In_419,In_3391);
xor U3644 (N_3644,In_408,In_2460);
nor U3645 (N_3645,In_4650,In_2634);
nor U3646 (N_3646,In_1844,In_4852);
xnor U3647 (N_3647,In_2274,In_4660);
xnor U3648 (N_3648,In_2392,In_95);
or U3649 (N_3649,In_2152,In_1805);
and U3650 (N_3650,In_4061,In_1390);
nor U3651 (N_3651,In_3081,In_4196);
nor U3652 (N_3652,In_764,In_1355);
or U3653 (N_3653,In_4649,In_274);
and U3654 (N_3654,In_2911,In_439);
xnor U3655 (N_3655,In_462,In_2223);
and U3656 (N_3656,In_1739,In_2417);
and U3657 (N_3657,In_787,In_1484);
and U3658 (N_3658,In_597,In_1424);
xnor U3659 (N_3659,In_4058,In_595);
xor U3660 (N_3660,In_1598,In_3004);
nor U3661 (N_3661,In_3580,In_4904);
and U3662 (N_3662,In_2571,In_1266);
nand U3663 (N_3663,In_4743,In_961);
nand U3664 (N_3664,In_937,In_1705);
nand U3665 (N_3665,In_3351,In_4931);
xor U3666 (N_3666,In_4913,In_3299);
and U3667 (N_3667,In_4431,In_4832);
and U3668 (N_3668,In_1388,In_3577);
xor U3669 (N_3669,In_3770,In_4012);
nand U3670 (N_3670,In_1543,In_4375);
and U3671 (N_3671,In_1119,In_3305);
or U3672 (N_3672,In_1797,In_4342);
xor U3673 (N_3673,In_8,In_4993);
and U3674 (N_3674,In_4856,In_755);
and U3675 (N_3675,In_700,In_4266);
nor U3676 (N_3676,In_2965,In_1743);
or U3677 (N_3677,In_985,In_4785);
or U3678 (N_3678,In_3106,In_1919);
nand U3679 (N_3679,In_3561,In_2822);
or U3680 (N_3680,In_2424,In_1823);
and U3681 (N_3681,In_2559,In_1397);
nor U3682 (N_3682,In_3077,In_3172);
nand U3683 (N_3683,In_4823,In_4578);
xor U3684 (N_3684,In_4411,In_1869);
or U3685 (N_3685,In_2782,In_1710);
xnor U3686 (N_3686,In_3153,In_3188);
and U3687 (N_3687,In_2060,In_11);
nor U3688 (N_3688,In_4989,In_3406);
and U3689 (N_3689,In_4937,In_2750);
xor U3690 (N_3690,In_3454,In_3680);
xnor U3691 (N_3691,In_419,In_429);
xnor U3692 (N_3692,In_1627,In_3377);
or U3693 (N_3693,In_701,In_4262);
nor U3694 (N_3694,In_1231,In_3497);
or U3695 (N_3695,In_1568,In_2520);
or U3696 (N_3696,In_2715,In_1956);
and U3697 (N_3697,In_0,In_2812);
xor U3698 (N_3698,In_2512,In_4361);
nand U3699 (N_3699,In_1014,In_2970);
nand U3700 (N_3700,In_306,In_4444);
nand U3701 (N_3701,In_4296,In_3774);
and U3702 (N_3702,In_1060,In_271);
xnor U3703 (N_3703,In_1046,In_2939);
and U3704 (N_3704,In_2052,In_3968);
nand U3705 (N_3705,In_1913,In_1764);
and U3706 (N_3706,In_1285,In_2991);
and U3707 (N_3707,In_2801,In_4033);
nor U3708 (N_3708,In_2830,In_2541);
nand U3709 (N_3709,In_1451,In_630);
xnor U3710 (N_3710,In_2186,In_2794);
nor U3711 (N_3711,In_3627,In_1026);
or U3712 (N_3712,In_360,In_1053);
and U3713 (N_3713,In_4816,In_757);
xor U3714 (N_3714,In_2313,In_3840);
or U3715 (N_3715,In_3644,In_1275);
xnor U3716 (N_3716,In_2091,In_4675);
and U3717 (N_3717,In_3887,In_1689);
or U3718 (N_3718,In_4520,In_3513);
xnor U3719 (N_3719,In_3122,In_4401);
nor U3720 (N_3720,In_1377,In_2883);
xnor U3721 (N_3721,In_2805,In_4867);
nor U3722 (N_3722,In_4583,In_4104);
nor U3723 (N_3723,In_799,In_4085);
nor U3724 (N_3724,In_855,In_2798);
or U3725 (N_3725,In_1013,In_1714);
nor U3726 (N_3726,In_910,In_2947);
xor U3727 (N_3727,In_2334,In_548);
and U3728 (N_3728,In_2663,In_1721);
nand U3729 (N_3729,In_4708,In_54);
xor U3730 (N_3730,In_518,In_3345);
nor U3731 (N_3731,In_2378,In_4553);
or U3732 (N_3732,In_83,In_601);
nand U3733 (N_3733,In_4481,In_3400);
or U3734 (N_3734,In_1853,In_4377);
or U3735 (N_3735,In_4582,In_2770);
nand U3736 (N_3736,In_1229,In_935);
nor U3737 (N_3737,In_381,In_4555);
nor U3738 (N_3738,In_421,In_4151);
and U3739 (N_3739,In_3659,In_1890);
or U3740 (N_3740,In_278,In_2499);
nor U3741 (N_3741,In_1107,In_969);
nor U3742 (N_3742,In_4407,In_3938);
and U3743 (N_3743,In_1646,In_888);
nand U3744 (N_3744,In_3918,In_1111);
nand U3745 (N_3745,In_4289,In_2298);
nand U3746 (N_3746,In_2304,In_2658);
nor U3747 (N_3747,In_2155,In_1104);
nor U3748 (N_3748,In_3060,In_361);
nor U3749 (N_3749,In_1687,In_4519);
nand U3750 (N_3750,In_3484,In_4990);
or U3751 (N_3751,In_4501,In_595);
and U3752 (N_3752,In_1837,In_4421);
and U3753 (N_3753,In_3004,In_849);
and U3754 (N_3754,In_3257,In_2790);
xor U3755 (N_3755,In_4617,In_3104);
or U3756 (N_3756,In_3956,In_3387);
nor U3757 (N_3757,In_677,In_3686);
nand U3758 (N_3758,In_936,In_2);
nor U3759 (N_3759,In_3413,In_2232);
nand U3760 (N_3760,In_4339,In_4018);
nand U3761 (N_3761,In_1997,In_253);
and U3762 (N_3762,In_435,In_3720);
and U3763 (N_3763,In_2501,In_4719);
and U3764 (N_3764,In_2489,In_4885);
and U3765 (N_3765,In_4144,In_4880);
and U3766 (N_3766,In_4731,In_1142);
nor U3767 (N_3767,In_218,In_1073);
nor U3768 (N_3768,In_2548,In_1302);
or U3769 (N_3769,In_2353,In_4069);
and U3770 (N_3770,In_3823,In_4256);
nand U3771 (N_3771,In_3473,In_1759);
or U3772 (N_3772,In_1652,In_2421);
xor U3773 (N_3773,In_4306,In_3959);
nor U3774 (N_3774,In_467,In_1740);
or U3775 (N_3775,In_3528,In_1462);
nor U3776 (N_3776,In_4364,In_2446);
nor U3777 (N_3777,In_850,In_647);
xnor U3778 (N_3778,In_3418,In_3403);
and U3779 (N_3779,In_213,In_3747);
xnor U3780 (N_3780,In_3562,In_3026);
nand U3781 (N_3781,In_1708,In_2153);
nand U3782 (N_3782,In_415,In_4178);
xor U3783 (N_3783,In_4126,In_1985);
or U3784 (N_3784,In_2955,In_3800);
or U3785 (N_3785,In_4002,In_1710);
or U3786 (N_3786,In_517,In_2940);
nand U3787 (N_3787,In_712,In_78);
xnor U3788 (N_3788,In_3081,In_4982);
nand U3789 (N_3789,In_4353,In_4950);
xnor U3790 (N_3790,In_2641,In_3461);
or U3791 (N_3791,In_2278,In_1826);
nand U3792 (N_3792,In_2804,In_1320);
and U3793 (N_3793,In_4677,In_370);
nand U3794 (N_3794,In_686,In_1788);
and U3795 (N_3795,In_679,In_2470);
xnor U3796 (N_3796,In_2701,In_230);
and U3797 (N_3797,In_2274,In_1104);
or U3798 (N_3798,In_2912,In_4786);
nor U3799 (N_3799,In_9,In_1661);
nand U3800 (N_3800,In_4532,In_1670);
nand U3801 (N_3801,In_4515,In_3685);
nand U3802 (N_3802,In_3474,In_2981);
or U3803 (N_3803,In_1752,In_2586);
nand U3804 (N_3804,In_930,In_1034);
xor U3805 (N_3805,In_1426,In_1467);
nand U3806 (N_3806,In_774,In_3178);
or U3807 (N_3807,In_4356,In_4567);
nand U3808 (N_3808,In_4747,In_841);
or U3809 (N_3809,In_2673,In_462);
nand U3810 (N_3810,In_3621,In_1789);
nand U3811 (N_3811,In_810,In_4121);
xor U3812 (N_3812,In_2807,In_4238);
nand U3813 (N_3813,In_2275,In_2053);
nor U3814 (N_3814,In_2756,In_1228);
xor U3815 (N_3815,In_122,In_4752);
nand U3816 (N_3816,In_3660,In_4001);
or U3817 (N_3817,In_14,In_2945);
nand U3818 (N_3818,In_4671,In_1653);
and U3819 (N_3819,In_429,In_2609);
and U3820 (N_3820,In_2673,In_2893);
and U3821 (N_3821,In_3399,In_389);
nor U3822 (N_3822,In_4621,In_234);
or U3823 (N_3823,In_1297,In_3762);
and U3824 (N_3824,In_453,In_3400);
nand U3825 (N_3825,In_4105,In_2723);
nand U3826 (N_3826,In_4297,In_308);
or U3827 (N_3827,In_4066,In_144);
nor U3828 (N_3828,In_3706,In_4040);
or U3829 (N_3829,In_4338,In_4640);
nor U3830 (N_3830,In_1535,In_3630);
nor U3831 (N_3831,In_1650,In_3827);
xnor U3832 (N_3832,In_4342,In_1308);
xor U3833 (N_3833,In_266,In_1261);
nor U3834 (N_3834,In_2768,In_1201);
nand U3835 (N_3835,In_814,In_4426);
and U3836 (N_3836,In_1237,In_2058);
and U3837 (N_3837,In_2282,In_108);
and U3838 (N_3838,In_153,In_336);
or U3839 (N_3839,In_2028,In_4471);
or U3840 (N_3840,In_1221,In_1512);
or U3841 (N_3841,In_35,In_3880);
nor U3842 (N_3842,In_2325,In_1258);
xnor U3843 (N_3843,In_3216,In_3829);
xor U3844 (N_3844,In_3312,In_176);
xor U3845 (N_3845,In_1667,In_1856);
nor U3846 (N_3846,In_2576,In_3609);
or U3847 (N_3847,In_4369,In_3625);
or U3848 (N_3848,In_4870,In_2454);
and U3849 (N_3849,In_1365,In_4357);
or U3850 (N_3850,In_4758,In_3609);
and U3851 (N_3851,In_1908,In_1237);
nor U3852 (N_3852,In_3625,In_4575);
nand U3853 (N_3853,In_399,In_853);
or U3854 (N_3854,In_585,In_2934);
and U3855 (N_3855,In_3597,In_3712);
or U3856 (N_3856,In_3399,In_3643);
or U3857 (N_3857,In_3814,In_1933);
xnor U3858 (N_3858,In_1721,In_1339);
nand U3859 (N_3859,In_347,In_4441);
or U3860 (N_3860,In_188,In_4772);
xor U3861 (N_3861,In_4497,In_2053);
nor U3862 (N_3862,In_3892,In_1757);
or U3863 (N_3863,In_830,In_4746);
xnor U3864 (N_3864,In_497,In_3163);
nand U3865 (N_3865,In_3736,In_1356);
and U3866 (N_3866,In_2243,In_1245);
and U3867 (N_3867,In_3285,In_3633);
and U3868 (N_3868,In_1563,In_1579);
or U3869 (N_3869,In_4459,In_463);
nand U3870 (N_3870,In_2431,In_527);
or U3871 (N_3871,In_1483,In_2448);
nor U3872 (N_3872,In_3436,In_1996);
nand U3873 (N_3873,In_1521,In_544);
xnor U3874 (N_3874,In_4635,In_866);
xnor U3875 (N_3875,In_2565,In_3575);
and U3876 (N_3876,In_3272,In_2350);
or U3877 (N_3877,In_4911,In_2315);
and U3878 (N_3878,In_3229,In_2476);
or U3879 (N_3879,In_1520,In_550);
nand U3880 (N_3880,In_3248,In_4458);
or U3881 (N_3881,In_797,In_3795);
nand U3882 (N_3882,In_1218,In_2321);
or U3883 (N_3883,In_22,In_2444);
xnor U3884 (N_3884,In_4318,In_4090);
nor U3885 (N_3885,In_373,In_2024);
or U3886 (N_3886,In_1928,In_1675);
nand U3887 (N_3887,In_3319,In_3758);
or U3888 (N_3888,In_4170,In_4503);
nor U3889 (N_3889,In_790,In_2908);
and U3890 (N_3890,In_1784,In_4884);
xor U3891 (N_3891,In_4608,In_482);
or U3892 (N_3892,In_4660,In_360);
nand U3893 (N_3893,In_2129,In_3342);
and U3894 (N_3894,In_1326,In_615);
and U3895 (N_3895,In_4369,In_666);
and U3896 (N_3896,In_1965,In_4014);
and U3897 (N_3897,In_46,In_4410);
and U3898 (N_3898,In_1930,In_1437);
nor U3899 (N_3899,In_1497,In_4004);
and U3900 (N_3900,In_1922,In_3034);
and U3901 (N_3901,In_2773,In_1721);
xnor U3902 (N_3902,In_628,In_669);
nand U3903 (N_3903,In_3528,In_219);
nor U3904 (N_3904,In_1508,In_4622);
and U3905 (N_3905,In_2448,In_862);
nor U3906 (N_3906,In_3848,In_3534);
nor U3907 (N_3907,In_1295,In_2988);
xnor U3908 (N_3908,In_3653,In_786);
xnor U3909 (N_3909,In_78,In_444);
or U3910 (N_3910,In_3651,In_3819);
nor U3911 (N_3911,In_3586,In_3218);
or U3912 (N_3912,In_4167,In_3385);
or U3913 (N_3913,In_831,In_4071);
nand U3914 (N_3914,In_4962,In_1209);
or U3915 (N_3915,In_4465,In_527);
nand U3916 (N_3916,In_3576,In_53);
and U3917 (N_3917,In_4311,In_1589);
nand U3918 (N_3918,In_1417,In_846);
nor U3919 (N_3919,In_4834,In_2894);
nand U3920 (N_3920,In_4159,In_3906);
nand U3921 (N_3921,In_3132,In_2406);
xnor U3922 (N_3922,In_1664,In_4622);
xor U3923 (N_3923,In_4239,In_2790);
or U3924 (N_3924,In_3786,In_1304);
nand U3925 (N_3925,In_3258,In_764);
nor U3926 (N_3926,In_4458,In_4130);
or U3927 (N_3927,In_3210,In_462);
or U3928 (N_3928,In_127,In_1280);
xnor U3929 (N_3929,In_1142,In_3051);
and U3930 (N_3930,In_2972,In_3838);
and U3931 (N_3931,In_987,In_2152);
nor U3932 (N_3932,In_1557,In_3417);
nor U3933 (N_3933,In_3503,In_1823);
nor U3934 (N_3934,In_4478,In_73);
or U3935 (N_3935,In_4627,In_780);
xnor U3936 (N_3936,In_916,In_2074);
nand U3937 (N_3937,In_2892,In_472);
or U3938 (N_3938,In_2518,In_733);
or U3939 (N_3939,In_2192,In_3092);
nand U3940 (N_3940,In_3515,In_174);
or U3941 (N_3941,In_4451,In_464);
xor U3942 (N_3942,In_1481,In_802);
nand U3943 (N_3943,In_2746,In_2712);
and U3944 (N_3944,In_2602,In_4013);
and U3945 (N_3945,In_4245,In_4656);
nor U3946 (N_3946,In_3033,In_2745);
and U3947 (N_3947,In_2054,In_3033);
xor U3948 (N_3948,In_4151,In_2460);
nand U3949 (N_3949,In_3818,In_2553);
nand U3950 (N_3950,In_3773,In_4271);
xnor U3951 (N_3951,In_3032,In_2871);
nor U3952 (N_3952,In_2371,In_600);
xnor U3953 (N_3953,In_4895,In_3536);
xor U3954 (N_3954,In_566,In_3178);
nor U3955 (N_3955,In_2650,In_503);
or U3956 (N_3956,In_2490,In_2982);
nor U3957 (N_3957,In_3661,In_1054);
or U3958 (N_3958,In_2128,In_3216);
xnor U3959 (N_3959,In_3120,In_2759);
nand U3960 (N_3960,In_1783,In_51);
and U3961 (N_3961,In_4900,In_1117);
or U3962 (N_3962,In_214,In_1658);
nor U3963 (N_3963,In_3093,In_2182);
nand U3964 (N_3964,In_3523,In_640);
nand U3965 (N_3965,In_1105,In_4292);
nor U3966 (N_3966,In_475,In_1090);
nand U3967 (N_3967,In_2273,In_3967);
or U3968 (N_3968,In_367,In_3054);
xnor U3969 (N_3969,In_4161,In_2843);
and U3970 (N_3970,In_3866,In_3760);
or U3971 (N_3971,In_915,In_4341);
nor U3972 (N_3972,In_675,In_2056);
and U3973 (N_3973,In_313,In_2635);
and U3974 (N_3974,In_116,In_4295);
xnor U3975 (N_3975,In_1277,In_2847);
xor U3976 (N_3976,In_766,In_4314);
xnor U3977 (N_3977,In_4369,In_792);
nor U3978 (N_3978,In_341,In_3093);
or U3979 (N_3979,In_1958,In_327);
or U3980 (N_3980,In_4961,In_1593);
nor U3981 (N_3981,In_3216,In_3028);
xnor U3982 (N_3982,In_538,In_2533);
or U3983 (N_3983,In_2909,In_3001);
nor U3984 (N_3984,In_3662,In_1366);
nor U3985 (N_3985,In_185,In_3936);
nor U3986 (N_3986,In_2547,In_1895);
nand U3987 (N_3987,In_4040,In_2957);
nand U3988 (N_3988,In_4371,In_3961);
or U3989 (N_3989,In_3509,In_3396);
nand U3990 (N_3990,In_3695,In_4070);
nor U3991 (N_3991,In_1750,In_4080);
nor U3992 (N_3992,In_2857,In_1113);
or U3993 (N_3993,In_3631,In_3723);
xor U3994 (N_3994,In_1439,In_176);
and U3995 (N_3995,In_2015,In_3950);
nor U3996 (N_3996,In_3745,In_4462);
xnor U3997 (N_3997,In_1587,In_4962);
nand U3998 (N_3998,In_3637,In_308);
or U3999 (N_3999,In_2737,In_4367);
nand U4000 (N_4000,In_3747,In_3466);
nand U4001 (N_4001,In_4249,In_334);
nor U4002 (N_4002,In_2646,In_785);
nor U4003 (N_4003,In_2821,In_168);
or U4004 (N_4004,In_2157,In_3715);
nand U4005 (N_4005,In_549,In_4657);
or U4006 (N_4006,In_1599,In_262);
xnor U4007 (N_4007,In_1971,In_3025);
nor U4008 (N_4008,In_797,In_859);
xor U4009 (N_4009,In_3919,In_3758);
or U4010 (N_4010,In_4160,In_595);
nor U4011 (N_4011,In_624,In_3);
xnor U4012 (N_4012,In_1529,In_654);
or U4013 (N_4013,In_4041,In_747);
xor U4014 (N_4014,In_4210,In_4317);
xor U4015 (N_4015,In_1307,In_3914);
xor U4016 (N_4016,In_2664,In_1057);
or U4017 (N_4017,In_2719,In_4084);
nand U4018 (N_4018,In_3409,In_4104);
and U4019 (N_4019,In_4822,In_4695);
nor U4020 (N_4020,In_1810,In_4356);
nand U4021 (N_4021,In_2546,In_971);
and U4022 (N_4022,In_2333,In_2235);
and U4023 (N_4023,In_4691,In_4426);
or U4024 (N_4024,In_174,In_1712);
and U4025 (N_4025,In_2179,In_4319);
or U4026 (N_4026,In_2339,In_4109);
nor U4027 (N_4027,In_4558,In_859);
nand U4028 (N_4028,In_2275,In_3941);
nand U4029 (N_4029,In_1334,In_3475);
or U4030 (N_4030,In_3014,In_332);
and U4031 (N_4031,In_2686,In_2056);
or U4032 (N_4032,In_4294,In_3324);
or U4033 (N_4033,In_705,In_690);
or U4034 (N_4034,In_3218,In_3612);
or U4035 (N_4035,In_1163,In_3682);
xor U4036 (N_4036,In_3867,In_2068);
nor U4037 (N_4037,In_1084,In_4612);
nor U4038 (N_4038,In_1570,In_4546);
and U4039 (N_4039,In_4917,In_3205);
or U4040 (N_4040,In_958,In_605);
xnor U4041 (N_4041,In_46,In_4426);
and U4042 (N_4042,In_4966,In_4718);
nand U4043 (N_4043,In_3536,In_4628);
nor U4044 (N_4044,In_3689,In_1044);
nand U4045 (N_4045,In_3147,In_4435);
xnor U4046 (N_4046,In_2469,In_3496);
xnor U4047 (N_4047,In_4304,In_3815);
xnor U4048 (N_4048,In_3099,In_4229);
and U4049 (N_4049,In_4309,In_4975);
nor U4050 (N_4050,In_2101,In_1748);
and U4051 (N_4051,In_886,In_4744);
nand U4052 (N_4052,In_778,In_1619);
and U4053 (N_4053,In_352,In_4763);
nor U4054 (N_4054,In_2985,In_772);
nand U4055 (N_4055,In_14,In_311);
xor U4056 (N_4056,In_2616,In_816);
and U4057 (N_4057,In_2838,In_1175);
xnor U4058 (N_4058,In_2887,In_2348);
and U4059 (N_4059,In_4660,In_4383);
and U4060 (N_4060,In_1851,In_2262);
and U4061 (N_4061,In_1362,In_3536);
xnor U4062 (N_4062,In_3467,In_414);
nand U4063 (N_4063,In_2284,In_2083);
nand U4064 (N_4064,In_4097,In_2667);
or U4065 (N_4065,In_1357,In_3306);
and U4066 (N_4066,In_2782,In_4045);
nand U4067 (N_4067,In_4558,In_56);
nor U4068 (N_4068,In_4309,In_1897);
nor U4069 (N_4069,In_2444,In_4717);
and U4070 (N_4070,In_1306,In_476);
or U4071 (N_4071,In_2027,In_2154);
nor U4072 (N_4072,In_1474,In_849);
nand U4073 (N_4073,In_4773,In_1805);
nor U4074 (N_4074,In_301,In_3075);
nand U4075 (N_4075,In_2556,In_631);
nand U4076 (N_4076,In_1445,In_1237);
nor U4077 (N_4077,In_2331,In_4808);
and U4078 (N_4078,In_3439,In_2717);
nand U4079 (N_4079,In_3334,In_2752);
nor U4080 (N_4080,In_1259,In_3891);
and U4081 (N_4081,In_4600,In_4689);
or U4082 (N_4082,In_4909,In_2761);
or U4083 (N_4083,In_1410,In_1918);
and U4084 (N_4084,In_1364,In_347);
nor U4085 (N_4085,In_4066,In_4289);
nor U4086 (N_4086,In_2280,In_3476);
xnor U4087 (N_4087,In_1011,In_3404);
nor U4088 (N_4088,In_2656,In_3504);
xnor U4089 (N_4089,In_728,In_944);
xnor U4090 (N_4090,In_4578,In_2486);
xor U4091 (N_4091,In_4264,In_3390);
nand U4092 (N_4092,In_2595,In_1679);
and U4093 (N_4093,In_2782,In_2980);
and U4094 (N_4094,In_1090,In_3572);
nor U4095 (N_4095,In_4353,In_3764);
or U4096 (N_4096,In_3904,In_2295);
nor U4097 (N_4097,In_1271,In_1510);
xor U4098 (N_4098,In_568,In_129);
nor U4099 (N_4099,In_1952,In_4647);
nor U4100 (N_4100,In_697,In_2335);
nand U4101 (N_4101,In_910,In_4398);
nand U4102 (N_4102,In_2899,In_4026);
or U4103 (N_4103,In_1939,In_1360);
or U4104 (N_4104,In_1060,In_2683);
nor U4105 (N_4105,In_2150,In_326);
nand U4106 (N_4106,In_2063,In_796);
nor U4107 (N_4107,In_1087,In_3441);
nand U4108 (N_4108,In_2756,In_2901);
nand U4109 (N_4109,In_1809,In_2725);
or U4110 (N_4110,In_1649,In_4902);
nand U4111 (N_4111,In_3240,In_233);
xnor U4112 (N_4112,In_319,In_2057);
xor U4113 (N_4113,In_4494,In_4164);
xnor U4114 (N_4114,In_632,In_454);
and U4115 (N_4115,In_2961,In_2637);
nand U4116 (N_4116,In_4899,In_2067);
xnor U4117 (N_4117,In_3497,In_4871);
nor U4118 (N_4118,In_3257,In_1328);
nor U4119 (N_4119,In_4402,In_2661);
or U4120 (N_4120,In_4848,In_1727);
xor U4121 (N_4121,In_2414,In_4767);
nor U4122 (N_4122,In_3989,In_90);
nand U4123 (N_4123,In_1962,In_2799);
xnor U4124 (N_4124,In_1653,In_2438);
xnor U4125 (N_4125,In_3234,In_3452);
and U4126 (N_4126,In_1774,In_389);
nor U4127 (N_4127,In_734,In_2164);
nand U4128 (N_4128,In_4840,In_4690);
or U4129 (N_4129,In_2780,In_1348);
xnor U4130 (N_4130,In_950,In_3210);
and U4131 (N_4131,In_4367,In_2490);
nor U4132 (N_4132,In_4596,In_1762);
and U4133 (N_4133,In_233,In_2631);
nand U4134 (N_4134,In_1618,In_1636);
or U4135 (N_4135,In_3798,In_3907);
nand U4136 (N_4136,In_2023,In_892);
nand U4137 (N_4137,In_4244,In_2695);
nand U4138 (N_4138,In_196,In_2239);
or U4139 (N_4139,In_2086,In_2795);
xnor U4140 (N_4140,In_4208,In_4341);
nand U4141 (N_4141,In_2537,In_3290);
xnor U4142 (N_4142,In_603,In_2764);
xor U4143 (N_4143,In_3820,In_737);
nand U4144 (N_4144,In_2124,In_88);
nand U4145 (N_4145,In_4576,In_2942);
nand U4146 (N_4146,In_4682,In_3087);
or U4147 (N_4147,In_3391,In_2377);
and U4148 (N_4148,In_1958,In_1402);
nand U4149 (N_4149,In_324,In_1269);
nor U4150 (N_4150,In_2591,In_3765);
xor U4151 (N_4151,In_4055,In_1597);
xnor U4152 (N_4152,In_481,In_4652);
nor U4153 (N_4153,In_263,In_1580);
or U4154 (N_4154,In_4723,In_2511);
xor U4155 (N_4155,In_1768,In_620);
or U4156 (N_4156,In_1075,In_3347);
xor U4157 (N_4157,In_2275,In_1135);
xnor U4158 (N_4158,In_3964,In_1178);
nor U4159 (N_4159,In_1376,In_3587);
nor U4160 (N_4160,In_1330,In_452);
xor U4161 (N_4161,In_4374,In_3041);
or U4162 (N_4162,In_1247,In_97);
or U4163 (N_4163,In_1294,In_1924);
nor U4164 (N_4164,In_1184,In_2211);
and U4165 (N_4165,In_2236,In_2943);
nor U4166 (N_4166,In_4388,In_1246);
nand U4167 (N_4167,In_4846,In_1748);
xor U4168 (N_4168,In_1262,In_164);
and U4169 (N_4169,In_4183,In_104);
xnor U4170 (N_4170,In_4723,In_4255);
and U4171 (N_4171,In_2479,In_2221);
nor U4172 (N_4172,In_1155,In_1275);
or U4173 (N_4173,In_36,In_4005);
and U4174 (N_4174,In_1762,In_4515);
nor U4175 (N_4175,In_3074,In_3163);
or U4176 (N_4176,In_1408,In_3409);
or U4177 (N_4177,In_104,In_3854);
nor U4178 (N_4178,In_752,In_2709);
nand U4179 (N_4179,In_1344,In_1426);
and U4180 (N_4180,In_2268,In_3156);
xor U4181 (N_4181,In_4556,In_444);
nand U4182 (N_4182,In_55,In_428);
nand U4183 (N_4183,In_1528,In_1374);
nor U4184 (N_4184,In_36,In_1633);
and U4185 (N_4185,In_580,In_2269);
nand U4186 (N_4186,In_51,In_1038);
xnor U4187 (N_4187,In_3086,In_1096);
nand U4188 (N_4188,In_4656,In_1987);
nand U4189 (N_4189,In_4863,In_2119);
xnor U4190 (N_4190,In_3263,In_896);
and U4191 (N_4191,In_2457,In_2591);
nor U4192 (N_4192,In_3457,In_1358);
or U4193 (N_4193,In_3018,In_4585);
nor U4194 (N_4194,In_1676,In_4224);
and U4195 (N_4195,In_3801,In_3122);
xnor U4196 (N_4196,In_1986,In_3171);
nand U4197 (N_4197,In_719,In_3699);
xor U4198 (N_4198,In_38,In_4296);
and U4199 (N_4199,In_2881,In_2987);
or U4200 (N_4200,In_1870,In_3139);
or U4201 (N_4201,In_4248,In_4170);
and U4202 (N_4202,In_2819,In_2732);
or U4203 (N_4203,In_1606,In_4945);
or U4204 (N_4204,In_4462,In_1479);
xnor U4205 (N_4205,In_2514,In_2554);
xor U4206 (N_4206,In_1603,In_4457);
and U4207 (N_4207,In_243,In_4998);
and U4208 (N_4208,In_2386,In_4586);
xor U4209 (N_4209,In_3146,In_1458);
xnor U4210 (N_4210,In_1364,In_3373);
nor U4211 (N_4211,In_1665,In_2946);
xnor U4212 (N_4212,In_4586,In_2852);
and U4213 (N_4213,In_2940,In_2392);
or U4214 (N_4214,In_3866,In_2415);
or U4215 (N_4215,In_1040,In_137);
nand U4216 (N_4216,In_4916,In_2185);
xnor U4217 (N_4217,In_3503,In_3637);
nor U4218 (N_4218,In_1088,In_1376);
xnor U4219 (N_4219,In_1980,In_1967);
or U4220 (N_4220,In_3030,In_1898);
xor U4221 (N_4221,In_2454,In_3014);
nand U4222 (N_4222,In_3784,In_424);
nand U4223 (N_4223,In_1568,In_491);
nor U4224 (N_4224,In_2277,In_2073);
nor U4225 (N_4225,In_4686,In_105);
nand U4226 (N_4226,In_2682,In_4596);
nor U4227 (N_4227,In_1082,In_702);
and U4228 (N_4228,In_1793,In_885);
xor U4229 (N_4229,In_2584,In_1450);
or U4230 (N_4230,In_3615,In_4987);
nand U4231 (N_4231,In_2142,In_370);
or U4232 (N_4232,In_2939,In_2015);
nand U4233 (N_4233,In_790,In_3951);
xor U4234 (N_4234,In_487,In_1048);
nor U4235 (N_4235,In_3900,In_3562);
nand U4236 (N_4236,In_1448,In_3326);
nand U4237 (N_4237,In_3257,In_3740);
and U4238 (N_4238,In_531,In_4110);
xnor U4239 (N_4239,In_2336,In_3756);
xnor U4240 (N_4240,In_361,In_2259);
nand U4241 (N_4241,In_1934,In_3470);
xnor U4242 (N_4242,In_2358,In_3708);
and U4243 (N_4243,In_1653,In_1888);
or U4244 (N_4244,In_1492,In_4304);
or U4245 (N_4245,In_2007,In_4039);
nor U4246 (N_4246,In_3689,In_1150);
nor U4247 (N_4247,In_1288,In_399);
and U4248 (N_4248,In_600,In_2751);
and U4249 (N_4249,In_2232,In_1755);
xnor U4250 (N_4250,In_2406,In_3510);
xnor U4251 (N_4251,In_2459,In_2908);
nand U4252 (N_4252,In_342,In_1589);
and U4253 (N_4253,In_649,In_1252);
xnor U4254 (N_4254,In_1987,In_1719);
nor U4255 (N_4255,In_1680,In_4373);
or U4256 (N_4256,In_1046,In_2053);
nand U4257 (N_4257,In_1806,In_1485);
or U4258 (N_4258,In_2583,In_3132);
nor U4259 (N_4259,In_2798,In_1969);
nor U4260 (N_4260,In_2394,In_414);
nand U4261 (N_4261,In_2940,In_1530);
nor U4262 (N_4262,In_1198,In_557);
nand U4263 (N_4263,In_704,In_1316);
nand U4264 (N_4264,In_1111,In_1398);
nand U4265 (N_4265,In_1702,In_1391);
and U4266 (N_4266,In_2200,In_1399);
and U4267 (N_4267,In_110,In_982);
nand U4268 (N_4268,In_1515,In_1534);
nor U4269 (N_4269,In_1170,In_3159);
nor U4270 (N_4270,In_2994,In_2690);
xor U4271 (N_4271,In_3836,In_2752);
xor U4272 (N_4272,In_2093,In_3413);
xnor U4273 (N_4273,In_644,In_333);
nand U4274 (N_4274,In_2850,In_3982);
nand U4275 (N_4275,In_688,In_27);
or U4276 (N_4276,In_3248,In_1087);
or U4277 (N_4277,In_3552,In_975);
and U4278 (N_4278,In_2585,In_586);
xnor U4279 (N_4279,In_2758,In_3060);
nand U4280 (N_4280,In_1175,In_3134);
nor U4281 (N_4281,In_4142,In_4066);
nor U4282 (N_4282,In_3812,In_1558);
nand U4283 (N_4283,In_4488,In_544);
and U4284 (N_4284,In_3744,In_850);
and U4285 (N_4285,In_3349,In_3123);
xnor U4286 (N_4286,In_2730,In_4620);
xor U4287 (N_4287,In_2693,In_2551);
nor U4288 (N_4288,In_4511,In_3258);
nand U4289 (N_4289,In_2900,In_2676);
xor U4290 (N_4290,In_1279,In_2559);
xor U4291 (N_4291,In_391,In_3190);
and U4292 (N_4292,In_3363,In_4031);
nand U4293 (N_4293,In_1385,In_616);
nand U4294 (N_4294,In_3045,In_1636);
or U4295 (N_4295,In_526,In_2824);
nor U4296 (N_4296,In_4917,In_2193);
xnor U4297 (N_4297,In_1535,In_4996);
nor U4298 (N_4298,In_1982,In_352);
nor U4299 (N_4299,In_985,In_1380);
nor U4300 (N_4300,In_4300,In_4845);
or U4301 (N_4301,In_63,In_4309);
nand U4302 (N_4302,In_4693,In_1180);
and U4303 (N_4303,In_503,In_4826);
xor U4304 (N_4304,In_4713,In_4103);
or U4305 (N_4305,In_4116,In_2020);
nand U4306 (N_4306,In_666,In_3363);
or U4307 (N_4307,In_4165,In_4706);
nand U4308 (N_4308,In_3243,In_1051);
and U4309 (N_4309,In_3527,In_190);
nand U4310 (N_4310,In_1247,In_747);
nand U4311 (N_4311,In_2987,In_2070);
and U4312 (N_4312,In_3644,In_148);
xnor U4313 (N_4313,In_2904,In_4593);
and U4314 (N_4314,In_4336,In_905);
nand U4315 (N_4315,In_2503,In_4526);
or U4316 (N_4316,In_1738,In_4300);
nand U4317 (N_4317,In_2771,In_1100);
nand U4318 (N_4318,In_2026,In_2308);
nor U4319 (N_4319,In_4301,In_2893);
xnor U4320 (N_4320,In_1399,In_1626);
or U4321 (N_4321,In_633,In_2287);
xor U4322 (N_4322,In_3595,In_2344);
and U4323 (N_4323,In_1725,In_3027);
and U4324 (N_4324,In_916,In_752);
nand U4325 (N_4325,In_4102,In_2282);
nor U4326 (N_4326,In_4709,In_695);
nor U4327 (N_4327,In_4387,In_941);
xor U4328 (N_4328,In_4798,In_590);
xor U4329 (N_4329,In_3075,In_1207);
or U4330 (N_4330,In_2583,In_4618);
nor U4331 (N_4331,In_1894,In_951);
xor U4332 (N_4332,In_4484,In_962);
or U4333 (N_4333,In_2188,In_4322);
nor U4334 (N_4334,In_3887,In_4992);
or U4335 (N_4335,In_60,In_2923);
nor U4336 (N_4336,In_3044,In_4090);
nor U4337 (N_4337,In_746,In_3625);
nand U4338 (N_4338,In_1172,In_2088);
nand U4339 (N_4339,In_4515,In_1560);
xor U4340 (N_4340,In_1582,In_3999);
or U4341 (N_4341,In_233,In_306);
nor U4342 (N_4342,In_4562,In_1213);
xnor U4343 (N_4343,In_4628,In_2181);
xnor U4344 (N_4344,In_4720,In_3915);
xor U4345 (N_4345,In_2269,In_4545);
nor U4346 (N_4346,In_4831,In_1384);
and U4347 (N_4347,In_1109,In_4227);
xor U4348 (N_4348,In_1927,In_4323);
nor U4349 (N_4349,In_4147,In_4492);
xor U4350 (N_4350,In_4445,In_964);
and U4351 (N_4351,In_1125,In_3400);
nand U4352 (N_4352,In_4668,In_1321);
xnor U4353 (N_4353,In_1359,In_2957);
nor U4354 (N_4354,In_4856,In_293);
nand U4355 (N_4355,In_2048,In_4926);
and U4356 (N_4356,In_3001,In_2469);
or U4357 (N_4357,In_2353,In_954);
nand U4358 (N_4358,In_1678,In_228);
nand U4359 (N_4359,In_859,In_2395);
xnor U4360 (N_4360,In_1719,In_4681);
or U4361 (N_4361,In_573,In_148);
nand U4362 (N_4362,In_2546,In_473);
or U4363 (N_4363,In_3128,In_1507);
or U4364 (N_4364,In_346,In_4381);
nand U4365 (N_4365,In_3699,In_2028);
and U4366 (N_4366,In_697,In_4299);
nor U4367 (N_4367,In_1659,In_11);
and U4368 (N_4368,In_3922,In_1451);
xnor U4369 (N_4369,In_587,In_61);
and U4370 (N_4370,In_999,In_1093);
nand U4371 (N_4371,In_518,In_452);
nor U4372 (N_4372,In_3895,In_3296);
xor U4373 (N_4373,In_384,In_3261);
nor U4374 (N_4374,In_3588,In_3108);
or U4375 (N_4375,In_321,In_1468);
and U4376 (N_4376,In_2100,In_3253);
xnor U4377 (N_4377,In_1339,In_4159);
nor U4378 (N_4378,In_3221,In_3630);
nor U4379 (N_4379,In_114,In_3130);
xnor U4380 (N_4380,In_4273,In_3129);
nor U4381 (N_4381,In_4105,In_4798);
nand U4382 (N_4382,In_1567,In_468);
and U4383 (N_4383,In_3854,In_3055);
and U4384 (N_4384,In_3826,In_3945);
nand U4385 (N_4385,In_2156,In_4100);
nor U4386 (N_4386,In_1128,In_4805);
and U4387 (N_4387,In_1230,In_159);
nand U4388 (N_4388,In_604,In_932);
nor U4389 (N_4389,In_4990,In_3353);
nor U4390 (N_4390,In_1407,In_1776);
and U4391 (N_4391,In_4564,In_3447);
or U4392 (N_4392,In_3509,In_2199);
or U4393 (N_4393,In_3976,In_446);
or U4394 (N_4394,In_1351,In_4996);
nand U4395 (N_4395,In_802,In_96);
nor U4396 (N_4396,In_2332,In_1762);
nand U4397 (N_4397,In_3933,In_134);
xnor U4398 (N_4398,In_811,In_694);
nor U4399 (N_4399,In_158,In_2771);
nor U4400 (N_4400,In_1371,In_59);
or U4401 (N_4401,In_4878,In_1083);
or U4402 (N_4402,In_4194,In_3852);
xnor U4403 (N_4403,In_347,In_4332);
nor U4404 (N_4404,In_4461,In_4444);
nor U4405 (N_4405,In_4234,In_2916);
and U4406 (N_4406,In_1473,In_4413);
or U4407 (N_4407,In_3951,In_1819);
xnor U4408 (N_4408,In_245,In_2246);
and U4409 (N_4409,In_43,In_782);
xnor U4410 (N_4410,In_2316,In_2314);
nand U4411 (N_4411,In_3261,In_4446);
nand U4412 (N_4412,In_4842,In_3951);
xnor U4413 (N_4413,In_3744,In_4857);
nand U4414 (N_4414,In_531,In_4590);
nor U4415 (N_4415,In_1969,In_3706);
nand U4416 (N_4416,In_778,In_3115);
nor U4417 (N_4417,In_851,In_4956);
and U4418 (N_4418,In_2535,In_1982);
nand U4419 (N_4419,In_1862,In_1631);
and U4420 (N_4420,In_922,In_1257);
xor U4421 (N_4421,In_3079,In_4138);
and U4422 (N_4422,In_2667,In_2995);
or U4423 (N_4423,In_4953,In_1635);
nor U4424 (N_4424,In_4244,In_2018);
xor U4425 (N_4425,In_1804,In_283);
and U4426 (N_4426,In_3715,In_3613);
nand U4427 (N_4427,In_3448,In_439);
and U4428 (N_4428,In_2306,In_828);
xor U4429 (N_4429,In_3204,In_1013);
or U4430 (N_4430,In_4013,In_3453);
xor U4431 (N_4431,In_4921,In_2267);
nand U4432 (N_4432,In_177,In_1836);
xnor U4433 (N_4433,In_229,In_3462);
or U4434 (N_4434,In_2622,In_1653);
xor U4435 (N_4435,In_3444,In_54);
or U4436 (N_4436,In_967,In_707);
nand U4437 (N_4437,In_213,In_3599);
nor U4438 (N_4438,In_4392,In_3146);
nand U4439 (N_4439,In_2121,In_685);
nor U4440 (N_4440,In_4269,In_4872);
xor U4441 (N_4441,In_1930,In_226);
or U4442 (N_4442,In_3747,In_740);
or U4443 (N_4443,In_829,In_2617);
or U4444 (N_4444,In_992,In_4951);
or U4445 (N_4445,In_3779,In_3800);
xor U4446 (N_4446,In_2274,In_924);
or U4447 (N_4447,In_461,In_4106);
xnor U4448 (N_4448,In_3153,In_220);
nor U4449 (N_4449,In_1225,In_4343);
xnor U4450 (N_4450,In_1070,In_3463);
or U4451 (N_4451,In_3102,In_290);
or U4452 (N_4452,In_907,In_4135);
nand U4453 (N_4453,In_4921,In_883);
or U4454 (N_4454,In_393,In_1897);
or U4455 (N_4455,In_1393,In_392);
nor U4456 (N_4456,In_4816,In_3873);
or U4457 (N_4457,In_435,In_4071);
and U4458 (N_4458,In_243,In_2973);
or U4459 (N_4459,In_3376,In_1134);
or U4460 (N_4460,In_3763,In_1797);
and U4461 (N_4461,In_4997,In_1823);
nor U4462 (N_4462,In_1420,In_126);
nor U4463 (N_4463,In_399,In_4553);
nand U4464 (N_4464,In_1304,In_3135);
nand U4465 (N_4465,In_1334,In_4945);
and U4466 (N_4466,In_327,In_1589);
and U4467 (N_4467,In_4483,In_4652);
or U4468 (N_4468,In_4711,In_4398);
and U4469 (N_4469,In_262,In_1218);
and U4470 (N_4470,In_4470,In_14);
xor U4471 (N_4471,In_305,In_3111);
and U4472 (N_4472,In_3730,In_4178);
xnor U4473 (N_4473,In_2080,In_4065);
nand U4474 (N_4474,In_3234,In_678);
or U4475 (N_4475,In_4829,In_1670);
and U4476 (N_4476,In_3344,In_1476);
nor U4477 (N_4477,In_4277,In_3925);
xnor U4478 (N_4478,In_2202,In_4492);
xor U4479 (N_4479,In_4375,In_746);
xnor U4480 (N_4480,In_2540,In_613);
xor U4481 (N_4481,In_104,In_2656);
nand U4482 (N_4482,In_112,In_3720);
or U4483 (N_4483,In_1426,In_1954);
nand U4484 (N_4484,In_2958,In_2641);
and U4485 (N_4485,In_4810,In_1396);
and U4486 (N_4486,In_2217,In_4361);
xor U4487 (N_4487,In_4909,In_3435);
nand U4488 (N_4488,In_4294,In_1160);
xnor U4489 (N_4489,In_1498,In_742);
nor U4490 (N_4490,In_4808,In_1901);
and U4491 (N_4491,In_2340,In_1437);
or U4492 (N_4492,In_354,In_149);
nand U4493 (N_4493,In_2595,In_4004);
and U4494 (N_4494,In_847,In_3805);
nor U4495 (N_4495,In_2396,In_1324);
and U4496 (N_4496,In_3955,In_4302);
nand U4497 (N_4497,In_2738,In_3729);
nor U4498 (N_4498,In_2510,In_486);
or U4499 (N_4499,In_2544,In_2179);
nor U4500 (N_4500,In_463,In_1164);
nor U4501 (N_4501,In_2961,In_2994);
or U4502 (N_4502,In_2473,In_3043);
and U4503 (N_4503,In_364,In_4071);
and U4504 (N_4504,In_4507,In_3449);
nand U4505 (N_4505,In_1861,In_3180);
nand U4506 (N_4506,In_1043,In_3693);
nand U4507 (N_4507,In_392,In_2745);
nor U4508 (N_4508,In_730,In_4582);
nor U4509 (N_4509,In_4842,In_1008);
nand U4510 (N_4510,In_2726,In_3756);
and U4511 (N_4511,In_2203,In_1986);
or U4512 (N_4512,In_4622,In_3166);
nand U4513 (N_4513,In_608,In_3686);
and U4514 (N_4514,In_403,In_2136);
or U4515 (N_4515,In_3112,In_1630);
and U4516 (N_4516,In_2318,In_925);
or U4517 (N_4517,In_217,In_3023);
nand U4518 (N_4518,In_801,In_4029);
and U4519 (N_4519,In_3351,In_1684);
or U4520 (N_4520,In_4803,In_3113);
or U4521 (N_4521,In_4892,In_1920);
and U4522 (N_4522,In_1315,In_2063);
or U4523 (N_4523,In_36,In_3271);
nand U4524 (N_4524,In_1940,In_889);
nand U4525 (N_4525,In_2419,In_4487);
and U4526 (N_4526,In_1027,In_2080);
or U4527 (N_4527,In_3004,In_1501);
xnor U4528 (N_4528,In_1280,In_1899);
or U4529 (N_4529,In_2254,In_2606);
xor U4530 (N_4530,In_3285,In_4071);
nand U4531 (N_4531,In_1922,In_1772);
xnor U4532 (N_4532,In_2871,In_2511);
and U4533 (N_4533,In_313,In_2369);
xor U4534 (N_4534,In_1982,In_3679);
xnor U4535 (N_4535,In_3102,In_559);
or U4536 (N_4536,In_1076,In_2884);
nand U4537 (N_4537,In_1736,In_3448);
and U4538 (N_4538,In_2905,In_2745);
or U4539 (N_4539,In_2900,In_3567);
or U4540 (N_4540,In_10,In_1901);
nand U4541 (N_4541,In_2326,In_3385);
and U4542 (N_4542,In_1980,In_1227);
nand U4543 (N_4543,In_3057,In_4763);
and U4544 (N_4544,In_2051,In_1411);
nand U4545 (N_4545,In_2958,In_2738);
xnor U4546 (N_4546,In_732,In_4341);
and U4547 (N_4547,In_3411,In_3394);
and U4548 (N_4548,In_1750,In_1092);
xor U4549 (N_4549,In_2459,In_2197);
xor U4550 (N_4550,In_3158,In_1340);
or U4551 (N_4551,In_297,In_3102);
nor U4552 (N_4552,In_2418,In_120);
and U4553 (N_4553,In_864,In_4993);
xnor U4554 (N_4554,In_1821,In_2521);
or U4555 (N_4555,In_1482,In_1);
and U4556 (N_4556,In_846,In_1662);
xnor U4557 (N_4557,In_4498,In_4998);
or U4558 (N_4558,In_4375,In_3299);
and U4559 (N_4559,In_443,In_185);
and U4560 (N_4560,In_1917,In_2008);
and U4561 (N_4561,In_1584,In_4468);
or U4562 (N_4562,In_2866,In_2085);
nor U4563 (N_4563,In_125,In_3107);
or U4564 (N_4564,In_1212,In_2545);
xor U4565 (N_4565,In_2870,In_3379);
nor U4566 (N_4566,In_3030,In_1636);
xnor U4567 (N_4567,In_3294,In_732);
nor U4568 (N_4568,In_4184,In_2863);
nor U4569 (N_4569,In_3360,In_2580);
nand U4570 (N_4570,In_654,In_14);
nand U4571 (N_4571,In_2678,In_751);
or U4572 (N_4572,In_3396,In_4708);
nand U4573 (N_4573,In_3600,In_2053);
xnor U4574 (N_4574,In_3784,In_2071);
xnor U4575 (N_4575,In_280,In_1414);
nor U4576 (N_4576,In_3502,In_1911);
and U4577 (N_4577,In_4018,In_1583);
nor U4578 (N_4578,In_3442,In_4656);
nand U4579 (N_4579,In_3408,In_3250);
xnor U4580 (N_4580,In_1369,In_1659);
or U4581 (N_4581,In_449,In_3984);
nand U4582 (N_4582,In_2033,In_72);
and U4583 (N_4583,In_1944,In_4551);
nand U4584 (N_4584,In_3559,In_1069);
nand U4585 (N_4585,In_654,In_4633);
nand U4586 (N_4586,In_3524,In_3680);
nor U4587 (N_4587,In_3429,In_2434);
nand U4588 (N_4588,In_4266,In_1369);
nand U4589 (N_4589,In_1790,In_2576);
or U4590 (N_4590,In_706,In_894);
and U4591 (N_4591,In_4111,In_778);
xor U4592 (N_4592,In_620,In_979);
xnor U4593 (N_4593,In_3350,In_3997);
or U4594 (N_4594,In_3515,In_2336);
xnor U4595 (N_4595,In_4452,In_1159);
xnor U4596 (N_4596,In_3388,In_4606);
and U4597 (N_4597,In_4680,In_3183);
nand U4598 (N_4598,In_2036,In_4901);
nor U4599 (N_4599,In_1796,In_3888);
nor U4600 (N_4600,In_3554,In_3889);
xor U4601 (N_4601,In_4410,In_206);
nor U4602 (N_4602,In_2392,In_4018);
nor U4603 (N_4603,In_3059,In_1278);
or U4604 (N_4604,In_2715,In_3931);
nor U4605 (N_4605,In_144,In_1264);
or U4606 (N_4606,In_2591,In_2350);
or U4607 (N_4607,In_2856,In_1707);
or U4608 (N_4608,In_502,In_1555);
nor U4609 (N_4609,In_299,In_4969);
and U4610 (N_4610,In_591,In_39);
and U4611 (N_4611,In_4892,In_696);
xor U4612 (N_4612,In_2246,In_612);
nand U4613 (N_4613,In_533,In_2828);
nor U4614 (N_4614,In_92,In_1680);
and U4615 (N_4615,In_3043,In_3794);
nand U4616 (N_4616,In_659,In_4984);
or U4617 (N_4617,In_2285,In_2666);
and U4618 (N_4618,In_870,In_3356);
xor U4619 (N_4619,In_3796,In_2595);
xnor U4620 (N_4620,In_1918,In_2494);
nand U4621 (N_4621,In_499,In_4990);
and U4622 (N_4622,In_1478,In_839);
or U4623 (N_4623,In_3246,In_2976);
and U4624 (N_4624,In_2769,In_2734);
nand U4625 (N_4625,In_4052,In_1401);
xor U4626 (N_4626,In_557,In_695);
or U4627 (N_4627,In_1060,In_2523);
nor U4628 (N_4628,In_2495,In_4290);
or U4629 (N_4629,In_2741,In_3983);
and U4630 (N_4630,In_1586,In_3093);
xor U4631 (N_4631,In_1702,In_1354);
or U4632 (N_4632,In_1945,In_4629);
nor U4633 (N_4633,In_1437,In_1145);
nand U4634 (N_4634,In_2137,In_218);
nand U4635 (N_4635,In_271,In_3801);
nor U4636 (N_4636,In_4152,In_1440);
xor U4637 (N_4637,In_226,In_3767);
and U4638 (N_4638,In_447,In_734);
and U4639 (N_4639,In_3491,In_4889);
nand U4640 (N_4640,In_1286,In_3351);
nand U4641 (N_4641,In_882,In_2841);
xnor U4642 (N_4642,In_2041,In_3367);
and U4643 (N_4643,In_3933,In_462);
and U4644 (N_4644,In_1931,In_4755);
nor U4645 (N_4645,In_4813,In_3204);
or U4646 (N_4646,In_447,In_1412);
and U4647 (N_4647,In_1872,In_3176);
and U4648 (N_4648,In_512,In_4693);
and U4649 (N_4649,In_779,In_3319);
xor U4650 (N_4650,In_1957,In_2330);
xnor U4651 (N_4651,In_4014,In_1641);
or U4652 (N_4652,In_4674,In_1335);
nand U4653 (N_4653,In_4502,In_281);
and U4654 (N_4654,In_2937,In_1970);
nand U4655 (N_4655,In_591,In_1536);
nor U4656 (N_4656,In_669,In_4921);
or U4657 (N_4657,In_2495,In_1129);
or U4658 (N_4658,In_2344,In_527);
nand U4659 (N_4659,In_3022,In_2958);
and U4660 (N_4660,In_2262,In_4074);
or U4661 (N_4661,In_2142,In_3383);
or U4662 (N_4662,In_418,In_2987);
nor U4663 (N_4663,In_1799,In_4371);
xor U4664 (N_4664,In_4853,In_1620);
nor U4665 (N_4665,In_304,In_2115);
and U4666 (N_4666,In_4907,In_3234);
xnor U4667 (N_4667,In_3289,In_3421);
nor U4668 (N_4668,In_423,In_1956);
xnor U4669 (N_4669,In_3107,In_1097);
nand U4670 (N_4670,In_2548,In_1843);
nor U4671 (N_4671,In_1454,In_565);
or U4672 (N_4672,In_386,In_4400);
nor U4673 (N_4673,In_3230,In_1291);
nor U4674 (N_4674,In_185,In_4357);
nand U4675 (N_4675,In_142,In_4862);
or U4676 (N_4676,In_4274,In_4569);
xnor U4677 (N_4677,In_2574,In_3956);
xnor U4678 (N_4678,In_232,In_2630);
nand U4679 (N_4679,In_4548,In_1678);
nor U4680 (N_4680,In_2386,In_610);
or U4681 (N_4681,In_2438,In_2532);
and U4682 (N_4682,In_2888,In_3428);
xnor U4683 (N_4683,In_3251,In_1995);
nand U4684 (N_4684,In_2208,In_4419);
or U4685 (N_4685,In_480,In_1407);
and U4686 (N_4686,In_244,In_4974);
and U4687 (N_4687,In_2673,In_1462);
xnor U4688 (N_4688,In_955,In_3102);
nor U4689 (N_4689,In_4893,In_4955);
nand U4690 (N_4690,In_2021,In_77);
nand U4691 (N_4691,In_2552,In_3320);
nand U4692 (N_4692,In_4318,In_2134);
or U4693 (N_4693,In_2316,In_4116);
nor U4694 (N_4694,In_4777,In_2137);
nor U4695 (N_4695,In_2745,In_4621);
xor U4696 (N_4696,In_565,In_3169);
or U4697 (N_4697,In_2734,In_1939);
nand U4698 (N_4698,In_522,In_2451);
xor U4699 (N_4699,In_1909,In_2199);
nor U4700 (N_4700,In_550,In_2427);
xnor U4701 (N_4701,In_3536,In_3684);
xor U4702 (N_4702,In_714,In_1159);
nand U4703 (N_4703,In_4372,In_1712);
and U4704 (N_4704,In_1382,In_588);
nand U4705 (N_4705,In_3268,In_4907);
xnor U4706 (N_4706,In_4777,In_3479);
xnor U4707 (N_4707,In_2540,In_2045);
or U4708 (N_4708,In_602,In_1596);
nor U4709 (N_4709,In_499,In_4888);
nor U4710 (N_4710,In_4978,In_4791);
nand U4711 (N_4711,In_4922,In_2339);
or U4712 (N_4712,In_983,In_4194);
nor U4713 (N_4713,In_1704,In_4474);
nand U4714 (N_4714,In_2016,In_493);
nand U4715 (N_4715,In_504,In_984);
xor U4716 (N_4716,In_3394,In_4737);
nor U4717 (N_4717,In_3564,In_3685);
nor U4718 (N_4718,In_1033,In_2470);
nor U4719 (N_4719,In_152,In_4720);
and U4720 (N_4720,In_4051,In_4770);
or U4721 (N_4721,In_4978,In_2225);
xor U4722 (N_4722,In_2976,In_593);
xnor U4723 (N_4723,In_547,In_3883);
nand U4724 (N_4724,In_4632,In_4045);
nor U4725 (N_4725,In_3633,In_2583);
and U4726 (N_4726,In_2720,In_4066);
nand U4727 (N_4727,In_1638,In_3394);
and U4728 (N_4728,In_3939,In_213);
and U4729 (N_4729,In_1915,In_163);
nor U4730 (N_4730,In_3883,In_4286);
nand U4731 (N_4731,In_3068,In_4074);
nor U4732 (N_4732,In_2022,In_4337);
or U4733 (N_4733,In_3886,In_134);
or U4734 (N_4734,In_4754,In_1564);
or U4735 (N_4735,In_2521,In_2152);
nor U4736 (N_4736,In_567,In_544);
xor U4737 (N_4737,In_658,In_684);
nand U4738 (N_4738,In_1695,In_1386);
nand U4739 (N_4739,In_4859,In_3156);
xnor U4740 (N_4740,In_882,In_4316);
xnor U4741 (N_4741,In_901,In_1991);
nand U4742 (N_4742,In_2935,In_753);
xnor U4743 (N_4743,In_1889,In_707);
xor U4744 (N_4744,In_4786,In_1082);
or U4745 (N_4745,In_4022,In_751);
xnor U4746 (N_4746,In_3382,In_3957);
and U4747 (N_4747,In_4448,In_3005);
xnor U4748 (N_4748,In_1282,In_244);
or U4749 (N_4749,In_3781,In_3897);
or U4750 (N_4750,In_3310,In_4835);
or U4751 (N_4751,In_4976,In_3818);
nor U4752 (N_4752,In_53,In_4828);
or U4753 (N_4753,In_1427,In_3285);
and U4754 (N_4754,In_1116,In_2459);
and U4755 (N_4755,In_1180,In_182);
and U4756 (N_4756,In_381,In_1715);
nor U4757 (N_4757,In_748,In_4841);
nor U4758 (N_4758,In_531,In_4681);
nand U4759 (N_4759,In_3452,In_4711);
or U4760 (N_4760,In_1198,In_4339);
xor U4761 (N_4761,In_802,In_2673);
nor U4762 (N_4762,In_3891,In_624);
and U4763 (N_4763,In_2428,In_3165);
nand U4764 (N_4764,In_4918,In_696);
nor U4765 (N_4765,In_4998,In_2647);
nor U4766 (N_4766,In_123,In_1042);
xnor U4767 (N_4767,In_677,In_3236);
nand U4768 (N_4768,In_1646,In_4764);
nand U4769 (N_4769,In_1103,In_873);
or U4770 (N_4770,In_2941,In_1744);
nor U4771 (N_4771,In_736,In_4241);
or U4772 (N_4772,In_1515,In_3214);
and U4773 (N_4773,In_4799,In_3398);
nand U4774 (N_4774,In_1002,In_2361);
or U4775 (N_4775,In_3321,In_3101);
nand U4776 (N_4776,In_1143,In_2156);
or U4777 (N_4777,In_1020,In_4669);
nand U4778 (N_4778,In_1159,In_2717);
or U4779 (N_4779,In_2081,In_485);
xor U4780 (N_4780,In_4325,In_2644);
and U4781 (N_4781,In_1473,In_2085);
nand U4782 (N_4782,In_1515,In_3127);
and U4783 (N_4783,In_544,In_3927);
nor U4784 (N_4784,In_4444,In_2230);
nand U4785 (N_4785,In_435,In_4101);
and U4786 (N_4786,In_1631,In_665);
xor U4787 (N_4787,In_4821,In_3057);
nor U4788 (N_4788,In_3421,In_2872);
nand U4789 (N_4789,In_1825,In_4689);
nand U4790 (N_4790,In_746,In_4802);
nor U4791 (N_4791,In_1014,In_2063);
or U4792 (N_4792,In_4368,In_4656);
or U4793 (N_4793,In_34,In_4793);
or U4794 (N_4794,In_969,In_3673);
or U4795 (N_4795,In_3328,In_199);
xnor U4796 (N_4796,In_213,In_2961);
nor U4797 (N_4797,In_2220,In_1231);
nand U4798 (N_4798,In_2940,In_4866);
nor U4799 (N_4799,In_532,In_4435);
xnor U4800 (N_4800,In_3888,In_4403);
or U4801 (N_4801,In_417,In_1308);
nand U4802 (N_4802,In_2577,In_1528);
and U4803 (N_4803,In_1850,In_4532);
nor U4804 (N_4804,In_515,In_1346);
and U4805 (N_4805,In_2795,In_953);
and U4806 (N_4806,In_481,In_3240);
and U4807 (N_4807,In_3109,In_2696);
xnor U4808 (N_4808,In_3909,In_585);
nor U4809 (N_4809,In_3757,In_2698);
and U4810 (N_4810,In_2312,In_4474);
and U4811 (N_4811,In_2783,In_1435);
or U4812 (N_4812,In_2118,In_1916);
or U4813 (N_4813,In_1903,In_2032);
xor U4814 (N_4814,In_1863,In_4740);
or U4815 (N_4815,In_1254,In_3710);
and U4816 (N_4816,In_2488,In_3808);
xnor U4817 (N_4817,In_4904,In_4802);
nor U4818 (N_4818,In_1489,In_156);
nand U4819 (N_4819,In_2013,In_1830);
or U4820 (N_4820,In_520,In_3912);
nand U4821 (N_4821,In_2359,In_279);
xor U4822 (N_4822,In_4396,In_2320);
nand U4823 (N_4823,In_1277,In_3589);
nand U4824 (N_4824,In_4375,In_4750);
nor U4825 (N_4825,In_3251,In_3930);
nor U4826 (N_4826,In_1731,In_967);
xnor U4827 (N_4827,In_4863,In_1915);
xnor U4828 (N_4828,In_1992,In_2571);
xor U4829 (N_4829,In_3334,In_2842);
nand U4830 (N_4830,In_109,In_3983);
and U4831 (N_4831,In_1293,In_1734);
and U4832 (N_4832,In_4230,In_4774);
and U4833 (N_4833,In_1007,In_2968);
nor U4834 (N_4834,In_3417,In_2518);
nand U4835 (N_4835,In_4320,In_4451);
xnor U4836 (N_4836,In_3670,In_4385);
nand U4837 (N_4837,In_3553,In_4938);
xnor U4838 (N_4838,In_4146,In_4910);
nor U4839 (N_4839,In_1774,In_2619);
nor U4840 (N_4840,In_1260,In_4832);
and U4841 (N_4841,In_1598,In_4437);
nand U4842 (N_4842,In_3696,In_639);
and U4843 (N_4843,In_515,In_99);
nor U4844 (N_4844,In_971,In_964);
nand U4845 (N_4845,In_2577,In_3715);
nor U4846 (N_4846,In_748,In_2051);
and U4847 (N_4847,In_4312,In_894);
or U4848 (N_4848,In_3578,In_3246);
and U4849 (N_4849,In_4376,In_3052);
nor U4850 (N_4850,In_1618,In_3546);
nand U4851 (N_4851,In_3556,In_2975);
or U4852 (N_4852,In_3214,In_3279);
or U4853 (N_4853,In_4108,In_2806);
or U4854 (N_4854,In_1747,In_480);
nand U4855 (N_4855,In_909,In_3098);
or U4856 (N_4856,In_4882,In_2030);
and U4857 (N_4857,In_2347,In_2371);
and U4858 (N_4858,In_802,In_4074);
nand U4859 (N_4859,In_507,In_155);
and U4860 (N_4860,In_3553,In_478);
nor U4861 (N_4861,In_3959,In_2059);
and U4862 (N_4862,In_4625,In_276);
or U4863 (N_4863,In_1409,In_1826);
nand U4864 (N_4864,In_780,In_4756);
and U4865 (N_4865,In_3689,In_3369);
nand U4866 (N_4866,In_1908,In_1798);
and U4867 (N_4867,In_1656,In_713);
nand U4868 (N_4868,In_2371,In_4080);
nor U4869 (N_4869,In_2988,In_4721);
or U4870 (N_4870,In_1074,In_121);
and U4871 (N_4871,In_1674,In_998);
nor U4872 (N_4872,In_3195,In_3932);
nand U4873 (N_4873,In_989,In_4962);
and U4874 (N_4874,In_3366,In_3853);
and U4875 (N_4875,In_2549,In_3553);
nor U4876 (N_4876,In_610,In_4383);
or U4877 (N_4877,In_225,In_4913);
nor U4878 (N_4878,In_2519,In_3959);
or U4879 (N_4879,In_211,In_2237);
or U4880 (N_4880,In_3366,In_3607);
nand U4881 (N_4881,In_2636,In_2334);
nor U4882 (N_4882,In_68,In_4166);
nor U4883 (N_4883,In_4893,In_4660);
or U4884 (N_4884,In_2110,In_3779);
and U4885 (N_4885,In_1457,In_101);
or U4886 (N_4886,In_4398,In_1308);
nand U4887 (N_4887,In_456,In_1682);
or U4888 (N_4888,In_1992,In_4459);
nor U4889 (N_4889,In_2468,In_1396);
nor U4890 (N_4890,In_4729,In_8);
nand U4891 (N_4891,In_329,In_4339);
nor U4892 (N_4892,In_1406,In_3480);
or U4893 (N_4893,In_650,In_1204);
nand U4894 (N_4894,In_2520,In_4875);
xor U4895 (N_4895,In_4827,In_1866);
nand U4896 (N_4896,In_1465,In_2729);
nand U4897 (N_4897,In_2528,In_4213);
and U4898 (N_4898,In_1401,In_3327);
xnor U4899 (N_4899,In_487,In_3767);
and U4900 (N_4900,In_2436,In_876);
xor U4901 (N_4901,In_1335,In_4122);
nor U4902 (N_4902,In_3310,In_204);
nor U4903 (N_4903,In_4054,In_603);
and U4904 (N_4904,In_1935,In_4326);
and U4905 (N_4905,In_1981,In_1311);
nand U4906 (N_4906,In_3009,In_1842);
or U4907 (N_4907,In_1336,In_1840);
nand U4908 (N_4908,In_3583,In_457);
xnor U4909 (N_4909,In_2330,In_1788);
or U4910 (N_4910,In_702,In_1965);
and U4911 (N_4911,In_2411,In_2577);
or U4912 (N_4912,In_608,In_4903);
and U4913 (N_4913,In_939,In_611);
nand U4914 (N_4914,In_893,In_3323);
and U4915 (N_4915,In_3331,In_2110);
nor U4916 (N_4916,In_4072,In_3457);
or U4917 (N_4917,In_152,In_3823);
or U4918 (N_4918,In_4019,In_4044);
xor U4919 (N_4919,In_2653,In_1143);
nor U4920 (N_4920,In_4155,In_3145);
or U4921 (N_4921,In_509,In_3699);
xnor U4922 (N_4922,In_3904,In_3373);
and U4923 (N_4923,In_3518,In_3043);
nand U4924 (N_4924,In_3313,In_4641);
or U4925 (N_4925,In_1829,In_4799);
nand U4926 (N_4926,In_4613,In_4430);
nand U4927 (N_4927,In_3552,In_3201);
nand U4928 (N_4928,In_837,In_260);
nor U4929 (N_4929,In_4829,In_64);
or U4930 (N_4930,In_2465,In_1813);
and U4931 (N_4931,In_3226,In_4633);
xnor U4932 (N_4932,In_3346,In_515);
or U4933 (N_4933,In_269,In_314);
or U4934 (N_4934,In_3769,In_3865);
nand U4935 (N_4935,In_189,In_1241);
nand U4936 (N_4936,In_3452,In_500);
or U4937 (N_4937,In_3045,In_2334);
nand U4938 (N_4938,In_2854,In_2268);
and U4939 (N_4939,In_2753,In_2979);
nor U4940 (N_4940,In_1008,In_2560);
xor U4941 (N_4941,In_1753,In_4272);
or U4942 (N_4942,In_1907,In_325);
and U4943 (N_4943,In_4337,In_3061);
or U4944 (N_4944,In_321,In_2255);
or U4945 (N_4945,In_1678,In_884);
xor U4946 (N_4946,In_2686,In_3684);
xnor U4947 (N_4947,In_1806,In_1117);
and U4948 (N_4948,In_4115,In_4279);
or U4949 (N_4949,In_3750,In_4052);
or U4950 (N_4950,In_1004,In_1508);
nand U4951 (N_4951,In_399,In_974);
or U4952 (N_4952,In_119,In_1678);
and U4953 (N_4953,In_3111,In_520);
nand U4954 (N_4954,In_1177,In_1309);
or U4955 (N_4955,In_2090,In_742);
and U4956 (N_4956,In_307,In_319);
or U4957 (N_4957,In_550,In_975);
and U4958 (N_4958,In_3754,In_4627);
or U4959 (N_4959,In_3642,In_1199);
xnor U4960 (N_4960,In_168,In_553);
nand U4961 (N_4961,In_3194,In_710);
nand U4962 (N_4962,In_4109,In_4349);
nand U4963 (N_4963,In_4944,In_1505);
or U4964 (N_4964,In_830,In_4395);
or U4965 (N_4965,In_1385,In_1087);
or U4966 (N_4966,In_3470,In_4365);
nand U4967 (N_4967,In_3590,In_2936);
nand U4968 (N_4968,In_3658,In_3139);
nand U4969 (N_4969,In_1736,In_1829);
or U4970 (N_4970,In_2572,In_1530);
nand U4971 (N_4971,In_272,In_3596);
and U4972 (N_4972,In_396,In_361);
or U4973 (N_4973,In_2703,In_4400);
and U4974 (N_4974,In_4385,In_1948);
xor U4975 (N_4975,In_1473,In_1774);
xor U4976 (N_4976,In_1418,In_2028);
xor U4977 (N_4977,In_1110,In_371);
nand U4978 (N_4978,In_2210,In_1534);
nand U4979 (N_4979,In_3840,In_26);
xor U4980 (N_4980,In_717,In_4109);
and U4981 (N_4981,In_2095,In_2676);
xor U4982 (N_4982,In_1485,In_4789);
or U4983 (N_4983,In_4578,In_1414);
nand U4984 (N_4984,In_1220,In_4056);
xnor U4985 (N_4985,In_2390,In_611);
nand U4986 (N_4986,In_1277,In_266);
or U4987 (N_4987,In_2485,In_1885);
nor U4988 (N_4988,In_3340,In_1067);
or U4989 (N_4989,In_2706,In_4485);
nand U4990 (N_4990,In_2067,In_1134);
nand U4991 (N_4991,In_2362,In_374);
and U4992 (N_4992,In_2869,In_2845);
nor U4993 (N_4993,In_3808,In_1095);
or U4994 (N_4994,In_4626,In_2009);
and U4995 (N_4995,In_2582,In_1726);
xor U4996 (N_4996,In_59,In_520);
nand U4997 (N_4997,In_3854,In_3350);
nor U4998 (N_4998,In_4366,In_572);
xor U4999 (N_4999,In_3331,In_143);
nand U5000 (N_5000,In_4759,In_1367);
or U5001 (N_5001,In_3790,In_3553);
nor U5002 (N_5002,In_2371,In_556);
xnor U5003 (N_5003,In_1683,In_3727);
nor U5004 (N_5004,In_436,In_4845);
xnor U5005 (N_5005,In_3919,In_3332);
and U5006 (N_5006,In_2584,In_1791);
xnor U5007 (N_5007,In_3393,In_4222);
and U5008 (N_5008,In_1663,In_4771);
or U5009 (N_5009,In_2738,In_1428);
or U5010 (N_5010,In_3481,In_3068);
xor U5011 (N_5011,In_3624,In_4872);
nor U5012 (N_5012,In_4320,In_2609);
xor U5013 (N_5013,In_4267,In_2162);
xnor U5014 (N_5014,In_2877,In_354);
nand U5015 (N_5015,In_567,In_3812);
nor U5016 (N_5016,In_2062,In_2907);
nand U5017 (N_5017,In_154,In_1471);
nor U5018 (N_5018,In_3533,In_450);
xnor U5019 (N_5019,In_3578,In_2954);
nand U5020 (N_5020,In_3574,In_2080);
xor U5021 (N_5021,In_1470,In_4262);
nand U5022 (N_5022,In_1642,In_2079);
and U5023 (N_5023,In_3005,In_2756);
and U5024 (N_5024,In_4965,In_774);
and U5025 (N_5025,In_3344,In_1486);
and U5026 (N_5026,In_2641,In_4241);
or U5027 (N_5027,In_2609,In_1546);
or U5028 (N_5028,In_2571,In_1246);
or U5029 (N_5029,In_543,In_1029);
nor U5030 (N_5030,In_998,In_4368);
nor U5031 (N_5031,In_3622,In_3413);
and U5032 (N_5032,In_840,In_119);
nor U5033 (N_5033,In_915,In_2874);
nand U5034 (N_5034,In_3257,In_3097);
xnor U5035 (N_5035,In_2872,In_4105);
or U5036 (N_5036,In_2347,In_3780);
nand U5037 (N_5037,In_1526,In_4826);
nand U5038 (N_5038,In_3254,In_3748);
or U5039 (N_5039,In_4413,In_4315);
and U5040 (N_5040,In_1964,In_2629);
and U5041 (N_5041,In_1995,In_2908);
or U5042 (N_5042,In_3021,In_2815);
xnor U5043 (N_5043,In_2900,In_3999);
and U5044 (N_5044,In_4349,In_2955);
and U5045 (N_5045,In_376,In_2572);
nor U5046 (N_5046,In_4224,In_4317);
and U5047 (N_5047,In_4117,In_3858);
nor U5048 (N_5048,In_814,In_2710);
xor U5049 (N_5049,In_4204,In_3536);
xnor U5050 (N_5050,In_713,In_3408);
or U5051 (N_5051,In_3578,In_4716);
and U5052 (N_5052,In_727,In_258);
nor U5053 (N_5053,In_1477,In_2055);
nand U5054 (N_5054,In_1373,In_3007);
nor U5055 (N_5055,In_1868,In_198);
nor U5056 (N_5056,In_1366,In_3929);
and U5057 (N_5057,In_3005,In_1922);
nand U5058 (N_5058,In_618,In_4639);
or U5059 (N_5059,In_3898,In_3037);
nand U5060 (N_5060,In_3081,In_3717);
nor U5061 (N_5061,In_2937,In_706);
and U5062 (N_5062,In_2314,In_1863);
nand U5063 (N_5063,In_2062,In_4632);
nor U5064 (N_5064,In_770,In_2698);
nand U5065 (N_5065,In_3113,In_2979);
nor U5066 (N_5066,In_3442,In_3329);
xnor U5067 (N_5067,In_4019,In_2880);
and U5068 (N_5068,In_3783,In_3956);
nor U5069 (N_5069,In_1923,In_4551);
or U5070 (N_5070,In_2494,In_4622);
nand U5071 (N_5071,In_3791,In_1953);
nor U5072 (N_5072,In_537,In_4733);
xnor U5073 (N_5073,In_2646,In_2149);
nand U5074 (N_5074,In_2869,In_1445);
or U5075 (N_5075,In_2103,In_1378);
xnor U5076 (N_5076,In_4969,In_890);
and U5077 (N_5077,In_4167,In_4193);
nor U5078 (N_5078,In_618,In_3250);
xor U5079 (N_5079,In_3628,In_2646);
xor U5080 (N_5080,In_865,In_4594);
and U5081 (N_5081,In_3956,In_4626);
nand U5082 (N_5082,In_1655,In_4276);
xor U5083 (N_5083,In_4207,In_2707);
and U5084 (N_5084,In_1562,In_93);
nor U5085 (N_5085,In_4357,In_367);
nand U5086 (N_5086,In_4308,In_3871);
and U5087 (N_5087,In_307,In_572);
nand U5088 (N_5088,In_3761,In_3424);
nor U5089 (N_5089,In_3952,In_4422);
or U5090 (N_5090,In_4837,In_1807);
and U5091 (N_5091,In_2960,In_1731);
xnor U5092 (N_5092,In_1778,In_32);
and U5093 (N_5093,In_1953,In_2260);
xor U5094 (N_5094,In_4951,In_4191);
nor U5095 (N_5095,In_4130,In_1244);
nor U5096 (N_5096,In_3750,In_3384);
xor U5097 (N_5097,In_4882,In_4904);
xnor U5098 (N_5098,In_4738,In_3804);
and U5099 (N_5099,In_440,In_215);
or U5100 (N_5100,In_4024,In_876);
nand U5101 (N_5101,In_901,In_3012);
xnor U5102 (N_5102,In_3728,In_2004);
xor U5103 (N_5103,In_886,In_2729);
or U5104 (N_5104,In_2965,In_1253);
nand U5105 (N_5105,In_1062,In_4666);
nor U5106 (N_5106,In_4314,In_2355);
and U5107 (N_5107,In_1353,In_380);
xor U5108 (N_5108,In_494,In_870);
nor U5109 (N_5109,In_3423,In_3477);
nor U5110 (N_5110,In_3952,In_2308);
xnor U5111 (N_5111,In_877,In_254);
or U5112 (N_5112,In_4452,In_333);
xnor U5113 (N_5113,In_3139,In_4549);
or U5114 (N_5114,In_502,In_1940);
xnor U5115 (N_5115,In_359,In_1027);
xnor U5116 (N_5116,In_4098,In_6);
nand U5117 (N_5117,In_4343,In_3830);
nor U5118 (N_5118,In_2488,In_971);
nor U5119 (N_5119,In_3661,In_4691);
xor U5120 (N_5120,In_563,In_2828);
and U5121 (N_5121,In_4316,In_2671);
nand U5122 (N_5122,In_1504,In_2692);
nand U5123 (N_5123,In_1182,In_1960);
nand U5124 (N_5124,In_3682,In_675);
xnor U5125 (N_5125,In_3857,In_4571);
nand U5126 (N_5126,In_914,In_4833);
nor U5127 (N_5127,In_1974,In_3702);
or U5128 (N_5128,In_1944,In_1709);
nand U5129 (N_5129,In_1021,In_4601);
and U5130 (N_5130,In_1226,In_2121);
nor U5131 (N_5131,In_497,In_2499);
nor U5132 (N_5132,In_1053,In_1359);
xor U5133 (N_5133,In_3322,In_3701);
or U5134 (N_5134,In_248,In_2088);
or U5135 (N_5135,In_2314,In_2932);
xnor U5136 (N_5136,In_4861,In_1425);
nor U5137 (N_5137,In_3437,In_27);
nand U5138 (N_5138,In_4941,In_2197);
or U5139 (N_5139,In_1465,In_983);
nand U5140 (N_5140,In_4520,In_4402);
nand U5141 (N_5141,In_4767,In_1906);
nand U5142 (N_5142,In_2810,In_248);
nor U5143 (N_5143,In_3635,In_3851);
nand U5144 (N_5144,In_274,In_2451);
nand U5145 (N_5145,In_1443,In_3240);
nand U5146 (N_5146,In_2350,In_2945);
nand U5147 (N_5147,In_1947,In_3638);
or U5148 (N_5148,In_2805,In_3123);
or U5149 (N_5149,In_4582,In_4916);
xnor U5150 (N_5150,In_4414,In_2424);
nor U5151 (N_5151,In_4990,In_1266);
nand U5152 (N_5152,In_2775,In_1231);
and U5153 (N_5153,In_920,In_733);
nor U5154 (N_5154,In_3450,In_1892);
or U5155 (N_5155,In_4030,In_963);
xnor U5156 (N_5156,In_1957,In_2354);
xor U5157 (N_5157,In_280,In_380);
or U5158 (N_5158,In_1657,In_3678);
xor U5159 (N_5159,In_162,In_1902);
nor U5160 (N_5160,In_3060,In_1409);
or U5161 (N_5161,In_2803,In_2489);
or U5162 (N_5162,In_3058,In_4983);
nor U5163 (N_5163,In_2734,In_1032);
nor U5164 (N_5164,In_4220,In_2525);
or U5165 (N_5165,In_4888,In_3142);
xor U5166 (N_5166,In_2968,In_3053);
and U5167 (N_5167,In_216,In_479);
or U5168 (N_5168,In_1052,In_4550);
nand U5169 (N_5169,In_1946,In_895);
xor U5170 (N_5170,In_4397,In_281);
and U5171 (N_5171,In_1131,In_2654);
nand U5172 (N_5172,In_3969,In_3179);
and U5173 (N_5173,In_4826,In_4574);
and U5174 (N_5174,In_1305,In_2620);
or U5175 (N_5175,In_4020,In_4472);
or U5176 (N_5176,In_3797,In_1917);
and U5177 (N_5177,In_228,In_361);
or U5178 (N_5178,In_634,In_1290);
nand U5179 (N_5179,In_3436,In_576);
nand U5180 (N_5180,In_4780,In_4491);
or U5181 (N_5181,In_3545,In_1749);
nand U5182 (N_5182,In_2709,In_1047);
and U5183 (N_5183,In_1007,In_2156);
nand U5184 (N_5184,In_1465,In_3736);
nand U5185 (N_5185,In_3928,In_3872);
and U5186 (N_5186,In_1691,In_2558);
and U5187 (N_5187,In_2575,In_2009);
or U5188 (N_5188,In_1429,In_2403);
nand U5189 (N_5189,In_2304,In_4318);
nor U5190 (N_5190,In_4640,In_1447);
xnor U5191 (N_5191,In_304,In_3644);
or U5192 (N_5192,In_2044,In_2795);
or U5193 (N_5193,In_3826,In_2755);
nand U5194 (N_5194,In_2222,In_798);
or U5195 (N_5195,In_2958,In_4863);
xor U5196 (N_5196,In_167,In_3858);
or U5197 (N_5197,In_311,In_357);
and U5198 (N_5198,In_3114,In_915);
and U5199 (N_5199,In_312,In_3686);
nor U5200 (N_5200,In_4635,In_971);
nand U5201 (N_5201,In_510,In_4349);
or U5202 (N_5202,In_4291,In_360);
nor U5203 (N_5203,In_3912,In_3392);
nand U5204 (N_5204,In_582,In_2340);
and U5205 (N_5205,In_2047,In_3634);
and U5206 (N_5206,In_875,In_2712);
nor U5207 (N_5207,In_4803,In_866);
nand U5208 (N_5208,In_1202,In_3657);
nor U5209 (N_5209,In_2244,In_4539);
nor U5210 (N_5210,In_160,In_475);
nand U5211 (N_5211,In_4911,In_2763);
and U5212 (N_5212,In_4898,In_218);
nand U5213 (N_5213,In_152,In_1731);
nand U5214 (N_5214,In_1821,In_36);
or U5215 (N_5215,In_4810,In_1927);
xnor U5216 (N_5216,In_2556,In_2435);
nor U5217 (N_5217,In_3237,In_1115);
nand U5218 (N_5218,In_3068,In_3152);
nand U5219 (N_5219,In_2385,In_1936);
or U5220 (N_5220,In_3838,In_4287);
and U5221 (N_5221,In_1450,In_2028);
nor U5222 (N_5222,In_4246,In_3403);
nand U5223 (N_5223,In_3739,In_1554);
nor U5224 (N_5224,In_3932,In_4864);
xor U5225 (N_5225,In_4719,In_4400);
nor U5226 (N_5226,In_3665,In_1397);
nand U5227 (N_5227,In_846,In_683);
xnor U5228 (N_5228,In_4466,In_100);
nand U5229 (N_5229,In_3071,In_2218);
nor U5230 (N_5230,In_3619,In_45);
nand U5231 (N_5231,In_902,In_3200);
xnor U5232 (N_5232,In_1399,In_1572);
or U5233 (N_5233,In_307,In_2588);
and U5234 (N_5234,In_4849,In_4437);
nor U5235 (N_5235,In_70,In_2637);
xor U5236 (N_5236,In_978,In_4355);
nor U5237 (N_5237,In_4025,In_3597);
nor U5238 (N_5238,In_3753,In_4654);
or U5239 (N_5239,In_4111,In_2614);
or U5240 (N_5240,In_2568,In_1631);
and U5241 (N_5241,In_3182,In_4383);
nor U5242 (N_5242,In_1932,In_665);
nor U5243 (N_5243,In_2390,In_4850);
and U5244 (N_5244,In_1576,In_980);
xor U5245 (N_5245,In_752,In_3187);
and U5246 (N_5246,In_2812,In_4596);
xor U5247 (N_5247,In_2854,In_1674);
nand U5248 (N_5248,In_2330,In_1292);
and U5249 (N_5249,In_2675,In_339);
or U5250 (N_5250,In_3599,In_1365);
or U5251 (N_5251,In_2133,In_158);
nand U5252 (N_5252,In_1452,In_2364);
or U5253 (N_5253,In_4956,In_1956);
and U5254 (N_5254,In_2790,In_4344);
or U5255 (N_5255,In_3930,In_2622);
xor U5256 (N_5256,In_4506,In_2904);
or U5257 (N_5257,In_905,In_3916);
or U5258 (N_5258,In_1255,In_3812);
nor U5259 (N_5259,In_2888,In_1513);
nor U5260 (N_5260,In_531,In_889);
xnor U5261 (N_5261,In_191,In_3622);
xor U5262 (N_5262,In_1483,In_1871);
and U5263 (N_5263,In_4852,In_3429);
xor U5264 (N_5264,In_2325,In_4031);
and U5265 (N_5265,In_1901,In_4787);
xnor U5266 (N_5266,In_3517,In_3770);
nor U5267 (N_5267,In_1120,In_4087);
and U5268 (N_5268,In_3041,In_849);
or U5269 (N_5269,In_3838,In_2338);
xor U5270 (N_5270,In_3686,In_1600);
nor U5271 (N_5271,In_3417,In_2522);
xor U5272 (N_5272,In_4404,In_1298);
and U5273 (N_5273,In_4278,In_2086);
and U5274 (N_5274,In_2834,In_4989);
nor U5275 (N_5275,In_1422,In_138);
nand U5276 (N_5276,In_1704,In_3632);
or U5277 (N_5277,In_4648,In_1588);
and U5278 (N_5278,In_4047,In_3579);
nand U5279 (N_5279,In_3092,In_4296);
nand U5280 (N_5280,In_4256,In_868);
nor U5281 (N_5281,In_755,In_3215);
and U5282 (N_5282,In_2802,In_3298);
xnor U5283 (N_5283,In_549,In_3477);
nand U5284 (N_5284,In_4423,In_1698);
xor U5285 (N_5285,In_148,In_4371);
xnor U5286 (N_5286,In_1917,In_4200);
xor U5287 (N_5287,In_4290,In_1462);
or U5288 (N_5288,In_2044,In_1843);
xor U5289 (N_5289,In_3937,In_3258);
or U5290 (N_5290,In_2300,In_1250);
xnor U5291 (N_5291,In_4606,In_2972);
and U5292 (N_5292,In_1772,In_799);
xor U5293 (N_5293,In_1741,In_4560);
or U5294 (N_5294,In_612,In_4233);
nand U5295 (N_5295,In_1975,In_4828);
nor U5296 (N_5296,In_3430,In_1467);
xor U5297 (N_5297,In_4576,In_4173);
xor U5298 (N_5298,In_4463,In_3036);
nand U5299 (N_5299,In_143,In_1883);
nand U5300 (N_5300,In_3553,In_935);
xnor U5301 (N_5301,In_2855,In_3261);
nand U5302 (N_5302,In_1852,In_3568);
and U5303 (N_5303,In_4371,In_2830);
xnor U5304 (N_5304,In_3917,In_2136);
nand U5305 (N_5305,In_562,In_3849);
nand U5306 (N_5306,In_1289,In_595);
nor U5307 (N_5307,In_4483,In_3154);
nand U5308 (N_5308,In_3393,In_3170);
nor U5309 (N_5309,In_4167,In_4882);
nand U5310 (N_5310,In_4594,In_4304);
xnor U5311 (N_5311,In_4771,In_1014);
xnor U5312 (N_5312,In_2128,In_309);
nand U5313 (N_5313,In_4764,In_1395);
and U5314 (N_5314,In_1911,In_116);
nor U5315 (N_5315,In_1706,In_756);
or U5316 (N_5316,In_4903,In_4136);
nor U5317 (N_5317,In_2394,In_2286);
and U5318 (N_5318,In_968,In_3195);
nand U5319 (N_5319,In_2822,In_4418);
or U5320 (N_5320,In_3420,In_1982);
nor U5321 (N_5321,In_1741,In_853);
or U5322 (N_5322,In_4556,In_4435);
nand U5323 (N_5323,In_2633,In_3574);
xnor U5324 (N_5324,In_3725,In_4160);
xnor U5325 (N_5325,In_3824,In_148);
nand U5326 (N_5326,In_3509,In_63);
or U5327 (N_5327,In_3679,In_1757);
nor U5328 (N_5328,In_1071,In_1179);
or U5329 (N_5329,In_2874,In_3513);
nand U5330 (N_5330,In_4999,In_3800);
or U5331 (N_5331,In_1738,In_2963);
nand U5332 (N_5332,In_1954,In_2774);
xor U5333 (N_5333,In_1978,In_1277);
xnor U5334 (N_5334,In_4389,In_2506);
and U5335 (N_5335,In_891,In_2236);
or U5336 (N_5336,In_389,In_3411);
and U5337 (N_5337,In_534,In_590);
or U5338 (N_5338,In_4095,In_4757);
xnor U5339 (N_5339,In_2307,In_4479);
xnor U5340 (N_5340,In_758,In_3910);
or U5341 (N_5341,In_1058,In_353);
or U5342 (N_5342,In_4657,In_18);
and U5343 (N_5343,In_2811,In_4909);
nand U5344 (N_5344,In_4211,In_350);
nor U5345 (N_5345,In_993,In_166);
or U5346 (N_5346,In_1955,In_2244);
and U5347 (N_5347,In_1756,In_3789);
or U5348 (N_5348,In_1177,In_1221);
nor U5349 (N_5349,In_2173,In_3671);
nor U5350 (N_5350,In_3269,In_2449);
and U5351 (N_5351,In_1334,In_3648);
nor U5352 (N_5352,In_1854,In_4421);
nand U5353 (N_5353,In_4565,In_1086);
nor U5354 (N_5354,In_4184,In_3043);
nand U5355 (N_5355,In_4319,In_3884);
nand U5356 (N_5356,In_2356,In_1403);
nor U5357 (N_5357,In_1997,In_2700);
xor U5358 (N_5358,In_3934,In_1810);
and U5359 (N_5359,In_468,In_1595);
xor U5360 (N_5360,In_4569,In_3753);
and U5361 (N_5361,In_2303,In_1212);
and U5362 (N_5362,In_964,In_1387);
xnor U5363 (N_5363,In_2339,In_1609);
or U5364 (N_5364,In_1298,In_2995);
and U5365 (N_5365,In_2905,In_3275);
and U5366 (N_5366,In_4885,In_3536);
nand U5367 (N_5367,In_499,In_73);
and U5368 (N_5368,In_2476,In_2024);
xnor U5369 (N_5369,In_3266,In_1838);
or U5370 (N_5370,In_4025,In_443);
nand U5371 (N_5371,In_3611,In_3482);
nand U5372 (N_5372,In_1180,In_2301);
and U5373 (N_5373,In_3425,In_3096);
and U5374 (N_5374,In_4595,In_1800);
and U5375 (N_5375,In_830,In_3180);
and U5376 (N_5376,In_4158,In_4200);
xnor U5377 (N_5377,In_4037,In_912);
nand U5378 (N_5378,In_3542,In_513);
xor U5379 (N_5379,In_1172,In_1246);
and U5380 (N_5380,In_2772,In_2285);
nand U5381 (N_5381,In_1115,In_4321);
nand U5382 (N_5382,In_4258,In_4582);
xnor U5383 (N_5383,In_1200,In_833);
or U5384 (N_5384,In_3297,In_3865);
or U5385 (N_5385,In_2270,In_1255);
or U5386 (N_5386,In_3265,In_1510);
nor U5387 (N_5387,In_4772,In_2424);
nor U5388 (N_5388,In_4912,In_2114);
nor U5389 (N_5389,In_1865,In_2580);
xnor U5390 (N_5390,In_4770,In_2609);
nor U5391 (N_5391,In_1005,In_3303);
nand U5392 (N_5392,In_501,In_127);
nand U5393 (N_5393,In_244,In_2771);
nand U5394 (N_5394,In_4851,In_2594);
and U5395 (N_5395,In_4796,In_3625);
or U5396 (N_5396,In_3130,In_510);
nand U5397 (N_5397,In_4584,In_2808);
xor U5398 (N_5398,In_1591,In_1441);
xor U5399 (N_5399,In_3147,In_1532);
nor U5400 (N_5400,In_2934,In_3887);
or U5401 (N_5401,In_4552,In_3014);
and U5402 (N_5402,In_4925,In_762);
or U5403 (N_5403,In_738,In_4185);
nor U5404 (N_5404,In_3295,In_58);
nand U5405 (N_5405,In_3490,In_2357);
or U5406 (N_5406,In_3398,In_4322);
nor U5407 (N_5407,In_1269,In_3729);
nor U5408 (N_5408,In_1079,In_2090);
xor U5409 (N_5409,In_3432,In_1953);
nor U5410 (N_5410,In_3020,In_3738);
xnor U5411 (N_5411,In_4671,In_286);
or U5412 (N_5412,In_1168,In_2857);
or U5413 (N_5413,In_4826,In_2850);
nand U5414 (N_5414,In_4582,In_4173);
or U5415 (N_5415,In_1019,In_3939);
nor U5416 (N_5416,In_709,In_2693);
or U5417 (N_5417,In_272,In_268);
nor U5418 (N_5418,In_1935,In_2848);
xnor U5419 (N_5419,In_423,In_30);
nor U5420 (N_5420,In_2331,In_367);
or U5421 (N_5421,In_584,In_3480);
xor U5422 (N_5422,In_571,In_3026);
xor U5423 (N_5423,In_4586,In_2439);
xnor U5424 (N_5424,In_3946,In_4608);
or U5425 (N_5425,In_2339,In_580);
xor U5426 (N_5426,In_3793,In_2925);
nor U5427 (N_5427,In_2593,In_4809);
nor U5428 (N_5428,In_2681,In_2028);
xor U5429 (N_5429,In_1234,In_1649);
nand U5430 (N_5430,In_1320,In_3817);
or U5431 (N_5431,In_2938,In_3694);
xnor U5432 (N_5432,In_3418,In_4165);
nor U5433 (N_5433,In_1536,In_1447);
and U5434 (N_5434,In_1903,In_3046);
nand U5435 (N_5435,In_4462,In_2130);
nor U5436 (N_5436,In_2055,In_1837);
nand U5437 (N_5437,In_3326,In_4632);
nand U5438 (N_5438,In_2645,In_2382);
or U5439 (N_5439,In_4062,In_1195);
and U5440 (N_5440,In_1204,In_2619);
and U5441 (N_5441,In_3308,In_4677);
or U5442 (N_5442,In_4122,In_2167);
and U5443 (N_5443,In_317,In_1346);
nand U5444 (N_5444,In_2602,In_1203);
xor U5445 (N_5445,In_3454,In_1189);
xnor U5446 (N_5446,In_1250,In_4060);
nand U5447 (N_5447,In_1273,In_4917);
and U5448 (N_5448,In_2754,In_799);
nand U5449 (N_5449,In_1563,In_56);
nand U5450 (N_5450,In_1582,In_531);
and U5451 (N_5451,In_796,In_2322);
or U5452 (N_5452,In_2573,In_1721);
xnor U5453 (N_5453,In_1507,In_48);
nand U5454 (N_5454,In_1360,In_12);
xor U5455 (N_5455,In_2201,In_4340);
nand U5456 (N_5456,In_4435,In_1372);
or U5457 (N_5457,In_2316,In_4582);
nor U5458 (N_5458,In_4750,In_3426);
or U5459 (N_5459,In_1105,In_1508);
and U5460 (N_5460,In_3651,In_104);
nand U5461 (N_5461,In_3192,In_4970);
and U5462 (N_5462,In_2576,In_4111);
xor U5463 (N_5463,In_2686,In_2069);
or U5464 (N_5464,In_98,In_4191);
xnor U5465 (N_5465,In_3372,In_1369);
and U5466 (N_5466,In_1896,In_2247);
xor U5467 (N_5467,In_3749,In_2692);
or U5468 (N_5468,In_1177,In_2768);
nor U5469 (N_5469,In_4475,In_4528);
and U5470 (N_5470,In_1314,In_4562);
or U5471 (N_5471,In_1735,In_4114);
nand U5472 (N_5472,In_1430,In_3471);
nand U5473 (N_5473,In_240,In_480);
and U5474 (N_5474,In_1286,In_2319);
nor U5475 (N_5475,In_4021,In_621);
nand U5476 (N_5476,In_1971,In_1411);
or U5477 (N_5477,In_4048,In_3663);
and U5478 (N_5478,In_2220,In_2311);
xnor U5479 (N_5479,In_3980,In_2188);
nand U5480 (N_5480,In_3542,In_4156);
and U5481 (N_5481,In_1630,In_583);
xnor U5482 (N_5482,In_339,In_2463);
and U5483 (N_5483,In_4534,In_4482);
and U5484 (N_5484,In_2407,In_2701);
nand U5485 (N_5485,In_3025,In_1875);
xnor U5486 (N_5486,In_4738,In_9);
nand U5487 (N_5487,In_2022,In_2803);
nand U5488 (N_5488,In_2344,In_4835);
and U5489 (N_5489,In_4213,In_3406);
and U5490 (N_5490,In_266,In_3072);
and U5491 (N_5491,In_1428,In_4360);
nand U5492 (N_5492,In_2234,In_2861);
nand U5493 (N_5493,In_3492,In_4458);
and U5494 (N_5494,In_4820,In_2639);
nor U5495 (N_5495,In_2019,In_109);
xnor U5496 (N_5496,In_2538,In_4739);
or U5497 (N_5497,In_780,In_4073);
or U5498 (N_5498,In_2498,In_4633);
xor U5499 (N_5499,In_2264,In_4066);
nand U5500 (N_5500,In_760,In_726);
xnor U5501 (N_5501,In_4579,In_1224);
and U5502 (N_5502,In_4044,In_2950);
nand U5503 (N_5503,In_441,In_1480);
nand U5504 (N_5504,In_2843,In_1132);
xnor U5505 (N_5505,In_4269,In_4975);
nor U5506 (N_5506,In_1541,In_1502);
and U5507 (N_5507,In_3368,In_4709);
xnor U5508 (N_5508,In_4036,In_9);
or U5509 (N_5509,In_4141,In_2519);
xor U5510 (N_5510,In_1636,In_3576);
nor U5511 (N_5511,In_2421,In_4810);
nor U5512 (N_5512,In_4862,In_2076);
nand U5513 (N_5513,In_2309,In_1984);
nand U5514 (N_5514,In_3184,In_398);
or U5515 (N_5515,In_3173,In_1297);
nor U5516 (N_5516,In_4373,In_3685);
nor U5517 (N_5517,In_612,In_908);
nor U5518 (N_5518,In_2437,In_3462);
nor U5519 (N_5519,In_4294,In_154);
xnor U5520 (N_5520,In_4973,In_4657);
xnor U5521 (N_5521,In_948,In_2510);
nand U5522 (N_5522,In_4914,In_2136);
or U5523 (N_5523,In_550,In_1350);
and U5524 (N_5524,In_383,In_2008);
nor U5525 (N_5525,In_2718,In_2369);
nor U5526 (N_5526,In_2548,In_1635);
or U5527 (N_5527,In_1604,In_2751);
and U5528 (N_5528,In_3253,In_0);
xnor U5529 (N_5529,In_2698,In_3490);
nor U5530 (N_5530,In_3098,In_984);
and U5531 (N_5531,In_405,In_3047);
and U5532 (N_5532,In_3175,In_1945);
or U5533 (N_5533,In_205,In_469);
and U5534 (N_5534,In_3595,In_3533);
nand U5535 (N_5535,In_2509,In_2933);
or U5536 (N_5536,In_1838,In_3941);
nand U5537 (N_5537,In_221,In_882);
and U5538 (N_5538,In_4522,In_1240);
xor U5539 (N_5539,In_4348,In_788);
xnor U5540 (N_5540,In_4809,In_2597);
nand U5541 (N_5541,In_4699,In_2440);
nor U5542 (N_5542,In_2506,In_2555);
nand U5543 (N_5543,In_1606,In_4646);
nand U5544 (N_5544,In_2100,In_424);
nor U5545 (N_5545,In_705,In_0);
nor U5546 (N_5546,In_3482,In_3456);
xnor U5547 (N_5547,In_2408,In_4864);
xnor U5548 (N_5548,In_3957,In_2343);
or U5549 (N_5549,In_4134,In_645);
and U5550 (N_5550,In_4395,In_14);
and U5551 (N_5551,In_3636,In_2761);
or U5552 (N_5552,In_2492,In_4683);
xor U5553 (N_5553,In_3178,In_3565);
nand U5554 (N_5554,In_244,In_623);
xor U5555 (N_5555,In_4058,In_1773);
and U5556 (N_5556,In_2301,In_971);
and U5557 (N_5557,In_3519,In_4536);
or U5558 (N_5558,In_1829,In_701);
xnor U5559 (N_5559,In_4521,In_298);
nor U5560 (N_5560,In_916,In_3630);
or U5561 (N_5561,In_2356,In_1158);
nor U5562 (N_5562,In_2867,In_2676);
xnor U5563 (N_5563,In_3010,In_1828);
or U5564 (N_5564,In_1967,In_3991);
nand U5565 (N_5565,In_3231,In_396);
nand U5566 (N_5566,In_2855,In_1542);
or U5567 (N_5567,In_4908,In_1856);
or U5568 (N_5568,In_4380,In_1100);
nand U5569 (N_5569,In_3918,In_2934);
or U5570 (N_5570,In_4470,In_1054);
or U5571 (N_5571,In_2859,In_680);
nor U5572 (N_5572,In_2102,In_3377);
xor U5573 (N_5573,In_2459,In_3776);
xor U5574 (N_5574,In_1238,In_2222);
and U5575 (N_5575,In_1556,In_4465);
nor U5576 (N_5576,In_4840,In_333);
or U5577 (N_5577,In_324,In_4180);
xnor U5578 (N_5578,In_798,In_2115);
or U5579 (N_5579,In_477,In_4233);
xor U5580 (N_5580,In_3763,In_3171);
nand U5581 (N_5581,In_2440,In_4015);
and U5582 (N_5582,In_3415,In_1710);
and U5583 (N_5583,In_4932,In_3003);
nor U5584 (N_5584,In_1163,In_2500);
xnor U5585 (N_5585,In_28,In_2924);
nand U5586 (N_5586,In_683,In_3629);
and U5587 (N_5587,In_4579,In_2112);
nor U5588 (N_5588,In_1472,In_419);
nand U5589 (N_5589,In_4619,In_2561);
nand U5590 (N_5590,In_4908,In_3421);
xor U5591 (N_5591,In_2297,In_684);
and U5592 (N_5592,In_1052,In_2757);
and U5593 (N_5593,In_1866,In_1321);
nor U5594 (N_5594,In_1611,In_2456);
or U5595 (N_5595,In_1817,In_2565);
and U5596 (N_5596,In_3947,In_3250);
and U5597 (N_5597,In_900,In_3624);
and U5598 (N_5598,In_17,In_1264);
nand U5599 (N_5599,In_2885,In_3833);
xnor U5600 (N_5600,In_930,In_243);
nand U5601 (N_5601,In_2566,In_3792);
nor U5602 (N_5602,In_1245,In_295);
xor U5603 (N_5603,In_1841,In_4971);
or U5604 (N_5604,In_2779,In_484);
nand U5605 (N_5605,In_1042,In_3147);
and U5606 (N_5606,In_190,In_3545);
and U5607 (N_5607,In_2744,In_2942);
xnor U5608 (N_5608,In_2622,In_1585);
nand U5609 (N_5609,In_1034,In_4225);
nand U5610 (N_5610,In_352,In_2958);
xnor U5611 (N_5611,In_1868,In_4360);
nand U5612 (N_5612,In_3959,In_1930);
and U5613 (N_5613,In_1002,In_3254);
xnor U5614 (N_5614,In_4543,In_86);
nor U5615 (N_5615,In_2850,In_4298);
nor U5616 (N_5616,In_4254,In_2178);
and U5617 (N_5617,In_1222,In_4904);
and U5618 (N_5618,In_2391,In_4897);
nand U5619 (N_5619,In_3101,In_248);
nor U5620 (N_5620,In_4107,In_4313);
nor U5621 (N_5621,In_1254,In_2152);
nor U5622 (N_5622,In_4164,In_3921);
nand U5623 (N_5623,In_247,In_4634);
xor U5624 (N_5624,In_2345,In_4410);
xnor U5625 (N_5625,In_3901,In_862);
nor U5626 (N_5626,In_3587,In_429);
xor U5627 (N_5627,In_735,In_1679);
or U5628 (N_5628,In_4837,In_2047);
and U5629 (N_5629,In_3767,In_7);
or U5630 (N_5630,In_4312,In_3699);
or U5631 (N_5631,In_764,In_3193);
nor U5632 (N_5632,In_4806,In_4673);
nand U5633 (N_5633,In_4724,In_2285);
nand U5634 (N_5634,In_2067,In_4356);
xor U5635 (N_5635,In_1640,In_779);
nand U5636 (N_5636,In_2783,In_3503);
nor U5637 (N_5637,In_3375,In_4729);
or U5638 (N_5638,In_3745,In_3286);
or U5639 (N_5639,In_2846,In_1218);
nand U5640 (N_5640,In_1299,In_3548);
or U5641 (N_5641,In_4639,In_2084);
and U5642 (N_5642,In_1265,In_1465);
xor U5643 (N_5643,In_2772,In_1884);
nand U5644 (N_5644,In_2716,In_2912);
and U5645 (N_5645,In_422,In_2639);
and U5646 (N_5646,In_888,In_1609);
nor U5647 (N_5647,In_1372,In_2037);
nor U5648 (N_5648,In_3563,In_3837);
xor U5649 (N_5649,In_2108,In_1824);
nor U5650 (N_5650,In_1290,In_2268);
and U5651 (N_5651,In_349,In_865);
nor U5652 (N_5652,In_4410,In_3363);
and U5653 (N_5653,In_4259,In_4765);
and U5654 (N_5654,In_3582,In_224);
and U5655 (N_5655,In_2640,In_1579);
nor U5656 (N_5656,In_1291,In_2338);
and U5657 (N_5657,In_4858,In_2256);
and U5658 (N_5658,In_2458,In_2434);
and U5659 (N_5659,In_3592,In_3799);
nand U5660 (N_5660,In_3467,In_443);
or U5661 (N_5661,In_2785,In_3057);
or U5662 (N_5662,In_2708,In_3293);
nor U5663 (N_5663,In_363,In_282);
and U5664 (N_5664,In_4698,In_4392);
nand U5665 (N_5665,In_4904,In_1331);
or U5666 (N_5666,In_2081,In_2528);
nand U5667 (N_5667,In_3727,In_745);
and U5668 (N_5668,In_611,In_3885);
nand U5669 (N_5669,In_25,In_2242);
xor U5670 (N_5670,In_4239,In_372);
nand U5671 (N_5671,In_4753,In_46);
xnor U5672 (N_5672,In_551,In_3954);
nand U5673 (N_5673,In_3509,In_1968);
xnor U5674 (N_5674,In_1614,In_945);
nor U5675 (N_5675,In_98,In_4730);
xnor U5676 (N_5676,In_3271,In_3150);
and U5677 (N_5677,In_2958,In_1284);
nand U5678 (N_5678,In_450,In_4198);
nand U5679 (N_5679,In_3870,In_3203);
and U5680 (N_5680,In_4141,In_2315);
and U5681 (N_5681,In_665,In_3289);
or U5682 (N_5682,In_1869,In_1167);
xnor U5683 (N_5683,In_1902,In_188);
or U5684 (N_5684,In_2617,In_3448);
nor U5685 (N_5685,In_1480,In_2738);
xnor U5686 (N_5686,In_2252,In_4574);
nand U5687 (N_5687,In_3977,In_3871);
xnor U5688 (N_5688,In_2226,In_4203);
xor U5689 (N_5689,In_3819,In_4435);
or U5690 (N_5690,In_2294,In_2084);
nand U5691 (N_5691,In_3753,In_671);
or U5692 (N_5692,In_4000,In_4945);
xnor U5693 (N_5693,In_4081,In_4335);
nor U5694 (N_5694,In_3507,In_1094);
or U5695 (N_5695,In_2894,In_18);
and U5696 (N_5696,In_3820,In_3543);
or U5697 (N_5697,In_1548,In_4333);
nand U5698 (N_5698,In_3904,In_824);
nor U5699 (N_5699,In_1329,In_2821);
nand U5700 (N_5700,In_4871,In_4007);
nor U5701 (N_5701,In_3650,In_3821);
xnor U5702 (N_5702,In_1202,In_2119);
xnor U5703 (N_5703,In_3761,In_4694);
xnor U5704 (N_5704,In_3131,In_4926);
nor U5705 (N_5705,In_3420,In_4988);
nor U5706 (N_5706,In_819,In_3106);
or U5707 (N_5707,In_4427,In_3764);
xor U5708 (N_5708,In_3851,In_4361);
and U5709 (N_5709,In_2916,In_2881);
nand U5710 (N_5710,In_636,In_569);
nand U5711 (N_5711,In_2253,In_3161);
or U5712 (N_5712,In_2713,In_118);
nor U5713 (N_5713,In_4497,In_3929);
nor U5714 (N_5714,In_3345,In_803);
xor U5715 (N_5715,In_4984,In_4703);
xnor U5716 (N_5716,In_1510,In_3882);
or U5717 (N_5717,In_2360,In_3781);
and U5718 (N_5718,In_3270,In_657);
xor U5719 (N_5719,In_611,In_3461);
and U5720 (N_5720,In_3621,In_2032);
or U5721 (N_5721,In_3822,In_3838);
nor U5722 (N_5722,In_1754,In_3271);
xor U5723 (N_5723,In_4898,In_2884);
nor U5724 (N_5724,In_2063,In_351);
nor U5725 (N_5725,In_6,In_687);
nand U5726 (N_5726,In_2198,In_2693);
nor U5727 (N_5727,In_3446,In_402);
xnor U5728 (N_5728,In_3409,In_3289);
nand U5729 (N_5729,In_4127,In_840);
and U5730 (N_5730,In_2969,In_2413);
and U5731 (N_5731,In_3386,In_4644);
and U5732 (N_5732,In_3401,In_2759);
and U5733 (N_5733,In_1748,In_2915);
or U5734 (N_5734,In_1844,In_4876);
nand U5735 (N_5735,In_353,In_2639);
xor U5736 (N_5736,In_2627,In_3974);
nand U5737 (N_5737,In_850,In_1604);
nand U5738 (N_5738,In_2328,In_4914);
xnor U5739 (N_5739,In_2876,In_2512);
nor U5740 (N_5740,In_2204,In_1017);
nand U5741 (N_5741,In_205,In_679);
nor U5742 (N_5742,In_4298,In_2847);
or U5743 (N_5743,In_1943,In_3676);
nand U5744 (N_5744,In_3924,In_3373);
xnor U5745 (N_5745,In_2312,In_425);
nand U5746 (N_5746,In_4393,In_3625);
xnor U5747 (N_5747,In_4820,In_1909);
nor U5748 (N_5748,In_4949,In_921);
nor U5749 (N_5749,In_3401,In_1022);
xor U5750 (N_5750,In_2904,In_696);
and U5751 (N_5751,In_2412,In_3193);
or U5752 (N_5752,In_2754,In_2057);
xor U5753 (N_5753,In_526,In_2413);
xor U5754 (N_5754,In_193,In_3963);
or U5755 (N_5755,In_4344,In_1355);
nand U5756 (N_5756,In_3724,In_3775);
and U5757 (N_5757,In_4771,In_4001);
xnor U5758 (N_5758,In_3683,In_2764);
or U5759 (N_5759,In_1731,In_4823);
xnor U5760 (N_5760,In_2424,In_1207);
or U5761 (N_5761,In_632,In_1644);
nor U5762 (N_5762,In_2185,In_3316);
and U5763 (N_5763,In_2615,In_4020);
and U5764 (N_5764,In_2326,In_4323);
nand U5765 (N_5765,In_4624,In_4976);
or U5766 (N_5766,In_3347,In_1780);
or U5767 (N_5767,In_508,In_3529);
xnor U5768 (N_5768,In_3149,In_4067);
xnor U5769 (N_5769,In_561,In_3211);
xnor U5770 (N_5770,In_3533,In_4483);
nor U5771 (N_5771,In_3386,In_18);
nand U5772 (N_5772,In_3537,In_3310);
xor U5773 (N_5773,In_1965,In_2979);
nor U5774 (N_5774,In_3379,In_3212);
xnor U5775 (N_5775,In_1840,In_945);
and U5776 (N_5776,In_3527,In_2959);
xor U5777 (N_5777,In_4254,In_4703);
nor U5778 (N_5778,In_2523,In_257);
nand U5779 (N_5779,In_3602,In_4136);
xnor U5780 (N_5780,In_2880,In_608);
and U5781 (N_5781,In_3669,In_2448);
nor U5782 (N_5782,In_1448,In_2473);
xnor U5783 (N_5783,In_2921,In_685);
and U5784 (N_5784,In_80,In_596);
and U5785 (N_5785,In_4298,In_76);
and U5786 (N_5786,In_925,In_2376);
nor U5787 (N_5787,In_1072,In_773);
xnor U5788 (N_5788,In_1001,In_1820);
nand U5789 (N_5789,In_2656,In_3933);
or U5790 (N_5790,In_4826,In_4159);
xnor U5791 (N_5791,In_3611,In_3053);
nand U5792 (N_5792,In_4728,In_1951);
and U5793 (N_5793,In_2195,In_3914);
xnor U5794 (N_5794,In_727,In_3378);
nand U5795 (N_5795,In_4239,In_1841);
nand U5796 (N_5796,In_3330,In_134);
or U5797 (N_5797,In_4695,In_4607);
xor U5798 (N_5798,In_3911,In_992);
and U5799 (N_5799,In_211,In_3914);
nand U5800 (N_5800,In_2897,In_2570);
nand U5801 (N_5801,In_4659,In_1102);
nor U5802 (N_5802,In_1797,In_3414);
nor U5803 (N_5803,In_1521,In_35);
nor U5804 (N_5804,In_959,In_3095);
or U5805 (N_5805,In_683,In_3969);
xor U5806 (N_5806,In_194,In_2290);
xor U5807 (N_5807,In_4213,In_4215);
nor U5808 (N_5808,In_972,In_4393);
nand U5809 (N_5809,In_4524,In_439);
nand U5810 (N_5810,In_555,In_2419);
xor U5811 (N_5811,In_2645,In_547);
xnor U5812 (N_5812,In_3211,In_3637);
xnor U5813 (N_5813,In_2069,In_2993);
or U5814 (N_5814,In_960,In_4236);
nand U5815 (N_5815,In_4989,In_703);
nand U5816 (N_5816,In_4104,In_4721);
or U5817 (N_5817,In_3379,In_1066);
or U5818 (N_5818,In_2159,In_801);
or U5819 (N_5819,In_54,In_593);
nand U5820 (N_5820,In_2465,In_3975);
or U5821 (N_5821,In_1288,In_4803);
nor U5822 (N_5822,In_971,In_2207);
xor U5823 (N_5823,In_2873,In_2961);
nor U5824 (N_5824,In_2118,In_1671);
xnor U5825 (N_5825,In_2548,In_3223);
nor U5826 (N_5826,In_2435,In_3992);
and U5827 (N_5827,In_1646,In_4578);
and U5828 (N_5828,In_4453,In_4113);
and U5829 (N_5829,In_1787,In_321);
nor U5830 (N_5830,In_4794,In_4736);
and U5831 (N_5831,In_1213,In_3203);
and U5832 (N_5832,In_816,In_2430);
nor U5833 (N_5833,In_2921,In_3486);
nor U5834 (N_5834,In_351,In_2279);
and U5835 (N_5835,In_3518,In_3414);
nand U5836 (N_5836,In_4491,In_2564);
nand U5837 (N_5837,In_3017,In_3003);
and U5838 (N_5838,In_3873,In_2063);
or U5839 (N_5839,In_611,In_201);
nand U5840 (N_5840,In_3561,In_2793);
and U5841 (N_5841,In_2888,In_1808);
nor U5842 (N_5842,In_4878,In_73);
nor U5843 (N_5843,In_1756,In_3414);
nor U5844 (N_5844,In_1221,In_4140);
and U5845 (N_5845,In_4613,In_2254);
nand U5846 (N_5846,In_3484,In_3905);
nor U5847 (N_5847,In_4739,In_221);
or U5848 (N_5848,In_4771,In_3633);
nand U5849 (N_5849,In_637,In_4740);
and U5850 (N_5850,In_2710,In_4077);
nor U5851 (N_5851,In_2904,In_1480);
nor U5852 (N_5852,In_251,In_4685);
or U5853 (N_5853,In_4604,In_3510);
nor U5854 (N_5854,In_1792,In_729);
xnor U5855 (N_5855,In_4068,In_2427);
nand U5856 (N_5856,In_1435,In_4402);
and U5857 (N_5857,In_2263,In_2179);
nand U5858 (N_5858,In_709,In_1348);
or U5859 (N_5859,In_2444,In_4464);
nand U5860 (N_5860,In_2473,In_3979);
xor U5861 (N_5861,In_1688,In_4347);
or U5862 (N_5862,In_1656,In_3610);
nor U5863 (N_5863,In_136,In_2132);
nand U5864 (N_5864,In_4093,In_1973);
nor U5865 (N_5865,In_2232,In_1270);
or U5866 (N_5866,In_3666,In_1575);
nand U5867 (N_5867,In_3777,In_4625);
and U5868 (N_5868,In_3580,In_1529);
xor U5869 (N_5869,In_793,In_2109);
and U5870 (N_5870,In_3442,In_2321);
or U5871 (N_5871,In_1082,In_1806);
nand U5872 (N_5872,In_4981,In_3741);
and U5873 (N_5873,In_474,In_3967);
and U5874 (N_5874,In_795,In_2694);
nand U5875 (N_5875,In_4691,In_4763);
xor U5876 (N_5876,In_4736,In_2720);
xor U5877 (N_5877,In_4766,In_692);
xor U5878 (N_5878,In_3218,In_4417);
and U5879 (N_5879,In_65,In_1647);
or U5880 (N_5880,In_2273,In_1772);
xor U5881 (N_5881,In_2548,In_461);
xnor U5882 (N_5882,In_1216,In_2624);
xor U5883 (N_5883,In_2926,In_2127);
xor U5884 (N_5884,In_2252,In_3139);
and U5885 (N_5885,In_2616,In_4320);
nor U5886 (N_5886,In_100,In_1361);
or U5887 (N_5887,In_2018,In_4953);
nor U5888 (N_5888,In_2404,In_2242);
nand U5889 (N_5889,In_4901,In_3034);
nand U5890 (N_5890,In_2116,In_473);
nor U5891 (N_5891,In_2663,In_3049);
or U5892 (N_5892,In_4537,In_3967);
xor U5893 (N_5893,In_3179,In_1871);
or U5894 (N_5894,In_2846,In_717);
and U5895 (N_5895,In_3391,In_3087);
nand U5896 (N_5896,In_3446,In_4004);
and U5897 (N_5897,In_2828,In_4189);
or U5898 (N_5898,In_4730,In_3604);
nand U5899 (N_5899,In_2447,In_1405);
xnor U5900 (N_5900,In_4281,In_224);
nor U5901 (N_5901,In_2666,In_2228);
xnor U5902 (N_5902,In_3120,In_81);
xnor U5903 (N_5903,In_4639,In_4345);
and U5904 (N_5904,In_4663,In_6);
and U5905 (N_5905,In_4187,In_2953);
nand U5906 (N_5906,In_2621,In_1807);
nand U5907 (N_5907,In_1090,In_707);
nor U5908 (N_5908,In_3557,In_2569);
nand U5909 (N_5909,In_1926,In_171);
nand U5910 (N_5910,In_2433,In_3910);
nor U5911 (N_5911,In_4819,In_3000);
or U5912 (N_5912,In_3125,In_3198);
nand U5913 (N_5913,In_460,In_2273);
xor U5914 (N_5914,In_3638,In_948);
xor U5915 (N_5915,In_2471,In_1489);
xnor U5916 (N_5916,In_2278,In_1399);
nor U5917 (N_5917,In_3856,In_2065);
nor U5918 (N_5918,In_2360,In_64);
nand U5919 (N_5919,In_4093,In_4480);
and U5920 (N_5920,In_3431,In_4176);
xor U5921 (N_5921,In_2336,In_2498);
and U5922 (N_5922,In_2238,In_2431);
nor U5923 (N_5923,In_1847,In_472);
xnor U5924 (N_5924,In_167,In_2271);
nor U5925 (N_5925,In_4191,In_1890);
nor U5926 (N_5926,In_4594,In_3388);
nor U5927 (N_5927,In_4019,In_3966);
xor U5928 (N_5928,In_1331,In_1757);
and U5929 (N_5929,In_4442,In_1472);
xnor U5930 (N_5930,In_425,In_3175);
nor U5931 (N_5931,In_2451,In_631);
xor U5932 (N_5932,In_1280,In_4985);
and U5933 (N_5933,In_3508,In_3523);
or U5934 (N_5934,In_2434,In_1797);
xnor U5935 (N_5935,In_120,In_1131);
and U5936 (N_5936,In_4947,In_2188);
and U5937 (N_5937,In_1317,In_576);
nand U5938 (N_5938,In_4559,In_3853);
or U5939 (N_5939,In_962,In_3363);
and U5940 (N_5940,In_4094,In_454);
or U5941 (N_5941,In_4844,In_4096);
xor U5942 (N_5942,In_4414,In_1235);
or U5943 (N_5943,In_1195,In_338);
or U5944 (N_5944,In_175,In_3567);
nor U5945 (N_5945,In_1988,In_4140);
xnor U5946 (N_5946,In_4054,In_3810);
and U5947 (N_5947,In_1010,In_1812);
nand U5948 (N_5948,In_2496,In_181);
and U5949 (N_5949,In_3094,In_2234);
or U5950 (N_5950,In_852,In_40);
nand U5951 (N_5951,In_1635,In_4443);
xor U5952 (N_5952,In_4264,In_4301);
xnor U5953 (N_5953,In_2013,In_3503);
nand U5954 (N_5954,In_4033,In_2264);
and U5955 (N_5955,In_1450,In_2626);
and U5956 (N_5956,In_2509,In_4718);
xnor U5957 (N_5957,In_53,In_3169);
xnor U5958 (N_5958,In_4890,In_994);
or U5959 (N_5959,In_528,In_2022);
and U5960 (N_5960,In_1539,In_1603);
nor U5961 (N_5961,In_2120,In_351);
and U5962 (N_5962,In_1963,In_1766);
nand U5963 (N_5963,In_4385,In_532);
and U5964 (N_5964,In_1990,In_2734);
and U5965 (N_5965,In_2201,In_4176);
and U5966 (N_5966,In_69,In_4878);
nand U5967 (N_5967,In_2316,In_3313);
nor U5968 (N_5968,In_165,In_455);
xnor U5969 (N_5969,In_2615,In_1531);
nand U5970 (N_5970,In_4769,In_815);
nor U5971 (N_5971,In_1496,In_2396);
and U5972 (N_5972,In_3651,In_3495);
xor U5973 (N_5973,In_2323,In_4619);
nor U5974 (N_5974,In_3955,In_979);
nand U5975 (N_5975,In_2416,In_1615);
nand U5976 (N_5976,In_3731,In_4928);
or U5977 (N_5977,In_1852,In_3039);
or U5978 (N_5978,In_1010,In_733);
nor U5979 (N_5979,In_3437,In_877);
nand U5980 (N_5980,In_2295,In_364);
nor U5981 (N_5981,In_1826,In_2835);
nand U5982 (N_5982,In_327,In_698);
nor U5983 (N_5983,In_4402,In_4745);
or U5984 (N_5984,In_3428,In_1588);
xor U5985 (N_5985,In_208,In_4480);
nor U5986 (N_5986,In_3116,In_2878);
xor U5987 (N_5987,In_4301,In_3074);
nand U5988 (N_5988,In_610,In_4263);
or U5989 (N_5989,In_4950,In_4367);
nand U5990 (N_5990,In_2693,In_4638);
and U5991 (N_5991,In_669,In_4065);
xor U5992 (N_5992,In_3035,In_1574);
nand U5993 (N_5993,In_464,In_3959);
nand U5994 (N_5994,In_3499,In_3526);
or U5995 (N_5995,In_1564,In_3763);
and U5996 (N_5996,In_2895,In_2894);
or U5997 (N_5997,In_2813,In_2141);
nor U5998 (N_5998,In_3375,In_1785);
nand U5999 (N_5999,In_1849,In_3473);
or U6000 (N_6000,In_857,In_4592);
nor U6001 (N_6001,In_1844,In_3787);
xor U6002 (N_6002,In_4723,In_1217);
nor U6003 (N_6003,In_1390,In_2112);
or U6004 (N_6004,In_4528,In_4370);
nand U6005 (N_6005,In_3202,In_687);
and U6006 (N_6006,In_2050,In_3476);
nand U6007 (N_6007,In_2785,In_3769);
nor U6008 (N_6008,In_3160,In_3252);
xnor U6009 (N_6009,In_41,In_4776);
and U6010 (N_6010,In_2326,In_256);
and U6011 (N_6011,In_3550,In_4295);
xor U6012 (N_6012,In_2462,In_2414);
xnor U6013 (N_6013,In_815,In_3716);
nor U6014 (N_6014,In_4623,In_3209);
nor U6015 (N_6015,In_2386,In_1562);
or U6016 (N_6016,In_1862,In_538);
or U6017 (N_6017,In_3977,In_2496);
xnor U6018 (N_6018,In_823,In_4930);
nor U6019 (N_6019,In_2178,In_2946);
nand U6020 (N_6020,In_2618,In_820);
or U6021 (N_6021,In_2173,In_4505);
nor U6022 (N_6022,In_649,In_2181);
and U6023 (N_6023,In_4192,In_1387);
or U6024 (N_6024,In_2332,In_957);
or U6025 (N_6025,In_3615,In_1676);
and U6026 (N_6026,In_2311,In_2481);
or U6027 (N_6027,In_1324,In_3335);
and U6028 (N_6028,In_3051,In_2402);
or U6029 (N_6029,In_3628,In_1473);
nor U6030 (N_6030,In_666,In_841);
nor U6031 (N_6031,In_4779,In_1055);
nand U6032 (N_6032,In_4229,In_2016);
nor U6033 (N_6033,In_3118,In_4936);
xor U6034 (N_6034,In_2644,In_2716);
nand U6035 (N_6035,In_4402,In_2343);
xor U6036 (N_6036,In_4650,In_4940);
xnor U6037 (N_6037,In_1192,In_1139);
nor U6038 (N_6038,In_4059,In_1056);
nor U6039 (N_6039,In_3533,In_623);
nor U6040 (N_6040,In_3360,In_2969);
and U6041 (N_6041,In_1640,In_4183);
nand U6042 (N_6042,In_4473,In_3329);
nand U6043 (N_6043,In_4533,In_4968);
or U6044 (N_6044,In_4677,In_2789);
nor U6045 (N_6045,In_555,In_3365);
or U6046 (N_6046,In_2805,In_1317);
or U6047 (N_6047,In_3392,In_1625);
nor U6048 (N_6048,In_968,In_2498);
xnor U6049 (N_6049,In_4015,In_485);
xnor U6050 (N_6050,In_1210,In_498);
xor U6051 (N_6051,In_4506,In_3326);
nor U6052 (N_6052,In_3059,In_3134);
or U6053 (N_6053,In_1266,In_4266);
xnor U6054 (N_6054,In_487,In_462);
or U6055 (N_6055,In_136,In_3165);
xnor U6056 (N_6056,In_2020,In_889);
or U6057 (N_6057,In_1568,In_1727);
xnor U6058 (N_6058,In_2994,In_2289);
and U6059 (N_6059,In_2835,In_4405);
xnor U6060 (N_6060,In_3102,In_2871);
and U6061 (N_6061,In_3702,In_2309);
xnor U6062 (N_6062,In_1587,In_1287);
xnor U6063 (N_6063,In_1383,In_862);
nand U6064 (N_6064,In_963,In_977);
or U6065 (N_6065,In_4531,In_3666);
or U6066 (N_6066,In_1801,In_2422);
nand U6067 (N_6067,In_2363,In_3421);
nand U6068 (N_6068,In_4108,In_750);
or U6069 (N_6069,In_3442,In_3042);
or U6070 (N_6070,In_4704,In_1208);
xor U6071 (N_6071,In_3100,In_1875);
or U6072 (N_6072,In_2257,In_2098);
or U6073 (N_6073,In_2681,In_2498);
and U6074 (N_6074,In_3693,In_157);
and U6075 (N_6075,In_4401,In_1877);
and U6076 (N_6076,In_1188,In_3647);
xor U6077 (N_6077,In_2991,In_3677);
xor U6078 (N_6078,In_281,In_1175);
nand U6079 (N_6079,In_4814,In_940);
xor U6080 (N_6080,In_4963,In_2506);
and U6081 (N_6081,In_4700,In_2538);
or U6082 (N_6082,In_1092,In_3207);
nand U6083 (N_6083,In_992,In_2060);
nor U6084 (N_6084,In_3574,In_4706);
nor U6085 (N_6085,In_2944,In_3971);
nor U6086 (N_6086,In_727,In_2931);
and U6087 (N_6087,In_1941,In_4067);
or U6088 (N_6088,In_2294,In_1597);
nor U6089 (N_6089,In_4328,In_3741);
or U6090 (N_6090,In_2048,In_2053);
nor U6091 (N_6091,In_2527,In_3927);
and U6092 (N_6092,In_2069,In_2798);
or U6093 (N_6093,In_518,In_3474);
and U6094 (N_6094,In_1160,In_2419);
nor U6095 (N_6095,In_3103,In_2257);
xor U6096 (N_6096,In_3846,In_846);
and U6097 (N_6097,In_1109,In_2217);
and U6098 (N_6098,In_1503,In_4803);
nor U6099 (N_6099,In_1056,In_3183);
nor U6100 (N_6100,In_2470,In_917);
nor U6101 (N_6101,In_2861,In_2954);
nor U6102 (N_6102,In_4609,In_4983);
nand U6103 (N_6103,In_4772,In_4860);
nand U6104 (N_6104,In_4553,In_969);
nor U6105 (N_6105,In_4306,In_2251);
and U6106 (N_6106,In_2439,In_1122);
or U6107 (N_6107,In_347,In_314);
and U6108 (N_6108,In_2944,In_1060);
nand U6109 (N_6109,In_4475,In_2951);
and U6110 (N_6110,In_4114,In_3502);
or U6111 (N_6111,In_4539,In_4731);
nor U6112 (N_6112,In_3901,In_1174);
nor U6113 (N_6113,In_2711,In_2501);
xnor U6114 (N_6114,In_2830,In_3187);
and U6115 (N_6115,In_1956,In_2227);
nand U6116 (N_6116,In_3953,In_3884);
nor U6117 (N_6117,In_2402,In_2720);
nor U6118 (N_6118,In_2850,In_4532);
xor U6119 (N_6119,In_678,In_1887);
or U6120 (N_6120,In_3381,In_2728);
nor U6121 (N_6121,In_3241,In_283);
and U6122 (N_6122,In_3795,In_18);
nand U6123 (N_6123,In_3379,In_3681);
xor U6124 (N_6124,In_3322,In_695);
xor U6125 (N_6125,In_3876,In_3051);
nand U6126 (N_6126,In_3290,In_543);
nor U6127 (N_6127,In_940,In_2217);
xnor U6128 (N_6128,In_1711,In_4548);
and U6129 (N_6129,In_119,In_2283);
and U6130 (N_6130,In_3451,In_2001);
nor U6131 (N_6131,In_3698,In_4502);
and U6132 (N_6132,In_3835,In_399);
xnor U6133 (N_6133,In_718,In_1175);
xor U6134 (N_6134,In_2834,In_4721);
and U6135 (N_6135,In_349,In_4966);
and U6136 (N_6136,In_1051,In_1109);
or U6137 (N_6137,In_136,In_1849);
nand U6138 (N_6138,In_625,In_439);
or U6139 (N_6139,In_975,In_4175);
or U6140 (N_6140,In_1638,In_2201);
nand U6141 (N_6141,In_1411,In_21);
or U6142 (N_6142,In_3542,In_531);
nand U6143 (N_6143,In_2243,In_3683);
nand U6144 (N_6144,In_979,In_2194);
nor U6145 (N_6145,In_4373,In_1446);
nand U6146 (N_6146,In_4923,In_813);
and U6147 (N_6147,In_3328,In_1364);
nand U6148 (N_6148,In_3986,In_1252);
xnor U6149 (N_6149,In_2282,In_2247);
or U6150 (N_6150,In_775,In_4197);
nand U6151 (N_6151,In_4557,In_1000);
or U6152 (N_6152,In_242,In_3188);
xor U6153 (N_6153,In_2680,In_2199);
nand U6154 (N_6154,In_2340,In_3728);
or U6155 (N_6155,In_2100,In_2845);
or U6156 (N_6156,In_3252,In_4701);
nor U6157 (N_6157,In_2886,In_1900);
or U6158 (N_6158,In_1366,In_2344);
nor U6159 (N_6159,In_2104,In_4768);
xor U6160 (N_6160,In_3443,In_3020);
and U6161 (N_6161,In_3087,In_4651);
nor U6162 (N_6162,In_1271,In_698);
nand U6163 (N_6163,In_4239,In_2430);
xnor U6164 (N_6164,In_2581,In_3233);
xnor U6165 (N_6165,In_3129,In_2974);
nor U6166 (N_6166,In_1451,In_3398);
or U6167 (N_6167,In_4918,In_3887);
or U6168 (N_6168,In_1017,In_1064);
nor U6169 (N_6169,In_3290,In_1441);
xnor U6170 (N_6170,In_358,In_547);
xor U6171 (N_6171,In_715,In_2692);
and U6172 (N_6172,In_2304,In_2041);
or U6173 (N_6173,In_268,In_541);
or U6174 (N_6174,In_1926,In_2651);
xnor U6175 (N_6175,In_3689,In_1973);
nor U6176 (N_6176,In_1891,In_4611);
xnor U6177 (N_6177,In_3883,In_4192);
and U6178 (N_6178,In_2044,In_1516);
xnor U6179 (N_6179,In_2048,In_2013);
and U6180 (N_6180,In_3113,In_2182);
xnor U6181 (N_6181,In_4479,In_3231);
xor U6182 (N_6182,In_1545,In_3087);
or U6183 (N_6183,In_1398,In_4547);
nand U6184 (N_6184,In_3921,In_4784);
xor U6185 (N_6185,In_4012,In_1732);
nor U6186 (N_6186,In_3405,In_1552);
nand U6187 (N_6187,In_1000,In_3192);
nor U6188 (N_6188,In_3782,In_726);
and U6189 (N_6189,In_4664,In_3371);
nand U6190 (N_6190,In_1874,In_321);
or U6191 (N_6191,In_4305,In_1530);
or U6192 (N_6192,In_2102,In_4543);
and U6193 (N_6193,In_3568,In_2551);
nor U6194 (N_6194,In_1661,In_2704);
nand U6195 (N_6195,In_1894,In_3826);
xnor U6196 (N_6196,In_417,In_930);
and U6197 (N_6197,In_1292,In_379);
and U6198 (N_6198,In_1518,In_3451);
nor U6199 (N_6199,In_4898,In_4757);
or U6200 (N_6200,In_4085,In_1679);
and U6201 (N_6201,In_1602,In_2740);
xnor U6202 (N_6202,In_4720,In_808);
and U6203 (N_6203,In_1024,In_4930);
nand U6204 (N_6204,In_4389,In_2242);
nor U6205 (N_6205,In_521,In_2629);
nand U6206 (N_6206,In_4225,In_4316);
nand U6207 (N_6207,In_752,In_3749);
nand U6208 (N_6208,In_4438,In_117);
or U6209 (N_6209,In_2054,In_232);
or U6210 (N_6210,In_2604,In_2801);
and U6211 (N_6211,In_2271,In_3169);
xor U6212 (N_6212,In_138,In_2154);
xnor U6213 (N_6213,In_4806,In_3057);
nand U6214 (N_6214,In_841,In_2790);
nand U6215 (N_6215,In_4682,In_759);
or U6216 (N_6216,In_914,In_1840);
nor U6217 (N_6217,In_2309,In_1976);
or U6218 (N_6218,In_3776,In_3918);
and U6219 (N_6219,In_1949,In_2334);
nor U6220 (N_6220,In_1885,In_3338);
and U6221 (N_6221,In_4053,In_1254);
nand U6222 (N_6222,In_1306,In_1128);
and U6223 (N_6223,In_3814,In_1238);
and U6224 (N_6224,In_2174,In_812);
or U6225 (N_6225,In_3653,In_3392);
nor U6226 (N_6226,In_4422,In_806);
xnor U6227 (N_6227,In_4277,In_2095);
nor U6228 (N_6228,In_2051,In_3007);
nor U6229 (N_6229,In_4539,In_2461);
nand U6230 (N_6230,In_4754,In_4314);
nand U6231 (N_6231,In_803,In_3323);
or U6232 (N_6232,In_3498,In_3765);
and U6233 (N_6233,In_3831,In_3654);
xor U6234 (N_6234,In_1330,In_547);
and U6235 (N_6235,In_1695,In_1601);
nand U6236 (N_6236,In_1092,In_4510);
and U6237 (N_6237,In_512,In_82);
nand U6238 (N_6238,In_499,In_655);
and U6239 (N_6239,In_592,In_902);
nor U6240 (N_6240,In_4277,In_4287);
nand U6241 (N_6241,In_1047,In_730);
xor U6242 (N_6242,In_4709,In_4849);
xor U6243 (N_6243,In_2899,In_3074);
and U6244 (N_6244,In_444,In_3851);
and U6245 (N_6245,In_2519,In_4308);
nand U6246 (N_6246,In_3074,In_2094);
nor U6247 (N_6247,In_3707,In_471);
nand U6248 (N_6248,In_4293,In_3279);
nand U6249 (N_6249,In_2209,In_4839);
nand U6250 (N_6250,In_4933,In_2878);
xor U6251 (N_6251,In_3317,In_2601);
nand U6252 (N_6252,In_1801,In_548);
and U6253 (N_6253,In_2055,In_441);
and U6254 (N_6254,In_1239,In_1663);
or U6255 (N_6255,In_1253,In_4253);
and U6256 (N_6256,In_874,In_4825);
xnor U6257 (N_6257,In_2822,In_4761);
nand U6258 (N_6258,In_547,In_3819);
and U6259 (N_6259,In_4218,In_2058);
nor U6260 (N_6260,In_326,In_4801);
xnor U6261 (N_6261,In_122,In_3658);
or U6262 (N_6262,In_3880,In_2595);
and U6263 (N_6263,In_729,In_2437);
and U6264 (N_6264,In_4196,In_345);
and U6265 (N_6265,In_682,In_3423);
xor U6266 (N_6266,In_1034,In_4956);
nand U6267 (N_6267,In_158,In_18);
nand U6268 (N_6268,In_2177,In_507);
nand U6269 (N_6269,In_1195,In_3823);
nand U6270 (N_6270,In_3915,In_4519);
nand U6271 (N_6271,In_884,In_749);
xor U6272 (N_6272,In_4503,In_4731);
xor U6273 (N_6273,In_240,In_1598);
or U6274 (N_6274,In_3594,In_4550);
xnor U6275 (N_6275,In_4267,In_2962);
or U6276 (N_6276,In_2783,In_1104);
or U6277 (N_6277,In_3056,In_1716);
nor U6278 (N_6278,In_2831,In_4398);
nand U6279 (N_6279,In_4485,In_285);
nand U6280 (N_6280,In_3236,In_4511);
or U6281 (N_6281,In_3847,In_3174);
xnor U6282 (N_6282,In_3761,In_1430);
nor U6283 (N_6283,In_2018,In_4955);
xnor U6284 (N_6284,In_3203,In_3654);
nand U6285 (N_6285,In_4549,In_438);
nand U6286 (N_6286,In_2903,In_4074);
nand U6287 (N_6287,In_2166,In_1906);
xor U6288 (N_6288,In_3185,In_2102);
xnor U6289 (N_6289,In_2215,In_395);
nor U6290 (N_6290,In_106,In_334);
nand U6291 (N_6291,In_2523,In_1155);
xnor U6292 (N_6292,In_3192,In_654);
nand U6293 (N_6293,In_3830,In_1771);
and U6294 (N_6294,In_566,In_3642);
xor U6295 (N_6295,In_531,In_1037);
and U6296 (N_6296,In_499,In_4226);
or U6297 (N_6297,In_4162,In_4897);
or U6298 (N_6298,In_2619,In_1196);
and U6299 (N_6299,In_4754,In_2364);
xnor U6300 (N_6300,In_4753,In_2364);
and U6301 (N_6301,In_897,In_1083);
nand U6302 (N_6302,In_3479,In_205);
and U6303 (N_6303,In_3711,In_4265);
and U6304 (N_6304,In_3808,In_4614);
xor U6305 (N_6305,In_1485,In_3297);
xnor U6306 (N_6306,In_3126,In_885);
xor U6307 (N_6307,In_2084,In_4324);
nand U6308 (N_6308,In_664,In_428);
nor U6309 (N_6309,In_4801,In_3630);
nand U6310 (N_6310,In_3645,In_278);
nor U6311 (N_6311,In_1324,In_218);
nor U6312 (N_6312,In_3448,In_4544);
or U6313 (N_6313,In_2427,In_3185);
nand U6314 (N_6314,In_877,In_914);
xor U6315 (N_6315,In_1726,In_1555);
nor U6316 (N_6316,In_4848,In_2265);
nor U6317 (N_6317,In_610,In_4047);
xnor U6318 (N_6318,In_902,In_1308);
or U6319 (N_6319,In_2514,In_3813);
nor U6320 (N_6320,In_4295,In_1181);
and U6321 (N_6321,In_262,In_1729);
nor U6322 (N_6322,In_1623,In_2583);
and U6323 (N_6323,In_4413,In_2758);
or U6324 (N_6324,In_1145,In_2175);
or U6325 (N_6325,In_4066,In_455);
nor U6326 (N_6326,In_3520,In_4242);
and U6327 (N_6327,In_3312,In_37);
nand U6328 (N_6328,In_4070,In_4139);
nand U6329 (N_6329,In_1039,In_2260);
and U6330 (N_6330,In_3619,In_1738);
and U6331 (N_6331,In_2088,In_4594);
nand U6332 (N_6332,In_115,In_761);
nor U6333 (N_6333,In_3626,In_2984);
xor U6334 (N_6334,In_617,In_4413);
nand U6335 (N_6335,In_3851,In_2594);
and U6336 (N_6336,In_3505,In_888);
nor U6337 (N_6337,In_3928,In_338);
xnor U6338 (N_6338,In_3901,In_559);
nor U6339 (N_6339,In_898,In_2052);
and U6340 (N_6340,In_2020,In_241);
and U6341 (N_6341,In_3785,In_3348);
nor U6342 (N_6342,In_4895,In_4986);
and U6343 (N_6343,In_1655,In_2687);
xor U6344 (N_6344,In_2623,In_3560);
xnor U6345 (N_6345,In_2067,In_859);
nor U6346 (N_6346,In_3889,In_530);
xor U6347 (N_6347,In_3945,In_222);
nor U6348 (N_6348,In_3736,In_501);
nand U6349 (N_6349,In_439,In_2612);
nand U6350 (N_6350,In_1575,In_2599);
nand U6351 (N_6351,In_57,In_1409);
xor U6352 (N_6352,In_109,In_98);
and U6353 (N_6353,In_4620,In_3348);
nor U6354 (N_6354,In_3105,In_4705);
nand U6355 (N_6355,In_4530,In_3420);
or U6356 (N_6356,In_2625,In_4956);
and U6357 (N_6357,In_3499,In_809);
and U6358 (N_6358,In_1268,In_3496);
xor U6359 (N_6359,In_2179,In_3341);
or U6360 (N_6360,In_2752,In_4000);
nor U6361 (N_6361,In_2708,In_1283);
nand U6362 (N_6362,In_4005,In_1506);
nand U6363 (N_6363,In_3519,In_3043);
or U6364 (N_6364,In_4215,In_4109);
or U6365 (N_6365,In_2692,In_3085);
nand U6366 (N_6366,In_1848,In_2435);
nand U6367 (N_6367,In_4865,In_884);
and U6368 (N_6368,In_4255,In_855);
nand U6369 (N_6369,In_2444,In_1772);
nor U6370 (N_6370,In_4809,In_2637);
nor U6371 (N_6371,In_4373,In_3626);
or U6372 (N_6372,In_2683,In_909);
and U6373 (N_6373,In_3557,In_1891);
or U6374 (N_6374,In_1671,In_4229);
xor U6375 (N_6375,In_2505,In_3692);
xnor U6376 (N_6376,In_684,In_2985);
xnor U6377 (N_6377,In_899,In_4202);
xnor U6378 (N_6378,In_180,In_453);
or U6379 (N_6379,In_3785,In_4879);
nand U6380 (N_6380,In_4465,In_2000);
nand U6381 (N_6381,In_1770,In_2240);
nor U6382 (N_6382,In_1464,In_1591);
nor U6383 (N_6383,In_2237,In_3115);
nor U6384 (N_6384,In_2119,In_1879);
or U6385 (N_6385,In_1793,In_3437);
xnor U6386 (N_6386,In_4526,In_2956);
or U6387 (N_6387,In_2327,In_1333);
nand U6388 (N_6388,In_1434,In_4627);
nor U6389 (N_6389,In_3611,In_3254);
nor U6390 (N_6390,In_4335,In_1411);
nand U6391 (N_6391,In_2819,In_3393);
and U6392 (N_6392,In_699,In_4134);
and U6393 (N_6393,In_2206,In_3589);
xor U6394 (N_6394,In_3403,In_1150);
xnor U6395 (N_6395,In_4558,In_947);
nand U6396 (N_6396,In_1501,In_3001);
or U6397 (N_6397,In_3336,In_4764);
and U6398 (N_6398,In_4129,In_1026);
xor U6399 (N_6399,In_133,In_2891);
or U6400 (N_6400,In_37,In_3651);
xor U6401 (N_6401,In_3459,In_858);
nor U6402 (N_6402,In_4010,In_1779);
or U6403 (N_6403,In_3920,In_1781);
nand U6404 (N_6404,In_73,In_2969);
or U6405 (N_6405,In_1801,In_2054);
nand U6406 (N_6406,In_2229,In_431);
or U6407 (N_6407,In_2022,In_1936);
or U6408 (N_6408,In_946,In_656);
nor U6409 (N_6409,In_3861,In_2171);
nand U6410 (N_6410,In_3038,In_3297);
nor U6411 (N_6411,In_3403,In_2957);
or U6412 (N_6412,In_2521,In_4739);
nand U6413 (N_6413,In_3045,In_2461);
and U6414 (N_6414,In_1133,In_129);
nand U6415 (N_6415,In_2298,In_1516);
or U6416 (N_6416,In_3526,In_1302);
xnor U6417 (N_6417,In_2459,In_2099);
xnor U6418 (N_6418,In_4230,In_1015);
and U6419 (N_6419,In_417,In_11);
and U6420 (N_6420,In_486,In_1814);
and U6421 (N_6421,In_3113,In_4180);
xor U6422 (N_6422,In_436,In_1936);
nor U6423 (N_6423,In_504,In_3261);
nor U6424 (N_6424,In_300,In_911);
xor U6425 (N_6425,In_3452,In_814);
nor U6426 (N_6426,In_1220,In_1080);
and U6427 (N_6427,In_4288,In_1527);
xnor U6428 (N_6428,In_407,In_81);
nand U6429 (N_6429,In_4857,In_385);
or U6430 (N_6430,In_1719,In_702);
or U6431 (N_6431,In_4137,In_2948);
or U6432 (N_6432,In_4094,In_2058);
nand U6433 (N_6433,In_2051,In_4733);
or U6434 (N_6434,In_4529,In_3974);
and U6435 (N_6435,In_685,In_3359);
nand U6436 (N_6436,In_4466,In_933);
nand U6437 (N_6437,In_3440,In_4967);
xor U6438 (N_6438,In_1209,In_1415);
and U6439 (N_6439,In_3059,In_292);
nand U6440 (N_6440,In_3298,In_108);
nand U6441 (N_6441,In_1836,In_4430);
nand U6442 (N_6442,In_3300,In_1141);
xor U6443 (N_6443,In_3076,In_4054);
and U6444 (N_6444,In_4167,In_2556);
xnor U6445 (N_6445,In_3901,In_3962);
xnor U6446 (N_6446,In_4229,In_77);
and U6447 (N_6447,In_333,In_2080);
nand U6448 (N_6448,In_2871,In_2661);
or U6449 (N_6449,In_4829,In_782);
nand U6450 (N_6450,In_2615,In_2512);
nand U6451 (N_6451,In_2814,In_3129);
nand U6452 (N_6452,In_2314,In_3718);
nand U6453 (N_6453,In_4421,In_540);
nor U6454 (N_6454,In_1895,In_984);
and U6455 (N_6455,In_2385,In_3102);
or U6456 (N_6456,In_1209,In_3597);
nor U6457 (N_6457,In_3845,In_62);
nand U6458 (N_6458,In_1588,In_4360);
xnor U6459 (N_6459,In_2316,In_3834);
or U6460 (N_6460,In_3507,In_3978);
and U6461 (N_6461,In_2888,In_1684);
xnor U6462 (N_6462,In_1048,In_111);
nand U6463 (N_6463,In_3666,In_2600);
nand U6464 (N_6464,In_750,In_1501);
or U6465 (N_6465,In_1299,In_793);
or U6466 (N_6466,In_3608,In_2194);
nand U6467 (N_6467,In_4847,In_2761);
and U6468 (N_6468,In_3240,In_4678);
xnor U6469 (N_6469,In_3540,In_1402);
or U6470 (N_6470,In_514,In_1182);
nor U6471 (N_6471,In_1568,In_2288);
nand U6472 (N_6472,In_2992,In_635);
xor U6473 (N_6473,In_765,In_4045);
nor U6474 (N_6474,In_2196,In_388);
nor U6475 (N_6475,In_440,In_2420);
xor U6476 (N_6476,In_3771,In_1006);
or U6477 (N_6477,In_1365,In_1245);
nand U6478 (N_6478,In_2919,In_111);
and U6479 (N_6479,In_4107,In_1033);
xnor U6480 (N_6480,In_3253,In_1568);
and U6481 (N_6481,In_4503,In_2852);
nor U6482 (N_6482,In_931,In_4788);
xor U6483 (N_6483,In_4444,In_3876);
and U6484 (N_6484,In_3731,In_2594);
and U6485 (N_6485,In_3013,In_4008);
nand U6486 (N_6486,In_914,In_4038);
xnor U6487 (N_6487,In_4082,In_1419);
or U6488 (N_6488,In_563,In_3531);
nor U6489 (N_6489,In_2945,In_1576);
nand U6490 (N_6490,In_201,In_4944);
nor U6491 (N_6491,In_3030,In_137);
and U6492 (N_6492,In_1437,In_3424);
nor U6493 (N_6493,In_315,In_1866);
nor U6494 (N_6494,In_941,In_75);
and U6495 (N_6495,In_1953,In_4313);
nor U6496 (N_6496,In_4332,In_315);
and U6497 (N_6497,In_3170,In_41);
and U6498 (N_6498,In_4621,In_1826);
nand U6499 (N_6499,In_2633,In_4417);
xnor U6500 (N_6500,In_4049,In_1540);
nor U6501 (N_6501,In_1215,In_1724);
xnor U6502 (N_6502,In_2163,In_2771);
and U6503 (N_6503,In_2652,In_3388);
or U6504 (N_6504,In_251,In_3339);
or U6505 (N_6505,In_3710,In_277);
nor U6506 (N_6506,In_1411,In_960);
and U6507 (N_6507,In_3853,In_4151);
xnor U6508 (N_6508,In_2736,In_84);
and U6509 (N_6509,In_3860,In_2461);
xor U6510 (N_6510,In_3147,In_109);
and U6511 (N_6511,In_2704,In_2266);
nor U6512 (N_6512,In_738,In_139);
xor U6513 (N_6513,In_3289,In_729);
xnor U6514 (N_6514,In_3935,In_4996);
or U6515 (N_6515,In_1096,In_2402);
xnor U6516 (N_6516,In_2641,In_1212);
and U6517 (N_6517,In_4603,In_4267);
nand U6518 (N_6518,In_998,In_3796);
and U6519 (N_6519,In_3549,In_598);
nand U6520 (N_6520,In_986,In_4544);
nor U6521 (N_6521,In_4831,In_3846);
xor U6522 (N_6522,In_2948,In_1665);
or U6523 (N_6523,In_1319,In_4106);
or U6524 (N_6524,In_742,In_3322);
or U6525 (N_6525,In_2748,In_2702);
nand U6526 (N_6526,In_1711,In_2227);
and U6527 (N_6527,In_300,In_4291);
nor U6528 (N_6528,In_3363,In_325);
xor U6529 (N_6529,In_2079,In_3830);
nor U6530 (N_6530,In_1014,In_1741);
nor U6531 (N_6531,In_4560,In_1628);
nor U6532 (N_6532,In_1180,In_899);
xor U6533 (N_6533,In_4064,In_4518);
nor U6534 (N_6534,In_1591,In_1165);
nand U6535 (N_6535,In_52,In_2654);
or U6536 (N_6536,In_4559,In_1431);
xnor U6537 (N_6537,In_2212,In_4948);
nor U6538 (N_6538,In_824,In_1088);
nor U6539 (N_6539,In_3768,In_4130);
and U6540 (N_6540,In_3699,In_3538);
and U6541 (N_6541,In_4879,In_4476);
xnor U6542 (N_6542,In_4028,In_299);
nand U6543 (N_6543,In_1518,In_1472);
nor U6544 (N_6544,In_4654,In_583);
or U6545 (N_6545,In_2825,In_4712);
and U6546 (N_6546,In_3131,In_2050);
xnor U6547 (N_6547,In_1610,In_3425);
or U6548 (N_6548,In_4823,In_2612);
xnor U6549 (N_6549,In_37,In_4495);
nand U6550 (N_6550,In_228,In_4507);
nor U6551 (N_6551,In_4597,In_1251);
and U6552 (N_6552,In_4377,In_1219);
nand U6553 (N_6553,In_4706,In_3939);
and U6554 (N_6554,In_2343,In_1430);
or U6555 (N_6555,In_2553,In_1987);
and U6556 (N_6556,In_4557,In_3751);
and U6557 (N_6557,In_1367,In_1423);
xor U6558 (N_6558,In_2710,In_3645);
nand U6559 (N_6559,In_1559,In_789);
nor U6560 (N_6560,In_1701,In_4893);
nand U6561 (N_6561,In_3225,In_1571);
or U6562 (N_6562,In_1431,In_4192);
xor U6563 (N_6563,In_4031,In_3897);
or U6564 (N_6564,In_3314,In_3563);
and U6565 (N_6565,In_776,In_1574);
nor U6566 (N_6566,In_4346,In_1781);
or U6567 (N_6567,In_2742,In_2309);
nor U6568 (N_6568,In_1061,In_3764);
and U6569 (N_6569,In_1438,In_4306);
or U6570 (N_6570,In_1486,In_2646);
or U6571 (N_6571,In_2079,In_196);
or U6572 (N_6572,In_4570,In_4580);
xnor U6573 (N_6573,In_4244,In_864);
nor U6574 (N_6574,In_2562,In_458);
nand U6575 (N_6575,In_1294,In_870);
or U6576 (N_6576,In_2999,In_2998);
nand U6577 (N_6577,In_4692,In_3991);
nand U6578 (N_6578,In_3164,In_1702);
or U6579 (N_6579,In_3619,In_1948);
xor U6580 (N_6580,In_1443,In_2753);
or U6581 (N_6581,In_2110,In_2489);
xor U6582 (N_6582,In_1692,In_1044);
xor U6583 (N_6583,In_2956,In_3040);
xnor U6584 (N_6584,In_2494,In_3570);
nand U6585 (N_6585,In_223,In_3040);
or U6586 (N_6586,In_1029,In_2218);
nor U6587 (N_6587,In_688,In_4753);
xnor U6588 (N_6588,In_1493,In_3897);
and U6589 (N_6589,In_895,In_3509);
nor U6590 (N_6590,In_1881,In_4571);
nor U6591 (N_6591,In_2626,In_2658);
or U6592 (N_6592,In_4529,In_2760);
nor U6593 (N_6593,In_236,In_782);
and U6594 (N_6594,In_4348,In_2681);
and U6595 (N_6595,In_624,In_3875);
and U6596 (N_6596,In_3679,In_1830);
nor U6597 (N_6597,In_382,In_3173);
or U6598 (N_6598,In_882,In_4906);
nand U6599 (N_6599,In_321,In_57);
nor U6600 (N_6600,In_2854,In_1019);
and U6601 (N_6601,In_683,In_2058);
nand U6602 (N_6602,In_1711,In_2548);
xor U6603 (N_6603,In_3417,In_2356);
xnor U6604 (N_6604,In_3232,In_2826);
nand U6605 (N_6605,In_3533,In_3027);
nor U6606 (N_6606,In_247,In_2200);
and U6607 (N_6607,In_4922,In_1162);
xor U6608 (N_6608,In_3003,In_2859);
or U6609 (N_6609,In_3868,In_269);
nor U6610 (N_6610,In_753,In_800);
nand U6611 (N_6611,In_2265,In_10);
xor U6612 (N_6612,In_4357,In_444);
nand U6613 (N_6613,In_2979,In_3824);
nand U6614 (N_6614,In_89,In_2665);
nand U6615 (N_6615,In_2915,In_3156);
nand U6616 (N_6616,In_4180,In_500);
xnor U6617 (N_6617,In_1965,In_3788);
nor U6618 (N_6618,In_3643,In_2272);
nor U6619 (N_6619,In_2369,In_829);
nor U6620 (N_6620,In_4194,In_4700);
xor U6621 (N_6621,In_4571,In_3005);
and U6622 (N_6622,In_387,In_3661);
and U6623 (N_6623,In_41,In_2396);
nand U6624 (N_6624,In_3939,In_4670);
and U6625 (N_6625,In_2166,In_711);
nor U6626 (N_6626,In_1360,In_2877);
or U6627 (N_6627,In_614,In_1358);
nor U6628 (N_6628,In_1359,In_1419);
xnor U6629 (N_6629,In_2668,In_357);
nor U6630 (N_6630,In_4059,In_4117);
and U6631 (N_6631,In_2935,In_761);
nor U6632 (N_6632,In_1833,In_4265);
and U6633 (N_6633,In_4929,In_633);
or U6634 (N_6634,In_4882,In_4914);
nand U6635 (N_6635,In_3134,In_3023);
and U6636 (N_6636,In_1169,In_3423);
xor U6637 (N_6637,In_4911,In_3205);
or U6638 (N_6638,In_3888,In_653);
or U6639 (N_6639,In_659,In_1469);
xor U6640 (N_6640,In_4993,In_515);
and U6641 (N_6641,In_1499,In_3095);
xnor U6642 (N_6642,In_287,In_11);
and U6643 (N_6643,In_1317,In_2666);
xor U6644 (N_6644,In_4753,In_1843);
or U6645 (N_6645,In_1182,In_1691);
nor U6646 (N_6646,In_664,In_3935);
or U6647 (N_6647,In_935,In_2250);
and U6648 (N_6648,In_3482,In_1002);
xor U6649 (N_6649,In_2770,In_4703);
nor U6650 (N_6650,In_4543,In_3718);
or U6651 (N_6651,In_3541,In_3408);
nor U6652 (N_6652,In_388,In_4926);
nor U6653 (N_6653,In_1993,In_3551);
nand U6654 (N_6654,In_3567,In_4009);
and U6655 (N_6655,In_151,In_3002);
nor U6656 (N_6656,In_515,In_2927);
or U6657 (N_6657,In_1564,In_4128);
nand U6658 (N_6658,In_119,In_1646);
nor U6659 (N_6659,In_2625,In_4274);
xor U6660 (N_6660,In_1108,In_3960);
or U6661 (N_6661,In_4792,In_2906);
nor U6662 (N_6662,In_965,In_4837);
and U6663 (N_6663,In_3387,In_1171);
nor U6664 (N_6664,In_88,In_514);
nand U6665 (N_6665,In_819,In_1434);
xor U6666 (N_6666,In_1632,In_4187);
nand U6667 (N_6667,In_3818,In_1063);
or U6668 (N_6668,In_507,In_3124);
or U6669 (N_6669,In_4161,In_2363);
xor U6670 (N_6670,In_4416,In_2185);
or U6671 (N_6671,In_4683,In_4415);
or U6672 (N_6672,In_3354,In_255);
nor U6673 (N_6673,In_123,In_909);
nor U6674 (N_6674,In_3917,In_1882);
nor U6675 (N_6675,In_2373,In_3035);
xnor U6676 (N_6676,In_4488,In_2708);
nor U6677 (N_6677,In_4325,In_1926);
and U6678 (N_6678,In_2021,In_4598);
xnor U6679 (N_6679,In_34,In_615);
nand U6680 (N_6680,In_2282,In_4072);
xnor U6681 (N_6681,In_2346,In_2813);
nand U6682 (N_6682,In_4900,In_1153);
nand U6683 (N_6683,In_2789,In_34);
and U6684 (N_6684,In_2531,In_3990);
and U6685 (N_6685,In_4380,In_2317);
xnor U6686 (N_6686,In_1841,In_537);
nor U6687 (N_6687,In_3732,In_1322);
or U6688 (N_6688,In_3790,In_3232);
nor U6689 (N_6689,In_1331,In_2238);
and U6690 (N_6690,In_4745,In_4706);
or U6691 (N_6691,In_1181,In_1402);
xnor U6692 (N_6692,In_651,In_4781);
xnor U6693 (N_6693,In_1037,In_973);
and U6694 (N_6694,In_1665,In_3449);
nor U6695 (N_6695,In_1712,In_3461);
and U6696 (N_6696,In_2910,In_2178);
and U6697 (N_6697,In_4999,In_3184);
and U6698 (N_6698,In_4301,In_3862);
xor U6699 (N_6699,In_705,In_896);
nand U6700 (N_6700,In_1673,In_3610);
xor U6701 (N_6701,In_657,In_1001);
or U6702 (N_6702,In_398,In_882);
xor U6703 (N_6703,In_2913,In_635);
and U6704 (N_6704,In_584,In_1587);
nand U6705 (N_6705,In_569,In_798);
xnor U6706 (N_6706,In_65,In_2076);
and U6707 (N_6707,In_1877,In_4709);
or U6708 (N_6708,In_4426,In_4028);
or U6709 (N_6709,In_3736,In_161);
nor U6710 (N_6710,In_1017,In_4853);
and U6711 (N_6711,In_2529,In_2393);
nand U6712 (N_6712,In_4159,In_3508);
and U6713 (N_6713,In_4918,In_1682);
or U6714 (N_6714,In_372,In_3975);
xnor U6715 (N_6715,In_3985,In_3092);
or U6716 (N_6716,In_3846,In_2482);
nor U6717 (N_6717,In_1697,In_2528);
nand U6718 (N_6718,In_409,In_3452);
nor U6719 (N_6719,In_1030,In_2225);
xnor U6720 (N_6720,In_3926,In_2413);
nand U6721 (N_6721,In_3416,In_2095);
nand U6722 (N_6722,In_1430,In_3806);
or U6723 (N_6723,In_1628,In_3289);
and U6724 (N_6724,In_1863,In_1580);
xor U6725 (N_6725,In_114,In_3449);
or U6726 (N_6726,In_2431,In_1728);
nand U6727 (N_6727,In_1016,In_1468);
or U6728 (N_6728,In_4027,In_4526);
nor U6729 (N_6729,In_4534,In_2011);
or U6730 (N_6730,In_1718,In_932);
nand U6731 (N_6731,In_114,In_1480);
nor U6732 (N_6732,In_3650,In_718);
xnor U6733 (N_6733,In_152,In_2177);
or U6734 (N_6734,In_1237,In_1325);
xor U6735 (N_6735,In_2394,In_4959);
and U6736 (N_6736,In_2635,In_4107);
nand U6737 (N_6737,In_275,In_3055);
nor U6738 (N_6738,In_1552,In_3500);
or U6739 (N_6739,In_903,In_1171);
nor U6740 (N_6740,In_2656,In_4323);
nor U6741 (N_6741,In_2682,In_478);
and U6742 (N_6742,In_2425,In_2337);
or U6743 (N_6743,In_2193,In_2460);
nor U6744 (N_6744,In_808,In_1388);
nand U6745 (N_6745,In_1992,In_153);
or U6746 (N_6746,In_3911,In_3723);
and U6747 (N_6747,In_3277,In_1680);
and U6748 (N_6748,In_161,In_117);
nor U6749 (N_6749,In_2463,In_1203);
xor U6750 (N_6750,In_615,In_2697);
nor U6751 (N_6751,In_1570,In_144);
and U6752 (N_6752,In_4951,In_545);
nand U6753 (N_6753,In_4077,In_2017);
xor U6754 (N_6754,In_4187,In_2513);
nor U6755 (N_6755,In_992,In_4106);
and U6756 (N_6756,In_1684,In_178);
or U6757 (N_6757,In_3655,In_4971);
nand U6758 (N_6758,In_228,In_358);
and U6759 (N_6759,In_1067,In_4139);
and U6760 (N_6760,In_491,In_4953);
or U6761 (N_6761,In_1323,In_1950);
or U6762 (N_6762,In_1819,In_4049);
nor U6763 (N_6763,In_248,In_2489);
xor U6764 (N_6764,In_3194,In_839);
xor U6765 (N_6765,In_145,In_2872);
xor U6766 (N_6766,In_1762,In_4462);
and U6767 (N_6767,In_328,In_3384);
or U6768 (N_6768,In_1607,In_1891);
or U6769 (N_6769,In_223,In_3284);
nor U6770 (N_6770,In_2835,In_2571);
and U6771 (N_6771,In_2325,In_1226);
and U6772 (N_6772,In_2684,In_1224);
or U6773 (N_6773,In_3978,In_4611);
and U6774 (N_6774,In_1923,In_3765);
nor U6775 (N_6775,In_711,In_1803);
xnor U6776 (N_6776,In_607,In_884);
nor U6777 (N_6777,In_2247,In_313);
or U6778 (N_6778,In_210,In_534);
xor U6779 (N_6779,In_911,In_846);
nor U6780 (N_6780,In_897,In_3019);
xor U6781 (N_6781,In_995,In_1422);
and U6782 (N_6782,In_3854,In_2101);
or U6783 (N_6783,In_3635,In_3552);
and U6784 (N_6784,In_1631,In_532);
and U6785 (N_6785,In_4297,In_4776);
xor U6786 (N_6786,In_3143,In_680);
and U6787 (N_6787,In_703,In_343);
and U6788 (N_6788,In_575,In_562);
xnor U6789 (N_6789,In_4872,In_420);
nand U6790 (N_6790,In_2286,In_2472);
xor U6791 (N_6791,In_2353,In_989);
xor U6792 (N_6792,In_1304,In_2855);
nand U6793 (N_6793,In_4797,In_3664);
nor U6794 (N_6794,In_1718,In_1527);
nor U6795 (N_6795,In_3511,In_4942);
xnor U6796 (N_6796,In_2884,In_4042);
nor U6797 (N_6797,In_4468,In_1301);
or U6798 (N_6798,In_3931,In_1304);
or U6799 (N_6799,In_1524,In_781);
or U6800 (N_6800,In_2435,In_3049);
xor U6801 (N_6801,In_801,In_950);
or U6802 (N_6802,In_639,In_2394);
or U6803 (N_6803,In_436,In_1790);
nand U6804 (N_6804,In_477,In_4490);
xor U6805 (N_6805,In_2420,In_2637);
nor U6806 (N_6806,In_723,In_1609);
and U6807 (N_6807,In_155,In_3752);
xor U6808 (N_6808,In_3734,In_4522);
nand U6809 (N_6809,In_2398,In_4888);
nor U6810 (N_6810,In_4038,In_839);
or U6811 (N_6811,In_1434,In_2710);
xor U6812 (N_6812,In_2953,In_4692);
xor U6813 (N_6813,In_4718,In_1279);
xnor U6814 (N_6814,In_597,In_892);
nand U6815 (N_6815,In_1602,In_4366);
and U6816 (N_6816,In_1942,In_987);
xnor U6817 (N_6817,In_299,In_4093);
nand U6818 (N_6818,In_2715,In_2183);
or U6819 (N_6819,In_761,In_3517);
nor U6820 (N_6820,In_627,In_4529);
xor U6821 (N_6821,In_921,In_4183);
nor U6822 (N_6822,In_4637,In_2749);
nor U6823 (N_6823,In_3191,In_937);
nor U6824 (N_6824,In_1345,In_1674);
nand U6825 (N_6825,In_2959,In_3677);
nor U6826 (N_6826,In_3345,In_45);
xnor U6827 (N_6827,In_2142,In_3776);
nand U6828 (N_6828,In_2371,In_4814);
and U6829 (N_6829,In_3404,In_4882);
nor U6830 (N_6830,In_4875,In_3013);
and U6831 (N_6831,In_2650,In_3058);
nand U6832 (N_6832,In_507,In_1764);
nor U6833 (N_6833,In_1051,In_135);
nand U6834 (N_6834,In_2616,In_4812);
or U6835 (N_6835,In_968,In_1154);
nor U6836 (N_6836,In_1344,In_2320);
xnor U6837 (N_6837,In_3547,In_1046);
and U6838 (N_6838,In_1660,In_3282);
or U6839 (N_6839,In_1578,In_1802);
nand U6840 (N_6840,In_4061,In_4817);
xnor U6841 (N_6841,In_354,In_1577);
and U6842 (N_6842,In_103,In_1126);
nor U6843 (N_6843,In_3944,In_2591);
or U6844 (N_6844,In_3653,In_120);
or U6845 (N_6845,In_4323,In_2856);
and U6846 (N_6846,In_3447,In_2050);
and U6847 (N_6847,In_3507,In_3231);
and U6848 (N_6848,In_3369,In_4263);
xnor U6849 (N_6849,In_1198,In_4935);
or U6850 (N_6850,In_4517,In_4421);
or U6851 (N_6851,In_811,In_3146);
nand U6852 (N_6852,In_1173,In_403);
nor U6853 (N_6853,In_419,In_4544);
nand U6854 (N_6854,In_2763,In_4326);
nor U6855 (N_6855,In_3113,In_263);
or U6856 (N_6856,In_164,In_3654);
nand U6857 (N_6857,In_2766,In_2609);
and U6858 (N_6858,In_3164,In_3750);
and U6859 (N_6859,In_4751,In_44);
and U6860 (N_6860,In_1461,In_4065);
or U6861 (N_6861,In_1332,In_3151);
xnor U6862 (N_6862,In_1017,In_3744);
nand U6863 (N_6863,In_2755,In_4786);
and U6864 (N_6864,In_1406,In_1903);
or U6865 (N_6865,In_3373,In_2697);
nor U6866 (N_6866,In_3842,In_3726);
xnor U6867 (N_6867,In_4430,In_4799);
nand U6868 (N_6868,In_1753,In_862);
xnor U6869 (N_6869,In_2593,In_300);
nor U6870 (N_6870,In_1534,In_1195);
xor U6871 (N_6871,In_3336,In_3669);
and U6872 (N_6872,In_132,In_4946);
xor U6873 (N_6873,In_3689,In_1201);
or U6874 (N_6874,In_767,In_258);
and U6875 (N_6875,In_4842,In_4819);
xor U6876 (N_6876,In_126,In_840);
xnor U6877 (N_6877,In_2386,In_1852);
or U6878 (N_6878,In_2668,In_1763);
nor U6879 (N_6879,In_1587,In_593);
and U6880 (N_6880,In_3480,In_3512);
nand U6881 (N_6881,In_2262,In_4332);
xor U6882 (N_6882,In_4115,In_3355);
or U6883 (N_6883,In_877,In_3658);
nand U6884 (N_6884,In_866,In_3573);
or U6885 (N_6885,In_3487,In_510);
nor U6886 (N_6886,In_4645,In_4649);
nor U6887 (N_6887,In_4144,In_4450);
nand U6888 (N_6888,In_1016,In_4029);
nand U6889 (N_6889,In_3137,In_2437);
nor U6890 (N_6890,In_3955,In_1653);
nor U6891 (N_6891,In_3038,In_3527);
and U6892 (N_6892,In_3827,In_2048);
or U6893 (N_6893,In_4595,In_828);
and U6894 (N_6894,In_3313,In_4292);
xnor U6895 (N_6895,In_3752,In_4012);
nand U6896 (N_6896,In_3310,In_1947);
nor U6897 (N_6897,In_4707,In_4553);
xor U6898 (N_6898,In_3646,In_1262);
nor U6899 (N_6899,In_4307,In_1306);
nor U6900 (N_6900,In_4546,In_4712);
xor U6901 (N_6901,In_1134,In_402);
xor U6902 (N_6902,In_1396,In_2539);
or U6903 (N_6903,In_2838,In_2957);
nand U6904 (N_6904,In_1107,In_431);
xor U6905 (N_6905,In_1181,In_4562);
nand U6906 (N_6906,In_4728,In_2623);
and U6907 (N_6907,In_4797,In_3502);
nand U6908 (N_6908,In_2714,In_3063);
nor U6909 (N_6909,In_2292,In_52);
nand U6910 (N_6910,In_3975,In_4385);
and U6911 (N_6911,In_2479,In_1606);
xor U6912 (N_6912,In_2579,In_2338);
xnor U6913 (N_6913,In_3707,In_4248);
nor U6914 (N_6914,In_3071,In_1069);
nand U6915 (N_6915,In_919,In_1662);
xor U6916 (N_6916,In_698,In_2527);
and U6917 (N_6917,In_2513,In_2271);
xor U6918 (N_6918,In_2442,In_3612);
and U6919 (N_6919,In_1271,In_167);
nand U6920 (N_6920,In_3358,In_2015);
xnor U6921 (N_6921,In_2635,In_2994);
and U6922 (N_6922,In_2913,In_999);
nand U6923 (N_6923,In_2511,In_3192);
and U6924 (N_6924,In_1826,In_4385);
and U6925 (N_6925,In_3263,In_2589);
xor U6926 (N_6926,In_1830,In_1705);
nand U6927 (N_6927,In_2227,In_1250);
xnor U6928 (N_6928,In_1594,In_2170);
xnor U6929 (N_6929,In_1152,In_4046);
nor U6930 (N_6930,In_602,In_2189);
xnor U6931 (N_6931,In_3095,In_133);
nand U6932 (N_6932,In_984,In_3156);
xor U6933 (N_6933,In_3316,In_2234);
nand U6934 (N_6934,In_2485,In_4340);
xor U6935 (N_6935,In_1232,In_3158);
xor U6936 (N_6936,In_4928,In_3088);
nor U6937 (N_6937,In_4733,In_2004);
and U6938 (N_6938,In_4829,In_3763);
nor U6939 (N_6939,In_2869,In_2946);
xnor U6940 (N_6940,In_2073,In_2177);
and U6941 (N_6941,In_746,In_2047);
nand U6942 (N_6942,In_425,In_399);
nand U6943 (N_6943,In_2833,In_1052);
or U6944 (N_6944,In_3161,In_3442);
nor U6945 (N_6945,In_3982,In_4248);
and U6946 (N_6946,In_419,In_529);
nand U6947 (N_6947,In_3062,In_4497);
xnor U6948 (N_6948,In_722,In_1699);
or U6949 (N_6949,In_796,In_973);
nand U6950 (N_6950,In_4284,In_3014);
nor U6951 (N_6951,In_4976,In_3659);
nor U6952 (N_6952,In_118,In_4142);
nor U6953 (N_6953,In_4205,In_1004);
nor U6954 (N_6954,In_3272,In_4877);
or U6955 (N_6955,In_4651,In_1751);
nor U6956 (N_6956,In_2824,In_1639);
nor U6957 (N_6957,In_3243,In_3367);
and U6958 (N_6958,In_1446,In_264);
or U6959 (N_6959,In_325,In_4046);
and U6960 (N_6960,In_4394,In_3710);
or U6961 (N_6961,In_477,In_3200);
nor U6962 (N_6962,In_1151,In_2199);
or U6963 (N_6963,In_2148,In_3718);
xor U6964 (N_6964,In_1719,In_4854);
nand U6965 (N_6965,In_268,In_3812);
xnor U6966 (N_6966,In_127,In_1882);
nor U6967 (N_6967,In_3957,In_4807);
or U6968 (N_6968,In_3353,In_3303);
nor U6969 (N_6969,In_1352,In_2032);
xor U6970 (N_6970,In_1788,In_2259);
and U6971 (N_6971,In_2169,In_1657);
nand U6972 (N_6972,In_895,In_566);
nand U6973 (N_6973,In_3636,In_1400);
nand U6974 (N_6974,In_3761,In_1552);
and U6975 (N_6975,In_2527,In_3871);
nand U6976 (N_6976,In_3683,In_985);
and U6977 (N_6977,In_4800,In_3047);
nand U6978 (N_6978,In_3435,In_705);
nand U6979 (N_6979,In_4926,In_3304);
nand U6980 (N_6980,In_963,In_3621);
or U6981 (N_6981,In_1624,In_1452);
xor U6982 (N_6982,In_976,In_13);
xnor U6983 (N_6983,In_500,In_1474);
nor U6984 (N_6984,In_2331,In_3043);
and U6985 (N_6985,In_1375,In_203);
xnor U6986 (N_6986,In_1840,In_4763);
nand U6987 (N_6987,In_1809,In_4958);
or U6988 (N_6988,In_2857,In_2421);
nor U6989 (N_6989,In_3498,In_3427);
nand U6990 (N_6990,In_499,In_2835);
or U6991 (N_6991,In_4812,In_3507);
xor U6992 (N_6992,In_3836,In_3779);
nand U6993 (N_6993,In_2189,In_3441);
xnor U6994 (N_6994,In_2647,In_2191);
nor U6995 (N_6995,In_597,In_2415);
xor U6996 (N_6996,In_3800,In_1466);
or U6997 (N_6997,In_1481,In_3961);
xor U6998 (N_6998,In_4452,In_3304);
xnor U6999 (N_6999,In_1082,In_3674);
xor U7000 (N_7000,In_4432,In_2120);
xnor U7001 (N_7001,In_922,In_2306);
and U7002 (N_7002,In_3875,In_3463);
xnor U7003 (N_7003,In_4474,In_4000);
or U7004 (N_7004,In_1538,In_2542);
nor U7005 (N_7005,In_3995,In_2749);
and U7006 (N_7006,In_3811,In_321);
or U7007 (N_7007,In_2760,In_1017);
or U7008 (N_7008,In_4357,In_3143);
nand U7009 (N_7009,In_1116,In_2952);
or U7010 (N_7010,In_1729,In_1947);
xor U7011 (N_7011,In_3814,In_4174);
nand U7012 (N_7012,In_370,In_3715);
xnor U7013 (N_7013,In_4753,In_4011);
nand U7014 (N_7014,In_3699,In_2652);
and U7015 (N_7015,In_2205,In_1215);
xnor U7016 (N_7016,In_459,In_2209);
xor U7017 (N_7017,In_4689,In_3231);
xnor U7018 (N_7018,In_1781,In_1549);
and U7019 (N_7019,In_1618,In_2957);
nand U7020 (N_7020,In_433,In_643);
and U7021 (N_7021,In_1362,In_4273);
nor U7022 (N_7022,In_1654,In_978);
xor U7023 (N_7023,In_535,In_1669);
nor U7024 (N_7024,In_2824,In_4373);
and U7025 (N_7025,In_631,In_2262);
or U7026 (N_7026,In_4644,In_516);
and U7027 (N_7027,In_135,In_47);
or U7028 (N_7028,In_2626,In_3182);
nand U7029 (N_7029,In_156,In_4688);
and U7030 (N_7030,In_4452,In_1377);
and U7031 (N_7031,In_3076,In_4074);
or U7032 (N_7032,In_633,In_1897);
nor U7033 (N_7033,In_1031,In_4278);
or U7034 (N_7034,In_3271,In_4279);
and U7035 (N_7035,In_1832,In_1510);
nand U7036 (N_7036,In_3496,In_698);
xor U7037 (N_7037,In_3332,In_4831);
or U7038 (N_7038,In_2103,In_4681);
nand U7039 (N_7039,In_1228,In_4267);
nand U7040 (N_7040,In_4473,In_4283);
or U7041 (N_7041,In_237,In_1522);
or U7042 (N_7042,In_431,In_154);
xor U7043 (N_7043,In_4862,In_2579);
nand U7044 (N_7044,In_3324,In_3302);
xor U7045 (N_7045,In_3351,In_1921);
nand U7046 (N_7046,In_1011,In_1010);
or U7047 (N_7047,In_1164,In_80);
and U7048 (N_7048,In_2600,In_1862);
xor U7049 (N_7049,In_3029,In_1914);
or U7050 (N_7050,In_3533,In_19);
xnor U7051 (N_7051,In_1042,In_4200);
or U7052 (N_7052,In_4039,In_3003);
and U7053 (N_7053,In_827,In_4945);
and U7054 (N_7054,In_2812,In_2779);
nor U7055 (N_7055,In_3993,In_958);
nand U7056 (N_7056,In_2815,In_3477);
nand U7057 (N_7057,In_2190,In_4897);
nor U7058 (N_7058,In_2125,In_3552);
nor U7059 (N_7059,In_3074,In_321);
nor U7060 (N_7060,In_4786,In_2462);
xor U7061 (N_7061,In_4097,In_91);
xnor U7062 (N_7062,In_2481,In_2051);
and U7063 (N_7063,In_2609,In_1460);
xor U7064 (N_7064,In_3160,In_3037);
xor U7065 (N_7065,In_1089,In_1209);
xnor U7066 (N_7066,In_4496,In_3818);
nand U7067 (N_7067,In_521,In_107);
or U7068 (N_7068,In_4318,In_3051);
or U7069 (N_7069,In_1019,In_4391);
xnor U7070 (N_7070,In_2356,In_1916);
and U7071 (N_7071,In_3310,In_4711);
or U7072 (N_7072,In_1314,In_1343);
nor U7073 (N_7073,In_939,In_2247);
and U7074 (N_7074,In_4655,In_3123);
nand U7075 (N_7075,In_4061,In_4675);
or U7076 (N_7076,In_1488,In_4294);
nor U7077 (N_7077,In_3430,In_4961);
or U7078 (N_7078,In_2444,In_3102);
or U7079 (N_7079,In_871,In_2775);
nor U7080 (N_7080,In_179,In_2759);
and U7081 (N_7081,In_3999,In_1234);
nand U7082 (N_7082,In_3316,In_1427);
nor U7083 (N_7083,In_4842,In_3186);
or U7084 (N_7084,In_4928,In_3912);
nand U7085 (N_7085,In_1727,In_1756);
or U7086 (N_7086,In_1383,In_378);
nand U7087 (N_7087,In_2473,In_886);
nand U7088 (N_7088,In_993,In_3509);
xor U7089 (N_7089,In_401,In_4225);
nand U7090 (N_7090,In_4615,In_4691);
xnor U7091 (N_7091,In_2787,In_2908);
xnor U7092 (N_7092,In_1960,In_3993);
xor U7093 (N_7093,In_2537,In_316);
or U7094 (N_7094,In_3018,In_3638);
xor U7095 (N_7095,In_1226,In_4783);
and U7096 (N_7096,In_2931,In_3641);
or U7097 (N_7097,In_2286,In_4960);
nor U7098 (N_7098,In_2821,In_4052);
nor U7099 (N_7099,In_2726,In_3099);
nand U7100 (N_7100,In_2014,In_4841);
or U7101 (N_7101,In_4213,In_4261);
or U7102 (N_7102,In_4730,In_3840);
nand U7103 (N_7103,In_2097,In_2118);
or U7104 (N_7104,In_1806,In_136);
nand U7105 (N_7105,In_238,In_835);
nor U7106 (N_7106,In_4333,In_1806);
and U7107 (N_7107,In_2836,In_807);
xor U7108 (N_7108,In_2219,In_2586);
xor U7109 (N_7109,In_3286,In_2907);
or U7110 (N_7110,In_3026,In_619);
and U7111 (N_7111,In_3272,In_795);
or U7112 (N_7112,In_3363,In_69);
and U7113 (N_7113,In_703,In_1714);
nor U7114 (N_7114,In_1321,In_2220);
nor U7115 (N_7115,In_579,In_274);
nor U7116 (N_7116,In_1432,In_2598);
and U7117 (N_7117,In_3373,In_3549);
and U7118 (N_7118,In_1057,In_1597);
nand U7119 (N_7119,In_953,In_801);
and U7120 (N_7120,In_3426,In_3943);
or U7121 (N_7121,In_4405,In_4085);
xnor U7122 (N_7122,In_2152,In_4939);
nand U7123 (N_7123,In_162,In_4796);
and U7124 (N_7124,In_1437,In_3303);
xor U7125 (N_7125,In_1343,In_1586);
nand U7126 (N_7126,In_3793,In_4637);
xnor U7127 (N_7127,In_1280,In_3002);
and U7128 (N_7128,In_4025,In_2000);
and U7129 (N_7129,In_494,In_141);
nor U7130 (N_7130,In_1083,In_3312);
and U7131 (N_7131,In_3064,In_2136);
xor U7132 (N_7132,In_1983,In_3188);
nor U7133 (N_7133,In_2040,In_388);
nand U7134 (N_7134,In_219,In_2655);
xor U7135 (N_7135,In_3693,In_3490);
and U7136 (N_7136,In_2956,In_3369);
xnor U7137 (N_7137,In_1110,In_4749);
nor U7138 (N_7138,In_2939,In_4821);
xor U7139 (N_7139,In_4745,In_461);
nor U7140 (N_7140,In_3721,In_4466);
or U7141 (N_7141,In_1381,In_529);
and U7142 (N_7142,In_4303,In_1056);
or U7143 (N_7143,In_1137,In_673);
and U7144 (N_7144,In_3414,In_3309);
or U7145 (N_7145,In_4576,In_1492);
nand U7146 (N_7146,In_2715,In_4952);
xnor U7147 (N_7147,In_3746,In_1749);
nor U7148 (N_7148,In_4934,In_1025);
xnor U7149 (N_7149,In_3126,In_3850);
nor U7150 (N_7150,In_2274,In_4765);
xor U7151 (N_7151,In_4228,In_4310);
xor U7152 (N_7152,In_1324,In_4701);
and U7153 (N_7153,In_2053,In_1462);
xnor U7154 (N_7154,In_1631,In_1659);
and U7155 (N_7155,In_191,In_2172);
and U7156 (N_7156,In_4062,In_3260);
or U7157 (N_7157,In_1362,In_4021);
nor U7158 (N_7158,In_1019,In_2246);
nand U7159 (N_7159,In_1250,In_3527);
nand U7160 (N_7160,In_4266,In_807);
nand U7161 (N_7161,In_4485,In_2076);
xnor U7162 (N_7162,In_4091,In_1658);
and U7163 (N_7163,In_310,In_1689);
and U7164 (N_7164,In_2743,In_4224);
and U7165 (N_7165,In_2788,In_2829);
and U7166 (N_7166,In_2323,In_3042);
and U7167 (N_7167,In_1713,In_3779);
or U7168 (N_7168,In_702,In_4924);
nand U7169 (N_7169,In_3475,In_3110);
xor U7170 (N_7170,In_325,In_2148);
nand U7171 (N_7171,In_3497,In_1788);
and U7172 (N_7172,In_2760,In_4893);
or U7173 (N_7173,In_3116,In_3315);
and U7174 (N_7174,In_2564,In_3938);
and U7175 (N_7175,In_3663,In_4749);
xor U7176 (N_7176,In_4313,In_1754);
nor U7177 (N_7177,In_933,In_3043);
nand U7178 (N_7178,In_137,In_2383);
nor U7179 (N_7179,In_692,In_3025);
nor U7180 (N_7180,In_4641,In_2079);
or U7181 (N_7181,In_3944,In_3560);
nand U7182 (N_7182,In_28,In_4442);
and U7183 (N_7183,In_735,In_661);
and U7184 (N_7184,In_1709,In_3345);
nand U7185 (N_7185,In_2578,In_1261);
and U7186 (N_7186,In_1185,In_1837);
nor U7187 (N_7187,In_4312,In_650);
nand U7188 (N_7188,In_4249,In_4163);
or U7189 (N_7189,In_1043,In_2489);
or U7190 (N_7190,In_3631,In_1265);
and U7191 (N_7191,In_1560,In_1195);
and U7192 (N_7192,In_2287,In_3052);
or U7193 (N_7193,In_1098,In_3041);
and U7194 (N_7194,In_2542,In_1633);
or U7195 (N_7195,In_2892,In_3489);
xor U7196 (N_7196,In_4530,In_2562);
or U7197 (N_7197,In_3543,In_3832);
nand U7198 (N_7198,In_2277,In_827);
and U7199 (N_7199,In_4570,In_2057);
or U7200 (N_7200,In_2983,In_313);
nor U7201 (N_7201,In_4582,In_1961);
and U7202 (N_7202,In_2272,In_2235);
nand U7203 (N_7203,In_3131,In_1861);
nor U7204 (N_7204,In_3378,In_4304);
nand U7205 (N_7205,In_4466,In_2323);
xnor U7206 (N_7206,In_2123,In_1480);
xnor U7207 (N_7207,In_4709,In_3465);
and U7208 (N_7208,In_3925,In_2234);
and U7209 (N_7209,In_4932,In_1714);
nor U7210 (N_7210,In_2222,In_1810);
nor U7211 (N_7211,In_3066,In_1565);
or U7212 (N_7212,In_2384,In_2523);
xnor U7213 (N_7213,In_3137,In_1712);
nand U7214 (N_7214,In_202,In_3408);
nor U7215 (N_7215,In_372,In_504);
and U7216 (N_7216,In_597,In_2455);
nand U7217 (N_7217,In_4961,In_2368);
xnor U7218 (N_7218,In_1433,In_3638);
xnor U7219 (N_7219,In_391,In_4587);
nand U7220 (N_7220,In_2612,In_1338);
and U7221 (N_7221,In_3666,In_3590);
and U7222 (N_7222,In_1457,In_1011);
nand U7223 (N_7223,In_4162,In_4572);
and U7224 (N_7224,In_1572,In_1485);
nand U7225 (N_7225,In_1592,In_3603);
nor U7226 (N_7226,In_2967,In_2089);
nand U7227 (N_7227,In_4768,In_1208);
and U7228 (N_7228,In_4095,In_2446);
nor U7229 (N_7229,In_4813,In_2020);
and U7230 (N_7230,In_2262,In_2504);
and U7231 (N_7231,In_2789,In_86);
and U7232 (N_7232,In_2628,In_1453);
xor U7233 (N_7233,In_2264,In_4095);
and U7234 (N_7234,In_2397,In_3140);
xnor U7235 (N_7235,In_4360,In_3996);
nor U7236 (N_7236,In_3088,In_2834);
nand U7237 (N_7237,In_2119,In_337);
xnor U7238 (N_7238,In_3397,In_1071);
and U7239 (N_7239,In_2333,In_3170);
nor U7240 (N_7240,In_612,In_3329);
nor U7241 (N_7241,In_3341,In_474);
and U7242 (N_7242,In_3537,In_2276);
and U7243 (N_7243,In_3542,In_3860);
nand U7244 (N_7244,In_2953,In_405);
xor U7245 (N_7245,In_3769,In_885);
and U7246 (N_7246,In_4610,In_469);
or U7247 (N_7247,In_482,In_476);
and U7248 (N_7248,In_1211,In_1388);
xor U7249 (N_7249,In_4153,In_219);
nand U7250 (N_7250,In_2615,In_238);
or U7251 (N_7251,In_4424,In_799);
xor U7252 (N_7252,In_3306,In_654);
xnor U7253 (N_7253,In_4208,In_3234);
nand U7254 (N_7254,In_3055,In_163);
or U7255 (N_7255,In_816,In_4491);
or U7256 (N_7256,In_4167,In_2489);
xor U7257 (N_7257,In_1162,In_1953);
xnor U7258 (N_7258,In_575,In_2338);
nor U7259 (N_7259,In_1117,In_2296);
xnor U7260 (N_7260,In_611,In_2709);
nor U7261 (N_7261,In_2298,In_3025);
nor U7262 (N_7262,In_4905,In_4819);
nand U7263 (N_7263,In_867,In_4056);
nand U7264 (N_7264,In_1973,In_4034);
xor U7265 (N_7265,In_3394,In_3729);
and U7266 (N_7266,In_3348,In_4088);
nand U7267 (N_7267,In_4305,In_1665);
nand U7268 (N_7268,In_2043,In_1283);
nor U7269 (N_7269,In_133,In_4959);
nand U7270 (N_7270,In_1102,In_1438);
or U7271 (N_7271,In_993,In_3422);
and U7272 (N_7272,In_4494,In_4148);
or U7273 (N_7273,In_4982,In_1042);
xnor U7274 (N_7274,In_3692,In_4322);
nand U7275 (N_7275,In_3959,In_55);
nand U7276 (N_7276,In_2201,In_328);
nand U7277 (N_7277,In_631,In_3208);
or U7278 (N_7278,In_2768,In_2432);
and U7279 (N_7279,In_3333,In_3353);
nand U7280 (N_7280,In_4875,In_3198);
nor U7281 (N_7281,In_220,In_4232);
xor U7282 (N_7282,In_4961,In_1742);
nand U7283 (N_7283,In_1332,In_1465);
or U7284 (N_7284,In_2887,In_4092);
or U7285 (N_7285,In_4713,In_2098);
or U7286 (N_7286,In_1119,In_160);
or U7287 (N_7287,In_1349,In_2135);
or U7288 (N_7288,In_3333,In_4465);
and U7289 (N_7289,In_1396,In_1051);
and U7290 (N_7290,In_543,In_790);
or U7291 (N_7291,In_4391,In_2528);
and U7292 (N_7292,In_1118,In_4421);
nor U7293 (N_7293,In_4740,In_4946);
xnor U7294 (N_7294,In_986,In_3525);
nor U7295 (N_7295,In_635,In_536);
nor U7296 (N_7296,In_1838,In_2630);
or U7297 (N_7297,In_1118,In_4606);
and U7298 (N_7298,In_4501,In_4405);
xor U7299 (N_7299,In_122,In_2542);
and U7300 (N_7300,In_4450,In_1943);
and U7301 (N_7301,In_2645,In_933);
and U7302 (N_7302,In_4194,In_4441);
or U7303 (N_7303,In_3871,In_3266);
nand U7304 (N_7304,In_4798,In_3726);
or U7305 (N_7305,In_2826,In_832);
or U7306 (N_7306,In_2696,In_1594);
xnor U7307 (N_7307,In_1366,In_3557);
xor U7308 (N_7308,In_473,In_2284);
xnor U7309 (N_7309,In_962,In_2505);
nor U7310 (N_7310,In_2295,In_4103);
xnor U7311 (N_7311,In_1015,In_2474);
xor U7312 (N_7312,In_4590,In_743);
and U7313 (N_7313,In_1385,In_308);
xor U7314 (N_7314,In_2847,In_3137);
nand U7315 (N_7315,In_1758,In_2973);
xor U7316 (N_7316,In_608,In_637);
and U7317 (N_7317,In_2264,In_1917);
nand U7318 (N_7318,In_1093,In_3261);
xor U7319 (N_7319,In_1362,In_2627);
xor U7320 (N_7320,In_2453,In_4662);
or U7321 (N_7321,In_3961,In_2406);
and U7322 (N_7322,In_3561,In_4273);
xor U7323 (N_7323,In_1933,In_562);
and U7324 (N_7324,In_3566,In_3268);
or U7325 (N_7325,In_3223,In_3388);
nor U7326 (N_7326,In_517,In_2387);
xnor U7327 (N_7327,In_3093,In_1198);
or U7328 (N_7328,In_3833,In_4751);
or U7329 (N_7329,In_3795,In_4795);
xnor U7330 (N_7330,In_3533,In_687);
or U7331 (N_7331,In_810,In_1378);
nand U7332 (N_7332,In_831,In_3440);
xor U7333 (N_7333,In_2762,In_4156);
nor U7334 (N_7334,In_633,In_3634);
nand U7335 (N_7335,In_4668,In_3959);
and U7336 (N_7336,In_3498,In_1437);
nand U7337 (N_7337,In_4691,In_71);
nor U7338 (N_7338,In_1762,In_2632);
xor U7339 (N_7339,In_2886,In_2668);
or U7340 (N_7340,In_1007,In_715);
xor U7341 (N_7341,In_1026,In_138);
nor U7342 (N_7342,In_135,In_2179);
and U7343 (N_7343,In_269,In_2275);
or U7344 (N_7344,In_4251,In_2061);
nand U7345 (N_7345,In_108,In_3385);
and U7346 (N_7346,In_567,In_1131);
or U7347 (N_7347,In_214,In_2463);
nor U7348 (N_7348,In_77,In_3055);
and U7349 (N_7349,In_4,In_3325);
nand U7350 (N_7350,In_4866,In_1148);
nand U7351 (N_7351,In_2244,In_4821);
or U7352 (N_7352,In_2669,In_429);
nor U7353 (N_7353,In_1915,In_1877);
xor U7354 (N_7354,In_1213,In_3707);
or U7355 (N_7355,In_2572,In_1960);
xor U7356 (N_7356,In_4000,In_4963);
nor U7357 (N_7357,In_3358,In_3729);
nor U7358 (N_7358,In_4983,In_2813);
and U7359 (N_7359,In_4562,In_228);
or U7360 (N_7360,In_3268,In_3900);
nand U7361 (N_7361,In_3141,In_3520);
xnor U7362 (N_7362,In_2328,In_363);
and U7363 (N_7363,In_1117,In_397);
nand U7364 (N_7364,In_1338,In_53);
nand U7365 (N_7365,In_3779,In_224);
or U7366 (N_7366,In_4839,In_4853);
xnor U7367 (N_7367,In_971,In_4597);
nor U7368 (N_7368,In_2627,In_4172);
nand U7369 (N_7369,In_127,In_4177);
xnor U7370 (N_7370,In_4479,In_2454);
nand U7371 (N_7371,In_1883,In_2958);
nand U7372 (N_7372,In_4178,In_2406);
or U7373 (N_7373,In_2375,In_3294);
or U7374 (N_7374,In_549,In_2254);
nor U7375 (N_7375,In_1632,In_3642);
nand U7376 (N_7376,In_3550,In_4667);
xnor U7377 (N_7377,In_99,In_3441);
xnor U7378 (N_7378,In_2543,In_1259);
nor U7379 (N_7379,In_4394,In_260);
nand U7380 (N_7380,In_768,In_451);
or U7381 (N_7381,In_421,In_4128);
or U7382 (N_7382,In_2409,In_3624);
xnor U7383 (N_7383,In_2415,In_3848);
or U7384 (N_7384,In_483,In_4990);
xnor U7385 (N_7385,In_4111,In_2296);
nand U7386 (N_7386,In_2081,In_4950);
xor U7387 (N_7387,In_609,In_3599);
and U7388 (N_7388,In_2907,In_2026);
nand U7389 (N_7389,In_2977,In_3579);
or U7390 (N_7390,In_4101,In_1752);
xnor U7391 (N_7391,In_2644,In_2548);
or U7392 (N_7392,In_2230,In_171);
or U7393 (N_7393,In_2346,In_4036);
or U7394 (N_7394,In_551,In_1468);
or U7395 (N_7395,In_834,In_2949);
xnor U7396 (N_7396,In_3782,In_3022);
and U7397 (N_7397,In_1017,In_3473);
or U7398 (N_7398,In_2162,In_3422);
nor U7399 (N_7399,In_4843,In_4001);
nand U7400 (N_7400,In_3603,In_3768);
or U7401 (N_7401,In_4107,In_3923);
xor U7402 (N_7402,In_2502,In_2009);
or U7403 (N_7403,In_2376,In_3282);
nand U7404 (N_7404,In_604,In_108);
or U7405 (N_7405,In_3729,In_4595);
xnor U7406 (N_7406,In_1491,In_2654);
and U7407 (N_7407,In_3675,In_3120);
nor U7408 (N_7408,In_4115,In_1583);
and U7409 (N_7409,In_4098,In_2760);
xor U7410 (N_7410,In_2450,In_2614);
and U7411 (N_7411,In_856,In_1199);
xnor U7412 (N_7412,In_1827,In_275);
xor U7413 (N_7413,In_3732,In_107);
and U7414 (N_7414,In_712,In_3750);
nor U7415 (N_7415,In_4261,In_2730);
or U7416 (N_7416,In_2896,In_4599);
nor U7417 (N_7417,In_3794,In_2597);
nand U7418 (N_7418,In_3387,In_2206);
and U7419 (N_7419,In_4889,In_3209);
xor U7420 (N_7420,In_1203,In_2930);
xnor U7421 (N_7421,In_3434,In_3412);
xnor U7422 (N_7422,In_4189,In_4954);
nand U7423 (N_7423,In_2314,In_719);
and U7424 (N_7424,In_2061,In_1490);
nand U7425 (N_7425,In_3331,In_788);
or U7426 (N_7426,In_4266,In_2274);
and U7427 (N_7427,In_323,In_2504);
and U7428 (N_7428,In_830,In_2140);
nand U7429 (N_7429,In_1689,In_1716);
and U7430 (N_7430,In_1899,In_3045);
nor U7431 (N_7431,In_1693,In_3245);
nand U7432 (N_7432,In_3399,In_3805);
or U7433 (N_7433,In_4269,In_2079);
nand U7434 (N_7434,In_118,In_627);
nand U7435 (N_7435,In_4543,In_2602);
xnor U7436 (N_7436,In_1702,In_1188);
nand U7437 (N_7437,In_1263,In_2575);
and U7438 (N_7438,In_2517,In_1275);
or U7439 (N_7439,In_2089,In_1184);
or U7440 (N_7440,In_2606,In_4379);
and U7441 (N_7441,In_4047,In_3704);
nor U7442 (N_7442,In_4728,In_1266);
nor U7443 (N_7443,In_3841,In_358);
or U7444 (N_7444,In_4628,In_1542);
or U7445 (N_7445,In_1204,In_1330);
nand U7446 (N_7446,In_2934,In_779);
or U7447 (N_7447,In_4691,In_4046);
xnor U7448 (N_7448,In_542,In_1203);
nor U7449 (N_7449,In_4706,In_2547);
nand U7450 (N_7450,In_3573,In_3470);
and U7451 (N_7451,In_2674,In_2741);
or U7452 (N_7452,In_3647,In_639);
or U7453 (N_7453,In_4970,In_3115);
nor U7454 (N_7454,In_166,In_4575);
nor U7455 (N_7455,In_4633,In_656);
nand U7456 (N_7456,In_3896,In_262);
or U7457 (N_7457,In_2576,In_1373);
and U7458 (N_7458,In_286,In_3751);
or U7459 (N_7459,In_3530,In_3491);
xor U7460 (N_7460,In_1130,In_3834);
nand U7461 (N_7461,In_3210,In_875);
and U7462 (N_7462,In_4329,In_232);
xnor U7463 (N_7463,In_3305,In_1831);
or U7464 (N_7464,In_310,In_1278);
nor U7465 (N_7465,In_1360,In_1073);
xor U7466 (N_7466,In_1284,In_2395);
nand U7467 (N_7467,In_1229,In_554);
xor U7468 (N_7468,In_4870,In_2841);
or U7469 (N_7469,In_3557,In_2069);
or U7470 (N_7470,In_4477,In_4553);
nand U7471 (N_7471,In_2294,In_510);
nor U7472 (N_7472,In_2247,In_2614);
or U7473 (N_7473,In_319,In_4004);
and U7474 (N_7474,In_3738,In_1479);
nand U7475 (N_7475,In_1473,In_1093);
xnor U7476 (N_7476,In_3350,In_3729);
or U7477 (N_7477,In_3369,In_4224);
or U7478 (N_7478,In_3756,In_4486);
or U7479 (N_7479,In_3756,In_656);
nor U7480 (N_7480,In_3523,In_4176);
nor U7481 (N_7481,In_4418,In_2029);
nand U7482 (N_7482,In_1172,In_1061);
or U7483 (N_7483,In_2940,In_3733);
and U7484 (N_7484,In_380,In_3791);
nor U7485 (N_7485,In_2724,In_4739);
and U7486 (N_7486,In_187,In_4211);
or U7487 (N_7487,In_4049,In_322);
xor U7488 (N_7488,In_4431,In_1716);
or U7489 (N_7489,In_4807,In_1127);
nand U7490 (N_7490,In_2107,In_2212);
or U7491 (N_7491,In_4423,In_4453);
and U7492 (N_7492,In_4419,In_942);
nand U7493 (N_7493,In_75,In_2306);
xor U7494 (N_7494,In_2029,In_442);
xnor U7495 (N_7495,In_2833,In_1917);
or U7496 (N_7496,In_4389,In_1320);
xnor U7497 (N_7497,In_1425,In_4940);
nor U7498 (N_7498,In_1599,In_821);
or U7499 (N_7499,In_972,In_1987);
and U7500 (N_7500,In_2785,In_813);
or U7501 (N_7501,In_3484,In_2086);
xnor U7502 (N_7502,In_2664,In_31);
nor U7503 (N_7503,In_313,In_15);
xor U7504 (N_7504,In_2962,In_991);
nand U7505 (N_7505,In_362,In_3938);
and U7506 (N_7506,In_4627,In_1167);
xor U7507 (N_7507,In_3307,In_1318);
nor U7508 (N_7508,In_2967,In_1039);
nor U7509 (N_7509,In_349,In_3908);
nand U7510 (N_7510,In_4274,In_2905);
and U7511 (N_7511,In_4349,In_442);
nor U7512 (N_7512,In_2254,In_3097);
xnor U7513 (N_7513,In_1876,In_2526);
nand U7514 (N_7514,In_1452,In_857);
nand U7515 (N_7515,In_988,In_1647);
and U7516 (N_7516,In_4102,In_3749);
xnor U7517 (N_7517,In_661,In_2616);
nand U7518 (N_7518,In_1223,In_4793);
xnor U7519 (N_7519,In_3087,In_3585);
nand U7520 (N_7520,In_2397,In_1723);
nand U7521 (N_7521,In_3019,In_2424);
nand U7522 (N_7522,In_3587,In_3570);
and U7523 (N_7523,In_4395,In_3677);
nor U7524 (N_7524,In_2824,In_3478);
nand U7525 (N_7525,In_3697,In_2617);
nand U7526 (N_7526,In_3190,In_2069);
and U7527 (N_7527,In_4122,In_2882);
or U7528 (N_7528,In_3847,In_2778);
nand U7529 (N_7529,In_1811,In_589);
xor U7530 (N_7530,In_2297,In_4642);
and U7531 (N_7531,In_4010,In_4473);
xnor U7532 (N_7532,In_3606,In_99);
nor U7533 (N_7533,In_3109,In_2547);
xnor U7534 (N_7534,In_1694,In_3225);
xor U7535 (N_7535,In_4142,In_2335);
or U7536 (N_7536,In_4034,In_1797);
nand U7537 (N_7537,In_4436,In_3603);
and U7538 (N_7538,In_4365,In_3466);
xor U7539 (N_7539,In_2487,In_2387);
nor U7540 (N_7540,In_1486,In_2203);
xor U7541 (N_7541,In_3080,In_2657);
and U7542 (N_7542,In_76,In_1638);
xnor U7543 (N_7543,In_1712,In_2814);
or U7544 (N_7544,In_1527,In_3937);
nand U7545 (N_7545,In_4981,In_3581);
and U7546 (N_7546,In_1648,In_3161);
nand U7547 (N_7547,In_1562,In_38);
nand U7548 (N_7548,In_11,In_3203);
nand U7549 (N_7549,In_2456,In_1708);
xnor U7550 (N_7550,In_3016,In_3098);
or U7551 (N_7551,In_572,In_3201);
xnor U7552 (N_7552,In_4918,In_2634);
and U7553 (N_7553,In_294,In_1400);
xor U7554 (N_7554,In_1990,In_1371);
and U7555 (N_7555,In_2100,In_4730);
nor U7556 (N_7556,In_2214,In_281);
nor U7557 (N_7557,In_3889,In_4169);
xnor U7558 (N_7558,In_900,In_3631);
or U7559 (N_7559,In_1682,In_3173);
and U7560 (N_7560,In_2600,In_4501);
nor U7561 (N_7561,In_623,In_2526);
nand U7562 (N_7562,In_4040,In_2184);
nand U7563 (N_7563,In_3278,In_4109);
nand U7564 (N_7564,In_4188,In_4780);
nor U7565 (N_7565,In_1256,In_1000);
nand U7566 (N_7566,In_992,In_2279);
xor U7567 (N_7567,In_1474,In_1357);
nor U7568 (N_7568,In_4710,In_1888);
and U7569 (N_7569,In_3173,In_4617);
nor U7570 (N_7570,In_908,In_3231);
nand U7571 (N_7571,In_245,In_863);
xor U7572 (N_7572,In_1480,In_1146);
nand U7573 (N_7573,In_4361,In_1705);
xnor U7574 (N_7574,In_4409,In_97);
nand U7575 (N_7575,In_727,In_554);
xor U7576 (N_7576,In_4864,In_1439);
xnor U7577 (N_7577,In_3978,In_999);
xnor U7578 (N_7578,In_3972,In_1660);
and U7579 (N_7579,In_3261,In_2569);
nor U7580 (N_7580,In_1586,In_1325);
nor U7581 (N_7581,In_2426,In_609);
or U7582 (N_7582,In_4055,In_3093);
or U7583 (N_7583,In_855,In_2805);
and U7584 (N_7584,In_2715,In_1740);
or U7585 (N_7585,In_1602,In_3485);
or U7586 (N_7586,In_4479,In_1335);
or U7587 (N_7587,In_2730,In_2505);
and U7588 (N_7588,In_4249,In_4793);
or U7589 (N_7589,In_2509,In_1086);
nor U7590 (N_7590,In_2093,In_1818);
nand U7591 (N_7591,In_1549,In_4293);
xor U7592 (N_7592,In_622,In_1174);
nor U7593 (N_7593,In_34,In_1955);
xor U7594 (N_7594,In_4539,In_1502);
xnor U7595 (N_7595,In_4322,In_1698);
and U7596 (N_7596,In_3132,In_1020);
nand U7597 (N_7597,In_1696,In_3962);
nand U7598 (N_7598,In_3161,In_4371);
and U7599 (N_7599,In_2189,In_4851);
nand U7600 (N_7600,In_2167,In_4611);
or U7601 (N_7601,In_2782,In_4262);
xnor U7602 (N_7602,In_561,In_68);
nand U7603 (N_7603,In_3237,In_76);
and U7604 (N_7604,In_41,In_2111);
xnor U7605 (N_7605,In_4464,In_1700);
nor U7606 (N_7606,In_4093,In_4106);
nor U7607 (N_7607,In_4536,In_1786);
and U7608 (N_7608,In_3014,In_507);
and U7609 (N_7609,In_3488,In_4114);
xnor U7610 (N_7610,In_1711,In_1338);
nand U7611 (N_7611,In_1867,In_331);
nand U7612 (N_7612,In_1119,In_4962);
or U7613 (N_7613,In_2570,In_3147);
nor U7614 (N_7614,In_4688,In_681);
nor U7615 (N_7615,In_566,In_969);
nor U7616 (N_7616,In_1206,In_1517);
nor U7617 (N_7617,In_4348,In_3862);
nor U7618 (N_7618,In_3306,In_1770);
nor U7619 (N_7619,In_4421,In_2591);
xnor U7620 (N_7620,In_3620,In_1049);
or U7621 (N_7621,In_1979,In_3481);
nor U7622 (N_7622,In_4978,In_780);
nor U7623 (N_7623,In_1018,In_4966);
nor U7624 (N_7624,In_2669,In_3700);
and U7625 (N_7625,In_1387,In_619);
nand U7626 (N_7626,In_3268,In_3161);
xor U7627 (N_7627,In_3506,In_3191);
or U7628 (N_7628,In_4207,In_814);
xor U7629 (N_7629,In_4589,In_758);
or U7630 (N_7630,In_579,In_4514);
nor U7631 (N_7631,In_2171,In_2556);
or U7632 (N_7632,In_3239,In_959);
and U7633 (N_7633,In_10,In_192);
and U7634 (N_7634,In_885,In_2948);
xor U7635 (N_7635,In_1471,In_4510);
nand U7636 (N_7636,In_1222,In_1436);
nor U7637 (N_7637,In_1926,In_3144);
xor U7638 (N_7638,In_989,In_4171);
and U7639 (N_7639,In_2881,In_2519);
nor U7640 (N_7640,In_4844,In_2224);
nor U7641 (N_7641,In_4879,In_2989);
or U7642 (N_7642,In_312,In_2642);
or U7643 (N_7643,In_1110,In_3374);
or U7644 (N_7644,In_2800,In_3599);
nand U7645 (N_7645,In_731,In_1390);
nand U7646 (N_7646,In_1035,In_1563);
or U7647 (N_7647,In_776,In_256);
and U7648 (N_7648,In_4722,In_4252);
and U7649 (N_7649,In_488,In_3781);
or U7650 (N_7650,In_4949,In_2569);
xnor U7651 (N_7651,In_2178,In_1760);
nor U7652 (N_7652,In_2365,In_4090);
nand U7653 (N_7653,In_3400,In_1297);
or U7654 (N_7654,In_1881,In_3983);
xnor U7655 (N_7655,In_1495,In_311);
nand U7656 (N_7656,In_2951,In_1132);
nor U7657 (N_7657,In_2647,In_2859);
nor U7658 (N_7658,In_3994,In_4781);
nand U7659 (N_7659,In_43,In_4445);
nor U7660 (N_7660,In_711,In_371);
or U7661 (N_7661,In_2276,In_4325);
xor U7662 (N_7662,In_2877,In_2945);
xnor U7663 (N_7663,In_423,In_2775);
nor U7664 (N_7664,In_2114,In_3310);
nand U7665 (N_7665,In_4944,In_3140);
nand U7666 (N_7666,In_1082,In_3301);
and U7667 (N_7667,In_2738,In_3990);
or U7668 (N_7668,In_4347,In_3511);
or U7669 (N_7669,In_1919,In_1474);
and U7670 (N_7670,In_4261,In_4456);
nand U7671 (N_7671,In_486,In_552);
and U7672 (N_7672,In_1521,In_801);
and U7673 (N_7673,In_549,In_2553);
and U7674 (N_7674,In_2613,In_162);
nand U7675 (N_7675,In_1620,In_4062);
and U7676 (N_7676,In_1542,In_923);
xnor U7677 (N_7677,In_4621,In_3167);
nand U7678 (N_7678,In_4549,In_4338);
xor U7679 (N_7679,In_2617,In_23);
xnor U7680 (N_7680,In_2816,In_2269);
or U7681 (N_7681,In_4073,In_3808);
and U7682 (N_7682,In_1075,In_2202);
nand U7683 (N_7683,In_2572,In_646);
nor U7684 (N_7684,In_3182,In_4663);
xnor U7685 (N_7685,In_2324,In_1258);
nor U7686 (N_7686,In_3717,In_3627);
xnor U7687 (N_7687,In_1905,In_2216);
xor U7688 (N_7688,In_2904,In_856);
nor U7689 (N_7689,In_1857,In_306);
nor U7690 (N_7690,In_1269,In_692);
xnor U7691 (N_7691,In_3979,In_4977);
or U7692 (N_7692,In_4044,In_261);
nor U7693 (N_7693,In_764,In_529);
and U7694 (N_7694,In_3476,In_2561);
and U7695 (N_7695,In_412,In_754);
nand U7696 (N_7696,In_1936,In_4806);
and U7697 (N_7697,In_4603,In_2987);
nor U7698 (N_7698,In_3580,In_4562);
nand U7699 (N_7699,In_3624,In_4179);
or U7700 (N_7700,In_1424,In_4902);
nor U7701 (N_7701,In_4018,In_552);
nand U7702 (N_7702,In_1121,In_3274);
nor U7703 (N_7703,In_1993,In_1884);
or U7704 (N_7704,In_922,In_2645);
and U7705 (N_7705,In_2022,In_2330);
nor U7706 (N_7706,In_3134,In_4591);
and U7707 (N_7707,In_4506,In_3219);
nand U7708 (N_7708,In_3853,In_1024);
and U7709 (N_7709,In_12,In_4693);
nand U7710 (N_7710,In_4886,In_3552);
or U7711 (N_7711,In_1840,In_3601);
nor U7712 (N_7712,In_367,In_1223);
or U7713 (N_7713,In_2581,In_3400);
nand U7714 (N_7714,In_3214,In_1589);
xnor U7715 (N_7715,In_1681,In_2412);
and U7716 (N_7716,In_1317,In_4893);
or U7717 (N_7717,In_2631,In_2658);
xor U7718 (N_7718,In_450,In_1675);
nor U7719 (N_7719,In_1475,In_3209);
and U7720 (N_7720,In_2414,In_1952);
nand U7721 (N_7721,In_2612,In_1736);
nand U7722 (N_7722,In_1461,In_4316);
and U7723 (N_7723,In_2274,In_725);
nand U7724 (N_7724,In_4638,In_4858);
nor U7725 (N_7725,In_3721,In_933);
nand U7726 (N_7726,In_4119,In_933);
or U7727 (N_7727,In_2524,In_3181);
nand U7728 (N_7728,In_2233,In_9);
nand U7729 (N_7729,In_1401,In_4527);
and U7730 (N_7730,In_309,In_3395);
xnor U7731 (N_7731,In_990,In_335);
xor U7732 (N_7732,In_1172,In_3134);
nor U7733 (N_7733,In_2763,In_4569);
or U7734 (N_7734,In_4149,In_987);
or U7735 (N_7735,In_4860,In_4630);
or U7736 (N_7736,In_3837,In_227);
nand U7737 (N_7737,In_3958,In_3003);
nor U7738 (N_7738,In_1723,In_4631);
and U7739 (N_7739,In_4079,In_289);
nand U7740 (N_7740,In_2327,In_1834);
and U7741 (N_7741,In_3186,In_1866);
nand U7742 (N_7742,In_2193,In_2753);
and U7743 (N_7743,In_4872,In_2374);
and U7744 (N_7744,In_3495,In_4405);
xnor U7745 (N_7745,In_4658,In_1564);
and U7746 (N_7746,In_219,In_4668);
nand U7747 (N_7747,In_940,In_4509);
and U7748 (N_7748,In_750,In_1244);
nand U7749 (N_7749,In_253,In_3496);
and U7750 (N_7750,In_3970,In_3571);
or U7751 (N_7751,In_3715,In_398);
and U7752 (N_7752,In_898,In_3155);
or U7753 (N_7753,In_485,In_4559);
and U7754 (N_7754,In_3421,In_4498);
nand U7755 (N_7755,In_4787,In_1787);
nor U7756 (N_7756,In_3767,In_601);
and U7757 (N_7757,In_416,In_2856);
or U7758 (N_7758,In_3129,In_3913);
or U7759 (N_7759,In_1058,In_2103);
nand U7760 (N_7760,In_890,In_2025);
xnor U7761 (N_7761,In_2249,In_99);
and U7762 (N_7762,In_11,In_4964);
or U7763 (N_7763,In_4212,In_4075);
xnor U7764 (N_7764,In_4576,In_3028);
xnor U7765 (N_7765,In_16,In_2462);
and U7766 (N_7766,In_701,In_365);
xor U7767 (N_7767,In_2879,In_2248);
xor U7768 (N_7768,In_3434,In_411);
nand U7769 (N_7769,In_2060,In_86);
xor U7770 (N_7770,In_4505,In_1903);
xnor U7771 (N_7771,In_4354,In_4082);
nand U7772 (N_7772,In_1805,In_696);
xnor U7773 (N_7773,In_4096,In_3697);
and U7774 (N_7774,In_1561,In_4253);
xor U7775 (N_7775,In_160,In_1882);
nor U7776 (N_7776,In_219,In_531);
or U7777 (N_7777,In_2357,In_1369);
nand U7778 (N_7778,In_2133,In_2576);
nor U7779 (N_7779,In_4574,In_1889);
nor U7780 (N_7780,In_968,In_1014);
or U7781 (N_7781,In_3032,In_1140);
nor U7782 (N_7782,In_2415,In_1172);
xor U7783 (N_7783,In_955,In_965);
or U7784 (N_7784,In_1150,In_2381);
and U7785 (N_7785,In_339,In_4347);
nand U7786 (N_7786,In_716,In_2157);
nor U7787 (N_7787,In_1350,In_1636);
nand U7788 (N_7788,In_3856,In_4131);
nand U7789 (N_7789,In_4228,In_70);
nand U7790 (N_7790,In_4027,In_260);
xnor U7791 (N_7791,In_113,In_4953);
xor U7792 (N_7792,In_339,In_2602);
xnor U7793 (N_7793,In_4411,In_1279);
nor U7794 (N_7794,In_4668,In_1099);
and U7795 (N_7795,In_2866,In_3181);
and U7796 (N_7796,In_4903,In_2343);
nor U7797 (N_7797,In_3572,In_3110);
nand U7798 (N_7798,In_1015,In_3369);
nand U7799 (N_7799,In_3846,In_109);
nand U7800 (N_7800,In_1171,In_3704);
and U7801 (N_7801,In_2869,In_774);
and U7802 (N_7802,In_4302,In_2232);
xor U7803 (N_7803,In_3695,In_245);
nor U7804 (N_7804,In_2298,In_4648);
and U7805 (N_7805,In_275,In_2442);
xor U7806 (N_7806,In_1804,In_652);
xor U7807 (N_7807,In_4132,In_3706);
nor U7808 (N_7808,In_3697,In_2523);
nand U7809 (N_7809,In_2612,In_3168);
or U7810 (N_7810,In_4872,In_1915);
xnor U7811 (N_7811,In_3807,In_2698);
and U7812 (N_7812,In_3665,In_881);
and U7813 (N_7813,In_1616,In_459);
nor U7814 (N_7814,In_2961,In_4469);
and U7815 (N_7815,In_914,In_26);
nor U7816 (N_7816,In_1461,In_4794);
nor U7817 (N_7817,In_1830,In_3650);
xnor U7818 (N_7818,In_2302,In_4007);
xor U7819 (N_7819,In_1735,In_2156);
and U7820 (N_7820,In_2865,In_3992);
xnor U7821 (N_7821,In_729,In_1096);
nor U7822 (N_7822,In_3824,In_4485);
xnor U7823 (N_7823,In_4040,In_3969);
and U7824 (N_7824,In_3224,In_175);
nand U7825 (N_7825,In_1655,In_2319);
xor U7826 (N_7826,In_3155,In_3373);
and U7827 (N_7827,In_3215,In_4152);
nand U7828 (N_7828,In_1290,In_4272);
and U7829 (N_7829,In_914,In_2994);
or U7830 (N_7830,In_3109,In_1066);
or U7831 (N_7831,In_4436,In_3662);
and U7832 (N_7832,In_63,In_4954);
nand U7833 (N_7833,In_1988,In_4437);
nand U7834 (N_7834,In_3760,In_4643);
xor U7835 (N_7835,In_3843,In_3791);
or U7836 (N_7836,In_4181,In_351);
xnor U7837 (N_7837,In_593,In_16);
and U7838 (N_7838,In_4352,In_2366);
nor U7839 (N_7839,In_2328,In_1658);
nand U7840 (N_7840,In_2257,In_2377);
nand U7841 (N_7841,In_1738,In_902);
xnor U7842 (N_7842,In_2091,In_977);
and U7843 (N_7843,In_1778,In_4945);
xnor U7844 (N_7844,In_437,In_1713);
nand U7845 (N_7845,In_755,In_3044);
nor U7846 (N_7846,In_1617,In_4659);
or U7847 (N_7847,In_1814,In_4022);
xor U7848 (N_7848,In_2547,In_348);
nor U7849 (N_7849,In_1668,In_465);
xor U7850 (N_7850,In_1363,In_1298);
or U7851 (N_7851,In_429,In_4403);
xor U7852 (N_7852,In_4266,In_627);
or U7853 (N_7853,In_550,In_2891);
and U7854 (N_7854,In_4833,In_4722);
nor U7855 (N_7855,In_4904,In_3939);
and U7856 (N_7856,In_3458,In_2742);
or U7857 (N_7857,In_2878,In_167);
nor U7858 (N_7858,In_1277,In_3060);
nand U7859 (N_7859,In_1605,In_3331);
or U7860 (N_7860,In_1606,In_1349);
and U7861 (N_7861,In_1725,In_285);
nand U7862 (N_7862,In_1622,In_2534);
nand U7863 (N_7863,In_3275,In_1822);
nand U7864 (N_7864,In_281,In_384);
and U7865 (N_7865,In_3584,In_818);
nand U7866 (N_7866,In_2455,In_291);
nand U7867 (N_7867,In_3138,In_906);
and U7868 (N_7868,In_1484,In_226);
nor U7869 (N_7869,In_1516,In_4024);
and U7870 (N_7870,In_3962,In_1496);
nand U7871 (N_7871,In_3262,In_1359);
xor U7872 (N_7872,In_2055,In_1292);
nand U7873 (N_7873,In_999,In_3860);
or U7874 (N_7874,In_2486,In_756);
and U7875 (N_7875,In_4866,In_1933);
and U7876 (N_7876,In_4860,In_2309);
and U7877 (N_7877,In_3730,In_2862);
nand U7878 (N_7878,In_839,In_2863);
nor U7879 (N_7879,In_4749,In_1673);
or U7880 (N_7880,In_371,In_1717);
and U7881 (N_7881,In_3734,In_1359);
or U7882 (N_7882,In_647,In_4092);
nand U7883 (N_7883,In_1946,In_2135);
nor U7884 (N_7884,In_4913,In_2117);
nor U7885 (N_7885,In_1985,In_4033);
or U7886 (N_7886,In_1730,In_71);
and U7887 (N_7887,In_4047,In_2602);
or U7888 (N_7888,In_981,In_4989);
nor U7889 (N_7889,In_4202,In_4351);
nand U7890 (N_7890,In_221,In_4043);
nand U7891 (N_7891,In_3593,In_4979);
nor U7892 (N_7892,In_312,In_1848);
and U7893 (N_7893,In_4294,In_4534);
nand U7894 (N_7894,In_1915,In_1589);
xor U7895 (N_7895,In_2355,In_3593);
and U7896 (N_7896,In_4903,In_1493);
nand U7897 (N_7897,In_3038,In_4929);
nand U7898 (N_7898,In_3761,In_2740);
nand U7899 (N_7899,In_2269,In_4883);
nand U7900 (N_7900,In_689,In_4687);
and U7901 (N_7901,In_3822,In_3457);
or U7902 (N_7902,In_3780,In_2692);
nand U7903 (N_7903,In_1043,In_578);
nand U7904 (N_7904,In_1635,In_1417);
or U7905 (N_7905,In_2495,In_3085);
or U7906 (N_7906,In_4735,In_2082);
nor U7907 (N_7907,In_4424,In_3320);
or U7908 (N_7908,In_2099,In_854);
xnor U7909 (N_7909,In_2113,In_589);
nand U7910 (N_7910,In_4035,In_2555);
xnor U7911 (N_7911,In_1676,In_681);
nand U7912 (N_7912,In_4097,In_1734);
and U7913 (N_7913,In_3724,In_1075);
or U7914 (N_7914,In_4166,In_1325);
or U7915 (N_7915,In_356,In_2624);
and U7916 (N_7916,In_2338,In_3408);
and U7917 (N_7917,In_505,In_2847);
and U7918 (N_7918,In_960,In_1059);
nor U7919 (N_7919,In_3970,In_4307);
or U7920 (N_7920,In_2750,In_4613);
nor U7921 (N_7921,In_463,In_3983);
or U7922 (N_7922,In_3674,In_587);
nor U7923 (N_7923,In_255,In_3857);
or U7924 (N_7924,In_3257,In_2921);
nor U7925 (N_7925,In_3107,In_3637);
and U7926 (N_7926,In_1379,In_1840);
or U7927 (N_7927,In_4348,In_3760);
nand U7928 (N_7928,In_4317,In_1734);
or U7929 (N_7929,In_4794,In_3422);
nor U7930 (N_7930,In_1281,In_4706);
and U7931 (N_7931,In_4566,In_882);
nand U7932 (N_7932,In_27,In_288);
and U7933 (N_7933,In_1646,In_1289);
or U7934 (N_7934,In_3988,In_1304);
xnor U7935 (N_7935,In_3897,In_4195);
and U7936 (N_7936,In_433,In_1290);
nor U7937 (N_7937,In_4505,In_308);
or U7938 (N_7938,In_2383,In_4419);
nand U7939 (N_7939,In_4659,In_3678);
nand U7940 (N_7940,In_4053,In_3879);
or U7941 (N_7941,In_1645,In_1425);
nor U7942 (N_7942,In_838,In_3109);
or U7943 (N_7943,In_687,In_2924);
nand U7944 (N_7944,In_4497,In_4596);
xor U7945 (N_7945,In_3454,In_1573);
or U7946 (N_7946,In_1858,In_3875);
or U7947 (N_7947,In_2797,In_1475);
xor U7948 (N_7948,In_3917,In_865);
nor U7949 (N_7949,In_413,In_3676);
xnor U7950 (N_7950,In_3482,In_4903);
nand U7951 (N_7951,In_4176,In_923);
or U7952 (N_7952,In_3914,In_3326);
or U7953 (N_7953,In_4364,In_3403);
or U7954 (N_7954,In_2113,In_1937);
nand U7955 (N_7955,In_3190,In_3937);
nor U7956 (N_7956,In_175,In_4114);
and U7957 (N_7957,In_156,In_1622);
nand U7958 (N_7958,In_1843,In_840);
nand U7959 (N_7959,In_3490,In_4322);
nor U7960 (N_7960,In_4631,In_4976);
or U7961 (N_7961,In_1316,In_2848);
nor U7962 (N_7962,In_2011,In_1519);
or U7963 (N_7963,In_736,In_4808);
xor U7964 (N_7964,In_1823,In_2979);
or U7965 (N_7965,In_2939,In_1314);
nand U7966 (N_7966,In_1249,In_4945);
nand U7967 (N_7967,In_4276,In_3245);
nand U7968 (N_7968,In_68,In_711);
and U7969 (N_7969,In_4771,In_2723);
nand U7970 (N_7970,In_2169,In_2213);
or U7971 (N_7971,In_3722,In_3444);
xnor U7972 (N_7972,In_2958,In_543);
and U7973 (N_7973,In_1772,In_691);
or U7974 (N_7974,In_3941,In_185);
nand U7975 (N_7975,In_969,In_3260);
nor U7976 (N_7976,In_3960,In_3445);
xor U7977 (N_7977,In_266,In_3261);
and U7978 (N_7978,In_1831,In_2784);
and U7979 (N_7979,In_3819,In_1026);
xnor U7980 (N_7980,In_930,In_312);
xor U7981 (N_7981,In_2373,In_3053);
and U7982 (N_7982,In_1728,In_2308);
nand U7983 (N_7983,In_323,In_931);
and U7984 (N_7984,In_909,In_1843);
and U7985 (N_7985,In_1383,In_577);
nand U7986 (N_7986,In_839,In_3140);
and U7987 (N_7987,In_1864,In_400);
nand U7988 (N_7988,In_2365,In_1992);
nand U7989 (N_7989,In_1684,In_336);
nand U7990 (N_7990,In_1625,In_4527);
nand U7991 (N_7991,In_4414,In_2071);
nand U7992 (N_7992,In_1737,In_647);
or U7993 (N_7993,In_2093,In_4314);
nor U7994 (N_7994,In_4164,In_3056);
or U7995 (N_7995,In_510,In_319);
and U7996 (N_7996,In_1187,In_970);
xor U7997 (N_7997,In_3564,In_3468);
and U7998 (N_7998,In_209,In_4829);
and U7999 (N_7999,In_3732,In_3841);
xnor U8000 (N_8000,In_2158,In_1253);
xor U8001 (N_8001,In_4511,In_3212);
nand U8002 (N_8002,In_308,In_735);
nand U8003 (N_8003,In_639,In_1447);
nor U8004 (N_8004,In_2328,In_4340);
xor U8005 (N_8005,In_337,In_1516);
nand U8006 (N_8006,In_2791,In_4865);
nand U8007 (N_8007,In_4926,In_757);
nand U8008 (N_8008,In_4775,In_899);
or U8009 (N_8009,In_544,In_1387);
or U8010 (N_8010,In_1744,In_4690);
nor U8011 (N_8011,In_1752,In_2415);
nand U8012 (N_8012,In_3764,In_446);
nor U8013 (N_8013,In_4043,In_2219);
or U8014 (N_8014,In_207,In_3332);
nor U8015 (N_8015,In_2474,In_4035);
nand U8016 (N_8016,In_1483,In_2650);
xor U8017 (N_8017,In_1548,In_2903);
nor U8018 (N_8018,In_487,In_2614);
nor U8019 (N_8019,In_189,In_631);
xnor U8020 (N_8020,In_3063,In_2367);
xnor U8021 (N_8021,In_3008,In_956);
xnor U8022 (N_8022,In_1886,In_3324);
xnor U8023 (N_8023,In_1466,In_3316);
nor U8024 (N_8024,In_3727,In_1531);
and U8025 (N_8025,In_850,In_2658);
or U8026 (N_8026,In_1790,In_2618);
nor U8027 (N_8027,In_4893,In_2528);
nor U8028 (N_8028,In_3427,In_3637);
or U8029 (N_8029,In_4316,In_4243);
and U8030 (N_8030,In_4534,In_102);
xor U8031 (N_8031,In_3175,In_3188);
xor U8032 (N_8032,In_4838,In_4593);
nand U8033 (N_8033,In_1487,In_4529);
nand U8034 (N_8034,In_1264,In_1832);
nand U8035 (N_8035,In_826,In_2799);
or U8036 (N_8036,In_4063,In_1669);
nand U8037 (N_8037,In_1112,In_4719);
nor U8038 (N_8038,In_4375,In_102);
and U8039 (N_8039,In_1856,In_1271);
xor U8040 (N_8040,In_3609,In_2558);
nor U8041 (N_8041,In_1479,In_2690);
xnor U8042 (N_8042,In_1490,In_4524);
and U8043 (N_8043,In_4630,In_4500);
and U8044 (N_8044,In_250,In_2896);
xnor U8045 (N_8045,In_3004,In_2345);
and U8046 (N_8046,In_1367,In_2822);
or U8047 (N_8047,In_242,In_4596);
nor U8048 (N_8048,In_2644,In_4830);
and U8049 (N_8049,In_4306,In_981);
nor U8050 (N_8050,In_1886,In_2735);
nand U8051 (N_8051,In_1767,In_916);
and U8052 (N_8052,In_1762,In_2768);
and U8053 (N_8053,In_736,In_1001);
xor U8054 (N_8054,In_3327,In_3492);
and U8055 (N_8055,In_2865,In_565);
and U8056 (N_8056,In_859,In_4391);
or U8057 (N_8057,In_901,In_2728);
nand U8058 (N_8058,In_4314,In_3662);
nor U8059 (N_8059,In_858,In_4007);
nor U8060 (N_8060,In_188,In_1740);
or U8061 (N_8061,In_926,In_4699);
or U8062 (N_8062,In_4461,In_2551);
xor U8063 (N_8063,In_236,In_1826);
or U8064 (N_8064,In_4665,In_1996);
xor U8065 (N_8065,In_4857,In_3628);
nor U8066 (N_8066,In_1121,In_4386);
xor U8067 (N_8067,In_2015,In_735);
or U8068 (N_8068,In_2036,In_1251);
and U8069 (N_8069,In_4727,In_1307);
nand U8070 (N_8070,In_683,In_3314);
xnor U8071 (N_8071,In_1151,In_4847);
nand U8072 (N_8072,In_4987,In_3874);
xor U8073 (N_8073,In_4,In_553);
and U8074 (N_8074,In_2700,In_3157);
nand U8075 (N_8075,In_4856,In_2536);
nor U8076 (N_8076,In_2241,In_4558);
xor U8077 (N_8077,In_2995,In_1803);
and U8078 (N_8078,In_3231,In_741);
and U8079 (N_8079,In_4563,In_3635);
nand U8080 (N_8080,In_3427,In_505);
nand U8081 (N_8081,In_2202,In_1468);
and U8082 (N_8082,In_2866,In_2670);
nand U8083 (N_8083,In_3139,In_2574);
xor U8084 (N_8084,In_3173,In_2453);
nor U8085 (N_8085,In_998,In_2855);
or U8086 (N_8086,In_4177,In_482);
nand U8087 (N_8087,In_4223,In_673);
or U8088 (N_8088,In_1869,In_3367);
or U8089 (N_8089,In_3618,In_451);
nand U8090 (N_8090,In_1458,In_1423);
or U8091 (N_8091,In_4792,In_4362);
or U8092 (N_8092,In_4663,In_3321);
or U8093 (N_8093,In_1085,In_2850);
or U8094 (N_8094,In_1598,In_1685);
or U8095 (N_8095,In_2557,In_2186);
nand U8096 (N_8096,In_1483,In_1060);
nor U8097 (N_8097,In_2166,In_99);
nor U8098 (N_8098,In_2749,In_3507);
and U8099 (N_8099,In_4160,In_3382);
or U8100 (N_8100,In_4512,In_3297);
or U8101 (N_8101,In_4807,In_228);
xnor U8102 (N_8102,In_2768,In_3668);
nand U8103 (N_8103,In_2729,In_1659);
nor U8104 (N_8104,In_1086,In_1115);
xor U8105 (N_8105,In_781,In_1443);
nor U8106 (N_8106,In_3530,In_4346);
and U8107 (N_8107,In_1988,In_3875);
xor U8108 (N_8108,In_4939,In_3945);
and U8109 (N_8109,In_429,In_669);
nor U8110 (N_8110,In_3479,In_927);
and U8111 (N_8111,In_4696,In_1283);
nor U8112 (N_8112,In_2020,In_2123);
and U8113 (N_8113,In_4536,In_4388);
and U8114 (N_8114,In_363,In_270);
xnor U8115 (N_8115,In_3232,In_4293);
nand U8116 (N_8116,In_1721,In_2403);
nand U8117 (N_8117,In_1179,In_537);
nor U8118 (N_8118,In_3825,In_2453);
nand U8119 (N_8119,In_3740,In_4608);
nand U8120 (N_8120,In_4041,In_2574);
xor U8121 (N_8121,In_2998,In_2973);
nand U8122 (N_8122,In_1883,In_4534);
nor U8123 (N_8123,In_3159,In_4511);
nand U8124 (N_8124,In_4014,In_4814);
and U8125 (N_8125,In_244,In_972);
nor U8126 (N_8126,In_2134,In_2111);
or U8127 (N_8127,In_1117,In_530);
nand U8128 (N_8128,In_1130,In_3003);
and U8129 (N_8129,In_2412,In_3141);
nand U8130 (N_8130,In_3037,In_799);
xnor U8131 (N_8131,In_1694,In_2122);
and U8132 (N_8132,In_2915,In_3448);
xor U8133 (N_8133,In_4042,In_1414);
nor U8134 (N_8134,In_2454,In_3625);
or U8135 (N_8135,In_4086,In_1289);
nand U8136 (N_8136,In_2566,In_2062);
and U8137 (N_8137,In_182,In_3083);
and U8138 (N_8138,In_2654,In_2994);
nor U8139 (N_8139,In_949,In_4460);
nand U8140 (N_8140,In_1612,In_4847);
xnor U8141 (N_8141,In_3195,In_2876);
and U8142 (N_8142,In_3456,In_4087);
and U8143 (N_8143,In_447,In_4428);
xnor U8144 (N_8144,In_2510,In_4577);
xor U8145 (N_8145,In_1137,In_4336);
and U8146 (N_8146,In_4387,In_3003);
xnor U8147 (N_8147,In_4519,In_3112);
xor U8148 (N_8148,In_4700,In_4551);
or U8149 (N_8149,In_2691,In_2950);
nand U8150 (N_8150,In_2161,In_4828);
xor U8151 (N_8151,In_273,In_4883);
nand U8152 (N_8152,In_2508,In_3187);
and U8153 (N_8153,In_167,In_215);
nor U8154 (N_8154,In_4731,In_2958);
xor U8155 (N_8155,In_3124,In_3407);
or U8156 (N_8156,In_848,In_3017);
nor U8157 (N_8157,In_2397,In_2157);
or U8158 (N_8158,In_2465,In_3095);
or U8159 (N_8159,In_1476,In_1178);
and U8160 (N_8160,In_4035,In_4832);
nor U8161 (N_8161,In_1250,In_1955);
nor U8162 (N_8162,In_1601,In_1620);
or U8163 (N_8163,In_2629,In_2122);
nand U8164 (N_8164,In_308,In_1747);
and U8165 (N_8165,In_3737,In_4878);
nand U8166 (N_8166,In_1,In_4993);
or U8167 (N_8167,In_1178,In_296);
nand U8168 (N_8168,In_3743,In_694);
and U8169 (N_8169,In_1725,In_4200);
and U8170 (N_8170,In_2039,In_4573);
or U8171 (N_8171,In_1233,In_2718);
and U8172 (N_8172,In_686,In_1811);
and U8173 (N_8173,In_4894,In_268);
or U8174 (N_8174,In_3552,In_3689);
or U8175 (N_8175,In_3013,In_3274);
nor U8176 (N_8176,In_1485,In_2292);
xnor U8177 (N_8177,In_130,In_3659);
nor U8178 (N_8178,In_2264,In_2248);
and U8179 (N_8179,In_1556,In_4808);
xnor U8180 (N_8180,In_2936,In_1436);
nand U8181 (N_8181,In_366,In_2659);
and U8182 (N_8182,In_4285,In_3788);
or U8183 (N_8183,In_1711,In_1494);
and U8184 (N_8184,In_3320,In_2446);
nor U8185 (N_8185,In_3267,In_2768);
or U8186 (N_8186,In_503,In_4758);
or U8187 (N_8187,In_3630,In_2557);
or U8188 (N_8188,In_1182,In_4986);
nand U8189 (N_8189,In_3203,In_2004);
and U8190 (N_8190,In_2243,In_1238);
xnor U8191 (N_8191,In_3191,In_4740);
nand U8192 (N_8192,In_3930,In_3789);
or U8193 (N_8193,In_721,In_3831);
or U8194 (N_8194,In_3508,In_4713);
nand U8195 (N_8195,In_3854,In_4879);
xnor U8196 (N_8196,In_4523,In_874);
or U8197 (N_8197,In_1837,In_4143);
nand U8198 (N_8198,In_4320,In_4090);
or U8199 (N_8199,In_3348,In_3478);
nand U8200 (N_8200,In_4689,In_4501);
nor U8201 (N_8201,In_2471,In_853);
xnor U8202 (N_8202,In_3566,In_2307);
nor U8203 (N_8203,In_4624,In_965);
or U8204 (N_8204,In_4933,In_4900);
or U8205 (N_8205,In_3903,In_379);
and U8206 (N_8206,In_2235,In_2150);
nand U8207 (N_8207,In_4510,In_170);
and U8208 (N_8208,In_1791,In_1477);
xnor U8209 (N_8209,In_1998,In_2738);
xnor U8210 (N_8210,In_649,In_978);
nor U8211 (N_8211,In_3557,In_3680);
nand U8212 (N_8212,In_2660,In_3804);
or U8213 (N_8213,In_2230,In_3996);
xnor U8214 (N_8214,In_4399,In_3374);
and U8215 (N_8215,In_4712,In_2406);
nand U8216 (N_8216,In_4999,In_1621);
nor U8217 (N_8217,In_734,In_882);
nand U8218 (N_8218,In_4970,In_3022);
or U8219 (N_8219,In_196,In_1672);
and U8220 (N_8220,In_938,In_3618);
and U8221 (N_8221,In_3985,In_138);
nand U8222 (N_8222,In_3718,In_2769);
nand U8223 (N_8223,In_620,In_3833);
nand U8224 (N_8224,In_4015,In_2350);
or U8225 (N_8225,In_3875,In_2334);
or U8226 (N_8226,In_3319,In_2531);
nand U8227 (N_8227,In_1533,In_1995);
and U8228 (N_8228,In_2540,In_1762);
nand U8229 (N_8229,In_4397,In_1336);
nor U8230 (N_8230,In_4645,In_2667);
xor U8231 (N_8231,In_4573,In_2643);
xor U8232 (N_8232,In_3925,In_825);
nor U8233 (N_8233,In_1563,In_1830);
nand U8234 (N_8234,In_3130,In_826);
nand U8235 (N_8235,In_681,In_1458);
and U8236 (N_8236,In_1548,In_3205);
nor U8237 (N_8237,In_867,In_1317);
nor U8238 (N_8238,In_108,In_1729);
xnor U8239 (N_8239,In_575,In_2661);
and U8240 (N_8240,In_1938,In_4568);
or U8241 (N_8241,In_1527,In_1788);
or U8242 (N_8242,In_1992,In_4295);
xnor U8243 (N_8243,In_1257,In_4518);
xor U8244 (N_8244,In_4056,In_3845);
nor U8245 (N_8245,In_4992,In_604);
or U8246 (N_8246,In_1403,In_1764);
nor U8247 (N_8247,In_4480,In_3330);
or U8248 (N_8248,In_3062,In_4623);
nor U8249 (N_8249,In_752,In_2323);
or U8250 (N_8250,In_789,In_2618);
nor U8251 (N_8251,In_1929,In_1808);
or U8252 (N_8252,In_733,In_3541);
and U8253 (N_8253,In_4499,In_1559);
nand U8254 (N_8254,In_2081,In_2355);
nand U8255 (N_8255,In_1412,In_531);
xnor U8256 (N_8256,In_496,In_3286);
xnor U8257 (N_8257,In_3062,In_3191);
nor U8258 (N_8258,In_2557,In_964);
nor U8259 (N_8259,In_1027,In_1483);
nand U8260 (N_8260,In_861,In_4933);
and U8261 (N_8261,In_1426,In_3657);
xnor U8262 (N_8262,In_1248,In_1030);
nor U8263 (N_8263,In_2684,In_2150);
and U8264 (N_8264,In_3828,In_3200);
nor U8265 (N_8265,In_3167,In_2852);
and U8266 (N_8266,In_425,In_1022);
or U8267 (N_8267,In_792,In_2009);
xor U8268 (N_8268,In_4538,In_664);
nand U8269 (N_8269,In_2012,In_2995);
or U8270 (N_8270,In_3351,In_2818);
or U8271 (N_8271,In_774,In_4146);
nand U8272 (N_8272,In_4152,In_994);
and U8273 (N_8273,In_1626,In_4761);
nor U8274 (N_8274,In_1719,In_1888);
and U8275 (N_8275,In_4903,In_2859);
or U8276 (N_8276,In_4295,In_1404);
nor U8277 (N_8277,In_1039,In_4620);
and U8278 (N_8278,In_611,In_3293);
nor U8279 (N_8279,In_1156,In_517);
xnor U8280 (N_8280,In_523,In_668);
nor U8281 (N_8281,In_3024,In_777);
xnor U8282 (N_8282,In_4143,In_3585);
or U8283 (N_8283,In_1892,In_156);
xnor U8284 (N_8284,In_499,In_3502);
nand U8285 (N_8285,In_4123,In_1779);
nor U8286 (N_8286,In_3152,In_4083);
nand U8287 (N_8287,In_1852,In_2799);
and U8288 (N_8288,In_4521,In_1096);
xor U8289 (N_8289,In_622,In_1675);
or U8290 (N_8290,In_4472,In_4510);
nor U8291 (N_8291,In_4072,In_3073);
and U8292 (N_8292,In_1615,In_3306);
xnor U8293 (N_8293,In_736,In_3200);
xnor U8294 (N_8294,In_1752,In_3545);
and U8295 (N_8295,In_1550,In_3378);
or U8296 (N_8296,In_3805,In_4269);
or U8297 (N_8297,In_3856,In_3313);
or U8298 (N_8298,In_3647,In_3393);
nor U8299 (N_8299,In_3313,In_2056);
or U8300 (N_8300,In_3601,In_4328);
and U8301 (N_8301,In_481,In_3646);
xnor U8302 (N_8302,In_1593,In_2976);
nor U8303 (N_8303,In_3167,In_1598);
or U8304 (N_8304,In_1868,In_3381);
xnor U8305 (N_8305,In_3522,In_1005);
xor U8306 (N_8306,In_2830,In_3268);
or U8307 (N_8307,In_2609,In_3663);
or U8308 (N_8308,In_3505,In_3880);
and U8309 (N_8309,In_2558,In_316);
nor U8310 (N_8310,In_3416,In_4321);
nor U8311 (N_8311,In_3252,In_4878);
nand U8312 (N_8312,In_2021,In_2924);
or U8313 (N_8313,In_3326,In_3430);
nand U8314 (N_8314,In_4328,In_3218);
or U8315 (N_8315,In_473,In_3142);
or U8316 (N_8316,In_4749,In_2373);
and U8317 (N_8317,In_4461,In_2052);
nand U8318 (N_8318,In_1766,In_2564);
or U8319 (N_8319,In_2711,In_2089);
xnor U8320 (N_8320,In_2580,In_2164);
xnor U8321 (N_8321,In_459,In_2548);
xnor U8322 (N_8322,In_170,In_743);
or U8323 (N_8323,In_4863,In_963);
and U8324 (N_8324,In_1790,In_4073);
xor U8325 (N_8325,In_2836,In_3038);
nand U8326 (N_8326,In_1440,In_3474);
or U8327 (N_8327,In_110,In_1750);
nand U8328 (N_8328,In_2413,In_822);
nor U8329 (N_8329,In_888,In_1340);
or U8330 (N_8330,In_2608,In_3546);
nor U8331 (N_8331,In_1908,In_368);
nor U8332 (N_8332,In_1807,In_2966);
xnor U8333 (N_8333,In_179,In_4737);
and U8334 (N_8334,In_233,In_3780);
and U8335 (N_8335,In_3213,In_987);
nand U8336 (N_8336,In_4895,In_1611);
nor U8337 (N_8337,In_861,In_2445);
nor U8338 (N_8338,In_3693,In_3743);
xor U8339 (N_8339,In_4393,In_2878);
or U8340 (N_8340,In_2140,In_2833);
nand U8341 (N_8341,In_4920,In_3612);
nand U8342 (N_8342,In_23,In_3410);
or U8343 (N_8343,In_3072,In_3049);
and U8344 (N_8344,In_4192,In_3652);
nor U8345 (N_8345,In_127,In_2577);
or U8346 (N_8346,In_4630,In_2604);
nor U8347 (N_8347,In_3329,In_2238);
nor U8348 (N_8348,In_1258,In_3088);
xnor U8349 (N_8349,In_4592,In_3114);
nand U8350 (N_8350,In_2524,In_3323);
and U8351 (N_8351,In_2747,In_975);
nor U8352 (N_8352,In_1350,In_604);
xor U8353 (N_8353,In_794,In_315);
nand U8354 (N_8354,In_406,In_3837);
or U8355 (N_8355,In_4388,In_4532);
nor U8356 (N_8356,In_2647,In_1032);
nand U8357 (N_8357,In_4865,In_2387);
nor U8358 (N_8358,In_3052,In_3147);
nor U8359 (N_8359,In_254,In_4140);
nand U8360 (N_8360,In_2764,In_4994);
or U8361 (N_8361,In_2298,In_2833);
or U8362 (N_8362,In_2057,In_3553);
nand U8363 (N_8363,In_578,In_4718);
or U8364 (N_8364,In_717,In_1428);
or U8365 (N_8365,In_1863,In_4743);
or U8366 (N_8366,In_1037,In_220);
xor U8367 (N_8367,In_4800,In_3633);
xnor U8368 (N_8368,In_4372,In_3965);
and U8369 (N_8369,In_1877,In_2557);
xnor U8370 (N_8370,In_3841,In_2896);
nor U8371 (N_8371,In_3629,In_1670);
or U8372 (N_8372,In_1987,In_3690);
or U8373 (N_8373,In_3675,In_1214);
or U8374 (N_8374,In_2665,In_3669);
or U8375 (N_8375,In_4715,In_4996);
nor U8376 (N_8376,In_4728,In_3628);
and U8377 (N_8377,In_4366,In_377);
nand U8378 (N_8378,In_1966,In_3029);
or U8379 (N_8379,In_431,In_3593);
nand U8380 (N_8380,In_2720,In_2632);
xor U8381 (N_8381,In_3200,In_3125);
xor U8382 (N_8382,In_1358,In_43);
xnor U8383 (N_8383,In_648,In_3074);
and U8384 (N_8384,In_2108,In_3014);
xor U8385 (N_8385,In_2564,In_68);
nor U8386 (N_8386,In_2988,In_1436);
or U8387 (N_8387,In_4334,In_774);
nand U8388 (N_8388,In_3198,In_4440);
and U8389 (N_8389,In_1798,In_2348);
nand U8390 (N_8390,In_171,In_3521);
and U8391 (N_8391,In_4688,In_3819);
or U8392 (N_8392,In_900,In_3861);
xnor U8393 (N_8393,In_4757,In_1790);
or U8394 (N_8394,In_2885,In_355);
xnor U8395 (N_8395,In_2584,In_3864);
xnor U8396 (N_8396,In_1144,In_1506);
nor U8397 (N_8397,In_2860,In_2884);
nor U8398 (N_8398,In_4762,In_3621);
or U8399 (N_8399,In_1342,In_3760);
nor U8400 (N_8400,In_2792,In_690);
xnor U8401 (N_8401,In_912,In_3315);
and U8402 (N_8402,In_399,In_3403);
xor U8403 (N_8403,In_2246,In_2470);
or U8404 (N_8404,In_4856,In_1995);
nor U8405 (N_8405,In_4204,In_4002);
xor U8406 (N_8406,In_2776,In_1423);
xnor U8407 (N_8407,In_3283,In_4013);
nand U8408 (N_8408,In_537,In_4968);
nor U8409 (N_8409,In_3183,In_80);
nand U8410 (N_8410,In_72,In_4617);
nand U8411 (N_8411,In_2813,In_200);
nand U8412 (N_8412,In_2375,In_718);
xnor U8413 (N_8413,In_2096,In_3401);
nor U8414 (N_8414,In_1130,In_665);
or U8415 (N_8415,In_377,In_1250);
and U8416 (N_8416,In_2426,In_3616);
nand U8417 (N_8417,In_4319,In_252);
or U8418 (N_8418,In_2801,In_1783);
nor U8419 (N_8419,In_1048,In_1920);
and U8420 (N_8420,In_1448,In_4609);
and U8421 (N_8421,In_1548,In_2324);
nand U8422 (N_8422,In_4167,In_1286);
nor U8423 (N_8423,In_4107,In_3517);
nor U8424 (N_8424,In_2426,In_1560);
or U8425 (N_8425,In_3464,In_3828);
nor U8426 (N_8426,In_4419,In_668);
nand U8427 (N_8427,In_4661,In_3897);
and U8428 (N_8428,In_1516,In_501);
and U8429 (N_8429,In_3033,In_2820);
and U8430 (N_8430,In_4274,In_3263);
and U8431 (N_8431,In_4701,In_4847);
nand U8432 (N_8432,In_841,In_4260);
and U8433 (N_8433,In_1635,In_323);
nor U8434 (N_8434,In_4324,In_1502);
or U8435 (N_8435,In_3377,In_3538);
nand U8436 (N_8436,In_4862,In_4363);
nand U8437 (N_8437,In_2852,In_4206);
or U8438 (N_8438,In_2124,In_1413);
nand U8439 (N_8439,In_4527,In_1783);
xnor U8440 (N_8440,In_1813,In_2299);
and U8441 (N_8441,In_1988,In_3492);
xor U8442 (N_8442,In_1810,In_4184);
nand U8443 (N_8443,In_1005,In_3989);
and U8444 (N_8444,In_3693,In_4285);
xnor U8445 (N_8445,In_4556,In_2932);
or U8446 (N_8446,In_4427,In_3737);
nor U8447 (N_8447,In_1683,In_2352);
nand U8448 (N_8448,In_3498,In_4814);
nand U8449 (N_8449,In_4825,In_2415);
nand U8450 (N_8450,In_417,In_3920);
or U8451 (N_8451,In_2320,In_1506);
and U8452 (N_8452,In_3082,In_1593);
or U8453 (N_8453,In_3826,In_3698);
or U8454 (N_8454,In_4993,In_4499);
nor U8455 (N_8455,In_4880,In_2942);
and U8456 (N_8456,In_4349,In_1967);
xor U8457 (N_8457,In_440,In_821);
or U8458 (N_8458,In_3549,In_4229);
and U8459 (N_8459,In_3547,In_2709);
and U8460 (N_8460,In_2419,In_4550);
or U8461 (N_8461,In_1422,In_1528);
nand U8462 (N_8462,In_4386,In_2684);
nor U8463 (N_8463,In_1149,In_4750);
or U8464 (N_8464,In_2580,In_456);
and U8465 (N_8465,In_4793,In_2437);
or U8466 (N_8466,In_2460,In_2846);
or U8467 (N_8467,In_3291,In_4776);
xnor U8468 (N_8468,In_161,In_454);
nand U8469 (N_8469,In_2978,In_2564);
or U8470 (N_8470,In_2078,In_2976);
nor U8471 (N_8471,In_3832,In_4978);
nand U8472 (N_8472,In_2913,In_1434);
or U8473 (N_8473,In_4165,In_1917);
xnor U8474 (N_8474,In_3282,In_3302);
nor U8475 (N_8475,In_3649,In_3468);
xor U8476 (N_8476,In_894,In_2006);
xor U8477 (N_8477,In_3620,In_814);
nor U8478 (N_8478,In_899,In_2754);
or U8479 (N_8479,In_2339,In_3365);
or U8480 (N_8480,In_2948,In_1168);
xor U8481 (N_8481,In_462,In_889);
nor U8482 (N_8482,In_3568,In_1224);
nor U8483 (N_8483,In_1473,In_631);
and U8484 (N_8484,In_1752,In_3394);
xnor U8485 (N_8485,In_1400,In_4595);
nand U8486 (N_8486,In_3363,In_3062);
xnor U8487 (N_8487,In_4865,In_2085);
xnor U8488 (N_8488,In_3068,In_860);
nand U8489 (N_8489,In_4286,In_1216);
or U8490 (N_8490,In_3419,In_438);
xnor U8491 (N_8491,In_4115,In_1908);
and U8492 (N_8492,In_2083,In_4488);
nor U8493 (N_8493,In_3651,In_624);
nor U8494 (N_8494,In_1385,In_1045);
nand U8495 (N_8495,In_3135,In_3681);
and U8496 (N_8496,In_3615,In_3929);
nand U8497 (N_8497,In_3791,In_3277);
xnor U8498 (N_8498,In_3679,In_3182);
nand U8499 (N_8499,In_750,In_3665);
and U8500 (N_8500,In_927,In_1504);
xor U8501 (N_8501,In_1626,In_1762);
nand U8502 (N_8502,In_1701,In_3535);
nand U8503 (N_8503,In_1087,In_3794);
xor U8504 (N_8504,In_2104,In_2734);
or U8505 (N_8505,In_624,In_2545);
or U8506 (N_8506,In_1111,In_1597);
nor U8507 (N_8507,In_422,In_2109);
or U8508 (N_8508,In_3861,In_1070);
and U8509 (N_8509,In_4708,In_803);
and U8510 (N_8510,In_2081,In_1980);
nor U8511 (N_8511,In_2695,In_207);
nor U8512 (N_8512,In_4522,In_2134);
and U8513 (N_8513,In_4555,In_1566);
nand U8514 (N_8514,In_2878,In_4514);
nor U8515 (N_8515,In_158,In_2563);
and U8516 (N_8516,In_4584,In_1486);
nand U8517 (N_8517,In_1145,In_3803);
xnor U8518 (N_8518,In_3552,In_4505);
nor U8519 (N_8519,In_3364,In_1405);
and U8520 (N_8520,In_1348,In_575);
nor U8521 (N_8521,In_1677,In_1974);
xor U8522 (N_8522,In_3014,In_4323);
nand U8523 (N_8523,In_2776,In_4418);
nand U8524 (N_8524,In_4526,In_4502);
nor U8525 (N_8525,In_4714,In_1049);
or U8526 (N_8526,In_4109,In_2570);
xnor U8527 (N_8527,In_2732,In_510);
and U8528 (N_8528,In_3071,In_4391);
or U8529 (N_8529,In_4803,In_383);
nor U8530 (N_8530,In_2410,In_1980);
xnor U8531 (N_8531,In_3928,In_3948);
xnor U8532 (N_8532,In_2296,In_627);
xnor U8533 (N_8533,In_409,In_749);
nand U8534 (N_8534,In_1390,In_2652);
and U8535 (N_8535,In_3405,In_1113);
nand U8536 (N_8536,In_1909,In_2507);
nand U8537 (N_8537,In_286,In_27);
nand U8538 (N_8538,In_1344,In_1436);
nor U8539 (N_8539,In_1102,In_4771);
and U8540 (N_8540,In_34,In_3016);
and U8541 (N_8541,In_3362,In_2425);
xnor U8542 (N_8542,In_1852,In_1633);
nor U8543 (N_8543,In_4953,In_2518);
nand U8544 (N_8544,In_1112,In_3387);
nand U8545 (N_8545,In_4852,In_2955);
nor U8546 (N_8546,In_2519,In_3433);
and U8547 (N_8547,In_4117,In_4600);
or U8548 (N_8548,In_4800,In_4311);
and U8549 (N_8549,In_3575,In_2970);
and U8550 (N_8550,In_4494,In_2416);
xor U8551 (N_8551,In_3239,In_4862);
nand U8552 (N_8552,In_4670,In_4324);
nand U8553 (N_8553,In_1853,In_3923);
or U8554 (N_8554,In_790,In_157);
nor U8555 (N_8555,In_459,In_762);
xnor U8556 (N_8556,In_4055,In_3732);
xor U8557 (N_8557,In_3842,In_2524);
nand U8558 (N_8558,In_1588,In_4568);
nand U8559 (N_8559,In_2804,In_2077);
and U8560 (N_8560,In_4842,In_3884);
xor U8561 (N_8561,In_2007,In_2850);
or U8562 (N_8562,In_3401,In_821);
xor U8563 (N_8563,In_1823,In_1098);
nand U8564 (N_8564,In_68,In_4459);
or U8565 (N_8565,In_1265,In_2139);
nand U8566 (N_8566,In_1223,In_1787);
and U8567 (N_8567,In_4685,In_4876);
nor U8568 (N_8568,In_3380,In_3457);
nand U8569 (N_8569,In_2538,In_4321);
and U8570 (N_8570,In_414,In_1023);
or U8571 (N_8571,In_3818,In_1322);
xor U8572 (N_8572,In_2242,In_2863);
nand U8573 (N_8573,In_4477,In_2576);
and U8574 (N_8574,In_483,In_4030);
and U8575 (N_8575,In_2251,In_955);
or U8576 (N_8576,In_2592,In_4648);
nand U8577 (N_8577,In_2782,In_4445);
or U8578 (N_8578,In_1007,In_4047);
and U8579 (N_8579,In_4744,In_255);
xnor U8580 (N_8580,In_4698,In_325);
xnor U8581 (N_8581,In_2774,In_2505);
or U8582 (N_8582,In_922,In_4242);
and U8583 (N_8583,In_941,In_546);
nor U8584 (N_8584,In_3412,In_3141);
nor U8585 (N_8585,In_435,In_2909);
nor U8586 (N_8586,In_4936,In_1178);
nor U8587 (N_8587,In_2111,In_2804);
or U8588 (N_8588,In_1705,In_3972);
nor U8589 (N_8589,In_1835,In_2747);
nor U8590 (N_8590,In_4016,In_1476);
or U8591 (N_8591,In_2513,In_4678);
and U8592 (N_8592,In_1849,In_2477);
or U8593 (N_8593,In_542,In_2857);
xor U8594 (N_8594,In_2937,In_4930);
xnor U8595 (N_8595,In_3787,In_518);
nand U8596 (N_8596,In_2155,In_3935);
xnor U8597 (N_8597,In_1276,In_3154);
or U8598 (N_8598,In_604,In_2045);
nand U8599 (N_8599,In_2726,In_3271);
xor U8600 (N_8600,In_1862,In_1240);
nand U8601 (N_8601,In_495,In_589);
or U8602 (N_8602,In_2275,In_3543);
or U8603 (N_8603,In_1268,In_4570);
nor U8604 (N_8604,In_312,In_1226);
or U8605 (N_8605,In_2923,In_4086);
xor U8606 (N_8606,In_275,In_3901);
xnor U8607 (N_8607,In_3186,In_2524);
nand U8608 (N_8608,In_793,In_4615);
or U8609 (N_8609,In_50,In_1272);
and U8610 (N_8610,In_1995,In_2414);
or U8611 (N_8611,In_863,In_780);
or U8612 (N_8612,In_31,In_3724);
nand U8613 (N_8613,In_2533,In_3908);
nand U8614 (N_8614,In_191,In_1687);
nor U8615 (N_8615,In_3675,In_3176);
nor U8616 (N_8616,In_3712,In_1938);
nor U8617 (N_8617,In_3561,In_2364);
xor U8618 (N_8618,In_4834,In_1699);
nor U8619 (N_8619,In_4595,In_784);
xor U8620 (N_8620,In_1107,In_436);
or U8621 (N_8621,In_4517,In_3666);
and U8622 (N_8622,In_571,In_3179);
or U8623 (N_8623,In_144,In_1940);
nand U8624 (N_8624,In_3195,In_1231);
nand U8625 (N_8625,In_1760,In_4258);
nor U8626 (N_8626,In_1537,In_956);
nor U8627 (N_8627,In_4870,In_4770);
or U8628 (N_8628,In_1613,In_1332);
nand U8629 (N_8629,In_4841,In_3431);
xnor U8630 (N_8630,In_3905,In_2511);
xor U8631 (N_8631,In_19,In_3332);
nor U8632 (N_8632,In_4026,In_4157);
and U8633 (N_8633,In_262,In_1900);
xor U8634 (N_8634,In_1189,In_2888);
or U8635 (N_8635,In_995,In_540);
or U8636 (N_8636,In_4556,In_4038);
and U8637 (N_8637,In_126,In_2031);
xnor U8638 (N_8638,In_992,In_3887);
and U8639 (N_8639,In_1871,In_3613);
xor U8640 (N_8640,In_862,In_4688);
nand U8641 (N_8641,In_1590,In_1307);
nor U8642 (N_8642,In_844,In_863);
and U8643 (N_8643,In_930,In_2779);
nand U8644 (N_8644,In_413,In_4314);
or U8645 (N_8645,In_3133,In_2050);
nor U8646 (N_8646,In_3863,In_2140);
or U8647 (N_8647,In_4663,In_141);
xnor U8648 (N_8648,In_4209,In_3554);
or U8649 (N_8649,In_2044,In_3561);
or U8650 (N_8650,In_2260,In_4712);
and U8651 (N_8651,In_3673,In_1845);
and U8652 (N_8652,In_1521,In_305);
or U8653 (N_8653,In_4135,In_4639);
and U8654 (N_8654,In_3649,In_293);
and U8655 (N_8655,In_1855,In_2839);
or U8656 (N_8656,In_1535,In_3010);
nor U8657 (N_8657,In_4129,In_3253);
nand U8658 (N_8658,In_2839,In_374);
and U8659 (N_8659,In_3625,In_1216);
nor U8660 (N_8660,In_4548,In_2929);
nand U8661 (N_8661,In_4715,In_2827);
and U8662 (N_8662,In_2785,In_1186);
nor U8663 (N_8663,In_2332,In_3362);
nand U8664 (N_8664,In_1401,In_1514);
or U8665 (N_8665,In_4707,In_2080);
xnor U8666 (N_8666,In_521,In_3826);
nor U8667 (N_8667,In_4598,In_4452);
and U8668 (N_8668,In_3993,In_996);
and U8669 (N_8669,In_273,In_108);
nor U8670 (N_8670,In_3300,In_310);
and U8671 (N_8671,In_1207,In_4443);
nand U8672 (N_8672,In_4346,In_1285);
nor U8673 (N_8673,In_353,In_1429);
xor U8674 (N_8674,In_3502,In_2163);
and U8675 (N_8675,In_4064,In_3770);
nand U8676 (N_8676,In_477,In_1441);
nand U8677 (N_8677,In_1227,In_150);
and U8678 (N_8678,In_3375,In_112);
and U8679 (N_8679,In_4565,In_433);
and U8680 (N_8680,In_2139,In_4031);
nor U8681 (N_8681,In_576,In_2538);
and U8682 (N_8682,In_3730,In_1720);
or U8683 (N_8683,In_2284,In_3124);
and U8684 (N_8684,In_1805,In_2445);
nor U8685 (N_8685,In_873,In_1788);
or U8686 (N_8686,In_3450,In_4906);
and U8687 (N_8687,In_2611,In_1684);
nand U8688 (N_8688,In_1015,In_4045);
nand U8689 (N_8689,In_1136,In_536);
and U8690 (N_8690,In_3871,In_3763);
nand U8691 (N_8691,In_3395,In_4941);
xor U8692 (N_8692,In_2280,In_3334);
or U8693 (N_8693,In_1631,In_2307);
xnor U8694 (N_8694,In_2775,In_4777);
xnor U8695 (N_8695,In_2348,In_2623);
and U8696 (N_8696,In_2918,In_3495);
or U8697 (N_8697,In_3041,In_4606);
xnor U8698 (N_8698,In_3998,In_4147);
and U8699 (N_8699,In_1577,In_3042);
xor U8700 (N_8700,In_4427,In_2634);
nor U8701 (N_8701,In_4990,In_3308);
and U8702 (N_8702,In_313,In_4982);
and U8703 (N_8703,In_333,In_1246);
nand U8704 (N_8704,In_3276,In_2059);
xor U8705 (N_8705,In_2841,In_2487);
nor U8706 (N_8706,In_3387,In_2554);
xor U8707 (N_8707,In_3875,In_297);
and U8708 (N_8708,In_2169,In_4302);
nand U8709 (N_8709,In_670,In_3005);
nor U8710 (N_8710,In_4711,In_4703);
nor U8711 (N_8711,In_2331,In_975);
nand U8712 (N_8712,In_1163,In_4589);
nand U8713 (N_8713,In_1302,In_2963);
and U8714 (N_8714,In_204,In_2112);
and U8715 (N_8715,In_1777,In_3314);
nand U8716 (N_8716,In_4259,In_4371);
xor U8717 (N_8717,In_2749,In_4920);
or U8718 (N_8718,In_554,In_354);
or U8719 (N_8719,In_2861,In_1555);
nand U8720 (N_8720,In_4695,In_1178);
nand U8721 (N_8721,In_763,In_983);
xor U8722 (N_8722,In_540,In_2782);
and U8723 (N_8723,In_2769,In_2860);
or U8724 (N_8724,In_847,In_629);
nor U8725 (N_8725,In_4324,In_3761);
and U8726 (N_8726,In_15,In_1122);
nor U8727 (N_8727,In_4438,In_2356);
nor U8728 (N_8728,In_1387,In_164);
and U8729 (N_8729,In_425,In_3997);
nand U8730 (N_8730,In_4505,In_4312);
nor U8731 (N_8731,In_4736,In_2645);
xnor U8732 (N_8732,In_464,In_3701);
xor U8733 (N_8733,In_2988,In_718);
xnor U8734 (N_8734,In_2342,In_4413);
xor U8735 (N_8735,In_1541,In_1340);
nor U8736 (N_8736,In_2566,In_3951);
xnor U8737 (N_8737,In_2477,In_4434);
and U8738 (N_8738,In_3127,In_483);
or U8739 (N_8739,In_1935,In_328);
or U8740 (N_8740,In_855,In_1032);
nor U8741 (N_8741,In_193,In_4255);
nor U8742 (N_8742,In_662,In_887);
and U8743 (N_8743,In_2760,In_2439);
or U8744 (N_8744,In_3220,In_3744);
nand U8745 (N_8745,In_2596,In_797);
nor U8746 (N_8746,In_1166,In_3793);
or U8747 (N_8747,In_1313,In_215);
or U8748 (N_8748,In_1230,In_395);
and U8749 (N_8749,In_1854,In_617);
nand U8750 (N_8750,In_4509,In_4032);
nand U8751 (N_8751,In_4234,In_2541);
xnor U8752 (N_8752,In_774,In_1007);
nor U8753 (N_8753,In_1462,In_1223);
or U8754 (N_8754,In_965,In_3542);
and U8755 (N_8755,In_4276,In_3126);
or U8756 (N_8756,In_1228,In_1025);
nand U8757 (N_8757,In_360,In_2162);
nand U8758 (N_8758,In_66,In_2026);
xnor U8759 (N_8759,In_241,In_2920);
or U8760 (N_8760,In_426,In_844);
nand U8761 (N_8761,In_3824,In_3988);
nor U8762 (N_8762,In_1717,In_4953);
nor U8763 (N_8763,In_1843,In_813);
or U8764 (N_8764,In_4182,In_2842);
and U8765 (N_8765,In_121,In_292);
nor U8766 (N_8766,In_4335,In_2692);
and U8767 (N_8767,In_2179,In_4669);
xnor U8768 (N_8768,In_1558,In_2268);
xnor U8769 (N_8769,In_1453,In_3980);
or U8770 (N_8770,In_2545,In_4800);
nand U8771 (N_8771,In_350,In_4236);
or U8772 (N_8772,In_4095,In_1237);
or U8773 (N_8773,In_4946,In_2663);
or U8774 (N_8774,In_2418,In_134);
or U8775 (N_8775,In_3708,In_2796);
or U8776 (N_8776,In_148,In_3495);
xnor U8777 (N_8777,In_2233,In_3195);
xnor U8778 (N_8778,In_3339,In_1283);
xor U8779 (N_8779,In_2507,In_3255);
xnor U8780 (N_8780,In_181,In_4529);
xnor U8781 (N_8781,In_259,In_1998);
xor U8782 (N_8782,In_3006,In_3513);
nand U8783 (N_8783,In_1430,In_4577);
and U8784 (N_8784,In_3160,In_4511);
nand U8785 (N_8785,In_3190,In_2224);
or U8786 (N_8786,In_379,In_1926);
nor U8787 (N_8787,In_2290,In_996);
nand U8788 (N_8788,In_3349,In_172);
nand U8789 (N_8789,In_2042,In_2935);
xor U8790 (N_8790,In_1918,In_335);
or U8791 (N_8791,In_499,In_1048);
xor U8792 (N_8792,In_574,In_2651);
and U8793 (N_8793,In_2180,In_2334);
nand U8794 (N_8794,In_3144,In_1189);
nand U8795 (N_8795,In_2081,In_927);
and U8796 (N_8796,In_2418,In_2749);
xor U8797 (N_8797,In_1784,In_1788);
xor U8798 (N_8798,In_4424,In_4016);
and U8799 (N_8799,In_2457,In_749);
xnor U8800 (N_8800,In_3129,In_1669);
xnor U8801 (N_8801,In_4030,In_4432);
nor U8802 (N_8802,In_712,In_4670);
nand U8803 (N_8803,In_2144,In_3791);
and U8804 (N_8804,In_237,In_2049);
and U8805 (N_8805,In_4235,In_4755);
xnor U8806 (N_8806,In_215,In_65);
nor U8807 (N_8807,In_3202,In_2906);
nor U8808 (N_8808,In_4322,In_2984);
nand U8809 (N_8809,In_2708,In_1099);
and U8810 (N_8810,In_792,In_3253);
and U8811 (N_8811,In_2611,In_4299);
xor U8812 (N_8812,In_3466,In_2952);
nand U8813 (N_8813,In_3105,In_2849);
xor U8814 (N_8814,In_2926,In_4123);
xnor U8815 (N_8815,In_4347,In_402);
and U8816 (N_8816,In_407,In_1165);
nand U8817 (N_8817,In_3589,In_1266);
nand U8818 (N_8818,In_2065,In_4128);
xor U8819 (N_8819,In_3084,In_788);
nor U8820 (N_8820,In_980,In_899);
xnor U8821 (N_8821,In_2855,In_693);
nand U8822 (N_8822,In_1284,In_311);
xor U8823 (N_8823,In_124,In_165);
and U8824 (N_8824,In_31,In_999);
nand U8825 (N_8825,In_1530,In_1128);
and U8826 (N_8826,In_552,In_4677);
or U8827 (N_8827,In_2725,In_4276);
or U8828 (N_8828,In_3876,In_160);
nand U8829 (N_8829,In_3134,In_3401);
and U8830 (N_8830,In_1003,In_4660);
nand U8831 (N_8831,In_4776,In_2528);
and U8832 (N_8832,In_4582,In_2809);
nand U8833 (N_8833,In_2869,In_410);
nor U8834 (N_8834,In_1009,In_169);
nand U8835 (N_8835,In_607,In_2385);
nor U8836 (N_8836,In_4108,In_3307);
nand U8837 (N_8837,In_1795,In_4474);
xor U8838 (N_8838,In_663,In_645);
nand U8839 (N_8839,In_4394,In_2193);
xnor U8840 (N_8840,In_1551,In_2474);
or U8841 (N_8841,In_680,In_3953);
or U8842 (N_8842,In_1152,In_2779);
nand U8843 (N_8843,In_783,In_863);
nor U8844 (N_8844,In_644,In_455);
and U8845 (N_8845,In_4757,In_3139);
nor U8846 (N_8846,In_2287,In_3833);
or U8847 (N_8847,In_3301,In_326);
nor U8848 (N_8848,In_1070,In_1435);
nand U8849 (N_8849,In_4426,In_2816);
and U8850 (N_8850,In_4108,In_3432);
xnor U8851 (N_8851,In_857,In_4825);
and U8852 (N_8852,In_3023,In_3989);
xor U8853 (N_8853,In_133,In_3688);
or U8854 (N_8854,In_2032,In_2680);
nand U8855 (N_8855,In_1575,In_1154);
nor U8856 (N_8856,In_974,In_3313);
nand U8857 (N_8857,In_1259,In_2764);
nand U8858 (N_8858,In_330,In_4418);
nand U8859 (N_8859,In_153,In_190);
nand U8860 (N_8860,In_933,In_1340);
xor U8861 (N_8861,In_1596,In_3148);
and U8862 (N_8862,In_3968,In_208);
or U8863 (N_8863,In_3524,In_1825);
or U8864 (N_8864,In_2918,In_820);
nand U8865 (N_8865,In_3989,In_4683);
and U8866 (N_8866,In_4856,In_1944);
and U8867 (N_8867,In_315,In_1526);
or U8868 (N_8868,In_1865,In_68);
and U8869 (N_8869,In_1329,In_860);
nor U8870 (N_8870,In_1713,In_2805);
xor U8871 (N_8871,In_4971,In_3684);
and U8872 (N_8872,In_114,In_204);
nand U8873 (N_8873,In_2559,In_2721);
xnor U8874 (N_8874,In_2410,In_2702);
or U8875 (N_8875,In_3062,In_2203);
and U8876 (N_8876,In_1139,In_1027);
nor U8877 (N_8877,In_2944,In_3381);
and U8878 (N_8878,In_2839,In_3607);
nor U8879 (N_8879,In_3113,In_3585);
nor U8880 (N_8880,In_4000,In_546);
or U8881 (N_8881,In_2583,In_845);
or U8882 (N_8882,In_4273,In_4646);
nor U8883 (N_8883,In_2343,In_2546);
nand U8884 (N_8884,In_1087,In_1444);
nor U8885 (N_8885,In_3287,In_1306);
and U8886 (N_8886,In_1113,In_252);
xor U8887 (N_8887,In_4207,In_4327);
and U8888 (N_8888,In_564,In_2281);
or U8889 (N_8889,In_4736,In_4619);
xnor U8890 (N_8890,In_2690,In_3136);
nor U8891 (N_8891,In_3957,In_3848);
nand U8892 (N_8892,In_4644,In_201);
or U8893 (N_8893,In_2248,In_1917);
or U8894 (N_8894,In_1532,In_1755);
and U8895 (N_8895,In_2328,In_4076);
nand U8896 (N_8896,In_2490,In_2234);
xnor U8897 (N_8897,In_4323,In_2834);
nor U8898 (N_8898,In_2926,In_2802);
or U8899 (N_8899,In_2253,In_4795);
xnor U8900 (N_8900,In_39,In_1559);
and U8901 (N_8901,In_3807,In_1943);
or U8902 (N_8902,In_4584,In_2537);
nand U8903 (N_8903,In_2477,In_3372);
nand U8904 (N_8904,In_2345,In_3770);
xor U8905 (N_8905,In_2237,In_3084);
or U8906 (N_8906,In_3203,In_4043);
xnor U8907 (N_8907,In_1132,In_198);
and U8908 (N_8908,In_1765,In_3523);
and U8909 (N_8909,In_862,In_4212);
and U8910 (N_8910,In_2802,In_3926);
or U8911 (N_8911,In_2368,In_3910);
or U8912 (N_8912,In_2409,In_3484);
nor U8913 (N_8913,In_769,In_3724);
and U8914 (N_8914,In_965,In_2654);
and U8915 (N_8915,In_2765,In_685);
or U8916 (N_8916,In_274,In_4365);
nor U8917 (N_8917,In_3373,In_262);
xor U8918 (N_8918,In_2218,In_4381);
nand U8919 (N_8919,In_2278,In_1556);
and U8920 (N_8920,In_2428,In_1795);
or U8921 (N_8921,In_2008,In_997);
xor U8922 (N_8922,In_4755,In_369);
nor U8923 (N_8923,In_2762,In_4252);
nand U8924 (N_8924,In_1596,In_3861);
and U8925 (N_8925,In_872,In_976);
and U8926 (N_8926,In_3233,In_1468);
and U8927 (N_8927,In_2243,In_1107);
and U8928 (N_8928,In_1572,In_1418);
nor U8929 (N_8929,In_4470,In_456);
xnor U8930 (N_8930,In_2476,In_284);
nand U8931 (N_8931,In_4261,In_4135);
or U8932 (N_8932,In_1881,In_2128);
nor U8933 (N_8933,In_1153,In_387);
nand U8934 (N_8934,In_1412,In_1344);
nor U8935 (N_8935,In_2929,In_1558);
xor U8936 (N_8936,In_133,In_4053);
and U8937 (N_8937,In_4906,In_3417);
nand U8938 (N_8938,In_869,In_1074);
xnor U8939 (N_8939,In_2832,In_2783);
nand U8940 (N_8940,In_2543,In_2899);
nand U8941 (N_8941,In_718,In_2703);
or U8942 (N_8942,In_2578,In_1205);
nand U8943 (N_8943,In_4419,In_4055);
and U8944 (N_8944,In_3855,In_3856);
and U8945 (N_8945,In_3380,In_913);
or U8946 (N_8946,In_4722,In_2841);
nor U8947 (N_8947,In_2946,In_3859);
and U8948 (N_8948,In_4686,In_3755);
nand U8949 (N_8949,In_2961,In_3782);
nor U8950 (N_8950,In_3016,In_292);
xnor U8951 (N_8951,In_1326,In_887);
and U8952 (N_8952,In_4986,In_1535);
and U8953 (N_8953,In_3317,In_4879);
or U8954 (N_8954,In_2025,In_3125);
or U8955 (N_8955,In_4816,In_1017);
xor U8956 (N_8956,In_3334,In_4054);
nand U8957 (N_8957,In_2999,In_3503);
xor U8958 (N_8958,In_1791,In_27);
nand U8959 (N_8959,In_4015,In_3685);
nand U8960 (N_8960,In_1674,In_1355);
and U8961 (N_8961,In_1037,In_927);
nor U8962 (N_8962,In_3448,In_6);
nand U8963 (N_8963,In_3925,In_375);
xor U8964 (N_8964,In_3416,In_215);
nor U8965 (N_8965,In_817,In_4559);
xor U8966 (N_8966,In_216,In_4418);
nor U8967 (N_8967,In_943,In_3793);
and U8968 (N_8968,In_4429,In_3338);
nor U8969 (N_8969,In_3160,In_3135);
nor U8970 (N_8970,In_387,In_1087);
and U8971 (N_8971,In_456,In_4725);
nand U8972 (N_8972,In_592,In_2118);
xor U8973 (N_8973,In_1560,In_1202);
and U8974 (N_8974,In_1078,In_735);
or U8975 (N_8975,In_1589,In_4995);
xor U8976 (N_8976,In_414,In_4533);
and U8977 (N_8977,In_133,In_2847);
xor U8978 (N_8978,In_1121,In_3150);
xnor U8979 (N_8979,In_3038,In_1462);
xnor U8980 (N_8980,In_4534,In_256);
nand U8981 (N_8981,In_256,In_346);
xor U8982 (N_8982,In_4577,In_2178);
nand U8983 (N_8983,In_1852,In_4660);
nor U8984 (N_8984,In_1586,In_468);
and U8985 (N_8985,In_1054,In_2900);
and U8986 (N_8986,In_3478,In_667);
nor U8987 (N_8987,In_4340,In_549);
nor U8988 (N_8988,In_4140,In_777);
or U8989 (N_8989,In_1015,In_4381);
nand U8990 (N_8990,In_1676,In_3650);
xor U8991 (N_8991,In_116,In_4244);
nand U8992 (N_8992,In_2510,In_1342);
or U8993 (N_8993,In_1442,In_3607);
nor U8994 (N_8994,In_170,In_4178);
nand U8995 (N_8995,In_1857,In_3778);
and U8996 (N_8996,In_359,In_1087);
or U8997 (N_8997,In_2657,In_1022);
and U8998 (N_8998,In_1501,In_2027);
xor U8999 (N_8999,In_833,In_4414);
nand U9000 (N_9000,In_4342,In_4075);
or U9001 (N_9001,In_3004,In_3056);
or U9002 (N_9002,In_4044,In_3824);
nor U9003 (N_9003,In_2373,In_243);
and U9004 (N_9004,In_2325,In_440);
xnor U9005 (N_9005,In_4024,In_4358);
nor U9006 (N_9006,In_1839,In_4563);
and U9007 (N_9007,In_1244,In_1595);
or U9008 (N_9008,In_4106,In_3740);
or U9009 (N_9009,In_4412,In_3208);
and U9010 (N_9010,In_1910,In_3045);
xor U9011 (N_9011,In_832,In_3614);
nand U9012 (N_9012,In_3799,In_319);
and U9013 (N_9013,In_2587,In_3034);
xnor U9014 (N_9014,In_2834,In_3288);
and U9015 (N_9015,In_1868,In_4334);
nand U9016 (N_9016,In_2870,In_2598);
nor U9017 (N_9017,In_4996,In_569);
and U9018 (N_9018,In_318,In_403);
or U9019 (N_9019,In_4588,In_2311);
and U9020 (N_9020,In_3003,In_3556);
nand U9021 (N_9021,In_2540,In_2652);
xnor U9022 (N_9022,In_1765,In_1968);
and U9023 (N_9023,In_3066,In_4813);
or U9024 (N_9024,In_3576,In_3263);
nand U9025 (N_9025,In_3498,In_506);
and U9026 (N_9026,In_3313,In_4118);
nor U9027 (N_9027,In_4309,In_1544);
or U9028 (N_9028,In_553,In_1904);
or U9029 (N_9029,In_1,In_2449);
or U9030 (N_9030,In_622,In_3566);
and U9031 (N_9031,In_3165,In_4007);
nand U9032 (N_9032,In_4703,In_687);
and U9033 (N_9033,In_227,In_1299);
and U9034 (N_9034,In_1074,In_3433);
and U9035 (N_9035,In_3446,In_2024);
xnor U9036 (N_9036,In_3374,In_1578);
xor U9037 (N_9037,In_3184,In_3484);
or U9038 (N_9038,In_2811,In_3152);
nor U9039 (N_9039,In_12,In_2679);
or U9040 (N_9040,In_2281,In_2261);
or U9041 (N_9041,In_56,In_689);
or U9042 (N_9042,In_4489,In_1996);
or U9043 (N_9043,In_4776,In_636);
xor U9044 (N_9044,In_3397,In_1503);
or U9045 (N_9045,In_1765,In_2510);
nand U9046 (N_9046,In_2963,In_4253);
nand U9047 (N_9047,In_3737,In_163);
nor U9048 (N_9048,In_451,In_4799);
xor U9049 (N_9049,In_4124,In_922);
or U9050 (N_9050,In_3609,In_1071);
or U9051 (N_9051,In_2987,In_4788);
xnor U9052 (N_9052,In_3603,In_863);
xor U9053 (N_9053,In_2249,In_1914);
or U9054 (N_9054,In_3045,In_3853);
nand U9055 (N_9055,In_1074,In_978);
nor U9056 (N_9056,In_213,In_2273);
or U9057 (N_9057,In_2044,In_631);
xor U9058 (N_9058,In_2232,In_45);
nor U9059 (N_9059,In_2449,In_3778);
or U9060 (N_9060,In_3684,In_4375);
nor U9061 (N_9061,In_2356,In_2354);
and U9062 (N_9062,In_1347,In_1584);
and U9063 (N_9063,In_2024,In_423);
or U9064 (N_9064,In_1190,In_1784);
nand U9065 (N_9065,In_422,In_2176);
nor U9066 (N_9066,In_1326,In_2585);
nand U9067 (N_9067,In_3126,In_4834);
nor U9068 (N_9068,In_1681,In_949);
and U9069 (N_9069,In_1281,In_732);
xor U9070 (N_9070,In_3823,In_4760);
or U9071 (N_9071,In_1239,In_500);
nor U9072 (N_9072,In_3652,In_1549);
xor U9073 (N_9073,In_2476,In_2407);
xnor U9074 (N_9074,In_1952,In_662);
or U9075 (N_9075,In_2488,In_67);
xnor U9076 (N_9076,In_3689,In_1609);
xnor U9077 (N_9077,In_3062,In_3573);
and U9078 (N_9078,In_2689,In_2395);
and U9079 (N_9079,In_1546,In_752);
and U9080 (N_9080,In_406,In_2742);
xnor U9081 (N_9081,In_64,In_1533);
or U9082 (N_9082,In_1802,In_3299);
nand U9083 (N_9083,In_4047,In_308);
and U9084 (N_9084,In_24,In_2814);
or U9085 (N_9085,In_2308,In_4527);
nor U9086 (N_9086,In_2285,In_2546);
xor U9087 (N_9087,In_3190,In_3216);
nand U9088 (N_9088,In_4260,In_2153);
nor U9089 (N_9089,In_4139,In_1869);
xnor U9090 (N_9090,In_908,In_4379);
or U9091 (N_9091,In_4893,In_1720);
and U9092 (N_9092,In_2673,In_824);
and U9093 (N_9093,In_4736,In_411);
nand U9094 (N_9094,In_702,In_620);
or U9095 (N_9095,In_4363,In_2120);
xor U9096 (N_9096,In_3629,In_50);
xnor U9097 (N_9097,In_462,In_2568);
nor U9098 (N_9098,In_2037,In_3536);
or U9099 (N_9099,In_2633,In_3509);
or U9100 (N_9100,In_3312,In_2018);
or U9101 (N_9101,In_399,In_2074);
nand U9102 (N_9102,In_1185,In_4969);
nand U9103 (N_9103,In_1023,In_4154);
nor U9104 (N_9104,In_571,In_4374);
nor U9105 (N_9105,In_851,In_2321);
and U9106 (N_9106,In_778,In_3090);
and U9107 (N_9107,In_1475,In_966);
and U9108 (N_9108,In_1894,In_2712);
and U9109 (N_9109,In_476,In_80);
nand U9110 (N_9110,In_3840,In_916);
xnor U9111 (N_9111,In_4679,In_4912);
or U9112 (N_9112,In_375,In_780);
and U9113 (N_9113,In_2674,In_879);
and U9114 (N_9114,In_338,In_1003);
or U9115 (N_9115,In_4213,In_1434);
nand U9116 (N_9116,In_2694,In_1777);
or U9117 (N_9117,In_2938,In_902);
and U9118 (N_9118,In_1240,In_4751);
or U9119 (N_9119,In_4683,In_2899);
nor U9120 (N_9120,In_3113,In_3666);
nand U9121 (N_9121,In_1828,In_2404);
nor U9122 (N_9122,In_856,In_3060);
and U9123 (N_9123,In_4642,In_1240);
nand U9124 (N_9124,In_2299,In_1665);
nand U9125 (N_9125,In_3159,In_2399);
xnor U9126 (N_9126,In_217,In_3369);
xnor U9127 (N_9127,In_1874,In_1025);
and U9128 (N_9128,In_557,In_3952);
nor U9129 (N_9129,In_1400,In_4127);
nand U9130 (N_9130,In_4214,In_4529);
nand U9131 (N_9131,In_502,In_3576);
and U9132 (N_9132,In_3675,In_1867);
xnor U9133 (N_9133,In_2697,In_4333);
or U9134 (N_9134,In_1519,In_4566);
or U9135 (N_9135,In_3058,In_4995);
or U9136 (N_9136,In_1436,In_1532);
xor U9137 (N_9137,In_4106,In_2453);
nor U9138 (N_9138,In_3700,In_4682);
or U9139 (N_9139,In_4330,In_1395);
or U9140 (N_9140,In_4281,In_3511);
nor U9141 (N_9141,In_2151,In_3052);
nand U9142 (N_9142,In_2006,In_1039);
xnor U9143 (N_9143,In_3958,In_1170);
or U9144 (N_9144,In_1369,In_1101);
nand U9145 (N_9145,In_3961,In_1863);
nor U9146 (N_9146,In_4852,In_4703);
nand U9147 (N_9147,In_1841,In_4224);
xnor U9148 (N_9148,In_136,In_2017);
or U9149 (N_9149,In_3354,In_1396);
nand U9150 (N_9150,In_2225,In_3890);
nor U9151 (N_9151,In_813,In_1083);
nand U9152 (N_9152,In_2007,In_3446);
nand U9153 (N_9153,In_1585,In_434);
nand U9154 (N_9154,In_424,In_1463);
or U9155 (N_9155,In_4406,In_528);
nor U9156 (N_9156,In_2364,In_4787);
nand U9157 (N_9157,In_2556,In_3237);
xnor U9158 (N_9158,In_3385,In_2442);
xnor U9159 (N_9159,In_3016,In_29);
xor U9160 (N_9160,In_3277,In_1418);
xnor U9161 (N_9161,In_1048,In_3762);
nand U9162 (N_9162,In_483,In_4697);
and U9163 (N_9163,In_1142,In_1892);
nand U9164 (N_9164,In_676,In_2806);
and U9165 (N_9165,In_4394,In_2680);
and U9166 (N_9166,In_1108,In_3693);
nand U9167 (N_9167,In_4355,In_208);
or U9168 (N_9168,In_2676,In_848);
xor U9169 (N_9169,In_2034,In_4703);
nand U9170 (N_9170,In_3504,In_3287);
and U9171 (N_9171,In_3795,In_2092);
xor U9172 (N_9172,In_3099,In_4307);
nand U9173 (N_9173,In_2612,In_4140);
nand U9174 (N_9174,In_4749,In_1604);
xor U9175 (N_9175,In_1808,In_4582);
or U9176 (N_9176,In_516,In_2143);
xor U9177 (N_9177,In_1741,In_286);
nor U9178 (N_9178,In_4049,In_470);
and U9179 (N_9179,In_1907,In_443);
xnor U9180 (N_9180,In_4838,In_4876);
and U9181 (N_9181,In_2529,In_2762);
and U9182 (N_9182,In_3808,In_2359);
nor U9183 (N_9183,In_2371,In_4033);
xnor U9184 (N_9184,In_2864,In_2975);
nor U9185 (N_9185,In_3904,In_3990);
xnor U9186 (N_9186,In_644,In_1159);
or U9187 (N_9187,In_3338,In_2486);
xor U9188 (N_9188,In_2474,In_228);
and U9189 (N_9189,In_2387,In_1558);
or U9190 (N_9190,In_760,In_4650);
xor U9191 (N_9191,In_1010,In_3699);
or U9192 (N_9192,In_518,In_3769);
nand U9193 (N_9193,In_4235,In_4005);
nor U9194 (N_9194,In_2769,In_630);
xor U9195 (N_9195,In_58,In_3825);
nand U9196 (N_9196,In_2838,In_4448);
nor U9197 (N_9197,In_1130,In_1799);
nand U9198 (N_9198,In_1887,In_4702);
nand U9199 (N_9199,In_3958,In_4223);
or U9200 (N_9200,In_4761,In_2511);
xnor U9201 (N_9201,In_4631,In_488);
or U9202 (N_9202,In_4337,In_3115);
xor U9203 (N_9203,In_1351,In_621);
nor U9204 (N_9204,In_3573,In_2152);
nand U9205 (N_9205,In_1951,In_3115);
and U9206 (N_9206,In_4434,In_4945);
or U9207 (N_9207,In_2435,In_1078);
and U9208 (N_9208,In_2134,In_213);
and U9209 (N_9209,In_2780,In_1706);
and U9210 (N_9210,In_2946,In_991);
and U9211 (N_9211,In_2459,In_746);
xor U9212 (N_9212,In_3029,In_3245);
or U9213 (N_9213,In_1428,In_4707);
xnor U9214 (N_9214,In_3059,In_2805);
or U9215 (N_9215,In_707,In_1810);
nor U9216 (N_9216,In_436,In_2585);
and U9217 (N_9217,In_25,In_1706);
and U9218 (N_9218,In_1130,In_4926);
xor U9219 (N_9219,In_4981,In_932);
or U9220 (N_9220,In_3059,In_1563);
or U9221 (N_9221,In_4739,In_4697);
or U9222 (N_9222,In_1465,In_3606);
nor U9223 (N_9223,In_650,In_3204);
xnor U9224 (N_9224,In_1438,In_2876);
and U9225 (N_9225,In_4373,In_96);
or U9226 (N_9226,In_811,In_2425);
nand U9227 (N_9227,In_3160,In_4010);
nor U9228 (N_9228,In_43,In_1599);
nand U9229 (N_9229,In_294,In_2813);
or U9230 (N_9230,In_4421,In_3976);
xnor U9231 (N_9231,In_4441,In_4153);
nor U9232 (N_9232,In_3075,In_4211);
or U9233 (N_9233,In_716,In_2282);
and U9234 (N_9234,In_1294,In_4041);
nor U9235 (N_9235,In_3617,In_3271);
xnor U9236 (N_9236,In_3865,In_3416);
xor U9237 (N_9237,In_2634,In_2275);
or U9238 (N_9238,In_3756,In_1979);
or U9239 (N_9239,In_225,In_1922);
or U9240 (N_9240,In_4534,In_502);
or U9241 (N_9241,In_971,In_3229);
or U9242 (N_9242,In_1781,In_4501);
xnor U9243 (N_9243,In_4830,In_4203);
or U9244 (N_9244,In_1197,In_820);
nor U9245 (N_9245,In_1391,In_202);
nor U9246 (N_9246,In_4226,In_813);
or U9247 (N_9247,In_775,In_493);
nand U9248 (N_9248,In_1629,In_1873);
xor U9249 (N_9249,In_2582,In_592);
xor U9250 (N_9250,In_716,In_1706);
and U9251 (N_9251,In_1907,In_1472);
xnor U9252 (N_9252,In_2550,In_1204);
xor U9253 (N_9253,In_1177,In_2101);
or U9254 (N_9254,In_1393,In_3864);
and U9255 (N_9255,In_977,In_937);
nor U9256 (N_9256,In_2865,In_939);
nand U9257 (N_9257,In_3413,In_3656);
nand U9258 (N_9258,In_1391,In_2365);
nor U9259 (N_9259,In_1420,In_1748);
xor U9260 (N_9260,In_1012,In_1469);
or U9261 (N_9261,In_954,In_360);
nand U9262 (N_9262,In_2482,In_4832);
nand U9263 (N_9263,In_4503,In_1864);
nor U9264 (N_9264,In_1419,In_3816);
nor U9265 (N_9265,In_1436,In_2104);
xor U9266 (N_9266,In_4933,In_2609);
and U9267 (N_9267,In_3726,In_716);
or U9268 (N_9268,In_2451,In_1851);
xnor U9269 (N_9269,In_185,In_1317);
xor U9270 (N_9270,In_3729,In_1102);
nand U9271 (N_9271,In_900,In_993);
and U9272 (N_9272,In_3037,In_2091);
and U9273 (N_9273,In_1360,In_492);
or U9274 (N_9274,In_843,In_4231);
and U9275 (N_9275,In_4934,In_1975);
nand U9276 (N_9276,In_4237,In_363);
xor U9277 (N_9277,In_1984,In_2172);
or U9278 (N_9278,In_4683,In_1982);
nand U9279 (N_9279,In_2970,In_3691);
and U9280 (N_9280,In_2468,In_3108);
nand U9281 (N_9281,In_3769,In_796);
xor U9282 (N_9282,In_4831,In_1005);
nand U9283 (N_9283,In_145,In_1003);
and U9284 (N_9284,In_1088,In_4314);
nor U9285 (N_9285,In_4919,In_4228);
and U9286 (N_9286,In_938,In_3713);
or U9287 (N_9287,In_2703,In_2818);
nor U9288 (N_9288,In_4092,In_2117);
and U9289 (N_9289,In_429,In_1294);
or U9290 (N_9290,In_4633,In_4588);
nor U9291 (N_9291,In_3909,In_4950);
or U9292 (N_9292,In_868,In_3893);
nand U9293 (N_9293,In_3276,In_348);
nor U9294 (N_9294,In_2249,In_2321);
xnor U9295 (N_9295,In_1828,In_1281);
nor U9296 (N_9296,In_3224,In_14);
or U9297 (N_9297,In_2713,In_3651);
xor U9298 (N_9298,In_1943,In_3765);
nand U9299 (N_9299,In_4244,In_2405);
nand U9300 (N_9300,In_2892,In_3123);
nor U9301 (N_9301,In_3515,In_1262);
or U9302 (N_9302,In_985,In_3062);
xor U9303 (N_9303,In_4149,In_533);
or U9304 (N_9304,In_3853,In_4590);
nor U9305 (N_9305,In_2434,In_3418);
or U9306 (N_9306,In_4637,In_504);
xor U9307 (N_9307,In_3705,In_3506);
or U9308 (N_9308,In_4418,In_4035);
or U9309 (N_9309,In_4776,In_4611);
nor U9310 (N_9310,In_2776,In_479);
and U9311 (N_9311,In_1312,In_381);
and U9312 (N_9312,In_3552,In_1882);
xnor U9313 (N_9313,In_275,In_4336);
or U9314 (N_9314,In_1772,In_535);
nor U9315 (N_9315,In_2078,In_4719);
nor U9316 (N_9316,In_1153,In_3565);
nand U9317 (N_9317,In_2296,In_2615);
nand U9318 (N_9318,In_1186,In_4429);
nor U9319 (N_9319,In_659,In_3073);
nand U9320 (N_9320,In_3478,In_1492);
nor U9321 (N_9321,In_3347,In_1113);
xor U9322 (N_9322,In_2457,In_1403);
xnor U9323 (N_9323,In_2457,In_1679);
or U9324 (N_9324,In_3093,In_969);
or U9325 (N_9325,In_2484,In_3047);
nand U9326 (N_9326,In_651,In_554);
xnor U9327 (N_9327,In_4967,In_864);
nor U9328 (N_9328,In_2073,In_1911);
xor U9329 (N_9329,In_1020,In_420);
xnor U9330 (N_9330,In_733,In_560);
or U9331 (N_9331,In_4200,In_3975);
and U9332 (N_9332,In_1092,In_874);
and U9333 (N_9333,In_4248,In_436);
xor U9334 (N_9334,In_4793,In_3679);
or U9335 (N_9335,In_4076,In_1532);
or U9336 (N_9336,In_4270,In_3581);
nor U9337 (N_9337,In_893,In_933);
nand U9338 (N_9338,In_154,In_623);
nand U9339 (N_9339,In_2108,In_2392);
nor U9340 (N_9340,In_4426,In_1300);
xor U9341 (N_9341,In_3217,In_88);
or U9342 (N_9342,In_3366,In_1438);
nand U9343 (N_9343,In_2790,In_2785);
and U9344 (N_9344,In_3843,In_1719);
xnor U9345 (N_9345,In_2023,In_1243);
and U9346 (N_9346,In_76,In_1899);
nor U9347 (N_9347,In_1976,In_2341);
and U9348 (N_9348,In_3716,In_424);
nand U9349 (N_9349,In_234,In_2537);
xor U9350 (N_9350,In_232,In_4105);
xnor U9351 (N_9351,In_120,In_4365);
nor U9352 (N_9352,In_943,In_2537);
or U9353 (N_9353,In_3580,In_3331);
or U9354 (N_9354,In_2638,In_3970);
nand U9355 (N_9355,In_2710,In_2667);
or U9356 (N_9356,In_13,In_988);
or U9357 (N_9357,In_636,In_578);
nor U9358 (N_9358,In_4452,In_3227);
nand U9359 (N_9359,In_4770,In_1993);
xnor U9360 (N_9360,In_3607,In_1304);
or U9361 (N_9361,In_3584,In_48);
xor U9362 (N_9362,In_677,In_2154);
nor U9363 (N_9363,In_1992,In_1218);
nor U9364 (N_9364,In_1470,In_1909);
xnor U9365 (N_9365,In_259,In_3732);
nand U9366 (N_9366,In_4006,In_2254);
and U9367 (N_9367,In_101,In_3624);
xor U9368 (N_9368,In_764,In_1907);
nor U9369 (N_9369,In_4591,In_588);
xor U9370 (N_9370,In_4983,In_4488);
nor U9371 (N_9371,In_4520,In_726);
nor U9372 (N_9372,In_4709,In_656);
or U9373 (N_9373,In_112,In_1170);
or U9374 (N_9374,In_2138,In_3200);
and U9375 (N_9375,In_719,In_1497);
and U9376 (N_9376,In_4162,In_4998);
nand U9377 (N_9377,In_2999,In_4458);
xor U9378 (N_9378,In_908,In_2820);
or U9379 (N_9379,In_2876,In_4261);
nand U9380 (N_9380,In_4657,In_2725);
nor U9381 (N_9381,In_4603,In_3240);
xnor U9382 (N_9382,In_4706,In_738);
nand U9383 (N_9383,In_4485,In_3185);
xnor U9384 (N_9384,In_4900,In_522);
and U9385 (N_9385,In_1336,In_3500);
or U9386 (N_9386,In_1702,In_379);
nor U9387 (N_9387,In_26,In_663);
nor U9388 (N_9388,In_982,In_4772);
nor U9389 (N_9389,In_2781,In_1697);
or U9390 (N_9390,In_1663,In_4096);
nor U9391 (N_9391,In_4187,In_138);
nand U9392 (N_9392,In_3728,In_1827);
or U9393 (N_9393,In_4668,In_2137);
xor U9394 (N_9394,In_1998,In_4295);
nand U9395 (N_9395,In_3783,In_1199);
and U9396 (N_9396,In_4016,In_2197);
nand U9397 (N_9397,In_1423,In_1183);
nor U9398 (N_9398,In_4709,In_2606);
and U9399 (N_9399,In_3731,In_4515);
or U9400 (N_9400,In_1530,In_1441);
nand U9401 (N_9401,In_4223,In_1097);
and U9402 (N_9402,In_356,In_2526);
nand U9403 (N_9403,In_2156,In_818);
or U9404 (N_9404,In_1944,In_4593);
or U9405 (N_9405,In_1043,In_2789);
nor U9406 (N_9406,In_2482,In_2422);
and U9407 (N_9407,In_4935,In_4197);
or U9408 (N_9408,In_770,In_1188);
and U9409 (N_9409,In_648,In_4811);
or U9410 (N_9410,In_4510,In_2326);
and U9411 (N_9411,In_1754,In_2647);
xor U9412 (N_9412,In_564,In_3079);
xor U9413 (N_9413,In_4212,In_3825);
and U9414 (N_9414,In_392,In_2630);
nor U9415 (N_9415,In_2094,In_1883);
or U9416 (N_9416,In_4916,In_4111);
and U9417 (N_9417,In_1772,In_723);
nor U9418 (N_9418,In_4027,In_3101);
or U9419 (N_9419,In_4116,In_311);
and U9420 (N_9420,In_839,In_1808);
nor U9421 (N_9421,In_3970,In_4854);
and U9422 (N_9422,In_3483,In_2152);
and U9423 (N_9423,In_4678,In_4071);
nand U9424 (N_9424,In_3373,In_4860);
and U9425 (N_9425,In_3337,In_315);
nand U9426 (N_9426,In_3709,In_4707);
or U9427 (N_9427,In_1116,In_1790);
nand U9428 (N_9428,In_1697,In_426);
and U9429 (N_9429,In_2904,In_442);
and U9430 (N_9430,In_1797,In_1741);
xor U9431 (N_9431,In_1749,In_1763);
or U9432 (N_9432,In_2834,In_2781);
nand U9433 (N_9433,In_312,In_3971);
xor U9434 (N_9434,In_3341,In_1515);
and U9435 (N_9435,In_3625,In_783);
or U9436 (N_9436,In_4510,In_1274);
nor U9437 (N_9437,In_1029,In_4047);
nand U9438 (N_9438,In_3306,In_1527);
and U9439 (N_9439,In_1873,In_3905);
nor U9440 (N_9440,In_2965,In_3080);
nand U9441 (N_9441,In_3148,In_3827);
and U9442 (N_9442,In_51,In_4880);
xor U9443 (N_9443,In_253,In_897);
nor U9444 (N_9444,In_2227,In_4996);
or U9445 (N_9445,In_1730,In_3383);
nor U9446 (N_9446,In_4072,In_968);
nor U9447 (N_9447,In_3583,In_3755);
xor U9448 (N_9448,In_3169,In_3700);
nand U9449 (N_9449,In_1191,In_3502);
xnor U9450 (N_9450,In_4370,In_4641);
xor U9451 (N_9451,In_3622,In_4302);
and U9452 (N_9452,In_3051,In_370);
xor U9453 (N_9453,In_1229,In_3516);
nand U9454 (N_9454,In_3065,In_155);
xor U9455 (N_9455,In_4983,In_2676);
nor U9456 (N_9456,In_1138,In_4899);
or U9457 (N_9457,In_2371,In_1769);
and U9458 (N_9458,In_3596,In_4937);
nand U9459 (N_9459,In_4108,In_3903);
nand U9460 (N_9460,In_863,In_345);
nand U9461 (N_9461,In_4236,In_2790);
xnor U9462 (N_9462,In_100,In_488);
xor U9463 (N_9463,In_3713,In_822);
or U9464 (N_9464,In_984,In_4470);
nand U9465 (N_9465,In_2488,In_343);
nor U9466 (N_9466,In_2785,In_3539);
or U9467 (N_9467,In_1559,In_4943);
nor U9468 (N_9468,In_1119,In_4324);
xor U9469 (N_9469,In_4021,In_1755);
and U9470 (N_9470,In_4300,In_305);
or U9471 (N_9471,In_376,In_4405);
or U9472 (N_9472,In_591,In_2477);
and U9473 (N_9473,In_1843,In_260);
or U9474 (N_9474,In_472,In_2424);
or U9475 (N_9475,In_957,In_524);
and U9476 (N_9476,In_2692,In_2056);
or U9477 (N_9477,In_2297,In_1830);
nand U9478 (N_9478,In_3913,In_229);
and U9479 (N_9479,In_1578,In_2673);
or U9480 (N_9480,In_1929,In_2570);
nor U9481 (N_9481,In_4064,In_4368);
nor U9482 (N_9482,In_865,In_3604);
xnor U9483 (N_9483,In_4974,In_2282);
xor U9484 (N_9484,In_979,In_2460);
nor U9485 (N_9485,In_2782,In_4242);
nor U9486 (N_9486,In_2543,In_4730);
and U9487 (N_9487,In_469,In_3004);
nand U9488 (N_9488,In_4607,In_2751);
nand U9489 (N_9489,In_2306,In_3667);
and U9490 (N_9490,In_4827,In_702);
xor U9491 (N_9491,In_4977,In_2726);
nor U9492 (N_9492,In_4302,In_263);
or U9493 (N_9493,In_2060,In_1933);
or U9494 (N_9494,In_3812,In_3120);
nand U9495 (N_9495,In_1456,In_1068);
nand U9496 (N_9496,In_709,In_2070);
and U9497 (N_9497,In_1295,In_2118);
nand U9498 (N_9498,In_4911,In_1093);
nor U9499 (N_9499,In_978,In_2936);
xnor U9500 (N_9500,In_805,In_4949);
or U9501 (N_9501,In_1419,In_2088);
or U9502 (N_9502,In_3530,In_3901);
and U9503 (N_9503,In_2671,In_720);
and U9504 (N_9504,In_517,In_1186);
and U9505 (N_9505,In_3851,In_257);
xnor U9506 (N_9506,In_1073,In_3391);
nor U9507 (N_9507,In_2344,In_2545);
xnor U9508 (N_9508,In_4132,In_475);
nor U9509 (N_9509,In_1433,In_111);
nand U9510 (N_9510,In_2037,In_2944);
nand U9511 (N_9511,In_3956,In_990);
nor U9512 (N_9512,In_4222,In_616);
and U9513 (N_9513,In_3656,In_1872);
xor U9514 (N_9514,In_418,In_3793);
or U9515 (N_9515,In_4391,In_3445);
nand U9516 (N_9516,In_1488,In_3184);
xor U9517 (N_9517,In_3893,In_1553);
xnor U9518 (N_9518,In_3529,In_4609);
and U9519 (N_9519,In_3757,In_2528);
xor U9520 (N_9520,In_3817,In_1568);
nor U9521 (N_9521,In_211,In_56);
nor U9522 (N_9522,In_4422,In_2312);
nor U9523 (N_9523,In_2840,In_2236);
nor U9524 (N_9524,In_2414,In_220);
nor U9525 (N_9525,In_721,In_1596);
xor U9526 (N_9526,In_4629,In_2693);
xor U9527 (N_9527,In_3260,In_2621);
xor U9528 (N_9528,In_3287,In_4647);
and U9529 (N_9529,In_2697,In_2304);
or U9530 (N_9530,In_16,In_736);
and U9531 (N_9531,In_2887,In_2510);
and U9532 (N_9532,In_2927,In_4984);
xnor U9533 (N_9533,In_1729,In_3322);
nand U9534 (N_9534,In_2966,In_230);
xnor U9535 (N_9535,In_3293,In_1320);
nor U9536 (N_9536,In_4899,In_4895);
xnor U9537 (N_9537,In_4319,In_3065);
xnor U9538 (N_9538,In_2319,In_3341);
nand U9539 (N_9539,In_4510,In_4241);
or U9540 (N_9540,In_3739,In_4607);
xor U9541 (N_9541,In_446,In_963);
nand U9542 (N_9542,In_2143,In_3698);
and U9543 (N_9543,In_2339,In_2686);
nand U9544 (N_9544,In_1630,In_3678);
or U9545 (N_9545,In_2450,In_505);
nor U9546 (N_9546,In_3748,In_939);
xor U9547 (N_9547,In_799,In_2210);
and U9548 (N_9548,In_1761,In_1198);
nand U9549 (N_9549,In_4081,In_3881);
xnor U9550 (N_9550,In_3523,In_1041);
or U9551 (N_9551,In_4073,In_3749);
or U9552 (N_9552,In_2847,In_2646);
or U9553 (N_9553,In_1532,In_4029);
and U9554 (N_9554,In_784,In_1449);
nand U9555 (N_9555,In_1029,In_1184);
xnor U9556 (N_9556,In_2442,In_4303);
nor U9557 (N_9557,In_1271,In_3169);
nor U9558 (N_9558,In_4982,In_711);
xor U9559 (N_9559,In_3422,In_1265);
nor U9560 (N_9560,In_3277,In_4479);
nand U9561 (N_9561,In_4281,In_350);
xnor U9562 (N_9562,In_4955,In_3162);
and U9563 (N_9563,In_1853,In_690);
nor U9564 (N_9564,In_2765,In_1771);
nand U9565 (N_9565,In_3986,In_1406);
and U9566 (N_9566,In_145,In_2607);
nand U9567 (N_9567,In_1691,In_3772);
and U9568 (N_9568,In_3257,In_4372);
and U9569 (N_9569,In_1626,In_2584);
nor U9570 (N_9570,In_186,In_1387);
or U9571 (N_9571,In_4744,In_344);
or U9572 (N_9572,In_1312,In_2110);
xnor U9573 (N_9573,In_794,In_2856);
nand U9574 (N_9574,In_4988,In_3851);
and U9575 (N_9575,In_3542,In_1234);
nor U9576 (N_9576,In_1060,In_1008);
nand U9577 (N_9577,In_2115,In_1706);
and U9578 (N_9578,In_1265,In_114);
and U9579 (N_9579,In_2773,In_1130);
nor U9580 (N_9580,In_4925,In_1998);
and U9581 (N_9581,In_4889,In_1698);
nor U9582 (N_9582,In_4550,In_4294);
nand U9583 (N_9583,In_2174,In_2364);
or U9584 (N_9584,In_2122,In_2219);
and U9585 (N_9585,In_1326,In_1138);
xnor U9586 (N_9586,In_2721,In_1529);
nand U9587 (N_9587,In_1130,In_2540);
nand U9588 (N_9588,In_3537,In_3279);
nand U9589 (N_9589,In_2988,In_2321);
or U9590 (N_9590,In_1375,In_448);
nand U9591 (N_9591,In_4543,In_1546);
xnor U9592 (N_9592,In_1182,In_2184);
xor U9593 (N_9593,In_282,In_2495);
xnor U9594 (N_9594,In_3603,In_491);
or U9595 (N_9595,In_3309,In_1375);
and U9596 (N_9596,In_1442,In_1644);
or U9597 (N_9597,In_1241,In_3955);
nand U9598 (N_9598,In_3410,In_3605);
nand U9599 (N_9599,In_46,In_1085);
or U9600 (N_9600,In_1789,In_3626);
and U9601 (N_9601,In_2706,In_2644);
or U9602 (N_9602,In_4867,In_434);
and U9603 (N_9603,In_4237,In_2391);
or U9604 (N_9604,In_1986,In_4925);
and U9605 (N_9605,In_3749,In_1704);
xnor U9606 (N_9606,In_4403,In_1031);
or U9607 (N_9607,In_4766,In_4265);
or U9608 (N_9608,In_23,In_2304);
and U9609 (N_9609,In_1464,In_368);
or U9610 (N_9610,In_4739,In_291);
or U9611 (N_9611,In_3505,In_1552);
nor U9612 (N_9612,In_4643,In_4349);
and U9613 (N_9613,In_3465,In_4837);
nand U9614 (N_9614,In_3598,In_4585);
or U9615 (N_9615,In_285,In_322);
and U9616 (N_9616,In_2093,In_3130);
and U9617 (N_9617,In_4634,In_1632);
or U9618 (N_9618,In_3032,In_3227);
nand U9619 (N_9619,In_2763,In_2758);
xor U9620 (N_9620,In_2046,In_2169);
xnor U9621 (N_9621,In_3125,In_764);
and U9622 (N_9622,In_2142,In_825);
or U9623 (N_9623,In_1191,In_1205);
nor U9624 (N_9624,In_2799,In_886);
nand U9625 (N_9625,In_104,In_3491);
nand U9626 (N_9626,In_671,In_1972);
nor U9627 (N_9627,In_1674,In_589);
xnor U9628 (N_9628,In_2254,In_120);
or U9629 (N_9629,In_4537,In_2282);
xor U9630 (N_9630,In_4555,In_1561);
nand U9631 (N_9631,In_4998,In_2811);
or U9632 (N_9632,In_4804,In_3654);
nor U9633 (N_9633,In_3981,In_553);
or U9634 (N_9634,In_3955,In_1123);
nand U9635 (N_9635,In_1671,In_916);
xor U9636 (N_9636,In_678,In_3500);
or U9637 (N_9637,In_1836,In_450);
nor U9638 (N_9638,In_2250,In_812);
and U9639 (N_9639,In_2935,In_3235);
nand U9640 (N_9640,In_4387,In_1901);
and U9641 (N_9641,In_2284,In_533);
and U9642 (N_9642,In_1139,In_4054);
nor U9643 (N_9643,In_87,In_3814);
or U9644 (N_9644,In_1811,In_3428);
and U9645 (N_9645,In_954,In_4457);
or U9646 (N_9646,In_2826,In_1658);
and U9647 (N_9647,In_357,In_3857);
or U9648 (N_9648,In_791,In_4119);
xor U9649 (N_9649,In_4480,In_2310);
and U9650 (N_9650,In_344,In_1057);
or U9651 (N_9651,In_4879,In_2086);
xor U9652 (N_9652,In_3730,In_2705);
or U9653 (N_9653,In_2980,In_4866);
and U9654 (N_9654,In_3067,In_3835);
or U9655 (N_9655,In_601,In_4331);
and U9656 (N_9656,In_651,In_1189);
nand U9657 (N_9657,In_4581,In_4228);
nor U9658 (N_9658,In_2882,In_47);
nand U9659 (N_9659,In_339,In_4869);
nand U9660 (N_9660,In_3766,In_3081);
nand U9661 (N_9661,In_4131,In_373);
and U9662 (N_9662,In_1727,In_2191);
and U9663 (N_9663,In_4105,In_4777);
or U9664 (N_9664,In_176,In_1314);
or U9665 (N_9665,In_1191,In_868);
nand U9666 (N_9666,In_103,In_1043);
nand U9667 (N_9667,In_4905,In_813);
nor U9668 (N_9668,In_345,In_4743);
and U9669 (N_9669,In_4978,In_3427);
or U9670 (N_9670,In_3604,In_1929);
or U9671 (N_9671,In_4077,In_4841);
and U9672 (N_9672,In_2882,In_3470);
nand U9673 (N_9673,In_1040,In_251);
nand U9674 (N_9674,In_2697,In_3840);
or U9675 (N_9675,In_1413,In_797);
nor U9676 (N_9676,In_3662,In_4340);
or U9677 (N_9677,In_3811,In_4429);
or U9678 (N_9678,In_1897,In_4837);
xnor U9679 (N_9679,In_4667,In_4771);
nor U9680 (N_9680,In_4513,In_2910);
and U9681 (N_9681,In_3039,In_1223);
or U9682 (N_9682,In_3575,In_1656);
and U9683 (N_9683,In_4264,In_3592);
nand U9684 (N_9684,In_3366,In_2910);
and U9685 (N_9685,In_1901,In_1303);
nor U9686 (N_9686,In_2669,In_2285);
xor U9687 (N_9687,In_2191,In_1369);
and U9688 (N_9688,In_2121,In_2254);
xor U9689 (N_9689,In_3113,In_3233);
and U9690 (N_9690,In_3384,In_1571);
xor U9691 (N_9691,In_1273,In_3139);
nand U9692 (N_9692,In_4158,In_2514);
xor U9693 (N_9693,In_4344,In_1229);
nor U9694 (N_9694,In_4358,In_1868);
xnor U9695 (N_9695,In_703,In_1086);
xor U9696 (N_9696,In_2802,In_3594);
nor U9697 (N_9697,In_2803,In_1340);
and U9698 (N_9698,In_4604,In_3910);
or U9699 (N_9699,In_2406,In_1838);
nand U9700 (N_9700,In_1811,In_3854);
nor U9701 (N_9701,In_4372,In_4504);
nand U9702 (N_9702,In_1885,In_765);
nand U9703 (N_9703,In_1274,In_2438);
or U9704 (N_9704,In_1688,In_2345);
nor U9705 (N_9705,In_4290,In_1818);
xor U9706 (N_9706,In_3753,In_1365);
xnor U9707 (N_9707,In_4202,In_4760);
nand U9708 (N_9708,In_4975,In_2716);
nand U9709 (N_9709,In_3379,In_1196);
or U9710 (N_9710,In_3904,In_4524);
nor U9711 (N_9711,In_776,In_3282);
nand U9712 (N_9712,In_2384,In_1955);
xor U9713 (N_9713,In_339,In_2372);
xnor U9714 (N_9714,In_1583,In_4489);
xnor U9715 (N_9715,In_26,In_2720);
or U9716 (N_9716,In_3250,In_3183);
nand U9717 (N_9717,In_4674,In_3011);
nor U9718 (N_9718,In_2042,In_329);
or U9719 (N_9719,In_3632,In_3186);
or U9720 (N_9720,In_187,In_3263);
and U9721 (N_9721,In_501,In_1412);
nor U9722 (N_9722,In_53,In_2819);
or U9723 (N_9723,In_2579,In_4313);
xnor U9724 (N_9724,In_2715,In_2669);
and U9725 (N_9725,In_4589,In_874);
or U9726 (N_9726,In_3868,In_4605);
nor U9727 (N_9727,In_2046,In_1875);
and U9728 (N_9728,In_786,In_4156);
nand U9729 (N_9729,In_4382,In_3337);
nor U9730 (N_9730,In_184,In_4127);
and U9731 (N_9731,In_410,In_569);
or U9732 (N_9732,In_695,In_3814);
xor U9733 (N_9733,In_1288,In_701);
and U9734 (N_9734,In_1628,In_215);
nand U9735 (N_9735,In_1013,In_3421);
nor U9736 (N_9736,In_3188,In_4012);
xnor U9737 (N_9737,In_3600,In_3921);
xor U9738 (N_9738,In_4083,In_4225);
or U9739 (N_9739,In_815,In_330);
or U9740 (N_9740,In_581,In_881);
nand U9741 (N_9741,In_195,In_3183);
and U9742 (N_9742,In_2731,In_3603);
nor U9743 (N_9743,In_60,In_4605);
or U9744 (N_9744,In_2903,In_4856);
nor U9745 (N_9745,In_2470,In_4691);
nand U9746 (N_9746,In_3649,In_3982);
or U9747 (N_9747,In_1354,In_2360);
and U9748 (N_9748,In_4467,In_2571);
nand U9749 (N_9749,In_4218,In_4972);
nand U9750 (N_9750,In_380,In_825);
and U9751 (N_9751,In_216,In_2710);
or U9752 (N_9752,In_2959,In_1303);
xnor U9753 (N_9753,In_3250,In_53);
xor U9754 (N_9754,In_1796,In_1507);
nand U9755 (N_9755,In_4223,In_2004);
or U9756 (N_9756,In_3473,In_1081);
xnor U9757 (N_9757,In_3384,In_885);
nand U9758 (N_9758,In_2040,In_879);
and U9759 (N_9759,In_2590,In_1484);
and U9760 (N_9760,In_4342,In_1538);
nor U9761 (N_9761,In_907,In_3784);
xor U9762 (N_9762,In_4288,In_3985);
or U9763 (N_9763,In_4747,In_2110);
nor U9764 (N_9764,In_1714,In_627);
and U9765 (N_9765,In_1349,In_4677);
nand U9766 (N_9766,In_4265,In_2347);
nor U9767 (N_9767,In_4725,In_37);
and U9768 (N_9768,In_4148,In_703);
or U9769 (N_9769,In_1274,In_3795);
xor U9770 (N_9770,In_3806,In_1347);
nand U9771 (N_9771,In_2836,In_582);
nor U9772 (N_9772,In_3454,In_699);
nand U9773 (N_9773,In_1943,In_1421);
nand U9774 (N_9774,In_3369,In_579);
nor U9775 (N_9775,In_31,In_3207);
nand U9776 (N_9776,In_4798,In_2648);
xnor U9777 (N_9777,In_1524,In_176);
or U9778 (N_9778,In_242,In_1071);
nor U9779 (N_9779,In_4730,In_2720);
or U9780 (N_9780,In_655,In_2464);
or U9781 (N_9781,In_1961,In_3635);
nand U9782 (N_9782,In_2261,In_406);
and U9783 (N_9783,In_2289,In_3989);
xnor U9784 (N_9784,In_1930,In_2401);
or U9785 (N_9785,In_947,In_4681);
nand U9786 (N_9786,In_759,In_2767);
nor U9787 (N_9787,In_4032,In_4538);
and U9788 (N_9788,In_3615,In_2309);
nor U9789 (N_9789,In_3287,In_3861);
xnor U9790 (N_9790,In_4040,In_4114);
nand U9791 (N_9791,In_1587,In_3308);
nor U9792 (N_9792,In_931,In_1561);
nor U9793 (N_9793,In_4733,In_2084);
xnor U9794 (N_9794,In_4901,In_3428);
nor U9795 (N_9795,In_2598,In_1876);
xor U9796 (N_9796,In_4428,In_2355);
xor U9797 (N_9797,In_4933,In_2350);
or U9798 (N_9798,In_4181,In_3212);
or U9799 (N_9799,In_4059,In_1117);
nand U9800 (N_9800,In_4404,In_4045);
nor U9801 (N_9801,In_1178,In_940);
nand U9802 (N_9802,In_2284,In_240);
xor U9803 (N_9803,In_2077,In_3911);
nand U9804 (N_9804,In_4235,In_1290);
or U9805 (N_9805,In_332,In_3794);
nor U9806 (N_9806,In_2558,In_3971);
nor U9807 (N_9807,In_2986,In_98);
xnor U9808 (N_9808,In_4677,In_3315);
or U9809 (N_9809,In_3552,In_4760);
or U9810 (N_9810,In_4136,In_221);
nand U9811 (N_9811,In_1963,In_866);
xnor U9812 (N_9812,In_4366,In_418);
nor U9813 (N_9813,In_1385,In_2147);
and U9814 (N_9814,In_2599,In_4253);
xor U9815 (N_9815,In_1058,In_4918);
xor U9816 (N_9816,In_322,In_472);
nand U9817 (N_9817,In_3845,In_1505);
xnor U9818 (N_9818,In_2638,In_3255);
nand U9819 (N_9819,In_292,In_614);
xor U9820 (N_9820,In_2089,In_356);
nor U9821 (N_9821,In_2756,In_1083);
nor U9822 (N_9822,In_1545,In_4430);
nor U9823 (N_9823,In_2241,In_2827);
and U9824 (N_9824,In_4512,In_4440);
or U9825 (N_9825,In_136,In_2049);
nor U9826 (N_9826,In_1014,In_903);
nor U9827 (N_9827,In_129,In_4066);
xor U9828 (N_9828,In_4675,In_2294);
nor U9829 (N_9829,In_796,In_329);
xnor U9830 (N_9830,In_4764,In_4188);
nand U9831 (N_9831,In_945,In_3060);
nand U9832 (N_9832,In_1966,In_2367);
or U9833 (N_9833,In_3249,In_2830);
and U9834 (N_9834,In_665,In_4507);
or U9835 (N_9835,In_4014,In_1079);
nand U9836 (N_9836,In_681,In_3489);
nand U9837 (N_9837,In_1554,In_1255);
nor U9838 (N_9838,In_478,In_1541);
nor U9839 (N_9839,In_3243,In_3503);
and U9840 (N_9840,In_4028,In_1256);
or U9841 (N_9841,In_4762,In_1504);
nand U9842 (N_9842,In_1407,In_3352);
xor U9843 (N_9843,In_4854,In_1425);
nor U9844 (N_9844,In_119,In_2922);
and U9845 (N_9845,In_3994,In_1716);
and U9846 (N_9846,In_1001,In_1112);
nand U9847 (N_9847,In_4874,In_3763);
xnor U9848 (N_9848,In_192,In_3550);
xor U9849 (N_9849,In_2909,In_280);
nor U9850 (N_9850,In_3446,In_2400);
nor U9851 (N_9851,In_3885,In_4330);
and U9852 (N_9852,In_1688,In_1217);
nor U9853 (N_9853,In_35,In_1883);
xor U9854 (N_9854,In_4465,In_756);
nor U9855 (N_9855,In_856,In_1707);
or U9856 (N_9856,In_2202,In_2336);
and U9857 (N_9857,In_2037,In_1779);
or U9858 (N_9858,In_4638,In_4410);
nand U9859 (N_9859,In_4622,In_3429);
or U9860 (N_9860,In_1892,In_2046);
xor U9861 (N_9861,In_1439,In_826);
nor U9862 (N_9862,In_3393,In_1632);
or U9863 (N_9863,In_2641,In_4564);
and U9864 (N_9864,In_1906,In_1721);
or U9865 (N_9865,In_1369,In_2333);
nor U9866 (N_9866,In_823,In_1138);
or U9867 (N_9867,In_3089,In_2358);
nand U9868 (N_9868,In_1266,In_1909);
and U9869 (N_9869,In_3363,In_1335);
and U9870 (N_9870,In_748,In_4725);
and U9871 (N_9871,In_3773,In_990);
nor U9872 (N_9872,In_848,In_3662);
xnor U9873 (N_9873,In_4235,In_3551);
nor U9874 (N_9874,In_20,In_4165);
and U9875 (N_9875,In_4436,In_1693);
or U9876 (N_9876,In_4878,In_4220);
nor U9877 (N_9877,In_2107,In_3518);
and U9878 (N_9878,In_717,In_1141);
nor U9879 (N_9879,In_1949,In_4516);
or U9880 (N_9880,In_2563,In_2514);
and U9881 (N_9881,In_3663,In_3828);
and U9882 (N_9882,In_4374,In_3218);
and U9883 (N_9883,In_3541,In_1459);
xnor U9884 (N_9884,In_2432,In_1212);
nor U9885 (N_9885,In_4360,In_3220);
or U9886 (N_9886,In_850,In_610);
and U9887 (N_9887,In_4933,In_2955);
nor U9888 (N_9888,In_4681,In_2904);
and U9889 (N_9889,In_2151,In_2888);
xor U9890 (N_9890,In_2351,In_2061);
or U9891 (N_9891,In_2743,In_1131);
nor U9892 (N_9892,In_4790,In_3835);
nand U9893 (N_9893,In_589,In_3331);
nand U9894 (N_9894,In_4958,In_2179);
xnor U9895 (N_9895,In_456,In_4238);
xnor U9896 (N_9896,In_4315,In_1726);
nor U9897 (N_9897,In_826,In_4456);
xnor U9898 (N_9898,In_1025,In_648);
nor U9899 (N_9899,In_1777,In_4300);
or U9900 (N_9900,In_4901,In_585);
nand U9901 (N_9901,In_4902,In_1319);
xnor U9902 (N_9902,In_3941,In_4921);
nand U9903 (N_9903,In_1915,In_1512);
and U9904 (N_9904,In_273,In_783);
nor U9905 (N_9905,In_1217,In_1743);
nor U9906 (N_9906,In_4850,In_48);
nand U9907 (N_9907,In_4756,In_50);
xnor U9908 (N_9908,In_1217,In_2115);
nor U9909 (N_9909,In_4725,In_2569);
nor U9910 (N_9910,In_1927,In_4205);
or U9911 (N_9911,In_1757,In_4263);
and U9912 (N_9912,In_1018,In_3605);
nand U9913 (N_9913,In_3760,In_3635);
nor U9914 (N_9914,In_2445,In_1594);
nor U9915 (N_9915,In_1603,In_4521);
xnor U9916 (N_9916,In_4186,In_2221);
nor U9917 (N_9917,In_4875,In_1873);
nand U9918 (N_9918,In_1126,In_4048);
or U9919 (N_9919,In_2551,In_3567);
nor U9920 (N_9920,In_2936,In_171);
nand U9921 (N_9921,In_4967,In_3284);
and U9922 (N_9922,In_10,In_1416);
or U9923 (N_9923,In_2161,In_1581);
nand U9924 (N_9924,In_4967,In_275);
nand U9925 (N_9925,In_1749,In_1651);
nand U9926 (N_9926,In_1791,In_2093);
nor U9927 (N_9927,In_3245,In_3935);
xor U9928 (N_9928,In_1057,In_4137);
and U9929 (N_9929,In_2811,In_1072);
nand U9930 (N_9930,In_826,In_3100);
nor U9931 (N_9931,In_1529,In_544);
nor U9932 (N_9932,In_1724,In_3813);
nand U9933 (N_9933,In_4464,In_4714);
nor U9934 (N_9934,In_1477,In_2735);
xor U9935 (N_9935,In_2679,In_4586);
nor U9936 (N_9936,In_3715,In_4153);
and U9937 (N_9937,In_4151,In_941);
xnor U9938 (N_9938,In_3594,In_2057);
and U9939 (N_9939,In_4970,In_4050);
nor U9940 (N_9940,In_4290,In_1552);
nand U9941 (N_9941,In_911,In_2686);
nand U9942 (N_9942,In_1884,In_1943);
nor U9943 (N_9943,In_2589,In_450);
and U9944 (N_9944,In_4432,In_2668);
nand U9945 (N_9945,In_2763,In_2048);
and U9946 (N_9946,In_2909,In_3937);
nand U9947 (N_9947,In_1088,In_4986);
and U9948 (N_9948,In_4173,In_1245);
nand U9949 (N_9949,In_4623,In_4632);
and U9950 (N_9950,In_38,In_587);
and U9951 (N_9951,In_3866,In_4264);
or U9952 (N_9952,In_2532,In_4773);
nor U9953 (N_9953,In_2914,In_2229);
and U9954 (N_9954,In_112,In_2173);
xor U9955 (N_9955,In_317,In_3437);
and U9956 (N_9956,In_4434,In_4837);
nor U9957 (N_9957,In_3670,In_3431);
and U9958 (N_9958,In_2890,In_4269);
or U9959 (N_9959,In_4822,In_108);
and U9960 (N_9960,In_3782,In_1632);
xnor U9961 (N_9961,In_2479,In_3981);
nor U9962 (N_9962,In_2768,In_14);
nor U9963 (N_9963,In_802,In_4788);
xor U9964 (N_9964,In_3367,In_1107);
xor U9965 (N_9965,In_2652,In_3469);
nor U9966 (N_9966,In_329,In_3425);
and U9967 (N_9967,In_2977,In_2309);
and U9968 (N_9968,In_3451,In_1583);
nor U9969 (N_9969,In_3183,In_4626);
xor U9970 (N_9970,In_910,In_3472);
xor U9971 (N_9971,In_4618,In_3417);
nand U9972 (N_9972,In_2092,In_1261);
nand U9973 (N_9973,In_2060,In_1774);
or U9974 (N_9974,In_1865,In_1408);
xnor U9975 (N_9975,In_2223,In_1848);
nor U9976 (N_9976,In_4030,In_2912);
or U9977 (N_9977,In_2895,In_1879);
and U9978 (N_9978,In_2378,In_2641);
xor U9979 (N_9979,In_1298,In_4561);
and U9980 (N_9980,In_1750,In_4687);
nor U9981 (N_9981,In_1636,In_2052);
xor U9982 (N_9982,In_3866,In_2479);
nand U9983 (N_9983,In_3812,In_1309);
and U9984 (N_9984,In_3554,In_3117);
and U9985 (N_9985,In_4508,In_2518);
nor U9986 (N_9986,In_2223,In_3840);
nor U9987 (N_9987,In_122,In_680);
or U9988 (N_9988,In_568,In_1367);
nor U9989 (N_9989,In_4083,In_263);
nand U9990 (N_9990,In_4541,In_3862);
xor U9991 (N_9991,In_4142,In_4446);
or U9992 (N_9992,In_2393,In_1323);
nor U9993 (N_9993,In_3175,In_23);
and U9994 (N_9994,In_2236,In_1909);
nor U9995 (N_9995,In_2895,In_2607);
xor U9996 (N_9996,In_2713,In_1948);
or U9997 (N_9997,In_4431,In_2656);
xor U9998 (N_9998,In_3275,In_439);
xnor U9999 (N_9999,In_3152,In_1583);
xnor U10000 (N_10000,N_2672,N_1274);
nand U10001 (N_10001,N_3925,N_1854);
nand U10002 (N_10002,N_7602,N_1420);
nand U10003 (N_10003,N_9746,N_3835);
or U10004 (N_10004,N_1713,N_6590);
or U10005 (N_10005,N_8324,N_6831);
xnor U10006 (N_10006,N_9367,N_9195);
or U10007 (N_10007,N_7222,N_2119);
nor U10008 (N_10008,N_9381,N_1810);
or U10009 (N_10009,N_9018,N_7201);
xnor U10010 (N_10010,N_7237,N_5455);
and U10011 (N_10011,N_900,N_1368);
nor U10012 (N_10012,N_2422,N_7058);
xnor U10013 (N_10013,N_3489,N_4948);
and U10014 (N_10014,N_5120,N_1291);
nand U10015 (N_10015,N_2569,N_9790);
nand U10016 (N_10016,N_1724,N_9371);
nor U10017 (N_10017,N_6046,N_7961);
nand U10018 (N_10018,N_4527,N_5728);
nor U10019 (N_10019,N_7018,N_9206);
and U10020 (N_10020,N_3104,N_1223);
nand U10021 (N_10021,N_919,N_7012);
xor U10022 (N_10022,N_161,N_6652);
nand U10023 (N_10023,N_5906,N_4469);
nor U10024 (N_10024,N_5016,N_1321);
or U10025 (N_10025,N_6268,N_1313);
xor U10026 (N_10026,N_7798,N_8970);
nor U10027 (N_10027,N_8217,N_3233);
xor U10028 (N_10028,N_9393,N_3607);
nor U10029 (N_10029,N_2163,N_3764);
and U10030 (N_10030,N_5939,N_4793);
xor U10031 (N_10031,N_2988,N_935);
nor U10032 (N_10032,N_6205,N_4556);
or U10033 (N_10033,N_9154,N_5741);
or U10034 (N_10034,N_95,N_3068);
nor U10035 (N_10035,N_8377,N_4043);
nor U10036 (N_10036,N_9428,N_1186);
nor U10037 (N_10037,N_9836,N_7215);
xor U10038 (N_10038,N_9952,N_2616);
nand U10039 (N_10039,N_2198,N_4292);
nor U10040 (N_10040,N_5571,N_7987);
or U10041 (N_10041,N_1714,N_3804);
nand U10042 (N_10042,N_9651,N_5577);
xor U10043 (N_10043,N_9288,N_1612);
nand U10044 (N_10044,N_8816,N_3945);
nand U10045 (N_10045,N_1793,N_6463);
or U10046 (N_10046,N_2041,N_6350);
xnor U10047 (N_10047,N_7642,N_3743);
xnor U10048 (N_10048,N_7354,N_7467);
nor U10049 (N_10049,N_7581,N_5951);
and U10050 (N_10050,N_1865,N_5627);
nor U10051 (N_10051,N_530,N_153);
nor U10052 (N_10052,N_9950,N_2493);
nand U10053 (N_10053,N_5042,N_53);
and U10054 (N_10054,N_5900,N_3491);
nor U10055 (N_10055,N_6497,N_9033);
nand U10056 (N_10056,N_163,N_885);
nand U10057 (N_10057,N_4392,N_1988);
or U10058 (N_10058,N_949,N_4156);
nand U10059 (N_10059,N_5838,N_2202);
xnor U10060 (N_10060,N_30,N_4311);
nand U10061 (N_10061,N_9189,N_8381);
or U10062 (N_10062,N_866,N_9917);
nor U10063 (N_10063,N_9242,N_7331);
or U10064 (N_10064,N_2221,N_2517);
and U10065 (N_10065,N_8955,N_9147);
nor U10066 (N_10066,N_2328,N_5987);
nand U10067 (N_10067,N_1893,N_442);
nor U10068 (N_10068,N_8658,N_1058);
nor U10069 (N_10069,N_587,N_7179);
nand U10070 (N_10070,N_5158,N_6687);
nor U10071 (N_10071,N_5148,N_1438);
nor U10072 (N_10072,N_7316,N_2767);
or U10073 (N_10073,N_9722,N_5108);
nand U10074 (N_10074,N_5256,N_3363);
nor U10075 (N_10075,N_678,N_1962);
and U10076 (N_10076,N_2206,N_3957);
or U10077 (N_10077,N_5129,N_1795);
xor U10078 (N_10078,N_4279,N_7944);
xnor U10079 (N_10079,N_1170,N_4443);
and U10080 (N_10080,N_8547,N_2568);
nor U10081 (N_10081,N_9920,N_1095);
nand U10082 (N_10082,N_1551,N_4174);
and U10083 (N_10083,N_8245,N_7119);
nor U10084 (N_10084,N_3094,N_3229);
and U10085 (N_10085,N_7950,N_9820);
nand U10086 (N_10086,N_3396,N_4909);
or U10087 (N_10087,N_4838,N_6611);
xnor U10088 (N_10088,N_7688,N_9126);
xor U10089 (N_10089,N_9134,N_1545);
nand U10090 (N_10090,N_8441,N_3189);
xnor U10091 (N_10091,N_3838,N_1237);
and U10092 (N_10092,N_1658,N_1760);
xor U10093 (N_10093,N_4489,N_1720);
nor U10094 (N_10094,N_6646,N_9323);
nand U10095 (N_10095,N_4275,N_680);
or U10096 (N_10096,N_3402,N_7823);
xnor U10097 (N_10097,N_45,N_9785);
or U10098 (N_10098,N_1176,N_792);
xnor U10099 (N_10099,N_3531,N_3300);
nand U10100 (N_10100,N_6902,N_3712);
xor U10101 (N_10101,N_5971,N_7868);
xnor U10102 (N_10102,N_9496,N_6018);
nand U10103 (N_10103,N_1045,N_5667);
nand U10104 (N_10104,N_7779,N_9934);
nand U10105 (N_10105,N_4518,N_3685);
and U10106 (N_10106,N_6088,N_9776);
nor U10107 (N_10107,N_7031,N_9404);
nand U10108 (N_10108,N_3534,N_4015);
nand U10109 (N_10109,N_9877,N_6345);
nor U10110 (N_10110,N_3322,N_7052);
nor U10111 (N_10111,N_1933,N_3387);
nor U10112 (N_10112,N_8841,N_1202);
nand U10113 (N_10113,N_5177,N_3254);
or U10114 (N_10114,N_6802,N_5657);
or U10115 (N_10115,N_5972,N_2310);
xnor U10116 (N_10116,N_1901,N_2900);
nor U10117 (N_10117,N_201,N_3959);
or U10118 (N_10118,N_3965,N_9554);
nor U10119 (N_10119,N_6025,N_5499);
and U10120 (N_10120,N_5468,N_9852);
nand U10121 (N_10121,N_1887,N_9417);
nand U10122 (N_10122,N_7223,N_423);
and U10123 (N_10123,N_2277,N_9841);
or U10124 (N_10124,N_6411,N_8232);
or U10125 (N_10125,N_6780,N_2696);
nand U10126 (N_10126,N_7909,N_2682);
nand U10127 (N_10127,N_3813,N_6840);
nor U10128 (N_10128,N_6850,N_1566);
nand U10129 (N_10129,N_4192,N_581);
or U10130 (N_10130,N_6891,N_9439);
nand U10131 (N_10131,N_8261,N_4308);
nor U10132 (N_10132,N_34,N_4103);
xnor U10133 (N_10133,N_5022,N_1514);
nand U10134 (N_10134,N_3049,N_4595);
nand U10135 (N_10135,N_5157,N_3983);
and U10136 (N_10136,N_3878,N_8801);
and U10137 (N_10137,N_6371,N_2986);
nand U10138 (N_10138,N_1035,N_8409);
xnor U10139 (N_10139,N_431,N_1452);
or U10140 (N_10140,N_6667,N_5918);
or U10141 (N_10141,N_7922,N_8253);
or U10142 (N_10142,N_4678,N_8842);
nand U10143 (N_10143,N_1794,N_6974);
and U10144 (N_10144,N_5990,N_7558);
or U10145 (N_10145,N_4792,N_4030);
nand U10146 (N_10146,N_4837,N_2182);
nand U10147 (N_10147,N_2944,N_5798);
nor U10148 (N_10148,N_2674,N_5562);
or U10149 (N_10149,N_9986,N_9320);
and U10150 (N_10150,N_1635,N_7572);
and U10151 (N_10151,N_64,N_3532);
nor U10152 (N_10152,N_9642,N_822);
xnor U10153 (N_10153,N_4369,N_3741);
xnor U10154 (N_10154,N_5373,N_7079);
nand U10155 (N_10155,N_7549,N_3120);
xnor U10156 (N_10156,N_6940,N_7797);
xor U10157 (N_10157,N_7208,N_3354);
and U10158 (N_10158,N_6766,N_2273);
nor U10159 (N_10159,N_8432,N_6030);
nand U10160 (N_10160,N_6063,N_446);
xor U10161 (N_10161,N_9310,N_1198);
or U10162 (N_10162,N_987,N_3435);
or U10163 (N_10163,N_5031,N_7173);
nand U10164 (N_10164,N_4362,N_7840);
xnor U10165 (N_10165,N_9679,N_1442);
and U10166 (N_10166,N_5843,N_8962);
and U10167 (N_10167,N_8230,N_7154);
or U10168 (N_10168,N_6991,N_4941);
xor U10169 (N_10169,N_3313,N_6420);
or U10170 (N_10170,N_4355,N_2800);
nor U10171 (N_10171,N_1173,N_2520);
and U10172 (N_10172,N_8083,N_6679);
and U10173 (N_10173,N_4516,N_8960);
and U10174 (N_10174,N_8934,N_1801);
xnor U10175 (N_10175,N_2430,N_7376);
or U10176 (N_10176,N_4132,N_5954);
and U10177 (N_10177,N_1864,N_4379);
xnor U10178 (N_10178,N_1337,N_5904);
nor U10179 (N_10179,N_3181,N_2385);
nor U10180 (N_10180,N_2720,N_7323);
and U10181 (N_10181,N_9041,N_7414);
xnor U10182 (N_10182,N_6271,N_5779);
nand U10183 (N_10183,N_7738,N_4214);
or U10184 (N_10184,N_1323,N_2439);
or U10185 (N_10185,N_3679,N_7406);
xnor U10186 (N_10186,N_7594,N_7404);
nor U10187 (N_10187,N_8267,N_1130);
or U10188 (N_10188,N_6035,N_1244);
and U10189 (N_10189,N_6932,N_9080);
nand U10190 (N_10190,N_3759,N_7311);
nor U10191 (N_10191,N_8176,N_6695);
and U10192 (N_10192,N_4503,N_3502);
or U10193 (N_10193,N_1390,N_8746);
nor U10194 (N_10194,N_2378,N_5644);
nor U10195 (N_10195,N_7678,N_7605);
xnor U10196 (N_10196,N_5655,N_2579);
xor U10197 (N_10197,N_2412,N_8480);
nor U10198 (N_10198,N_1536,N_6134);
xor U10199 (N_10199,N_9044,N_4223);
xor U10200 (N_10200,N_3516,N_1968);
xor U10201 (N_10201,N_1266,N_9477);
nor U10202 (N_10202,N_9083,N_9284);
or U10203 (N_10203,N_105,N_1593);
nor U10204 (N_10204,N_3087,N_9394);
and U10205 (N_10205,N_1428,N_2689);
or U10206 (N_10206,N_280,N_2731);
and U10207 (N_10207,N_1603,N_6860);
or U10208 (N_10208,N_4317,N_9379);
or U10209 (N_10209,N_3521,N_6503);
xor U10210 (N_10210,N_1596,N_6790);
xor U10211 (N_10211,N_6630,N_4973);
or U10212 (N_10212,N_4217,N_4294);
and U10213 (N_10213,N_7141,N_2225);
xnor U10214 (N_10214,N_5212,N_4890);
nor U10215 (N_10215,N_4680,N_590);
and U10216 (N_10216,N_300,N_5066);
xnor U10217 (N_10217,N_4861,N_9185);
nand U10218 (N_10218,N_9475,N_6150);
nand U10219 (N_10219,N_8513,N_5163);
xnor U10220 (N_10220,N_762,N_1026);
xor U10221 (N_10221,N_9494,N_7622);
or U10222 (N_10222,N_8391,N_4552);
nand U10223 (N_10223,N_5605,N_5492);
nor U10224 (N_10224,N_1333,N_7117);
nand U10225 (N_10225,N_9817,N_2455);
and U10226 (N_10226,N_2686,N_8206);
nand U10227 (N_10227,N_1624,N_6935);
nand U10228 (N_10228,N_1791,N_5982);
nand U10229 (N_10229,N_2706,N_6622);
nand U10230 (N_10230,N_4044,N_3618);
nand U10231 (N_10231,N_3298,N_975);
nand U10232 (N_10232,N_5382,N_9916);
nand U10233 (N_10233,N_1505,N_9434);
or U10234 (N_10234,N_1064,N_2442);
xnor U10235 (N_10235,N_7802,N_2364);
nand U10236 (N_10236,N_3921,N_9429);
nand U10237 (N_10237,N_7607,N_3606);
nand U10238 (N_10238,N_930,N_8259);
nor U10239 (N_10239,N_6725,N_9566);
nor U10240 (N_10240,N_8285,N_1446);
nor U10241 (N_10241,N_1383,N_3836);
and U10242 (N_10242,N_8941,N_8758);
and U10243 (N_10243,N_1370,N_5710);
nand U10244 (N_10244,N_5343,N_9029);
xor U10245 (N_10245,N_5725,N_6793);
and U10246 (N_10246,N_9876,N_8881);
nor U10247 (N_10247,N_7280,N_8007);
and U10248 (N_10248,N_3698,N_9015);
and U10249 (N_10249,N_7300,N_6635);
nand U10250 (N_10250,N_8454,N_6617);
xor U10251 (N_10251,N_5857,N_3433);
nor U10252 (N_10252,N_964,N_4849);
xor U10253 (N_10253,N_8202,N_728);
nand U10254 (N_10254,N_436,N_2826);
and U10255 (N_10255,N_9303,N_5764);
nand U10256 (N_10256,N_8527,N_9060);
nand U10257 (N_10257,N_2427,N_2852);
nand U10258 (N_10258,N_3978,N_5955);
xnor U10259 (N_10259,N_1060,N_4583);
xnor U10260 (N_10260,N_8976,N_3259);
and U10261 (N_10261,N_6381,N_863);
or U10262 (N_10262,N_4148,N_7664);
and U10263 (N_10263,N_7281,N_9214);
or U10264 (N_10264,N_8444,N_4900);
xnor U10265 (N_10265,N_9598,N_3503);
xor U10266 (N_10266,N_9692,N_6762);
or U10267 (N_10267,N_9944,N_5340);
nand U10268 (N_10268,N_8016,N_3112);
nand U10269 (N_10269,N_6825,N_571);
or U10270 (N_10270,N_2700,N_8251);
and U10271 (N_10271,N_8753,N_1703);
or U10272 (N_10272,N_6151,N_9431);
and U10273 (N_10273,N_7461,N_1028);
xor U10274 (N_10274,N_5994,N_2236);
and U10275 (N_10275,N_6255,N_715);
xor U10276 (N_10276,N_4025,N_6696);
xor U10277 (N_10277,N_1093,N_903);
or U10278 (N_10278,N_6884,N_1777);
nor U10279 (N_10279,N_8477,N_5181);
nand U10280 (N_10280,N_2240,N_3816);
or U10281 (N_10281,N_2037,N_8902);
and U10282 (N_10282,N_670,N_2080);
nand U10283 (N_10283,N_8281,N_9939);
and U10284 (N_10284,N_6224,N_8191);
or U10285 (N_10285,N_1640,N_6147);
and U10286 (N_10286,N_1056,N_5919);
or U10287 (N_10287,N_8370,N_3639);
and U10288 (N_10288,N_2046,N_4955);
xnor U10289 (N_10289,N_5606,N_4466);
nand U10290 (N_10290,N_9529,N_3237);
xnor U10291 (N_10291,N_3217,N_2088);
xor U10292 (N_10292,N_7303,N_8598);
and U10293 (N_10293,N_1102,N_698);
nand U10294 (N_10294,N_8482,N_9666);
xnor U10295 (N_10295,N_1388,N_7442);
nand U10296 (N_10296,N_3885,N_2538);
xor U10297 (N_10297,N_250,N_6480);
nor U10298 (N_10298,N_7927,N_2460);
or U10299 (N_10299,N_5176,N_5043);
or U10300 (N_10300,N_9095,N_7537);
or U10301 (N_10301,N_3117,N_6426);
nand U10302 (N_10302,N_8306,N_8378);
or U10303 (N_10303,N_1554,N_1577);
and U10304 (N_10304,N_6355,N_9601);
or U10305 (N_10305,N_3522,N_2334);
or U10306 (N_10306,N_6299,N_5705);
and U10307 (N_10307,N_9864,N_653);
nor U10308 (N_10308,N_6783,N_372);
and U10309 (N_10309,N_2681,N_6698);
and U10310 (N_10310,N_9525,N_2213);
xor U10311 (N_10311,N_1645,N_1386);
xor U10312 (N_10312,N_9948,N_9592);
and U10313 (N_10313,N_2913,N_4698);
nand U10314 (N_10314,N_8108,N_9549);
nand U10315 (N_10315,N_9299,N_6619);
nand U10316 (N_10316,N_1105,N_7039);
nand U10317 (N_10317,N_370,N_239);
nor U10318 (N_10318,N_1969,N_152);
xnor U10319 (N_10319,N_8028,N_7546);
and U10320 (N_10320,N_6072,N_7648);
and U10321 (N_10321,N_8362,N_3127);
nand U10322 (N_10322,N_6859,N_1487);
or U10323 (N_10323,N_8994,N_5740);
nor U10324 (N_10324,N_3557,N_5103);
nand U10325 (N_10325,N_2670,N_2001);
and U10326 (N_10326,N_2023,N_5143);
xnor U10327 (N_10327,N_6903,N_2584);
or U10328 (N_10328,N_3798,N_7197);
nor U10329 (N_10329,N_1262,N_9714);
nand U10330 (N_10330,N_9341,N_2070);
nand U10331 (N_10331,N_936,N_2224);
nor U10332 (N_10332,N_9838,N_7574);
xor U10333 (N_10333,N_323,N_9168);
and U10334 (N_10334,N_3533,N_3670);
nand U10335 (N_10335,N_6005,N_1678);
and U10336 (N_10336,N_1844,N_2630);
nand U10337 (N_10337,N_7974,N_17);
and U10338 (N_10338,N_8386,N_4018);
xor U10339 (N_10339,N_4615,N_4730);
and U10340 (N_10340,N_2139,N_5200);
nor U10341 (N_10341,N_6591,N_1157);
nand U10342 (N_10342,N_2489,N_6244);
nand U10343 (N_10343,N_3873,N_813);
nor U10344 (N_10344,N_9520,N_8868);
nand U10345 (N_10345,N_205,N_8874);
and U10346 (N_10346,N_6526,N_5882);
nand U10347 (N_10347,N_7464,N_7832);
nand U10348 (N_10348,N_6736,N_3960);
nor U10349 (N_10349,N_636,N_8866);
nor U10350 (N_10350,N_3968,N_2739);
nand U10351 (N_10351,N_5563,N_6614);
or U10352 (N_10352,N_6518,N_6111);
nor U10353 (N_10353,N_9268,N_8105);
or U10354 (N_10354,N_6894,N_4324);
and U10355 (N_10355,N_4638,N_8484);
xnor U10356 (N_10356,N_8905,N_2234);
xor U10357 (N_10357,N_9249,N_6259);
and U10358 (N_10358,N_8857,N_4335);
nand U10359 (N_10359,N_6867,N_8805);
nand U10360 (N_10360,N_8294,N_737);
or U10361 (N_10361,N_2264,N_9064);
and U10362 (N_10362,N_6776,N_1427);
xnor U10363 (N_10363,N_3182,N_9845);
xnor U10364 (N_10364,N_8783,N_2887);
nand U10365 (N_10365,N_1089,N_5805);
nand U10366 (N_10366,N_9472,N_9133);
or U10367 (N_10367,N_614,N_2220);
nand U10368 (N_10368,N_3343,N_1851);
and U10369 (N_10369,N_8468,N_5953);
or U10370 (N_10370,N_2744,N_9031);
nand U10371 (N_10371,N_3486,N_7431);
or U10372 (N_10372,N_1936,N_9207);
xnor U10373 (N_10373,N_9996,N_9359);
or U10374 (N_10374,N_1314,N_7737);
nor U10375 (N_10375,N_2166,N_7518);
xnor U10376 (N_10376,N_8160,N_7011);
and U10377 (N_10377,N_3981,N_9806);
and U10378 (N_10378,N_5858,N_4681);
and U10379 (N_10379,N_6814,N_4841);
or U10380 (N_10380,N_9114,N_2146);
nor U10381 (N_10381,N_20,N_1985);
xor U10382 (N_10382,N_1842,N_960);
or U10383 (N_10383,N_9724,N_4999);
or U10384 (N_10384,N_6997,N_6418);
xor U10385 (N_10385,N_9582,N_5684);
nand U10386 (N_10386,N_4962,N_2861);
or U10387 (N_10387,N_60,N_734);
nor U10388 (N_10388,N_7385,N_6785);
xor U10389 (N_10389,N_3169,N_293);
and U10390 (N_10390,N_4901,N_6848);
nand U10391 (N_10391,N_1905,N_9690);
nand U10392 (N_10392,N_9823,N_5826);
nand U10393 (N_10393,N_2649,N_8461);
xor U10394 (N_10394,N_9291,N_5626);
nand U10395 (N_10395,N_8609,N_1238);
nor U10396 (N_10396,N_3512,N_9077);
nand U10397 (N_10397,N_1124,N_1354);
nor U10398 (N_10398,N_3875,N_4045);
and U10399 (N_10399,N_200,N_2548);
nor U10400 (N_10400,N_3766,N_6367);
nor U10401 (N_10401,N_988,N_8396);
or U10402 (N_10402,N_7878,N_230);
nand U10403 (N_10403,N_6678,N_4415);
nor U10404 (N_10404,N_2192,N_6880);
and U10405 (N_10405,N_5559,N_2177);
nor U10406 (N_10406,N_5012,N_8789);
nor U10407 (N_10407,N_8578,N_5734);
and U10408 (N_10408,N_6399,N_1459);
and U10409 (N_10409,N_2884,N_5364);
nand U10410 (N_10410,N_9059,N_172);
or U10411 (N_10411,N_2076,N_9336);
and U10412 (N_10412,N_9966,N_7920);
or U10413 (N_10413,N_4884,N_8924);
and U10414 (N_10414,N_3819,N_8161);
nor U10415 (N_10415,N_8595,N_1391);
and U10416 (N_10416,N_2624,N_7796);
nand U10417 (N_10417,N_9935,N_6094);
xnor U10418 (N_10418,N_7369,N_2938);
xnor U10419 (N_10419,N_2771,N_4927);
nor U10420 (N_10420,N_9192,N_9608);
and U10421 (N_10421,N_3567,N_2824);
xor U10422 (N_10422,N_7524,N_5665);
nor U10423 (N_10423,N_8893,N_1680);
nand U10424 (N_10424,N_9631,N_2063);
nor U10425 (N_10425,N_963,N_7040);
xnor U10426 (N_10426,N_6349,N_9686);
xnor U10427 (N_10427,N_8530,N_5489);
nand U10428 (N_10428,N_270,N_1350);
xnor U10429 (N_10429,N_6099,N_5548);
nand U10430 (N_10430,N_7116,N_946);
or U10431 (N_10431,N_3197,N_2457);
nand U10432 (N_10432,N_1860,N_7207);
nand U10433 (N_10433,N_4546,N_8743);
nand U10434 (N_10434,N_1445,N_8951);
nor U10435 (N_10435,N_796,N_4989);
nand U10436 (N_10436,N_9383,N_4567);
and U10437 (N_10437,N_2976,N_7067);
or U10438 (N_10438,N_4474,N_6765);
or U10439 (N_10439,N_8124,N_4601);
xor U10440 (N_10440,N_4716,N_4700);
and U10441 (N_10441,N_8626,N_3572);
nor U10442 (N_10442,N_1627,N_7761);
xnor U10443 (N_10443,N_497,N_5417);
or U10444 (N_10444,N_5718,N_770);
nor U10445 (N_10445,N_1464,N_2332);
and U10446 (N_10446,N_8063,N_7060);
or U10447 (N_10447,N_7349,N_7722);
xnor U10448 (N_10448,N_750,N_9687);
nand U10449 (N_10449,N_2226,N_438);
nor U10450 (N_10450,N_3966,N_3635);
and U10451 (N_10451,N_8811,N_9758);
or U10452 (N_10452,N_3504,N_1482);
nor U10453 (N_10453,N_9344,N_9363);
nor U10454 (N_10454,N_8077,N_6798);
nand U10455 (N_10455,N_9648,N_9158);
or U10456 (N_10456,N_6174,N_9204);
or U10457 (N_10457,N_906,N_2204);
nand U10458 (N_10458,N_2935,N_2582);
or U10459 (N_10459,N_6298,N_9617);
or U10460 (N_10460,N_4671,N_3923);
nor U10461 (N_10461,N_6359,N_1139);
and U10462 (N_10462,N_4189,N_8721);
xor U10463 (N_10463,N_7482,N_274);
nand U10464 (N_10464,N_9880,N_6842);
and U10465 (N_10465,N_1435,N_2003);
nor U10466 (N_10466,N_1841,N_9016);
nor U10467 (N_10467,N_1717,N_8701);
and U10468 (N_10468,N_5604,N_1053);
nand U10469 (N_10469,N_4748,N_7361);
nor U10470 (N_10470,N_6753,N_8804);
nand U10471 (N_10471,N_5888,N_985);
xor U10472 (N_10472,N_6612,N_5395);
or U10473 (N_10473,N_79,N_6801);
or U10474 (N_10474,N_4936,N_6358);
and U10475 (N_10475,N_8825,N_1524);
nand U10476 (N_10476,N_8313,N_7611);
nand U10477 (N_10477,N_9965,N_7843);
and U10478 (N_10478,N_4404,N_9334);
nand U10479 (N_10479,N_2526,N_9091);
nor U10480 (N_10480,N_4811,N_1142);
xnor U10481 (N_10481,N_4391,N_5753);
nand U10482 (N_10482,N_2144,N_4077);
and U10483 (N_10483,N_5254,N_1357);
or U10484 (N_10484,N_8776,N_1516);
nand U10485 (N_10485,N_3370,N_7585);
nor U10486 (N_10486,N_2009,N_6050);
and U10487 (N_10487,N_1533,N_8489);
nand U10488 (N_10488,N_2563,N_1707);
nor U10489 (N_10489,N_3781,N_544);
nor U10490 (N_10490,N_154,N_7366);
nand U10491 (N_10491,N_5532,N_9868);
xnor U10492 (N_10492,N_2788,N_3481);
and U10493 (N_10493,N_6507,N_7983);
nor U10494 (N_10494,N_7899,N_740);
nor U10495 (N_10495,N_4542,N_3938);
xor U10496 (N_10496,N_4490,N_335);
xnor U10497 (N_10497,N_3391,N_6839);
and U10498 (N_10498,N_8583,N_2289);
or U10499 (N_10499,N_976,N_6653);
xor U10500 (N_10500,N_4816,N_7310);
nand U10501 (N_10501,N_9725,N_3317);
or U10502 (N_10502,N_3004,N_7334);
nor U10503 (N_10503,N_6338,N_9269);
or U10504 (N_10504,N_6486,N_7876);
nor U10505 (N_10505,N_1136,N_6362);
and U10506 (N_10506,N_5799,N_4218);
and U10507 (N_10507,N_5261,N_2250);
and U10508 (N_10508,N_3682,N_5476);
nor U10509 (N_10509,N_6330,N_8154);
nand U10510 (N_10510,N_4194,N_6686);
xnor U10511 (N_10511,N_2636,N_8695);
and U10512 (N_10512,N_6703,N_4422);
xor U10513 (N_10513,N_5768,N_9832);
nor U10514 (N_10514,N_4150,N_3397);
nor U10515 (N_10515,N_8367,N_6768);
or U10516 (N_10516,N_4460,N_2372);
nor U10517 (N_10517,N_1955,N_9246);
and U10518 (N_10518,N_7240,N_1282);
nor U10519 (N_10519,N_5003,N_7996);
or U10520 (N_10520,N_4677,N_7707);
nand U10521 (N_10521,N_115,N_3024);
xor U10522 (N_10522,N_8034,N_4857);
xor U10523 (N_10523,N_3642,N_6374);
nand U10524 (N_10524,N_7851,N_3305);
and U10525 (N_10525,N_9442,N_6058);
or U10526 (N_10526,N_8299,N_9156);
or U10527 (N_10527,N_2479,N_1751);
nand U10528 (N_10528,N_9127,N_6238);
or U10529 (N_10529,N_3100,N_2469);
or U10530 (N_10530,N_7837,N_3671);
and U10531 (N_10531,N_3003,N_354);
xnor U10532 (N_10532,N_7817,N_905);
nand U10533 (N_10533,N_9304,N_4885);
nor U10534 (N_10534,N_7907,N_2725);
or U10535 (N_10535,N_717,N_8283);
and U10536 (N_10536,N_8446,N_5062);
nand U10537 (N_10537,N_5247,N_3508);
or U10538 (N_10538,N_1254,N_159);
nand U10539 (N_10539,N_2205,N_4207);
or U10540 (N_10540,N_3047,N_3703);
nand U10541 (N_10541,N_1944,N_5406);
or U10542 (N_10542,N_5393,N_8133);
xnor U10543 (N_10543,N_6745,N_4676);
and U10544 (N_10544,N_9049,N_3107);
xnor U10545 (N_10545,N_3043,N_62);
nor U10546 (N_10546,N_5018,N_8946);
nand U10547 (N_10547,N_5234,N_6067);
xnor U10548 (N_10548,N_6960,N_2137);
nand U10549 (N_10549,N_6657,N_1853);
xnor U10550 (N_10550,N_927,N_3332);
and U10551 (N_10551,N_9165,N_9079);
nand U10552 (N_10552,N_4157,N_5403);
xor U10553 (N_10553,N_505,N_5026);
and U10554 (N_10554,N_9337,N_6521);
and U10555 (N_10555,N_495,N_1937);
xor U10556 (N_10556,N_8241,N_6158);
or U10557 (N_10557,N_9867,N_5866);
or U10558 (N_10558,N_1250,N_2160);
xnor U10559 (N_10559,N_1377,N_7499);
nor U10560 (N_10560,N_7653,N_3115);
or U10561 (N_10561,N_3152,N_3824);
nor U10562 (N_10562,N_7778,N_145);
xor U10563 (N_10563,N_8687,N_7142);
xor U10564 (N_10564,N_752,N_4301);
xnor U10565 (N_10565,N_6162,N_937);
nor U10566 (N_10566,N_2280,N_9819);
or U10567 (N_10567,N_4163,N_9452);
or U10568 (N_10568,N_5637,N_6654);
and U10569 (N_10569,N_7985,N_4351);
or U10570 (N_10570,N_2930,N_6325);
or U10571 (N_10571,N_7473,N_7054);
xor U10572 (N_10572,N_9775,N_5631);
nor U10573 (N_10573,N_2934,N_5568);
nor U10574 (N_10574,N_3162,N_7150);
nand U10575 (N_10575,N_3431,N_4953);
or U10576 (N_10576,N_7619,N_6452);
nor U10577 (N_10577,N_8221,N_1052);
xnor U10578 (N_10578,N_7398,N_212);
and U10579 (N_10579,N_118,N_8222);
nand U10580 (N_10580,N_8334,N_5362);
xnor U10581 (N_10581,N_6572,N_6317);
and U10582 (N_10582,N_4720,N_1356);
nand U10583 (N_10583,N_4235,N_329);
or U10584 (N_10584,N_5054,N_1183);
xor U10585 (N_10585,N_5367,N_3702);
xor U10586 (N_10586,N_1694,N_1838);
or U10587 (N_10587,N_4541,N_7428);
or U10588 (N_10588,N_9345,N_7535);
xnor U10589 (N_10589,N_9879,N_2266);
and U10590 (N_10590,N_803,N_7147);
and U10591 (N_10591,N_1242,N_4417);
nor U10592 (N_10592,N_46,N_2834);
or U10593 (N_10593,N_1004,N_6375);
and U10594 (N_10594,N_4461,N_4634);
nor U10595 (N_10595,N_5293,N_4115);
or U10596 (N_10596,N_4104,N_5376);
nor U10597 (N_10597,N_5794,N_4902);
nand U10598 (N_10598,N_6879,N_2962);
nand U10599 (N_10599,N_8449,N_6112);
nand U10600 (N_10600,N_7380,N_4633);
and U10601 (N_10601,N_2084,N_9712);
nor U10602 (N_10602,N_7801,N_2183);
and U10603 (N_10603,N_3211,N_2603);
nand U10604 (N_10604,N_327,N_5319);
nand U10605 (N_10605,N_3140,N_6055);
nor U10606 (N_10606,N_3543,N_313);
or U10607 (N_10607,N_7387,N_4667);
and U10608 (N_10608,N_1908,N_1318);
xnor U10609 (N_10609,N_6242,N_6575);
nor U10610 (N_10610,N_3829,N_3931);
or U10611 (N_10611,N_2723,N_3186);
nor U10612 (N_10612,N_3715,N_8337);
nand U10613 (N_10613,N_7734,N_7506);
and U10614 (N_10614,N_6354,N_4920);
and U10615 (N_10615,N_9640,N_3949);
xor U10616 (N_10616,N_2470,N_8806);
nor U10617 (N_10617,N_6217,N_2879);
or U10618 (N_10618,N_6208,N_8376);
or U10619 (N_10619,N_6144,N_4361);
and U10620 (N_10620,N_2741,N_5441);
and U10621 (N_10621,N_7759,N_5976);
nor U10622 (N_10622,N_6387,N_466);
or U10623 (N_10623,N_9658,N_4874);
xor U10624 (N_10624,N_3713,N_4219);
and U10625 (N_10625,N_8260,N_7363);
and U10626 (N_10626,N_4852,N_1231);
xnor U10627 (N_10627,N_264,N_7273);
and U10628 (N_10628,N_2919,N_1802);
and U10629 (N_10629,N_1351,N_5375);
xor U10630 (N_10630,N_4435,N_7695);
nand U10631 (N_10631,N_4886,N_1453);
and U10632 (N_10632,N_5235,N_5890);
xor U10633 (N_10633,N_6984,N_4568);
or U10634 (N_10634,N_4967,N_5738);
nand U10635 (N_10635,N_9628,N_9427);
nor U10636 (N_10636,N_5930,N_4446);
or U10637 (N_10637,N_4140,N_3158);
or U10638 (N_10638,N_4644,N_851);
nor U10639 (N_10639,N_4477,N_2283);
nand U10640 (N_10640,N_6951,N_6000);
nor U10641 (N_10641,N_1138,N_9102);
and U10642 (N_10642,N_4256,N_3753);
xnor U10643 (N_10643,N_1657,N_8277);
xnor U10644 (N_10644,N_6292,N_5775);
nand U10645 (N_10645,N_4585,N_7402);
nand U10646 (N_10646,N_8662,N_891);
nand U10647 (N_10647,N_3701,N_3240);
and U10648 (N_10648,N_6648,N_6669);
and U10649 (N_10649,N_8653,N_1473);
xnor U10650 (N_10650,N_4453,N_5613);
xnor U10651 (N_10651,N_9137,N_282);
nand U10652 (N_10652,N_3148,N_5767);
or U10653 (N_10653,N_1716,N_3016);
nand U10654 (N_10654,N_5208,N_7791);
or U10655 (N_10655,N_1820,N_4467);
nor U10656 (N_10656,N_1484,N_9201);
or U10657 (N_10657,N_4260,N_8047);
or U10658 (N_10658,N_5889,N_203);
nand U10659 (N_10659,N_2370,N_5192);
nor U10660 (N_10660,N_1348,N_3840);
nand U10661 (N_10661,N_4124,N_5850);
or U10662 (N_10662,N_4385,N_4805);
nand U10663 (N_10663,N_2684,N_5482);
nand U10664 (N_10664,N_6501,N_7603);
or U10665 (N_10665,N_5961,N_23);
and U10666 (N_10666,N_8602,N_834);
nor U10667 (N_10667,N_8846,N_9277);
xor U10668 (N_10668,N_225,N_4062);
xnor U10669 (N_10669,N_6624,N_3942);
xnor U10670 (N_10670,N_2075,N_1210);
or U10671 (N_10671,N_7757,N_831);
or U10672 (N_10672,N_2839,N_6851);
and U10673 (N_10673,N_7038,N_910);
and U10674 (N_10674,N_1207,N_855);
or U10675 (N_10675,N_6539,N_9361);
xnor U10676 (N_10676,N_6618,N_8213);
nand U10677 (N_10677,N_782,N_1579);
xor U10678 (N_10678,N_3950,N_3154);
and U10679 (N_10679,N_228,N_5916);
nand U10680 (N_10680,N_8520,N_8781);
or U10681 (N_10681,N_6412,N_7371);
xnor U10682 (N_10682,N_2606,N_3348);
or U10683 (N_10683,N_1369,N_4709);
nand U10684 (N_10684,N_6161,N_3042);
nand U10685 (N_10685,N_969,N_1253);
nand U10686 (N_10686,N_5695,N_0);
or U10687 (N_10687,N_3652,N_6198);
nor U10688 (N_10688,N_1950,N_3789);
or U10689 (N_10689,N_8650,N_6327);
or U10690 (N_10690,N_6252,N_1808);
nand U10691 (N_10691,N_9565,N_3545);
and U10692 (N_10692,N_1246,N_9524);
or U10693 (N_10693,N_2676,N_6971);
and U10694 (N_10694,N_4211,N_429);
nor U10695 (N_10695,N_6647,N_2434);
nor U10696 (N_10696,N_3622,N_3794);
nor U10697 (N_10697,N_6858,N_9422);
or U10698 (N_10698,N_4712,N_4245);
nor U10699 (N_10699,N_5047,N_7401);
or U10700 (N_10700,N_2733,N_8474);
and U10701 (N_10701,N_6841,N_1872);
xor U10702 (N_10702,N_3071,N_735);
xnor U10703 (N_10703,N_9769,N_8199);
nor U10704 (N_10704,N_8794,N_5146);
nor U10705 (N_10705,N_1070,N_8208);
and U10706 (N_10706,N_1994,N_5115);
nor U10707 (N_10707,N_4095,N_3728);
or U10708 (N_10708,N_4725,N_6562);
or U10709 (N_10709,N_2131,N_648);
xnor U10710 (N_10710,N_9085,N_444);
nor U10711 (N_10711,N_1631,N_3487);
nor U10712 (N_10712,N_3770,N_7189);
nor U10713 (N_10713,N_347,N_355);
xnor U10714 (N_10714,N_6103,N_9275);
nand U10715 (N_10715,N_9501,N_5126);
or U10716 (N_10716,N_4544,N_3676);
or U10717 (N_10717,N_7421,N_5737);
or U10718 (N_10718,N_1358,N_2643);
nor U10719 (N_10719,N_2209,N_810);
and U10720 (N_10720,N_6172,N_8761);
nand U10721 (N_10721,N_8425,N_9150);
and U10722 (N_10722,N_5301,N_1530);
and U10723 (N_10723,N_1389,N_5659);
nand U10724 (N_10724,N_7212,N_5190);
nor U10725 (N_10725,N_2821,N_7204);
nor U10726 (N_10726,N_4158,N_3124);
xor U10727 (N_10727,N_5486,N_9226);
xnor U10728 (N_10728,N_3078,N_7884);
nor U10729 (N_10729,N_7455,N_4997);
xnor U10730 (N_10730,N_5617,N_6090);
nor U10731 (N_10731,N_9998,N_4248);
and U10732 (N_10732,N_1091,N_6136);
and U10733 (N_10733,N_2846,N_8345);
nand U10734 (N_10734,N_3340,N_2292);
or U10735 (N_10735,N_2862,N_7175);
nor U10736 (N_10736,N_9231,N_8389);
nand U10737 (N_10737,N_1661,N_7245);
nand U10738 (N_10738,N_4827,N_5709);
nor U10739 (N_10739,N_4774,N_7488);
nor U10740 (N_10740,N_5681,N_6747);
nor U10741 (N_10741,N_4631,N_2172);
nand U10742 (N_10742,N_6331,N_5330);
and U10743 (N_10743,N_7396,N_5942);
nor U10744 (N_10744,N_1041,N_5321);
nor U10745 (N_10745,N_1209,N_3250);
and U10746 (N_10746,N_3037,N_3547);
and U10747 (N_10747,N_1299,N_2094);
xor U10748 (N_10748,N_2853,N_2639);
and U10749 (N_10749,N_9055,N_4624);
or U10750 (N_10750,N_947,N_4693);
or U10751 (N_10751,N_2138,N_6347);
or U10752 (N_10752,N_3005,N_3859);
or U10753 (N_10753,N_2097,N_5761);
and U10754 (N_10754,N_6655,N_3360);
nor U10755 (N_10755,N_4856,N_2102);
nor U10756 (N_10756,N_7627,N_6257);
and U10757 (N_10757,N_6499,N_6351);
nand U10758 (N_10758,N_6165,N_1729);
and U10759 (N_10759,N_3569,N_8017);
nand U10760 (N_10760,N_7749,N_7293);
xor U10761 (N_10761,N_6274,N_9420);
nand U10762 (N_10762,N_9522,N_3690);
xnor U10763 (N_10763,N_1496,N_8631);
xnor U10764 (N_10764,N_6771,N_7096);
and U10765 (N_10765,N_5603,N_7693);
xnor U10766 (N_10766,N_9087,N_7586);
nand U10767 (N_10767,N_1295,N_5056);
nor U10768 (N_10768,N_9217,N_8149);
and U10769 (N_10769,N_4597,N_5530);
xor U10770 (N_10770,N_9105,N_4587);
xnor U10771 (N_10771,N_2754,N_1552);
and U10772 (N_10772,N_6114,N_6705);
xnor U10773 (N_10773,N_8188,N_4505);
nand U10774 (N_10774,N_5149,N_4640);
nor U10775 (N_10775,N_3371,N_7176);
or U10776 (N_10776,N_5223,N_7026);
nand U10777 (N_10777,N_4550,N_7523);
and U10778 (N_10778,N_4153,N_5703);
nor U10779 (N_10779,N_9140,N_3814);
xor U10780 (N_10780,N_1109,N_4572);
nor U10781 (N_10781,N_687,N_5013);
and U10782 (N_10782,N_9042,N_7644);
nand U10783 (N_10783,N_6700,N_4376);
xnor U10784 (N_10784,N_2501,N_2737);
xnor U10785 (N_10785,N_6791,N_7526);
xor U10786 (N_10786,N_6741,N_5019);
nand U10787 (N_10787,N_1405,N_9068);
nand U10788 (N_10788,N_3123,N_49);
nand U10789 (N_10789,N_8608,N_3784);
nand U10790 (N_10790,N_5630,N_38);
xnor U10791 (N_10791,N_4675,N_4724);
xor U10792 (N_10792,N_1776,N_4872);
nand U10793 (N_10793,N_3684,N_531);
and U10794 (N_10794,N_9430,N_5791);
nor U10795 (N_10795,N_7988,N_1761);
nand U10796 (N_10796,N_875,N_5453);
or U10797 (N_10797,N_4084,N_9532);
xnor U10798 (N_10798,N_2377,N_9191);
and U10799 (N_10799,N_2473,N_9552);
or U10800 (N_10800,N_3324,N_6583);
nor U10801 (N_10801,N_7755,N_6315);
and U10802 (N_10802,N_7249,N_5198);
nor U10803 (N_10803,N_624,N_1167);
nand U10804 (N_10804,N_9223,N_4282);
and U10805 (N_10805,N_5484,N_6901);
nor U10806 (N_10806,N_2067,N_5411);
nand U10807 (N_10807,N_1688,N_8502);
nand U10808 (N_10808,N_9757,N_5944);
xnor U10809 (N_10809,N_2869,N_7528);
xor U10810 (N_10810,N_8997,N_9828);
or U10811 (N_10811,N_794,N_785);
or U10812 (N_10812,N_1491,N_2201);
xor U10813 (N_10813,N_6627,N_6693);
and U10814 (N_10814,N_1898,N_2632);
nor U10815 (N_10815,N_7187,N_7056);
xnor U10816 (N_10816,N_7808,N_5153);
nor U10817 (N_10817,N_1889,N_8977);
nand U10818 (N_10818,N_4596,N_2362);
nor U10819 (N_10819,N_7108,N_4265);
xor U10820 (N_10820,N_9292,N_9600);
or U10821 (N_10821,N_8800,N_4428);
and U10822 (N_10822,N_6959,N_8439);
and U10823 (N_10823,N_6260,N_2115);
or U10824 (N_10824,N_9444,N_3863);
and U10825 (N_10825,N_5434,N_7405);
nand U10826 (N_10826,N_797,N_1191);
nor U10827 (N_10827,N_7826,N_6558);
xnor U10828 (N_10828,N_2319,N_3329);
nand U10829 (N_10829,N_6405,N_1460);
or U10830 (N_10830,N_4041,N_2969);
nor U10831 (N_10831,N_4116,N_4228);
or U10832 (N_10832,N_623,N_9028);
nor U10833 (N_10833,N_2614,N_6691);
and U10834 (N_10834,N_4090,N_4500);
xor U10835 (N_10835,N_8654,N_8173);
or U10836 (N_10836,N_3319,N_3185);
or U10837 (N_10837,N_683,N_8600);
nand U10838 (N_10838,N_6003,N_2724);
xnor U10839 (N_10839,N_9644,N_7784);
nor U10840 (N_10840,N_7490,N_2029);
or U10841 (N_10841,N_5863,N_3449);
or U10842 (N_10842,N_3128,N_2351);
xor U10843 (N_10843,N_1581,N_2585);
nand U10844 (N_10844,N_9357,N_8963);
or U10845 (N_10845,N_9946,N_6837);
or U10846 (N_10846,N_3893,N_5937);
xor U10847 (N_10847,N_6989,N_7307);
and U10848 (N_10848,N_706,N_7790);
and U10849 (N_10849,N_9003,N_3356);
or U10850 (N_10850,N_9933,N_596);
nand U10851 (N_10851,N_5722,N_2384);
and U10852 (N_10852,N_3940,N_5576);
nand U10853 (N_10853,N_5209,N_3297);
nor U10854 (N_10854,N_8809,N_8323);
xnor U10855 (N_10855,N_2032,N_6552);
and U10856 (N_10856,N_9928,N_462);
or U10857 (N_10857,N_1048,N_2407);
and U10858 (N_10858,N_3758,N_2570);
and U10859 (N_10859,N_6995,N_3933);
xnor U10860 (N_10860,N_5973,N_3179);
nor U10861 (N_10861,N_4371,N_8909);
xor U10862 (N_10862,N_8991,N_4889);
or U10863 (N_10863,N_1376,N_6856);
nand U10864 (N_10864,N_4935,N_4131);
or U10865 (N_10865,N_876,N_9910);
nand U10866 (N_10866,N_4309,N_7304);
nor U10867 (N_10867,N_8123,N_1292);
and U10868 (N_10868,N_1683,N_9145);
xnor U10869 (N_10869,N_9074,N_6132);
and U10870 (N_10870,N_7333,N_9113);
xor U10871 (N_10871,N_5268,N_5349);
and U10872 (N_10872,N_4912,N_3514);
or U10873 (N_10873,N_4017,N_4880);
nand U10874 (N_10874,N_828,N_448);
and U10875 (N_10875,N_1180,N_6927);
nand U10876 (N_10876,N_1881,N_2510);
or U10877 (N_10877,N_2566,N_2661);
or U10878 (N_10878,N_1813,N_4957);
nand U10879 (N_10879,N_8748,N_5927);
xnor U10880 (N_10880,N_532,N_4481);
and U10881 (N_10881,N_39,N_7186);
or U10882 (N_10882,N_8490,N_141);
or U10883 (N_10883,N_8005,N_1074);
nor U10884 (N_10884,N_9750,N_2656);
nor U10885 (N_10885,N_2318,N_2666);
and U10886 (N_10886,N_1829,N_7305);
nand U10887 (N_10887,N_4699,N_3720);
xnor U10888 (N_10888,N_1084,N_5097);
xor U10889 (N_10889,N_8359,N_5195);
and U10890 (N_10890,N_5692,N_6204);
and U10891 (N_10891,N_6982,N_1480);
xnor U10892 (N_10892,N_720,N_8219);
nand U10893 (N_10893,N_9728,N_5231);
nor U10894 (N_10894,N_9459,N_9347);
nand U10895 (N_10895,N_5202,N_818);
nor U10896 (N_10896,N_139,N_4137);
or U10897 (N_10897,N_4813,N_3680);
or U10898 (N_10898,N_9890,N_6026);
or U10899 (N_10899,N_7009,N_533);
or U10900 (N_10900,N_5386,N_9579);
nor U10901 (N_10901,N_2149,N_7329);
or U10902 (N_10902,N_5378,N_4283);
and U10903 (N_10903,N_1557,N_3050);
xor U10904 (N_10904,N_2269,N_3303);
nor U10905 (N_10905,N_7828,N_4610);
xnor U10906 (N_10906,N_5770,N_7655);
and U10907 (N_10907,N_7576,N_3096);
and U10908 (N_10908,N_4642,N_1510);
nand U10909 (N_10909,N_1086,N_5438);
nand U10910 (N_10910,N_1935,N_6464);
nor U10911 (N_10911,N_3581,N_9377);
nand U10912 (N_10912,N_3640,N_2305);
and U10913 (N_10913,N_1137,N_6156);
xnor U10914 (N_10914,N_1633,N_404);
nor U10915 (N_10915,N_2966,N_6711);
or U10916 (N_10916,N_8402,N_412);
or U10917 (N_10917,N_2890,N_2841);
xnor U10918 (N_10918,N_9023,N_8526);
xnor U10919 (N_10919,N_7106,N_8603);
nand U10920 (N_10920,N_1924,N_4253);
nor U10921 (N_10921,N_6077,N_8832);
nand U10922 (N_10922,N_2865,N_8379);
or U10923 (N_10923,N_5350,N_1986);
and U10924 (N_10924,N_899,N_2081);
xnor U10925 (N_10925,N_8214,N_4438);
or U10926 (N_10926,N_3452,N_5232);
xor U10927 (N_10927,N_6584,N_6602);
or U10928 (N_10928,N_160,N_8829);
nand U10929 (N_10929,N_6167,N_3493);
nand U10930 (N_10930,N_9536,N_9556);
and U10931 (N_10931,N_5654,N_207);
and U10932 (N_10932,N_3434,N_5263);
xor U10933 (N_10933,N_5723,N_1249);
and U10934 (N_10934,N_1529,N_1947);
nor U10935 (N_10935,N_4535,N_9354);
xnor U10936 (N_10936,N_6610,N_7043);
or U10937 (N_10937,N_439,N_3805);
nand U10938 (N_10938,N_8979,N_9471);
xnor U10939 (N_10939,N_1293,N_3825);
xor U10940 (N_10940,N_6251,N_9396);
xor U10941 (N_10941,N_3724,N_2849);
and U10942 (N_10942,N_9530,N_2578);
nand U10943 (N_10943,N_4257,N_4755);
nand U10944 (N_10944,N_3167,N_686);
and U10945 (N_10945,N_9251,N_7657);
nand U10946 (N_10946,N_3072,N_5675);
or U10947 (N_10947,N_2525,N_3089);
nand U10948 (N_10948,N_4832,N_672);
and U10949 (N_10949,N_8659,N_1866);
nor U10950 (N_10950,N_8792,N_1788);
or U10951 (N_10951,N_6579,N_3620);
nand U10952 (N_10952,N_3506,N_275);
and U10953 (N_10953,N_5090,N_9791);
nand U10954 (N_10954,N_6565,N_2648);
nand U10955 (N_10955,N_3336,N_9486);
nor U10956 (N_10956,N_1651,N_2805);
and U10957 (N_10957,N_958,N_3014);
xor U10958 (N_10958,N_4571,N_5731);
xnor U10959 (N_10959,N_9210,N_3165);
and U10960 (N_10960,N_467,N_8826);
and U10961 (N_10961,N_6634,N_5211);
or U10962 (N_10962,N_6460,N_7977);
and U10963 (N_10963,N_1133,N_1172);
xnor U10964 (N_10964,N_7344,N_1190);
xnor U10965 (N_10965,N_5933,N_5747);
or U10966 (N_10966,N_8318,N_8355);
and U10967 (N_10967,N_6488,N_90);
or U10968 (N_10968,N_1647,N_3754);
xor U10969 (N_10969,N_3800,N_6231);
or U10970 (N_10970,N_232,N_5663);
or U10971 (N_10971,N_7726,N_1983);
nand U10972 (N_10972,N_9342,N_5825);
nand U10973 (N_10973,N_979,N_7423);
or U10974 (N_10974,N_7225,N_755);
xor U10975 (N_10975,N_849,N_5187);
nand U10976 (N_10976,N_4288,N_8120);
nand U10977 (N_10977,N_4539,N_3561);
nand U10978 (N_10978,N_5456,N_6038);
and U10979 (N_10979,N_7769,N_4187);
xor U10980 (N_10980,N_4230,N_5809);
or U10981 (N_10981,N_7050,N_5045);
nand U10982 (N_10982,N_7795,N_240);
xnor U10983 (N_10983,N_7127,N_167);
xnor U10984 (N_10984,N_8838,N_7313);
or U10985 (N_10985,N_5105,N_2694);
and U10986 (N_10986,N_6273,N_7807);
and U10987 (N_10987,N_7758,N_4547);
nor U10988 (N_10988,N_8987,N_606);
nand U10989 (N_10989,N_5935,N_6194);
or U10990 (N_10990,N_4144,N_6508);
xnor U10991 (N_10991,N_841,N_3266);
nor U10992 (N_10992,N_3616,N_7550);
nand U10993 (N_10993,N_2255,N_7811);
xor U10994 (N_10994,N_6807,N_492);
xnor U10995 (N_10995,N_1996,N_4147);
xor U10996 (N_10996,N_6416,N_4762);
or U10997 (N_10997,N_3518,N_5542);
and U10998 (N_10998,N_4632,N_7860);
nor U10999 (N_10999,N_932,N_1826);
nor U11000 (N_11000,N_547,N_55);
nand U11001 (N_11001,N_6980,N_1397);
or U11002 (N_11002,N_8159,N_7781);
or U11003 (N_11003,N_9609,N_1740);
or U11004 (N_11004,N_1725,N_6943);
and U11005 (N_11005,N_3653,N_5384);
nand U11006 (N_11006,N_3289,N_6002);
xor U11007 (N_11007,N_9262,N_9958);
and U11008 (N_11008,N_8072,N_8568);
or U11009 (N_11009,N_9197,N_1509);
nor U11010 (N_11010,N_7019,N_1433);
nand U11011 (N_11011,N_8265,N_9647);
and U11012 (N_11012,N_688,N_1878);
and U11013 (N_11013,N_9627,N_1559);
and U11014 (N_11014,N_7575,N_4306);
nand U11015 (N_11015,N_9097,N_4679);
nor U11016 (N_11016,N_3936,N_7651);
xor U11017 (N_11017,N_2642,N_19);
or U11018 (N_11018,N_5443,N_4512);
nor U11019 (N_11019,N_696,N_4781);
nor U11020 (N_11020,N_9252,N_3646);
nor U11021 (N_11021,N_1913,N_7420);
or U11022 (N_11022,N_8039,N_8471);
nor U11023 (N_11023,N_2745,N_4648);
nor U11024 (N_11024,N_8754,N_1367);
nor U11025 (N_11025,N_3350,N_4336);
and U11026 (N_11026,N_1911,N_2924);
nand U11027 (N_11027,N_709,N_4456);
nor U11028 (N_11028,N_3252,N_6928);
nor U11029 (N_11029,N_457,N_7094);
nand U11030 (N_11030,N_827,N_566);
nand U11031 (N_11031,N_248,N_5852);
or U11032 (N_11032,N_2677,N_6671);
xnor U11033 (N_11033,N_2732,N_459);
or U11034 (N_11034,N_5304,N_5945);
and U11035 (N_11035,N_1068,N_2323);
xor U11036 (N_11036,N_2581,N_6595);
xor U11037 (N_11037,N_9861,N_3883);
or U11038 (N_11038,N_8189,N_5575);
and U11039 (N_11039,N_4325,N_7076);
xnor U11040 (N_11040,N_3550,N_2736);
or U11041 (N_11041,N_6125,N_8856);
and U11042 (N_11042,N_7341,N_5029);
and U11043 (N_11043,N_210,N_3649);
and U11044 (N_11044,N_8672,N_4242);
xnor U11045 (N_11045,N_6964,N_425);
and U11046 (N_11046,N_4159,N_3315);
and U11047 (N_11047,N_2644,N_6628);
nor U11048 (N_11048,N_3203,N_8553);
nand U11049 (N_11049,N_3527,N_1251);
or U11050 (N_11050,N_3261,N_5743);
and U11051 (N_11051,N_8886,N_9514);
nand U11052 (N_11052,N_2959,N_1149);
xnor U11053 (N_11053,N_5896,N_2940);
or U11054 (N_11054,N_1964,N_2329);
xor U11055 (N_11055,N_637,N_2345);
xor U11056 (N_11056,N_2126,N_443);
or U11057 (N_11057,N_2476,N_3074);
nor U11058 (N_11058,N_8435,N_5283);
nand U11059 (N_11059,N_8967,N_8460);
and U11060 (N_11060,N_1735,N_8903);
nor U11061 (N_11061,N_2381,N_7814);
or U11062 (N_11062,N_6728,N_7254);
or U11063 (N_11063,N_8543,N_9499);
and U11064 (N_11064,N_6570,N_8089);
xor U11065 (N_11065,N_6006,N_7016);
nand U11066 (N_11066,N_5792,N_1401);
xor U11067 (N_11067,N_273,N_4662);
nand U11068 (N_11068,N_7444,N_2547);
nand U11069 (N_11069,N_99,N_819);
and U11070 (N_11070,N_3821,N_3641);
and U11071 (N_11071,N_9694,N_8284);
xnor U11072 (N_11072,N_6119,N_8091);
xnor U11073 (N_11073,N_6321,N_9186);
nand U11074 (N_11074,N_5420,N_3575);
xnor U11075 (N_11075,N_5974,N_7146);
nand U11076 (N_11076,N_4365,N_9727);
nor U11077 (N_11077,N_9982,N_3398);
nand U11078 (N_11078,N_9358,N_29);
xnor U11079 (N_11079,N_8844,N_8445);
and U11080 (N_11080,N_1547,N_5110);
xnor U11081 (N_11081,N_8112,N_6772);
nand U11082 (N_11082,N_2231,N_864);
nand U11083 (N_11083,N_4528,N_1979);
nand U11084 (N_11084,N_1236,N_1604);
nand U11085 (N_11085,N_2271,N_3213);
xor U11086 (N_11086,N_4388,N_6484);
and U11087 (N_11087,N_1585,N_5317);
and U11088 (N_11088,N_8995,N_1952);
nand U11089 (N_11089,N_3993,N_9587);
or U11090 (N_11090,N_9132,N_9364);
or U11091 (N_11091,N_5008,N_7241);
xor U11092 (N_11092,N_3911,N_6918);
xor U11093 (N_11093,N_1119,N_584);
or U11094 (N_11094,N_6740,N_853);
and U11095 (N_11095,N_1361,N_9193);
nor U11096 (N_11096,N_7560,N_2253);
nor U11097 (N_11097,N_9294,N_7636);
or U11098 (N_11098,N_6623,N_233);
or U11099 (N_11099,N_3648,N_7650);
and U11100 (N_11100,N_4639,N_8119);
and U11101 (N_11101,N_6752,N_411);
and U11102 (N_11102,N_4471,N_2383);
xor U11103 (N_11103,N_8812,N_2560);
or U11104 (N_11104,N_9847,N_669);
or U11105 (N_11105,N_1618,N_2452);
and U11106 (N_11106,N_6042,N_3194);
nor U11107 (N_11107,N_4497,N_7785);
xor U11108 (N_11108,N_44,N_4241);
and U11109 (N_11109,N_4674,N_5869);
nor U11110 (N_11110,N_9142,N_5981);
nand U11111 (N_11111,N_6413,N_8504);
and U11112 (N_11112,N_2222,N_570);
or U11113 (N_11113,N_6256,N_9837);
nand U11114 (N_11114,N_2015,N_2621);
xnor U11115 (N_11115,N_4142,N_3548);
and U11116 (N_11116,N_1927,N_8663);
or U11117 (N_11117,N_4896,N_8361);
nor U11118 (N_11118,N_1211,N_7219);
xnor U11119 (N_11119,N_6432,N_9082);
and U11120 (N_11120,N_261,N_1690);
nand U11121 (N_11121,N_8272,N_5893);
xor U11122 (N_11122,N_6775,N_1806);
nand U11123 (N_11123,N_2859,N_8836);
or U11124 (N_11124,N_9683,N_9980);
xnor U11125 (N_11125,N_8289,N_509);
xor U11126 (N_11126,N_510,N_1884);
and U11127 (N_11127,N_5522,N_3583);
xnor U11128 (N_11128,N_9382,N_8493);
xnor U11129 (N_11129,N_2371,N_5952);
and U11130 (N_11130,N_4990,N_2932);
nor U11131 (N_11131,N_5788,N_7696);
nor U11132 (N_11132,N_521,N_9072);
or U11133 (N_11133,N_4204,N_2688);
nor U11134 (N_11134,N_1644,N_4688);
nand U11135 (N_11135,N_6236,N_9513);
nor U11136 (N_11136,N_7534,N_8700);
and U11137 (N_11137,N_1406,N_8316);
xnor U11138 (N_11138,N_1235,N_445);
or U11139 (N_11139,N_366,N_8060);
or U11140 (N_11140,N_4006,N_1329);
nor U11141 (N_11141,N_121,N_3855);
and U11142 (N_11142,N_3334,N_8462);
nand U11143 (N_11143,N_9213,N_3976);
or U11144 (N_11144,N_6985,N_463);
nor U11145 (N_11145,N_469,N_5189);
nand U11146 (N_11146,N_8229,N_2124);
and U11147 (N_11147,N_5697,N_9051);
xnor U11148 (N_11148,N_8622,N_9538);
or U11149 (N_11149,N_8833,N_4819);
nand U11150 (N_11150,N_5329,N_5151);
nand U11151 (N_11151,N_6665,N_122);
nand U11152 (N_11152,N_4021,N_3619);
nand U11153 (N_11153,N_8197,N_3793);
and U11154 (N_11154,N_7008,N_8254);
nand U11155 (N_11155,N_4409,N_382);
xnor U11156 (N_11156,N_8931,N_3407);
and U11157 (N_11157,N_1303,N_1394);
nand U11158 (N_11158,N_8339,N_2134);
nor U11159 (N_11159,N_4765,N_9620);
xor U11160 (N_11160,N_4551,N_3984);
and U11161 (N_11161,N_9474,N_7590);
xnor U11162 (N_11162,N_5137,N_6467);
nor U11163 (N_11163,N_2703,N_8459);
nor U11164 (N_11164,N_3973,N_1959);
nor U11165 (N_11165,N_2856,N_5017);
nand U11166 (N_11166,N_8684,N_3909);
nor U11167 (N_11167,N_2360,N_4064);
or U11168 (N_11168,N_4739,N_2897);
nand U11169 (N_11169,N_4635,N_8724);
xor U11170 (N_11170,N_6731,N_7686);
xor U11171 (N_11171,N_6336,N_7543);
nor U11172 (N_11172,N_5514,N_3039);
xnor U11173 (N_11173,N_5950,N_3624);
xnor U11174 (N_11174,N_1116,N_7976);
xnor U11175 (N_11175,N_1247,N_2752);
and U11176 (N_11176,N_4341,N_3842);
and U11177 (N_11177,N_5372,N_9293);
xnor U11178 (N_11178,N_8649,N_9751);
and U11179 (N_11179,N_6075,N_786);
and U11180 (N_11180,N_1243,N_5688);
nor U11181 (N_11181,N_2423,N_7699);
or U11182 (N_11182,N_2313,N_4121);
and U11183 (N_11183,N_1430,N_7315);
and U11184 (N_11184,N_5095,N_3955);
or U11185 (N_11185,N_6779,N_5286);
nand U11186 (N_11186,N_9535,N_9822);
xnor U11187 (N_11187,N_173,N_3711);
or U11188 (N_11188,N_2403,N_989);
or U11189 (N_11189,N_8884,N_6091);
and U11190 (N_11190,N_1859,N_6365);
xnor U11191 (N_11191,N_1702,N_1304);
nor U11192 (N_11192,N_7774,N_263);
and U11193 (N_11193,N_5691,N_578);
or U11194 (N_11194,N_1669,N_1543);
xor U11195 (N_11195,N_8636,N_3900);
xnor U11196 (N_11196,N_3757,N_4395);
nand U11197 (N_11197,N_1404,N_8420);
and U11198 (N_11198,N_6953,N_5834);
and U11199 (N_11199,N_390,N_7182);
xor U11200 (N_11200,N_8406,N_3919);
nor U11201 (N_11201,N_2511,N_4316);
or U11202 (N_11202,N_1580,N_1507);
or U11203 (N_11203,N_3788,N_6229);
and U11204 (N_11204,N_8340,N_339);
nor U11205 (N_11205,N_9160,N_1733);
or U11206 (N_11206,N_4450,N_6095);
nor U11207 (N_11207,N_4802,N_7621);
or U11208 (N_11208,N_5241,N_2478);
nand U11209 (N_11209,N_2698,N_8058);
or U11210 (N_11210,N_5355,N_434);
and U11211 (N_11211,N_3174,N_7568);
nor U11212 (N_11212,N_4118,N_473);
and U11213 (N_11213,N_2592,N_475);
nor U11214 (N_11214,N_582,N_229);
and U11215 (N_11215,N_1963,N_8185);
nor U11216 (N_11216,N_7105,N_6688);
or U11217 (N_11217,N_1544,N_6019);
nand U11218 (N_11218,N_5555,N_7873);
and U11219 (N_11219,N_8064,N_3692);
nand U11220 (N_11220,N_3216,N_2574);
or U11221 (N_11221,N_3740,N_7002);
or U11222 (N_11222,N_307,N_2972);
and U11223 (N_11223,N_8311,N_2599);
and U11224 (N_11224,N_1938,N_369);
nand U11225 (N_11225,N_6767,N_9176);
and U11226 (N_11226,N_5780,N_3876);
nor U11227 (N_11227,N_9123,N_9709);
or U11228 (N_11228,N_9881,N_8904);
nand U11229 (N_11229,N_1413,N_2087);
or U11230 (N_11230,N_6492,N_146);
nand U11231 (N_11231,N_5500,N_4845);
nand U11232 (N_11232,N_6170,N_9766);
nor U11233 (N_11233,N_5795,N_8889);
and U11234 (N_11234,N_1519,N_4846);
nand U11235 (N_11235,N_9655,N_5701);
xor U11236 (N_11236,N_5922,N_7629);
or U11237 (N_11237,N_1063,N_1489);
and U11238 (N_11238,N_7812,N_8855);
nand U11239 (N_11239,N_4660,N_5064);
or U11240 (N_11240,N_6677,N_9012);
nand U11241 (N_11241,N_3119,N_4231);
or U11242 (N_11242,N_588,N_1392);
nand U11243 (N_11243,N_3953,N_1809);
nor U11244 (N_11244,N_7713,N_9199);
xor U11245 (N_11245,N_1024,N_9991);
and U11246 (N_11246,N_5871,N_659);
or U11247 (N_11247,N_6596,N_7593);
nand U11248 (N_11248,N_360,N_1711);
nor U11249 (N_11249,N_8006,N_8117);
xor U11250 (N_11250,N_7637,N_3592);
or U11251 (N_11251,N_6604,N_3891);
nand U11252 (N_11252,N_3286,N_1803);
xnor U11253 (N_11253,N_9528,N_3666);
xnor U11254 (N_11254,N_5998,N_315);
or U11255 (N_11255,N_8473,N_592);
nand U11256 (N_11256,N_1495,N_420);
nand U11257 (N_11257,N_553,N_8153);
nor U11258 (N_11258,N_3439,N_8181);
and U11259 (N_11259,N_8211,N_5030);
and U11260 (N_11260,N_6438,N_1517);
xor U11261 (N_11261,N_195,N_2537);
and U11262 (N_11262,N_489,N_8438);
nand U11263 (N_11263,N_6059,N_7668);
and U11264 (N_11264,N_3746,N_2267);
and U11265 (N_11265,N_6290,N_8643);
nor U11266 (N_11266,N_9372,N_6744);
xnor U11267 (N_11267,N_4619,N_6462);
xor U11268 (N_11268,N_2401,N_1686);
nor U11269 (N_11269,N_1322,N_4295);
nor U11270 (N_11270,N_865,N_6799);
xnor U11271 (N_11271,N_2013,N_1239);
or U11272 (N_11272,N_572,N_2790);
or U11273 (N_11273,N_326,N_4457);
xor U11274 (N_11274,N_4938,N_9723);
xnor U11275 (N_11275,N_7708,N_6185);
nand U11276 (N_11276,N_7059,N_3051);
xor U11277 (N_11277,N_5902,N_9397);
nand U11278 (N_11278,N_4945,N_8525);
and U11279 (N_11279,N_8003,N_3786);
and U11280 (N_11280,N_941,N_9325);
nand U11281 (N_11281,N_2843,N_5673);
nand U11282 (N_11282,N_9061,N_7294);
nand U11283 (N_11283,N_6864,N_9219);
or U11284 (N_11284,N_3220,N_3473);
or U11285 (N_11285,N_9455,N_4732);
nor U11286 (N_11286,N_6282,N_8671);
nand U11287 (N_11287,N_3762,N_1468);
xor U11288 (N_11288,N_8015,N_4299);
or U11289 (N_11289,N_6929,N_7268);
nand U11290 (N_11290,N_5832,N_1822);
or U11291 (N_11291,N_4918,N_2781);
nor U11292 (N_11292,N_4462,N_6773);
nand U11293 (N_11293,N_6944,N_9797);
nand U11294 (N_11294,N_7321,N_4329);
xnor U11295 (N_11295,N_1910,N_1478);
and U11296 (N_11296,N_2468,N_882);
and U11297 (N_11297,N_3628,N_5727);
or U11298 (N_11298,N_2692,N_7399);
nand U11299 (N_11299,N_6309,N_7214);
nand U11300 (N_11300,N_9409,N_9330);
nor U11301 (N_11301,N_2395,N_9663);
xnor U11302 (N_11302,N_6443,N_7810);
and U11303 (N_11303,N_2770,N_8985);
and U11304 (N_11304,N_7919,N_9495);
or U11305 (N_11305,N_5371,N_3399);
nor U11306 (N_11306,N_9438,N_5265);
and U11307 (N_11307,N_7426,N_5846);
and U11308 (N_11308,N_4645,N_2155);
and U11309 (N_11309,N_9413,N_5309);
and U11310 (N_11310,N_8322,N_8312);
xor U11311 (N_11311,N_6941,N_2232);
and U11312 (N_11312,N_1681,N_93);
or U11313 (N_11313,N_5175,N_3989);
nand U11314 (N_11314,N_2424,N_5279);
nor U11315 (N_11315,N_1381,N_8588);
and U11316 (N_11316,N_3562,N_337);
nor U11317 (N_11317,N_8660,N_9798);
and U11318 (N_11318,N_4307,N_6249);
xnor U11319 (N_11319,N_8535,N_2565);
nor U11320 (N_11320,N_701,N_5102);
nor U11321 (N_11321,N_6846,N_9636);
nand U11322 (N_11322,N_652,N_8347);
xnor U11323 (N_11323,N_9510,N_4154);
and U11324 (N_11324,N_8973,N_8755);
xor U11325 (N_11325,N_3914,N_476);
or U11326 (N_11326,N_6689,N_4485);
or U11327 (N_11327,N_6278,N_6872);
or U11328 (N_11328,N_5327,N_8550);
nor U11329 (N_11329,N_573,N_2926);
xnor U11330 (N_11330,N_4297,N_3245);
nand U11331 (N_11331,N_1129,N_8956);
or U11332 (N_11332,N_8615,N_7289);
and U11333 (N_11333,N_8770,N_7555);
and U11334 (N_11334,N_9255,N_6183);
nor U11335 (N_11335,N_9862,N_2288);
and U11336 (N_11336,N_4742,N_1443);
nor U11337 (N_11337,N_4298,N_7078);
nand U11338 (N_11338,N_6806,N_86);
nand U11339 (N_11339,N_4858,N_1380);
or U11340 (N_11340,N_6280,N_6495);
nand U11341 (N_11341,N_5507,N_7498);
or U11342 (N_11342,N_3437,N_730);
nor U11343 (N_11343,N_8090,N_2545);
xnor U11344 (N_11344,N_5539,N_4749);
and U11345 (N_11345,N_9216,N_7181);
xnor U11346 (N_11346,N_4421,N_7943);
and U11347 (N_11347,N_8470,N_7723);
and U11348 (N_11348,N_8696,N_488);
or U11349 (N_11349,N_9859,N_4854);
or U11350 (N_11350,N_3896,N_197);
nor U11351 (N_11351,N_7027,N_2421);
or U11352 (N_11352,N_5436,N_7751);
xor U11353 (N_11353,N_7616,N_2507);
or U11354 (N_11354,N_5282,N_5036);
nor U11355 (N_11355,N_9973,N_7510);
xor U11356 (N_11356,N_1570,N_7478);
xnor U11357 (N_11357,N_4098,N_7508);
nor U11358 (N_11358,N_6832,N_7397);
and U11359 (N_11359,N_6900,N_4135);
nand U11360 (N_11360,N_2474,N_452);
nor U11361 (N_11361,N_6965,N_4343);
nor U11362 (N_11362,N_607,N_9786);
xnor U11363 (N_11363,N_7416,N_8109);
nor U11364 (N_11364,N_998,N_3586);
xor U11365 (N_11365,N_4611,N_1588);
xnor U11366 (N_11366,N_809,N_2405);
or U11367 (N_11367,N_5934,N_773);
and U11368 (N_11368,N_5885,N_3342);
nand U11369 (N_11369,N_662,N_2341);
xnor U11370 (N_11370,N_2300,N_9911);
xnor U11371 (N_11371,N_1800,N_4863);
or U11372 (N_11372,N_2325,N_5125);
or U11373 (N_11373,N_7373,N_5580);
and U11374 (N_11374,N_1638,N_7981);
xnor U11375 (N_11375,N_5811,N_4127);
xor U11376 (N_11376,N_7126,N_9695);
xnor U11377 (N_11377,N_9225,N_8287);
and U11378 (N_11378,N_9260,N_5171);
and U11379 (N_11379,N_6138,N_6826);
or U11380 (N_11380,N_8487,N_5621);
and U11381 (N_11381,N_8303,N_2775);
xnor U11382 (N_11382,N_3870,N_1606);
nor U11383 (N_11383,N_6874,N_9990);
and U11384 (N_11384,N_7438,N_9490);
nand U11385 (N_11385,N_832,N_8503);
nor U11386 (N_11386,N_3858,N_527);
nand U11387 (N_11387,N_4713,N_71);
or U11388 (N_11388,N_2159,N_3946);
nand U11389 (N_11389,N_6726,N_7184);
nand U11390 (N_11390,N_7905,N_188);
xor U11391 (N_11391,N_9697,N_5622);
xor U11392 (N_11392,N_2937,N_1987);
nand U11393 (N_11393,N_3918,N_4564);
nand U11394 (N_11394,N_6190,N_8798);
nor U11395 (N_11395,N_5774,N_4433);
and U11396 (N_11396,N_6459,N_6303);
xor U11397 (N_11397,N_1799,N_5797);
or U11398 (N_11398,N_9316,N_3092);
or U11399 (N_11399,N_3571,N_3675);
xnor U11400 (N_11400,N_1044,N_4074);
or U11401 (N_11401,N_4419,N_3705);
xnor U11402 (N_11402,N_2340,N_545);
nand U11403 (N_11403,N_634,N_7960);
nor U11404 (N_11404,N_6803,N_8317);
or U11405 (N_11405,N_5142,N_5052);
xor U11406 (N_11406,N_8847,N_7918);
and U11407 (N_11407,N_6533,N_2726);
or U11408 (N_11408,N_6580,N_3714);
nor U11409 (N_11409,N_9717,N_5730);
nand U11410 (N_11410,N_3535,N_6560);
and U11411 (N_11411,N_42,N_6168);
and U11412 (N_11412,N_5845,N_5033);
nor U11413 (N_11413,N_5242,N_9398);
and U11414 (N_11414,N_4578,N_8440);
and U11415 (N_11415,N_4928,N_4871);
nor U11416 (N_11416,N_6476,N_2375);
and U11417 (N_11417,N_4616,N_3264);
or U11418 (N_11418,N_8871,N_7933);
nor U11419 (N_11419,N_1050,N_1120);
or U11420 (N_11420,N_5754,N_763);
nand U11421 (N_11421,N_8467,N_220);
nand U11422 (N_11422,N_679,N_3196);
nand U11423 (N_11423,N_2691,N_5599);
nor U11424 (N_11424,N_6239,N_35);
and U11425 (N_11425,N_3963,N_5597);
and U11426 (N_11426,N_1511,N_6620);
xor U11427 (N_11427,N_8733,N_6061);
nor U11428 (N_11428,N_3450,N_4035);
nand U11429 (N_11429,N_483,N_9283);
nor U11430 (N_11430,N_6758,N_1075);
or U11431 (N_11431,N_5357,N_5907);
nor U11432 (N_11432,N_4831,N_5298);
nor U11433 (N_11433,N_1372,N_1623);
or U11434 (N_11434,N_1710,N_5579);
nor U11435 (N_11435,N_6253,N_9220);
nor U11436 (N_11436,N_496,N_8356);
or U11437 (N_11437,N_1513,N_7419);
or U11438 (N_11438,N_5118,N_7162);
nor U11439 (N_11439,N_8585,N_9116);
and U11440 (N_11440,N_8492,N_364);
nand U11441 (N_11441,N_6563,N_8592);
nor U11442 (N_11442,N_4416,N_2872);
nand U11443 (N_11443,N_6384,N_8062);
nand U11444 (N_11444,N_4012,N_4758);
or U11445 (N_11445,N_3693,N_6897);
nor U11446 (N_11446,N_8495,N_2719);
nand U11447 (N_11447,N_6483,N_3175);
xnor U11448 (N_11448,N_1780,N_8775);
and U11449 (N_11449,N_8780,N_7450);
nor U11450 (N_11450,N_9058,N_7403);
and U11451 (N_11451,N_6264,N_3219);
and U11452 (N_11452,N_4033,N_1785);
and U11453 (N_11453,N_7047,N_3647);
nand U11454 (N_11454,N_6108,N_2039);
nor U11455 (N_11455,N_216,N_8456);
nand U11456 (N_11456,N_2482,N_625);
and U11457 (N_11457,N_5227,N_7925);
and U11458 (N_11458,N_806,N_237);
nand U11459 (N_11459,N_9773,N_4961);
and U11460 (N_11460,N_3406,N_9386);
and U11461 (N_11461,N_7258,N_5668);
xor U11462 (N_11462,N_2077,N_2295);
xor U11463 (N_11463,N_2064,N_1815);
nand U11464 (N_11464,N_8273,N_6721);
xnor U11465 (N_11465,N_9414,N_8421);
or U11466 (N_11466,N_6302,N_7335);
and U11467 (N_11467,N_3772,N_4711);
xor U11468 (N_11468,N_8357,N_6883);
xor U11469 (N_11469,N_7979,N_3228);
xnor U11470 (N_11470,N_5504,N_1135);
or U11471 (N_11471,N_8351,N_6440);
nor U11472 (N_11472,N_1625,N_6394);
or U11473 (N_11473,N_3395,N_5048);
nand U11474 (N_11474,N_9963,N_6962);
nand U11475 (N_11475,N_8476,N_7057);
and U11476 (N_11476,N_7538,N_727);
or U11477 (N_11477,N_7633,N_9726);
xnor U11478 (N_11478,N_5717,N_7171);
or U11479 (N_11479,N_4073,N_8713);
xor U11480 (N_11480,N_1001,N_2105);
nor U11481 (N_11481,N_3307,N_3045);
nor U11482 (N_11482,N_8288,N_3538);
or U11483 (N_11483,N_6966,N_6809);
nor U11484 (N_11484,N_9037,N_2179);
nand U11485 (N_11485,N_7194,N_5991);
or U11486 (N_11486,N_1422,N_7610);
nor U11487 (N_11487,N_1705,N_1240);
and U11488 (N_11488,N_9480,N_5089);
nand U11489 (N_11489,N_2086,N_764);
nand U11490 (N_11490,N_8014,N_7144);
nor U11491 (N_11491,N_2158,N_7743);
and U11492 (N_11492,N_3222,N_6029);
xnor U11493 (N_11493,N_3288,N_2485);
xnor U11494 (N_11494,N_565,N_6154);
xnor U11495 (N_11495,N_7041,N_7612);
nand U11496 (N_11496,N_689,N_4860);
nor U11497 (N_11497,N_9120,N_2920);
nand U11498 (N_11498,N_8968,N_3346);
xnor U11499 (N_11499,N_7880,N_6538);
xor U11500 (N_11500,N_3774,N_3546);
nand U11501 (N_11501,N_1738,N_3262);
or U11502 (N_11502,N_1765,N_1668);
xnor U11503 (N_11503,N_3367,N_9473);
or U11504 (N_11504,N_665,N_2242);
nor U11505 (N_11505,N_7051,N_6357);
nand U11506 (N_11506,N_7638,N_2982);
nor U11507 (N_11507,N_2016,N_5497);
nor U11508 (N_11508,N_8539,N_4161);
xnor U11509 (N_11509,N_413,N_8374);
and U11510 (N_11510,N_9904,N_673);
and U11511 (N_11511,N_9994,N_4560);
xnor U11512 (N_11512,N_6178,N_9332);
or U11513 (N_11513,N_9440,N_4799);
nor U11514 (N_11514,N_3276,N_4562);
xor U11515 (N_11515,N_5405,N_9247);
nor U11516 (N_11516,N_6685,N_3553);
nor U11517 (N_11517,N_7157,N_1712);
nand U11518 (N_11518,N_3820,N_3837);
nor U11519 (N_11519,N_3373,N_9177);
and U11520 (N_11520,N_5070,N_3067);
nand U11521 (N_11521,N_9738,N_6694);
or U11522 (N_11522,N_2480,N_6453);
nand U11523 (N_11523,N_3066,N_833);
and U11524 (N_11524,N_309,N_9290);
nor U11525 (N_11525,N_8424,N_5260);
and U11526 (N_11526,N_6366,N_7384);
and U11527 (N_11527,N_9253,N_2055);
or U11528 (N_11528,N_3485,N_8085);
or U11529 (N_11529,N_4251,N_8137);
nand U11530 (N_11530,N_9782,N_3765);
xor U11531 (N_11531,N_4478,N_2867);
or U11532 (N_11532,N_9922,N_8597);
xnor U11533 (N_11533,N_287,N_7152);
nor U11534 (N_11534,N_6324,N_2433);
and U11535 (N_11535,N_650,N_886);
nand U11536 (N_11536,N_2561,N_4629);
nor U11537 (N_11537,N_3834,N_7548);
xor U11538 (N_11538,N_6746,N_5612);
xnor U11539 (N_11539,N_3719,N_149);
nor U11540 (N_11540,N_896,N_3941);
or U11541 (N_11541,N_5672,N_8791);
or U11542 (N_11542,N_1975,N_5733);
and U11543 (N_11543,N_5553,N_616);
or U11544 (N_11544,N_8405,N_9622);
nand U11545 (N_11545,N_2145,N_5113);
xnor U11546 (N_11546,N_6683,N_8508);
nor U11547 (N_11547,N_7110,N_9907);
and U11548 (N_11548,N_4007,N_716);
nor U11549 (N_11549,N_8223,N_7709);
nand U11550 (N_11550,N_8916,N_777);
or U11551 (N_11551,N_3985,N_3114);
nor U11552 (N_11552,N_9162,N_2857);
nor U11553 (N_11553,N_4085,N_6127);
or U11554 (N_11554,N_6455,N_2336);
xor U11555 (N_11555,N_334,N_2245);
nor U11556 (N_11556,N_2317,N_2730);
xnor U11557 (N_11557,N_283,N_9891);
or U11558 (N_11558,N_9995,N_4870);
xor U11559 (N_11559,N_4775,N_7505);
or U11560 (N_11560,N_3997,N_7491);
xnor U11561 (N_11561,N_4756,N_2912);
nand U11562 (N_11562,N_767,N_8315);
nor U11563 (N_11563,N_2229,N_7163);
nor U11564 (N_11564,N_2996,N_7368);
xnor U11565 (N_11565,N_110,N_9084);
nor U11566 (N_11566,N_8292,N_8325);
nand U11567 (N_11567,N_251,N_2464);
or U11568 (N_11568,N_9913,N_7485);
nand U11569 (N_11569,N_5755,N_4333);
xnor U11570 (N_11570,N_3230,N_7833);
xor U11571 (N_11571,N_5363,N_2631);
nor U11572 (N_11572,N_1418,N_4464);
xor U11573 (N_11573,N_1230,N_8528);
and U11574 (N_11574,N_2655,N_948);
and U11575 (N_11575,N_8067,N_3311);
and U11576 (N_11576,N_6275,N_6805);
or U11577 (N_11577,N_3621,N_3874);
and U11578 (N_11578,N_9635,N_4559);
xnor U11579 (N_11579,N_5851,N_7088);
xnor U11580 (N_11580,N_8387,N_5505);
xnor U11581 (N_11581,N_6471,N_7641);
or U11582 (N_11582,N_5521,N_8879);
nor U11583 (N_11583,N_7937,N_7957);
nor U11584 (N_11584,N_8,N_1342);
nand U11585 (N_11585,N_3150,N_3164);
nor U11586 (N_11586,N_1896,N_3095);
xnor U11587 (N_11587,N_2010,N_7809);
nand U11588 (N_11588,N_6502,N_2942);
or U11589 (N_11589,N_9166,N_7230);
and U11590 (N_11590,N_6124,N_1499);
or U11591 (N_11591,N_4016,N_2894);
nand U11592 (N_11592,N_7322,N_486);
nand U11593 (N_11593,N_7747,N_112);
or U11594 (N_11594,N_8212,N_47);
xor U11595 (N_11595,N_8171,N_2968);
or U11596 (N_11596,N_2417,N_428);
or U11597 (N_11597,N_5536,N_1034);
or U11598 (N_11598,N_4620,N_7608);
and U11599 (N_11599,N_4125,N_5014);
nor U11600 (N_11600,N_8888,N_4337);
or U11601 (N_11601,N_1882,N_1768);
nor U11602 (N_11602,N_3103,N_3828);
or U11603 (N_11603,N_8538,N_8574);
and U11604 (N_11604,N_8061,N_1114);
or U11605 (N_11605,N_2709,N_3507);
xor U11606 (N_11606,N_6121,N_7053);
and U11607 (N_11607,N_199,N_8971);
nor U11608 (N_11608,N_7476,N_2492);
or U11609 (N_11609,N_2883,N_7454);
xnor U11610 (N_11610,N_8384,N_3630);
and U11611 (N_11611,N_3063,N_3608);
or U11612 (N_11612,N_1107,N_9454);
or U11613 (N_11613,N_6141,N_8787);
nor U11614 (N_11614,N_4226,N_9005);
nand U11615 (N_11615,N_5464,N_8082);
xnor U11616 (N_11616,N_464,N_4303);
nand U11617 (N_11617,N_1754,N_211);
nand U11618 (N_11618,N_2866,N_4575);
xor U11619 (N_11619,N_1332,N_9002);
xor U11620 (N_11620,N_621,N_157);
and U11621 (N_11621,N_56,N_8773);
nand U11622 (N_11622,N_3570,N_342);
xnor U11623 (N_11623,N_4236,N_4383);
nor U11624 (N_11624,N_2735,N_7777);
xor U11625 (N_11625,N_6008,N_4613);
xnor U11626 (N_11626,N_4867,N_6209);
nor U11627 (N_11627,N_4882,N_9328);
nor U11628 (N_11628,N_2881,N_1958);
and U11629 (N_11629,N_3706,N_4411);
nor U11630 (N_11630,N_8569,N_238);
nand U11631 (N_11631,N_9661,N_7971);
or U11632 (N_11632,N_6422,N_4397);
xnor U11633 (N_11633,N_1857,N_1946);
or U11634 (N_11634,N_1541,N_4003);
nor U11635 (N_11635,N_3306,N_5002);
or U11636 (N_11636,N_3943,N_824);
or U11637 (N_11637,N_2647,N_247);
nand U11638 (N_11638,N_5332,N_7857);
nand U11639 (N_11639,N_2650,N_5706);
xnor U11640 (N_11640,N_4502,N_2487);
xnor U11641 (N_11641,N_8009,N_9667);
nor U11642 (N_11642,N_5633,N_8026);
and U11643 (N_11643,N_2125,N_2244);
or U11644 (N_11644,N_4356,N_8873);
nand U11645 (N_11645,N_4291,N_8565);
and U11646 (N_11646,N_4753,N_2795);
xnor U11647 (N_11647,N_15,N_4926);
xor U11648 (N_11648,N_6296,N_5310);
nand U11649 (N_11649,N_9038,N_8126);
nand U11650 (N_11650,N_4191,N_9368);
or U11651 (N_11651,N_2874,N_5949);
xnor U11652 (N_11652,N_9014,N_3073);
xor U11653 (N_11653,N_6751,N_7375);
and U11654 (N_11654,N_4198,N_4836);
or U11655 (N_11655,N_5124,N_9482);
and U11656 (N_11656,N_226,N_9047);
nor U11657 (N_11657,N_723,N_148);
nand U11658 (N_11658,N_7183,N_793);
xnor U11659 (N_11659,N_3629,N_4921);
or U11660 (N_11660,N_7631,N_2562);
xnor U11661 (N_11661,N_4406,N_9075);
xnor U11662 (N_11662,N_3752,N_3996);
xor U11663 (N_11663,N_3791,N_1520);
xnor U11664 (N_11664,N_6191,N_9772);
nand U11665 (N_11665,N_5065,N_7952);
nor U11666 (N_11666,N_6415,N_5141);
nand U11667 (N_11667,N_6862,N_9036);
or U11668 (N_11668,N_1175,N_4817);
or U11669 (N_11669,N_1290,N_5566);
or U11670 (N_11670,N_5258,N_8414);
and U11671 (N_11671,N_6009,N_2618);
nor U11672 (N_11672,N_4839,N_4167);
or U11673 (N_11673,N_540,N_6670);
nor U11674 (N_11674,N_3166,N_3890);
nand U11675 (N_11675,N_8716,N_1763);
nand U11676 (N_11676,N_9390,N_9273);
and U11677 (N_11677,N_1941,N_3451);
and U11678 (N_11678,N_8834,N_861);
and U11679 (N_11679,N_7866,N_8536);
nand U11680 (N_11680,N_9243,N_3415);
nand U11681 (N_11681,N_1804,N_1432);
xor U11682 (N_11682,N_3323,N_1127);
nor U11683 (N_11683,N_8623,N_1030);
or U11684 (N_11684,N_6816,N_3246);
or U11685 (N_11685,N_4267,N_8139);
xnor U11686 (N_11686,N_4782,N_5354);
or U11687 (N_11687,N_6892,N_8867);
or U11688 (N_11688,N_1395,N_6182);
nor U11689 (N_11689,N_3472,N_2985);
and U11690 (N_11690,N_7167,N_3812);
nand U11691 (N_11691,N_9198,N_3270);
or U11692 (N_11692,N_7956,N_8326);
or U11693 (N_11693,N_8647,N_8698);
or U11694 (N_11694,N_1007,N_8930);
xor U11695 (N_11695,N_993,N_2312);
and U11696 (N_11696,N_1196,N_2307);
xnor U11697 (N_11697,N_952,N_1165);
and U11698 (N_11698,N_5084,N_651);
nor U11699 (N_11699,N_902,N_6016);
nor U11700 (N_11700,N_4440,N_599);
and U11701 (N_11701,N_5116,N_7794);
nand U11702 (N_11702,N_6382,N_4331);
xor U11703 (N_11703,N_5573,N_7131);
nand U11704 (N_11704,N_633,N_3426);
nand U11705 (N_11705,N_1518,N_6568);
nor U11706 (N_11706,N_1378,N_9811);
xnor U11707 (N_11707,N_6307,N_5098);
and U11708 (N_11708,N_5640,N_973);
xor U11709 (N_11709,N_8750,N_28);
or U11710 (N_11710,N_5664,N_9232);
nor U11711 (N_11711,N_8577,N_9465);
xor U11712 (N_11712,N_8182,N_7652);
xnor U11713 (N_11713,N_7908,N_7459);
and U11714 (N_11714,N_815,N_6509);
nor U11715 (N_11715,N_666,N_3320);
xor U11716 (N_11716,N_8227,N_6675);
or U11717 (N_11717,N_8670,N_5274);
or U11718 (N_11718,N_8572,N_1891);
and U11719 (N_11719,N_2426,N_997);
xnor U11720 (N_11720,N_5383,N_878);
or U11721 (N_11721,N_6193,N_401);
and U11722 (N_11722,N_3205,N_4170);
xnor U11723 (N_11723,N_9780,N_6377);
xnor U11724 (N_11724,N_5068,N_2040);
nand U11725 (N_11725,N_4046,N_4810);
nor U11726 (N_11726,N_6344,N_9742);
xor U11727 (N_11727,N_9526,N_3520);
and U11728 (N_11728,N_6645,N_3721);
xnor U11729 (N_11729,N_4346,N_4606);
xor U11730 (N_11730,N_4651,N_2947);
nor U11731 (N_11731,N_1587,N_1316);
and U11732 (N_11732,N_5816,N_1441);
or U11733 (N_11733,N_8571,N_9875);
or U11734 (N_11734,N_2324,N_6433);
nor U11735 (N_11735,N_3992,N_2854);
nand U11736 (N_11736,N_9462,N_3787);
and U11737 (N_11737,N_5038,N_3674);
nor U11738 (N_11738,N_7469,N_3098);
and U11739 (N_11739,N_5683,N_2396);
and U11740 (N_11740,N_974,N_9391);
xnor U11741 (N_11741,N_4833,N_1345);
xnor U11742 (N_11742,N_6915,N_4393);
nor U11743 (N_11743,N_6906,N_3101);
or U11744 (N_11744,N_7565,N_5428);
nand U11745 (N_11745,N_8518,N_2557);
nand U11746 (N_11746,N_9734,N_5179);
nor U11747 (N_11747,N_7745,N_8891);
nor U11748 (N_11748,N_5908,N_5704);
nand U11749 (N_11749,N_6938,N_8512);
and U11750 (N_11750,N_6397,N_9629);
and U11751 (N_11751,N_9689,N_5887);
and U11752 (N_11752,N_6485,N_8431);
nand U11753 (N_11753,N_2217,N_5720);
nor U11754 (N_11754,N_843,N_9376);
and U11755 (N_11755,N_9919,N_5288);
and U11756 (N_11756,N_8704,N_8706);
xnor U11757 (N_11757,N_586,N_3400);
nand U11758 (N_11758,N_1555,N_142);
and U11759 (N_11759,N_5700,N_4272);
nor U11760 (N_11760,N_2257,N_850);
xnor U11761 (N_11761,N_9700,N_7034);
xor U11762 (N_11762,N_6096,N_5287);
nand U11763 (N_11763,N_8778,N_244);
and U11764 (N_11764,N_4420,N_9032);
xor U11765 (N_11765,N_1672,N_8231);
nor U11766 (N_11766,N_8625,N_3010);
and U11767 (N_11767,N_9405,N_5999);
or U11768 (N_11768,N_4243,N_5812);
and U11769 (N_11769,N_8225,N_398);
nand U11770 (N_11770,N_4262,N_9);
or U11771 (N_11771,N_3442,N_144);
xnor U11772 (N_11772,N_7346,N_4145);
nor U11773 (N_11773,N_7021,N_9329);
or U11774 (N_11774,N_5913,N_5983);
and U11775 (N_11775,N_1821,N_7760);
xnor U11776 (N_11776,N_5432,N_3083);
or U11777 (N_11777,N_5032,N_1490);
and U11778 (N_11778,N_140,N_8984);
or U11779 (N_11779,N_5977,N_5639);
nand U11780 (N_11780,N_9305,N_2291);
xnor U11781 (N_11781,N_771,N_6992);
nor U11782 (N_11782,N_694,N_9007);
or U11783 (N_11783,N_6314,N_9849);
xor U11784 (N_11784,N_3479,N_6041);
nor U11785 (N_11785,N_5333,N_1909);
or U11786 (N_11786,N_5397,N_7121);
xor U11787 (N_11787,N_1025,N_9011);
and U11788 (N_11788,N_1564,N_6409);
nor U11789 (N_11789,N_4352,N_7355);
and U11790 (N_11790,N_5240,N_54);
and U11791 (N_11791,N_7532,N_2605);
xnor U11792 (N_11792,N_7155,N_6592);
and U11793 (N_11793,N_8343,N_6760);
nand U11794 (N_11794,N_8042,N_5719);
nand U11795 (N_11795,N_4078,N_8021);
nand U11796 (N_11796,N_3888,N_6898);
nor U11797 (N_11797,N_6312,N_567);
and U11798 (N_11798,N_852,N_2022);
or U11799 (N_11799,N_3085,N_2311);
xor U11800 (N_11800,N_1494,N_4593);
or U11801 (N_11801,N_5041,N_6800);
or U11802 (N_11802,N_1311,N_5361);
and U11803 (N_11803,N_4042,N_9089);
xnor U11804 (N_11804,N_5783,N_8699);
xor U11805 (N_11805,N_3032,N_9827);
nor U11806 (N_11806,N_3425,N_5677);
xnor U11807 (N_11807,N_2121,N_5259);
nor U11808 (N_11808,N_1605,N_9968);
nand U11809 (N_11809,N_2048,N_8582);
xnor U11810 (N_11810,N_3688,N_4754);
or U11811 (N_11811,N_9244,N_1456);
nor U11812 (N_11812,N_2895,N_608);
nor U11813 (N_11813,N_1855,N_6561);
and U11814 (N_11814,N_6219,N_7449);
and U11815 (N_11815,N_3554,N_787);
or U11816 (N_11816,N_1951,N_658);
nand U11817 (N_11817,N_5638,N_9340);
nor U11818 (N_11818,N_525,N_3961);
or U11819 (N_11819,N_6578,N_3868);
and U11820 (N_11820,N_7203,N_9551);
xor U11821 (N_11821,N_2176,N_2008);
or U11822 (N_11822,N_1479,N_5594);
nand U11823 (N_11823,N_9632,N_9161);
xnor U11824 (N_11824,N_6983,N_8081);
nor U11825 (N_11825,N_4913,N_2608);
nand U11826 (N_11826,N_2848,N_702);
nor U11827 (N_11827,N_7036,N_7386);
xor U11828 (N_11828,N_7556,N_2667);
or U11829 (N_11829,N_2840,N_4691);
nor U11830 (N_11830,N_2050,N_4122);
nand U11831 (N_11831,N_8022,N_3988);
nand U11832 (N_11832,N_2917,N_6970);
nor U11833 (N_11833,N_3139,N_2471);
and U11834 (N_11834,N_7752,N_6199);
and U11835 (N_11835,N_348,N_3659);
xor U11836 (N_11836,N_2060,N_8676);
and U11837 (N_11837,N_2446,N_6641);
or U11838 (N_11838,N_2314,N_4405);
nor U11839 (N_11839,N_470,N_3544);
xor U11840 (N_11840,N_2308,N_7792);
xnor U11841 (N_11841,N_7660,N_4979);
and U11842 (N_11842,N_1880,N_2627);
or U11843 (N_11843,N_5431,N_1228);
xor U11844 (N_11844,N_9710,N_7284);
nor U11845 (N_11845,N_9671,N_1305);
xnor U11846 (N_11846,N_6297,N_4037);
xnor U11847 (N_11847,N_780,N_3954);
nand U11848 (N_11848,N_7111,N_4618);
nand U11849 (N_11849,N_6922,N_2190);
or U11850 (N_11850,N_6078,N_9681);
xor U11851 (N_11851,N_601,N_8038);
nand U11852 (N_11852,N_3299,N_5646);
nor U11853 (N_11853,N_4834,N_7509);
nand U11854 (N_11854,N_2369,N_8581);
nand U11855 (N_11855,N_962,N_1033);
nor U11856 (N_11856,N_783,N_2508);
and U11857 (N_11857,N_8194,N_4196);
or U11858 (N_11858,N_6135,N_7700);
nor U11859 (N_11859,N_4855,N_498);
or U11860 (N_11860,N_9597,N_1273);
and U11861 (N_11861,N_9311,N_4048);
and U11862 (N_11862,N_8048,N_9200);
nand U11863 (N_11863,N_6582,N_3831);
xnor U11864 (N_11864,N_6554,N_8150);
nor U11865 (N_11865,N_4723,N_4160);
nor U11866 (N_11866,N_5457,N_2435);
xnor U11867 (N_11867,N_3526,N_2298);
xor U11868 (N_11868,N_1012,N_8448);
nand U11869 (N_11869,N_7582,N_9895);
nor U11870 (N_11870,N_7541,N_5883);
xnor U11871 (N_11871,N_562,N_2465);
or U11872 (N_11872,N_6169,N_2891);
nand U11873 (N_11873,N_579,N_3428);
or U11874 (N_11874,N_7748,N_2393);
xor U11875 (N_11875,N_3294,N_9241);
or U11876 (N_11876,N_1088,N_5624);
or U11877 (N_11877,N_5088,N_7500);
nand U11878 (N_11878,N_4772,N_7567);
or U11879 (N_11879,N_1660,N_3969);
nor U11880 (N_11880,N_3605,N_3811);
or U11881 (N_11881,N_7267,N_4683);
xnor U11882 (N_11882,N_6727,N_3915);
nor U11883 (N_11883,N_3204,N_132);
and U11884 (N_11884,N_1737,N_6086);
nand U11885 (N_11885,N_7251,N_3093);
nor U11886 (N_11886,N_9470,N_807);
and U11887 (N_11887,N_4482,N_4796);
xnor U11888 (N_11888,N_8066,N_3302);
nor U11889 (N_11889,N_7566,N_5875);
nor U11890 (N_11890,N_7435,N_6969);
xnor U11891 (N_11891,N_2044,N_7875);
or U11892 (N_11892,N_7844,N_5670);
xor U11893 (N_11893,N_5368,N_6625);
nor U11894 (N_11894,N_5864,N_695);
xor U11895 (N_11895,N_7164,N_7456);
and U11896 (N_11896,N_3198,N_7689);
xor U11897 (N_11897,N_2382,N_2626);
xnor U11898 (N_11898,N_6632,N_2967);
nor U11899 (N_11899,N_959,N_7584);
nor U11900 (N_11900,N_9604,N_1161);
nand U11901 (N_11901,N_2915,N_9285);
nand U11902 (N_11902,N_2760,N_6477);
xnor U11903 (N_11903,N_8737,N_2141);
or U11904 (N_11904,N_6855,N_52);
and U11905 (N_11905,N_1601,N_1399);
nand U11906 (N_11906,N_9467,N_2898);
and U11907 (N_11907,N_8346,N_6847);
xor U11908 (N_11908,N_5394,N_6184);
nand U11909 (N_11909,N_2746,N_3860);
and U11910 (N_11910,N_9638,N_9967);
xnor U11911 (N_11911,N_2363,N_9888);
nand U11912 (N_11912,N_8892,N_9673);
and U11913 (N_11913,N_176,N_3944);
or U11914 (N_11914,N_2803,N_1194);
or U11915 (N_11915,N_2980,N_524);
or U11916 (N_11916,N_5314,N_7902);
nand U11917 (N_11917,N_7552,N_2274);
and U11918 (N_11918,N_4823,N_2309);
nand U11919 (N_11919,N_4647,N_2005);
and U11920 (N_11920,N_2265,N_5300);
nand U11921 (N_11921,N_1338,N_6293);
nor U11922 (N_11922,N_8019,N_7336);
and U11923 (N_11923,N_1340,N_1061);
or U11924 (N_11924,N_1531,N_7037);
nand U11925 (N_11925,N_2665,N_6968);
nor U11926 (N_11926,N_5598,N_1363);
xnor U11927 (N_11927,N_845,N_241);
nor U11928 (N_11928,N_4670,N_8729);
and U11929 (N_11929,N_9534,N_4506);
nor U11930 (N_11930,N_1699,N_1398);
and U11931 (N_11931,N_6692,N_9512);
and U11932 (N_11932,N_9448,N_7968);
nand U11933 (N_11933,N_8558,N_305);
or U11934 (N_11934,N_8032,N_8728);
and U11935 (N_11935,N_5253,N_5204);
nand U11936 (N_11936,N_9764,N_4507);
xnor U11937 (N_11937,N_9626,N_5023);
xnor U11938 (N_11938,N_5173,N_1465);
xnor U11939 (N_11939,N_2514,N_2091);
nor U11940 (N_11940,N_1100,N_8264);
and U11941 (N_11941,N_7953,N_7861);
nor U11942 (N_11942,N_5501,N_8167);
or U11943 (N_11943,N_3662,N_2143);
nand U11944 (N_11944,N_9594,N_4968);
xor U11945 (N_11945,N_8927,N_2983);
nor U11946 (N_11946,N_6126,N_7849);
or U11947 (N_11947,N_2601,N_4091);
nand U11948 (N_11948,N_5239,N_3416);
and U11949 (N_11949,N_8705,N_4531);
xor U11950 (N_11950,N_2949,N_2400);
nor U11951 (N_11951,N_4063,N_2784);
xnor U11952 (N_11952,N_5842,N_8422);
nor U11953 (N_11953,N_9155,N_6281);
nand U11954 (N_11954,N_1258,N_6534);
and U11955 (N_11955,N_8741,N_7114);
or U11956 (N_11956,N_8614,N_2796);
or U11957 (N_11957,N_9803,N_5588);
and U11958 (N_11958,N_1415,N_4367);
nor U11959 (N_11959,N_9959,N_9567);
nand U11960 (N_11960,N_6952,N_227);
xor U11961 (N_11961,N_5004,N_8106);
xnor U11962 (N_11962,N_3668,N_6543);
and U11963 (N_11963,N_629,N_5099);
nand U11964 (N_11964,N_966,N_3939);
xnor U11965 (N_11965,N_8270,N_6838);
nand U11966 (N_11966,N_2499,N_2577);
nand U11967 (N_11967,N_1298,N_3202);
nand U11968 (N_11968,N_6642,N_5771);
and U11969 (N_11969,N_6643,N_4685);
or U11970 (N_11970,N_2073,N_2748);
or U11971 (N_11971,N_1067,N_6724);
or U11972 (N_11972,N_8717,N_5645);
nand U11973 (N_11973,N_332,N_3505);
nor U11974 (N_11974,N_9737,N_6391);
and U11975 (N_11975,N_736,N_5550);
xnor U11976 (N_11976,N_817,N_3980);
xnor U11977 (N_11977,N_8548,N_4910);
nor U11978 (N_11978,N_7910,N_2429);
xnor U11979 (N_11979,N_1772,N_6999);
xnor U11980 (N_11980,N_5508,N_4210);
nand U11981 (N_11981,N_4582,N_1171);
and U11982 (N_11982,N_888,N_8479);
xor U11983 (N_11983,N_6361,N_7793);
and U11984 (N_11984,N_8793,N_9149);
or U11985 (N_11985,N_3542,N_3987);
or U11986 (N_11986,N_2929,N_8617);
or U11987 (N_11987,N_6368,N_1676);
or U11988 (N_11988,N_1036,N_1248);
xnor U11989 (N_11989,N_3255,N_374);
nor U11990 (N_11990,N_9850,N_2964);
nor U11991 (N_11991,N_9833,N_8095);
and U11992 (N_11992,N_5814,N_2653);
xnor U11993 (N_11993,N_895,N_9753);
nand U11994 (N_11994,N_3389,N_1076);
nand U11995 (N_11995,N_3357,N_2367);
xor U11996 (N_11996,N_1309,N_8301);
nor U11997 (N_11997,N_8560,N_2118);
or U11998 (N_11998,N_8247,N_9645);
and U11999 (N_11999,N_3017,N_6996);
and U12000 (N_12000,N_4726,N_6656);
xnor U12001 (N_12001,N_5895,N_4168);
or U12002 (N_12002,N_5808,N_7358);
nand U12003 (N_12003,N_5419,N_6417);
nor U12004 (N_12004,N_5479,N_6876);
xor U12005 (N_12005,N_7472,N_1021);
and U12006 (N_12006,N_7046,N_2783);
xor U12007 (N_12007,N_5249,N_8989);
xnor U12008 (N_12008,N_4401,N_776);
and U12009 (N_12009,N_3806,N_8939);
nor U12010 (N_12010,N_6031,N_1670);
nand U12011 (N_12011,N_9239,N_7606);
or U12012 (N_12012,N_9403,N_2399);
nand U12013 (N_12013,N_3365,N_8719);
or U12014 (N_12014,N_7595,N_9605);
or U12015 (N_12015,N_9485,N_7279);
nor U12016 (N_12016,N_2078,N_3667);
and U12017 (N_12017,N_2590,N_8911);
nand U12018 (N_12018,N_7104,N_8949);
xnor U12019 (N_12019,N_190,N_5515);
nand U12020 (N_12020,N_4996,N_3105);
and U12021 (N_12021,N_6187,N_8455);
nor U12022 (N_12022,N_1481,N_1374);
and U12023 (N_12023,N_7674,N_1233);
or U12024 (N_12024,N_3386,N_9989);
or U12025 (N_12025,N_3046,N_4363);
and U12026 (N_12026,N_1696,N_9327);
nor U12027 (N_12027,N_9270,N_8632);
or U12028 (N_12028,N_996,N_4946);
nor U12029 (N_12029,N_4655,N_7231);
nand U12030 (N_12030,N_2831,N_8332);
and U12031 (N_12031,N_6956,N_2999);
xor U12032 (N_12032,N_6015,N_2810);
nor U12033 (N_12033,N_3401,N_1583);
nand U12034 (N_12034,N_8584,N_371);
or U12035 (N_12035,N_4686,N_8822);
and U12036 (N_12036,N_9813,N_6835);
or U12037 (N_12037,N_5589,N_4692);
or U12038 (N_12038,N_2984,N_5813);
and U12039 (N_12039,N_198,N_4607);
xnor U12040 (N_12040,N_2051,N_1610);
nor U12041 (N_12041,N_8655,N_6910);
and U12042 (N_12042,N_4444,N_3420);
xor U12043 (N_12043,N_3589,N_549);
or U12044 (N_12044,N_8075,N_1656);
nand U12045 (N_12045,N_7069,N_4804);
and U12046 (N_12046,N_3231,N_4185);
and U12047 (N_12047,N_6356,N_5246);
xnor U12048 (N_12048,N_6812,N_7112);
and U12049 (N_12049,N_4353,N_4800);
nor U12050 (N_12050,N_5837,N_5968);
nor U12051 (N_12051,N_8899,N_6512);
nand U12052 (N_12052,N_7822,N_5495);
nor U12053 (N_12053,N_4247,N_9721);
nand U12054 (N_12054,N_8795,N_699);
nor U12055 (N_12055,N_7020,N_7654);
nor U12056 (N_12056,N_3064,N_2392);
nand U12057 (N_12057,N_3080,N_8255);
nand U12058 (N_12058,N_1451,N_4978);
nor U12059 (N_12059,N_6553,N_5610);
and U12060 (N_12060,N_8562,N_8944);
and U12061 (N_12061,N_5123,N_3200);
nand U12062 (N_12062,N_1634,N_2387);
nand U12063 (N_12063,N_2066,N_504);
nor U12064 (N_12064,N_7433,N_4736);
xor U12065 (N_12065,N_748,N_4952);
nor U12066 (N_12066,N_5467,N_1862);
nor U12067 (N_12067,N_6697,N_3496);
or U12068 (N_12068,N_3362,N_1981);
xnor U12069 (N_12069,N_3736,N_1982);
nor U12070 (N_12070,N_9739,N_2099);
and U12071 (N_12071,N_8226,N_3802);
or U12072 (N_12072,N_6392,N_2714);
nand U12073 (N_12073,N_6571,N_8590);
nor U12074 (N_12074,N_4777,N_8411);
and U12075 (N_12075,N_4293,N_6525);
and U12076 (N_12076,N_9356,N_2611);
and U12077 (N_12077,N_4584,N_5796);
or U12078 (N_12078,N_508,N_9669);
nor U12079 (N_12079,N_289,N_2361);
and U12080 (N_12080,N_3129,N_7924);
nor U12081 (N_12081,N_5194,N_4213);
and U12082 (N_12082,N_3280,N_6076);
or U12083 (N_12083,N_4752,N_1611);
nor U12084 (N_12084,N_4992,N_1385);
and U12085 (N_12085,N_8697,N_8094);
or U12086 (N_12086,N_6250,N_7563);
xnor U12087 (N_12087,N_5061,N_6113);
and U12088 (N_12088,N_479,N_8146);
xnor U12089 (N_12089,N_1973,N_1731);
nor U12090 (N_12090,N_8685,N_3251);
and U12091 (N_12091,N_6666,N_926);
and U12092 (N_12092,N_336,N_4875);
nand U12093 (N_12093,N_3524,N_1679);
nand U12094 (N_12094,N_1080,N_7896);
and U12095 (N_12095,N_7100,N_9558);
xor U12096 (N_12096,N_2928,N_9925);
nor U12097 (N_12097,N_2657,N_7989);
or U12098 (N_12098,N_5481,N_9050);
xnor U12099 (N_12099,N_8689,N_9215);
nor U12100 (N_12100,N_5923,N_7);
xor U12101 (N_12101,N_3403,N_9517);
and U12102 (N_12102,N_243,N_4783);
nor U12103 (N_12103,N_4764,N_7973);
and U12104 (N_12104,N_2443,N_3882);
xnor U12105 (N_12105,N_1787,N_6794);
nand U12106 (N_12106,N_1279,N_943);
nand U12107 (N_12107,N_9322,N_8025);
nor U12108 (N_12108,N_9624,N_5815);
nand U12109 (N_12109,N_8559,N_8027);
and U12110 (N_12110,N_5322,N_3187);
nand U12111 (N_12111,N_3631,N_6810);
or U12112 (N_12112,N_5213,N_7958);
nor U12113 (N_12113,N_6436,N_1104);
or U12114 (N_12114,N_6390,N_7493);
nor U12115 (N_12115,N_2233,N_5152);
nand U12116 (N_12116,N_6,N_6101);
and U12117 (N_12117,N_3537,N_88);
xnor U12118 (N_12118,N_4364,N_4184);
or U12119 (N_12119,N_1148,N_4508);
nor U12120 (N_12120,N_7803,N_7283);
or U12121 (N_12121,N_6520,N_40);
or U12122 (N_12122,N_2773,N_5757);
and U12123 (N_12123,N_9281,N_4770);
nor U12124 (N_12124,N_385,N_5138);
or U12125 (N_12125,N_4806,N_4410);
or U12126 (N_12126,N_2256,N_7220);
and U12127 (N_12127,N_5509,N_4345);
and U12128 (N_12128,N_7917,N_7891);
or U12129 (N_12129,N_708,N_8517);
xor U12130 (N_12130,N_5275,N_3979);
and U12131 (N_12131,N_7679,N_9343);
xnor U12132 (N_12132,N_4843,N_2053);
and U12133 (N_12133,N_3061,N_6528);
nand U12134 (N_12134,N_9296,N_6788);
nand U12135 (N_12135,N_705,N_3482);
or U12136 (N_12136,N_8624,N_3295);
and U12137 (N_12137,N_8433,N_5197);
nor U12138 (N_12138,N_3081,N_2707);
or U12139 (N_12139,N_7658,N_2793);
nand U12140 (N_12140,N_6045,N_2210);
nor U12141 (N_12141,N_6222,N_6650);
xor U12142 (N_12142,N_9141,N_8056);
nor U12143 (N_12143,N_5266,N_1400);
or U12144 (N_12144,N_2211,N_5057);
nor U12145 (N_12145,N_5308,N_5230);
nor U12146 (N_12146,N_1153,N_5180);
nor U12147 (N_12147,N_3380,N_8416);
xor U12148 (N_12148,N_5647,N_2285);
nor U12149 (N_12149,N_5359,N_768);
and U12150 (N_12150,N_2596,N_4776);
xor U12151 (N_12151,N_8969,N_8887);
and U12152 (N_12152,N_4076,N_3687);
xnor U12153 (N_12153,N_8486,N_529);
nand U12154 (N_12154,N_3967,N_7772);
nand U12155 (N_12155,N_8606,N_3497);
nor U12156 (N_12156,N_356,N_6877);
xor U12157 (N_12157,N_9553,N_3710);
nand U12158 (N_12158,N_9389,N_8076);
nand U12159 (N_12159,N_3337,N_7120);
nor U12160 (N_12160,N_4594,N_231);
xnor U12161 (N_12161,N_9585,N_6441);
xor U12162 (N_12162,N_2960,N_8983);
xnor U12163 (N_12163,N_6179,N_6445);
xnor U12164 (N_12164,N_4514,N_2532);
nand U12165 (N_12165,N_3208,N_1883);
nor U12166 (N_12166,N_3138,N_8390);
and U12167 (N_12167,N_3803,N_1764);
or U12168 (N_12168,N_8849,N_5517);
nor U12169 (N_12169,N_6516,N_5096);
nor U12170 (N_12170,N_9930,N_4180);
or U12171 (N_12171,N_5225,N_4689);
xor U12172 (N_12172,N_8549,N_7869);
nor U12173 (N_12173,N_7998,N_8488);
xor U12174 (N_12174,N_2491,N_306);
nor U12175 (N_12175,N_246,N_5679);
nand U12176 (N_12176,N_7763,N_4786);
nor U12177 (N_12177,N_7370,N_5531);
or U12178 (N_12178,N_1352,N_2380);
xnor U12179 (N_12179,N_7544,N_5914);
xnor U12180 (N_12180,N_9774,N_9707);
nand U12181 (N_12181,N_7913,N_9096);
and U12182 (N_12182,N_21,N_3810);
xor U12183 (N_12183,N_2019,N_1355);
xor U12184 (N_12184,N_8453,N_1867);
nor U12185 (N_12185,N_7980,N_6853);
nor U12186 (N_12186,N_7730,N_5995);
nand U12187 (N_12187,N_4767,N_5450);
nand U12188 (N_12188,N_499,N_7082);
or U12189 (N_12189,N_2838,N_7856);
and U12190 (N_12190,N_9637,N_6396);
or U12191 (N_12191,N_4432,N_5458);
nor U12192 (N_12192,N_5365,N_5353);
nor U12193 (N_12193,N_9464,N_2715);
or U12194 (N_12194,N_4665,N_377);
nor U12195 (N_12195,N_2445,N_7545);
and U12196 (N_12196,N_9760,N_9309);
xor U12197 (N_12197,N_1162,N_5821);
and U12198 (N_12198,N_7017,N_4434);
nor U12199 (N_12199,N_7383,N_908);
xnor U12200 (N_12200,N_2955,N_591);
nand U12201 (N_12201,N_8542,N_5101);
nand U12202 (N_12202,N_2659,N_4013);
xnor U12203 (N_12203,N_8586,N_320);
and U12204 (N_12204,N_8540,N_4715);
xor U12205 (N_12205,N_8922,N_6117);
or U12206 (N_12206,N_1977,N_2481);
or U12207 (N_12207,N_2069,N_1447);
nor U12208 (N_12208,N_4704,N_1336);
nand U12209 (N_12209,N_9388,N_3887);
and U12210 (N_12210,N_5316,N_3525);
or U12211 (N_12211,N_2296,N_563);
nand U12212 (N_12212,N_7501,N_3192);
and U12213 (N_12213,N_6828,N_4702);
nand U12214 (N_12214,N_3099,N_9878);
xnor U12215 (N_12215,N_5524,N_8338);
nand U12216 (N_12216,N_7391,N_8400);
nand U12217 (N_12217,N_8249,N_1934);
xor U12218 (N_12218,N_3731,N_6319);
and U12219 (N_12219,N_6631,N_3422);
xnor U12220 (N_12220,N_1286,N_3906);
xor U12221 (N_12221,N_7218,N_3054);
xor U12222 (N_12222,N_5643,N_1974);
or U12223 (N_12223,N_5586,N_5714);
and U12224 (N_12224,N_2014,N_3290);
nor U12225 (N_12225,N_9896,N_5602);
nor U12226 (N_12226,N_4151,N_2889);
or U12227 (N_12227,N_5264,N_155);
and U12228 (N_12228,N_9355,N_6937);
and U12229 (N_12229,N_2021,N_6530);
and U12230 (N_12230,N_3777,N_3551);
xor U12231 (N_12231,N_1500,N_4431);
or U12232 (N_12232,N_5424,N_2366);
and U12233 (N_12233,N_3133,N_304);
nor U12234 (N_12234,N_8681,N_4455);
or U12235 (N_12235,N_913,N_7846);
nand U12236 (N_12236,N_8506,N_3853);
and U12237 (N_12237,N_4829,N_63);
or U12238 (N_12238,N_465,N_9460);
nand U12239 (N_12239,N_1728,N_6139);
or U12240 (N_12240,N_5433,N_6764);
nor U12241 (N_12241,N_9834,N_1449);
or U12242 (N_12242,N_3475,N_6254);
xor U12243 (N_12243,N_234,N_5447);
nor U12244 (N_12244,N_3163,N_3285);
nand U12245 (N_12245,N_9506,N_2792);
xor U12246 (N_12246,N_6431,N_8763);
nor U12247 (N_12247,N_7003,N_409);
or U12248 (N_12248,N_8621,N_6470);
and U12249 (N_12249,N_7540,N_6164);
and U12250 (N_12250,N_5389,N_314);
xor U12251 (N_12251,N_7244,N_3379);
nor U12252 (N_12252,N_3732,N_3778);
xor U12253 (N_12253,N_6410,N_5810);
nand U12254 (N_12254,N_642,N_400);
nor U12255 (N_12255,N_8827,N_6129);
or U12256 (N_12256,N_820,N_3916);
and U12257 (N_12257,N_3934,N_9092);
nand U12258 (N_12258,N_7514,N_9445);
xnor U12259 (N_12259,N_961,N_9418);
nor U12260 (N_12260,N_3121,N_611);
nand U12261 (N_12261,N_7533,N_7806);
nand U12262 (N_12262,N_5035,N_8996);
and U12263 (N_12263,N_6294,N_7732);
and U12264 (N_12264,N_7138,N_5131);
xor U12265 (N_12265,N_2893,N_7948);
nor U12266 (N_12266,N_9237,N_6240);
nand U12267 (N_12267,N_626,N_5841);
xnor U12268 (N_12268,N_4708,N_929);
nor U12269 (N_12269,N_6211,N_2957);
xnor U12270 (N_12270,N_2249,N_9705);
xor U12271 (N_12271,N_722,N_9755);
nor U12272 (N_12272,N_2851,N_2167);
xor U12273 (N_12273,N_9678,N_3239);
xnor U12274 (N_12274,N_7415,N_558);
and U12275 (N_12275,N_4982,N_2068);
nor U12276 (N_12276,N_4600,N_915);
nand U12277 (N_12277,N_1450,N_1160);
or U12278 (N_12278,N_4947,N_386);
nor U12279 (N_12279,N_5625,N_2120);
and U12280 (N_12280,N_8556,N_7677);
nand U12281 (N_12281,N_8360,N_5963);
or U12282 (N_12282,N_4605,N_8363);
nor U12283 (N_12283,N_5556,N_5986);
xnor U12284 (N_12284,N_9375,N_760);
nand U12285 (N_12285,N_7673,N_766);
and U12286 (N_12286,N_5370,N_127);
or U12287 (N_12287,N_3009,N_9035);
nor U12288 (N_12288,N_3001,N_9652);
and U12289 (N_12289,N_8164,N_6603);
nor U12290 (N_12290,N_2825,N_1412);
nand U12291 (N_12291,N_5218,N_7800);
nand U12292 (N_12292,N_8759,N_5632);
or U12293 (N_12293,N_8096,N_3894);
and U12294 (N_12294,N_3132,N_346);
xnor U12295 (N_12295,N_5827,N_8475);
or U12296 (N_12296,N_9313,N_2287);
nor U12297 (N_12297,N_7118,N_8814);
xnor U12298 (N_12298,N_5454,N_108);
xor U12299 (N_12299,N_3275,N_1019);
nand U12300 (N_12300,N_6506,N_7458);
and U12301 (N_12301,N_9886,N_5392);
and U12302 (N_12302,N_7853,N_9227);
nand U12303 (N_12303,N_6934,N_2549);
nor U12304 (N_12304,N_9446,N_1609);
and U12305 (N_12305,N_5948,N_2110);
nor U12306 (N_12306,N_8404,N_643);
nor U12307 (N_12307,N_8327,N_1663);
xnor U12308 (N_12308,N_8869,N_5150);
or U12309 (N_12309,N_67,N_1919);
nand U12310 (N_12310,N_6337,N_5425);
or U12311 (N_12311,N_7000,N_1069);
xor U12312 (N_12312,N_9063,N_295);
or U12313 (N_12313,N_8114,N_2294);
xor U12314 (N_12314,N_6600,N_2101);
nor U12315 (N_12315,N_1002,N_2701);
xor U12316 (N_12316,N_2816,N_8505);
or U12317 (N_12317,N_3948,N_5892);
or U12318 (N_12318,N_460,N_9515);
nor U12319 (N_12319,N_3625,N_517);
nor U12320 (N_12320,N_5366,N_6866);
and U12321 (N_12321,N_9812,N_7656);
nor U12322 (N_12322,N_8851,N_5408);
or U12323 (N_12323,N_1899,N_3700);
nor U12324 (N_12324,N_739,N_4188);
xnor U12325 (N_12325,N_3111,N_4735);
nand U12326 (N_12326,N_877,N_9488);
nand U12327 (N_12327,N_8297,N_8880);
and U12328 (N_12328,N_1586,N_2028);
or U12329 (N_12329,N_9312,N_6754);
xnor U12330 (N_12330,N_2586,N_1885);
nand U12331 (N_12331,N_3826,N_3414);
or U12332 (N_12332,N_8912,N_9298);
and U12333 (N_12333,N_8815,N_6639);
and U12334 (N_12334,N_3062,N_1320);
nor U12335 (N_12335,N_6585,N_4974);
and U12336 (N_12336,N_2595,N_136);
and U12337 (N_12337,N_8732,N_4650);
or U12338 (N_12338,N_4695,N_4350);
and U12339 (N_12339,N_7714,N_7579);
and U12340 (N_12340,N_8177,N_1758);
xor U12341 (N_12341,N_4487,N_3991);
nand U12342 (N_12342,N_1771,N_7196);
nand U12343 (N_12343,N_5711,N_8023);
nand U12344 (N_12344,N_6022,N_3366);
nor U12345 (N_12345,N_317,N_8282);
nor U12346 (N_12346,N_7900,N_9545);
nand U12347 (N_12347,N_177,N_1287);
or U12348 (N_12348,N_6976,N_98);
nor U12349 (N_12349,N_4588,N_405);
and U12350 (N_12350,N_5546,N_3555);
or U12351 (N_12351,N_4128,N_9778);
nand U12352 (N_12352,N_9650,N_2721);
nand U12353 (N_12353,N_8464,N_6466);
nand U12354 (N_12354,N_1359,N_2786);
or U12355 (N_12355,N_9674,N_1289);
nor U12356 (N_12356,N_8862,N_7591);
or U12357 (N_12357,N_7682,N_5547);
xnor U12358 (N_12358,N_7694,N_5130);
or U12359 (N_12359,N_8442,N_3982);
nor U12360 (N_12360,N_5926,N_1326);
or U12361 (N_12361,N_1347,N_5437);
xor U12362 (N_12362,N_5063,N_7578);
nand U12363 (N_12363,N_7883,N_9749);
nand U12364 (N_12364,N_1185,N_8537);
nand U12365 (N_12365,N_2552,N_1628);
nor U12366 (N_12366,N_7393,N_2868);
xnor U12367 (N_12367,N_2111,N_7762);
xnor U12368 (N_12368,N_1087,N_5629);
nor U12369 (N_12369,N_6613,N_931);
and U12370 (N_12370,N_8919,N_3033);
and U12371 (N_12371,N_6246,N_654);
xor U12372 (N_12372,N_7470,N_8275);
xnor U12373 (N_12373,N_7818,N_1874);
nand U12374 (N_12374,N_1038,N_5092);
nor U12375 (N_12375,N_4975,N_2004);
nand U12376 (N_12376,N_8803,N_3361);
xnor U12377 (N_12377,N_4203,N_6755);
nand U12378 (N_12378,N_2946,N_6813);
and U12379 (N_12379,N_9183,N_9653);
nor U12380 (N_12380,N_1101,N_8642);
nand U12381 (N_12381,N_8319,N_3075);
nand U12382 (N_12382,N_5294,N_4881);
and U12383 (N_12383,N_5236,N_7102);
and U12384 (N_12384,N_9040,N_7573);
or U12385 (N_12385,N_917,N_1561);
and U12386 (N_12386,N_4498,N_6519);
nand U12387 (N_12387,N_6360,N_9136);
and U12388 (N_12388,N_9326,N_9586);
and U12389 (N_12389,N_5569,N_328);
and U12390 (N_12390,N_4534,N_5585);
nor U12391 (N_12391,N_3994,N_4278);
xnor U12392 (N_12392,N_2038,N_8567);
xor U12393 (N_12393,N_2961,N_1907);
xnor U12394 (N_12394,N_4413,N_8546);
nand U12395 (N_12395,N_1205,N_8669);
xor U12396 (N_12396,N_7852,N_9263);
xnor U12397 (N_12397,N_4249,N_2451);
nor U12398 (N_12398,N_9936,N_5121);
nand U12399 (N_12399,N_5352,N_5828);
nand U12400 (N_12400,N_5666,N_7232);
nor U12401 (N_12401,N_9493,N_7178);
nand U12402 (N_12402,N_7813,N_835);
and U12403 (N_12403,N_5649,N_5686);
xor U12404 (N_12404,N_2628,N_7345);
nand U12405 (N_12405,N_4483,N_9138);
xor U12406 (N_12406,N_7613,N_6068);
and U12407 (N_12407,N_4812,N_9680);
and U12408 (N_12408,N_2664,N_9649);
or U12409 (N_12409,N_6817,N_8308);
and U12410 (N_12410,N_2180,N_7006);
or U12411 (N_12411,N_9121,N_9885);
nor U12412 (N_12412,N_288,N_4932);
and U12413 (N_12413,N_5104,N_6786);
and U12414 (N_12414,N_2034,N_319);
nand U12415 (N_12415,N_1614,N_1016);
xor U12416 (N_12416,N_9578,N_5452);
nand U12417 (N_12417,N_5726,N_4068);
or U12418 (N_12418,N_6027,N_1792);
nor U12419 (N_12419,N_6821,N_1926);
xnor U12420 (N_12420,N_7557,N_1701);
nand U12421 (N_12421,N_5044,N_4876);
and U12422 (N_12422,N_5898,N_2462);
xnor U12423 (N_12423,N_2675,N_9071);
nand U12424 (N_12424,N_4402,N_2531);
and U12425 (N_12425,N_7085,N_2218);
xor U12426 (N_12426,N_6542,N_2513);
and U12427 (N_12427,N_3281,N_6080);
nor U12428 (N_12428,N_8726,N_5716);
or U12429 (N_12429,N_5122,N_7475);
xnor U12430 (N_12430,N_5071,N_5028);
xnor U12431 (N_12431,N_2011,N_7048);
nand U12432 (N_12432,N_1092,N_2461);
xnor U12433 (N_12433,N_4454,N_281);
nand U12434 (N_12434,N_967,N_8238);
nor U12435 (N_12435,N_6701,N_3445);
xor U12436 (N_12436,N_284,N_7716);
nor U12437 (N_12437,N_3459,N_169);
nand U12438 (N_12438,N_7089,N_713);
xor U12439 (N_12439,N_7457,N_9961);
and U12440 (N_12440,N_3318,N_8418);
nand U12441 (N_12441,N_751,N_3986);
and U12442 (N_12442,N_9625,N_164);
nand U12443 (N_12443,N_9447,N_9010);
nor U12444 (N_12444,N_6820,N_4258);
or U12445 (N_12445,N_6305,N_2438);
or U12446 (N_12446,N_5980,N_7923);
xnor U12447 (N_12447,N_1984,N_7659);
nand U12448 (N_12448,N_373,N_2432);
and U12449 (N_12449,N_8101,N_1708);
xor U12450 (N_12450,N_2394,N_5011);
xor U12451 (N_12451,N_1582,N_5345);
nor U12452 (N_12452,N_3349,N_2290);
nand U12453 (N_12453,N_8802,N_4491);
xor U12454 (N_12454,N_4271,N_5360);
or U12455 (N_12455,N_5439,N_5989);
or U12456 (N_12456,N_7815,N_2350);
nor U12457 (N_12457,N_1741,N_5490);
or U12458 (N_12458,N_5641,N_1542);
nor U12459 (N_12459,N_61,N_9451);
or U12460 (N_12460,N_9282,N_4603);
and U12461 (N_12461,N_3084,N_2235);
and U12462 (N_12462,N_5380,N_7497);
xnor U12463 (N_12463,N_6243,N_65);
xor U12464 (N_12464,N_6110,N_7628);
nand U12465 (N_12465,N_4959,N_2178);
or U12466 (N_12466,N_2558,N_2801);
and U12467 (N_12467,N_7441,N_9208);
xor U12468 (N_12468,N_387,N_6963);
or U12469 (N_12469,N_9616,N_27);
or U12470 (N_12470,N_8648,N_1846);
xor U12471 (N_12471,N_8611,N_485);
and U12472 (N_12472,N_7466,N_5786);
nand U12473 (N_12473,N_6601,N_6889);
and U12474 (N_12474,N_1169,N_185);
nand U12475 (N_12475,N_823,N_6737);
nor U12476 (N_12476,N_8011,N_8736);
xnor U12477 (N_12477,N_3193,N_2899);
xnor U12478 (N_12478,N_2153,N_7277);
or U12479 (N_12479,N_2991,N_5172);
nor U12480 (N_12480,N_2089,N_8368);
and U12481 (N_12481,N_7101,N_3920);
nor U12482 (N_12482,N_6609,N_8209);
nor U12483 (N_12483,N_5669,N_4728);
xnor U12484 (N_12484,N_1824,N_3147);
nand U12485 (N_12485,N_6954,N_9088);
xor U12486 (N_12486,N_5166,N_9574);
and U12487 (N_12487,N_1993,N_4014);
xor U12488 (N_12488,N_5848,N_6389);
nor U12489 (N_12489,N_924,N_9484);
nor U12490 (N_12490,N_7443,N_9076);
and U12491 (N_12491,N_3279,N_3419);
and U12492 (N_12492,N_4985,N_9783);
and U12493 (N_12493,N_175,N_1009);
and U12494 (N_12494,N_9863,N_3183);
xnor U12495 (N_12495,N_468,N_9254);
nor U12496 (N_12496,N_873,N_4049);
xnor U12497 (N_12497,N_1301,N_3060);
xor U12498 (N_12498,N_2989,N_9301);
or U12499 (N_12499,N_3528,N_7964);
xor U12500 (N_12500,N_1123,N_4100);
and U12501 (N_12501,N_8309,N_9101);
nor U12502 (N_12502,N_8147,N_7066);
and U12503 (N_12503,N_4359,N_9024);
and U12504 (N_12504,N_2995,N_8959);
or U12505 (N_12505,N_9107,N_4492);
nand U12506 (N_12506,N_6819,N_9949);
nor U12507 (N_12507,N_8057,N_9971);
nand U12508 (N_12508,N_8074,N_3465);
xor U12509 (N_12509,N_4637,N_1062);
nor U12510 (N_12510,N_2797,N_6435);
nand U12511 (N_12511,N_2817,N_4179);
nor U12512 (N_12512,N_8258,N_1212);
xnor U12513 (N_12513,N_3474,N_7350);
or U12514 (N_12514,N_2193,N_3558);
or U12515 (N_12515,N_3539,N_1324);
and U12516 (N_12516,N_1131,N_7829);
and U12517 (N_12517,N_4470,N_6037);
or U12518 (N_12518,N_5461,N_4883);
xor U12519 (N_12519,N_5765,N_3626);
or U12520 (N_12520,N_4907,N_6133);
xnor U12521 (N_12521,N_6545,N_6873);
and U12522 (N_12522,N_2749,N_6491);
nand U12523 (N_12523,N_1066,N_8472);
nand U12524 (N_12524,N_9731,N_8500);
nor U12525 (N_12525,N_7848,N_3889);
and U12526 (N_12526,N_1723,N_8961);
nand U12527 (N_12527,N_4513,N_8051);
and U12528 (N_12528,N_3478,N_3460);
nand U12529 (N_12529,N_7626,N_972);
nor U12530 (N_12530,N_2062,N_5751);
xnor U12531 (N_12531,N_6408,N_9943);
nand U12532 (N_12532,N_5970,N_2740);
nor U12533 (N_12533,N_7915,N_2902);
and U12534 (N_12534,N_5305,N_2475);
nor U12535 (N_12535,N_4060,N_3745);
nor U12536 (N_12536,N_2301,N_700);
xor U12537 (N_12537,N_9997,N_174);
nor U12538 (N_12538,N_266,N_6448);
or U12539 (N_12539,N_7125,N_2263);
and U12540 (N_12540,N_9984,N_6975);
xor U12541 (N_12541,N_6216,N_3681);
nor U12542 (N_12542,N_8807,N_8099);
xor U12543 (N_12543,N_8694,N_7270);
xor U12544 (N_12544,N_3207,N_5228);
nand U12545 (N_12545,N_9953,N_7129);
xor U12546 (N_12546,N_5445,N_4386);
nand U12547 (N_12547,N_769,N_3585);
nand U12548 (N_12548,N_1055,N_5872);
xor U12549 (N_12549,N_6843,N_2284);
or U12550 (N_12550,N_9350,N_3748);
nand U12551 (N_12551,N_8734,N_3578);
or U12552 (N_12552,N_1163,N_1181);
nor U12553 (N_12553,N_7292,N_2858);
xnor U12554 (N_12554,N_4244,N_631);
nor U12555 (N_12555,N_3364,N_2660);
nand U12556 (N_12556,N_4237,N_2622);
nor U12557 (N_12557,N_77,N_8321);
nor U12558 (N_12558,N_1097,N_6334);
nor U12559 (N_12559,N_3511,N_5554);
nor U12560 (N_12560,N_7754,N_4061);
xor U12561 (N_12561,N_3913,N_1461);
or U12562 (N_12562,N_2945,N_481);
nand U12563 (N_12563,N_5251,N_970);
xor U12564 (N_12564,N_9412,N_3651);
xor U12565 (N_12565,N_217,N_3441);
nor U12566 (N_12566,N_7932,N_2416);
or U12567 (N_12567,N_808,N_8113);
xor U12568 (N_12568,N_8859,N_9564);
and U12569 (N_12569,N_6171,N_8990);
nor U12570 (N_12570,N_6212,N_4171);
xnor U12571 (N_12571,N_1226,N_9457);
or U12572 (N_12572,N_5313,N_424);
nor U12573 (N_12573,N_7434,N_9865);
or U12574 (N_12574,N_7029,N_4515);
nand U12575 (N_12575,N_2963,N_5356);
nor U12576 (N_12576,N_732,N_5390);
nand U12577 (N_12577,N_6401,N_1424);
nor U12578 (N_12578,N_5702,N_7306);
and U12579 (N_12579,N_4993,N_3191);
nor U12580 (N_12580,N_5510,N_859);
nand U12581 (N_12581,N_426,N_5059);
nor U12582 (N_12582,N_8690,N_7874);
or U12583 (N_12583,N_8144,N_2559);
nor U12584 (N_12584,N_5803,N_5423);
or U12585 (N_12585,N_2315,N_7166);
and U12586 (N_12586,N_3609,N_6339);
and U12587 (N_12587,N_1178,N_4);
and U12588 (N_12588,N_4284,N_871);
xor U12589 (N_12589,N_3595,N_7075);
and U12590 (N_12590,N_4318,N_4604);
nor U12591 (N_12591,N_1615,N_5634);
nand U12592 (N_12592,N_8635,N_8677);
nand U12593 (N_12593,N_7348,N_6458);
nor U12594 (N_12594,N_9261,N_7343);
nand U12595 (N_12595,N_2847,N_8752);
xor U12596 (N_12596,N_2200,N_5608);
nand U12597 (N_12597,N_5854,N_1365);
and U12598 (N_12598,N_1467,N_8708);
nor U12599 (N_12599,N_8103,N_8250);
and U12600 (N_12600,N_8628,N_5835);
xor U12601 (N_12601,N_4139,N_367);
xnor U12602 (N_12602,N_7061,N_889);
and U12603 (N_12603,N_3201,N_8986);
xnor U12604 (N_12604,N_7577,N_7531);
nand U12605 (N_12605,N_838,N_2449);
and U12606 (N_12606,N_6987,N_5689);
and U12607 (N_12607,N_8429,N_6914);
xnor U12608 (N_12608,N_6348,N_3265);
nor U12609 (N_12609,N_1789,N_2822);
nor U12610 (N_12610,N_9300,N_5938);
and U12611 (N_12611,N_1455,N_8936);
or U12612 (N_12612,N_2850,N_6074);
or U12613 (N_12613,N_2711,N_8243);
xor U12614 (N_12614,N_2373,N_8982);
and U12615 (N_12615,N_5975,N_9129);
nor U12616 (N_12616,N_8365,N_2390);
nor U12617 (N_12617,N_6573,N_9542);
and U12618 (N_12618,N_3556,N_5139);
and U12619 (N_12619,N_4200,N_8972);
nor U12620 (N_12620,N_2258,N_5388);
nand U12621 (N_12621,N_3600,N_4919);
nand U12622 (N_12622,N_8764,N_2002);
and U12623 (N_12623,N_9203,N_7377);
nand U12624 (N_12624,N_2640,N_9570);
nand U12625 (N_12625,N_6376,N_5191);
or U12626 (N_12626,N_5552,N_7624);
and U12627 (N_12627,N_4769,N_76);
xnor U12628 (N_12628,N_4212,N_3241);
or U12629 (N_12629,N_1915,N_5398);
nand U12630 (N_12630,N_7994,N_5529);
nor U12631 (N_12631,N_2161,N_8772);
nor U12632 (N_12632,N_7701,N_3244);
xnor U12633 (N_12633,N_5222,N_7502);
or U12634 (N_12634,N_1118,N_8004);
or U12635 (N_12635,N_3588,N_7705);
xor U12636 (N_12636,N_7765,N_7589);
nand U12637 (N_12637,N_799,N_310);
nand U12638 (N_12638,N_774,N_7786);
and U12639 (N_12639,N_9844,N_5748);
nor U12640 (N_12640,N_4344,N_5379);
or U12641 (N_12641,N_1572,N_8925);
and U12642 (N_12642,N_8988,N_9546);
nor U12643 (N_12643,N_3325,N_7667);
xor U12644 (N_12644,N_646,N_6442);
nand U12645 (N_12645,N_9824,N_7838);
nor U12646 (N_12646,N_2171,N_4888);
or U12647 (N_12647,N_3744,N_7520);
xor U12648 (N_12648,N_8073,N_6494);
or U12649 (N_12649,N_2909,N_2973);
or U12650 (N_12650,N_134,N_7299);
nor U12651 (N_12651,N_8693,N_5074);
nand U12652 (N_12652,N_6200,N_3560);
and U12653 (N_12653,N_9317,N_3864);
nand U12654 (N_12654,N_761,N_350);
xnor U12655 (N_12655,N_5184,N_2299);
nand U12656 (N_12656,N_1241,N_51);
xor U12657 (N_12657,N_2352,N_6919);
and U12658 (N_12658,N_4530,N_4784);
and U12659 (N_12659,N_3212,N_620);
nor U12660 (N_12660,N_7571,N_6977);
and U12661 (N_12661,N_6383,N_5477);
nor U12662 (N_12662,N_1082,N_4038);
or U12663 (N_12663,N_2092,N_8675);
nand U12664 (N_12664,N_8190,N_392);
and U12665 (N_12665,N_8436,N_9898);
nor U12666 (N_12666,N_7865,N_816);
nor U12667 (N_12667,N_4183,N_3904);
nor U12668 (N_12668,N_6576,N_6674);
nor U12669 (N_12669,N_6673,N_6214);
or U12670 (N_12670,N_8952,N_5480);
nor U12671 (N_12671,N_2575,N_6087);
or U12672 (N_12672,N_9274,N_6404);
nor U12673 (N_12673,N_5374,N_4930);
and U12674 (N_12674,N_1280,N_8618);
nor U12675 (N_12675,N_8531,N_4054);
xnor U12676 (N_12676,N_5652,N_5909);
nor U12677 (N_12677,N_8948,N_3867);
and U12678 (N_12678,N_5962,N_3059);
nor U12679 (N_12679,N_9794,N_2971);
xnor U12680 (N_12680,N_8024,N_8162);
nor U12681 (N_12681,N_2098,N_8929);
xnor U12682 (N_12682,N_4842,N_3283);
or U12683 (N_12683,N_4865,N_2753);
or U12684 (N_12684,N_4690,N_7872);
and U12685 (N_12685,N_9122,N_5537);
or U12686 (N_12686,N_9770,N_5248);
nor U12687 (N_12687,N_368,N_8710);
nor U12688 (N_12688,N_8100,N_2302);
and U12689 (N_12689,N_8296,N_1151);
nor U12690 (N_12690,N_9224,N_5278);
and U12691 (N_12691,N_5413,N_2683);
or U12692 (N_12692,N_2751,N_5085);
nand U12693 (N_12693,N_1697,N_4193);
xnor U12694 (N_12694,N_3034,N_5732);
xnor U12695 (N_12695,N_2414,N_3717);
and U12696 (N_12696,N_1521,N_5276);
xnor U12697 (N_12697,N_6313,N_1957);
xor U12698 (N_12698,N_9378,N_8092);
nand U12699 (N_12699,N_2762,N_5680);
nor U12700 (N_12700,N_3910,N_410);
nor U12701 (N_12701,N_7495,N_130);
and U12702 (N_12702,N_8524,N_4791);
nor U12703 (N_12703,N_7536,N_6594);
or U12704 (N_12704,N_9163,N_5465);
xor U12705 (N_12705,N_4703,N_9491);
xnor U12706 (N_12706,N_5651,N_6048);
xnor U12707 (N_12707,N_2096,N_437);
nor U12708 (N_12708,N_3090,N_6672);
and U12709 (N_12709,N_7935,N_7071);
and U12710 (N_12710,N_4274,N_6402);
or U12711 (N_12711,N_87,N_2551);
nand U12712 (N_12712,N_4071,N_365);
nor U12713 (N_12713,N_617,N_1805);
nand U12714 (N_12714,N_8966,N_2877);
nand U12715 (N_12715,N_1364,N_1744);
nand U12716 (N_12716,N_6734,N_6017);
and U12717 (N_12717,N_1918,N_180);
xor U12718 (N_12718,N_6778,N_4785);
and U12719 (N_12719,N_9086,N_5358);
or U12720 (N_12720,N_8020,N_984);
or U12721 (N_12721,N_8093,N_4424);
and U12722 (N_12722,N_3935,N_6735);
nand U12723 (N_12723,N_8407,N_9169);
nor U12724 (N_12724,N_3975,N_4081);
or U12725 (N_12725,N_5807,N_2512);
xnor U12726 (N_12726,N_318,N_1457);
and U12727 (N_12727,N_6140,N_2981);
or U12728 (N_12728,N_6511,N_4548);
or U12729 (N_12729,N_5351,N_4966);
nand U12730 (N_12730,N_7756,N_7507);
nor U12731 (N_12731,N_7217,N_8712);
nand U12732 (N_12732,N_9497,N_3235);
nand U12733 (N_12733,N_4657,N_9787);
nor U12734 (N_12734,N_8589,N_2759);
and U12735 (N_12735,N_4285,N_5793);
nand U12736 (N_12736,N_7264,N_1971);
nor U12737 (N_12737,N_6028,N_8820);
xor U12738 (N_12738,N_1897,N_6863);
nor U12739 (N_12739,N_9507,N_3335);
nand U12740 (N_12740,N_7665,N_982);
nor U12741 (N_12741,N_9171,N_7992);
nand U12742 (N_12742,N_4029,N_7063);
xnor U12743 (N_12743,N_2502,N_5410);
nand U12744 (N_12744,N_9518,N_609);
and U12745 (N_12745,N_8563,N_9463);
nand U12746 (N_12746,N_7367,N_6593);
or U12747 (N_12747,N_8373,N_4384);
or U12748 (N_12748,N_8981,N_7447);
nor U12749 (N_12749,N_9962,N_4414);
nor U12750 (N_12750,N_2544,N_9370);
or U12751 (N_12751,N_6472,N_2026);
nor U12752 (N_12752,N_3413,N_2409);
and U12753 (N_12753,N_4673,N_6946);
nand U12754 (N_12754,N_8667,N_2542);
xnor U12755 (N_12755,N_9483,N_994);
or U12756 (N_12756,N_950,N_1775);
nor U12757 (N_12757,N_3225,N_1483);
nand U12758 (N_12758,N_5010,N_4903);
nor U12759 (N_12759,N_3818,N_9561);
or U12760 (N_12760,N_9360,N_2600);
nand U12761 (N_12761,N_259,N_7746);
or U12762 (N_12762,N_6159,N_7453);
xnor U12763 (N_12763,N_186,N_7395);
nand U12764 (N_12764,N_1111,N_1990);
or U12765 (N_12765,N_8767,N_2104);
and U12766 (N_12766,N_6925,N_6265);
nor U12767 (N_12767,N_8291,N_1873);
xor U12768 (N_12768,N_4988,N_8901);
nor U12769 (N_12769,N_1078,N_615);
and U12770 (N_12770,N_3436,N_1339);
nor U12771 (N_12771,N_135,N_286);
or U12772 (N_12772,N_2472,N_7319);
xnor U12773 (N_12773,N_4322,N_9610);
nand U12774 (N_12774,N_945,N_278);
nor U12775 (N_12775,N_4080,N_8808);
nor U12776 (N_12776,N_103,N_9691);
nor U12777 (N_12777,N_3015,N_6196);
and U12778 (N_12778,N_749,N_7159);
xnor U12779 (N_12779,N_1732,N_6181);
or U12780 (N_12780,N_2855,N_5884);
or U12781 (N_12781,N_9519,N_7697);
nor U12782 (N_12782,N_9196,N_24);
xnor U12783 (N_12783,N_7525,N_59);
xor U12784 (N_12784,N_66,N_4480);
xnor U12785 (N_12785,N_3339,N_4224);
nand U12786 (N_12786,N_7302,N_9125);
nand U12787 (N_12787,N_2219,N_983);
or U12788 (N_12788,N_6829,N_5001);
or U12789 (N_12789,N_3383,N_3707);
nand U12790 (N_12790,N_8848,N_5877);
or U12791 (N_12791,N_7072,N_8509);
xor U12792 (N_12792,N_8333,N_9805);
nand U12793 (N_12793,N_8352,N_9711);
nand U12794 (N_12794,N_8148,N_5401);
and U12795 (N_12795,N_4760,N_8593);
and U12796 (N_12796,N_4969,N_8235);
nand U12797 (N_12797,N_7023,N_2629);
nand U12798 (N_12798,N_2103,N_9795);
nand U12799 (N_12799,N_7087,N_9202);
xor U12800 (N_12800,N_3385,N_6556);
nand U12801 (N_12801,N_6092,N_5776);
nor U12802 (N_12802,N_3405,N_222);
xnor U12803 (N_12803,N_9021,N_791);
and U12804 (N_12804,N_6157,N_6756);
xor U12805 (N_12805,N_4808,N_560);
nand U12806 (N_12806,N_2107,N_6226);
nand U12807 (N_12807,N_5967,N_3484);
and U12808 (N_12808,N_9938,N_4302);
nor U12809 (N_12809,N_2591,N_1693);
nand U12810 (N_12810,N_8175,N_6607);
and U12811 (N_12811,N_4598,N_3750);
nor U12812 (N_12812,N_7272,N_2534);
and U12813 (N_12813,N_8305,N_4746);
nand U12814 (N_12814,N_8186,N_8554);
xnor U12815 (N_12815,N_6177,N_50);
xnor U12816 (N_12816,N_3019,N_2662);
and U12817 (N_12817,N_6369,N_5216);
and U12818 (N_12818,N_4520,N_1046);
xor U12819 (N_12819,N_478,N_1592);
xnor U12820 (N_12820,N_171,N_125);
nand U12821 (N_12821,N_2,N_7963);
nand U12822 (N_12822,N_2467,N_655);
or U12823 (N_12823,N_3610,N_7614);
nand U12824 (N_12824,N_1550,N_2637);
nand U12825 (N_12825,N_1018,N_7410);
or U12826 (N_12826,N_1043,N_836);
and U12827 (N_12827,N_196,N_2958);
nor U12828 (N_12828,N_2789,N_3480);
or U12829 (N_12829,N_7512,N_9720);
xor U12830 (N_12830,N_9732,N_9801);
nand U12831 (N_12831,N_4511,N_6730);
and U12832 (N_12832,N_8204,N_9956);
or U12833 (N_12833,N_3382,N_1666);
xnor U12834 (N_12834,N_746,N_7191);
xnor U12835 (N_12835,N_2197,N_1718);
nand U12836 (N_12836,N_7035,N_1848);
nand U12837 (N_12837,N_8141,N_8762);
xnor U12838 (N_12838,N_3763,N_8142);
and U12839 (N_12839,N_1362,N_7670);
or U12840 (N_12840,N_109,N_3106);
or U12841 (N_12841,N_6318,N_5307);
and U12842 (N_12842,N_9618,N_2024);
and U12843 (N_12843,N_1953,N_1639);
xor U12844 (N_12844,N_4027,N_7080);
and U12845 (N_12845,N_4628,N_618);
or U12846 (N_12846,N_9612,N_9066);
xor U12847 (N_12847,N_1920,N_4058);
nor U12848 (N_12848,N_82,N_2503);
or U12849 (N_12849,N_5412,N_6173);
xnor U12850 (N_12850,N_1626,N_7372);
nor U12851 (N_12851,N_8845,N_9030);
nand U12852 (N_12852,N_5119,N_477);
and U12853 (N_12853,N_5328,N_9905);
nand U12854 (N_12854,N_291,N_2722);
nor U12855 (N_12855,N_2992,N_1317);
nand U12856 (N_12856,N_2304,N_6263);
xnor U12857 (N_12857,N_3599,N_4803);
or U12858 (N_12858,N_4862,N_2923);
or U12859 (N_12859,N_9914,N_9221);
and U12860 (N_12860,N_8252,N_6454);
and U12861 (N_12861,N_9670,N_7250);
nand U12862 (N_12862,N_5271,N_9164);
or U12863 (N_12863,N_4625,N_1832);
and U12864 (N_12864,N_5561,N_1206);
xnor U12865 (N_12865,N_726,N_9504);
or U12866 (N_12866,N_8947,N_1113);
xnor U12867 (N_12867,N_8917,N_8157);
and U12868 (N_12868,N_9730,N_1349);
or U12869 (N_12869,N_242,N_3155);
nand U12870 (N_12870,N_7553,N_3795);
or U12871 (N_12871,N_3030,N_3048);
and U12872 (N_12872,N_7954,N_4701);
or U12873 (N_12873,N_934,N_8777);
nand U12874 (N_12874,N_6270,N_6514);
xor U12875 (N_12875,N_6052,N_1858);
or U12876 (N_12876,N_3739,N_6931);
nand U12877 (N_12877,N_2135,N_4357);
xnor U12878 (N_12878,N_8428,N_6569);
and U12879 (N_12879,N_1402,N_9754);
or U12880 (N_12880,N_6024,N_7151);
nor U12881 (N_12881,N_9643,N_7389);
nor U12882 (N_12882,N_3756,N_292);
or U12883 (N_12883,N_4795,N_4682);
or U12884 (N_12884,N_5523,N_4252);
nand U12885 (N_12885,N_7295,N_6988);
nor U12886 (N_12886,N_8782,N_5306);
and U12887 (N_12887,N_2129,N_4495);
or U12888 (N_12888,N_3430,N_2251);
or U12889 (N_12889,N_3188,N_8501);
nand U12890 (N_12890,N_6870,N_1037);
xnor U12891 (N_12891,N_147,N_3394);
nor U12892 (N_12892,N_363,N_7445);
xnor U12893 (N_12893,N_3328,N_4591);
nor U12894 (N_12894,N_9399,N_294);
nand U12895 (N_12895,N_3517,N_2950);
nor U12896 (N_12896,N_5824,N_4093);
nor U12897 (N_12897,N_811,N_8638);
or U12898 (N_12898,N_500,N_9932);
or U12899 (N_12899,N_4020,N_5724);
nand U12900 (N_12900,N_640,N_6739);
or U12901 (N_12901,N_9860,N_6845);
or U12902 (N_12902,N_9212,N_330);
nor U12903 (N_12903,N_3077,N_2402);
xor U12904 (N_12904,N_5855,N_1637);
xnor U12905 (N_12905,N_8766,N_8001);
nor U12906 (N_12906,N_5220,N_8115);
or U12907 (N_12907,N_2112,N_2494);
nor U12908 (N_12908,N_4797,N_1421);
or U12909 (N_12909,N_3769,N_9540);
nand U12910 (N_12910,N_376,N_267);
nand U12911 (N_12911,N_5623,N_4524);
nor U12912 (N_12912,N_5943,N_3857);
xor U12913 (N_12913,N_8843,N_9302);
and U12914 (N_12914,N_5516,N_8310);
or U12915 (N_12915,N_8129,N_3515);
or U12916 (N_12916,N_2888,N_6913);
xnor U12917 (N_12917,N_2030,N_158);
and U12918 (N_12918,N_7906,N_8170);
and U12919 (N_12919,N_5912,N_2504);
nor U12920 (N_12920,N_206,N_8274);
nor U12921 (N_12921,N_7494,N_1416);
xor U12922 (N_12922,N_7492,N_1440);
nand U12923 (N_12923,N_75,N_1965);
nand U12924 (N_12924,N_7951,N_3153);
nor U12925 (N_12925,N_9257,N_4958);
xor U12926 (N_12926,N_91,N_1682);
and U12927 (N_12927,N_1182,N_8262);
xnor U12928 (N_12928,N_4312,N_7014);
or U12929 (N_12929,N_2571,N_2195);
xor U12930 (N_12930,N_1684,N_6706);
nor U12931 (N_12931,N_8882,N_2450);
or U12932 (N_12932,N_5182,N_5416);
nand U12933 (N_12933,N_9324,N_1940);
or U12934 (N_12934,N_5284,N_3645);
nand U12935 (N_12935,N_7136,N_1219);
nor U12936 (N_12936,N_2952,N_613);
nand U12937 (N_12937,N_235,N_7717);
nand U12938 (N_12938,N_8637,N_802);
xnor U12939 (N_12939,N_2541,N_312);
or U12940 (N_12940,N_9993,N_9034);
or U12941 (N_12941,N_6517,N_9503);
xor U12942 (N_12942,N_9111,N_43);
nor U12943 (N_12943,N_4773,N_9735);
nand U12944 (N_12944,N_4374,N_4177);
nor U12945 (N_12945,N_2593,N_4348);
xor U12946 (N_12946,N_920,N_5127);
or U12947 (N_12947,N_5396,N_9611);
nand U12948 (N_12948,N_6311,N_9278);
nor U12949 (N_12949,N_7409,N_6225);
and U12950 (N_12950,N_514,N_7645);
and U12951 (N_12951,N_4646,N_6994);
and U12952 (N_12952,N_8143,N_6854);
nor U12953 (N_12953,N_3157,N_6300);
and U12954 (N_12954,N_6146,N_4545);
nor U12955 (N_12955,N_8923,N_2965);
or U12956 (N_12956,N_2556,N_6089);
nand U12957 (N_12957,N_4602,N_742);
and U12958 (N_12958,N_3655,N_3110);
and U12959 (N_12959,N_2787,N_9657);
nand U12960 (N_12960,N_6490,N_3052);
or U12961 (N_12961,N_2483,N_4940);
nand U12962 (N_12962,N_6990,N_1715);
or U12963 (N_12963,N_3463,N_671);
and U12964 (N_12964,N_9443,N_7888);
and U12965 (N_12965,N_3596,N_5093);
or U12966 (N_12966,N_4533,N_7598);
nor U12967 (N_12967,N_9476,N_119);
or U12968 (N_12968,N_3799,N_3809);
xnor U12969 (N_12969,N_3602,N_3611);
and U12970 (N_12970,N_7213,N_9468);
xnor U12971 (N_12971,N_1492,N_6733);
and U12972 (N_12972,N_8935,N_5839);
xor U12973 (N_12973,N_8870,N_1215);
nand U12974 (N_12974,N_9716,N_5789);
nand U12975 (N_12975,N_1020,N_5399);
nand U12976 (N_12976,N_8302,N_3895);
nor U12977 (N_12977,N_6007,N_7123);
or U12978 (N_12978,N_7661,N_3310);
and U12979 (N_12979,N_4075,N_1594);
nand U12980 (N_12980,N_6010,N_74);
xnor U12981 (N_12981,N_8068,N_447);
nand U12982 (N_12982,N_8341,N_6888);
nor U12983 (N_12983,N_1278,N_8237);
xor U12984 (N_12984,N_6904,N_3845);
or U12985 (N_12985,N_9573,N_3683);
nor U12986 (N_12986,N_7342,N_513);
xnor U12987 (N_12987,N_7266,N_8443);
or U12988 (N_12988,N_4976,N_8224);
nand U12989 (N_12989,N_6235,N_4136);
nand U12990 (N_12990,N_8165,N_6122);
or U12991 (N_12991,N_5818,N_3271);
and U12992 (N_12992,N_4488,N_2456);
and U12993 (N_12993,N_2620,N_4372);
or U12994 (N_12994,N_9718,N_8469);
nor U12995 (N_12995,N_4114,N_6444);
or U12996 (N_12996,N_8821,N_6329);
and U12997 (N_12997,N_8878,N_6871);
xnor U12998 (N_12998,N_779,N_5442);
xor U12999 (N_12999,N_5237,N_7044);
or U13000 (N_13000,N_3694,N_9533);
or U13001 (N_13001,N_2910,N_6895);
nand U13002 (N_13002,N_9903,N_3656);
or U13003 (N_13003,N_4942,N_6014);
and U13004 (N_13004,N_2837,N_8980);
nand U13005 (N_13005,N_6266,N_3540);
xor U13006 (N_13006,N_6482,N_3727);
and U13007 (N_13007,N_3902,N_2818);
and U13008 (N_13008,N_6425,N_4024);
or U13009 (N_13009,N_5072,N_2823);
and U13010 (N_13010,N_515,N_7855);
nand U13011 (N_13011,N_7432,N_2555);
xnor U13012 (N_13012,N_9387,N_6247);
nand U13013 (N_13013,N_6704,N_1296);
nor U13014 (N_13014,N_2573,N_9157);
xor U13015 (N_13015,N_4261,N_2979);
nand U13016 (N_13016,N_7847,N_224);
nor U13017 (N_13017,N_4445,N_2680);
or U13018 (N_13018,N_9039,N_41);
nand U13019 (N_13019,N_2978,N_916);
nor U13020 (N_13020,N_7440,N_1375);
nor U13021 (N_13021,N_2916,N_2151);
nand U13022 (N_13022,N_7547,N_8463);
nor U13023 (N_13023,N_4718,N_1706);
nand U13024 (N_13024,N_7407,N_2260);
nand U13025 (N_13025,N_5238,N_6044);
xor U13026 (N_13026,N_3458,N_272);
nand U13027 (N_13027,N_3455,N_7253);
nand U13028 (N_13028,N_7174,N_9715);
nand U13029 (N_13029,N_6056,N_2042);
nand U13030 (N_13030,N_7199,N_3372);
and U13031 (N_13031,N_7206,N_1830);
nor U13032 (N_13032,N_308,N_399);
xnor U13033 (N_13033,N_3901,N_1144);
xnor U13034 (N_13034,N_9349,N_3519);
and U13035 (N_13035,N_2777,N_8203);
xor U13036 (N_13036,N_2127,N_8216);
and U13037 (N_13037,N_3776,N_2406);
xnor U13038 (N_13038,N_2668,N_1790);
xnor U13039 (N_13039,N_8372,N_6430);
nor U13040 (N_13040,N_5518,N_8640);
nor U13041 (N_13041,N_3995,N_4273);
and U13042 (N_13042,N_249,N_2203);
xor U13043 (N_13043,N_4220,N_3161);
and U13044 (N_13044,N_2173,N_1886);
or U13045 (N_13045,N_5221,N_3438);
and U13046 (N_13046,N_6175,N_8320);
or U13047 (N_13047,N_2346,N_5178);
xor U13048 (N_13048,N_890,N_8423);
or U13049 (N_13049,N_5,N_7767);
xnor U13050 (N_13050,N_9853,N_5459);
nand U13051 (N_13051,N_6034,N_73);
and U13052 (N_13052,N_1930,N_1655);
or U13053 (N_13053,N_9054,N_7195);
xor U13054 (N_13054,N_7124,N_6769);
xor U13055 (N_13055,N_595,N_1613);
xor U13056 (N_13056,N_9365,N_92);
nand U13057 (N_13057,N_8768,N_6267);
and U13058 (N_13058,N_2763,N_2829);
nor U13059 (N_13059,N_9571,N_569);
xor U13060 (N_13060,N_6824,N_733);
nand U13061 (N_13061,N_5430,N_7107);
or U13062 (N_13062,N_5083,N_8122);
and U13063 (N_13063,N_128,N_3673);
and U13064 (N_13064,N_3293,N_2500);
or U13065 (N_13065,N_638,N_9874);
nand U13066 (N_13066,N_2791,N_3697);
or U13067 (N_13067,N_7269,N_9840);
and U13068 (N_13068,N_6213,N_8330);
nor U13069 (N_13069,N_7934,N_7314);
xor U13070 (N_13070,N_4493,N_9144);
xor U13071 (N_13071,N_4960,N_9004);
or U13072 (N_13072,N_5656,N_5925);
and U13073 (N_13073,N_546,N_8207);
and U13074 (N_13074,N_3928,N_978);
nor U13075 (N_13075,N_4719,N_2216);
xnor U13076 (N_13076,N_1154,N_8375);
xor U13077 (N_13077,N_3227,N_5653);
nor U13078 (N_13078,N_2453,N_1675);
or U13079 (N_13079,N_8751,N_5790);
xor U13080 (N_13080,N_6153,N_3930);
nand U13081 (N_13081,N_3822,N_8078);
and U13082 (N_13082,N_1431,N_4176);
or U13083 (N_13083,N_2708,N_1504);
or U13084 (N_13084,N_7740,N_2827);
or U13085 (N_13085,N_9069,N_7486);
and U13086 (N_13086,N_9575,N_8749);
nand U13087 (N_13087,N_9906,N_4000);
xnor U13088 (N_13088,N_5199,N_7835);
nor U13089 (N_13089,N_6372,N_676);
xor U13090 (N_13090,N_5067,N_9978);
or U13091 (N_13091,N_7362,N_4744);
nor U13092 (N_13092,N_4939,N_6155);
xnor U13093 (N_13093,N_2448,N_4423);
or U13094 (N_13094,N_9380,N_9606);
or U13095 (N_13095,N_7820,N_4113);
and U13096 (N_13096,N_538,N_2903);
and U13097 (N_13097,N_6546,N_8765);
or U13098 (N_13098,N_7265,N_4830);
nand U13099 (N_13099,N_3579,N_4088);
xnor U13100 (N_13100,N_1474,N_4630);
xor U13101 (N_13101,N_1961,N_8110);
xor U13102 (N_13102,N_3709,N_731);
and U13103 (N_13103,N_9321,N_2331);
and U13104 (N_13104,N_417,N_1704);
or U13105 (N_13105,N_9112,N_9856);
or U13106 (N_13106,N_8678,N_3958);
nand U13107 (N_13107,N_265,N_8220);
xor U13108 (N_13108,N_1155,N_8958);
nand U13109 (N_13109,N_6388,N_3536);
nand U13110 (N_13110,N_7263,N_3199);
xnor U13111 (N_13111,N_6757,N_630);
nand U13112 (N_13112,N_3632,N_6304);
nor U13113 (N_13113,N_9424,N_4092);
nand U13114 (N_13114,N_4425,N_3761);
nor U13115 (N_13115,N_5978,N_7190);
xor U13116 (N_13116,N_6644,N_482);
nor U13117 (N_13117,N_9527,N_4199);
nor U13118 (N_13118,N_2093,N_414);
xnor U13119 (N_13119,N_3347,N_3027);
and U13120 (N_13120,N_4859,N_8661);
nand U13121 (N_13121,N_880,N_2488);
nor U13122 (N_13122,N_2441,N_4848);
nand U13123 (N_13123,N_3269,N_7122);
or U13124 (N_13124,N_6202,N_5600);
or U13125 (N_13125,N_7728,N_1823);
nand U13126 (N_13126,N_9676,N_2948);
or U13127 (N_13127,N_8163,N_3852);
nor U13128 (N_13128,N_9851,N_9589);
and U13129 (N_13129,N_9902,N_432);
or U13130 (N_13130,N_9960,N_3273);
and U13131 (N_13131,N_6702,N_6774);
or U13132 (N_13132,N_3282,N_7210);
or U13133 (N_13133,N_2778,N_7712);
or U13134 (N_13134,N_9781,N_2743);
nor U13135 (N_13135,N_2687,N_1334);
nor U13136 (N_13136,N_340,N_1602);
or U13137 (N_13137,N_7771,N_8953);
nor U13138 (N_13138,N_7032,N_9437);
nand U13139 (N_13139,N_9233,N_7451);
nand U13140 (N_13140,N_6439,N_9170);
and U13141 (N_13141,N_8483,N_5471);
xor U13142 (N_13142,N_7161,N_604);
and U13143 (N_13143,N_4468,N_7690);
xor U13144 (N_13144,N_4577,N_5342);
or U13145 (N_13145,N_8457,N_860);
nand U13146 (N_13146,N_7374,N_9318);
nor U13147 (N_13147,N_1925,N_5391);
xor U13148 (N_13148,N_8784,N_4729);
xor U13149 (N_13149,N_4589,N_1673);
or U13150 (N_13150,N_4649,N_7949);
or U13151 (N_13151,N_3937,N_3058);
nand U13152 (N_13152,N_5473,N_7153);
and U13153 (N_13153,N_7298,N_7511);
xnor U13154 (N_13154,N_8178,N_6340);
and U13155 (N_13155,N_7242,N_5593);
and U13156 (N_13156,N_2466,N_2404);
or U13157 (N_13157,N_7804,N_1906);
nor U13158 (N_13158,N_3069,N_9238);
nor U13159 (N_13159,N_1752,N_5964);
nor U13160 (N_13160,N_2184,N_3501);
nand U13161 (N_13161,N_8564,N_83);
or U13162 (N_13162,N_3779,N_3844);
and U13163 (N_13163,N_2140,N_7145);
or U13164 (N_13164,N_4375,N_2207);
nor U13165 (N_13165,N_3446,N_3529);
nor U13166 (N_13166,N_1261,N_6262);
or U13167 (N_13167,N_1072,N_6450);
and U13168 (N_13168,N_9402,N_1972);
nor U13169 (N_13169,N_4526,N_6341);
xnor U13170 (N_13170,N_9543,N_3729);
nand U13171 (N_13171,N_3170,N_8348);
nor U13172 (N_13172,N_1654,N_1032);
nand U13173 (N_13173,N_1121,N_1145);
nand U13174 (N_13174,N_3470,N_9435);
nor U13175 (N_13175,N_6716,N_8668);
and U13176 (N_13176,N_1227,N_4954);
nand U13177 (N_13177,N_1014,N_8774);
nor U13178 (N_13178,N_5781,N_9684);
nand U13179 (N_13179,N_8824,N_1150);
nor U13180 (N_13180,N_4032,N_1650);
nor U13181 (N_13181,N_9945,N_8239);
xnor U13182 (N_13182,N_3654,N_4532);
nor U13183 (N_13183,N_4394,N_7600);
and U13184 (N_13184,N_89,N_9909);
xnor U13185 (N_13185,N_4328,N_9924);
nand U13186 (N_13186,N_6967,N_5662);
nor U13187 (N_13187,N_7086,N_1106);
and U13188 (N_13188,N_453,N_3013);
nand U13189 (N_13189,N_7436,N_6942);
xnor U13190 (N_13190,N_7632,N_6446);
and U13191 (N_13191,N_3247,N_5609);
nor U13192 (N_13192,N_3177,N_2619);
or U13193 (N_13193,N_4807,N_3210);
xor U13194 (N_13194,N_4820,N_9704);
xnor U13195 (N_13195,N_301,N_4877);
and U13196 (N_13196,N_7669,N_4119);
nor U13197 (N_13197,N_3613,N_4403);
or U13198 (N_13198,N_5880,N_8371);
xnor U13199 (N_13199,N_7530,N_1256);
nor U13200 (N_13200,N_4499,N_170);
or U13201 (N_13201,N_5901,N_5164);
nand U13202 (N_13202,N_4787,N_1393);
xor U13203 (N_13203,N_738,N_6496);
nor U13204 (N_13204,N_7676,N_5069);
nor U13205 (N_13205,N_1214,N_4898);
nand U13206 (N_13206,N_5025,N_6743);
nor U13207 (N_13207,N_3168,N_5462);
nor U13208 (N_13208,N_2411,N_5618);
nor U13209 (N_13209,N_6933,N_5111);
and U13210 (N_13210,N_9108,N_3492);
nand U13211 (N_13211,N_2196,N_4521);
xor U13212 (N_13212,N_2742,N_5591);
nand U13213 (N_13213,N_6449,N_9664);
or U13214 (N_13214,N_3156,N_4338);
or U13215 (N_13215,N_3091,N_4566);
and U13216 (N_13216,N_449,N_4592);
xor U13217 (N_13217,N_1257,N_5957);
xnor U13218 (N_13218,N_9348,N_5549);
xor U13219 (N_13219,N_9081,N_1029);
xnor U13220 (N_13220,N_3195,N_5377);
or U13221 (N_13221,N_3768,N_5000);
and U13222 (N_13222,N_2842,N_8522);
and U13223 (N_13223,N_1868,N_4484);
and U13224 (N_13224,N_1128,N_7766);
xor U13225 (N_13225,N_4023,N_4950);
and U13226 (N_13226,N_7479,N_2757);
xnor U13227 (N_13227,N_1047,N_8408);
or U13228 (N_13228,N_5277,N_9693);
nor U13229 (N_13229,N_9205,N_6908);
and U13230 (N_13230,N_3236,N_4995);
or U13231 (N_13231,N_3393,N_4866);
nand U13232 (N_13232,N_3696,N_1463);
xnor U13233 (N_13233,N_6322,N_5830);
or U13234 (N_13234,N_8978,N_4656);
nand U13235 (N_13235,N_2420,N_9698);
nand U13236 (N_13236,N_9511,N_4553);
and U13237 (N_13237,N_8722,N_9194);
and U13238 (N_13238,N_2074,N_9607);
and U13239 (N_13239,N_3755,N_5140);
and U13240 (N_13240,N_6386,N_3841);
xnor U13241 (N_13241,N_7671,N_8145);
nand U13242 (N_13242,N_6082,N_4001);
nand U13243 (N_13243,N_6926,N_3886);
and U13244 (N_13244,N_9665,N_4354);
and U13245 (N_13245,N_2147,N_6131);
nand U13246 (N_13246,N_2755,N_2330);
nor U13247 (N_13247,N_9118,N_5331);
nor U13248 (N_13248,N_2339,N_5021);
nand U13249 (N_13249,N_2164,N_2761);
nor U13250 (N_13250,N_3125,N_2085);
and U13251 (N_13251,N_3057,N_9747);
xnor U13252 (N_13252,N_6782,N_1485);
xnor U13253 (N_13253,N_1662,N_756);
nand U13254 (N_13254,N_1687,N_8059);
and U13255 (N_13255,N_7986,N_4809);
xor U13256 (N_13256,N_9020,N_4609);
nand U13257 (N_13257,N_2117,N_2729);
nand U13258 (N_13258,N_9531,N_6469);
nand U13259 (N_13259,N_1756,N_7561);
and U13260 (N_13260,N_675,N_2437);
or U13261 (N_13261,N_3429,N_5543);
and U13262 (N_13262,N_1275,N_9762);
and U13263 (N_13263,N_4768,N_6353);
or U13264 (N_13264,N_519,N_6370);
nand U13265 (N_13265,N_3974,N_7975);
xnor U13266 (N_13266,N_4897,N_3663);
and U13267 (N_13267,N_5538,N_6333);
nand U13268 (N_13268,N_2931,N_9425);
nor U13269 (N_13269,N_7353,N_7400);
xor U13270 (N_13270,N_6732,N_4057);
nor U13271 (N_13271,N_1849,N_9174);
and U13272 (N_13272,N_2133,N_1444);
nor U13273 (N_13273,N_9509,N_7007);
and U13274 (N_13274,N_9073,N_2321);
xnor U13275 (N_13275,N_1652,N_6550);
nand U13276 (N_13276,N_5823,N_84);
xnor U13277 (N_13277,N_9577,N_397);
and U13278 (N_13278,N_3734,N_2533);
xnor U13279 (N_13279,N_1197,N_5772);
and U13280 (N_13280,N_2673,N_7768);
or U13281 (N_13281,N_1096,N_5076);
nand U13282 (N_13282,N_290,N_9562);
nand U13283 (N_13283,N_8937,N_8938);
and U13284 (N_13284,N_7617,N_4426);
nor U13285 (N_13285,N_585,N_7172);
nor U13286 (N_13286,N_5073,N_9319);
nand U13287 (N_13287,N_5168,N_4970);
or U13288 (N_13288,N_6784,N_3552);
or U13289 (N_13289,N_5541,N_8136);
or U13290 (N_13290,N_1458,N_7681);
or U13291 (N_13291,N_1895,N_1168);
or U13292 (N_13292,N_6636,N_189);
and U13293 (N_13293,N_8511,N_2122);
xor U13294 (N_13294,N_7931,N_3159);
xnor U13295 (N_13295,N_6640,N_745);
and U13296 (N_13296,N_7347,N_6659);
or U13297 (N_13297,N_8875,N_2175);
nand U13298 (N_13298,N_5769,N_2348);
nand U13299 (N_13299,N_299,N_5312);
nand U13300 (N_13300,N_1271,N_8029);
xnor U13301 (N_13301,N_416,N_4697);
xnor U13302 (N_13302,N_3338,N_4227);
or U13303 (N_13303,N_8127,N_2436);
nand U13304 (N_13304,N_5590,N_8860);
nand U13305 (N_13305,N_9614,N_1695);
xor U13306 (N_13306,N_440,N_703);
nor U13307 (N_13307,N_3587,N_3513);
nor U13308 (N_13308,N_9897,N_359);
and U13309 (N_13309,N_5426,N_1817);
xnor U13310 (N_13310,N_6285,N_5979);
nor U13311 (N_13311,N_597,N_1671);
nand U13312 (N_13312,N_4280,N_4779);
and U13313 (N_13313,N_3862,N_4314);
nor U13314 (N_13314,N_3964,N_3444);
nand U13315 (N_13315,N_1847,N_6708);
and U13316 (N_13316,N_4825,N_6551);
xnor U13317 (N_13317,N_3843,N_1085);
and U13318 (N_13318,N_4853,N_2779);
nand U13319 (N_13319,N_2509,N_5876);
and U13320 (N_13320,N_1528,N_151);
nor U13321 (N_13321,N_635,N_7736);
nand U13322 (N_13322,N_7947,N_721);
nand U13323 (N_13323,N_3006,N_4149);
xor U13324 (N_13324,N_9048,N_3856);
nor U13325 (N_13325,N_3355,N_4086);
or U13326 (N_13326,N_1685,N_5924);
and U13327 (N_13327,N_2043,N_1189);
and U13328 (N_13328,N_380,N_3801);
nor U13329 (N_13329,N_8810,N_1115);
or U13330 (N_13330,N_13,N_4387);
xor U13331 (N_13331,N_7278,N_6763);
and U13332 (N_13332,N_5784,N_8529);
nand U13333 (N_13333,N_9947,N_4039);
nand U13334 (N_13334,N_4696,N_9271);
xnor U13335 (N_13335,N_8897,N_2904);
or U13336 (N_13336,N_7042,N_8579);
nand U13337 (N_13337,N_9937,N_9719);
nand U13338 (N_13338,N_1916,N_3971);
nor U13339 (N_13339,N_6166,N_8510);
nor U13340 (N_13340,N_1073,N_5252);
xnor U13341 (N_13341,N_4441,N_7309);
xor U13342 (N_13342,N_8201,N_894);
nor U13343 (N_13343,N_3905,N_9265);
and U13344 (N_13344,N_7724,N_6473);
nand U13345 (N_13345,N_2994,N_6385);
xor U13346 (N_13346,N_6586,N_1425);
or U13347 (N_13347,N_5806,N_9056);
nor U13348 (N_13348,N_256,N_7170);
nor U13349 (N_13349,N_991,N_8069);
xor U13350 (N_13350,N_1879,N_7711);
and U13351 (N_13351,N_7297,N_3634);
xor U13352 (N_13352,N_5488,N_2090);
and U13353 (N_13353,N_9119,N_7516);
xor U13354 (N_13354,N_1892,N_503);
nor U13355 (N_13355,N_2136,N_1508);
and U13356 (N_13356,N_6598,N_7984);
or U13357 (N_13357,N_4458,N_9026);
and U13358 (N_13358,N_1535,N_5860);
and U13359 (N_13359,N_8757,N_4847);
and U13360 (N_13360,N_3053,N_7286);
xor U13361 (N_13361,N_3733,N_2974);
nand U13362 (N_13362,N_1648,N_2515);
nand U13363 (N_13363,N_490,N_6233);
xnor U13364 (N_13364,N_1419,N_9662);
xnor U13365 (N_13365,N_7083,N_5607);
nand U13366 (N_13366,N_4525,N_8686);
xor U13367 (N_13367,N_8738,N_6531);
nor U13368 (N_13368,N_8052,N_1143);
and U13369 (N_13369,N_6310,N_204);
nor U13370 (N_13370,N_7879,N_6834);
xor U13371 (N_13371,N_3972,N_9093);
and U13372 (N_13372,N_6621,N_5528);
nor U13373 (N_13373,N_4705,N_257);
and U13374 (N_13374,N_131,N_8328);
nand U13375 (N_13375,N_8412,N_8403);
nor U13376 (N_13376,N_6792,N_9736);
nand U13377 (N_13377,N_1005,N_1783);
xor U13378 (N_13378,N_5527,N_7149);
xor U13379 (N_13379,N_2142,N_8382);
nor U13380 (N_13380,N_7417,N_826);
and U13381 (N_13381,N_1742,N_2727);
xnor U13382 (N_13382,N_1475,N_6237);
xnor U13383 (N_13383,N_2191,N_8992);
or U13384 (N_13384,N_4522,N_7739);
xnor U13385 (N_13385,N_9887,N_5463);
or U13386 (N_13386,N_758,N_3722);
and U13387 (N_13387,N_8080,N_3018);
xnor U13388 (N_13388,N_6346,N_8993);
or U13389 (N_13389,N_5169,N_1659);
nand U13390 (N_13390,N_5470,N_343);
xor U13391 (N_13391,N_48,N_1569);
nand U13392 (N_13392,N_1493,N_7816);
nor U13393 (N_13393,N_5269,N_7065);
nor U13394 (N_13394,N_7978,N_6379);
nor U13395 (N_13395,N_2072,N_6844);
or U13396 (N_13396,N_179,N_9492);
xor U13397 (N_13397,N_2977,N_1540);
and U13398 (N_13398,N_4766,N_8419);
or U13399 (N_13399,N_1870,N_8336);
and U13400 (N_13400,N_3226,N_9796);
and U13401 (N_13401,N_4319,N_3808);
and U13402 (N_13402,N_1620,N_1590);
nor U13403 (N_13403,N_1522,N_3614);
xnor U13404 (N_13404,N_143,N_8065);
xor U13405 (N_13405,N_1834,N_9248);
nand U13406 (N_13406,N_3970,N_4835);
nor U13407 (N_13407,N_2506,N_4751);
xnor U13408 (N_13408,N_4390,N_795);
xor U13409 (N_13409,N_2057,N_7168);
and U13410 (N_13410,N_6818,N_6047);
and U13411 (N_13411,N_1409,N_2663);
or U13412 (N_13412,N_5787,N_8999);
xor U13413 (N_13413,N_6589,N_5421);
and U13414 (N_13414,N_9560,N_1344);
nand U13415 (N_13415,N_5203,N_8818);
and U13416 (N_13416,N_6796,N_7091);
nor U13417 (N_13417,N_7867,N_743);
or U13418 (N_13418,N_6950,N_4143);
and U13419 (N_13419,N_7010,N_6380);
nand U13420 (N_13420,N_2170,N_8195);
and U13421 (N_13421,N_7529,N_8037);
or U13422 (N_13422,N_1863,N_1193);
or U13423 (N_13423,N_9563,N_9555);
xor U13424 (N_13424,N_9008,N_5565);
xor U13425 (N_13425,N_3488,N_8594);
xnor U13426 (N_13426,N_9025,N_7741);
nor U13427 (N_13427,N_2886,N_4040);
nand U13428 (N_13428,N_1448,N_6921);
nor U13429 (N_13429,N_2936,N_1589);
nand U13430 (N_13430,N_6128,N_9768);
xor U13431 (N_13431,N_6651,N_4501);
and U13432 (N_13432,N_6306,N_7312);
and U13433 (N_13433,N_1094,N_4917);
or U13434 (N_13434,N_4574,N_4155);
nand U13435 (N_13435,N_8205,N_3392);
xnor U13436 (N_13436,N_6057,N_6286);
or U13437 (N_13437,N_5285,N_9103);
nor U13438 (N_13438,N_9633,N_3907);
or U13439 (N_13439,N_6527,N_57);
and U13440 (N_13440,N_862,N_8395);
and U13441 (N_13441,N_4661,N_8975);
xnor U13442 (N_13442,N_5051,N_3221);
nor U13443 (N_13443,N_7098,N_9235);
xnor U13444 (N_13444,N_389,N_2832);
nand U13445 (N_13445,N_102,N_1330);
nor U13446 (N_13446,N_7946,N_2444);
nor U13447 (N_13447,N_9046,N_3258);
xor U13448 (N_13448,N_7097,N_9884);
and U13449 (N_13449,N_1054,N_4818);
xnor U13450 (N_13450,N_990,N_8107);
nor U13451 (N_13451,N_6548,N_4738);
xnor U13452 (N_13452,N_3351,N_3999);
xor U13453 (N_13453,N_9184,N_6457);
or U13454 (N_13454,N_944,N_22);
nor U13455 (N_13455,N_2860,N_4538);
xnor U13456 (N_13456,N_6500,N_6878);
or U13457 (N_13457,N_4914,N_8674);
nor U13458 (N_13458,N_1423,N_7211);
nor U13459 (N_13459,N_1943,N_2214);
and U13460 (N_13460,N_7647,N_9415);
nor U13461 (N_13461,N_7789,N_5154);
or U13462 (N_13462,N_5870,N_5540);
xor U13463 (N_13463,N_6343,N_3565);
xnor U13464 (N_13464,N_245,N_7158);
and U13465 (N_13465,N_980,N_5418);
xor U13466 (N_13466,N_8964,N_2905);
nor U13467 (N_13467,N_11,N_7239);
nor U13468 (N_13468,N_1512,N_7939);
nor U13469 (N_13469,N_7921,N_9266);
xnor U13470 (N_13470,N_8354,N_9842);
xor U13471 (N_13471,N_9977,N_3418);
nand U13472 (N_13472,N_1538,N_8926);
nand U13473 (N_13473,N_3872,N_1560);
xor U13474 (N_13474,N_3490,N_8010);
nand U13475 (N_13475,N_4181,N_5078);
and U13476 (N_13476,N_3126,N_1195);
or U13477 (N_13477,N_1563,N_7836);
and U13478 (N_13478,N_8771,N_2693);
and U13479 (N_13479,N_2769,N_3604);
and U13480 (N_13480,N_2386,N_1877);
nor U13481 (N_13481,N_9808,N_5682);
and U13482 (N_13482,N_2505,N_3304);
xor U13483 (N_13483,N_1410,N_9572);
xor U13484 (N_13484,N_2911,N_3026);
nand U13485 (N_13485,N_9539,N_6993);
xor U13486 (N_13486,N_4580,N_5881);
nor U13487 (N_13487,N_117,N_8398);
xnor U13488 (N_13488,N_9124,N_754);
or U13489 (N_13489,N_6852,N_2230);
nor U13490 (N_13490,N_690,N_1649);
and U13491 (N_13491,N_1366,N_5674);
xor U13492 (N_13492,N_3388,N_2997);
or U13493 (N_13493,N_81,N_772);
or U13494 (N_13494,N_9744,N_1466);
or U13495 (N_13495,N_2718,N_3284);
nor U13496 (N_13496,N_3691,N_1027);
nor U13497 (N_13497,N_8633,N_5491);
xor U13498 (N_13498,N_1796,N_3708);
and U13499 (N_13499,N_3021,N_7583);
nand U13500 (N_13500,N_5348,N_7148);
or U13501 (N_13501,N_1748,N_1991);
xor U13502 (N_13502,N_9289,N_2521);
nand U13503 (N_13503,N_6363,N_9855);
and U13504 (N_13504,N_4087,N_3384);
and U13505 (N_13505,N_6104,N_7257);
nand U13506 (N_13506,N_1811,N_2148);
and U13507 (N_13507,N_4380,N_4130);
or U13508 (N_13508,N_5635,N_6564);
nand U13509 (N_13509,N_9152,N_9297);
xor U13510 (N_13510,N_5186,N_1945);
nand U13511 (N_13511,N_8688,N_7275);
nor U13512 (N_13512,N_5584,N_4313);
nor U13513 (N_13513,N_6335,N_2710);
xor U13514 (N_13514,N_9469,N_7995);
and U13515 (N_13515,N_9256,N_2128);
nor U13516 (N_13516,N_8044,N_8914);
xor U13517 (N_13517,N_9568,N_8908);
nor U13518 (N_13518,N_8742,N_1234);
xnor U13519 (N_13519,N_9599,N_7787);
nand U13520 (N_13520,N_5744,N_5708);
and U13521 (N_13521,N_7437,N_5217);
or U13522 (N_13522,N_7381,N_3623);
xnor U13523 (N_13523,N_2322,N_8680);
or U13524 (N_13524,N_2794,N_1527);
nor U13525 (N_13525,N_8070,N_5544);
xnor U13526 (N_13526,N_6972,N_4944);
nor U13527 (N_13527,N_3880,N_8616);
or U13528 (N_13528,N_4472,N_7156);
nand U13529 (N_13529,N_3378,N_992);
nand U13530 (N_13530,N_6605,N_3028);
or U13531 (N_13531,N_9419,N_8380);
nor U13532 (N_13532,N_6549,N_8198);
and U13533 (N_13533,N_3783,N_4069);
nand U13534 (N_13534,N_3792,N_3257);
and U13535 (N_13535,N_8491,N_3464);
nand U13536 (N_13536,N_4259,N_8645);
and U13537 (N_13537,N_3243,N_840);
nor U13538 (N_13538,N_2130,N_2286);
xnor U13539 (N_13539,N_4399,N_555);
or U13540 (N_13540,N_7055,N_9706);
nand U13541 (N_13541,N_5917,N_844);
and U13542 (N_13542,N_5959,N_5205);
and U13543 (N_13543,N_9900,N_9117);
xor U13544 (N_13544,N_8896,N_6192);
and U13545 (N_13545,N_7776,N_3815);
or U13546 (N_13546,N_2970,N_4537);
and U13547 (N_13547,N_714,N_408);
xnor U13548 (N_13548,N_8451,N_1949);
xor U13549 (N_13549,N_5595,N_5281);
and U13550 (N_13550,N_9843,N_3568);
xnor U13551 (N_13551,N_2880,N_7604);
nand U13552 (N_13552,N_3453,N_7587);
nor U13553 (N_13553,N_6316,N_3790);
nor U13554 (N_13554,N_58,N_1268);
or U13555 (N_13555,N_542,N_2717);
nand U13556 (N_13556,N_3664,N_2169);
xnor U13557 (N_13557,N_981,N_8397);
and U13558 (N_13558,N_5746,N_4554);
or U13559 (N_13559,N_3577,N_8043);
or U13560 (N_13560,N_5299,N_2617);
or U13561 (N_13561,N_2428,N_6749);
nand U13562 (N_13562,N_331,N_4986);
xor U13563 (N_13563,N_5020,N_16);
and U13564 (N_13564,N_6777,N_6849);
and U13565 (N_13565,N_8702,N_6478);
nor U13566 (N_13566,N_5077,N_5117);
and U13567 (N_13567,N_2658,N_5315);
or U13568 (N_13568,N_7886,N_8307);
or U13569 (N_13569,N_7248,N_2259);
nand U13570 (N_13570,N_4964,N_986);
nand U13571 (N_13571,N_7990,N_3025);
nand U13572 (N_13572,N_649,N_9846);
or U13573 (N_13573,N_3206,N_9094);
nand U13574 (N_13574,N_2734,N_2355);
and U13575 (N_13575,N_4400,N_7198);
nor U13576 (N_13576,N_1353,N_6406);
or U13577 (N_13577,N_4166,N_7430);
or U13578 (N_13578,N_3627,N_3827);
and U13579 (N_13579,N_4727,N_6120);
and U13580 (N_13580,N_4931,N_7234);
xnor U13581 (N_13581,N_6326,N_2243);
nand U13582 (N_13582,N_4899,N_7045);
or U13583 (N_13583,N_1049,N_6373);
or U13584 (N_13584,N_2320,N_7912);
nor U13585 (N_13585,N_5201,N_8369);
nand U13586 (N_13586,N_8691,N_7646);
or U13587 (N_13587,N_9580,N_4826);
xor U13588 (N_13588,N_3234,N_4067);
nand U13589 (N_13589,N_494,N_5485);
or U13590 (N_13590,N_4162,N_804);
or U13591 (N_13591,N_559,N_6663);
and U13592 (N_13592,N_1203,N_5449);
and U13593 (N_13593,N_6197,N_3932);
and U13594 (N_13594,N_5534,N_6245);
and U13595 (N_13595,N_5295,N_556);
xor U13596 (N_13596,N_765,N_9591);
nand U13597 (N_13597,N_2943,N_7357);
nor U13598 (N_13598,N_8155,N_6474);
xnor U13599 (N_13599,N_4778,N_8465);
and U13600 (N_13600,N_2368,N_6352);
or U13601 (N_13601,N_5109,N_7135);
nand U13602 (N_13602,N_1888,N_9901);
xor U13603 (N_13603,N_3947,N_7474);
nand U13604 (N_13604,N_1327,N_1382);
and U13605 (N_13605,N_258,N_9899);
nand U13606 (N_13606,N_6916,N_1503);
nand U13607 (N_13607,N_1188,N_480);
nand U13608 (N_13608,N_2020,N_6808);
nand U13609 (N_13609,N_9765,N_2536);
nand U13610 (N_13610,N_260,N_5862);
nor U13611 (N_13611,N_9941,N_8566);
and U13612 (N_13612,N_1840,N_156);
or U13613 (N_13613,N_8295,N_9743);
nor U13614 (N_13614,N_3142,N_4083);
xor U13615 (N_13615,N_8740,N_5581);
or U13616 (N_13616,N_6522,N_8830);
xor U13617 (N_13617,N_2833,N_7324);
xor U13618 (N_13618,N_668,N_8300);
xnor U13619 (N_13619,N_4164,N_7160);
nor U13620 (N_13620,N_5969,N_5006);
and U13621 (N_13621,N_6532,N_2645);
nand U13622 (N_13622,N_9969,N_9660);
or U13623 (N_13623,N_4096,N_6289);
xnor U13624 (N_13624,N_8111,N_884);
and U13625 (N_13625,N_5135,N_6574);
xor U13626 (N_13626,N_575,N_5040);
and U13627 (N_13627,N_7139,N_4321);
nor U13628 (N_13628,N_6152,N_3877);
nand U13629 (N_13629,N_1429,N_9426);
or U13630 (N_13630,N_7229,N_3292);
and U13631 (N_13631,N_341,N_1922);
nand U13632 (N_13632,N_80,N_644);
or U13633 (N_13633,N_2956,N_7271);
and U13634 (N_13634,N_2641,N_3352);
nor U13635 (N_13635,N_7411,N_7521);
nand U13636 (N_13636,N_2785,N_1730);
nand U13637 (N_13637,N_357,N_9222);
or U13638 (N_13638,N_940,N_1159);
nor U13639 (N_13639,N_5429,N_9001);
nand U13640 (N_13640,N_3644,N_4225);
nor U13641 (N_13641,N_1225,N_5853);
or U13642 (N_13642,N_8192,N_9685);
xnor U13643 (N_13643,N_8837,N_6261);
nor U13644 (N_13644,N_5369,N_5760);
xor U13645 (N_13645,N_2012,N_8933);
or U13646 (N_13646,N_3747,N_2031);
or U13647 (N_13647,N_4238,N_1294);
nor U13648 (N_13648,N_6664,N_8883);
xnor U13649 (N_13649,N_276,N_4743);
and U13650 (N_13650,N_5174,N_4304);
or U13651 (N_13651,N_6599,N_3530);
nand U13652 (N_13652,N_7675,N_9209);
and U13653 (N_13653,N_36,N_1567);
or U13654 (N_13654,N_1217,N_2774);
nand U13655 (N_13655,N_6923,N_269);
nand U13656 (N_13656,N_4202,N_441);
nand U13657 (N_13657,N_4276,N_3603);
nand U13658 (N_13658,N_3427,N_5400);
nand U13659 (N_13659,N_3817,N_3456);
nor U13660 (N_13660,N_4933,N_7462);
nor U13661 (N_13661,N_9985,N_2017);
or U13662 (N_13662,N_4706,N_4573);
xor U13663 (N_13663,N_9411,N_2061);
and U13664 (N_13664,N_316,N_9752);
xnor U13665 (N_13665,N_6083,N_8358);
nor U13666 (N_13666,N_8646,N_5027);
nor U13667 (N_13667,N_1199,N_6633);
xor U13668 (N_13668,N_2415,N_6258);
and U13669 (N_13669,N_2033,N_8895);
and U13670 (N_13670,N_8605,N_1665);
or U13671 (N_13671,N_9799,N_5773);
xnor U13672 (N_13672,N_9613,N_1757);
nor U13673 (N_13673,N_7074,N_2914);
and U13674 (N_13674,N_4864,N_9339);
and U13675 (N_13675,N_353,N_9135);
and U13676 (N_13676,N_9131,N_1562);
nand U13677 (N_13677,N_4622,N_3326);
or U13678 (N_13678,N_1472,N_8756);
and U13679 (N_13679,N_1276,N_8158);
xor U13680 (N_13680,N_7033,N_7093);
nand U13681 (N_13681,N_8591,N_4543);
xnor U13682 (N_13682,N_5080,N_6939);
nand U13683 (N_13683,N_219,N_3861);
or U13684 (N_13684,N_2712,N_8817);
nor U13685 (N_13685,N_3218,N_4652);
xnor U13686 (N_13686,N_1534,N_4576);
and U13687 (N_13687,N_8965,N_5742);
or U13688 (N_13688,N_4925,N_5318);
and U13689 (N_13689,N_5079,N_5402);
and U13690 (N_13690,N_1786,N_846);
and U13691 (N_13691,N_6714,N_6073);
or U13692 (N_13692,N_1619,N_1767);
xor U13693 (N_13693,N_4022,N_5658);
and U13694 (N_13694,N_1152,N_2333);
and U13695 (N_13695,N_8130,N_1998);
nand U13696 (N_13696,N_9810,N_2239);
or U13697 (N_13697,N_657,N_2337);
xnor U13698 (N_13698,N_461,N_7618);
nand U13699 (N_13699,N_2927,N_3242);
nand U13700 (N_13700,N_7427,N_921);
xnor U13701 (N_13701,N_3601,N_5219);
nand U13702 (N_13702,N_7720,N_551);
or U13703 (N_13703,N_3912,N_5273);
or U13704 (N_13704,N_4745,N_1270);
nor U13705 (N_13705,N_209,N_9883);
nor U13706 (N_13706,N_928,N_1709);
or U13707 (N_13707,N_1099,N_5592);
or U13708 (N_13708,N_3669,N_1384);
or U13709 (N_13709,N_133,N_2780);
and U13710 (N_13710,N_4731,N_856);
or U13711 (N_13711,N_9173,N_8426);
nor U13712 (N_13712,N_7073,N_8921);
nand U13713 (N_13713,N_5766,N_1525);
and U13714 (N_13714,N_2000,N_4277);
or U13715 (N_13715,N_554,N_5519);
nand U13716 (N_13716,N_9818,N_6781);
nand U13717 (N_13717,N_8723,N_825);
or U13718 (N_13718,N_451,N_3358);
and U13719 (N_13719,N_1759,N_3374);
nor U13720 (N_13720,N_2272,N_5897);
nand U13721 (N_13721,N_7889,N_5873);
nand U13722 (N_13722,N_6510,N_518);
xnor U13723 (N_13723,N_8516,N_7562);
nand U13724 (N_13724,N_6332,N_6882);
and U13725 (N_13725,N_3330,N_5050);
xnor U13726 (N_13726,N_6896,N_6378);
nand U13727 (N_13727,N_302,N_3180);
nand U13728 (N_13728,N_4079,N_7291);
xor U13729 (N_13729,N_5422,N_1439);
nand U13730 (N_13730,N_1599,N_2458);
and U13731 (N_13731,N_2871,N_8269);
nand U13732 (N_13732,N_1403,N_4101);
xor U13733 (N_13733,N_9872,N_6070);
nor U13734 (N_13734,N_7188,N_858);
nor U13735 (N_13735,N_5932,N_6936);
xnor U13736 (N_13736,N_9264,N_3749);
xnor U13737 (N_13737,N_4759,N_8727);
and U13738 (N_13738,N_6566,N_5921);
and U13739 (N_13739,N_2669,N_622);
or U13740 (N_13740,N_4053,N_5291);
nor U13741 (N_13741,N_297,N_2878);
nor U13742 (N_13742,N_5215,N_4496);
xnor U13743 (N_13743,N_255,N_4289);
xor U13744 (N_13744,N_6220,N_4349);
or U13745 (N_13745,N_918,N_4892);
or U13746 (N_13746,N_4636,N_5165);
nand U13747 (N_13747,N_1488,N_7894);
xor U13748 (N_13748,N_512,N_111);
nand U13749 (N_13749,N_4290,N_857);
and U13750 (N_13750,N_1277,N_2953);
nand U13751 (N_13751,N_4233,N_5758);
and U13752 (N_13752,N_3742,N_395);
and U13753 (N_13753,N_2425,N_4476);
or U13754 (N_13754,N_4891,N_7448);
xor U13755 (N_13755,N_9576,N_9761);
nand U13756 (N_13756,N_8298,N_4908);
or U13757 (N_13757,N_1184,N_3686);
xnor U13758 (N_13758,N_4627,N_7592);
and U13759 (N_13759,N_5034,N_7799);
nor U13760 (N_13760,N_938,N_1284);
xor U13761 (N_13761,N_7128,N_516);
xor U13762 (N_13762,N_4991,N_8651);
and U13763 (N_13763,N_5707,N_3278);
xor U13764 (N_13764,N_7133,N_5678);
nor U13765 (N_13765,N_3760,N_8140);
xor U13766 (N_13766,N_2349,N_2306);
xnor U13767 (N_13767,N_6097,N_4047);
xor U13768 (N_13768,N_537,N_2083);
and U13769 (N_13769,N_8898,N_7320);
and U13770 (N_13770,N_3917,N_9596);
nand U13771 (N_13771,N_6481,N_33);
nand U13772 (N_13772,N_2279,N_577);
nor U13773 (N_13773,N_9000,N_3035);
and U13774 (N_13774,N_7965,N_9106);
xor U13775 (N_13775,N_1325,N_8104);
nor U13776 (N_13776,N_5046,N_1379);
nor U13777 (N_13777,N_8831,N_2918);
nand U13778 (N_13778,N_5145,N_5060);
or U13779 (N_13779,N_3633,N_8523);
xor U13780 (N_13780,N_2071,N_965);
or U13781 (N_13781,N_6276,N_5513);
and U13782 (N_13782,N_8652,N_2374);
nor U13783 (N_13783,N_2199,N_6540);
nor U13784 (N_13784,N_805,N_5759);
nand U13785 (N_13785,N_6998,N_7169);
nand U13786 (N_13786,N_2413,N_6188);
or U13787 (N_13787,N_4987,N_1272);
xor U13788 (N_13788,N_6567,N_5414);
xnor U13789 (N_13789,N_5244,N_3498);
xnor U13790 (N_13790,N_9800,N_7940);
or U13791 (N_13791,N_9882,N_8174);
nand U13792 (N_13792,N_5762,N_1059);
xnor U13793 (N_13793,N_187,N_5290);
and U13794 (N_13794,N_2998,N_2768);
nand U13795 (N_13795,N_8604,N_5407);
or U13796 (N_13796,N_7821,N_4972);
nor U13797 (N_13797,N_2993,N_2809);
xor U13798 (N_13798,N_7870,N_1939);
nand U13799 (N_13799,N_4621,N_7077);
xnor U13800 (N_13800,N_9279,N_8596);
nand U13801 (N_13801,N_6036,N_7483);
and U13802 (N_13802,N_6342,N_8236);
or U13803 (N_13803,N_5341,N_5698);
xor U13804 (N_13804,N_2844,N_9362);
or U13805 (N_13805,N_2389,N_2025);
xor U13806 (N_13806,N_6505,N_3209);
or U13807 (N_13807,N_893,N_2716);
and U13808 (N_13808,N_8942,N_867);
xor U13809 (N_13809,N_3178,N_2344);
or U13810 (N_13810,N_9453,N_4009);
nand U13811 (N_13811,N_3564,N_8928);
nand U13812 (N_13812,N_9078,N_506);
xor U13813 (N_13813,N_2836,N_5660);
nand U13814 (N_13814,N_6176,N_3232);
nor U13815 (N_13815,N_1140,N_7864);
or U13816 (N_13816,N_1179,N_7068);
nor U13817 (N_13817,N_3929,N_9352);
nand U13818 (N_13818,N_3145,N_548);
and U13819 (N_13819,N_7365,N_2228);
nor U13820 (N_13820,N_3580,N_7202);
nor U13821 (N_13821,N_8138,N_8943);
or U13822 (N_13822,N_7246,N_7064);
or U13823 (N_13823,N_8040,N_1245);
nor U13824 (N_13824,N_3079,N_4658);
xor U13825 (N_13825,N_2806,N_4368);
xnor U13826 (N_13826,N_1999,N_8541);
nand U13827 (N_13827,N_4373,N_2463);
and U13828 (N_13828,N_7327,N_3151);
nand U13829 (N_13829,N_9830,N_7351);
xnor U13830 (N_13830,N_1506,N_3353);
and U13831 (N_13831,N_9987,N_2045);
or U13832 (N_13832,N_4643,N_2765);
and U13833 (N_13833,N_5745,N_4475);
xor U13834 (N_13834,N_120,N_1436);
or U13835 (N_13835,N_7247,N_8200);
or U13836 (N_13836,N_4065,N_1537);
and U13837 (N_13837,N_2408,N_9179);
xor U13838 (N_13838,N_9406,N_6690);
xnor U13839 (N_13839,N_8013,N_137);
nand U13840 (N_13840,N_1727,N_9287);
and U13841 (N_13841,N_1653,N_7850);
xnor U13842 (N_13842,N_3007,N_8735);
and U13843 (N_13843,N_5440,N_7252);
xor U13844 (N_13844,N_3704,N_1966);
nor U13845 (N_13845,N_5082,N_501);
nor U13846 (N_13846,N_418,N_2343);
xor U13847 (N_13847,N_3375,N_9858);
or U13848 (N_13848,N_3922,N_854);
nor U13849 (N_13849,N_4473,N_8193);
nand U13850 (N_13850,N_5650,N_711);
and U13851 (N_13851,N_9957,N_8350);
nor U13852 (N_13852,N_8278,N_1373);
or U13853 (N_13853,N_4120,N_9423);
nor U13854 (N_13854,N_528,N_9763);
and U13855 (N_13855,N_759,N_3268);
or U13856 (N_13856,N_8576,N_5920);
xnor U13857 (N_13857,N_1617,N_435);
xnor U13858 (N_13858,N_262,N_1023);
or U13859 (N_13859,N_2633,N_6105);
nor U13860 (N_13860,N_2496,N_2338);
and U13861 (N_13861,N_4347,N_8910);
and U13862 (N_13862,N_5721,N_9942);
or U13863 (N_13863,N_1200,N_324);
nor U13864 (N_13864,N_812,N_8861);
nor U13865 (N_13865,N_8256,N_6013);
or U13866 (N_13866,N_3108,N_7392);
and U13867 (N_13867,N_2018,N_5715);
nor U13868 (N_13868,N_1470,N_1011);
xnor U13869 (N_13869,N_5756,N_8534);
nor U13870 (N_13870,N_7941,N_1288);
xnor U13871 (N_13871,N_8555,N_9295);
and U13872 (N_13872,N_116,N_7379);
or U13873 (N_13873,N_1989,N_1221);
nor U13874 (N_13874,N_4929,N_9979);
xor U13875 (N_13875,N_821,N_1501);
or U13876 (N_13876,N_3253,N_7025);
and U13877 (N_13877,N_5502,N_999);
nor U13878 (N_13878,N_3055,N_1902);
and U13879 (N_13879,N_6649,N_641);
nand U13880 (N_13880,N_520,N_8665);
nor U13881 (N_13881,N_5346,N_1869);
nand U13882 (N_13882,N_977,N_6393);
xnor U13883 (N_13883,N_6945,N_6504);
nor U13884 (N_13884,N_1753,N_6804);
or U13885 (N_13885,N_8610,N_536);
nor U13886 (N_13886,N_5984,N_5940);
xnor U13887 (N_13887,N_5270,N_957);
nand U13888 (N_13888,N_6557,N_9230);
nand U13889 (N_13889,N_4342,N_4052);
nor U13890 (N_13890,N_663,N_2873);
nand U13891 (N_13891,N_2007,N_3510);
nor U13892 (N_13892,N_2518,N_8393);
or U13893 (N_13893,N_8745,N_3377);
nand U13894 (N_13894,N_5899,N_450);
xor U13895 (N_13895,N_1778,N_6949);
or U13896 (N_13896,N_2685,N_1071);
or U13897 (N_13897,N_697,N_8413);
xnor U13898 (N_13898,N_3643,N_2484);
xor U13899 (N_13899,N_72,N_168);
or U13900 (N_13900,N_6513,N_1600);
and U13901 (N_13901,N_3215,N_4152);
or U13902 (N_13902,N_5894,N_4439);
and U13903 (N_13903,N_3144,N_2036);
or U13904 (N_13904,N_7901,N_3926);
nand U13905 (N_13905,N_5750,N_3650);
or U13906 (N_13906,N_1408,N_4358);
and U13907 (N_13907,N_4138,N_7788);
nand U13908 (N_13908,N_8437,N_600);
nor U13909 (N_13909,N_2418,N_4895);
or U13910 (N_13910,N_4788,N_3136);
xnor U13911 (N_13911,N_4586,N_303);
or U13912 (N_13912,N_8998,N_8000);
nand U13913 (N_13913,N_3137,N_9052);
and U13914 (N_13914,N_7727,N_178);
nand U13915 (N_13915,N_955,N_8885);
or U13916 (N_13916,N_1220,N_5381);
nand U13917 (N_13917,N_4814,N_2495);
nor U13918 (N_13918,N_311,N_6717);
nand U13919 (N_13919,N_8053,N_5448);
nand U13920 (N_13920,N_7200,N_8018);
nand U13921 (N_13921,N_660,N_3854);
nand U13922 (N_13922,N_9067,N_7542);
nor U13923 (N_13923,N_6079,N_7882);
nor U13924 (N_13924,N_3998,N_3846);
xor U13925 (N_13925,N_9098,N_8819);
nand U13926 (N_13926,N_5185,N_8314);
or U13927 (N_13927,N_8954,N_1719);
xnor U13928 (N_13928,N_5671,N_2764);
xor U13929 (N_13929,N_5444,N_8557);
nor U13930 (N_13930,N_1921,N_2440);
nand U13931 (N_13931,N_9182,N_4722);
and U13932 (N_13932,N_393,N_7704);
or U13933 (N_13933,N_3847,N_9090);
or U13934 (N_13934,N_4234,N_2875);
nand U13935 (N_13935,N_6064,N_3423);
nand U13936 (N_13936,N_5905,N_7942);
nand U13937 (N_13937,N_8945,N_685);
nor U13938 (N_13938,N_37,N_3122);
nor U13939 (N_13939,N_165,N_4126);
and U13940 (N_13940,N_1876,N_2157);
nor U13941 (N_13941,N_9745,N_5936);
or U13942 (N_13942,N_358,N_8116);
nand U13943 (N_13943,N_5243,N_8890);
or U13944 (N_13944,N_7092,N_874);
or U13945 (N_13945,N_31,N_5736);
or U13946 (N_13946,N_7725,N_2123);
nor U13947 (N_13947,N_1252,N_6093);
nand U13948 (N_13948,N_4398,N_9988);
or U13949 (N_13949,N_6447,N_5840);
xnor U13950 (N_13950,N_9802,N_9521);
nand U13951 (N_13951,N_6815,N_9699);
and U13952 (N_13952,N_7702,N_4264);
or U13953 (N_13953,N_956,N_1630);
and U13954 (N_13954,N_729,N_1875);
xor U13955 (N_13955,N_8497,N_4536);
xnor U13956 (N_13956,N_5849,N_3141);
nand U13957 (N_13957,N_7137,N_8570);
xnor U13958 (N_13958,N_954,N_1477);
nor U13959 (N_13959,N_1837,N_1015);
xor U13960 (N_13960,N_3260,N_9456);
xor U13961 (N_13961,N_3011,N_1523);
nor U13962 (N_13962,N_6419,N_1360);
xor U13963 (N_13963,N_2615,N_3566);
xnor U13964 (N_13964,N_1224,N_1553);
xor U13965 (N_13965,N_564,N_7132);
or U13966 (N_13966,N_3417,N_1929);
and U13967 (N_13967,N_693,N_8639);
nor U13968 (N_13968,N_7596,N_511);
nand U13969 (N_13969,N_4517,N_6523);
or U13970 (N_13970,N_1828,N_4878);
xor U13971 (N_13971,N_8853,N_6272);
or U13972 (N_13972,N_9788,N_5661);
and U13973 (N_13973,N_4937,N_6066);
nor U13974 (N_13974,N_4599,N_2604);
or U13975 (N_13975,N_8703,N_9333);
and U13976 (N_13976,N_939,N_3443);
nor U13977 (N_13977,N_9918,N_6961);
and U13978 (N_13978,N_4663,N_1814);
and U13979 (N_13979,N_9416,N_1568);
nor U13980 (N_13980,N_3903,N_5648);
or U13981 (N_13981,N_3462,N_8135);
nor U13982 (N_13982,N_4287,N_4216);
or U13983 (N_13983,N_6713,N_9654);
xnor U13984 (N_13984,N_6012,N_7569);
xor U13985 (N_13985,N_5081,N_2109);
xor U13986 (N_13986,N_7936,N_1576);
nand U13987 (N_13987,N_4821,N_6287);
or U13988 (N_13988,N_4270,N_8629);
xor U13989 (N_13989,N_9964,N_6195);
nand U13990 (N_13990,N_7970,N_9109);
or U13991 (N_13991,N_9741,N_8731);
nand U13992 (N_13992,N_1836,N_9019);
nor U13993 (N_13993,N_3897,N_4750);
nor U13994 (N_13994,N_8850,N_129);
nand U13995 (N_13995,N_1643,N_7460);
nand U13996 (N_13996,N_4437,N_612);
and U13997 (N_13997,N_8747,N_6544);
nor U13998 (N_13998,N_4178,N_3190);
and U13999 (N_13999,N_5339,N_898);
or U14000 (N_14000,N_7827,N_3466);
nand U14001 (N_14001,N_2876,N_3223);
nor U14002 (N_14002,N_2527,N_8545);
or U14003 (N_14003,N_8760,N_9789);
xnor U14004 (N_14004,N_6040,N_4175);
xnor U14005 (N_14005,N_7049,N_2567);
xor U14006 (N_14006,N_7885,N_7328);
nand U14007 (N_14007,N_3780,N_3977);
nand U14008 (N_14008,N_32,N_4396);
xor U14009 (N_14009,N_5075,N_2812);
nor U14010 (N_14010,N_8102,N_5114);
or U14011 (N_14011,N_6723,N_4109);
or U14012 (N_14012,N_9259,N_3871);
or U14013 (N_14013,N_3029,N_4687);
xor U14014 (N_14014,N_5387,N_8045);
nor U14015 (N_14015,N_150,N_8561);
or U14016 (N_14016,N_6637,N_869);
nand U14017 (N_14017,N_6577,N_5956);
and U14018 (N_14018,N_2654,N_2713);
nor U14019 (N_14019,N_8907,N_3574);
and U14020 (N_14020,N_4102,N_2431);
or U14021 (N_14021,N_322,N_1134);
or U14022 (N_14022,N_9366,N_8184);
nor U14023 (N_14023,N_2690,N_2059);
and U14024 (N_14024,N_3773,N_8071);
or U14025 (N_14025,N_6684,N_138);
nand U14026 (N_14026,N_4206,N_4561);
and U14027 (N_14027,N_3767,N_9548);
nor U14028 (N_14028,N_4668,N_6986);
or U14029 (N_14029,N_4463,N_1629);
nand U14030 (N_14030,N_9458,N_5829);
or U14031 (N_14031,N_5210,N_1734);
or U14032 (N_14032,N_6234,N_375);
and U14033 (N_14033,N_3421,N_4923);
xnor U14034 (N_14034,N_6291,N_6836);
or U14035 (N_14035,N_1931,N_9641);
nand U14036 (N_14036,N_8399,N_539);
and U14037 (N_14037,N_6115,N_2454);
nor U14038 (N_14038,N_2303,N_1312);
nor U14039 (N_14039,N_647,N_9814);
or U14040 (N_14040,N_6893,N_7228);
nand U14041 (N_14041,N_1890,N_5642);
nor U14042 (N_14042,N_3176,N_8233);
or U14043 (N_14043,N_1677,N_396);
and U14044 (N_14044,N_3314,N_3584);
xor U14045 (N_14045,N_8036,N_4977);
nor U14046 (N_14046,N_5868,N_7916);
nand U14047 (N_14047,N_1546,N_7640);
nand U14048 (N_14048,N_1770,N_5752);
xnor U14049 (N_14049,N_1502,N_9581);
and U14050 (N_14050,N_362,N_6857);
or U14051 (N_14051,N_1839,N_1558);
nand U14052 (N_14052,N_9999,N_6421);
xnor U14053 (N_14053,N_9621,N_5833);
nor U14054 (N_14054,N_487,N_9602);
nand U14055 (N_14055,N_493,N_107);
nor U14056 (N_14056,N_3509,N_3296);
nand U14057 (N_14057,N_6277,N_3173);
xor U14058 (N_14058,N_3381,N_1773);
nor U14059 (N_14059,N_8033,N_1816);
or U14060 (N_14060,N_7967,N_9639);
or U14061 (N_14061,N_4798,N_9857);
nand U14062 (N_14062,N_1743,N_2634);
or U14063 (N_14063,N_5763,N_9070);
or U14064 (N_14064,N_4255,N_1692);
or U14065 (N_14065,N_2550,N_1017);
nand U14066 (N_14066,N_9584,N_3866);
xor U14067 (N_14067,N_3952,N_9043);
nand U14068 (N_14068,N_2049,N_4436);
and U14069 (N_14069,N_4794,N_6515);
and U14070 (N_14070,N_7259,N_1632);
and U14071 (N_14071,N_3345,N_8210);
and U14072 (N_14072,N_8134,N_7103);
nor U14073 (N_14073,N_3082,N_9374);
nand U14074 (N_14074,N_4028,N_6709);
nor U14075 (N_14075,N_1781,N_1);
nand U14076 (N_14076,N_455,N_2602);
and U14077 (N_14077,N_9646,N_9835);
xor U14078 (N_14078,N_6608,N_7731);
nor U14079 (N_14079,N_5941,N_4911);
nand U14080 (N_14080,N_1187,N_3638);
nor U14081 (N_14081,N_70,N_2835);
xnor U14082 (N_14082,N_1132,N_1595);
or U14083 (N_14083,N_4780,N_2583);
xnor U14084 (N_14084,N_7698,N_4339);
xnor U14085 (N_14085,N_4182,N_9351);
nor U14086 (N_14086,N_8187,N_6218);
and U14087 (N_14087,N_6789,N_9450);
and U14088 (N_14088,N_534,N_1335);
and U14089 (N_14089,N_912,N_321);
nand U14090 (N_14090,N_4201,N_7991);
xnor U14091 (N_14091,N_8131,N_192);
and U14092 (N_14092,N_5326,N_96);
nor U14093 (N_14093,N_7422,N_1051);
and U14094 (N_14094,N_904,N_7733);
nand U14095 (N_14095,N_8532,N_5965);
and U14096 (N_14096,N_1642,N_7340);
or U14097 (N_14097,N_4983,N_3593);
xnor U14098 (N_14098,N_6797,N_798);
nor U14099 (N_14099,N_3899,N_7609);
or U14100 (N_14100,N_8242,N_7356);
xor U14101 (N_14101,N_9590,N_7972);
and U14102 (N_14102,N_7819,N_4737);
nand U14103 (N_14103,N_3830,N_7109);
xnor U14104 (N_14104,N_2901,N_6920);
xor U14105 (N_14105,N_6398,N_6227);
nor U14106 (N_14106,N_9315,N_8664);
nand U14107 (N_14107,N_1213,N_1755);
nand U14108 (N_14108,N_7081,N_1229);
nor U14109 (N_14109,N_5574,N_594);
nand U14110 (N_14110,N_352,N_9659);
nor U14111 (N_14111,N_1306,N_6284);
nand U14112 (N_14112,N_5801,N_5435);
or U14113 (N_14113,N_3171,N_3483);
and U14114 (N_14114,N_1031,N_3411);
nor U14115 (N_14115,N_7274,N_3130);
xnor U14116 (N_14116,N_1255,N_9955);
nand U14117 (N_14117,N_3301,N_6770);
xor U14118 (N_14118,N_5226,N_5696);
nand U14119 (N_14119,N_4694,N_9541);
xnor U14120 (N_14120,N_3097,N_1548);
nor U14121 (N_14121,N_3368,N_8573);
nor U14122 (N_14122,N_7099,N_7030);
xor U14123 (N_14123,N_744,N_2975);
xor U14124 (N_14124,N_7770,N_3272);
xnor U14125 (N_14125,N_1833,N_3312);
and U14126 (N_14126,N_9593,N_2297);
nor U14127 (N_14127,N_6886,N_2524);
xor U14128 (N_14128,N_8183,N_1942);
xnor U14129 (N_14129,N_3440,N_6718);
or U14130 (N_14130,N_2212,N_1371);
and U14131 (N_14131,N_3549,N_1174);
and U14132 (N_14132,N_6559,N_7630);
or U14133 (N_14133,N_4117,N_6912);
nor U14134 (N_14134,N_5739,N_6160);
nand U14135 (N_14135,N_8335,N_8828);
or U14136 (N_14136,N_9777,N_2252);
xor U14137 (N_14137,N_4486,N_5777);
and U14138 (N_14138,N_3884,N_2174);
nor U14139 (N_14139,N_333,N_6149);
nor U14140 (N_14140,N_2564,N_8863);
xor U14141 (N_14141,N_6241,N_3076);
and U14142 (N_14142,N_3102,N_7966);
or U14143 (N_14143,N_5511,N_4381);
or U14144 (N_14144,N_8913,N_2922);
nor U14145 (N_14145,N_8619,N_9854);
xnor U14146 (N_14146,N_6978,N_1126);
or U14147 (N_14147,N_2116,N_6207);
and U14148 (N_14148,N_3134,N_471);
xnor U14149 (N_14149,N_5159,N_1698);
nor U14150 (N_14150,N_5257,N_8228);
nand U14151 (N_14151,N_1281,N_1807);
xnor U14152 (N_14152,N_8450,N_1691);
nor U14153 (N_14153,N_2254,N_4873);
and U14154 (N_14154,N_2588,N_848);
nor U14155 (N_14155,N_3677,N_907);
xor U14156 (N_14156,N_5469,N_9104);
nor U14157 (N_14157,N_2215,N_7959);
nor U14158 (N_14158,N_1784,N_6130);
nand U14159 (N_14159,N_1079,N_381);
nor U14160 (N_14160,N_3785,N_2276);
nor U14161 (N_14161,N_9702,N_6729);
nand U14162 (N_14162,N_6588,N_5134);
xor U14163 (N_14163,N_5475,N_7639);
or U14164 (N_14164,N_8714,N_5128);
and U14165 (N_14165,N_296,N_3751);
and U14166 (N_14166,N_8575,N_4209);
and U14167 (N_14167,N_5311,N_3088);
nor U14168 (N_14168,N_8481,N_1900);
nand U14169 (N_14169,N_1300,N_8166);
xor U14170 (N_14170,N_6423,N_4246);
xnor U14171 (N_14171,N_2553,N_3224);
nor U14172 (N_14172,N_9234,N_8613);
xnor U14173 (N_14173,N_8179,N_4684);
nand U14174 (N_14174,N_2241,N_1498);
nor U14175 (N_14175,N_2702,N_1232);
nor U14176 (N_14176,N_9569,N_8950);
nand U14177 (N_14177,N_9481,N_3771);
nor U14178 (N_14178,N_4569,N_4916);
or U14179 (N_14179,N_3065,N_6861);
nor U14180 (N_14180,N_2194,N_7243);
and U14181 (N_14181,N_1995,N_6465);
nor U14182 (N_14182,N_193,N_8280);
or U14183 (N_14183,N_5144,N_9767);
and U14184 (N_14184,N_5996,N_9062);
nor U14185 (N_14185,N_1825,N_7599);
xor U14186 (N_14186,N_113,N_7782);
and U14187 (N_14187,N_7515,N_3617);
and U14188 (N_14188,N_5303,N_7185);
nand U14189 (N_14189,N_1526,N_7378);
xor U14190 (N_14190,N_1997,N_951);
nor U14191 (N_14191,N_4366,N_3832);
xor U14192 (N_14192,N_7881,N_2638);
or U14193 (N_14193,N_8813,N_9369);
or U14194 (N_14194,N_847,N_5545);
nor U14195 (N_14195,N_6668,N_4300);
or U14196 (N_14196,N_7871,N_3020);
xnor U14197 (N_14197,N_8601,N_8152);
xor U14198 (N_14198,N_1917,N_7382);
or U14199 (N_14199,N_7620,N_6715);
xor U14200 (N_14200,N_184,N_9869);
or U14201 (N_14201,N_5874,N_2156);
nand U14202 (N_14202,N_6587,N_8957);
xor U14203 (N_14203,N_7672,N_5415);
or U14204 (N_14204,N_4822,N_4924);
and U14205 (N_14205,N_4761,N_6084);
and U14206 (N_14206,N_3796,N_3327);
nor U14207 (N_14207,N_1726,N_1689);
or U14208 (N_14208,N_2747,N_4221);
nor U14209 (N_14209,N_2612,N_5155);
nand U14210 (N_14210,N_7710,N_628);
nor U14211 (N_14211,N_4112,N_1722);
or U14212 (N_14212,N_2154,N_5578);
or U14213 (N_14213,N_5337,N_9972);
xor U14214 (N_14214,N_9839,N_7424);
xnor U14215 (N_14215,N_5460,N_2497);
nand U14216 (N_14216,N_2610,N_8276);
or U14217 (N_14217,N_2798,N_6069);
nor U14218 (N_14218,N_1407,N_3031);
nor U14219 (N_14219,N_325,N_4869);
and U14220 (N_14220,N_1636,N_778);
and U14221 (N_14221,N_7134,N_5903);
xor U14222 (N_14222,N_8620,N_9487);
or U14223 (N_14223,N_4108,N_6909);
nand U14224 (N_14224,N_7084,N_2185);
or U14225 (N_14225,N_4377,N_8877);
nor U14226 (N_14226,N_7588,N_4205);
or U14227 (N_14227,N_3149,N_4879);
nor U14228 (N_14228,N_5619,N_4763);
xor U14229 (N_14229,N_7623,N_3256);
nor U14230 (N_14230,N_2941,N_2208);
or U14231 (N_14231,N_1607,N_7408);
or U14232 (N_14232,N_872,N_6228);
and U14233 (N_14233,N_6487,N_3000);
nand U14234 (N_14234,N_9308,N_8169);
xor U14235 (N_14235,N_2152,N_1856);
and U14236 (N_14236,N_7446,N_3499);
or U14237 (N_14237,N_6955,N_2543);
or U14238 (N_14238,N_6143,N_3500);
or U14239 (N_14239,N_6407,N_5831);
and U14240 (N_14240,N_4581,N_6098);
nand U14241 (N_14241,N_6456,N_1166);
xor U14242 (N_14242,N_1894,N_4981);
nand U14243 (N_14243,N_9373,N_6053);
nor U14244 (N_14244,N_1090,N_5614);
or U14245 (N_14245,N_3590,N_2419);
nor U14246 (N_14246,N_5520,N_8331);
or U14247 (N_14247,N_7394,N_4549);
nor U14248 (N_14248,N_6062,N_2058);
nand U14249 (N_14249,N_6328,N_9099);
nand U14250 (N_14250,N_3447,N_4906);
or U14251 (N_14251,N_7703,N_605);
nor U14252 (N_14252,N_9280,N_298);
nand U14253 (N_14253,N_2079,N_8118);
or U14254 (N_14254,N_4105,N_1782);
nand U14255 (N_14255,N_6535,N_4382);
nand U14256 (N_14256,N_6081,N_100);
or U14257 (N_14257,N_5183,N_2906);
nand U14258 (N_14258,N_1667,N_3924);
and U14259 (N_14259,N_5819,N_9603);
nor U14260 (N_14260,N_2802,N_9821);
and U14261 (N_14261,N_3287,N_6403);
or U14262 (N_14262,N_9870,N_8329);
nand U14263 (N_14263,N_5960,N_5820);
xor U14264 (N_14264,N_2609,N_661);
nor U14265 (N_14265,N_9807,N_2882);
nand U14266 (N_14266,N_6890,N_8401);
and U14267 (N_14267,N_9951,N_8679);
xnor U14268 (N_14268,N_7005,N_5567);
nor U14269 (N_14269,N_3573,N_2519);
xnor U14270 (N_14270,N_2772,N_7352);
or U14271 (N_14271,N_2819,N_7193);
nor U14272 (N_14272,N_1264,N_9848);
nor U14273 (N_14273,N_114,N_2635);
and U14274 (N_14274,N_4558,N_8656);
nor U14275 (N_14275,N_789,N_3291);
nand U14276 (N_14276,N_2811,N_4868);
nand U14277 (N_14277,N_8392,N_4059);
and U14278 (N_14278,N_8682,N_8974);
nor U14279 (N_14279,N_4141,N_4612);
or U14280 (N_14280,N_2535,N_2820);
nand U14281 (N_14281,N_535,N_5847);
or U14282 (N_14282,N_3848,N_8240);
nand U14283 (N_14283,N_7841,N_9829);
nor U14284 (N_14284,N_2347,N_8128);
nor U14285 (N_14285,N_3432,N_5478);
nor U14286 (N_14286,N_419,N_1216);
and U14287 (N_14287,N_6427,N_5947);
and U14288 (N_14288,N_7115,N_8692);
xnor U14289 (N_14289,N_18,N_4757);
nor U14290 (N_14290,N_3849,N_6761);
xor U14291 (N_14291,N_1003,N_4519);
or U14292 (N_14292,N_2391,N_6662);
nand U14293 (N_14293,N_5446,N_8279);
or U14294 (N_14294,N_933,N_2921);
xnor U14295 (N_14295,N_4905,N_6118);
and U14296 (N_14296,N_433,N_4844);
nor U14297 (N_14297,N_5572,N_9804);
nand U14298 (N_14298,N_3523,N_879);
or U14299 (N_14299,N_9178,N_4641);
and U14300 (N_14300,N_3782,N_3597);
nor U14301 (N_14301,N_9630,N_6032);
nor U14302 (N_14302,N_6479,N_5009);
and U14303 (N_14303,N_3951,N_7729);
nor U14304 (N_14304,N_5512,N_1147);
nand U14305 (N_14305,N_7615,N_8739);
nor U14306 (N_14306,N_9229,N_719);
nand U14307 (N_14307,N_8168,N_2342);
or U14308 (N_14308,N_9346,N_9180);
xor U14309 (N_14309,N_8304,N_338);
and U14310 (N_14310,N_2704,N_9983);
xor U14311 (N_14311,N_2678,N_6905);
xnor U14312 (N_14312,N_7496,N_4133);
xor U14313 (N_14313,N_4565,N_7236);
and U14314 (N_14314,N_593,N_4330);
or U14315 (N_14315,N_8666,N_7928);
nand U14316 (N_14316,N_8458,N_656);
nand U14317 (N_14317,N_1747,N_7539);
nor U14318 (N_14318,N_6615,N_1766);
xnor U14319 (N_14319,N_7892,N_8349);
nand U14320 (N_14320,N_2939,N_2238);
or U14321 (N_14321,N_842,N_3494);
or U14322 (N_14322,N_2896,N_674);
nor U14323 (N_14323,N_4340,N_7390);
nor U14324 (N_14324,N_3990,N_1414);
and U14325 (N_14325,N_8715,N_4026);
nand U14326 (N_14326,N_5162,N_1112);
xnor U14327 (N_14327,N_9045,N_1426);
nor U14328 (N_14328,N_8940,N_4523);
xnor U14329 (N_14329,N_4654,N_682);
or U14330 (N_14330,N_8466,N_7914);
nor U14331 (N_14331,N_8920,N_7824);
or U14332 (N_14332,N_6958,N_5206);
nor U14333 (N_14333,N_8707,N_9921);
or U14334 (N_14334,N_69,N_9272);
nand U14335 (N_14335,N_6107,N_7750);
xor U14336 (N_14336,N_5628,N_8519);
nand U14337 (N_14337,N_2954,N_9401);
xor U14338 (N_14338,N_472,N_541);
xor U14339 (N_14339,N_522,N_9825);
nor U14340 (N_14340,N_5427,N_9027);
nand U14341 (N_14341,N_5551,N_9550);
or U14342 (N_14342,N_5409,N_598);
or U14343 (N_14343,N_5255,N_2261);
nand U14344 (N_14344,N_4452,N_7015);
nand U14345 (N_14345,N_427,N_4963);
or U14346 (N_14346,N_7177,N_4669);
or U14347 (N_14347,N_2281,N_1396);
xnor U14348 (N_14348,N_7332,N_502);
and U14349 (N_14349,N_741,N_9748);
nor U14350 (N_14350,N_7635,N_2695);
xnor U14351 (N_14351,N_6023,N_6221);
and U14352 (N_14352,N_6364,N_8452);
and U14353 (N_14353,N_9784,N_78);
nand U14354 (N_14354,N_5611,N_9408);
nand U14355 (N_14355,N_1819,N_1565);
or U14356 (N_14356,N_126,N_2546);
nor U14357 (N_14357,N_1976,N_9017);
nand U14358 (N_14358,N_7519,N_3467);
xnor U14359 (N_14359,N_7692,N_7192);
or U14360 (N_14360,N_5596,N_8008);
or U14361 (N_14361,N_7487,N_4332);
nand U14362 (N_14362,N_5292,N_7680);
nand U14363 (N_14363,N_5147,N_3344);
and U14364 (N_14364,N_9392,N_3);
nor U14365 (N_14365,N_7683,N_4479);
and U14366 (N_14366,N_6537,N_4672);
nand U14367 (N_14367,N_3143,N_3737);
nor U14368 (N_14368,N_3308,N_7597);
and U14369 (N_14369,N_97,N_3036);
or U14370 (N_14370,N_7691,N_1222);
nand U14371 (N_14371,N_4240,N_5735);
or U14372 (N_14372,N_7261,N_7205);
xor U14373 (N_14373,N_2065,N_3408);
nand U14374 (N_14374,N_8151,N_5966);
nand U14375 (N_14375,N_6917,N_7666);
or U14376 (N_14376,N_6875,N_5785);
and U14377 (N_14377,N_5867,N_9976);
nand U14378 (N_14378,N_3086,N_2316);
and U14379 (N_14379,N_9167,N_6947);
nor U14380 (N_14380,N_6930,N_162);
nor U14381 (N_14381,N_971,N_6004);
and U14382 (N_14382,N_4429,N_6911);
nor U14383 (N_14383,N_1746,N_1674);
nand U14384 (N_14384,N_868,N_8344);
and U14385 (N_14385,N_3012,N_182);
nand U14386 (N_14386,N_7764,N_9188);
and U14387 (N_14387,N_8718,N_6555);
or U14388 (N_14388,N_4510,N_9100);
or U14389 (N_14389,N_1812,N_2807);
or U14390 (N_14390,N_1574,N_4296);
nor U14391 (N_14391,N_5107,N_403);
or U14392 (N_14392,N_6924,N_790);
nor U14393 (N_14393,N_6020,N_7330);
nand U14394 (N_14394,N_8478,N_6660);
and U14395 (N_14395,N_7564,N_922);
xnor U14396 (N_14396,N_3184,N_7238);
or U14397 (N_14397,N_7339,N_8865);
and U14398 (N_14398,N_3457,N_3657);
nor U14399 (N_14399,N_887,N_5233);
xor U14400 (N_14400,N_3248,N_8434);
or U14401 (N_14401,N_3598,N_8132);
nor U14402 (N_14402,N_1904,N_6887);
nand U14403 (N_14403,N_6907,N_4190);
nand U14404 (N_14404,N_7930,N_2892);
xnor U14405 (N_14405,N_7559,N_2699);
nor U14406 (N_14406,N_2679,N_3321);
nand U14407 (N_14407,N_1641,N_1928);
nor U14408 (N_14408,N_5170,N_7022);
or U14409 (N_14409,N_8839,N_2270);
or U14410 (N_14410,N_6100,N_775);
or U14411 (N_14411,N_8521,N_6145);
xnor U14412 (N_14412,N_9981,N_124);
nor U14413 (N_14413,N_4146,N_7831);
and U14414 (N_14414,N_1861,N_4815);
and U14415 (N_14415,N_7489,N_214);
nor U14416 (N_14416,N_7718,N_5494);
nand U14417 (N_14417,N_8388,N_3541);
xor U14418 (N_14418,N_1108,N_4326);
and U14419 (N_14419,N_4070,N_12);
and U14420 (N_14420,N_8587,N_2246);
and U14421 (N_14421,N_8796,N_830);
or U14422 (N_14422,N_5267,N_5616);
xor U14423 (N_14423,N_9940,N_6434);
nor U14424 (N_14424,N_7898,N_215);
or U14425 (N_14425,N_4430,N_7687);
nor U14426 (N_14426,N_5404,N_7070);
xor U14427 (N_14427,N_9353,N_3898);
and U14428 (N_14428,N_8196,N_4055);
nand U14429 (N_14429,N_2580,N_1000);
and U14430 (N_14430,N_8054,N_3723);
or U14431 (N_14431,N_6658,N_6885);
nor U14432 (N_14432,N_2248,N_3591);
nor U14433 (N_14433,N_3369,N_1914);
nand U14434 (N_14434,N_6085,N_7982);
and U14435 (N_14435,N_4050,N_3665);
nand U14436 (N_14436,N_4407,N_1992);
xor U14437 (N_14437,N_1042,N_704);
nand U14438 (N_14438,N_5558,N_1497);
nand U14439 (N_14439,N_5483,N_9433);
and U14440 (N_14440,N_9656,N_9009);
nor U14441 (N_14441,N_1083,N_5533);
or U14442 (N_14442,N_7625,N_5836);
nor U14443 (N_14443,N_1269,N_7911);
nand U14444 (N_14444,N_2990,N_550);
nand U14445 (N_14445,N_3962,N_3735);
xnor U14446 (N_14446,N_4965,N_4943);
and U14447 (N_14447,N_1208,N_4956);
or U14448 (N_14448,N_8799,N_5493);
or U14449 (N_14449,N_9831,N_645);
xnor U14450 (N_14450,N_1328,N_4051);
xor U14451 (N_14451,N_3495,N_2594);
nor U14452 (N_14452,N_4590,N_6461);
xor U14453 (N_14453,N_1954,N_1259);
or U14454 (N_14454,N_1539,N_3409);
or U14455 (N_14455,N_1831,N_7224);
and U14456 (N_14456,N_1192,N_4851);
xnor U14457 (N_14457,N_7221,N_4980);
and U14458 (N_14458,N_1597,N_788);
nor U14459 (N_14459,N_9115,N_4824);
or U14460 (N_14460,N_1556,N_8366);
or U14461 (N_14461,N_6475,N_7276);
nor U14462 (N_14462,N_6021,N_1515);
and U14463 (N_14463,N_474,N_1845);
and U14464 (N_14464,N_7143,N_2646);
nand U14465 (N_14465,N_9498,N_6269);
xnor U14466 (N_14466,N_1039,N_4327);
xnor U14467 (N_14467,N_4828,N_2813);
and U14468 (N_14468,N_5196,N_602);
nor U14469 (N_14469,N_3469,N_1008);
nor U14470 (N_14470,N_6606,N_1967);
nor U14471 (N_14471,N_7130,N_9250);
and U14472 (N_14472,N_5385,N_5324);
or U14473 (N_14473,N_6308,N_9006);
nor U14474 (N_14474,N_6676,N_6707);
nand U14475 (N_14475,N_6823,N_8514);
xnor U14476 (N_14476,N_574,N_2186);
or U14477 (N_14477,N_458,N_2247);
or U14478 (N_14478,N_383,N_4442);
or U14479 (N_14479,N_3615,N_7338);
nor U14480 (N_14480,N_8932,N_9159);
nor U14481 (N_14481,N_8268,N_6323);
and U14482 (N_14482,N_8864,N_7780);
xor U14483 (N_14483,N_8627,N_5800);
or U14484 (N_14484,N_8257,N_8049);
or U14485 (N_14485,N_2082,N_2987);
or U14486 (N_14486,N_2165,N_2035);
and U14487 (N_14487,N_2863,N_7999);
or U14488 (N_14488,N_3576,N_7325);
nor U14489 (N_14489,N_9923,N_3716);
xnor U14490 (N_14490,N_4717,N_8417);
nor U14491 (N_14491,N_8012,N_580);
nor U14492 (N_14492,N_4056,N_1263);
xnor U14493 (N_14493,N_8494,N_2623);
and U14494 (N_14494,N_8785,N_4664);
nand U14495 (N_14495,N_3468,N_9929);
xor U14496 (N_14496,N_6581,N_781);
nor U14497 (N_14497,N_7095,N_2607);
nor U14498 (N_14498,N_9139,N_1204);
or U14499 (N_14499,N_4066,N_25);
nand U14500 (N_14500,N_8779,N_4266);
and U14501 (N_14501,N_9505,N_5161);
or U14502 (N_14502,N_6215,N_9623);
nand U14503 (N_14503,N_4111,N_5302);
or U14504 (N_14504,N_6186,N_3461);
xor U14505 (N_14505,N_9187,N_379);
and U14506 (N_14506,N_8872,N_5136);
or U14507 (N_14507,N_691,N_3263);
nor U14508 (N_14508,N_9927,N_4173);
nor U14509 (N_14509,N_1762,N_710);
nand U14510 (N_14510,N_2845,N_3637);
and U14511 (N_14511,N_6065,N_6001);
and U14512 (N_14512,N_6051,N_6428);
or U14513 (N_14513,N_1948,N_3927);
nor U14514 (N_14514,N_9708,N_1437);
xor U14515 (N_14515,N_9400,N_4106);
nand U14516 (N_14516,N_8035,N_9245);
nand U14517 (N_14517,N_8002,N_4418);
and U14518 (N_14518,N_8918,N_3471);
and U14519 (N_14519,N_5015,N_6180);
nand U14520 (N_14520,N_2597,N_9559);
nand U14521 (N_14521,N_5712,N_9912);
nor U14522 (N_14522,N_2459,N_213);
and U14523 (N_14523,N_4459,N_4626);
xor U14524 (N_14524,N_3563,N_1476);
nand U14525 (N_14525,N_3678,N_3725);
or U14526 (N_14526,N_6279,N_6638);
nor U14527 (N_14527,N_7877,N_1411);
xor U14528 (N_14528,N_4254,N_2095);
nor U14529 (N_14529,N_1065,N_1307);
and U14530 (N_14530,N_3865,N_9713);
and U14531 (N_14531,N_892,N_5100);
and U14532 (N_14532,N_7001,N_610);
xor U14533 (N_14533,N_7643,N_7028);
nand U14534 (N_14534,N_2181,N_2864);
xor U14535 (N_14535,N_2652,N_208);
xnor U14536 (N_14536,N_4197,N_8286);
or U14537 (N_14537,N_194,N_7226);
or U14538 (N_14538,N_1297,N_1308);
or U14539 (N_14539,N_7890,N_6189);
and U14540 (N_14540,N_9672,N_7929);
or U14541 (N_14541,N_909,N_8711);
nand U14542 (N_14542,N_9461,N_8657);
and U14543 (N_14543,N_2398,N_5245);
xor U14544 (N_14544,N_421,N_2587);
and U14545 (N_14545,N_181,N_9703);
nand U14546 (N_14546,N_4097,N_2168);
nand U14547 (N_14547,N_9502,N_1912);
or U14548 (N_14548,N_4263,N_7685);
nor U14549 (N_14549,N_814,N_9384);
or U14550 (N_14550,N_7296,N_5878);
nor U14551 (N_14551,N_9489,N_1265);
nor U14552 (N_14552,N_8797,N_1608);
nor U14553 (N_14553,N_1827,N_7513);
nand U14554 (N_14554,N_4801,N_5988);
and U14555 (N_14555,N_9547,N_2486);
or U14556 (N_14556,N_8121,N_5334);
nor U14557 (N_14557,N_3131,N_2808);
or U14558 (N_14558,N_4408,N_5879);
xnor U14559 (N_14559,N_837,N_5582);
xnor U14560 (N_14560,N_7993,N_5087);
nand U14561 (N_14561,N_1156,N_5224);
nor U14562 (N_14562,N_6011,N_2815);
or U14563 (N_14563,N_26,N_7318);
xor U14564 (N_14564,N_8246,N_870);
xor U14565 (N_14565,N_7897,N_4110);
and U14566 (N_14566,N_8580,N_4334);
nor U14567 (N_14567,N_7285,N_5685);
or U14568 (N_14568,N_6616,N_7359);
or U14569 (N_14569,N_724,N_9701);
and U14570 (N_14570,N_5250,N_6710);
nor U14571 (N_14571,N_6541,N_6750);
xor U14572 (N_14572,N_9954,N_897);
nand U14573 (N_14573,N_2529,N_1664);
and U14574 (N_14574,N_2528,N_6210);
nor U14575 (N_14575,N_5560,N_6232);
nand U14576 (N_14576,N_1346,N_9172);
nor U14577 (N_14577,N_4734,N_2268);
nand U14578 (N_14578,N_6722,N_6795);
xor U14579 (N_14579,N_6524,N_5865);
nand U14580 (N_14580,N_5676,N_883);
xor U14581 (N_14581,N_3612,N_9893);
or U14582 (N_14582,N_394,N_7262);
xor U14583 (N_14583,N_8342,N_5039);
or U14584 (N_14584,N_9175,N_5167);
nor U14585 (N_14585,N_7719,N_7227);
nand U14586 (N_14586,N_7287,N_5474);
or U14587 (N_14587,N_7862,N_1486);
nand U14588 (N_14588,N_6682,N_5931);
nand U14589 (N_14589,N_6109,N_7735);
and U14590 (N_14590,N_7413,N_491);
xor U14591 (N_14591,N_3274,N_3658);
or U14592 (N_14592,N_6719,N_6699);
xor U14593 (N_14593,N_7337,N_7288);
nor U14594 (N_14594,N_1158,N_589);
xor U14595 (N_14595,N_4269,N_881);
and U14596 (N_14596,N_9466,N_5997);
and U14597 (N_14597,N_4123,N_2804);
nand U14598 (N_14598,N_9615,N_9022);
nor U14599 (N_14599,N_5844,N_5049);
or U14600 (N_14600,N_191,N_5946);
xor U14601 (N_14601,N_712,N_2870);
xor U14602 (N_14602,N_5557,N_9595);
xnor U14603 (N_14603,N_7830,N_6738);
xnor U14604 (N_14604,N_603,N_5985);
nor U14605 (N_14605,N_104,N_1843);
xor U14606 (N_14606,N_7845,N_8290);
or U14607 (N_14607,N_3316,N_5451);
or U14608 (N_14608,N_4082,N_7290);
xnor U14609 (N_14609,N_484,N_6827);
and U14610 (N_14610,N_2907,N_800);
nand U14611 (N_14611,N_2756,N_5699);
and U14612 (N_14612,N_4099,N_5690);
nand U14613 (N_14613,N_2728,N_2047);
or U14614 (N_14614,N_1871,N_6536);
nand U14615 (N_14615,N_3041,N_85);
nor U14616 (N_14616,N_3672,N_4555);
nor U14617 (N_14617,N_1462,N_7282);
and U14618 (N_14618,N_9314,N_106);
and U14619 (N_14619,N_2830,N_2106);
and U14620 (N_14620,N_7140,N_6043);
nand U14621 (N_14621,N_2885,N_384);
xnor U14622 (N_14622,N_456,N_2933);
nand U14623 (N_14623,N_9779,N_6301);
and U14624 (N_14624,N_7468,N_221);
or U14625 (N_14625,N_7938,N_9153);
xnor U14626 (N_14626,N_9146,N_7522);
xor U14627 (N_14627,N_3718,N_8709);
and U14628 (N_14628,N_3660,N_9792);
nand U14629 (N_14629,N_6400,N_8544);
nand U14630 (N_14630,N_667,N_4320);
nand U14631 (N_14631,N_1417,N_5570);
xnor U14632 (N_14632,N_3477,N_430);
and U14633 (N_14633,N_3116,N_1343);
and U14634 (N_14634,N_6223,N_2776);
xor U14635 (N_14635,N_1932,N_5636);
xor U14636 (N_14636,N_2490,N_2951);
xnor U14637 (N_14637,N_5338,N_1103);
or U14638 (N_14638,N_7527,N_8507);
nor U14639 (N_14639,N_9537,N_1923);
and U14640 (N_14640,N_378,N_7301);
and U14641 (N_14641,N_7895,N_5503);
nor U14642 (N_14642,N_3879,N_747);
or U14643 (N_14643,N_9065,N_4250);
or U14644 (N_14644,N_5496,N_1549);
and U14645 (N_14645,N_8769,N_2766);
and U14646 (N_14646,N_5817,N_236);
and U14647 (N_14647,N_2187,N_5958);
and U14648 (N_14648,N_9759,N_4004);
nor U14649 (N_14649,N_1434,N_4887);
and U14650 (N_14650,N_9992,N_9190);
and U14651 (N_14651,N_6248,N_5822);
or U14652 (N_14652,N_344,N_5325);
xor U14653 (N_14653,N_6106,N_4165);
nor U14654 (N_14654,N_1616,N_4707);
nor U14655 (N_14655,N_3118,N_7317);
nand U14656 (N_14656,N_9307,N_1532);
nand U14657 (N_14657,N_8499,N_4002);
and U14658 (N_14658,N_4509,N_9331);
nand U14659 (N_14659,N_8098,N_8031);
nand U14660 (N_14660,N_9866,N_5106);
nand U14661 (N_14661,N_3113,N_757);
nor U14662 (N_14662,N_5156,N_8906);
or U14663 (N_14663,N_402,N_5620);
xnor U14664 (N_14664,N_9432,N_4949);
and U14665 (N_14665,N_4134,N_9793);
and U14666 (N_14666,N_6071,N_3056);
nor U14667 (N_14667,N_8730,N_5587);
or U14668 (N_14668,N_277,N_9449);
nand U14669 (N_14669,N_166,N_5005);
xor U14670 (N_14670,N_8394,N_4215);
xnor U14671 (N_14671,N_5335,N_4239);
nor U14672 (N_14672,N_5214,N_345);
and U14673 (N_14673,N_6049,N_5749);
and U14674 (N_14674,N_4850,N_7863);
and U14675 (N_14675,N_2908,N_4747);
nor U14676 (N_14676,N_6437,N_202);
and U14677 (N_14677,N_9771,N_901);
or U14678 (N_14678,N_8552,N_7634);
and U14679 (N_14679,N_3376,N_692);
nand U14680 (N_14680,N_3661,N_9583);
xnor U14681 (N_14681,N_7663,N_3807);
nor U14682 (N_14682,N_4031,N_7504);
and U14683 (N_14683,N_1578,N_7113);
xor U14684 (N_14684,N_7825,N_8271);
xor U14685 (N_14685,N_1006,N_4010);
nor U14686 (N_14686,N_9181,N_123);
and U14687 (N_14687,N_4465,N_94);
nand U14688 (N_14688,N_6468,N_4305);
nand U14689 (N_14689,N_4840,N_7783);
xnor U14690 (N_14690,N_6137,N_9441);
nand U14691 (N_14691,N_8835,N_5024);
or U14692 (N_14692,N_801,N_4169);
xnor U14693 (N_14693,N_6142,N_619);
nand U14694 (N_14694,N_8293,N_9110);
xnor U14695 (N_14695,N_7962,N_1125);
xor U14696 (N_14696,N_8852,N_9931);
nor U14697 (N_14697,N_6283,N_9508);
and U14698 (N_14698,N_4714,N_4005);
xnor U14699 (N_14699,N_7903,N_4412);
nand U14700 (N_14700,N_8599,N_6288);
and U14701 (N_14701,N_5094,N_561);
xor U14702 (N_14702,N_8041,N_3689);
or U14703 (N_14703,N_7904,N_9688);
nand U14704 (N_14704,N_6948,N_2516);
and U14705 (N_14705,N_5037,N_1721);
or U14706 (N_14706,N_3726,N_6881);
and U14707 (N_14707,N_9211,N_7715);
nor U14708 (N_14708,N_1201,N_6033);
nand U14709 (N_14709,N_6054,N_4011);
or U14710 (N_14710,N_5193,N_753);
or U14711 (N_14711,N_9975,N_5910);
xor U14712 (N_14712,N_4915,N_4893);
nor U14713 (N_14713,N_9148,N_5993);
xnor U14714 (N_14714,N_5133,N_7945);
or U14715 (N_14715,N_2613,N_10);
xor U14716 (N_14716,N_1591,N_2522);
nor U14717 (N_14717,N_7649,N_3869);
and U14718 (N_14718,N_1956,N_3636);
xnor U14719 (N_14719,N_271,N_9218);
nor U14720 (N_14720,N_6395,N_2358);
xnor U14721 (N_14721,N_3238,N_1749);
nand U14722 (N_14722,N_677,N_925);
or U14723 (N_14723,N_684,N_7216);
or U14724 (N_14724,N_5583,N_8720);
and U14725 (N_14725,N_968,N_1598);
nor U14726 (N_14726,N_8634,N_8079);
or U14727 (N_14727,N_5466,N_2188);
xor U14728 (N_14728,N_8823,N_8234);
nand U14729 (N_14729,N_6201,N_4894);
or U14730 (N_14730,N_1040,N_5207);
nand U14731 (N_14731,N_5086,N_3331);
nand U14732 (N_14732,N_7742,N_718);
xor U14733 (N_14733,N_9557,N_9675);
nand U14734 (N_14734,N_6414,N_3040);
and U14735 (N_14735,N_1970,N_5992);
nor U14736 (N_14736,N_1571,N_2150);
nor U14737 (N_14737,N_2335,N_7744);
xnor U14738 (N_14738,N_9696,N_8612);
and U14739 (N_14739,N_7955,N_254);
and U14740 (N_14740,N_507,N_3699);
xor U14741 (N_14741,N_9151,N_8125);
nor U14742 (N_14742,N_1010,N_2388);
xor U14743 (N_14743,N_914,N_422);
and U14744 (N_14744,N_5297,N_5053);
nor U14745 (N_14745,N_3424,N_2530);
xor U14746 (N_14746,N_9970,N_252);
nor U14747 (N_14747,N_101,N_1285);
nand U14748 (N_14748,N_4449,N_4971);
nor U14749 (N_14749,N_3775,N_2162);
xnor U14750 (N_14750,N_6039,N_2576);
and U14751 (N_14751,N_5694,N_2738);
xor U14752 (N_14752,N_415,N_2799);
nand U14753 (N_14753,N_4107,N_3109);
nand U14754 (N_14754,N_3267,N_4504);
xor U14755 (N_14755,N_3044,N_3070);
nand U14756 (N_14756,N_1769,N_7969);
nand U14757 (N_14757,N_1818,N_4323);
and U14758 (N_14758,N_9826,N_6493);
and U14759 (N_14759,N_7570,N_4019);
or U14760 (N_14760,N_8485,N_391);
and U14761 (N_14761,N_9815,N_5861);
nor U14762 (N_14762,N_6320,N_4789);
or U14763 (N_14763,N_6680,N_1573);
nor U14764 (N_14764,N_2814,N_4186);
nor U14765 (N_14765,N_2539,N_9523);
or U14766 (N_14766,N_923,N_1081);
nand U14767 (N_14767,N_1850,N_8427);
or U14768 (N_14768,N_1057,N_2598);
nand U14769 (N_14769,N_253,N_4494);
xor U14770 (N_14770,N_6868,N_8097);
xor U14771 (N_14771,N_183,N_7388);
nor U14772 (N_14772,N_2589,N_7308);
and U14773 (N_14773,N_6123,N_9619);
xnor U14774 (N_14774,N_3146,N_223);
and U14775 (N_14775,N_5336,N_4570);
or U14776 (N_14776,N_5915,N_6822);
and U14777 (N_14777,N_9516,N_9500);
and U14778 (N_14778,N_5535,N_3839);
xnor U14779 (N_14779,N_2262,N_2056);
or U14780 (N_14780,N_4232,N_5713);
or U14781 (N_14781,N_1331,N_2278);
or U14782 (N_14782,N_2353,N_2282);
nand U14783 (N_14783,N_942,N_526);
nand U14784 (N_14784,N_5272,N_8030);
xnor U14785 (N_14785,N_9407,N_9740);
xnor U14786 (N_14786,N_3594,N_3559);
or U14787 (N_14787,N_279,N_9410);
and U14788 (N_14788,N_3797,N_285);
or U14789 (N_14789,N_4208,N_8263);
nand U14790 (N_14790,N_7209,N_2925);
and U14791 (N_14791,N_8084,N_1315);
nand U14792 (N_14792,N_3333,N_1774);
xor U14793 (N_14793,N_6230,N_543);
nand U14794 (N_14794,N_5886,N_1267);
nand U14795 (N_14795,N_6869,N_8447);
or U14796 (N_14796,N_2293,N_5007);
xnor U14797 (N_14797,N_8046,N_7997);
or U14798 (N_14798,N_6626,N_6979);
nor U14799 (N_14799,N_5091,N_3454);
and U14800 (N_14800,N_5911,N_8498);
nor U14801 (N_14801,N_1098,N_6742);
nand U14802 (N_14802,N_406,N_4447);
and U14803 (N_14803,N_2625,N_5229);
and U14804 (N_14804,N_7463,N_7465);
xor U14805 (N_14805,N_7364,N_6720);
nand U14806 (N_14806,N_5112,N_7439);
nand U14807 (N_14807,N_627,N_5804);
nor U14808 (N_14808,N_8894,N_9634);
and U14809 (N_14809,N_5055,N_4557);
xnor U14810 (N_14810,N_4370,N_7858);
nand U14811 (N_14811,N_8353,N_1798);
nand U14812 (N_14812,N_3038,N_1797);
and U14813 (N_14813,N_4904,N_4427);
nor U14814 (N_14814,N_8786,N_3008);
nor U14815 (N_14815,N_3002,N_1387);
and U14816 (N_14816,N_6429,N_1622);
and U14817 (N_14817,N_4540,N_7013);
or U14818 (N_14818,N_1750,N_2705);
nand U14819 (N_14819,N_5160,N_1835);
xor U14820 (N_14820,N_7412,N_639);
xnor U14821 (N_14821,N_7090,N_5289);
nand U14822 (N_14822,N_5859,N_2376);
nor U14823 (N_14823,N_4389,N_2237);
nor U14824 (N_14824,N_6206,N_7165);
nand U14825 (N_14825,N_4666,N_2447);
nor U14826 (N_14826,N_349,N_4998);
or U14827 (N_14827,N_2365,N_3892);
nand U14828 (N_14828,N_7773,N_829);
or U14829 (N_14829,N_2651,N_9130);
or U14830 (N_14830,N_4195,N_9871);
and U14831 (N_14831,N_6547,N_4740);
nor U14832 (N_14832,N_8430,N_9677);
and U14833 (N_14833,N_9335,N_68);
xor U14834 (N_14834,N_5778,N_7418);
xor U14835 (N_14835,N_7517,N_6957);
nor U14836 (N_14836,N_2758,N_6787);
xnor U14837 (N_14837,N_4653,N_3160);
xor U14838 (N_14838,N_6981,N_6899);
and U14839 (N_14839,N_351,N_361);
nand U14840 (N_14840,N_7554,N_5782);
nor U14841 (N_14841,N_2108,N_8364);
or U14842 (N_14842,N_995,N_6116);
nor U14843 (N_14843,N_1177,N_911);
and U14844 (N_14844,N_9682,N_9889);
nand U14845 (N_14845,N_9276,N_4089);
or U14846 (N_14846,N_2227,N_5729);
or U14847 (N_14847,N_4733,N_5262);
or U14848 (N_14848,N_6203,N_8218);
or U14849 (N_14849,N_5526,N_7842);
or U14850 (N_14850,N_7235,N_1022);
and U14851 (N_14851,N_6451,N_7503);
nor U14852 (N_14852,N_3956,N_8156);
xnor U14853 (N_14853,N_8641,N_7601);
nand U14854 (N_14854,N_4094,N_7684);
or U14855 (N_14855,N_3695,N_8383);
and U14856 (N_14856,N_2113,N_8244);
or U14857 (N_14857,N_8055,N_1164);
or U14858 (N_14858,N_4281,N_5347);
nand U14859 (N_14859,N_2354,N_1584);
nor U14860 (N_14860,N_5188,N_3410);
nor U14861 (N_14861,N_8415,N_4222);
xnor U14862 (N_14862,N_583,N_3214);
nand U14863 (N_14863,N_2523,N_632);
or U14864 (N_14864,N_1469,N_6759);
xor U14865 (N_14865,N_3023,N_3730);
or U14866 (N_14866,N_5525,N_5058);
or U14867 (N_14867,N_6295,N_6489);
or U14868 (N_14868,N_2054,N_3908);
nor U14869 (N_14869,N_6661,N_454);
nand U14870 (N_14870,N_6163,N_4710);
nand U14871 (N_14871,N_1852,N_8630);
nand U14872 (N_14872,N_8683,N_1302);
nor U14873 (N_14873,N_953,N_3833);
xnor U14874 (N_14874,N_2052,N_8180);
nand U14875 (N_14875,N_4617,N_7481);
and U14876 (N_14876,N_7471,N_4608);
nand U14877 (N_14877,N_7854,N_7662);
nor U14878 (N_14878,N_5323,N_7926);
xnor U14879 (N_14879,N_8788,N_1454);
nor U14880 (N_14880,N_5891,N_2572);
nand U14881 (N_14881,N_2750,N_8496);
and U14882 (N_14882,N_7180,N_3851);
nand U14883 (N_14883,N_664,N_4563);
xor U14884 (N_14884,N_2100,N_8050);
nor U14885 (N_14885,N_839,N_8248);
or U14886 (N_14886,N_6811,N_7887);
and U14887 (N_14887,N_6498,N_6830);
xnor U14888 (N_14888,N_4451,N_9013);
nor U14889 (N_14889,N_1575,N_3476);
and U14890 (N_14890,N_1779,N_9733);
nor U14891 (N_14891,N_557,N_3390);
xor U14892 (N_14892,N_784,N_9816);
xor U14893 (N_14893,N_7004,N_9894);
nor U14894 (N_14894,N_218,N_8900);
and U14895 (N_14895,N_9385,N_4036);
nor U14896 (N_14896,N_2498,N_4922);
xnor U14897 (N_14897,N_2540,N_7260);
xor U14898 (N_14898,N_2671,N_5615);
xnor U14899 (N_14899,N_1077,N_4229);
and U14900 (N_14900,N_4310,N_4579);
nor U14901 (N_14901,N_1122,N_8533);
xnor U14902 (N_14902,N_8087,N_8086);
and U14903 (N_14903,N_7706,N_3341);
xor U14904 (N_14904,N_8876,N_1310);
nor U14905 (N_14905,N_8915,N_6865);
or U14906 (N_14906,N_5506,N_4741);
or U14907 (N_14907,N_5344,N_8744);
and U14908 (N_14908,N_5498,N_5280);
and U14909 (N_14909,N_5487,N_9926);
nand U14910 (N_14910,N_7024,N_4721);
nor U14911 (N_14911,N_8088,N_2828);
nand U14912 (N_14912,N_4448,N_5802);
xor U14913 (N_14913,N_1646,N_2027);
xnor U14914 (N_14914,N_9974,N_3172);
nand U14915 (N_14915,N_9544,N_5320);
or U14916 (N_14916,N_268,N_407);
and U14917 (N_14917,N_1117,N_7839);
nor U14918 (N_14918,N_3249,N_2114);
nand U14919 (N_14919,N_5856,N_568);
xor U14920 (N_14920,N_5928,N_4623);
nand U14921 (N_14921,N_3359,N_8551);
xnor U14922 (N_14922,N_2379,N_7360);
or U14923 (N_14923,N_5687,N_9478);
nor U14924 (N_14924,N_2410,N_576);
or U14925 (N_14925,N_2327,N_707);
and U14926 (N_14926,N_1745,N_7893);
nor U14927 (N_14927,N_4286,N_9236);
nand U14928 (N_14928,N_7256,N_1013);
or U14929 (N_14929,N_9395,N_3448);
or U14930 (N_14930,N_2477,N_6629);
xnor U14931 (N_14931,N_4994,N_8644);
nor U14932 (N_14932,N_8854,N_3277);
nor U14933 (N_14933,N_8673,N_4172);
nor U14934 (N_14934,N_6148,N_8172);
xor U14935 (N_14935,N_3850,N_9057);
nand U14936 (N_14936,N_9729,N_2006);
nand U14937 (N_14937,N_9053,N_4360);
nor U14938 (N_14938,N_3135,N_8385);
or U14939 (N_14939,N_2275,N_1341);
xor U14940 (N_14940,N_9873,N_8790);
xnor U14941 (N_14941,N_9286,N_9240);
and U14942 (N_14942,N_6748,N_1319);
and U14943 (N_14943,N_9479,N_4529);
nand U14944 (N_14944,N_5132,N_7425);
nand U14945 (N_14945,N_6712,N_1110);
and U14946 (N_14946,N_1260,N_1960);
or U14947 (N_14947,N_523,N_725);
nor U14948 (N_14948,N_4614,N_7753);
nand U14949 (N_14949,N_4315,N_1739);
xnor U14950 (N_14950,N_9756,N_3582);
nor U14951 (N_14951,N_8266,N_7551);
xor U14952 (N_14952,N_1218,N_6973);
nor U14953 (N_14953,N_2189,N_2697);
nand U14954 (N_14954,N_9421,N_9128);
and U14955 (N_14955,N_681,N_9258);
and U14956 (N_14956,N_7859,N_7805);
nand U14957 (N_14957,N_1141,N_9306);
or U14958 (N_14958,N_7233,N_5564);
and U14959 (N_14959,N_7477,N_8607);
or U14960 (N_14960,N_7452,N_1980);
nor U14961 (N_14961,N_9915,N_7834);
nand U14962 (N_14962,N_3309,N_2326);
and U14963 (N_14963,N_2357,N_3738);
or U14964 (N_14964,N_8410,N_6424);
or U14965 (N_14965,N_7480,N_2782);
nor U14966 (N_14966,N_388,N_3881);
and U14967 (N_14967,N_4984,N_552);
xor U14968 (N_14968,N_9143,N_4771);
and U14969 (N_14969,N_4378,N_7062);
nor U14970 (N_14970,N_7484,N_3412);
or U14971 (N_14971,N_9228,N_2554);
nor U14972 (N_14972,N_7721,N_3404);
and U14973 (N_14973,N_4790,N_8840);
or U14974 (N_14974,N_14,N_4659);
nor U14975 (N_14975,N_4129,N_1471);
xor U14976 (N_14976,N_4934,N_9892);
nor U14977 (N_14977,N_2359,N_1736);
or U14978 (N_14978,N_5601,N_8515);
or U14979 (N_14979,N_5296,N_6597);
nand U14980 (N_14980,N_9668,N_1283);
and U14981 (N_14981,N_1978,N_1621);
xnor U14982 (N_14982,N_6681,N_4008);
and U14983 (N_14983,N_6529,N_2223);
xnor U14984 (N_14984,N_5929,N_9908);
nor U14985 (N_14985,N_4072,N_1700);
and U14986 (N_14986,N_6833,N_5472);
and U14987 (N_14987,N_6060,N_3022);
or U14988 (N_14988,N_7580,N_4034);
and U14989 (N_14989,N_7326,N_5693);
and U14990 (N_14990,N_6102,N_3823);
nor U14991 (N_14991,N_7255,N_8215);
nand U14992 (N_14992,N_1146,N_4951);
and U14993 (N_14993,N_4268,N_9267);
nor U14994 (N_14994,N_2132,N_9436);
nand U14995 (N_14995,N_9809,N_2397);
xor U14996 (N_14996,N_9338,N_7429);
and U14997 (N_14997,N_9588,N_1903);
nand U14998 (N_14998,N_7775,N_8858);
nand U14999 (N_14999,N_2356,N_8725);
or U15000 (N_15000,N_9533,N_9745);
nand U15001 (N_15001,N_9171,N_2376);
or U15002 (N_15002,N_819,N_1091);
nor U15003 (N_15003,N_5374,N_5676);
xnor U15004 (N_15004,N_8740,N_1872);
xor U15005 (N_15005,N_5035,N_9745);
or U15006 (N_15006,N_3754,N_8745);
xnor U15007 (N_15007,N_3452,N_1302);
nor U15008 (N_15008,N_9926,N_500);
nand U15009 (N_15009,N_8230,N_263);
nor U15010 (N_15010,N_2146,N_8048);
xnor U15011 (N_15011,N_5071,N_8740);
xnor U15012 (N_15012,N_9531,N_4231);
and U15013 (N_15013,N_5703,N_8021);
and U15014 (N_15014,N_7967,N_5152);
xor U15015 (N_15015,N_3156,N_2191);
nand U15016 (N_15016,N_3913,N_8484);
nand U15017 (N_15017,N_2391,N_5795);
nand U15018 (N_15018,N_7275,N_4464);
xnor U15019 (N_15019,N_5970,N_4604);
or U15020 (N_15020,N_5117,N_4636);
xor U15021 (N_15021,N_6422,N_9292);
or U15022 (N_15022,N_7585,N_4793);
xor U15023 (N_15023,N_3490,N_2923);
nor U15024 (N_15024,N_6878,N_477);
and U15025 (N_15025,N_2893,N_3844);
nor U15026 (N_15026,N_7415,N_2793);
or U15027 (N_15027,N_8720,N_7462);
and U15028 (N_15028,N_5487,N_4773);
and U15029 (N_15029,N_4794,N_2537);
or U15030 (N_15030,N_1983,N_3374);
and U15031 (N_15031,N_5165,N_4747);
nand U15032 (N_15032,N_1782,N_8843);
xnor U15033 (N_15033,N_2672,N_1411);
xnor U15034 (N_15034,N_8724,N_8082);
nor U15035 (N_15035,N_5984,N_4069);
and U15036 (N_15036,N_5830,N_4823);
xor U15037 (N_15037,N_4141,N_5448);
and U15038 (N_15038,N_9994,N_7781);
or U15039 (N_15039,N_9685,N_4346);
nand U15040 (N_15040,N_7850,N_1405);
nand U15041 (N_15041,N_1090,N_127);
nor U15042 (N_15042,N_8080,N_3813);
nand U15043 (N_15043,N_9788,N_5066);
or U15044 (N_15044,N_2738,N_7183);
nor U15045 (N_15045,N_6144,N_128);
nand U15046 (N_15046,N_4130,N_755);
xor U15047 (N_15047,N_6460,N_185);
and U15048 (N_15048,N_5956,N_910);
and U15049 (N_15049,N_8331,N_7853);
nand U15050 (N_15050,N_7076,N_1797);
xnor U15051 (N_15051,N_5788,N_2696);
and U15052 (N_15052,N_6221,N_7568);
nand U15053 (N_15053,N_4827,N_5501);
and U15054 (N_15054,N_6571,N_9583);
xnor U15055 (N_15055,N_5695,N_3322);
nand U15056 (N_15056,N_1034,N_2468);
and U15057 (N_15057,N_4356,N_5560);
xor U15058 (N_15058,N_1535,N_522);
xnor U15059 (N_15059,N_3878,N_3261);
nor U15060 (N_15060,N_447,N_279);
xor U15061 (N_15061,N_3883,N_7088);
xor U15062 (N_15062,N_1874,N_6438);
nand U15063 (N_15063,N_7565,N_4244);
nand U15064 (N_15064,N_3199,N_2741);
xor U15065 (N_15065,N_4196,N_7614);
nand U15066 (N_15066,N_6522,N_8000);
and U15067 (N_15067,N_8207,N_7932);
or U15068 (N_15068,N_5823,N_8111);
and U15069 (N_15069,N_9138,N_8784);
nor U15070 (N_15070,N_5247,N_9853);
nor U15071 (N_15071,N_2290,N_7540);
nand U15072 (N_15072,N_2472,N_2063);
nor U15073 (N_15073,N_5351,N_5044);
nand U15074 (N_15074,N_9741,N_4562);
or U15075 (N_15075,N_5616,N_8319);
xnor U15076 (N_15076,N_8767,N_6316);
nand U15077 (N_15077,N_4124,N_7454);
nand U15078 (N_15078,N_904,N_9814);
or U15079 (N_15079,N_7018,N_3490);
xor U15080 (N_15080,N_8353,N_5957);
and U15081 (N_15081,N_3525,N_9156);
nor U15082 (N_15082,N_2040,N_7937);
xnor U15083 (N_15083,N_6209,N_4208);
or U15084 (N_15084,N_5977,N_2428);
nand U15085 (N_15085,N_9341,N_5499);
xnor U15086 (N_15086,N_6942,N_9468);
xor U15087 (N_15087,N_794,N_2178);
nand U15088 (N_15088,N_8606,N_6687);
xnor U15089 (N_15089,N_8694,N_4621);
nor U15090 (N_15090,N_5922,N_7889);
and U15091 (N_15091,N_6251,N_6364);
nand U15092 (N_15092,N_7837,N_3169);
nand U15093 (N_15093,N_3370,N_2360);
nor U15094 (N_15094,N_4854,N_3357);
and U15095 (N_15095,N_572,N_4598);
nand U15096 (N_15096,N_6028,N_9158);
xnor U15097 (N_15097,N_7745,N_4027);
xnor U15098 (N_15098,N_5976,N_9145);
xnor U15099 (N_15099,N_7956,N_7000);
and U15100 (N_15100,N_1052,N_429);
or U15101 (N_15101,N_4873,N_779);
and U15102 (N_15102,N_4671,N_4225);
and U15103 (N_15103,N_1300,N_3813);
nor U15104 (N_15104,N_467,N_4687);
xnor U15105 (N_15105,N_681,N_4756);
and U15106 (N_15106,N_7386,N_8278);
and U15107 (N_15107,N_6452,N_2523);
or U15108 (N_15108,N_2601,N_868);
xor U15109 (N_15109,N_7455,N_5610);
nor U15110 (N_15110,N_7356,N_3147);
or U15111 (N_15111,N_7620,N_4183);
xnor U15112 (N_15112,N_2825,N_6887);
and U15113 (N_15113,N_7999,N_486);
nor U15114 (N_15114,N_2433,N_1368);
xnor U15115 (N_15115,N_8173,N_2528);
nor U15116 (N_15116,N_8591,N_8272);
and U15117 (N_15117,N_2998,N_4528);
and U15118 (N_15118,N_8297,N_3205);
xnor U15119 (N_15119,N_945,N_2650);
and U15120 (N_15120,N_9192,N_4813);
nand U15121 (N_15121,N_7282,N_9711);
and U15122 (N_15122,N_4735,N_9783);
or U15123 (N_15123,N_4485,N_3535);
nor U15124 (N_15124,N_5573,N_8150);
and U15125 (N_15125,N_9545,N_7604);
or U15126 (N_15126,N_5307,N_6711);
nor U15127 (N_15127,N_1014,N_2277);
nor U15128 (N_15128,N_282,N_6837);
nor U15129 (N_15129,N_7075,N_2337);
or U15130 (N_15130,N_4365,N_8934);
xnor U15131 (N_15131,N_548,N_6538);
or U15132 (N_15132,N_1934,N_7827);
or U15133 (N_15133,N_6186,N_7286);
and U15134 (N_15134,N_9972,N_3653);
or U15135 (N_15135,N_6276,N_644);
and U15136 (N_15136,N_3140,N_8299);
nand U15137 (N_15137,N_3121,N_5382);
xor U15138 (N_15138,N_9553,N_324);
nor U15139 (N_15139,N_6017,N_9108);
nand U15140 (N_15140,N_7801,N_9868);
nor U15141 (N_15141,N_447,N_5645);
or U15142 (N_15142,N_7331,N_975);
nand U15143 (N_15143,N_7237,N_5956);
nor U15144 (N_15144,N_4080,N_8135);
nand U15145 (N_15145,N_3564,N_9323);
nor U15146 (N_15146,N_424,N_2769);
nand U15147 (N_15147,N_4323,N_6596);
or U15148 (N_15148,N_9300,N_1965);
or U15149 (N_15149,N_2831,N_5633);
nor U15150 (N_15150,N_7254,N_6779);
nand U15151 (N_15151,N_1106,N_2257);
and U15152 (N_15152,N_3423,N_789);
xor U15153 (N_15153,N_1011,N_4801);
and U15154 (N_15154,N_955,N_7183);
or U15155 (N_15155,N_9270,N_7607);
and U15156 (N_15156,N_24,N_6691);
nand U15157 (N_15157,N_5722,N_4450);
and U15158 (N_15158,N_3437,N_698);
or U15159 (N_15159,N_5971,N_2783);
or U15160 (N_15160,N_596,N_6366);
nor U15161 (N_15161,N_1704,N_3247);
xor U15162 (N_15162,N_8619,N_4015);
xnor U15163 (N_15163,N_2596,N_6598);
nand U15164 (N_15164,N_692,N_3672);
nor U15165 (N_15165,N_1444,N_8956);
nand U15166 (N_15166,N_9649,N_6559);
nand U15167 (N_15167,N_5403,N_5683);
nand U15168 (N_15168,N_2026,N_7774);
and U15169 (N_15169,N_919,N_5047);
and U15170 (N_15170,N_6988,N_6771);
xnor U15171 (N_15171,N_6896,N_7078);
nor U15172 (N_15172,N_590,N_3061);
and U15173 (N_15173,N_6328,N_4647);
and U15174 (N_15174,N_8355,N_4030);
nor U15175 (N_15175,N_7352,N_7284);
xor U15176 (N_15176,N_8939,N_7540);
nor U15177 (N_15177,N_7143,N_6153);
xor U15178 (N_15178,N_8127,N_5479);
nor U15179 (N_15179,N_4244,N_6195);
nand U15180 (N_15180,N_9260,N_8349);
nand U15181 (N_15181,N_5385,N_3235);
nor U15182 (N_15182,N_8304,N_9622);
or U15183 (N_15183,N_881,N_4740);
or U15184 (N_15184,N_9825,N_5445);
nor U15185 (N_15185,N_7324,N_818);
or U15186 (N_15186,N_7980,N_72);
xor U15187 (N_15187,N_10,N_5246);
xnor U15188 (N_15188,N_2246,N_6336);
xor U15189 (N_15189,N_5268,N_6106);
or U15190 (N_15190,N_2252,N_9628);
or U15191 (N_15191,N_6151,N_9593);
nor U15192 (N_15192,N_4073,N_2032);
and U15193 (N_15193,N_4283,N_3609);
and U15194 (N_15194,N_1101,N_6306);
nand U15195 (N_15195,N_2707,N_2525);
or U15196 (N_15196,N_3876,N_2245);
nor U15197 (N_15197,N_3835,N_7889);
nor U15198 (N_15198,N_5379,N_2371);
xor U15199 (N_15199,N_4637,N_5869);
xnor U15200 (N_15200,N_1937,N_1983);
and U15201 (N_15201,N_5885,N_1460);
nand U15202 (N_15202,N_8266,N_6355);
or U15203 (N_15203,N_2816,N_585);
and U15204 (N_15204,N_6273,N_5707);
or U15205 (N_15205,N_4796,N_357);
xor U15206 (N_15206,N_2183,N_9158);
or U15207 (N_15207,N_9593,N_592);
nor U15208 (N_15208,N_7977,N_1214);
nor U15209 (N_15209,N_4382,N_2664);
xor U15210 (N_15210,N_4878,N_9394);
nand U15211 (N_15211,N_266,N_6355);
nand U15212 (N_15212,N_5015,N_9002);
xnor U15213 (N_15213,N_4101,N_4986);
nor U15214 (N_15214,N_3128,N_9151);
nor U15215 (N_15215,N_4854,N_2954);
or U15216 (N_15216,N_5892,N_6303);
nand U15217 (N_15217,N_1927,N_8083);
xnor U15218 (N_15218,N_9596,N_6753);
or U15219 (N_15219,N_1308,N_5588);
nand U15220 (N_15220,N_8840,N_9585);
nand U15221 (N_15221,N_1695,N_5365);
or U15222 (N_15222,N_8377,N_909);
or U15223 (N_15223,N_7216,N_8956);
and U15224 (N_15224,N_1498,N_2689);
nor U15225 (N_15225,N_8262,N_8285);
and U15226 (N_15226,N_3149,N_3739);
nor U15227 (N_15227,N_7333,N_2254);
and U15228 (N_15228,N_802,N_7976);
nand U15229 (N_15229,N_8286,N_6697);
and U15230 (N_15230,N_8530,N_2328);
and U15231 (N_15231,N_8958,N_3722);
nand U15232 (N_15232,N_7597,N_4420);
nor U15233 (N_15233,N_5058,N_1122);
and U15234 (N_15234,N_6927,N_3533);
and U15235 (N_15235,N_6055,N_1931);
and U15236 (N_15236,N_6768,N_4059);
nand U15237 (N_15237,N_6946,N_9156);
or U15238 (N_15238,N_8416,N_9663);
nand U15239 (N_15239,N_3270,N_7897);
nor U15240 (N_15240,N_878,N_2752);
nor U15241 (N_15241,N_722,N_350);
or U15242 (N_15242,N_8936,N_9125);
xnor U15243 (N_15243,N_7918,N_3691);
and U15244 (N_15244,N_5838,N_1093);
or U15245 (N_15245,N_6043,N_861);
nand U15246 (N_15246,N_1048,N_6011);
nand U15247 (N_15247,N_1429,N_6356);
nor U15248 (N_15248,N_938,N_5138);
nand U15249 (N_15249,N_2978,N_1542);
xor U15250 (N_15250,N_5503,N_5656);
nor U15251 (N_15251,N_4294,N_1698);
nor U15252 (N_15252,N_2818,N_2023);
xor U15253 (N_15253,N_3582,N_82);
xor U15254 (N_15254,N_5302,N_5710);
xnor U15255 (N_15255,N_7171,N_168);
nand U15256 (N_15256,N_2721,N_7246);
nor U15257 (N_15257,N_7997,N_7958);
and U15258 (N_15258,N_3675,N_3032);
xnor U15259 (N_15259,N_4401,N_623);
xor U15260 (N_15260,N_1507,N_4410);
nor U15261 (N_15261,N_8869,N_820);
or U15262 (N_15262,N_5126,N_8265);
xnor U15263 (N_15263,N_7454,N_3572);
nand U15264 (N_15264,N_2299,N_3302);
or U15265 (N_15265,N_7764,N_9606);
xor U15266 (N_15266,N_3977,N_134);
xor U15267 (N_15267,N_1569,N_9441);
nor U15268 (N_15268,N_6366,N_9245);
nand U15269 (N_15269,N_5067,N_4601);
or U15270 (N_15270,N_9003,N_5265);
nor U15271 (N_15271,N_971,N_4153);
and U15272 (N_15272,N_9349,N_8533);
or U15273 (N_15273,N_6069,N_9640);
xor U15274 (N_15274,N_4385,N_1173);
nand U15275 (N_15275,N_5542,N_1287);
and U15276 (N_15276,N_8237,N_1927);
nor U15277 (N_15277,N_2580,N_696);
nand U15278 (N_15278,N_9884,N_4793);
or U15279 (N_15279,N_5690,N_4343);
or U15280 (N_15280,N_8449,N_5111);
and U15281 (N_15281,N_6962,N_7488);
nor U15282 (N_15282,N_3625,N_5246);
nor U15283 (N_15283,N_1699,N_1602);
or U15284 (N_15284,N_5438,N_3505);
nor U15285 (N_15285,N_994,N_3981);
xnor U15286 (N_15286,N_1361,N_1227);
xnor U15287 (N_15287,N_1374,N_3575);
or U15288 (N_15288,N_4783,N_3124);
or U15289 (N_15289,N_5722,N_2283);
nand U15290 (N_15290,N_2460,N_8090);
xnor U15291 (N_15291,N_3075,N_2053);
and U15292 (N_15292,N_2102,N_6945);
or U15293 (N_15293,N_5962,N_5683);
or U15294 (N_15294,N_3001,N_784);
nand U15295 (N_15295,N_4071,N_2095);
or U15296 (N_15296,N_8566,N_8529);
or U15297 (N_15297,N_4625,N_7733);
nor U15298 (N_15298,N_3324,N_7581);
nor U15299 (N_15299,N_9401,N_2553);
nor U15300 (N_15300,N_5516,N_6047);
xor U15301 (N_15301,N_6568,N_2893);
nand U15302 (N_15302,N_3196,N_5277);
and U15303 (N_15303,N_955,N_2061);
nand U15304 (N_15304,N_356,N_8316);
xnor U15305 (N_15305,N_3444,N_7360);
and U15306 (N_15306,N_7848,N_3829);
nor U15307 (N_15307,N_3291,N_1213);
nand U15308 (N_15308,N_5252,N_2628);
or U15309 (N_15309,N_940,N_9884);
or U15310 (N_15310,N_5946,N_9340);
nand U15311 (N_15311,N_7830,N_1458);
and U15312 (N_15312,N_6749,N_3194);
nand U15313 (N_15313,N_896,N_8678);
or U15314 (N_15314,N_685,N_2105);
and U15315 (N_15315,N_8766,N_4787);
nand U15316 (N_15316,N_8557,N_5947);
or U15317 (N_15317,N_4553,N_2254);
nand U15318 (N_15318,N_3895,N_1507);
or U15319 (N_15319,N_4772,N_9870);
nand U15320 (N_15320,N_8843,N_8192);
xor U15321 (N_15321,N_2877,N_9172);
nand U15322 (N_15322,N_8287,N_1592);
nand U15323 (N_15323,N_4584,N_260);
xor U15324 (N_15324,N_9918,N_7727);
or U15325 (N_15325,N_4352,N_945);
and U15326 (N_15326,N_6449,N_3978);
xnor U15327 (N_15327,N_5394,N_4745);
xor U15328 (N_15328,N_553,N_6348);
nand U15329 (N_15329,N_165,N_8932);
and U15330 (N_15330,N_1361,N_3526);
or U15331 (N_15331,N_400,N_1348);
and U15332 (N_15332,N_6466,N_7184);
and U15333 (N_15333,N_5823,N_6632);
xor U15334 (N_15334,N_5361,N_1672);
nand U15335 (N_15335,N_5874,N_4275);
or U15336 (N_15336,N_5515,N_7802);
nand U15337 (N_15337,N_6128,N_2590);
xor U15338 (N_15338,N_9627,N_2914);
and U15339 (N_15339,N_4143,N_4278);
and U15340 (N_15340,N_2428,N_769);
xnor U15341 (N_15341,N_365,N_1259);
or U15342 (N_15342,N_9516,N_4178);
and U15343 (N_15343,N_1337,N_7245);
xor U15344 (N_15344,N_7728,N_5318);
nand U15345 (N_15345,N_8543,N_1619);
xnor U15346 (N_15346,N_3119,N_6714);
nor U15347 (N_15347,N_4501,N_2670);
nand U15348 (N_15348,N_7341,N_9354);
xor U15349 (N_15349,N_7734,N_1215);
nand U15350 (N_15350,N_5109,N_6505);
and U15351 (N_15351,N_5743,N_7073);
or U15352 (N_15352,N_4347,N_931);
nor U15353 (N_15353,N_9461,N_9068);
and U15354 (N_15354,N_6571,N_4070);
nor U15355 (N_15355,N_1839,N_8450);
xnor U15356 (N_15356,N_2207,N_3366);
and U15357 (N_15357,N_3210,N_9109);
and U15358 (N_15358,N_2559,N_6792);
and U15359 (N_15359,N_1806,N_7421);
or U15360 (N_15360,N_7299,N_1340);
nand U15361 (N_15361,N_6894,N_2985);
xnor U15362 (N_15362,N_7282,N_639);
nand U15363 (N_15363,N_6268,N_987);
nand U15364 (N_15364,N_5029,N_7245);
nand U15365 (N_15365,N_8857,N_660);
and U15366 (N_15366,N_358,N_1916);
nor U15367 (N_15367,N_4578,N_6213);
nor U15368 (N_15368,N_5914,N_7784);
xnor U15369 (N_15369,N_4457,N_9175);
or U15370 (N_15370,N_3507,N_2227);
nand U15371 (N_15371,N_3399,N_1891);
xnor U15372 (N_15372,N_8594,N_5110);
nand U15373 (N_15373,N_219,N_1013);
nor U15374 (N_15374,N_2438,N_3520);
xnor U15375 (N_15375,N_4879,N_1812);
and U15376 (N_15376,N_6665,N_7335);
xor U15377 (N_15377,N_2109,N_5276);
or U15378 (N_15378,N_9440,N_1590);
or U15379 (N_15379,N_739,N_4215);
xnor U15380 (N_15380,N_6887,N_9871);
xor U15381 (N_15381,N_4290,N_7724);
nand U15382 (N_15382,N_2850,N_2110);
or U15383 (N_15383,N_951,N_5724);
nand U15384 (N_15384,N_5213,N_8796);
and U15385 (N_15385,N_4208,N_1502);
xor U15386 (N_15386,N_5648,N_1812);
or U15387 (N_15387,N_6933,N_3682);
nand U15388 (N_15388,N_2696,N_167);
or U15389 (N_15389,N_2046,N_7530);
or U15390 (N_15390,N_6029,N_2743);
xor U15391 (N_15391,N_6237,N_4563);
nand U15392 (N_15392,N_6352,N_5299);
and U15393 (N_15393,N_7775,N_459);
xnor U15394 (N_15394,N_2641,N_4082);
and U15395 (N_15395,N_8207,N_6430);
xor U15396 (N_15396,N_1401,N_5181);
or U15397 (N_15397,N_5382,N_9422);
or U15398 (N_15398,N_3953,N_7163);
and U15399 (N_15399,N_8226,N_4167);
xnor U15400 (N_15400,N_4513,N_2031);
nand U15401 (N_15401,N_9091,N_815);
xor U15402 (N_15402,N_80,N_887);
and U15403 (N_15403,N_4418,N_9014);
nor U15404 (N_15404,N_4030,N_3164);
nor U15405 (N_15405,N_2875,N_7574);
or U15406 (N_15406,N_1348,N_4801);
xnor U15407 (N_15407,N_5272,N_9536);
nand U15408 (N_15408,N_8532,N_4704);
or U15409 (N_15409,N_1037,N_4845);
or U15410 (N_15410,N_6153,N_3119);
and U15411 (N_15411,N_7578,N_3624);
nand U15412 (N_15412,N_2811,N_8216);
nor U15413 (N_15413,N_463,N_600);
and U15414 (N_15414,N_9824,N_49);
and U15415 (N_15415,N_7,N_4612);
or U15416 (N_15416,N_8766,N_6704);
nor U15417 (N_15417,N_6123,N_5304);
xor U15418 (N_15418,N_4429,N_7303);
or U15419 (N_15419,N_4235,N_1201);
nand U15420 (N_15420,N_5507,N_814);
xnor U15421 (N_15421,N_8198,N_5546);
nor U15422 (N_15422,N_4663,N_1048);
nor U15423 (N_15423,N_2238,N_5452);
and U15424 (N_15424,N_3473,N_835);
nand U15425 (N_15425,N_7020,N_9192);
nor U15426 (N_15426,N_8443,N_522);
nor U15427 (N_15427,N_185,N_8563);
nor U15428 (N_15428,N_8989,N_8518);
nor U15429 (N_15429,N_6564,N_8256);
nor U15430 (N_15430,N_2322,N_8497);
nand U15431 (N_15431,N_5951,N_8273);
xnor U15432 (N_15432,N_1082,N_4966);
or U15433 (N_15433,N_3194,N_1293);
and U15434 (N_15434,N_2219,N_674);
nor U15435 (N_15435,N_653,N_2075);
and U15436 (N_15436,N_8570,N_8441);
nor U15437 (N_15437,N_8123,N_2843);
xor U15438 (N_15438,N_4725,N_6149);
nor U15439 (N_15439,N_3909,N_4961);
or U15440 (N_15440,N_8573,N_4980);
and U15441 (N_15441,N_431,N_8088);
nand U15442 (N_15442,N_5063,N_9336);
or U15443 (N_15443,N_4878,N_7067);
and U15444 (N_15444,N_4352,N_8916);
and U15445 (N_15445,N_5431,N_4047);
xnor U15446 (N_15446,N_4586,N_4474);
and U15447 (N_15447,N_5026,N_3023);
nor U15448 (N_15448,N_9597,N_5041);
nand U15449 (N_15449,N_8099,N_2311);
or U15450 (N_15450,N_5594,N_3600);
or U15451 (N_15451,N_2956,N_987);
xnor U15452 (N_15452,N_9078,N_275);
xor U15453 (N_15453,N_2417,N_3475);
or U15454 (N_15454,N_2660,N_3043);
and U15455 (N_15455,N_5543,N_9819);
or U15456 (N_15456,N_1372,N_936);
nor U15457 (N_15457,N_4341,N_2417);
xor U15458 (N_15458,N_2567,N_9821);
and U15459 (N_15459,N_972,N_5715);
nor U15460 (N_15460,N_1309,N_8138);
and U15461 (N_15461,N_2098,N_4030);
nor U15462 (N_15462,N_6069,N_8147);
nor U15463 (N_15463,N_291,N_8064);
or U15464 (N_15464,N_6569,N_113);
nand U15465 (N_15465,N_9294,N_1148);
nor U15466 (N_15466,N_2149,N_8829);
xor U15467 (N_15467,N_5450,N_6072);
nand U15468 (N_15468,N_7104,N_3484);
and U15469 (N_15469,N_1133,N_8632);
nand U15470 (N_15470,N_5167,N_6238);
xor U15471 (N_15471,N_4363,N_437);
nand U15472 (N_15472,N_6682,N_4137);
nand U15473 (N_15473,N_991,N_1390);
nor U15474 (N_15474,N_5801,N_527);
xnor U15475 (N_15475,N_2756,N_726);
nor U15476 (N_15476,N_8581,N_5812);
or U15477 (N_15477,N_3941,N_8938);
nand U15478 (N_15478,N_5759,N_9678);
or U15479 (N_15479,N_3818,N_6372);
nor U15480 (N_15480,N_8120,N_9407);
nand U15481 (N_15481,N_6558,N_1493);
and U15482 (N_15482,N_8904,N_9734);
and U15483 (N_15483,N_4159,N_7940);
and U15484 (N_15484,N_3516,N_6395);
or U15485 (N_15485,N_532,N_2694);
and U15486 (N_15486,N_4887,N_7297);
nor U15487 (N_15487,N_7524,N_453);
nand U15488 (N_15488,N_2848,N_4841);
or U15489 (N_15489,N_620,N_7111);
nand U15490 (N_15490,N_691,N_1690);
xor U15491 (N_15491,N_7714,N_6497);
or U15492 (N_15492,N_2037,N_5636);
nor U15493 (N_15493,N_9417,N_81);
nand U15494 (N_15494,N_4594,N_678);
nand U15495 (N_15495,N_3785,N_2198);
nand U15496 (N_15496,N_5530,N_9702);
xor U15497 (N_15497,N_4856,N_3541);
and U15498 (N_15498,N_2569,N_1767);
xor U15499 (N_15499,N_1008,N_1383);
and U15500 (N_15500,N_4111,N_9053);
and U15501 (N_15501,N_9432,N_1917);
xnor U15502 (N_15502,N_2238,N_5594);
or U15503 (N_15503,N_5769,N_5968);
nor U15504 (N_15504,N_6698,N_738);
nand U15505 (N_15505,N_8842,N_7111);
and U15506 (N_15506,N_273,N_1584);
or U15507 (N_15507,N_4500,N_1875);
or U15508 (N_15508,N_89,N_1553);
nor U15509 (N_15509,N_6898,N_6533);
nor U15510 (N_15510,N_9485,N_4458);
and U15511 (N_15511,N_7001,N_6755);
or U15512 (N_15512,N_9996,N_4470);
and U15513 (N_15513,N_4124,N_3209);
or U15514 (N_15514,N_4568,N_5826);
nand U15515 (N_15515,N_4382,N_2561);
nand U15516 (N_15516,N_9890,N_7667);
xnor U15517 (N_15517,N_2405,N_8096);
nand U15518 (N_15518,N_6613,N_5417);
or U15519 (N_15519,N_6466,N_6873);
or U15520 (N_15520,N_9661,N_2299);
or U15521 (N_15521,N_6989,N_8633);
nand U15522 (N_15522,N_8798,N_6222);
nor U15523 (N_15523,N_6151,N_7438);
or U15524 (N_15524,N_9865,N_1811);
or U15525 (N_15525,N_8456,N_7702);
nor U15526 (N_15526,N_1949,N_8708);
nor U15527 (N_15527,N_2260,N_6115);
xnor U15528 (N_15528,N_7048,N_3917);
and U15529 (N_15529,N_4422,N_2417);
nand U15530 (N_15530,N_4747,N_2089);
xnor U15531 (N_15531,N_8039,N_9712);
xor U15532 (N_15532,N_2461,N_4483);
nor U15533 (N_15533,N_4052,N_9508);
nor U15534 (N_15534,N_3454,N_7618);
xor U15535 (N_15535,N_3493,N_8249);
nand U15536 (N_15536,N_1122,N_7986);
and U15537 (N_15537,N_4704,N_9790);
and U15538 (N_15538,N_7066,N_1435);
xor U15539 (N_15539,N_3856,N_920);
or U15540 (N_15540,N_2635,N_5897);
xor U15541 (N_15541,N_9589,N_7190);
xnor U15542 (N_15542,N_4377,N_8405);
xnor U15543 (N_15543,N_3141,N_2526);
nand U15544 (N_15544,N_5280,N_7372);
nor U15545 (N_15545,N_89,N_9161);
xor U15546 (N_15546,N_8972,N_3597);
xor U15547 (N_15547,N_8126,N_5736);
nor U15548 (N_15548,N_8501,N_714);
xor U15549 (N_15549,N_8329,N_7301);
nand U15550 (N_15550,N_1552,N_851);
xor U15551 (N_15551,N_5586,N_1098);
and U15552 (N_15552,N_6045,N_5446);
xnor U15553 (N_15553,N_5582,N_4476);
xor U15554 (N_15554,N_8627,N_3207);
nor U15555 (N_15555,N_2395,N_9127);
and U15556 (N_15556,N_5652,N_9243);
nor U15557 (N_15557,N_899,N_377);
or U15558 (N_15558,N_1823,N_5918);
xnor U15559 (N_15559,N_8400,N_9439);
or U15560 (N_15560,N_5261,N_9932);
xor U15561 (N_15561,N_1901,N_7340);
xnor U15562 (N_15562,N_5177,N_3387);
xor U15563 (N_15563,N_2560,N_3631);
nand U15564 (N_15564,N_7449,N_6147);
nor U15565 (N_15565,N_4584,N_5596);
nor U15566 (N_15566,N_4324,N_727);
xnor U15567 (N_15567,N_7323,N_5707);
and U15568 (N_15568,N_5482,N_4126);
xnor U15569 (N_15569,N_5237,N_7023);
xor U15570 (N_15570,N_3664,N_2555);
or U15571 (N_15571,N_4918,N_3931);
xor U15572 (N_15572,N_7535,N_7211);
or U15573 (N_15573,N_7843,N_2356);
or U15574 (N_15574,N_9670,N_4276);
and U15575 (N_15575,N_9774,N_85);
and U15576 (N_15576,N_5051,N_2142);
xor U15577 (N_15577,N_9397,N_203);
and U15578 (N_15578,N_5884,N_2103);
nor U15579 (N_15579,N_1880,N_9191);
nand U15580 (N_15580,N_2393,N_9632);
nor U15581 (N_15581,N_7302,N_9311);
and U15582 (N_15582,N_9172,N_6489);
xnor U15583 (N_15583,N_4044,N_198);
and U15584 (N_15584,N_4925,N_5969);
or U15585 (N_15585,N_3845,N_2848);
or U15586 (N_15586,N_5440,N_7367);
nor U15587 (N_15587,N_5315,N_4910);
nor U15588 (N_15588,N_9523,N_5110);
and U15589 (N_15589,N_6846,N_6527);
or U15590 (N_15590,N_6569,N_3315);
or U15591 (N_15591,N_5964,N_7929);
or U15592 (N_15592,N_6848,N_1269);
xnor U15593 (N_15593,N_62,N_4368);
nor U15594 (N_15594,N_6792,N_9480);
nor U15595 (N_15595,N_8996,N_9962);
xor U15596 (N_15596,N_7643,N_3084);
xnor U15597 (N_15597,N_8124,N_4668);
and U15598 (N_15598,N_4923,N_861);
or U15599 (N_15599,N_8299,N_1710);
nor U15600 (N_15600,N_5649,N_7118);
nand U15601 (N_15601,N_7766,N_7790);
or U15602 (N_15602,N_5768,N_9811);
nand U15603 (N_15603,N_7115,N_8606);
nor U15604 (N_15604,N_1239,N_6846);
xnor U15605 (N_15605,N_9258,N_2429);
and U15606 (N_15606,N_5670,N_6131);
nand U15607 (N_15607,N_320,N_2180);
nor U15608 (N_15608,N_4532,N_7611);
nand U15609 (N_15609,N_1788,N_7405);
or U15610 (N_15610,N_5227,N_7786);
xnor U15611 (N_15611,N_8501,N_7220);
or U15612 (N_15612,N_4029,N_3330);
and U15613 (N_15613,N_8109,N_3626);
or U15614 (N_15614,N_7386,N_5337);
or U15615 (N_15615,N_3159,N_7039);
xor U15616 (N_15616,N_6688,N_7011);
xnor U15617 (N_15617,N_3602,N_8849);
nand U15618 (N_15618,N_824,N_1061);
nand U15619 (N_15619,N_2662,N_9206);
xor U15620 (N_15620,N_4328,N_8177);
nor U15621 (N_15621,N_815,N_7425);
and U15622 (N_15622,N_9529,N_5587);
xor U15623 (N_15623,N_868,N_84);
and U15624 (N_15624,N_782,N_3938);
nand U15625 (N_15625,N_7599,N_5648);
and U15626 (N_15626,N_8071,N_5587);
nand U15627 (N_15627,N_2659,N_8857);
or U15628 (N_15628,N_9014,N_48);
nand U15629 (N_15629,N_8022,N_9261);
xor U15630 (N_15630,N_8595,N_8584);
nor U15631 (N_15631,N_9958,N_4837);
and U15632 (N_15632,N_4378,N_7386);
and U15633 (N_15633,N_8265,N_1225);
and U15634 (N_15634,N_7537,N_6405);
or U15635 (N_15635,N_1459,N_8366);
nand U15636 (N_15636,N_3796,N_7786);
xor U15637 (N_15637,N_765,N_2697);
and U15638 (N_15638,N_7804,N_8922);
nor U15639 (N_15639,N_3761,N_5280);
xor U15640 (N_15640,N_2894,N_4370);
nor U15641 (N_15641,N_2546,N_1102);
xnor U15642 (N_15642,N_4770,N_5893);
nor U15643 (N_15643,N_467,N_7312);
nor U15644 (N_15644,N_7103,N_3940);
nand U15645 (N_15645,N_7487,N_9214);
and U15646 (N_15646,N_5347,N_1041);
nand U15647 (N_15647,N_1459,N_4800);
nor U15648 (N_15648,N_949,N_676);
nor U15649 (N_15649,N_9398,N_3383);
nand U15650 (N_15650,N_5181,N_6311);
xnor U15651 (N_15651,N_1868,N_56);
or U15652 (N_15652,N_8664,N_2171);
and U15653 (N_15653,N_7760,N_260);
xnor U15654 (N_15654,N_5457,N_216);
nand U15655 (N_15655,N_7528,N_6457);
or U15656 (N_15656,N_6174,N_5732);
xor U15657 (N_15657,N_1404,N_8999);
nor U15658 (N_15658,N_8759,N_2620);
nor U15659 (N_15659,N_3348,N_5904);
nor U15660 (N_15660,N_5828,N_7755);
nand U15661 (N_15661,N_7877,N_7534);
nor U15662 (N_15662,N_3295,N_8904);
and U15663 (N_15663,N_525,N_8088);
nand U15664 (N_15664,N_8330,N_7740);
nor U15665 (N_15665,N_537,N_4096);
nand U15666 (N_15666,N_8955,N_7956);
or U15667 (N_15667,N_6612,N_5367);
or U15668 (N_15668,N_6990,N_1886);
nand U15669 (N_15669,N_5370,N_3294);
or U15670 (N_15670,N_9553,N_430);
or U15671 (N_15671,N_6388,N_2481);
xor U15672 (N_15672,N_7882,N_7384);
or U15673 (N_15673,N_6062,N_1493);
nor U15674 (N_15674,N_2665,N_8561);
nor U15675 (N_15675,N_2123,N_7961);
xnor U15676 (N_15676,N_7835,N_4632);
nand U15677 (N_15677,N_4343,N_1397);
or U15678 (N_15678,N_288,N_4270);
nand U15679 (N_15679,N_6837,N_1171);
or U15680 (N_15680,N_9522,N_9259);
or U15681 (N_15681,N_3952,N_8446);
nand U15682 (N_15682,N_5525,N_2688);
and U15683 (N_15683,N_1560,N_302);
nand U15684 (N_15684,N_8873,N_1975);
or U15685 (N_15685,N_1068,N_3012);
xnor U15686 (N_15686,N_4783,N_8141);
xnor U15687 (N_15687,N_5136,N_201);
or U15688 (N_15688,N_6128,N_9743);
nor U15689 (N_15689,N_641,N_5384);
and U15690 (N_15690,N_8734,N_4050);
xor U15691 (N_15691,N_1534,N_2133);
nor U15692 (N_15692,N_7376,N_7291);
or U15693 (N_15693,N_3584,N_9845);
or U15694 (N_15694,N_4497,N_6002);
or U15695 (N_15695,N_705,N_5743);
and U15696 (N_15696,N_5414,N_7751);
or U15697 (N_15697,N_4274,N_4527);
nand U15698 (N_15698,N_3171,N_9949);
nand U15699 (N_15699,N_7688,N_1817);
nor U15700 (N_15700,N_8209,N_4147);
nand U15701 (N_15701,N_8248,N_9580);
nand U15702 (N_15702,N_2108,N_2591);
xnor U15703 (N_15703,N_554,N_1141);
xnor U15704 (N_15704,N_2163,N_2860);
xor U15705 (N_15705,N_838,N_9440);
xnor U15706 (N_15706,N_1702,N_1245);
or U15707 (N_15707,N_4284,N_5694);
or U15708 (N_15708,N_6104,N_2341);
and U15709 (N_15709,N_3262,N_2742);
nand U15710 (N_15710,N_86,N_1073);
and U15711 (N_15711,N_8086,N_7377);
and U15712 (N_15712,N_4136,N_8960);
or U15713 (N_15713,N_4892,N_9020);
or U15714 (N_15714,N_7567,N_6193);
and U15715 (N_15715,N_2926,N_4588);
xor U15716 (N_15716,N_4426,N_8553);
and U15717 (N_15717,N_2313,N_8477);
nand U15718 (N_15718,N_3510,N_3740);
nand U15719 (N_15719,N_7093,N_1092);
and U15720 (N_15720,N_4550,N_1295);
xor U15721 (N_15721,N_9070,N_3675);
or U15722 (N_15722,N_3769,N_4996);
xor U15723 (N_15723,N_1854,N_3097);
or U15724 (N_15724,N_7927,N_6137);
and U15725 (N_15725,N_1471,N_3836);
nor U15726 (N_15726,N_3524,N_2995);
and U15727 (N_15727,N_5563,N_9097);
xor U15728 (N_15728,N_5409,N_1674);
or U15729 (N_15729,N_7295,N_9909);
or U15730 (N_15730,N_999,N_8585);
xnor U15731 (N_15731,N_2554,N_5013);
xnor U15732 (N_15732,N_4529,N_1549);
xor U15733 (N_15733,N_9496,N_2855);
xnor U15734 (N_15734,N_2305,N_8504);
and U15735 (N_15735,N_918,N_7817);
nand U15736 (N_15736,N_121,N_836);
or U15737 (N_15737,N_3895,N_9076);
nand U15738 (N_15738,N_3158,N_7216);
nand U15739 (N_15739,N_5921,N_6921);
and U15740 (N_15740,N_6119,N_8080);
or U15741 (N_15741,N_2590,N_578);
nand U15742 (N_15742,N_4677,N_7845);
nor U15743 (N_15743,N_3626,N_5638);
and U15744 (N_15744,N_3080,N_4720);
or U15745 (N_15745,N_2955,N_1102);
and U15746 (N_15746,N_2799,N_4230);
and U15747 (N_15747,N_260,N_7107);
nor U15748 (N_15748,N_7481,N_3261);
and U15749 (N_15749,N_2032,N_4454);
nor U15750 (N_15750,N_6069,N_6881);
and U15751 (N_15751,N_266,N_2855);
xor U15752 (N_15752,N_8914,N_7667);
or U15753 (N_15753,N_1137,N_2967);
nor U15754 (N_15754,N_5733,N_8067);
nand U15755 (N_15755,N_281,N_7669);
and U15756 (N_15756,N_2642,N_723);
xor U15757 (N_15757,N_7485,N_3074);
nand U15758 (N_15758,N_1404,N_4818);
or U15759 (N_15759,N_8117,N_1595);
or U15760 (N_15760,N_1583,N_7486);
or U15761 (N_15761,N_6737,N_9783);
nor U15762 (N_15762,N_1578,N_7452);
xor U15763 (N_15763,N_9504,N_424);
nor U15764 (N_15764,N_4306,N_8226);
nor U15765 (N_15765,N_436,N_6238);
xnor U15766 (N_15766,N_5673,N_4319);
and U15767 (N_15767,N_902,N_4516);
or U15768 (N_15768,N_7986,N_2569);
and U15769 (N_15769,N_7007,N_9362);
and U15770 (N_15770,N_2019,N_8806);
nand U15771 (N_15771,N_5637,N_8118);
nand U15772 (N_15772,N_9504,N_9076);
nor U15773 (N_15773,N_7127,N_2074);
and U15774 (N_15774,N_9565,N_6729);
nor U15775 (N_15775,N_3270,N_8331);
and U15776 (N_15776,N_5686,N_4122);
xor U15777 (N_15777,N_3114,N_3038);
or U15778 (N_15778,N_6051,N_4826);
xor U15779 (N_15779,N_2558,N_2842);
nand U15780 (N_15780,N_8966,N_1563);
and U15781 (N_15781,N_1567,N_2580);
or U15782 (N_15782,N_9503,N_2407);
nand U15783 (N_15783,N_9170,N_5944);
and U15784 (N_15784,N_1025,N_4624);
xnor U15785 (N_15785,N_5388,N_8387);
nand U15786 (N_15786,N_9218,N_3291);
nor U15787 (N_15787,N_7993,N_8571);
nand U15788 (N_15788,N_3673,N_4449);
or U15789 (N_15789,N_1070,N_6790);
nand U15790 (N_15790,N_7022,N_1473);
and U15791 (N_15791,N_170,N_747);
nor U15792 (N_15792,N_725,N_8567);
nand U15793 (N_15793,N_397,N_542);
or U15794 (N_15794,N_8375,N_8652);
nand U15795 (N_15795,N_7086,N_1151);
and U15796 (N_15796,N_7391,N_7871);
and U15797 (N_15797,N_9666,N_2111);
and U15798 (N_15798,N_7894,N_6358);
and U15799 (N_15799,N_3432,N_6989);
nand U15800 (N_15800,N_2655,N_6613);
nor U15801 (N_15801,N_2757,N_4892);
nand U15802 (N_15802,N_4212,N_4498);
nand U15803 (N_15803,N_3527,N_5348);
and U15804 (N_15804,N_3111,N_5529);
and U15805 (N_15805,N_401,N_5449);
and U15806 (N_15806,N_2404,N_7968);
and U15807 (N_15807,N_8567,N_8130);
xor U15808 (N_15808,N_2574,N_1467);
nand U15809 (N_15809,N_6313,N_9586);
xor U15810 (N_15810,N_693,N_2657);
or U15811 (N_15811,N_8808,N_6524);
and U15812 (N_15812,N_179,N_9320);
nand U15813 (N_15813,N_5270,N_9732);
nand U15814 (N_15814,N_7801,N_4324);
xnor U15815 (N_15815,N_1766,N_9645);
nor U15816 (N_15816,N_2429,N_3546);
and U15817 (N_15817,N_9559,N_127);
xnor U15818 (N_15818,N_9757,N_5428);
xor U15819 (N_15819,N_2388,N_1145);
and U15820 (N_15820,N_5500,N_5802);
and U15821 (N_15821,N_3963,N_1215);
nor U15822 (N_15822,N_9361,N_5790);
or U15823 (N_15823,N_6835,N_8552);
xor U15824 (N_15824,N_8163,N_5122);
or U15825 (N_15825,N_9606,N_6431);
and U15826 (N_15826,N_2730,N_6618);
or U15827 (N_15827,N_1286,N_810);
nor U15828 (N_15828,N_9753,N_4364);
nand U15829 (N_15829,N_3510,N_6645);
nor U15830 (N_15830,N_8762,N_5692);
nor U15831 (N_15831,N_2888,N_3259);
and U15832 (N_15832,N_9754,N_2179);
xnor U15833 (N_15833,N_3093,N_2860);
nor U15834 (N_15834,N_6863,N_7444);
and U15835 (N_15835,N_2675,N_6112);
and U15836 (N_15836,N_7594,N_3433);
or U15837 (N_15837,N_4121,N_7574);
nand U15838 (N_15838,N_8134,N_6903);
or U15839 (N_15839,N_8284,N_2412);
nand U15840 (N_15840,N_4882,N_541);
and U15841 (N_15841,N_9434,N_7055);
nand U15842 (N_15842,N_7664,N_3791);
nor U15843 (N_15843,N_8031,N_368);
xor U15844 (N_15844,N_5797,N_6104);
nand U15845 (N_15845,N_9034,N_1247);
or U15846 (N_15846,N_5531,N_3716);
and U15847 (N_15847,N_3621,N_464);
nor U15848 (N_15848,N_5502,N_1340);
and U15849 (N_15849,N_8981,N_5859);
nand U15850 (N_15850,N_4975,N_9145);
nor U15851 (N_15851,N_7695,N_2556);
xor U15852 (N_15852,N_8136,N_8204);
or U15853 (N_15853,N_4247,N_7219);
nand U15854 (N_15854,N_3598,N_5868);
xnor U15855 (N_15855,N_3313,N_4723);
or U15856 (N_15856,N_5907,N_9129);
and U15857 (N_15857,N_6766,N_5932);
nand U15858 (N_15858,N_2390,N_3048);
nand U15859 (N_15859,N_7434,N_1009);
nor U15860 (N_15860,N_2193,N_846);
nor U15861 (N_15861,N_859,N_5334);
xnor U15862 (N_15862,N_3682,N_8757);
or U15863 (N_15863,N_3454,N_3376);
nor U15864 (N_15864,N_2382,N_8683);
and U15865 (N_15865,N_2610,N_1991);
nor U15866 (N_15866,N_7431,N_5485);
nand U15867 (N_15867,N_9471,N_5531);
and U15868 (N_15868,N_4428,N_8658);
and U15869 (N_15869,N_2040,N_3836);
and U15870 (N_15870,N_280,N_1118);
or U15871 (N_15871,N_9240,N_9868);
nor U15872 (N_15872,N_4287,N_5909);
nor U15873 (N_15873,N_1517,N_7964);
nor U15874 (N_15874,N_7060,N_8986);
or U15875 (N_15875,N_8126,N_3815);
nor U15876 (N_15876,N_6218,N_3896);
and U15877 (N_15877,N_1198,N_9875);
and U15878 (N_15878,N_9384,N_6539);
nor U15879 (N_15879,N_8530,N_6216);
and U15880 (N_15880,N_301,N_1621);
and U15881 (N_15881,N_2893,N_2658);
nor U15882 (N_15882,N_7619,N_6222);
nor U15883 (N_15883,N_1572,N_4006);
and U15884 (N_15884,N_4099,N_6520);
and U15885 (N_15885,N_1542,N_9600);
nand U15886 (N_15886,N_710,N_54);
and U15887 (N_15887,N_658,N_5559);
xor U15888 (N_15888,N_2415,N_1819);
and U15889 (N_15889,N_5122,N_8816);
xor U15890 (N_15890,N_8475,N_3196);
and U15891 (N_15891,N_8071,N_7313);
nand U15892 (N_15892,N_4281,N_1002);
and U15893 (N_15893,N_2362,N_7639);
nor U15894 (N_15894,N_4904,N_5600);
or U15895 (N_15895,N_4785,N_6851);
xnor U15896 (N_15896,N_2877,N_7967);
and U15897 (N_15897,N_4524,N_6190);
or U15898 (N_15898,N_6424,N_2178);
nor U15899 (N_15899,N_9620,N_1281);
or U15900 (N_15900,N_94,N_1279);
or U15901 (N_15901,N_7797,N_5230);
nand U15902 (N_15902,N_6630,N_9060);
nor U15903 (N_15903,N_1814,N_1076);
or U15904 (N_15904,N_6191,N_6497);
nand U15905 (N_15905,N_7487,N_8500);
or U15906 (N_15906,N_4142,N_8012);
nand U15907 (N_15907,N_8824,N_4054);
xor U15908 (N_15908,N_1341,N_8020);
nand U15909 (N_15909,N_5844,N_4617);
nor U15910 (N_15910,N_2181,N_8571);
xnor U15911 (N_15911,N_7569,N_3878);
nand U15912 (N_15912,N_1307,N_5460);
nand U15913 (N_15913,N_1194,N_5498);
xor U15914 (N_15914,N_210,N_9979);
nand U15915 (N_15915,N_5937,N_4044);
and U15916 (N_15916,N_2228,N_3839);
or U15917 (N_15917,N_7085,N_1186);
xor U15918 (N_15918,N_1798,N_4686);
nor U15919 (N_15919,N_4902,N_5639);
and U15920 (N_15920,N_1633,N_2920);
nand U15921 (N_15921,N_4127,N_9049);
xnor U15922 (N_15922,N_5882,N_1748);
xor U15923 (N_15923,N_3978,N_1753);
and U15924 (N_15924,N_2612,N_8634);
xnor U15925 (N_15925,N_9836,N_1848);
nor U15926 (N_15926,N_1678,N_8523);
or U15927 (N_15927,N_708,N_890);
and U15928 (N_15928,N_5057,N_9914);
xnor U15929 (N_15929,N_5902,N_9717);
and U15930 (N_15930,N_7213,N_5780);
nor U15931 (N_15931,N_5361,N_6426);
and U15932 (N_15932,N_2947,N_8610);
or U15933 (N_15933,N_6443,N_4599);
nand U15934 (N_15934,N_3059,N_3168);
nor U15935 (N_15935,N_5083,N_4918);
or U15936 (N_15936,N_8088,N_6460);
xnor U15937 (N_15937,N_1388,N_7271);
nor U15938 (N_15938,N_4997,N_7450);
and U15939 (N_15939,N_2343,N_1467);
nand U15940 (N_15940,N_8898,N_870);
nand U15941 (N_15941,N_96,N_39);
or U15942 (N_15942,N_9120,N_6088);
and U15943 (N_15943,N_7912,N_9220);
and U15944 (N_15944,N_8765,N_3645);
xor U15945 (N_15945,N_9790,N_5773);
or U15946 (N_15946,N_9563,N_2949);
xor U15947 (N_15947,N_6344,N_5876);
nor U15948 (N_15948,N_1270,N_3777);
or U15949 (N_15949,N_4881,N_3695);
xnor U15950 (N_15950,N_3516,N_404);
nand U15951 (N_15951,N_5031,N_2733);
nand U15952 (N_15952,N_6548,N_9267);
and U15953 (N_15953,N_528,N_3911);
xnor U15954 (N_15954,N_6213,N_8893);
nor U15955 (N_15955,N_4104,N_7155);
and U15956 (N_15956,N_6716,N_9766);
or U15957 (N_15957,N_8056,N_6357);
nand U15958 (N_15958,N_2285,N_5306);
xnor U15959 (N_15959,N_1190,N_6466);
nor U15960 (N_15960,N_2407,N_5087);
xor U15961 (N_15961,N_1211,N_4526);
xor U15962 (N_15962,N_5684,N_2394);
nor U15963 (N_15963,N_9546,N_7866);
or U15964 (N_15964,N_1158,N_2716);
xnor U15965 (N_15965,N_8556,N_860);
nand U15966 (N_15966,N_6605,N_3258);
nand U15967 (N_15967,N_184,N_1033);
or U15968 (N_15968,N_2020,N_265);
nor U15969 (N_15969,N_7451,N_7912);
nor U15970 (N_15970,N_3020,N_4497);
and U15971 (N_15971,N_7043,N_7479);
and U15972 (N_15972,N_3940,N_5496);
xor U15973 (N_15973,N_6668,N_9865);
nand U15974 (N_15974,N_27,N_8010);
and U15975 (N_15975,N_8930,N_6132);
and U15976 (N_15976,N_1548,N_1107);
nand U15977 (N_15977,N_1387,N_4937);
or U15978 (N_15978,N_2762,N_7695);
nor U15979 (N_15979,N_7020,N_3671);
and U15980 (N_15980,N_9779,N_9055);
and U15981 (N_15981,N_3222,N_5799);
nand U15982 (N_15982,N_639,N_526);
nor U15983 (N_15983,N_7759,N_2501);
nand U15984 (N_15984,N_4395,N_2660);
nor U15985 (N_15985,N_4314,N_5277);
xnor U15986 (N_15986,N_9008,N_9355);
or U15987 (N_15987,N_8516,N_1665);
and U15988 (N_15988,N_5533,N_4563);
xnor U15989 (N_15989,N_8208,N_3017);
and U15990 (N_15990,N_612,N_2245);
xor U15991 (N_15991,N_1490,N_9769);
and U15992 (N_15992,N_9069,N_9777);
nand U15993 (N_15993,N_6613,N_2968);
nand U15994 (N_15994,N_3112,N_1454);
and U15995 (N_15995,N_1496,N_4569);
nand U15996 (N_15996,N_6939,N_2471);
xnor U15997 (N_15997,N_8032,N_2497);
nand U15998 (N_15998,N_9449,N_6479);
or U15999 (N_15999,N_2971,N_2541);
or U16000 (N_16000,N_9127,N_1564);
nor U16001 (N_16001,N_612,N_4997);
nand U16002 (N_16002,N_4870,N_9962);
or U16003 (N_16003,N_9731,N_339);
nor U16004 (N_16004,N_9080,N_4277);
nand U16005 (N_16005,N_3697,N_412);
nand U16006 (N_16006,N_2490,N_8538);
or U16007 (N_16007,N_333,N_3547);
or U16008 (N_16008,N_182,N_1737);
and U16009 (N_16009,N_8691,N_936);
nand U16010 (N_16010,N_6555,N_8009);
nor U16011 (N_16011,N_1828,N_1613);
and U16012 (N_16012,N_1449,N_4363);
or U16013 (N_16013,N_5062,N_823);
and U16014 (N_16014,N_5650,N_8999);
xnor U16015 (N_16015,N_7914,N_4641);
and U16016 (N_16016,N_5314,N_6344);
or U16017 (N_16017,N_3562,N_5229);
nor U16018 (N_16018,N_3081,N_3986);
xor U16019 (N_16019,N_8586,N_3444);
and U16020 (N_16020,N_4157,N_5622);
nand U16021 (N_16021,N_5979,N_2877);
xnor U16022 (N_16022,N_2773,N_688);
nor U16023 (N_16023,N_4929,N_4281);
nor U16024 (N_16024,N_9577,N_7441);
nand U16025 (N_16025,N_897,N_3885);
and U16026 (N_16026,N_8152,N_8408);
and U16027 (N_16027,N_6234,N_9278);
or U16028 (N_16028,N_9921,N_9648);
xnor U16029 (N_16029,N_3809,N_9136);
or U16030 (N_16030,N_4066,N_5111);
xor U16031 (N_16031,N_5847,N_7510);
or U16032 (N_16032,N_2131,N_2073);
nand U16033 (N_16033,N_398,N_7458);
or U16034 (N_16034,N_9812,N_8775);
or U16035 (N_16035,N_5516,N_484);
xnor U16036 (N_16036,N_806,N_2850);
and U16037 (N_16037,N_3079,N_379);
nand U16038 (N_16038,N_334,N_6367);
nand U16039 (N_16039,N_2212,N_1853);
or U16040 (N_16040,N_9841,N_3672);
nor U16041 (N_16041,N_9688,N_9560);
xor U16042 (N_16042,N_952,N_286);
and U16043 (N_16043,N_8996,N_1784);
or U16044 (N_16044,N_1815,N_3169);
and U16045 (N_16045,N_650,N_9371);
and U16046 (N_16046,N_1569,N_238);
or U16047 (N_16047,N_7732,N_3064);
and U16048 (N_16048,N_4215,N_5469);
nor U16049 (N_16049,N_9978,N_9866);
nand U16050 (N_16050,N_387,N_1688);
or U16051 (N_16051,N_6196,N_6165);
or U16052 (N_16052,N_7778,N_6438);
and U16053 (N_16053,N_9815,N_51);
xnor U16054 (N_16054,N_4866,N_3540);
xnor U16055 (N_16055,N_5006,N_2488);
xnor U16056 (N_16056,N_1636,N_1735);
or U16057 (N_16057,N_7162,N_8273);
nand U16058 (N_16058,N_3652,N_8614);
nor U16059 (N_16059,N_2447,N_9231);
and U16060 (N_16060,N_5300,N_6960);
nand U16061 (N_16061,N_555,N_6868);
nand U16062 (N_16062,N_6968,N_9896);
or U16063 (N_16063,N_6362,N_8911);
or U16064 (N_16064,N_6728,N_5580);
nand U16065 (N_16065,N_3742,N_9089);
xor U16066 (N_16066,N_7897,N_5233);
and U16067 (N_16067,N_2090,N_6606);
nand U16068 (N_16068,N_9531,N_3066);
nand U16069 (N_16069,N_3690,N_8783);
and U16070 (N_16070,N_5429,N_4945);
or U16071 (N_16071,N_5278,N_9106);
xnor U16072 (N_16072,N_9460,N_3782);
or U16073 (N_16073,N_6502,N_1664);
nand U16074 (N_16074,N_94,N_3030);
xnor U16075 (N_16075,N_8950,N_7843);
nor U16076 (N_16076,N_2030,N_4145);
or U16077 (N_16077,N_8343,N_2368);
xnor U16078 (N_16078,N_8417,N_1386);
xor U16079 (N_16079,N_4545,N_1469);
nand U16080 (N_16080,N_7392,N_9729);
nor U16081 (N_16081,N_6340,N_6102);
or U16082 (N_16082,N_2310,N_9294);
and U16083 (N_16083,N_815,N_9423);
xnor U16084 (N_16084,N_3668,N_492);
and U16085 (N_16085,N_4558,N_8791);
nor U16086 (N_16086,N_145,N_5005);
and U16087 (N_16087,N_483,N_6179);
or U16088 (N_16088,N_13,N_3180);
nand U16089 (N_16089,N_3977,N_2531);
or U16090 (N_16090,N_1730,N_9867);
nor U16091 (N_16091,N_189,N_8524);
nand U16092 (N_16092,N_8290,N_2598);
nand U16093 (N_16093,N_5982,N_7602);
and U16094 (N_16094,N_5622,N_2480);
nor U16095 (N_16095,N_6220,N_4956);
xnor U16096 (N_16096,N_5828,N_4620);
nand U16097 (N_16097,N_176,N_6468);
or U16098 (N_16098,N_194,N_9128);
and U16099 (N_16099,N_9963,N_117);
xor U16100 (N_16100,N_198,N_2063);
xor U16101 (N_16101,N_1895,N_7269);
and U16102 (N_16102,N_5368,N_9559);
and U16103 (N_16103,N_8458,N_6222);
nor U16104 (N_16104,N_7668,N_7716);
and U16105 (N_16105,N_1269,N_1526);
xnor U16106 (N_16106,N_8200,N_5728);
or U16107 (N_16107,N_8048,N_9934);
xor U16108 (N_16108,N_8614,N_9682);
xor U16109 (N_16109,N_2835,N_4735);
xor U16110 (N_16110,N_20,N_1640);
xor U16111 (N_16111,N_240,N_7499);
xnor U16112 (N_16112,N_6800,N_5180);
and U16113 (N_16113,N_8519,N_4387);
nand U16114 (N_16114,N_9221,N_4390);
nor U16115 (N_16115,N_7652,N_3769);
and U16116 (N_16116,N_7146,N_7160);
xnor U16117 (N_16117,N_8502,N_2921);
or U16118 (N_16118,N_7011,N_9731);
or U16119 (N_16119,N_3565,N_2929);
nor U16120 (N_16120,N_9623,N_4754);
nand U16121 (N_16121,N_9806,N_5195);
or U16122 (N_16122,N_7603,N_8116);
nand U16123 (N_16123,N_7470,N_1429);
and U16124 (N_16124,N_6658,N_3977);
or U16125 (N_16125,N_2531,N_5731);
nand U16126 (N_16126,N_2301,N_8641);
xnor U16127 (N_16127,N_6344,N_6420);
nand U16128 (N_16128,N_6357,N_2538);
nor U16129 (N_16129,N_9412,N_4296);
nand U16130 (N_16130,N_365,N_8530);
nor U16131 (N_16131,N_5484,N_7282);
xor U16132 (N_16132,N_9260,N_5931);
xor U16133 (N_16133,N_3435,N_5246);
nor U16134 (N_16134,N_5231,N_8737);
or U16135 (N_16135,N_1159,N_1974);
nor U16136 (N_16136,N_3860,N_1799);
and U16137 (N_16137,N_2373,N_7226);
or U16138 (N_16138,N_593,N_7904);
nor U16139 (N_16139,N_7824,N_5384);
xnor U16140 (N_16140,N_9918,N_3409);
or U16141 (N_16141,N_4611,N_2181);
nor U16142 (N_16142,N_1885,N_5715);
and U16143 (N_16143,N_4806,N_4122);
or U16144 (N_16144,N_8475,N_5842);
and U16145 (N_16145,N_6266,N_6996);
nand U16146 (N_16146,N_2860,N_2323);
nand U16147 (N_16147,N_1399,N_1509);
or U16148 (N_16148,N_8744,N_9243);
nand U16149 (N_16149,N_4321,N_1256);
nor U16150 (N_16150,N_1406,N_7928);
xor U16151 (N_16151,N_7029,N_3276);
xor U16152 (N_16152,N_7002,N_1372);
and U16153 (N_16153,N_1980,N_7428);
nor U16154 (N_16154,N_4231,N_2694);
and U16155 (N_16155,N_2083,N_942);
nand U16156 (N_16156,N_6651,N_9626);
nand U16157 (N_16157,N_6834,N_2363);
xor U16158 (N_16158,N_4335,N_8946);
xor U16159 (N_16159,N_8071,N_3988);
and U16160 (N_16160,N_423,N_9585);
xor U16161 (N_16161,N_9468,N_2420);
or U16162 (N_16162,N_7696,N_5575);
or U16163 (N_16163,N_9086,N_5996);
or U16164 (N_16164,N_7465,N_8212);
or U16165 (N_16165,N_5716,N_4119);
or U16166 (N_16166,N_8275,N_3560);
xor U16167 (N_16167,N_6249,N_9439);
nor U16168 (N_16168,N_2573,N_2670);
or U16169 (N_16169,N_7831,N_561);
or U16170 (N_16170,N_8339,N_3394);
and U16171 (N_16171,N_7269,N_747);
and U16172 (N_16172,N_391,N_5911);
or U16173 (N_16173,N_5786,N_2640);
nor U16174 (N_16174,N_9557,N_5585);
nor U16175 (N_16175,N_2841,N_3871);
nor U16176 (N_16176,N_2239,N_3723);
nor U16177 (N_16177,N_4432,N_8260);
or U16178 (N_16178,N_5360,N_3054);
nand U16179 (N_16179,N_5138,N_481);
or U16180 (N_16180,N_9491,N_1552);
or U16181 (N_16181,N_5542,N_6466);
xnor U16182 (N_16182,N_6186,N_7251);
and U16183 (N_16183,N_3616,N_9826);
xnor U16184 (N_16184,N_1635,N_7244);
or U16185 (N_16185,N_8498,N_1211);
and U16186 (N_16186,N_9827,N_7644);
xnor U16187 (N_16187,N_4870,N_6950);
nand U16188 (N_16188,N_6818,N_758);
nand U16189 (N_16189,N_1440,N_2231);
xor U16190 (N_16190,N_805,N_499);
nor U16191 (N_16191,N_5920,N_3758);
nor U16192 (N_16192,N_4601,N_2208);
xnor U16193 (N_16193,N_5289,N_7013);
nor U16194 (N_16194,N_923,N_5520);
xnor U16195 (N_16195,N_5596,N_8937);
xor U16196 (N_16196,N_4703,N_9240);
or U16197 (N_16197,N_8030,N_6345);
or U16198 (N_16198,N_5787,N_5784);
xnor U16199 (N_16199,N_1319,N_3286);
nor U16200 (N_16200,N_5876,N_6792);
or U16201 (N_16201,N_3743,N_1414);
xor U16202 (N_16202,N_4531,N_2053);
nor U16203 (N_16203,N_9041,N_2081);
nor U16204 (N_16204,N_1248,N_6284);
and U16205 (N_16205,N_2042,N_831);
nand U16206 (N_16206,N_3243,N_9665);
xnor U16207 (N_16207,N_5056,N_8444);
nor U16208 (N_16208,N_6148,N_8705);
xor U16209 (N_16209,N_6502,N_4720);
xor U16210 (N_16210,N_1588,N_8779);
nor U16211 (N_16211,N_9915,N_6405);
nor U16212 (N_16212,N_547,N_17);
and U16213 (N_16213,N_816,N_1595);
nand U16214 (N_16214,N_8771,N_3713);
and U16215 (N_16215,N_5239,N_1476);
or U16216 (N_16216,N_1634,N_1580);
nand U16217 (N_16217,N_3870,N_8924);
nand U16218 (N_16218,N_1663,N_2509);
and U16219 (N_16219,N_8927,N_762);
nor U16220 (N_16220,N_5593,N_2236);
nor U16221 (N_16221,N_6207,N_5428);
nand U16222 (N_16222,N_484,N_5949);
and U16223 (N_16223,N_8673,N_1797);
xnor U16224 (N_16224,N_1071,N_8234);
nand U16225 (N_16225,N_6450,N_8844);
nand U16226 (N_16226,N_7,N_4144);
xor U16227 (N_16227,N_1547,N_5174);
and U16228 (N_16228,N_7171,N_1700);
or U16229 (N_16229,N_848,N_3424);
xnor U16230 (N_16230,N_6157,N_2736);
and U16231 (N_16231,N_591,N_3294);
or U16232 (N_16232,N_3181,N_6426);
xnor U16233 (N_16233,N_3960,N_1216);
nand U16234 (N_16234,N_4431,N_6304);
nor U16235 (N_16235,N_4089,N_4522);
or U16236 (N_16236,N_9289,N_866);
nand U16237 (N_16237,N_4125,N_4118);
xor U16238 (N_16238,N_8043,N_998);
nor U16239 (N_16239,N_4220,N_6133);
xor U16240 (N_16240,N_9146,N_5802);
nand U16241 (N_16241,N_2326,N_6686);
nand U16242 (N_16242,N_8324,N_8091);
or U16243 (N_16243,N_2049,N_7603);
nand U16244 (N_16244,N_3270,N_7499);
or U16245 (N_16245,N_6779,N_1543);
or U16246 (N_16246,N_8142,N_4531);
nand U16247 (N_16247,N_9302,N_5265);
nor U16248 (N_16248,N_2411,N_3247);
nand U16249 (N_16249,N_6662,N_4513);
nor U16250 (N_16250,N_2627,N_6116);
xor U16251 (N_16251,N_5203,N_7065);
and U16252 (N_16252,N_2932,N_7290);
xnor U16253 (N_16253,N_2155,N_1881);
nor U16254 (N_16254,N_4788,N_6465);
nand U16255 (N_16255,N_99,N_7547);
and U16256 (N_16256,N_9799,N_3385);
nand U16257 (N_16257,N_3468,N_3788);
nor U16258 (N_16258,N_6826,N_2920);
xnor U16259 (N_16259,N_1109,N_8344);
nor U16260 (N_16260,N_4357,N_7687);
and U16261 (N_16261,N_5293,N_1397);
and U16262 (N_16262,N_6040,N_9171);
and U16263 (N_16263,N_2799,N_2326);
and U16264 (N_16264,N_1846,N_8604);
nor U16265 (N_16265,N_5178,N_7604);
or U16266 (N_16266,N_6293,N_7993);
or U16267 (N_16267,N_5167,N_8393);
or U16268 (N_16268,N_7568,N_7456);
and U16269 (N_16269,N_390,N_3049);
or U16270 (N_16270,N_9716,N_6853);
and U16271 (N_16271,N_1627,N_2867);
nor U16272 (N_16272,N_9773,N_8560);
or U16273 (N_16273,N_7499,N_8480);
and U16274 (N_16274,N_8754,N_1179);
or U16275 (N_16275,N_9047,N_7411);
nand U16276 (N_16276,N_1213,N_4911);
and U16277 (N_16277,N_5814,N_6832);
and U16278 (N_16278,N_3816,N_6335);
and U16279 (N_16279,N_3854,N_6461);
xor U16280 (N_16280,N_4064,N_936);
and U16281 (N_16281,N_3394,N_2579);
and U16282 (N_16282,N_6348,N_842);
or U16283 (N_16283,N_9277,N_7190);
and U16284 (N_16284,N_3729,N_8137);
or U16285 (N_16285,N_5682,N_5318);
nor U16286 (N_16286,N_1542,N_9603);
nor U16287 (N_16287,N_5203,N_5915);
or U16288 (N_16288,N_6804,N_7136);
nand U16289 (N_16289,N_8510,N_279);
xnor U16290 (N_16290,N_5080,N_8738);
nand U16291 (N_16291,N_4322,N_2590);
xor U16292 (N_16292,N_4525,N_4838);
nor U16293 (N_16293,N_4257,N_8061);
xnor U16294 (N_16294,N_57,N_1308);
nand U16295 (N_16295,N_4871,N_4004);
and U16296 (N_16296,N_5117,N_8398);
xnor U16297 (N_16297,N_9209,N_5958);
and U16298 (N_16298,N_4174,N_1640);
or U16299 (N_16299,N_6998,N_1137);
xor U16300 (N_16300,N_3136,N_4332);
and U16301 (N_16301,N_6771,N_7561);
or U16302 (N_16302,N_5031,N_3017);
xor U16303 (N_16303,N_9712,N_8503);
nor U16304 (N_16304,N_7244,N_5570);
nand U16305 (N_16305,N_5465,N_8892);
nand U16306 (N_16306,N_6490,N_6902);
or U16307 (N_16307,N_666,N_701);
nor U16308 (N_16308,N_9447,N_6872);
or U16309 (N_16309,N_7877,N_7012);
nor U16310 (N_16310,N_1047,N_7100);
nand U16311 (N_16311,N_5957,N_6056);
nor U16312 (N_16312,N_1819,N_4358);
xor U16313 (N_16313,N_6955,N_4533);
or U16314 (N_16314,N_7420,N_1288);
nand U16315 (N_16315,N_7339,N_362);
nor U16316 (N_16316,N_3481,N_1892);
xnor U16317 (N_16317,N_5453,N_8251);
nor U16318 (N_16318,N_5006,N_8562);
xor U16319 (N_16319,N_9759,N_764);
nand U16320 (N_16320,N_7261,N_1948);
xnor U16321 (N_16321,N_226,N_6069);
and U16322 (N_16322,N_7510,N_2343);
or U16323 (N_16323,N_454,N_6648);
nor U16324 (N_16324,N_4079,N_1412);
nand U16325 (N_16325,N_687,N_4782);
and U16326 (N_16326,N_6717,N_9644);
or U16327 (N_16327,N_9943,N_7799);
nor U16328 (N_16328,N_6859,N_9280);
nor U16329 (N_16329,N_6067,N_4334);
nand U16330 (N_16330,N_8202,N_6079);
nor U16331 (N_16331,N_8105,N_8541);
or U16332 (N_16332,N_5047,N_8748);
xor U16333 (N_16333,N_4787,N_5837);
xor U16334 (N_16334,N_7286,N_4754);
nand U16335 (N_16335,N_4922,N_9663);
xnor U16336 (N_16336,N_3324,N_1918);
nor U16337 (N_16337,N_3307,N_4727);
nand U16338 (N_16338,N_3155,N_1575);
or U16339 (N_16339,N_8256,N_3005);
nand U16340 (N_16340,N_2828,N_6762);
or U16341 (N_16341,N_733,N_5521);
or U16342 (N_16342,N_8551,N_1793);
or U16343 (N_16343,N_2149,N_2594);
or U16344 (N_16344,N_4932,N_8420);
nand U16345 (N_16345,N_940,N_3341);
and U16346 (N_16346,N_5051,N_2076);
nor U16347 (N_16347,N_3270,N_5483);
nand U16348 (N_16348,N_2933,N_4166);
and U16349 (N_16349,N_153,N_891);
nor U16350 (N_16350,N_8423,N_7188);
or U16351 (N_16351,N_5325,N_9907);
or U16352 (N_16352,N_2686,N_5674);
and U16353 (N_16353,N_2751,N_5194);
xor U16354 (N_16354,N_4325,N_9467);
and U16355 (N_16355,N_999,N_1618);
or U16356 (N_16356,N_7132,N_4805);
nor U16357 (N_16357,N_6645,N_8030);
or U16358 (N_16358,N_7956,N_6339);
and U16359 (N_16359,N_1053,N_3056);
nand U16360 (N_16360,N_7030,N_4940);
nand U16361 (N_16361,N_6956,N_7313);
nand U16362 (N_16362,N_3102,N_2408);
nor U16363 (N_16363,N_535,N_5468);
nand U16364 (N_16364,N_9436,N_8931);
or U16365 (N_16365,N_5682,N_5576);
or U16366 (N_16366,N_4848,N_7342);
xor U16367 (N_16367,N_6434,N_5434);
nand U16368 (N_16368,N_877,N_2707);
nor U16369 (N_16369,N_4524,N_8738);
nand U16370 (N_16370,N_7190,N_4934);
xnor U16371 (N_16371,N_1170,N_2609);
and U16372 (N_16372,N_4897,N_4106);
and U16373 (N_16373,N_3471,N_9911);
and U16374 (N_16374,N_8153,N_9026);
xor U16375 (N_16375,N_2226,N_3327);
nor U16376 (N_16376,N_3226,N_202);
or U16377 (N_16377,N_8787,N_3974);
nor U16378 (N_16378,N_4848,N_4639);
or U16379 (N_16379,N_9548,N_5501);
nor U16380 (N_16380,N_4639,N_9677);
xnor U16381 (N_16381,N_3016,N_6654);
and U16382 (N_16382,N_3952,N_6119);
xor U16383 (N_16383,N_4806,N_5169);
xor U16384 (N_16384,N_7049,N_108);
nand U16385 (N_16385,N_5094,N_854);
nor U16386 (N_16386,N_6381,N_5338);
and U16387 (N_16387,N_3281,N_8755);
or U16388 (N_16388,N_9163,N_3446);
or U16389 (N_16389,N_8952,N_7628);
nor U16390 (N_16390,N_7812,N_9522);
nand U16391 (N_16391,N_6794,N_3015);
xor U16392 (N_16392,N_4511,N_3028);
xor U16393 (N_16393,N_5035,N_1407);
xnor U16394 (N_16394,N_3170,N_8715);
nor U16395 (N_16395,N_697,N_5161);
or U16396 (N_16396,N_8731,N_8700);
xnor U16397 (N_16397,N_1860,N_9862);
xor U16398 (N_16398,N_8453,N_7761);
and U16399 (N_16399,N_5513,N_9387);
nor U16400 (N_16400,N_5237,N_8760);
xor U16401 (N_16401,N_8962,N_7639);
and U16402 (N_16402,N_3156,N_9382);
nor U16403 (N_16403,N_7095,N_3840);
nand U16404 (N_16404,N_7105,N_8924);
or U16405 (N_16405,N_2247,N_8817);
xor U16406 (N_16406,N_2922,N_9729);
xor U16407 (N_16407,N_2657,N_9394);
nand U16408 (N_16408,N_5669,N_7588);
and U16409 (N_16409,N_3401,N_8537);
nor U16410 (N_16410,N_5885,N_8300);
xor U16411 (N_16411,N_3846,N_2087);
xor U16412 (N_16412,N_1588,N_4441);
xor U16413 (N_16413,N_2112,N_3666);
nor U16414 (N_16414,N_9019,N_3209);
nand U16415 (N_16415,N_622,N_8458);
nand U16416 (N_16416,N_8289,N_4100);
or U16417 (N_16417,N_4633,N_4048);
nor U16418 (N_16418,N_3625,N_8721);
or U16419 (N_16419,N_9850,N_274);
or U16420 (N_16420,N_8626,N_868);
xnor U16421 (N_16421,N_719,N_8215);
xor U16422 (N_16422,N_8642,N_8246);
or U16423 (N_16423,N_9062,N_6263);
nand U16424 (N_16424,N_6581,N_4007);
nand U16425 (N_16425,N_181,N_5466);
nand U16426 (N_16426,N_5342,N_1231);
or U16427 (N_16427,N_8014,N_6704);
and U16428 (N_16428,N_9765,N_3712);
xor U16429 (N_16429,N_5032,N_8081);
or U16430 (N_16430,N_5389,N_7297);
nand U16431 (N_16431,N_3112,N_5667);
nand U16432 (N_16432,N_6345,N_8721);
and U16433 (N_16433,N_7869,N_6478);
or U16434 (N_16434,N_7501,N_7286);
nand U16435 (N_16435,N_9667,N_7336);
or U16436 (N_16436,N_2856,N_1871);
nand U16437 (N_16437,N_788,N_1681);
nand U16438 (N_16438,N_3742,N_1401);
and U16439 (N_16439,N_3459,N_8058);
nand U16440 (N_16440,N_4391,N_5841);
or U16441 (N_16441,N_1651,N_1819);
xnor U16442 (N_16442,N_4217,N_5050);
nor U16443 (N_16443,N_5361,N_2716);
xnor U16444 (N_16444,N_3732,N_1492);
nor U16445 (N_16445,N_6765,N_2960);
nor U16446 (N_16446,N_5764,N_7475);
nand U16447 (N_16447,N_5644,N_4744);
nor U16448 (N_16448,N_6892,N_5432);
xor U16449 (N_16449,N_6662,N_7532);
nand U16450 (N_16450,N_8153,N_7706);
xor U16451 (N_16451,N_1724,N_1735);
nand U16452 (N_16452,N_1708,N_885);
nand U16453 (N_16453,N_5815,N_1130);
and U16454 (N_16454,N_6256,N_6163);
or U16455 (N_16455,N_7680,N_347);
nor U16456 (N_16456,N_4519,N_3905);
nand U16457 (N_16457,N_3426,N_3702);
nor U16458 (N_16458,N_7804,N_4909);
or U16459 (N_16459,N_7595,N_2529);
xor U16460 (N_16460,N_2064,N_7735);
nor U16461 (N_16461,N_2701,N_6415);
nand U16462 (N_16462,N_6676,N_7910);
nor U16463 (N_16463,N_5707,N_1449);
and U16464 (N_16464,N_8791,N_1119);
and U16465 (N_16465,N_3226,N_7369);
nand U16466 (N_16466,N_2129,N_2877);
nor U16467 (N_16467,N_9858,N_3676);
and U16468 (N_16468,N_9173,N_150);
nor U16469 (N_16469,N_7326,N_60);
nor U16470 (N_16470,N_9973,N_5730);
nor U16471 (N_16471,N_9898,N_3277);
xnor U16472 (N_16472,N_6657,N_3443);
xor U16473 (N_16473,N_5276,N_2552);
xor U16474 (N_16474,N_6276,N_1781);
xnor U16475 (N_16475,N_6796,N_8385);
or U16476 (N_16476,N_9268,N_5511);
and U16477 (N_16477,N_5786,N_6975);
nor U16478 (N_16478,N_7046,N_9407);
nand U16479 (N_16479,N_2992,N_5479);
nor U16480 (N_16480,N_2997,N_5611);
nand U16481 (N_16481,N_5327,N_8271);
nor U16482 (N_16482,N_9250,N_698);
nand U16483 (N_16483,N_893,N_8612);
and U16484 (N_16484,N_1118,N_2898);
nor U16485 (N_16485,N_2718,N_1932);
xnor U16486 (N_16486,N_519,N_8680);
nor U16487 (N_16487,N_508,N_9014);
nand U16488 (N_16488,N_1923,N_3519);
xnor U16489 (N_16489,N_4014,N_819);
and U16490 (N_16490,N_5482,N_6918);
nor U16491 (N_16491,N_5935,N_3321);
nand U16492 (N_16492,N_1168,N_583);
and U16493 (N_16493,N_553,N_4014);
nand U16494 (N_16494,N_9801,N_2996);
or U16495 (N_16495,N_1592,N_9417);
and U16496 (N_16496,N_211,N_2733);
or U16497 (N_16497,N_7621,N_6539);
and U16498 (N_16498,N_8791,N_7723);
or U16499 (N_16499,N_9013,N_5729);
xnor U16500 (N_16500,N_346,N_9728);
xnor U16501 (N_16501,N_1149,N_6849);
and U16502 (N_16502,N_4575,N_124);
xor U16503 (N_16503,N_9917,N_5669);
nor U16504 (N_16504,N_7295,N_8931);
nand U16505 (N_16505,N_6861,N_24);
nor U16506 (N_16506,N_199,N_9463);
nand U16507 (N_16507,N_9641,N_1413);
nor U16508 (N_16508,N_5455,N_7581);
xor U16509 (N_16509,N_8082,N_2353);
nor U16510 (N_16510,N_5541,N_2944);
xnor U16511 (N_16511,N_6840,N_711);
nor U16512 (N_16512,N_8808,N_9733);
and U16513 (N_16513,N_8307,N_3781);
nor U16514 (N_16514,N_9378,N_6082);
nor U16515 (N_16515,N_7711,N_78);
nor U16516 (N_16516,N_5257,N_3226);
nor U16517 (N_16517,N_7711,N_7544);
xnor U16518 (N_16518,N_3819,N_3787);
xnor U16519 (N_16519,N_4932,N_314);
nor U16520 (N_16520,N_7539,N_5052);
xnor U16521 (N_16521,N_3189,N_1921);
nand U16522 (N_16522,N_7810,N_2919);
and U16523 (N_16523,N_6087,N_5364);
and U16524 (N_16524,N_4203,N_3462);
or U16525 (N_16525,N_9310,N_8445);
xnor U16526 (N_16526,N_5567,N_5615);
nor U16527 (N_16527,N_6989,N_9383);
or U16528 (N_16528,N_2970,N_6339);
nand U16529 (N_16529,N_4238,N_934);
nor U16530 (N_16530,N_623,N_5428);
xnor U16531 (N_16531,N_894,N_5264);
nand U16532 (N_16532,N_3684,N_5336);
xnor U16533 (N_16533,N_7264,N_2453);
xnor U16534 (N_16534,N_1598,N_8518);
nor U16535 (N_16535,N_7124,N_7085);
and U16536 (N_16536,N_5648,N_9965);
nand U16537 (N_16537,N_3465,N_6810);
nand U16538 (N_16538,N_1821,N_5392);
xor U16539 (N_16539,N_4209,N_9057);
or U16540 (N_16540,N_2288,N_7079);
and U16541 (N_16541,N_97,N_1895);
xnor U16542 (N_16542,N_1583,N_7796);
and U16543 (N_16543,N_5077,N_2907);
nand U16544 (N_16544,N_8255,N_1276);
and U16545 (N_16545,N_1115,N_6611);
xnor U16546 (N_16546,N_4019,N_5169);
nand U16547 (N_16547,N_1944,N_886);
nand U16548 (N_16548,N_9495,N_4769);
nand U16549 (N_16549,N_7421,N_1626);
nor U16550 (N_16550,N_7153,N_5125);
or U16551 (N_16551,N_194,N_2950);
nand U16552 (N_16552,N_7594,N_9108);
or U16553 (N_16553,N_2613,N_2219);
nand U16554 (N_16554,N_990,N_5472);
or U16555 (N_16555,N_2613,N_6155);
or U16556 (N_16556,N_9333,N_3203);
nand U16557 (N_16557,N_5314,N_100);
xor U16558 (N_16558,N_3752,N_2800);
nand U16559 (N_16559,N_5291,N_6483);
nand U16560 (N_16560,N_9139,N_4901);
or U16561 (N_16561,N_9432,N_5095);
and U16562 (N_16562,N_5355,N_3167);
and U16563 (N_16563,N_452,N_9254);
nor U16564 (N_16564,N_1293,N_2986);
or U16565 (N_16565,N_6484,N_1129);
nand U16566 (N_16566,N_28,N_2467);
nand U16567 (N_16567,N_3844,N_9834);
nor U16568 (N_16568,N_3589,N_7112);
nand U16569 (N_16569,N_6625,N_670);
or U16570 (N_16570,N_2035,N_1831);
nor U16571 (N_16571,N_407,N_2704);
or U16572 (N_16572,N_1447,N_6670);
nand U16573 (N_16573,N_7303,N_6396);
nor U16574 (N_16574,N_9233,N_820);
and U16575 (N_16575,N_9949,N_7889);
nor U16576 (N_16576,N_4063,N_2112);
or U16577 (N_16577,N_4631,N_8367);
and U16578 (N_16578,N_6628,N_1007);
nor U16579 (N_16579,N_6351,N_6960);
nand U16580 (N_16580,N_4901,N_4382);
xor U16581 (N_16581,N_1138,N_5755);
and U16582 (N_16582,N_2845,N_7);
or U16583 (N_16583,N_5515,N_2885);
nand U16584 (N_16584,N_6501,N_9999);
nor U16585 (N_16585,N_6614,N_4330);
and U16586 (N_16586,N_1788,N_7033);
xnor U16587 (N_16587,N_1589,N_3442);
nor U16588 (N_16588,N_814,N_7555);
nand U16589 (N_16589,N_1046,N_5698);
and U16590 (N_16590,N_5582,N_885);
or U16591 (N_16591,N_4296,N_8767);
or U16592 (N_16592,N_4718,N_6496);
nor U16593 (N_16593,N_2783,N_3793);
nor U16594 (N_16594,N_1253,N_9463);
nand U16595 (N_16595,N_7919,N_523);
and U16596 (N_16596,N_5664,N_7318);
nand U16597 (N_16597,N_2440,N_7795);
or U16598 (N_16598,N_6730,N_7542);
or U16599 (N_16599,N_6772,N_3976);
xnor U16600 (N_16600,N_4293,N_8422);
or U16601 (N_16601,N_1682,N_5657);
xnor U16602 (N_16602,N_5472,N_1147);
and U16603 (N_16603,N_3387,N_8691);
xnor U16604 (N_16604,N_502,N_5413);
or U16605 (N_16605,N_9252,N_2856);
nor U16606 (N_16606,N_7124,N_3739);
nand U16607 (N_16607,N_6518,N_3773);
xor U16608 (N_16608,N_573,N_5651);
nand U16609 (N_16609,N_4117,N_7340);
nor U16610 (N_16610,N_288,N_6662);
and U16611 (N_16611,N_7455,N_7745);
xnor U16612 (N_16612,N_7072,N_8165);
or U16613 (N_16613,N_3050,N_4317);
nand U16614 (N_16614,N_8881,N_7370);
xnor U16615 (N_16615,N_3911,N_1020);
nand U16616 (N_16616,N_5745,N_8624);
xnor U16617 (N_16617,N_5460,N_7028);
or U16618 (N_16618,N_8426,N_4146);
nor U16619 (N_16619,N_9320,N_2799);
xor U16620 (N_16620,N_9651,N_1113);
nor U16621 (N_16621,N_8281,N_8176);
and U16622 (N_16622,N_9231,N_2320);
xor U16623 (N_16623,N_9189,N_8787);
and U16624 (N_16624,N_6967,N_8396);
nor U16625 (N_16625,N_1835,N_3482);
nor U16626 (N_16626,N_5334,N_662);
nor U16627 (N_16627,N_646,N_3431);
xnor U16628 (N_16628,N_3397,N_63);
nand U16629 (N_16629,N_541,N_3615);
nand U16630 (N_16630,N_4511,N_7212);
and U16631 (N_16631,N_6914,N_4027);
or U16632 (N_16632,N_7322,N_2517);
xor U16633 (N_16633,N_5266,N_3528);
xor U16634 (N_16634,N_4507,N_3171);
nor U16635 (N_16635,N_1529,N_9015);
nand U16636 (N_16636,N_2762,N_2201);
or U16637 (N_16637,N_4515,N_3501);
nand U16638 (N_16638,N_4390,N_7757);
and U16639 (N_16639,N_8444,N_4443);
nand U16640 (N_16640,N_6452,N_3576);
and U16641 (N_16641,N_5289,N_2412);
nor U16642 (N_16642,N_6402,N_8271);
nor U16643 (N_16643,N_2908,N_5079);
or U16644 (N_16644,N_7494,N_906);
and U16645 (N_16645,N_7492,N_9702);
nand U16646 (N_16646,N_8694,N_637);
and U16647 (N_16647,N_8066,N_7907);
and U16648 (N_16648,N_3392,N_2160);
and U16649 (N_16649,N_6517,N_2812);
nand U16650 (N_16650,N_3024,N_8257);
nand U16651 (N_16651,N_3141,N_2978);
or U16652 (N_16652,N_6625,N_4126);
nand U16653 (N_16653,N_1553,N_1387);
xnor U16654 (N_16654,N_1930,N_1234);
and U16655 (N_16655,N_6259,N_9857);
nor U16656 (N_16656,N_1311,N_1812);
and U16657 (N_16657,N_7526,N_843);
or U16658 (N_16658,N_9879,N_612);
and U16659 (N_16659,N_9120,N_7928);
or U16660 (N_16660,N_3445,N_1009);
or U16661 (N_16661,N_1192,N_8998);
or U16662 (N_16662,N_7838,N_1135);
nand U16663 (N_16663,N_4802,N_61);
nand U16664 (N_16664,N_7965,N_2011);
or U16665 (N_16665,N_6578,N_3797);
and U16666 (N_16666,N_4252,N_9469);
nor U16667 (N_16667,N_4282,N_4622);
and U16668 (N_16668,N_2939,N_8172);
xor U16669 (N_16669,N_7353,N_9972);
or U16670 (N_16670,N_126,N_5876);
or U16671 (N_16671,N_4476,N_2255);
or U16672 (N_16672,N_4525,N_8365);
and U16673 (N_16673,N_6891,N_1875);
nand U16674 (N_16674,N_5658,N_6612);
nor U16675 (N_16675,N_4030,N_116);
or U16676 (N_16676,N_2124,N_3277);
nor U16677 (N_16677,N_1923,N_1447);
and U16678 (N_16678,N_1594,N_3411);
and U16679 (N_16679,N_1400,N_7446);
and U16680 (N_16680,N_8417,N_9292);
and U16681 (N_16681,N_8827,N_4581);
and U16682 (N_16682,N_1229,N_1500);
nand U16683 (N_16683,N_4600,N_5641);
or U16684 (N_16684,N_5929,N_9230);
and U16685 (N_16685,N_113,N_6957);
nor U16686 (N_16686,N_1308,N_9787);
xnor U16687 (N_16687,N_4568,N_7675);
nand U16688 (N_16688,N_4911,N_8472);
or U16689 (N_16689,N_8787,N_8204);
nand U16690 (N_16690,N_5734,N_8931);
and U16691 (N_16691,N_2753,N_2484);
and U16692 (N_16692,N_1682,N_1916);
nor U16693 (N_16693,N_8654,N_6109);
xor U16694 (N_16694,N_3837,N_9236);
nand U16695 (N_16695,N_7838,N_8890);
or U16696 (N_16696,N_7922,N_8592);
or U16697 (N_16697,N_1914,N_2924);
xnor U16698 (N_16698,N_3749,N_1862);
xor U16699 (N_16699,N_6526,N_298);
nor U16700 (N_16700,N_1780,N_2936);
xnor U16701 (N_16701,N_860,N_7591);
nand U16702 (N_16702,N_3406,N_6970);
nor U16703 (N_16703,N_5985,N_7759);
nor U16704 (N_16704,N_9138,N_8749);
and U16705 (N_16705,N_2202,N_1855);
nand U16706 (N_16706,N_919,N_3220);
nor U16707 (N_16707,N_2142,N_726);
or U16708 (N_16708,N_2967,N_6996);
xor U16709 (N_16709,N_6867,N_39);
or U16710 (N_16710,N_1364,N_4994);
or U16711 (N_16711,N_722,N_3178);
and U16712 (N_16712,N_9125,N_3311);
nand U16713 (N_16713,N_1284,N_1749);
or U16714 (N_16714,N_3936,N_4021);
nand U16715 (N_16715,N_8571,N_8396);
nand U16716 (N_16716,N_7563,N_457);
nand U16717 (N_16717,N_3621,N_9837);
or U16718 (N_16718,N_9050,N_259);
and U16719 (N_16719,N_1614,N_1003);
nor U16720 (N_16720,N_3729,N_5430);
xor U16721 (N_16721,N_5415,N_6457);
or U16722 (N_16722,N_4104,N_3543);
nand U16723 (N_16723,N_5055,N_2354);
nand U16724 (N_16724,N_4830,N_9352);
or U16725 (N_16725,N_1869,N_9938);
and U16726 (N_16726,N_4616,N_1993);
and U16727 (N_16727,N_111,N_6561);
nor U16728 (N_16728,N_5742,N_5333);
or U16729 (N_16729,N_8936,N_7458);
xor U16730 (N_16730,N_9698,N_2730);
and U16731 (N_16731,N_8470,N_6793);
xnor U16732 (N_16732,N_5736,N_1557);
xor U16733 (N_16733,N_4381,N_9957);
xor U16734 (N_16734,N_7635,N_3987);
and U16735 (N_16735,N_3926,N_9956);
nand U16736 (N_16736,N_1664,N_1613);
or U16737 (N_16737,N_6506,N_3009);
nor U16738 (N_16738,N_9268,N_5195);
nand U16739 (N_16739,N_7337,N_2383);
nor U16740 (N_16740,N_1405,N_7913);
nor U16741 (N_16741,N_352,N_9738);
and U16742 (N_16742,N_1130,N_3671);
or U16743 (N_16743,N_9642,N_5598);
and U16744 (N_16744,N_3357,N_1677);
and U16745 (N_16745,N_7681,N_7628);
or U16746 (N_16746,N_9655,N_8499);
and U16747 (N_16747,N_5848,N_6860);
xor U16748 (N_16748,N_9427,N_6530);
xnor U16749 (N_16749,N_7161,N_5247);
nor U16750 (N_16750,N_1613,N_5917);
and U16751 (N_16751,N_2481,N_2452);
nor U16752 (N_16752,N_5385,N_4687);
nand U16753 (N_16753,N_2295,N_5213);
or U16754 (N_16754,N_8585,N_3385);
xnor U16755 (N_16755,N_4495,N_4812);
and U16756 (N_16756,N_3477,N_1232);
or U16757 (N_16757,N_3465,N_9799);
xor U16758 (N_16758,N_2130,N_8302);
nor U16759 (N_16759,N_1402,N_8628);
xnor U16760 (N_16760,N_8478,N_8632);
and U16761 (N_16761,N_2924,N_464);
or U16762 (N_16762,N_2549,N_3862);
nand U16763 (N_16763,N_8331,N_574);
or U16764 (N_16764,N_7977,N_6806);
nand U16765 (N_16765,N_3326,N_2467);
xor U16766 (N_16766,N_3363,N_9677);
nand U16767 (N_16767,N_7376,N_2011);
nand U16768 (N_16768,N_3531,N_1228);
xor U16769 (N_16769,N_8272,N_3686);
nor U16770 (N_16770,N_1654,N_7101);
nor U16771 (N_16771,N_3172,N_6785);
and U16772 (N_16772,N_4328,N_7342);
or U16773 (N_16773,N_2858,N_9839);
nand U16774 (N_16774,N_9114,N_7404);
or U16775 (N_16775,N_9823,N_8728);
or U16776 (N_16776,N_6480,N_4415);
nor U16777 (N_16777,N_6752,N_7272);
nand U16778 (N_16778,N_6467,N_6432);
nor U16779 (N_16779,N_1361,N_5912);
nor U16780 (N_16780,N_5880,N_9587);
nand U16781 (N_16781,N_9733,N_1491);
xor U16782 (N_16782,N_8285,N_5324);
or U16783 (N_16783,N_3798,N_5191);
nor U16784 (N_16784,N_4136,N_8467);
nand U16785 (N_16785,N_8633,N_6446);
and U16786 (N_16786,N_9912,N_8560);
nor U16787 (N_16787,N_2803,N_8764);
xnor U16788 (N_16788,N_8357,N_1148);
nand U16789 (N_16789,N_255,N_2729);
or U16790 (N_16790,N_8712,N_810);
and U16791 (N_16791,N_7498,N_3663);
and U16792 (N_16792,N_5732,N_5232);
nand U16793 (N_16793,N_6169,N_7255);
and U16794 (N_16794,N_4904,N_125);
xnor U16795 (N_16795,N_7264,N_1315);
or U16796 (N_16796,N_2830,N_2086);
and U16797 (N_16797,N_9826,N_659);
nor U16798 (N_16798,N_9747,N_4148);
or U16799 (N_16799,N_7018,N_8232);
nand U16800 (N_16800,N_717,N_9591);
nand U16801 (N_16801,N_4008,N_1146);
nor U16802 (N_16802,N_2341,N_6525);
nor U16803 (N_16803,N_9831,N_7844);
xor U16804 (N_16804,N_1859,N_3281);
nand U16805 (N_16805,N_449,N_9452);
xnor U16806 (N_16806,N_6254,N_5409);
nor U16807 (N_16807,N_9758,N_6415);
xor U16808 (N_16808,N_4916,N_1744);
or U16809 (N_16809,N_6315,N_7059);
xnor U16810 (N_16810,N_2056,N_913);
nor U16811 (N_16811,N_1633,N_4428);
and U16812 (N_16812,N_9524,N_9112);
and U16813 (N_16813,N_7451,N_3269);
nor U16814 (N_16814,N_257,N_3216);
xor U16815 (N_16815,N_8906,N_3582);
and U16816 (N_16816,N_4884,N_1922);
nand U16817 (N_16817,N_2908,N_9400);
or U16818 (N_16818,N_3758,N_597);
or U16819 (N_16819,N_5612,N_9445);
xor U16820 (N_16820,N_6913,N_642);
or U16821 (N_16821,N_3578,N_6921);
nand U16822 (N_16822,N_2674,N_1542);
xnor U16823 (N_16823,N_7245,N_4007);
nand U16824 (N_16824,N_805,N_7420);
and U16825 (N_16825,N_1854,N_1410);
or U16826 (N_16826,N_9988,N_2826);
and U16827 (N_16827,N_582,N_4745);
nor U16828 (N_16828,N_9491,N_947);
nand U16829 (N_16829,N_824,N_795);
nand U16830 (N_16830,N_4672,N_9728);
or U16831 (N_16831,N_6658,N_6657);
xnor U16832 (N_16832,N_734,N_6174);
xor U16833 (N_16833,N_3107,N_2421);
or U16834 (N_16834,N_416,N_3762);
nor U16835 (N_16835,N_1940,N_2620);
nor U16836 (N_16836,N_5365,N_3566);
and U16837 (N_16837,N_2596,N_4707);
xor U16838 (N_16838,N_3406,N_7630);
or U16839 (N_16839,N_9621,N_8084);
nor U16840 (N_16840,N_2766,N_4071);
and U16841 (N_16841,N_87,N_4332);
xor U16842 (N_16842,N_2863,N_9755);
xnor U16843 (N_16843,N_5967,N_2900);
nand U16844 (N_16844,N_3946,N_1582);
xor U16845 (N_16845,N_7448,N_6338);
or U16846 (N_16846,N_4788,N_7378);
and U16847 (N_16847,N_555,N_1892);
and U16848 (N_16848,N_6063,N_5264);
nand U16849 (N_16849,N_1440,N_6788);
and U16850 (N_16850,N_563,N_6029);
nand U16851 (N_16851,N_1406,N_2053);
xnor U16852 (N_16852,N_5832,N_8980);
nand U16853 (N_16853,N_4295,N_8804);
and U16854 (N_16854,N_6899,N_6827);
nor U16855 (N_16855,N_8486,N_5667);
nor U16856 (N_16856,N_8009,N_8076);
xnor U16857 (N_16857,N_6192,N_3238);
and U16858 (N_16858,N_841,N_9437);
or U16859 (N_16859,N_8756,N_5677);
nand U16860 (N_16860,N_8920,N_1928);
or U16861 (N_16861,N_547,N_1978);
nand U16862 (N_16862,N_6126,N_5576);
and U16863 (N_16863,N_1563,N_1821);
or U16864 (N_16864,N_2622,N_9243);
and U16865 (N_16865,N_4655,N_2428);
or U16866 (N_16866,N_9211,N_1503);
nor U16867 (N_16867,N_8566,N_3016);
nand U16868 (N_16868,N_3636,N_9490);
nor U16869 (N_16869,N_3252,N_3103);
or U16870 (N_16870,N_3240,N_3873);
nand U16871 (N_16871,N_5212,N_3181);
or U16872 (N_16872,N_3998,N_886);
and U16873 (N_16873,N_8915,N_406);
xnor U16874 (N_16874,N_5304,N_5658);
xnor U16875 (N_16875,N_6894,N_3042);
and U16876 (N_16876,N_6160,N_9732);
or U16877 (N_16877,N_1742,N_3538);
xnor U16878 (N_16878,N_3811,N_9446);
nor U16879 (N_16879,N_2706,N_907);
or U16880 (N_16880,N_4196,N_5052);
nor U16881 (N_16881,N_8713,N_6024);
and U16882 (N_16882,N_9961,N_8282);
xor U16883 (N_16883,N_3697,N_4346);
and U16884 (N_16884,N_5986,N_2411);
nor U16885 (N_16885,N_4209,N_7183);
or U16886 (N_16886,N_3823,N_8321);
nand U16887 (N_16887,N_1832,N_7186);
nand U16888 (N_16888,N_2725,N_6090);
xor U16889 (N_16889,N_5259,N_6080);
and U16890 (N_16890,N_705,N_901);
nand U16891 (N_16891,N_2045,N_550);
or U16892 (N_16892,N_3668,N_106);
xor U16893 (N_16893,N_426,N_8262);
xor U16894 (N_16894,N_8390,N_6241);
or U16895 (N_16895,N_3632,N_241);
xor U16896 (N_16896,N_2254,N_5875);
nand U16897 (N_16897,N_9007,N_2022);
or U16898 (N_16898,N_8971,N_7357);
or U16899 (N_16899,N_792,N_2689);
nor U16900 (N_16900,N_8471,N_1215);
nand U16901 (N_16901,N_4886,N_7852);
nand U16902 (N_16902,N_4288,N_5600);
nor U16903 (N_16903,N_7835,N_6615);
and U16904 (N_16904,N_9049,N_2780);
or U16905 (N_16905,N_694,N_4670);
or U16906 (N_16906,N_5418,N_5125);
or U16907 (N_16907,N_2474,N_2817);
nand U16908 (N_16908,N_2449,N_1015);
nand U16909 (N_16909,N_7741,N_1720);
and U16910 (N_16910,N_3795,N_2221);
and U16911 (N_16911,N_484,N_7563);
and U16912 (N_16912,N_2880,N_7843);
or U16913 (N_16913,N_6922,N_2461);
or U16914 (N_16914,N_4730,N_7374);
nor U16915 (N_16915,N_7474,N_4028);
and U16916 (N_16916,N_7669,N_4229);
nor U16917 (N_16917,N_8917,N_5921);
nor U16918 (N_16918,N_9519,N_6581);
nor U16919 (N_16919,N_1514,N_7748);
or U16920 (N_16920,N_8414,N_9408);
nor U16921 (N_16921,N_9223,N_5380);
or U16922 (N_16922,N_3114,N_9357);
and U16923 (N_16923,N_4491,N_9688);
xnor U16924 (N_16924,N_8775,N_8432);
xor U16925 (N_16925,N_2649,N_9487);
or U16926 (N_16926,N_3078,N_6571);
or U16927 (N_16927,N_5600,N_4328);
xnor U16928 (N_16928,N_116,N_8870);
nor U16929 (N_16929,N_429,N_9249);
xor U16930 (N_16930,N_684,N_9269);
or U16931 (N_16931,N_3384,N_6746);
xnor U16932 (N_16932,N_8121,N_413);
xor U16933 (N_16933,N_388,N_4929);
nand U16934 (N_16934,N_5763,N_3018);
nand U16935 (N_16935,N_1801,N_641);
or U16936 (N_16936,N_3633,N_2035);
and U16937 (N_16937,N_7553,N_1454);
and U16938 (N_16938,N_995,N_3218);
nor U16939 (N_16939,N_7960,N_4014);
nand U16940 (N_16940,N_9414,N_6899);
nor U16941 (N_16941,N_4299,N_5665);
nand U16942 (N_16942,N_1523,N_2050);
nor U16943 (N_16943,N_5530,N_1456);
or U16944 (N_16944,N_6408,N_3257);
nor U16945 (N_16945,N_8556,N_8899);
nor U16946 (N_16946,N_7307,N_6916);
nor U16947 (N_16947,N_6472,N_2833);
and U16948 (N_16948,N_9773,N_7897);
nor U16949 (N_16949,N_1108,N_7757);
xnor U16950 (N_16950,N_7261,N_5867);
or U16951 (N_16951,N_1112,N_6426);
xor U16952 (N_16952,N_5542,N_4785);
xor U16953 (N_16953,N_6031,N_1295);
nand U16954 (N_16954,N_4139,N_9597);
nor U16955 (N_16955,N_86,N_6020);
xnor U16956 (N_16956,N_7808,N_2007);
or U16957 (N_16957,N_3926,N_143);
nor U16958 (N_16958,N_6090,N_7589);
xnor U16959 (N_16959,N_6584,N_344);
xor U16960 (N_16960,N_1200,N_2746);
xnor U16961 (N_16961,N_5169,N_9231);
xor U16962 (N_16962,N_418,N_590);
or U16963 (N_16963,N_4738,N_8159);
or U16964 (N_16964,N_8540,N_1386);
xor U16965 (N_16965,N_1041,N_5989);
nor U16966 (N_16966,N_6387,N_3973);
and U16967 (N_16967,N_8386,N_7379);
xor U16968 (N_16968,N_6717,N_3092);
nand U16969 (N_16969,N_5141,N_8434);
xnor U16970 (N_16970,N_7866,N_288);
or U16971 (N_16971,N_9940,N_3020);
or U16972 (N_16972,N_3231,N_9276);
nand U16973 (N_16973,N_8223,N_6115);
or U16974 (N_16974,N_5840,N_5015);
and U16975 (N_16975,N_608,N_1228);
nor U16976 (N_16976,N_1747,N_9115);
and U16977 (N_16977,N_6223,N_1843);
nor U16978 (N_16978,N_7578,N_5907);
nor U16979 (N_16979,N_545,N_3855);
nor U16980 (N_16980,N_2890,N_9252);
and U16981 (N_16981,N_499,N_527);
nand U16982 (N_16982,N_7518,N_6804);
xor U16983 (N_16983,N_6656,N_2047);
and U16984 (N_16984,N_1716,N_3069);
nor U16985 (N_16985,N_2484,N_8865);
nand U16986 (N_16986,N_3433,N_1110);
and U16987 (N_16987,N_465,N_8968);
or U16988 (N_16988,N_8962,N_2373);
and U16989 (N_16989,N_69,N_2020);
nor U16990 (N_16990,N_8613,N_4293);
nand U16991 (N_16991,N_9156,N_8172);
and U16992 (N_16992,N_3002,N_3783);
xor U16993 (N_16993,N_83,N_9068);
nor U16994 (N_16994,N_6747,N_231);
and U16995 (N_16995,N_2323,N_7044);
or U16996 (N_16996,N_996,N_470);
xnor U16997 (N_16997,N_956,N_2705);
xnor U16998 (N_16998,N_2921,N_9586);
and U16999 (N_16999,N_161,N_4108);
nand U17000 (N_17000,N_1348,N_9802);
and U17001 (N_17001,N_1434,N_8418);
xnor U17002 (N_17002,N_5244,N_8917);
nor U17003 (N_17003,N_9580,N_5268);
and U17004 (N_17004,N_8666,N_2796);
or U17005 (N_17005,N_3371,N_1318);
or U17006 (N_17006,N_8857,N_7747);
xor U17007 (N_17007,N_5189,N_7464);
and U17008 (N_17008,N_5305,N_6469);
or U17009 (N_17009,N_995,N_7278);
or U17010 (N_17010,N_5455,N_6930);
or U17011 (N_17011,N_345,N_6734);
or U17012 (N_17012,N_8400,N_6885);
nor U17013 (N_17013,N_4892,N_2006);
xor U17014 (N_17014,N_9214,N_9857);
nor U17015 (N_17015,N_2156,N_1601);
and U17016 (N_17016,N_1782,N_6297);
nand U17017 (N_17017,N_3826,N_7163);
and U17018 (N_17018,N_762,N_2567);
nand U17019 (N_17019,N_837,N_8281);
xnor U17020 (N_17020,N_443,N_4751);
and U17021 (N_17021,N_5367,N_1308);
nor U17022 (N_17022,N_3238,N_1771);
or U17023 (N_17023,N_1202,N_972);
or U17024 (N_17024,N_8447,N_7726);
or U17025 (N_17025,N_4560,N_8806);
or U17026 (N_17026,N_3079,N_3793);
and U17027 (N_17027,N_6306,N_9414);
nor U17028 (N_17028,N_8068,N_1184);
nand U17029 (N_17029,N_3871,N_4488);
or U17030 (N_17030,N_9742,N_7998);
xnor U17031 (N_17031,N_6362,N_1602);
or U17032 (N_17032,N_3104,N_6906);
xor U17033 (N_17033,N_9531,N_4919);
nand U17034 (N_17034,N_2724,N_5510);
and U17035 (N_17035,N_1061,N_4211);
xor U17036 (N_17036,N_7648,N_4360);
nand U17037 (N_17037,N_9329,N_7451);
and U17038 (N_17038,N_2955,N_2212);
or U17039 (N_17039,N_1056,N_4674);
nor U17040 (N_17040,N_5461,N_2397);
or U17041 (N_17041,N_2278,N_630);
or U17042 (N_17042,N_6593,N_1866);
nor U17043 (N_17043,N_9508,N_7148);
nand U17044 (N_17044,N_6243,N_8732);
nor U17045 (N_17045,N_5170,N_7277);
nor U17046 (N_17046,N_1626,N_7848);
nand U17047 (N_17047,N_3806,N_3900);
nor U17048 (N_17048,N_8164,N_2298);
nor U17049 (N_17049,N_172,N_5673);
nor U17050 (N_17050,N_4859,N_8296);
or U17051 (N_17051,N_7293,N_3712);
nand U17052 (N_17052,N_3834,N_2485);
and U17053 (N_17053,N_1516,N_9897);
or U17054 (N_17054,N_1975,N_6861);
and U17055 (N_17055,N_905,N_5766);
nor U17056 (N_17056,N_3706,N_9998);
and U17057 (N_17057,N_7909,N_7138);
and U17058 (N_17058,N_4261,N_5937);
and U17059 (N_17059,N_7210,N_3644);
xor U17060 (N_17060,N_3664,N_4523);
and U17061 (N_17061,N_9923,N_5557);
xnor U17062 (N_17062,N_3855,N_8169);
nand U17063 (N_17063,N_7182,N_1724);
nor U17064 (N_17064,N_6480,N_9578);
nor U17065 (N_17065,N_8374,N_9436);
or U17066 (N_17066,N_8587,N_564);
or U17067 (N_17067,N_1007,N_5709);
nand U17068 (N_17068,N_3294,N_4568);
nand U17069 (N_17069,N_4411,N_6497);
and U17070 (N_17070,N_4039,N_3797);
nor U17071 (N_17071,N_3592,N_5912);
nand U17072 (N_17072,N_3034,N_2234);
nand U17073 (N_17073,N_2269,N_3825);
or U17074 (N_17074,N_8384,N_5139);
nor U17075 (N_17075,N_9241,N_1185);
nand U17076 (N_17076,N_2513,N_1015);
and U17077 (N_17077,N_3250,N_8053);
and U17078 (N_17078,N_5763,N_5176);
and U17079 (N_17079,N_7881,N_7760);
or U17080 (N_17080,N_4702,N_9155);
and U17081 (N_17081,N_1675,N_8427);
nand U17082 (N_17082,N_933,N_2557);
nor U17083 (N_17083,N_6952,N_7332);
xnor U17084 (N_17084,N_6099,N_8655);
or U17085 (N_17085,N_5597,N_5378);
nand U17086 (N_17086,N_6836,N_3009);
nor U17087 (N_17087,N_3186,N_8973);
nor U17088 (N_17088,N_5668,N_944);
xnor U17089 (N_17089,N_832,N_1203);
or U17090 (N_17090,N_1237,N_5547);
nand U17091 (N_17091,N_3134,N_8709);
and U17092 (N_17092,N_2195,N_1818);
nand U17093 (N_17093,N_2255,N_6246);
nor U17094 (N_17094,N_1696,N_604);
nor U17095 (N_17095,N_1876,N_7313);
nand U17096 (N_17096,N_1753,N_9626);
or U17097 (N_17097,N_8682,N_5926);
or U17098 (N_17098,N_8888,N_265);
xnor U17099 (N_17099,N_1721,N_8011);
or U17100 (N_17100,N_1519,N_7752);
nor U17101 (N_17101,N_2344,N_942);
or U17102 (N_17102,N_1487,N_7837);
nand U17103 (N_17103,N_4027,N_1903);
nor U17104 (N_17104,N_6618,N_5730);
or U17105 (N_17105,N_9256,N_6498);
nor U17106 (N_17106,N_8018,N_5013);
or U17107 (N_17107,N_3844,N_2430);
nor U17108 (N_17108,N_9977,N_7519);
nor U17109 (N_17109,N_3142,N_7634);
or U17110 (N_17110,N_9599,N_4878);
or U17111 (N_17111,N_3085,N_7911);
and U17112 (N_17112,N_6308,N_9806);
xnor U17113 (N_17113,N_421,N_7088);
nor U17114 (N_17114,N_1355,N_433);
and U17115 (N_17115,N_2574,N_9524);
xnor U17116 (N_17116,N_4639,N_4319);
or U17117 (N_17117,N_74,N_6439);
or U17118 (N_17118,N_5338,N_1351);
and U17119 (N_17119,N_8909,N_3034);
xor U17120 (N_17120,N_3780,N_8848);
xnor U17121 (N_17121,N_7975,N_4279);
nor U17122 (N_17122,N_5790,N_7237);
nor U17123 (N_17123,N_3304,N_7361);
nand U17124 (N_17124,N_5518,N_577);
nand U17125 (N_17125,N_6357,N_2174);
xnor U17126 (N_17126,N_2573,N_3238);
or U17127 (N_17127,N_8513,N_6363);
nand U17128 (N_17128,N_7261,N_2562);
and U17129 (N_17129,N_9063,N_1875);
nand U17130 (N_17130,N_9457,N_3987);
nand U17131 (N_17131,N_1035,N_5362);
nor U17132 (N_17132,N_6226,N_1663);
nor U17133 (N_17133,N_8163,N_7323);
or U17134 (N_17134,N_881,N_1712);
nor U17135 (N_17135,N_6929,N_9674);
nor U17136 (N_17136,N_6951,N_5934);
or U17137 (N_17137,N_4691,N_7611);
nand U17138 (N_17138,N_5941,N_4560);
or U17139 (N_17139,N_4435,N_649);
xnor U17140 (N_17140,N_5749,N_8797);
xor U17141 (N_17141,N_7884,N_7027);
nor U17142 (N_17142,N_4061,N_1796);
and U17143 (N_17143,N_9670,N_7256);
nor U17144 (N_17144,N_9957,N_1563);
nor U17145 (N_17145,N_9286,N_236);
xor U17146 (N_17146,N_9490,N_3202);
nand U17147 (N_17147,N_1341,N_4723);
or U17148 (N_17148,N_9415,N_1129);
nor U17149 (N_17149,N_49,N_4152);
xor U17150 (N_17150,N_2160,N_1154);
nor U17151 (N_17151,N_523,N_8997);
and U17152 (N_17152,N_9044,N_2263);
nor U17153 (N_17153,N_2193,N_531);
nand U17154 (N_17154,N_1769,N_3256);
nand U17155 (N_17155,N_600,N_9959);
nor U17156 (N_17156,N_1634,N_4908);
nor U17157 (N_17157,N_3436,N_8909);
or U17158 (N_17158,N_5482,N_4957);
or U17159 (N_17159,N_1383,N_8072);
and U17160 (N_17160,N_2634,N_6156);
and U17161 (N_17161,N_9887,N_3263);
xor U17162 (N_17162,N_507,N_1865);
nor U17163 (N_17163,N_8832,N_9003);
nor U17164 (N_17164,N_8654,N_898);
and U17165 (N_17165,N_9365,N_7138);
nand U17166 (N_17166,N_1683,N_1414);
or U17167 (N_17167,N_7987,N_4133);
and U17168 (N_17168,N_858,N_9783);
and U17169 (N_17169,N_1931,N_7719);
nand U17170 (N_17170,N_2373,N_6177);
nor U17171 (N_17171,N_7303,N_4879);
or U17172 (N_17172,N_9724,N_3413);
nor U17173 (N_17173,N_8151,N_4855);
and U17174 (N_17174,N_5903,N_8916);
xnor U17175 (N_17175,N_6247,N_814);
nand U17176 (N_17176,N_7325,N_839);
or U17177 (N_17177,N_64,N_6923);
xnor U17178 (N_17178,N_8931,N_5197);
nand U17179 (N_17179,N_522,N_1859);
nor U17180 (N_17180,N_5313,N_3201);
nor U17181 (N_17181,N_6298,N_9657);
and U17182 (N_17182,N_2206,N_7778);
or U17183 (N_17183,N_6878,N_9112);
nand U17184 (N_17184,N_3308,N_1578);
xor U17185 (N_17185,N_2282,N_9382);
xnor U17186 (N_17186,N_574,N_120);
nor U17187 (N_17187,N_6683,N_6771);
or U17188 (N_17188,N_3222,N_6872);
or U17189 (N_17189,N_5994,N_1614);
and U17190 (N_17190,N_2318,N_8225);
nand U17191 (N_17191,N_3654,N_1522);
xnor U17192 (N_17192,N_1609,N_5203);
nor U17193 (N_17193,N_2617,N_5236);
or U17194 (N_17194,N_479,N_1069);
xnor U17195 (N_17195,N_1751,N_3461);
nor U17196 (N_17196,N_6218,N_1215);
nor U17197 (N_17197,N_9161,N_4998);
or U17198 (N_17198,N_6805,N_1731);
and U17199 (N_17199,N_3008,N_726);
nand U17200 (N_17200,N_470,N_9741);
and U17201 (N_17201,N_852,N_9);
nor U17202 (N_17202,N_9883,N_369);
nor U17203 (N_17203,N_3625,N_2856);
or U17204 (N_17204,N_3474,N_3294);
nand U17205 (N_17205,N_7604,N_7362);
nand U17206 (N_17206,N_8269,N_5025);
and U17207 (N_17207,N_8309,N_1655);
or U17208 (N_17208,N_8208,N_4670);
xnor U17209 (N_17209,N_5224,N_3293);
and U17210 (N_17210,N_9326,N_6611);
and U17211 (N_17211,N_2629,N_341);
or U17212 (N_17212,N_379,N_8816);
and U17213 (N_17213,N_5570,N_7093);
or U17214 (N_17214,N_4958,N_973);
xnor U17215 (N_17215,N_197,N_265);
xnor U17216 (N_17216,N_465,N_8439);
nand U17217 (N_17217,N_8379,N_2771);
xor U17218 (N_17218,N_2669,N_1665);
nand U17219 (N_17219,N_373,N_7250);
or U17220 (N_17220,N_9514,N_1736);
and U17221 (N_17221,N_8101,N_4892);
nor U17222 (N_17222,N_1194,N_3467);
xnor U17223 (N_17223,N_669,N_3185);
xor U17224 (N_17224,N_8530,N_7818);
nor U17225 (N_17225,N_1054,N_477);
xor U17226 (N_17226,N_8508,N_1590);
and U17227 (N_17227,N_1610,N_8116);
or U17228 (N_17228,N_3547,N_9253);
xnor U17229 (N_17229,N_3294,N_8837);
nand U17230 (N_17230,N_881,N_7890);
and U17231 (N_17231,N_4155,N_6153);
xor U17232 (N_17232,N_8674,N_8515);
nand U17233 (N_17233,N_3022,N_5619);
nor U17234 (N_17234,N_2029,N_1234);
or U17235 (N_17235,N_2724,N_645);
and U17236 (N_17236,N_1066,N_8338);
or U17237 (N_17237,N_7207,N_6957);
nand U17238 (N_17238,N_5521,N_3259);
and U17239 (N_17239,N_4863,N_4138);
or U17240 (N_17240,N_3899,N_3904);
xnor U17241 (N_17241,N_488,N_3634);
xnor U17242 (N_17242,N_5845,N_7679);
nor U17243 (N_17243,N_306,N_7044);
xnor U17244 (N_17244,N_7408,N_9087);
nor U17245 (N_17245,N_894,N_4137);
nor U17246 (N_17246,N_7154,N_6529);
nand U17247 (N_17247,N_4910,N_6033);
xnor U17248 (N_17248,N_4819,N_4129);
nand U17249 (N_17249,N_4191,N_7026);
nand U17250 (N_17250,N_6766,N_5618);
nor U17251 (N_17251,N_2770,N_8483);
and U17252 (N_17252,N_2632,N_6193);
and U17253 (N_17253,N_9607,N_5654);
and U17254 (N_17254,N_9134,N_4177);
nand U17255 (N_17255,N_7910,N_2191);
and U17256 (N_17256,N_9114,N_3242);
and U17257 (N_17257,N_6398,N_452);
nor U17258 (N_17258,N_9604,N_8328);
nor U17259 (N_17259,N_4076,N_7070);
and U17260 (N_17260,N_426,N_5261);
or U17261 (N_17261,N_7021,N_5096);
nand U17262 (N_17262,N_8642,N_5782);
or U17263 (N_17263,N_2359,N_7734);
or U17264 (N_17264,N_771,N_1060);
nor U17265 (N_17265,N_855,N_5003);
and U17266 (N_17266,N_4168,N_3979);
or U17267 (N_17267,N_7968,N_4593);
nand U17268 (N_17268,N_7102,N_3884);
nand U17269 (N_17269,N_7544,N_1924);
nand U17270 (N_17270,N_3507,N_7292);
xnor U17271 (N_17271,N_3438,N_172);
nand U17272 (N_17272,N_7901,N_1756);
nor U17273 (N_17273,N_6064,N_2644);
and U17274 (N_17274,N_9699,N_5930);
nand U17275 (N_17275,N_2583,N_7322);
nand U17276 (N_17276,N_2400,N_4249);
xor U17277 (N_17277,N_2786,N_4241);
nor U17278 (N_17278,N_7278,N_3098);
and U17279 (N_17279,N_8602,N_6042);
xor U17280 (N_17280,N_616,N_2900);
and U17281 (N_17281,N_8275,N_4046);
or U17282 (N_17282,N_2687,N_6864);
and U17283 (N_17283,N_2985,N_4393);
nand U17284 (N_17284,N_4551,N_1116);
and U17285 (N_17285,N_3241,N_1770);
and U17286 (N_17286,N_2985,N_4635);
xnor U17287 (N_17287,N_5116,N_3629);
xnor U17288 (N_17288,N_4742,N_5452);
and U17289 (N_17289,N_473,N_5832);
xor U17290 (N_17290,N_1912,N_8824);
xor U17291 (N_17291,N_5202,N_4043);
or U17292 (N_17292,N_7281,N_9559);
and U17293 (N_17293,N_7451,N_77);
xor U17294 (N_17294,N_3429,N_8215);
nor U17295 (N_17295,N_8916,N_6563);
and U17296 (N_17296,N_3453,N_5739);
nor U17297 (N_17297,N_8224,N_8816);
nor U17298 (N_17298,N_2390,N_4747);
nor U17299 (N_17299,N_5110,N_179);
nor U17300 (N_17300,N_1727,N_2160);
nor U17301 (N_17301,N_4882,N_7474);
nand U17302 (N_17302,N_6765,N_1192);
nor U17303 (N_17303,N_3296,N_40);
or U17304 (N_17304,N_5980,N_6114);
and U17305 (N_17305,N_7356,N_4126);
nand U17306 (N_17306,N_8870,N_5671);
and U17307 (N_17307,N_9533,N_9345);
nand U17308 (N_17308,N_4413,N_664);
and U17309 (N_17309,N_3946,N_8074);
or U17310 (N_17310,N_553,N_3881);
nor U17311 (N_17311,N_5730,N_4026);
or U17312 (N_17312,N_4617,N_1441);
xnor U17313 (N_17313,N_9500,N_673);
xnor U17314 (N_17314,N_8410,N_4679);
nand U17315 (N_17315,N_9840,N_9398);
xnor U17316 (N_17316,N_7177,N_1617);
nor U17317 (N_17317,N_7805,N_8213);
or U17318 (N_17318,N_5503,N_5390);
xor U17319 (N_17319,N_7813,N_7132);
nand U17320 (N_17320,N_1739,N_6561);
nand U17321 (N_17321,N_3410,N_6068);
or U17322 (N_17322,N_4787,N_8492);
nor U17323 (N_17323,N_155,N_8247);
xnor U17324 (N_17324,N_7845,N_4575);
or U17325 (N_17325,N_8588,N_8904);
nor U17326 (N_17326,N_7173,N_8067);
xnor U17327 (N_17327,N_8317,N_8829);
nand U17328 (N_17328,N_3571,N_9045);
and U17329 (N_17329,N_5358,N_7655);
xor U17330 (N_17330,N_9844,N_4212);
and U17331 (N_17331,N_1071,N_5939);
nand U17332 (N_17332,N_8537,N_5072);
nand U17333 (N_17333,N_4190,N_5204);
or U17334 (N_17334,N_6129,N_8667);
nor U17335 (N_17335,N_817,N_771);
nor U17336 (N_17336,N_1259,N_7728);
nor U17337 (N_17337,N_1569,N_3512);
xor U17338 (N_17338,N_5815,N_6345);
nor U17339 (N_17339,N_8727,N_1663);
nor U17340 (N_17340,N_4048,N_586);
and U17341 (N_17341,N_166,N_5826);
xnor U17342 (N_17342,N_701,N_7390);
or U17343 (N_17343,N_8612,N_8120);
and U17344 (N_17344,N_200,N_9506);
nor U17345 (N_17345,N_2240,N_2933);
or U17346 (N_17346,N_1176,N_9288);
nand U17347 (N_17347,N_6787,N_8984);
or U17348 (N_17348,N_5514,N_8166);
and U17349 (N_17349,N_2324,N_5179);
and U17350 (N_17350,N_9580,N_8758);
nor U17351 (N_17351,N_1649,N_7676);
or U17352 (N_17352,N_9545,N_9057);
nor U17353 (N_17353,N_9682,N_940);
or U17354 (N_17354,N_8897,N_797);
or U17355 (N_17355,N_9100,N_7720);
xor U17356 (N_17356,N_1724,N_2605);
and U17357 (N_17357,N_879,N_6466);
or U17358 (N_17358,N_992,N_1903);
or U17359 (N_17359,N_6014,N_2648);
nor U17360 (N_17360,N_9079,N_2072);
xnor U17361 (N_17361,N_1339,N_9663);
xnor U17362 (N_17362,N_2248,N_3498);
nor U17363 (N_17363,N_9056,N_7014);
and U17364 (N_17364,N_6764,N_9632);
and U17365 (N_17365,N_8809,N_2930);
nor U17366 (N_17366,N_128,N_957);
and U17367 (N_17367,N_3945,N_7607);
or U17368 (N_17368,N_8575,N_6222);
or U17369 (N_17369,N_6966,N_1203);
nand U17370 (N_17370,N_4186,N_7838);
nand U17371 (N_17371,N_7530,N_9020);
xor U17372 (N_17372,N_9174,N_2157);
or U17373 (N_17373,N_1484,N_8075);
and U17374 (N_17374,N_6937,N_3818);
or U17375 (N_17375,N_1131,N_6451);
xnor U17376 (N_17376,N_5794,N_6012);
or U17377 (N_17377,N_9854,N_7109);
xnor U17378 (N_17378,N_6507,N_5325);
xnor U17379 (N_17379,N_5499,N_1899);
nand U17380 (N_17380,N_7913,N_6551);
xor U17381 (N_17381,N_69,N_9595);
xnor U17382 (N_17382,N_2245,N_7808);
nor U17383 (N_17383,N_1737,N_9792);
xnor U17384 (N_17384,N_5761,N_6495);
and U17385 (N_17385,N_6587,N_6410);
nor U17386 (N_17386,N_3346,N_6547);
and U17387 (N_17387,N_8595,N_2795);
or U17388 (N_17388,N_5878,N_3495);
or U17389 (N_17389,N_6151,N_4182);
xor U17390 (N_17390,N_8945,N_4482);
nor U17391 (N_17391,N_127,N_8201);
xor U17392 (N_17392,N_5319,N_7616);
nor U17393 (N_17393,N_5514,N_2221);
xor U17394 (N_17394,N_6135,N_6982);
xnor U17395 (N_17395,N_9285,N_9964);
xnor U17396 (N_17396,N_5566,N_1312);
nand U17397 (N_17397,N_5947,N_1608);
nor U17398 (N_17398,N_7841,N_7187);
xnor U17399 (N_17399,N_1213,N_3066);
nand U17400 (N_17400,N_2661,N_3852);
xor U17401 (N_17401,N_3246,N_1302);
and U17402 (N_17402,N_9415,N_1447);
xnor U17403 (N_17403,N_7407,N_3044);
nand U17404 (N_17404,N_2832,N_5628);
and U17405 (N_17405,N_4368,N_2815);
xor U17406 (N_17406,N_5976,N_1730);
xnor U17407 (N_17407,N_4887,N_8142);
nand U17408 (N_17408,N_4522,N_3681);
xnor U17409 (N_17409,N_8093,N_9895);
nand U17410 (N_17410,N_4310,N_944);
xnor U17411 (N_17411,N_2073,N_3025);
nand U17412 (N_17412,N_3091,N_3223);
or U17413 (N_17413,N_4431,N_9431);
nand U17414 (N_17414,N_1082,N_2372);
nor U17415 (N_17415,N_5657,N_2649);
xnor U17416 (N_17416,N_621,N_6898);
or U17417 (N_17417,N_4347,N_7570);
nor U17418 (N_17418,N_4332,N_4728);
and U17419 (N_17419,N_8975,N_3490);
nand U17420 (N_17420,N_1826,N_1783);
or U17421 (N_17421,N_4263,N_9533);
nand U17422 (N_17422,N_9889,N_8399);
nand U17423 (N_17423,N_8843,N_3156);
or U17424 (N_17424,N_2067,N_3915);
xnor U17425 (N_17425,N_580,N_7473);
nor U17426 (N_17426,N_811,N_9082);
or U17427 (N_17427,N_2115,N_3676);
or U17428 (N_17428,N_8153,N_7223);
xor U17429 (N_17429,N_7808,N_55);
or U17430 (N_17430,N_2144,N_7832);
xor U17431 (N_17431,N_9648,N_6290);
xor U17432 (N_17432,N_9647,N_804);
xnor U17433 (N_17433,N_4221,N_5460);
nand U17434 (N_17434,N_9749,N_3475);
nand U17435 (N_17435,N_3097,N_6480);
nor U17436 (N_17436,N_5592,N_5109);
xnor U17437 (N_17437,N_9647,N_8243);
or U17438 (N_17438,N_2225,N_459);
and U17439 (N_17439,N_8534,N_8540);
xor U17440 (N_17440,N_8599,N_5751);
nand U17441 (N_17441,N_953,N_401);
and U17442 (N_17442,N_1890,N_7811);
or U17443 (N_17443,N_7630,N_1212);
nand U17444 (N_17444,N_4878,N_4894);
nand U17445 (N_17445,N_7167,N_8990);
or U17446 (N_17446,N_5708,N_9842);
nor U17447 (N_17447,N_3766,N_9725);
xor U17448 (N_17448,N_7375,N_3366);
or U17449 (N_17449,N_1774,N_9743);
nor U17450 (N_17450,N_1083,N_9179);
nand U17451 (N_17451,N_7369,N_2860);
and U17452 (N_17452,N_2323,N_2182);
nand U17453 (N_17453,N_6321,N_4440);
nand U17454 (N_17454,N_2908,N_1236);
or U17455 (N_17455,N_3840,N_5230);
and U17456 (N_17456,N_7936,N_4564);
and U17457 (N_17457,N_3788,N_8333);
and U17458 (N_17458,N_812,N_5648);
xor U17459 (N_17459,N_1700,N_8348);
xnor U17460 (N_17460,N_1474,N_1240);
xnor U17461 (N_17461,N_8690,N_4222);
nand U17462 (N_17462,N_1305,N_5910);
nor U17463 (N_17463,N_6387,N_9389);
xnor U17464 (N_17464,N_1392,N_3105);
nand U17465 (N_17465,N_5664,N_7001);
xnor U17466 (N_17466,N_3651,N_2245);
nand U17467 (N_17467,N_7514,N_9279);
nand U17468 (N_17468,N_5893,N_7929);
xnor U17469 (N_17469,N_6897,N_2186);
or U17470 (N_17470,N_5913,N_9538);
nand U17471 (N_17471,N_1619,N_6420);
or U17472 (N_17472,N_238,N_8503);
or U17473 (N_17473,N_6315,N_9637);
and U17474 (N_17474,N_3152,N_7518);
nor U17475 (N_17475,N_2123,N_5088);
nand U17476 (N_17476,N_1572,N_7971);
xnor U17477 (N_17477,N_5270,N_487);
nor U17478 (N_17478,N_3336,N_8748);
nand U17479 (N_17479,N_1269,N_8282);
and U17480 (N_17480,N_9866,N_8387);
and U17481 (N_17481,N_2826,N_9024);
xnor U17482 (N_17482,N_9274,N_9376);
and U17483 (N_17483,N_6421,N_9043);
and U17484 (N_17484,N_9151,N_8699);
nand U17485 (N_17485,N_8856,N_454);
or U17486 (N_17486,N_984,N_2263);
or U17487 (N_17487,N_9289,N_2780);
and U17488 (N_17488,N_7134,N_6110);
nand U17489 (N_17489,N_5986,N_1634);
nor U17490 (N_17490,N_9815,N_307);
or U17491 (N_17491,N_6789,N_9718);
or U17492 (N_17492,N_7201,N_8990);
nor U17493 (N_17493,N_1350,N_4356);
and U17494 (N_17494,N_3818,N_4797);
nand U17495 (N_17495,N_8008,N_9684);
nand U17496 (N_17496,N_8240,N_7887);
nand U17497 (N_17497,N_7750,N_9210);
nor U17498 (N_17498,N_3125,N_2361);
nor U17499 (N_17499,N_2789,N_6220);
or U17500 (N_17500,N_1165,N_7873);
xnor U17501 (N_17501,N_1982,N_7691);
and U17502 (N_17502,N_9405,N_2333);
xnor U17503 (N_17503,N_2275,N_2415);
xnor U17504 (N_17504,N_1516,N_9789);
or U17505 (N_17505,N_6076,N_2748);
nand U17506 (N_17506,N_8482,N_1150);
nand U17507 (N_17507,N_5849,N_6354);
nor U17508 (N_17508,N_5955,N_1522);
or U17509 (N_17509,N_1060,N_8192);
xor U17510 (N_17510,N_6766,N_3391);
nand U17511 (N_17511,N_1908,N_9896);
xnor U17512 (N_17512,N_8931,N_4366);
xor U17513 (N_17513,N_3474,N_3334);
and U17514 (N_17514,N_838,N_7251);
or U17515 (N_17515,N_5563,N_5461);
or U17516 (N_17516,N_6255,N_9350);
xnor U17517 (N_17517,N_1748,N_9713);
xnor U17518 (N_17518,N_3498,N_2714);
and U17519 (N_17519,N_3707,N_5518);
or U17520 (N_17520,N_1988,N_221);
nand U17521 (N_17521,N_639,N_2161);
nor U17522 (N_17522,N_2228,N_7228);
nand U17523 (N_17523,N_5360,N_1844);
nor U17524 (N_17524,N_6422,N_3825);
xnor U17525 (N_17525,N_9225,N_438);
and U17526 (N_17526,N_9793,N_4666);
nor U17527 (N_17527,N_8889,N_6426);
nand U17528 (N_17528,N_9300,N_656);
nor U17529 (N_17529,N_8053,N_5877);
xor U17530 (N_17530,N_1610,N_9651);
xor U17531 (N_17531,N_1149,N_8419);
and U17532 (N_17532,N_309,N_918);
nor U17533 (N_17533,N_878,N_1246);
and U17534 (N_17534,N_149,N_1511);
nand U17535 (N_17535,N_7085,N_773);
nor U17536 (N_17536,N_8174,N_2617);
and U17537 (N_17537,N_1534,N_9782);
nor U17538 (N_17538,N_9951,N_6115);
nor U17539 (N_17539,N_1442,N_8578);
or U17540 (N_17540,N_1668,N_3955);
nor U17541 (N_17541,N_2880,N_8048);
and U17542 (N_17542,N_6120,N_4175);
or U17543 (N_17543,N_2816,N_6954);
xor U17544 (N_17544,N_5692,N_3755);
nor U17545 (N_17545,N_4232,N_5097);
nand U17546 (N_17546,N_4216,N_4071);
nand U17547 (N_17547,N_3747,N_9819);
xnor U17548 (N_17548,N_4478,N_5259);
xnor U17549 (N_17549,N_2709,N_4421);
nand U17550 (N_17550,N_786,N_6125);
nor U17551 (N_17551,N_3560,N_2058);
xnor U17552 (N_17552,N_6447,N_9764);
and U17553 (N_17553,N_1547,N_706);
xor U17554 (N_17554,N_3453,N_2442);
and U17555 (N_17555,N_7299,N_8683);
nand U17556 (N_17556,N_680,N_5688);
or U17557 (N_17557,N_9817,N_786);
nand U17558 (N_17558,N_9105,N_2162);
and U17559 (N_17559,N_1824,N_7467);
or U17560 (N_17560,N_7267,N_6588);
nor U17561 (N_17561,N_1109,N_8714);
and U17562 (N_17562,N_249,N_7578);
xor U17563 (N_17563,N_9752,N_9988);
or U17564 (N_17564,N_5626,N_5864);
nand U17565 (N_17565,N_4207,N_4505);
xnor U17566 (N_17566,N_990,N_8571);
nor U17567 (N_17567,N_5186,N_600);
xor U17568 (N_17568,N_5991,N_3500);
xnor U17569 (N_17569,N_1112,N_9070);
xor U17570 (N_17570,N_2978,N_2318);
or U17571 (N_17571,N_8696,N_6494);
xor U17572 (N_17572,N_5009,N_64);
and U17573 (N_17573,N_3073,N_9849);
xor U17574 (N_17574,N_7823,N_7917);
and U17575 (N_17575,N_5419,N_5822);
or U17576 (N_17576,N_2936,N_3907);
or U17577 (N_17577,N_9367,N_271);
nand U17578 (N_17578,N_2923,N_3001);
nand U17579 (N_17579,N_5590,N_4995);
and U17580 (N_17580,N_7751,N_9012);
xnor U17581 (N_17581,N_225,N_8964);
and U17582 (N_17582,N_2379,N_4707);
nor U17583 (N_17583,N_9194,N_2692);
or U17584 (N_17584,N_4330,N_9444);
nor U17585 (N_17585,N_4661,N_1785);
nand U17586 (N_17586,N_8225,N_8480);
or U17587 (N_17587,N_3065,N_7803);
nand U17588 (N_17588,N_5375,N_872);
or U17589 (N_17589,N_2431,N_9814);
and U17590 (N_17590,N_294,N_609);
and U17591 (N_17591,N_3505,N_3204);
nor U17592 (N_17592,N_9321,N_5147);
xor U17593 (N_17593,N_7098,N_1614);
nor U17594 (N_17594,N_7139,N_4650);
nand U17595 (N_17595,N_3900,N_5152);
nor U17596 (N_17596,N_195,N_309);
and U17597 (N_17597,N_9307,N_2895);
and U17598 (N_17598,N_2931,N_7088);
or U17599 (N_17599,N_3126,N_2064);
xnor U17600 (N_17600,N_4236,N_664);
and U17601 (N_17601,N_4745,N_9888);
xor U17602 (N_17602,N_4951,N_9703);
nand U17603 (N_17603,N_7378,N_1643);
nor U17604 (N_17604,N_6823,N_4100);
and U17605 (N_17605,N_286,N_7121);
nand U17606 (N_17606,N_1422,N_5029);
nand U17607 (N_17607,N_4449,N_435);
xnor U17608 (N_17608,N_3383,N_3649);
nor U17609 (N_17609,N_809,N_5718);
and U17610 (N_17610,N_5762,N_5753);
nor U17611 (N_17611,N_4389,N_7307);
or U17612 (N_17612,N_1042,N_1527);
nor U17613 (N_17613,N_813,N_6797);
xor U17614 (N_17614,N_1369,N_8132);
and U17615 (N_17615,N_1490,N_3464);
or U17616 (N_17616,N_4959,N_2047);
nor U17617 (N_17617,N_8420,N_1363);
nor U17618 (N_17618,N_201,N_5545);
or U17619 (N_17619,N_6189,N_9373);
xnor U17620 (N_17620,N_3796,N_2421);
nor U17621 (N_17621,N_5889,N_4847);
and U17622 (N_17622,N_3699,N_3832);
nand U17623 (N_17623,N_7051,N_56);
or U17624 (N_17624,N_700,N_8862);
nand U17625 (N_17625,N_9705,N_6490);
and U17626 (N_17626,N_4721,N_745);
or U17627 (N_17627,N_8185,N_9705);
and U17628 (N_17628,N_7741,N_2600);
nor U17629 (N_17629,N_355,N_315);
xnor U17630 (N_17630,N_5080,N_6582);
and U17631 (N_17631,N_4595,N_5792);
xnor U17632 (N_17632,N_2,N_3628);
or U17633 (N_17633,N_8437,N_9176);
or U17634 (N_17634,N_3258,N_8212);
or U17635 (N_17635,N_7467,N_9698);
xnor U17636 (N_17636,N_3499,N_8429);
xor U17637 (N_17637,N_9563,N_5328);
xnor U17638 (N_17638,N_1188,N_4490);
or U17639 (N_17639,N_318,N_8695);
nand U17640 (N_17640,N_2105,N_3096);
nor U17641 (N_17641,N_4882,N_3816);
and U17642 (N_17642,N_2174,N_1871);
and U17643 (N_17643,N_3068,N_3709);
and U17644 (N_17644,N_7126,N_3602);
nor U17645 (N_17645,N_6161,N_9340);
nor U17646 (N_17646,N_816,N_5247);
nor U17647 (N_17647,N_2203,N_4019);
nor U17648 (N_17648,N_9288,N_9041);
or U17649 (N_17649,N_2974,N_6018);
nand U17650 (N_17650,N_4097,N_254);
or U17651 (N_17651,N_9055,N_4589);
nor U17652 (N_17652,N_7812,N_6121);
or U17653 (N_17653,N_1571,N_3159);
nand U17654 (N_17654,N_5194,N_6422);
or U17655 (N_17655,N_9006,N_6040);
or U17656 (N_17656,N_6383,N_2578);
or U17657 (N_17657,N_8666,N_3220);
and U17658 (N_17658,N_9417,N_1719);
xor U17659 (N_17659,N_1622,N_2217);
nor U17660 (N_17660,N_4152,N_894);
nand U17661 (N_17661,N_1818,N_1564);
nor U17662 (N_17662,N_2892,N_4940);
nor U17663 (N_17663,N_4345,N_9106);
xnor U17664 (N_17664,N_3674,N_3970);
and U17665 (N_17665,N_5154,N_5234);
nand U17666 (N_17666,N_2420,N_134);
nor U17667 (N_17667,N_5334,N_9460);
and U17668 (N_17668,N_2247,N_3950);
xnor U17669 (N_17669,N_448,N_6504);
and U17670 (N_17670,N_5759,N_6876);
nor U17671 (N_17671,N_5211,N_8112);
nor U17672 (N_17672,N_3296,N_8087);
xor U17673 (N_17673,N_1028,N_9499);
xnor U17674 (N_17674,N_1937,N_678);
and U17675 (N_17675,N_8072,N_9936);
nand U17676 (N_17676,N_2011,N_4606);
xnor U17677 (N_17677,N_9684,N_4179);
or U17678 (N_17678,N_9848,N_208);
nand U17679 (N_17679,N_784,N_9792);
and U17680 (N_17680,N_922,N_2781);
nor U17681 (N_17681,N_1556,N_4852);
or U17682 (N_17682,N_9294,N_8174);
or U17683 (N_17683,N_217,N_4405);
nand U17684 (N_17684,N_6001,N_3347);
nor U17685 (N_17685,N_8515,N_4595);
and U17686 (N_17686,N_4382,N_2523);
xor U17687 (N_17687,N_2460,N_2270);
or U17688 (N_17688,N_6488,N_8463);
nor U17689 (N_17689,N_9190,N_9837);
and U17690 (N_17690,N_3583,N_2586);
xnor U17691 (N_17691,N_6613,N_9458);
and U17692 (N_17692,N_906,N_965);
or U17693 (N_17693,N_7114,N_7879);
or U17694 (N_17694,N_8112,N_6113);
nand U17695 (N_17695,N_5412,N_7428);
xnor U17696 (N_17696,N_2027,N_8857);
xor U17697 (N_17697,N_9574,N_6329);
and U17698 (N_17698,N_3717,N_2639);
nor U17699 (N_17699,N_7343,N_3230);
nor U17700 (N_17700,N_8690,N_3278);
and U17701 (N_17701,N_6552,N_9074);
and U17702 (N_17702,N_3911,N_4002);
nor U17703 (N_17703,N_7044,N_1576);
xnor U17704 (N_17704,N_6112,N_5517);
nor U17705 (N_17705,N_1366,N_3418);
and U17706 (N_17706,N_9903,N_6880);
and U17707 (N_17707,N_5110,N_6348);
and U17708 (N_17708,N_7541,N_7837);
or U17709 (N_17709,N_858,N_3424);
or U17710 (N_17710,N_8708,N_4533);
nor U17711 (N_17711,N_6443,N_8536);
nand U17712 (N_17712,N_5039,N_9999);
nand U17713 (N_17713,N_4630,N_5012);
nor U17714 (N_17714,N_7843,N_7097);
and U17715 (N_17715,N_3347,N_2665);
or U17716 (N_17716,N_2795,N_1998);
nand U17717 (N_17717,N_2159,N_4950);
or U17718 (N_17718,N_2024,N_5428);
or U17719 (N_17719,N_4216,N_7370);
nand U17720 (N_17720,N_6309,N_2473);
xnor U17721 (N_17721,N_8248,N_8735);
nor U17722 (N_17722,N_5533,N_2865);
xor U17723 (N_17723,N_7825,N_5928);
and U17724 (N_17724,N_3918,N_2530);
nor U17725 (N_17725,N_4808,N_6288);
xnor U17726 (N_17726,N_3336,N_5976);
nor U17727 (N_17727,N_8525,N_5383);
xnor U17728 (N_17728,N_8630,N_2664);
nand U17729 (N_17729,N_9458,N_9982);
or U17730 (N_17730,N_5658,N_7608);
xnor U17731 (N_17731,N_4935,N_7507);
or U17732 (N_17732,N_9770,N_6254);
or U17733 (N_17733,N_838,N_9422);
xnor U17734 (N_17734,N_5153,N_2280);
nor U17735 (N_17735,N_4701,N_810);
or U17736 (N_17736,N_4721,N_787);
nor U17737 (N_17737,N_6697,N_7770);
nor U17738 (N_17738,N_9656,N_542);
nor U17739 (N_17739,N_9640,N_4019);
nand U17740 (N_17740,N_9183,N_4193);
or U17741 (N_17741,N_8326,N_4333);
or U17742 (N_17742,N_1861,N_692);
or U17743 (N_17743,N_8186,N_870);
and U17744 (N_17744,N_6192,N_4738);
nand U17745 (N_17745,N_3336,N_7763);
and U17746 (N_17746,N_6211,N_6651);
and U17747 (N_17747,N_9906,N_1359);
or U17748 (N_17748,N_4481,N_403);
or U17749 (N_17749,N_7306,N_291);
or U17750 (N_17750,N_4420,N_256);
or U17751 (N_17751,N_57,N_4708);
xnor U17752 (N_17752,N_175,N_3628);
or U17753 (N_17753,N_1519,N_9171);
xor U17754 (N_17754,N_5755,N_5536);
nand U17755 (N_17755,N_5105,N_4697);
nand U17756 (N_17756,N_7963,N_2957);
xor U17757 (N_17757,N_4836,N_2771);
nand U17758 (N_17758,N_53,N_4840);
xor U17759 (N_17759,N_8628,N_2503);
nor U17760 (N_17760,N_3754,N_8596);
xor U17761 (N_17761,N_6892,N_5551);
nor U17762 (N_17762,N_4202,N_1165);
nor U17763 (N_17763,N_1515,N_2317);
nor U17764 (N_17764,N_3076,N_5109);
and U17765 (N_17765,N_7346,N_8168);
xor U17766 (N_17766,N_7460,N_7016);
nor U17767 (N_17767,N_7409,N_6463);
and U17768 (N_17768,N_9714,N_1737);
and U17769 (N_17769,N_7738,N_9019);
or U17770 (N_17770,N_3015,N_6720);
nor U17771 (N_17771,N_8192,N_8749);
or U17772 (N_17772,N_1908,N_4962);
nor U17773 (N_17773,N_330,N_9747);
or U17774 (N_17774,N_5927,N_6638);
nand U17775 (N_17775,N_471,N_7011);
nand U17776 (N_17776,N_7647,N_7193);
xnor U17777 (N_17777,N_4527,N_3687);
xor U17778 (N_17778,N_9243,N_9524);
xnor U17779 (N_17779,N_3656,N_1504);
nand U17780 (N_17780,N_6373,N_151);
and U17781 (N_17781,N_7571,N_5602);
nor U17782 (N_17782,N_1326,N_1537);
and U17783 (N_17783,N_6081,N_9644);
and U17784 (N_17784,N_1461,N_947);
or U17785 (N_17785,N_5612,N_263);
or U17786 (N_17786,N_3988,N_9303);
xnor U17787 (N_17787,N_8281,N_9380);
and U17788 (N_17788,N_2846,N_366);
nand U17789 (N_17789,N_9237,N_8234);
and U17790 (N_17790,N_9100,N_6424);
xor U17791 (N_17791,N_1014,N_464);
nor U17792 (N_17792,N_2538,N_7975);
xnor U17793 (N_17793,N_6293,N_747);
xnor U17794 (N_17794,N_1219,N_7751);
xor U17795 (N_17795,N_3343,N_6458);
and U17796 (N_17796,N_3130,N_7560);
and U17797 (N_17797,N_4973,N_3260);
xnor U17798 (N_17798,N_1555,N_7146);
xnor U17799 (N_17799,N_6402,N_4344);
xor U17800 (N_17800,N_5776,N_7307);
nand U17801 (N_17801,N_9395,N_3898);
nand U17802 (N_17802,N_4118,N_5898);
nand U17803 (N_17803,N_6011,N_5465);
xor U17804 (N_17804,N_2817,N_2512);
nor U17805 (N_17805,N_8915,N_1373);
or U17806 (N_17806,N_2127,N_8567);
and U17807 (N_17807,N_3746,N_9529);
and U17808 (N_17808,N_1784,N_4528);
nor U17809 (N_17809,N_3410,N_7890);
or U17810 (N_17810,N_8604,N_4587);
or U17811 (N_17811,N_2170,N_1385);
nor U17812 (N_17812,N_4568,N_6616);
nor U17813 (N_17813,N_2553,N_6749);
and U17814 (N_17814,N_7941,N_7894);
nand U17815 (N_17815,N_2716,N_8841);
and U17816 (N_17816,N_4862,N_5903);
or U17817 (N_17817,N_3345,N_7387);
and U17818 (N_17818,N_555,N_4011);
nand U17819 (N_17819,N_2703,N_3693);
nand U17820 (N_17820,N_2368,N_4806);
and U17821 (N_17821,N_4335,N_4246);
nand U17822 (N_17822,N_2157,N_5654);
or U17823 (N_17823,N_9628,N_698);
or U17824 (N_17824,N_4866,N_4981);
nand U17825 (N_17825,N_2039,N_5486);
and U17826 (N_17826,N_4215,N_5478);
xor U17827 (N_17827,N_479,N_4895);
nor U17828 (N_17828,N_8659,N_5801);
and U17829 (N_17829,N_3020,N_5107);
nand U17830 (N_17830,N_4973,N_7953);
xor U17831 (N_17831,N_8456,N_2023);
nor U17832 (N_17832,N_14,N_370);
or U17833 (N_17833,N_512,N_7232);
nor U17834 (N_17834,N_7756,N_2681);
nand U17835 (N_17835,N_150,N_4591);
nand U17836 (N_17836,N_1360,N_9403);
or U17837 (N_17837,N_4861,N_6045);
or U17838 (N_17838,N_361,N_8430);
xnor U17839 (N_17839,N_5851,N_7621);
xnor U17840 (N_17840,N_8657,N_6802);
xor U17841 (N_17841,N_3911,N_4064);
xor U17842 (N_17842,N_2720,N_1088);
xor U17843 (N_17843,N_135,N_9041);
nand U17844 (N_17844,N_9975,N_9978);
and U17845 (N_17845,N_6084,N_5174);
nand U17846 (N_17846,N_5148,N_6214);
nor U17847 (N_17847,N_6955,N_801);
nand U17848 (N_17848,N_696,N_6419);
or U17849 (N_17849,N_3219,N_2064);
xnor U17850 (N_17850,N_8520,N_8323);
or U17851 (N_17851,N_492,N_8578);
nor U17852 (N_17852,N_9440,N_1494);
or U17853 (N_17853,N_623,N_1347);
or U17854 (N_17854,N_3129,N_8395);
nor U17855 (N_17855,N_6868,N_1807);
xor U17856 (N_17856,N_1423,N_8432);
nand U17857 (N_17857,N_4414,N_6422);
nand U17858 (N_17858,N_1195,N_6584);
nor U17859 (N_17859,N_9341,N_6658);
or U17860 (N_17860,N_6177,N_7470);
and U17861 (N_17861,N_8688,N_686);
nand U17862 (N_17862,N_2918,N_7485);
and U17863 (N_17863,N_5457,N_4447);
nand U17864 (N_17864,N_8723,N_5491);
nand U17865 (N_17865,N_7945,N_839);
or U17866 (N_17866,N_1004,N_4981);
or U17867 (N_17867,N_892,N_9131);
and U17868 (N_17868,N_9770,N_8069);
or U17869 (N_17869,N_2572,N_2868);
nor U17870 (N_17870,N_7227,N_6923);
and U17871 (N_17871,N_1692,N_1224);
xor U17872 (N_17872,N_700,N_4292);
and U17873 (N_17873,N_6850,N_7167);
nor U17874 (N_17874,N_4014,N_1604);
and U17875 (N_17875,N_6575,N_3364);
or U17876 (N_17876,N_8637,N_3745);
or U17877 (N_17877,N_2707,N_8381);
xor U17878 (N_17878,N_9537,N_7797);
or U17879 (N_17879,N_8693,N_5688);
nor U17880 (N_17880,N_1607,N_7760);
xor U17881 (N_17881,N_4812,N_2481);
and U17882 (N_17882,N_48,N_9186);
and U17883 (N_17883,N_5232,N_4713);
nand U17884 (N_17884,N_2527,N_8280);
nand U17885 (N_17885,N_3987,N_605);
or U17886 (N_17886,N_232,N_4299);
xor U17887 (N_17887,N_9278,N_1284);
nor U17888 (N_17888,N_933,N_9378);
or U17889 (N_17889,N_1348,N_4227);
xor U17890 (N_17890,N_7847,N_9488);
nand U17891 (N_17891,N_2210,N_1449);
xor U17892 (N_17892,N_8675,N_1122);
nor U17893 (N_17893,N_9297,N_3862);
nand U17894 (N_17894,N_151,N_7942);
nor U17895 (N_17895,N_3781,N_3794);
or U17896 (N_17896,N_4376,N_346);
nor U17897 (N_17897,N_3566,N_5694);
or U17898 (N_17898,N_3957,N_9759);
nor U17899 (N_17899,N_2584,N_4037);
and U17900 (N_17900,N_228,N_4352);
xor U17901 (N_17901,N_8339,N_3242);
and U17902 (N_17902,N_8236,N_4391);
nor U17903 (N_17903,N_6679,N_342);
and U17904 (N_17904,N_4331,N_3736);
or U17905 (N_17905,N_2613,N_3632);
nand U17906 (N_17906,N_2130,N_6707);
xor U17907 (N_17907,N_6958,N_294);
and U17908 (N_17908,N_6486,N_2986);
or U17909 (N_17909,N_6759,N_9670);
xor U17910 (N_17910,N_9294,N_7802);
nor U17911 (N_17911,N_2726,N_6272);
and U17912 (N_17912,N_4370,N_6216);
nor U17913 (N_17913,N_4757,N_6442);
nor U17914 (N_17914,N_7728,N_8497);
nor U17915 (N_17915,N_2552,N_3622);
nand U17916 (N_17916,N_5352,N_9107);
xnor U17917 (N_17917,N_1363,N_1487);
nand U17918 (N_17918,N_5082,N_51);
and U17919 (N_17919,N_619,N_2595);
nand U17920 (N_17920,N_1886,N_4306);
nand U17921 (N_17921,N_7319,N_1444);
and U17922 (N_17922,N_4610,N_634);
and U17923 (N_17923,N_9888,N_9579);
nor U17924 (N_17924,N_6810,N_6509);
or U17925 (N_17925,N_7454,N_3568);
nor U17926 (N_17926,N_9791,N_5757);
nand U17927 (N_17927,N_3392,N_7845);
or U17928 (N_17928,N_5038,N_7888);
and U17929 (N_17929,N_1698,N_1554);
nand U17930 (N_17930,N_6371,N_8398);
and U17931 (N_17931,N_6114,N_1203);
or U17932 (N_17932,N_1461,N_4258);
xnor U17933 (N_17933,N_4965,N_5882);
nand U17934 (N_17934,N_4672,N_4942);
nand U17935 (N_17935,N_2981,N_9588);
xor U17936 (N_17936,N_6253,N_5777);
nand U17937 (N_17937,N_652,N_8788);
nor U17938 (N_17938,N_141,N_5629);
or U17939 (N_17939,N_6001,N_247);
nand U17940 (N_17940,N_1052,N_1298);
or U17941 (N_17941,N_3605,N_7042);
and U17942 (N_17942,N_5101,N_4073);
and U17943 (N_17943,N_672,N_1239);
or U17944 (N_17944,N_7474,N_3384);
and U17945 (N_17945,N_8851,N_6800);
nor U17946 (N_17946,N_6325,N_3793);
xor U17947 (N_17947,N_1910,N_9746);
xnor U17948 (N_17948,N_9144,N_3404);
and U17949 (N_17949,N_3454,N_6758);
nand U17950 (N_17950,N_9497,N_7032);
nand U17951 (N_17951,N_7945,N_122);
and U17952 (N_17952,N_2650,N_5529);
or U17953 (N_17953,N_1071,N_6446);
xor U17954 (N_17954,N_8662,N_8840);
nor U17955 (N_17955,N_422,N_2496);
and U17956 (N_17956,N_2578,N_6675);
and U17957 (N_17957,N_2160,N_6054);
xnor U17958 (N_17958,N_8916,N_2426);
xor U17959 (N_17959,N_8035,N_2442);
xor U17960 (N_17960,N_620,N_7523);
and U17961 (N_17961,N_2677,N_8601);
xnor U17962 (N_17962,N_9152,N_3620);
or U17963 (N_17963,N_9720,N_9705);
or U17964 (N_17964,N_7089,N_4816);
xnor U17965 (N_17965,N_4086,N_6461);
or U17966 (N_17966,N_7542,N_5208);
nand U17967 (N_17967,N_560,N_3913);
and U17968 (N_17968,N_9964,N_7735);
nand U17969 (N_17969,N_375,N_519);
nor U17970 (N_17970,N_6555,N_9462);
and U17971 (N_17971,N_9186,N_9976);
nand U17972 (N_17972,N_4882,N_7986);
and U17973 (N_17973,N_71,N_6075);
xnor U17974 (N_17974,N_3304,N_7884);
nand U17975 (N_17975,N_2835,N_4353);
xor U17976 (N_17976,N_5635,N_3681);
xnor U17977 (N_17977,N_7490,N_2063);
nor U17978 (N_17978,N_5660,N_281);
or U17979 (N_17979,N_880,N_5307);
xor U17980 (N_17980,N_6171,N_8347);
and U17981 (N_17981,N_2022,N_6973);
or U17982 (N_17982,N_7141,N_322);
nor U17983 (N_17983,N_9747,N_9338);
nand U17984 (N_17984,N_5690,N_8729);
nor U17985 (N_17985,N_1487,N_285);
or U17986 (N_17986,N_3097,N_5282);
or U17987 (N_17987,N_8689,N_2688);
and U17988 (N_17988,N_4958,N_4021);
and U17989 (N_17989,N_1991,N_6667);
nor U17990 (N_17990,N_1298,N_4751);
xnor U17991 (N_17991,N_3956,N_8302);
nor U17992 (N_17992,N_9434,N_3631);
xor U17993 (N_17993,N_430,N_7484);
or U17994 (N_17994,N_2609,N_7493);
nor U17995 (N_17995,N_9105,N_38);
nor U17996 (N_17996,N_1026,N_8132);
nor U17997 (N_17997,N_9968,N_5041);
xor U17998 (N_17998,N_5881,N_1992);
nor U17999 (N_17999,N_3755,N_5176);
xnor U18000 (N_18000,N_4561,N_956);
xor U18001 (N_18001,N_1064,N_1281);
nand U18002 (N_18002,N_6540,N_1612);
xor U18003 (N_18003,N_8880,N_1100);
nand U18004 (N_18004,N_8179,N_2558);
nand U18005 (N_18005,N_52,N_2297);
nand U18006 (N_18006,N_3504,N_7728);
nor U18007 (N_18007,N_3234,N_3117);
nor U18008 (N_18008,N_1526,N_8947);
xnor U18009 (N_18009,N_1477,N_3098);
nor U18010 (N_18010,N_2717,N_1844);
nor U18011 (N_18011,N_4714,N_6503);
nor U18012 (N_18012,N_19,N_4933);
nand U18013 (N_18013,N_1489,N_8632);
nand U18014 (N_18014,N_7396,N_8060);
nand U18015 (N_18015,N_8398,N_3777);
and U18016 (N_18016,N_5965,N_8728);
or U18017 (N_18017,N_8608,N_3035);
or U18018 (N_18018,N_5180,N_2170);
xnor U18019 (N_18019,N_311,N_5251);
and U18020 (N_18020,N_1214,N_3160);
nand U18021 (N_18021,N_8064,N_7155);
and U18022 (N_18022,N_3430,N_8888);
nor U18023 (N_18023,N_7875,N_2930);
nand U18024 (N_18024,N_7862,N_85);
nor U18025 (N_18025,N_8594,N_5922);
or U18026 (N_18026,N_984,N_1936);
nor U18027 (N_18027,N_4715,N_4397);
or U18028 (N_18028,N_399,N_3381);
nor U18029 (N_18029,N_6079,N_8573);
or U18030 (N_18030,N_9288,N_8852);
or U18031 (N_18031,N_2318,N_2692);
or U18032 (N_18032,N_4258,N_7219);
nor U18033 (N_18033,N_3358,N_5715);
xnor U18034 (N_18034,N_3244,N_9088);
nor U18035 (N_18035,N_6840,N_1852);
and U18036 (N_18036,N_4106,N_5354);
nor U18037 (N_18037,N_6875,N_2529);
or U18038 (N_18038,N_4649,N_2119);
nand U18039 (N_18039,N_1170,N_8467);
nor U18040 (N_18040,N_3185,N_8066);
or U18041 (N_18041,N_3462,N_1684);
nand U18042 (N_18042,N_2366,N_892);
nor U18043 (N_18043,N_8700,N_515);
and U18044 (N_18044,N_798,N_9225);
and U18045 (N_18045,N_9914,N_845);
nor U18046 (N_18046,N_5859,N_3989);
nand U18047 (N_18047,N_832,N_783);
nor U18048 (N_18048,N_4001,N_9980);
xnor U18049 (N_18049,N_4956,N_2555);
or U18050 (N_18050,N_1481,N_4133);
nor U18051 (N_18051,N_1362,N_4425);
nor U18052 (N_18052,N_8732,N_1042);
and U18053 (N_18053,N_4478,N_6443);
or U18054 (N_18054,N_8977,N_3045);
xor U18055 (N_18055,N_9228,N_9384);
nand U18056 (N_18056,N_4409,N_7693);
and U18057 (N_18057,N_5075,N_5006);
xor U18058 (N_18058,N_2389,N_264);
nor U18059 (N_18059,N_1071,N_8298);
and U18060 (N_18060,N_6818,N_7823);
xnor U18061 (N_18061,N_6552,N_8647);
xor U18062 (N_18062,N_8510,N_4426);
and U18063 (N_18063,N_7520,N_5112);
and U18064 (N_18064,N_4596,N_7991);
nand U18065 (N_18065,N_2532,N_7868);
nor U18066 (N_18066,N_5155,N_3568);
or U18067 (N_18067,N_9579,N_4386);
xor U18068 (N_18068,N_5224,N_5966);
nor U18069 (N_18069,N_165,N_6120);
nor U18070 (N_18070,N_8015,N_9140);
or U18071 (N_18071,N_9498,N_3972);
nand U18072 (N_18072,N_1829,N_6497);
and U18073 (N_18073,N_533,N_163);
xor U18074 (N_18074,N_1206,N_7839);
nand U18075 (N_18075,N_2363,N_7143);
nor U18076 (N_18076,N_8398,N_4767);
nand U18077 (N_18077,N_7725,N_7799);
nor U18078 (N_18078,N_6499,N_2668);
nor U18079 (N_18079,N_3376,N_5467);
or U18080 (N_18080,N_7402,N_5099);
nand U18081 (N_18081,N_1187,N_8508);
xor U18082 (N_18082,N_2364,N_8610);
and U18083 (N_18083,N_1666,N_5048);
or U18084 (N_18084,N_7072,N_2451);
nor U18085 (N_18085,N_5446,N_3775);
and U18086 (N_18086,N_987,N_9880);
nor U18087 (N_18087,N_714,N_9341);
xor U18088 (N_18088,N_3787,N_6474);
and U18089 (N_18089,N_7788,N_1293);
or U18090 (N_18090,N_7438,N_2931);
and U18091 (N_18091,N_9978,N_5333);
or U18092 (N_18092,N_9416,N_3374);
xor U18093 (N_18093,N_8058,N_9322);
and U18094 (N_18094,N_2865,N_2675);
or U18095 (N_18095,N_5843,N_2111);
or U18096 (N_18096,N_8711,N_8797);
and U18097 (N_18097,N_465,N_803);
nor U18098 (N_18098,N_7736,N_4389);
xor U18099 (N_18099,N_7894,N_6842);
or U18100 (N_18100,N_2175,N_6425);
nor U18101 (N_18101,N_338,N_7736);
and U18102 (N_18102,N_1460,N_6362);
and U18103 (N_18103,N_5173,N_5441);
xnor U18104 (N_18104,N_5582,N_9903);
or U18105 (N_18105,N_1301,N_1816);
nand U18106 (N_18106,N_9295,N_2988);
nor U18107 (N_18107,N_9516,N_5293);
nor U18108 (N_18108,N_1567,N_7443);
and U18109 (N_18109,N_7557,N_7003);
xor U18110 (N_18110,N_7760,N_2428);
or U18111 (N_18111,N_7374,N_2321);
and U18112 (N_18112,N_7092,N_6704);
and U18113 (N_18113,N_2659,N_8913);
xor U18114 (N_18114,N_4567,N_744);
or U18115 (N_18115,N_9381,N_5066);
and U18116 (N_18116,N_7824,N_7287);
nand U18117 (N_18117,N_1299,N_5027);
or U18118 (N_18118,N_9328,N_5686);
and U18119 (N_18119,N_5813,N_5741);
or U18120 (N_18120,N_4424,N_6595);
nand U18121 (N_18121,N_4109,N_4790);
or U18122 (N_18122,N_661,N_6910);
nand U18123 (N_18123,N_5968,N_6990);
and U18124 (N_18124,N_6321,N_8405);
nor U18125 (N_18125,N_7751,N_2515);
nand U18126 (N_18126,N_5987,N_9665);
or U18127 (N_18127,N_5013,N_8338);
nor U18128 (N_18128,N_350,N_9961);
and U18129 (N_18129,N_2322,N_6707);
and U18130 (N_18130,N_3186,N_8757);
nand U18131 (N_18131,N_7918,N_5653);
nor U18132 (N_18132,N_8866,N_3779);
xnor U18133 (N_18133,N_2752,N_6213);
xor U18134 (N_18134,N_7144,N_8376);
xor U18135 (N_18135,N_4343,N_2375);
and U18136 (N_18136,N_5944,N_257);
and U18137 (N_18137,N_8158,N_625);
or U18138 (N_18138,N_864,N_5096);
nor U18139 (N_18139,N_8165,N_1229);
nor U18140 (N_18140,N_7093,N_9970);
nand U18141 (N_18141,N_2713,N_7285);
nor U18142 (N_18142,N_7734,N_5601);
nand U18143 (N_18143,N_1477,N_8732);
nand U18144 (N_18144,N_2364,N_7613);
nand U18145 (N_18145,N_1587,N_5562);
nor U18146 (N_18146,N_9660,N_3023);
nor U18147 (N_18147,N_5110,N_7008);
nor U18148 (N_18148,N_2986,N_8258);
nand U18149 (N_18149,N_6870,N_4539);
nand U18150 (N_18150,N_2628,N_5827);
nand U18151 (N_18151,N_3150,N_3291);
nand U18152 (N_18152,N_2172,N_6631);
xor U18153 (N_18153,N_876,N_4654);
nor U18154 (N_18154,N_3301,N_7861);
or U18155 (N_18155,N_1604,N_643);
nand U18156 (N_18156,N_1324,N_1310);
or U18157 (N_18157,N_5307,N_5632);
nor U18158 (N_18158,N_7427,N_4688);
nor U18159 (N_18159,N_36,N_1194);
or U18160 (N_18160,N_763,N_8401);
nand U18161 (N_18161,N_9192,N_5721);
and U18162 (N_18162,N_1408,N_3899);
or U18163 (N_18163,N_7855,N_3991);
nand U18164 (N_18164,N_9771,N_4071);
nand U18165 (N_18165,N_1124,N_1379);
or U18166 (N_18166,N_9416,N_6095);
nor U18167 (N_18167,N_1581,N_9493);
and U18168 (N_18168,N_4541,N_1855);
xor U18169 (N_18169,N_9084,N_1335);
xnor U18170 (N_18170,N_9818,N_9578);
or U18171 (N_18171,N_8915,N_8546);
xor U18172 (N_18172,N_592,N_7189);
and U18173 (N_18173,N_8217,N_6177);
and U18174 (N_18174,N_1780,N_2656);
and U18175 (N_18175,N_928,N_9906);
nor U18176 (N_18176,N_871,N_4401);
and U18177 (N_18177,N_202,N_2105);
nor U18178 (N_18178,N_533,N_2601);
xnor U18179 (N_18179,N_2619,N_8695);
or U18180 (N_18180,N_7594,N_4756);
and U18181 (N_18181,N_7201,N_1122);
xor U18182 (N_18182,N_7890,N_555);
xnor U18183 (N_18183,N_5393,N_7835);
and U18184 (N_18184,N_4199,N_7533);
and U18185 (N_18185,N_4838,N_4461);
nor U18186 (N_18186,N_1795,N_3525);
and U18187 (N_18187,N_8979,N_6603);
xnor U18188 (N_18188,N_2533,N_4007);
or U18189 (N_18189,N_2611,N_2879);
nand U18190 (N_18190,N_3776,N_4836);
and U18191 (N_18191,N_525,N_1347);
or U18192 (N_18192,N_2152,N_8640);
and U18193 (N_18193,N_7015,N_9706);
xnor U18194 (N_18194,N_7117,N_7339);
or U18195 (N_18195,N_6371,N_3692);
and U18196 (N_18196,N_6642,N_250);
nor U18197 (N_18197,N_8161,N_4793);
nor U18198 (N_18198,N_8499,N_2470);
or U18199 (N_18199,N_7867,N_3407);
nor U18200 (N_18200,N_2493,N_9122);
and U18201 (N_18201,N_5613,N_5208);
nor U18202 (N_18202,N_9483,N_7310);
nor U18203 (N_18203,N_4710,N_8668);
and U18204 (N_18204,N_5052,N_4607);
xnor U18205 (N_18205,N_890,N_9962);
xor U18206 (N_18206,N_4247,N_5010);
nand U18207 (N_18207,N_5205,N_2301);
nand U18208 (N_18208,N_1662,N_5992);
nand U18209 (N_18209,N_7730,N_4355);
nor U18210 (N_18210,N_2033,N_8264);
nand U18211 (N_18211,N_5836,N_1332);
or U18212 (N_18212,N_8509,N_3273);
xnor U18213 (N_18213,N_7786,N_8329);
or U18214 (N_18214,N_8126,N_201);
nand U18215 (N_18215,N_2086,N_7887);
nand U18216 (N_18216,N_9530,N_8511);
nor U18217 (N_18217,N_8506,N_6508);
nand U18218 (N_18218,N_7584,N_1385);
nor U18219 (N_18219,N_4541,N_9938);
nor U18220 (N_18220,N_9809,N_2840);
xor U18221 (N_18221,N_2708,N_8256);
and U18222 (N_18222,N_5867,N_3798);
xnor U18223 (N_18223,N_5962,N_7693);
xor U18224 (N_18224,N_5100,N_8734);
and U18225 (N_18225,N_8714,N_2432);
nor U18226 (N_18226,N_1522,N_1569);
and U18227 (N_18227,N_1837,N_8030);
nor U18228 (N_18228,N_1974,N_6316);
xnor U18229 (N_18229,N_1643,N_5997);
nand U18230 (N_18230,N_2449,N_2724);
nand U18231 (N_18231,N_4777,N_3946);
and U18232 (N_18232,N_7789,N_1043);
nand U18233 (N_18233,N_8366,N_243);
xnor U18234 (N_18234,N_3408,N_3527);
and U18235 (N_18235,N_15,N_393);
or U18236 (N_18236,N_8251,N_9478);
or U18237 (N_18237,N_5185,N_457);
nor U18238 (N_18238,N_78,N_6057);
or U18239 (N_18239,N_6973,N_7688);
xor U18240 (N_18240,N_5630,N_9396);
nor U18241 (N_18241,N_3883,N_6957);
xor U18242 (N_18242,N_5687,N_6523);
or U18243 (N_18243,N_5486,N_9734);
nand U18244 (N_18244,N_8789,N_3827);
nand U18245 (N_18245,N_8407,N_2105);
or U18246 (N_18246,N_144,N_4102);
or U18247 (N_18247,N_6639,N_52);
xor U18248 (N_18248,N_9041,N_1373);
xnor U18249 (N_18249,N_5401,N_8127);
nor U18250 (N_18250,N_6273,N_1081);
or U18251 (N_18251,N_3572,N_3289);
nor U18252 (N_18252,N_914,N_1969);
xor U18253 (N_18253,N_6164,N_2980);
nor U18254 (N_18254,N_5286,N_317);
nand U18255 (N_18255,N_3043,N_7615);
or U18256 (N_18256,N_1104,N_7658);
nand U18257 (N_18257,N_7870,N_325);
or U18258 (N_18258,N_4259,N_1649);
xor U18259 (N_18259,N_5644,N_6036);
nor U18260 (N_18260,N_2946,N_9578);
nand U18261 (N_18261,N_460,N_72);
or U18262 (N_18262,N_5077,N_3279);
nand U18263 (N_18263,N_6091,N_1876);
nand U18264 (N_18264,N_659,N_3936);
nor U18265 (N_18265,N_1956,N_2857);
nand U18266 (N_18266,N_4704,N_7454);
and U18267 (N_18267,N_4254,N_985);
nand U18268 (N_18268,N_1209,N_9834);
and U18269 (N_18269,N_5382,N_237);
nand U18270 (N_18270,N_1778,N_2948);
nand U18271 (N_18271,N_8874,N_1758);
nor U18272 (N_18272,N_7490,N_551);
xor U18273 (N_18273,N_9148,N_9638);
and U18274 (N_18274,N_736,N_4947);
nor U18275 (N_18275,N_7254,N_9555);
xor U18276 (N_18276,N_3897,N_7428);
xnor U18277 (N_18277,N_2963,N_6390);
or U18278 (N_18278,N_8867,N_5867);
and U18279 (N_18279,N_3187,N_9696);
or U18280 (N_18280,N_6691,N_4701);
nor U18281 (N_18281,N_472,N_344);
or U18282 (N_18282,N_4930,N_1429);
xnor U18283 (N_18283,N_4825,N_5503);
or U18284 (N_18284,N_4702,N_348);
or U18285 (N_18285,N_2969,N_9524);
nor U18286 (N_18286,N_3870,N_2934);
xnor U18287 (N_18287,N_7484,N_9793);
xor U18288 (N_18288,N_4618,N_3066);
nor U18289 (N_18289,N_3152,N_496);
xor U18290 (N_18290,N_5884,N_8460);
xor U18291 (N_18291,N_866,N_17);
nor U18292 (N_18292,N_5666,N_4977);
or U18293 (N_18293,N_7222,N_6577);
and U18294 (N_18294,N_3678,N_1075);
and U18295 (N_18295,N_7703,N_2781);
and U18296 (N_18296,N_7178,N_2188);
xor U18297 (N_18297,N_1000,N_1031);
nand U18298 (N_18298,N_8043,N_1062);
nor U18299 (N_18299,N_5281,N_3387);
nor U18300 (N_18300,N_5853,N_2620);
or U18301 (N_18301,N_2764,N_8330);
and U18302 (N_18302,N_5468,N_6504);
xnor U18303 (N_18303,N_1662,N_4286);
nand U18304 (N_18304,N_6544,N_4567);
or U18305 (N_18305,N_3080,N_1153);
and U18306 (N_18306,N_371,N_4193);
nor U18307 (N_18307,N_452,N_4442);
and U18308 (N_18308,N_9519,N_9187);
nor U18309 (N_18309,N_4918,N_3609);
or U18310 (N_18310,N_277,N_3663);
and U18311 (N_18311,N_2893,N_8924);
xnor U18312 (N_18312,N_7039,N_6754);
nor U18313 (N_18313,N_5064,N_4274);
nor U18314 (N_18314,N_5190,N_6390);
nor U18315 (N_18315,N_436,N_8898);
nor U18316 (N_18316,N_2552,N_1372);
xnor U18317 (N_18317,N_6285,N_5698);
or U18318 (N_18318,N_1996,N_8854);
or U18319 (N_18319,N_9850,N_2858);
xor U18320 (N_18320,N_4006,N_5617);
xnor U18321 (N_18321,N_1952,N_8418);
nor U18322 (N_18322,N_9812,N_5178);
or U18323 (N_18323,N_310,N_3164);
nand U18324 (N_18324,N_864,N_8753);
nor U18325 (N_18325,N_6235,N_9254);
and U18326 (N_18326,N_9054,N_533);
and U18327 (N_18327,N_5059,N_2302);
nor U18328 (N_18328,N_4163,N_9716);
nor U18329 (N_18329,N_1439,N_5780);
xor U18330 (N_18330,N_369,N_4569);
nand U18331 (N_18331,N_1697,N_9557);
xnor U18332 (N_18332,N_290,N_4997);
nand U18333 (N_18333,N_4048,N_2891);
and U18334 (N_18334,N_8923,N_4849);
or U18335 (N_18335,N_2359,N_3303);
xor U18336 (N_18336,N_6897,N_465);
or U18337 (N_18337,N_8250,N_5185);
or U18338 (N_18338,N_5582,N_4704);
xnor U18339 (N_18339,N_1260,N_7668);
xnor U18340 (N_18340,N_1202,N_4288);
or U18341 (N_18341,N_6849,N_8938);
nand U18342 (N_18342,N_8419,N_5431);
nor U18343 (N_18343,N_3914,N_7462);
or U18344 (N_18344,N_2611,N_1572);
or U18345 (N_18345,N_9262,N_1319);
xnor U18346 (N_18346,N_1099,N_7117);
or U18347 (N_18347,N_1367,N_6065);
or U18348 (N_18348,N_7472,N_7595);
nand U18349 (N_18349,N_2091,N_8233);
and U18350 (N_18350,N_9742,N_701);
or U18351 (N_18351,N_3219,N_9400);
nand U18352 (N_18352,N_7937,N_8598);
xnor U18353 (N_18353,N_3896,N_8586);
and U18354 (N_18354,N_6053,N_7607);
and U18355 (N_18355,N_1636,N_3202);
nand U18356 (N_18356,N_3550,N_6882);
nor U18357 (N_18357,N_3962,N_9863);
nand U18358 (N_18358,N_9143,N_322);
nand U18359 (N_18359,N_1284,N_4339);
nand U18360 (N_18360,N_283,N_9186);
xor U18361 (N_18361,N_7912,N_7953);
or U18362 (N_18362,N_917,N_5571);
nor U18363 (N_18363,N_4975,N_7636);
xor U18364 (N_18364,N_5082,N_8978);
or U18365 (N_18365,N_8586,N_8649);
nand U18366 (N_18366,N_6324,N_2613);
and U18367 (N_18367,N_7191,N_3735);
or U18368 (N_18368,N_9697,N_1972);
and U18369 (N_18369,N_7732,N_8208);
xnor U18370 (N_18370,N_9580,N_7730);
xor U18371 (N_18371,N_4663,N_2976);
nor U18372 (N_18372,N_507,N_7010);
nand U18373 (N_18373,N_3638,N_9622);
nor U18374 (N_18374,N_9183,N_8653);
and U18375 (N_18375,N_9162,N_7366);
and U18376 (N_18376,N_8945,N_4801);
xnor U18377 (N_18377,N_6800,N_1223);
nand U18378 (N_18378,N_2736,N_6393);
nand U18379 (N_18379,N_777,N_1823);
xor U18380 (N_18380,N_753,N_8076);
and U18381 (N_18381,N_8307,N_5919);
nor U18382 (N_18382,N_2312,N_279);
nand U18383 (N_18383,N_5669,N_3671);
nand U18384 (N_18384,N_2514,N_8094);
xnor U18385 (N_18385,N_9609,N_771);
nor U18386 (N_18386,N_3346,N_3545);
nand U18387 (N_18387,N_4465,N_5183);
and U18388 (N_18388,N_1809,N_1387);
and U18389 (N_18389,N_8213,N_1453);
or U18390 (N_18390,N_4884,N_9236);
xnor U18391 (N_18391,N_3309,N_6114);
nand U18392 (N_18392,N_6507,N_4909);
or U18393 (N_18393,N_8539,N_8360);
and U18394 (N_18394,N_2962,N_2621);
nor U18395 (N_18395,N_2155,N_3261);
and U18396 (N_18396,N_5185,N_1147);
nand U18397 (N_18397,N_2385,N_4122);
or U18398 (N_18398,N_5951,N_6207);
or U18399 (N_18399,N_9193,N_9674);
or U18400 (N_18400,N_7919,N_3340);
and U18401 (N_18401,N_7413,N_7907);
xnor U18402 (N_18402,N_420,N_9630);
nand U18403 (N_18403,N_5021,N_4584);
nand U18404 (N_18404,N_851,N_4817);
or U18405 (N_18405,N_8591,N_7142);
nand U18406 (N_18406,N_5916,N_9214);
nand U18407 (N_18407,N_3504,N_3449);
nand U18408 (N_18408,N_1606,N_4829);
nor U18409 (N_18409,N_6946,N_9689);
or U18410 (N_18410,N_8079,N_5549);
nand U18411 (N_18411,N_6554,N_3103);
xor U18412 (N_18412,N_4936,N_5057);
xor U18413 (N_18413,N_5266,N_4745);
or U18414 (N_18414,N_7280,N_6819);
nand U18415 (N_18415,N_8927,N_9881);
or U18416 (N_18416,N_4452,N_4802);
nor U18417 (N_18417,N_4627,N_9279);
or U18418 (N_18418,N_5869,N_5372);
nor U18419 (N_18419,N_8225,N_414);
nor U18420 (N_18420,N_8488,N_7002);
nand U18421 (N_18421,N_5097,N_5638);
and U18422 (N_18422,N_66,N_8760);
nand U18423 (N_18423,N_3573,N_9669);
nand U18424 (N_18424,N_7080,N_3125);
or U18425 (N_18425,N_3335,N_4034);
or U18426 (N_18426,N_4811,N_7787);
nand U18427 (N_18427,N_883,N_2789);
nor U18428 (N_18428,N_4252,N_2874);
nor U18429 (N_18429,N_3558,N_1634);
nand U18430 (N_18430,N_9454,N_8234);
nand U18431 (N_18431,N_6927,N_2519);
xor U18432 (N_18432,N_3327,N_9281);
or U18433 (N_18433,N_8060,N_1803);
xnor U18434 (N_18434,N_2469,N_9718);
or U18435 (N_18435,N_3097,N_9781);
nor U18436 (N_18436,N_4293,N_829);
nand U18437 (N_18437,N_1308,N_103);
nor U18438 (N_18438,N_8754,N_4785);
nand U18439 (N_18439,N_2807,N_7775);
xor U18440 (N_18440,N_8292,N_2029);
nand U18441 (N_18441,N_3806,N_5224);
nand U18442 (N_18442,N_1419,N_988);
or U18443 (N_18443,N_411,N_6884);
or U18444 (N_18444,N_835,N_3239);
or U18445 (N_18445,N_521,N_9314);
or U18446 (N_18446,N_9157,N_8241);
xor U18447 (N_18447,N_7938,N_3042);
nand U18448 (N_18448,N_1689,N_4995);
xnor U18449 (N_18449,N_6562,N_6362);
xnor U18450 (N_18450,N_4831,N_7217);
and U18451 (N_18451,N_311,N_9915);
xor U18452 (N_18452,N_8769,N_5063);
and U18453 (N_18453,N_9487,N_4879);
and U18454 (N_18454,N_8285,N_6065);
or U18455 (N_18455,N_1883,N_1996);
or U18456 (N_18456,N_8525,N_1682);
nor U18457 (N_18457,N_6977,N_1364);
nor U18458 (N_18458,N_750,N_4989);
and U18459 (N_18459,N_7030,N_3076);
xnor U18460 (N_18460,N_5500,N_3847);
nor U18461 (N_18461,N_9812,N_3943);
xor U18462 (N_18462,N_8402,N_3204);
and U18463 (N_18463,N_8159,N_8040);
nor U18464 (N_18464,N_336,N_6359);
or U18465 (N_18465,N_6714,N_4974);
xnor U18466 (N_18466,N_2666,N_6966);
nand U18467 (N_18467,N_2436,N_9738);
nor U18468 (N_18468,N_6822,N_5712);
nand U18469 (N_18469,N_5484,N_9581);
or U18470 (N_18470,N_6839,N_7111);
or U18471 (N_18471,N_7129,N_1575);
nor U18472 (N_18472,N_4577,N_9472);
nor U18473 (N_18473,N_7191,N_6259);
or U18474 (N_18474,N_9979,N_5921);
xnor U18475 (N_18475,N_4249,N_7540);
or U18476 (N_18476,N_6411,N_4581);
or U18477 (N_18477,N_1993,N_6558);
xor U18478 (N_18478,N_8279,N_2363);
nor U18479 (N_18479,N_2844,N_9036);
nand U18480 (N_18480,N_5125,N_1728);
nand U18481 (N_18481,N_7292,N_6706);
and U18482 (N_18482,N_19,N_2682);
nand U18483 (N_18483,N_1229,N_2387);
xnor U18484 (N_18484,N_119,N_4804);
and U18485 (N_18485,N_1613,N_6103);
nand U18486 (N_18486,N_9392,N_7877);
nor U18487 (N_18487,N_4261,N_6801);
xnor U18488 (N_18488,N_6426,N_7522);
xnor U18489 (N_18489,N_2949,N_7881);
nand U18490 (N_18490,N_3605,N_1693);
or U18491 (N_18491,N_2525,N_8867);
or U18492 (N_18492,N_620,N_9117);
nand U18493 (N_18493,N_7158,N_2435);
and U18494 (N_18494,N_9492,N_6738);
nand U18495 (N_18495,N_1601,N_6477);
nand U18496 (N_18496,N_5608,N_3997);
nor U18497 (N_18497,N_6055,N_778);
or U18498 (N_18498,N_6495,N_8809);
or U18499 (N_18499,N_806,N_589);
xor U18500 (N_18500,N_2249,N_4139);
xnor U18501 (N_18501,N_8137,N_7517);
xor U18502 (N_18502,N_6842,N_6480);
and U18503 (N_18503,N_6711,N_7603);
xnor U18504 (N_18504,N_3573,N_2358);
or U18505 (N_18505,N_3189,N_783);
or U18506 (N_18506,N_89,N_3246);
or U18507 (N_18507,N_5689,N_7407);
xnor U18508 (N_18508,N_5170,N_2907);
or U18509 (N_18509,N_2799,N_3828);
xor U18510 (N_18510,N_7479,N_4221);
nand U18511 (N_18511,N_6918,N_5257);
nor U18512 (N_18512,N_5915,N_6801);
or U18513 (N_18513,N_5487,N_5522);
or U18514 (N_18514,N_607,N_5551);
or U18515 (N_18515,N_3729,N_9333);
nor U18516 (N_18516,N_6081,N_4348);
nor U18517 (N_18517,N_3297,N_5247);
nand U18518 (N_18518,N_5152,N_2492);
nor U18519 (N_18519,N_7820,N_5945);
or U18520 (N_18520,N_8707,N_4833);
nand U18521 (N_18521,N_7145,N_858);
or U18522 (N_18522,N_217,N_2723);
and U18523 (N_18523,N_7767,N_7648);
and U18524 (N_18524,N_6834,N_4349);
nor U18525 (N_18525,N_6491,N_9613);
or U18526 (N_18526,N_4230,N_4162);
nand U18527 (N_18527,N_9094,N_9264);
and U18528 (N_18528,N_9415,N_4138);
nor U18529 (N_18529,N_6556,N_6990);
xor U18530 (N_18530,N_9595,N_5026);
and U18531 (N_18531,N_2506,N_6208);
nor U18532 (N_18532,N_873,N_2072);
nand U18533 (N_18533,N_1653,N_9394);
nor U18534 (N_18534,N_1254,N_2908);
or U18535 (N_18535,N_6946,N_8740);
nand U18536 (N_18536,N_9468,N_9778);
and U18537 (N_18537,N_509,N_5726);
nor U18538 (N_18538,N_9277,N_2970);
or U18539 (N_18539,N_3646,N_3498);
and U18540 (N_18540,N_7928,N_5335);
and U18541 (N_18541,N_9831,N_9884);
nand U18542 (N_18542,N_6243,N_5881);
xor U18543 (N_18543,N_8241,N_1179);
and U18544 (N_18544,N_6169,N_9947);
xor U18545 (N_18545,N_2840,N_9662);
xnor U18546 (N_18546,N_8464,N_7071);
xor U18547 (N_18547,N_3010,N_8312);
and U18548 (N_18548,N_279,N_464);
nor U18549 (N_18549,N_2315,N_6719);
or U18550 (N_18550,N_8579,N_4264);
nand U18551 (N_18551,N_8006,N_8803);
and U18552 (N_18552,N_9523,N_7410);
and U18553 (N_18553,N_1675,N_3169);
nand U18554 (N_18554,N_6156,N_474);
or U18555 (N_18555,N_9564,N_9203);
nor U18556 (N_18556,N_8065,N_1807);
xnor U18557 (N_18557,N_418,N_8494);
and U18558 (N_18558,N_4534,N_5553);
or U18559 (N_18559,N_5497,N_513);
nor U18560 (N_18560,N_845,N_7126);
nor U18561 (N_18561,N_4121,N_8533);
or U18562 (N_18562,N_5702,N_7944);
nor U18563 (N_18563,N_227,N_2747);
nand U18564 (N_18564,N_2195,N_475);
and U18565 (N_18565,N_1544,N_5021);
and U18566 (N_18566,N_5570,N_5320);
or U18567 (N_18567,N_227,N_2277);
xnor U18568 (N_18568,N_8265,N_7664);
nand U18569 (N_18569,N_7097,N_2411);
xnor U18570 (N_18570,N_3659,N_8381);
and U18571 (N_18571,N_980,N_5936);
nand U18572 (N_18572,N_1453,N_9495);
or U18573 (N_18573,N_8061,N_1287);
nor U18574 (N_18574,N_8967,N_7391);
xor U18575 (N_18575,N_6741,N_5484);
nand U18576 (N_18576,N_6012,N_1134);
or U18577 (N_18577,N_2205,N_1444);
nor U18578 (N_18578,N_2502,N_5952);
nand U18579 (N_18579,N_3166,N_8655);
xor U18580 (N_18580,N_7229,N_392);
nor U18581 (N_18581,N_9475,N_7201);
or U18582 (N_18582,N_5666,N_9434);
or U18583 (N_18583,N_7614,N_6114);
and U18584 (N_18584,N_2366,N_1042);
and U18585 (N_18585,N_5668,N_982);
nand U18586 (N_18586,N_4381,N_3624);
nand U18587 (N_18587,N_8001,N_3210);
xor U18588 (N_18588,N_5192,N_3683);
nor U18589 (N_18589,N_1211,N_4429);
and U18590 (N_18590,N_3475,N_5884);
and U18591 (N_18591,N_9727,N_1890);
nand U18592 (N_18592,N_7206,N_79);
or U18593 (N_18593,N_2787,N_6979);
xor U18594 (N_18594,N_7816,N_1329);
nand U18595 (N_18595,N_3834,N_5771);
xnor U18596 (N_18596,N_9895,N_4213);
and U18597 (N_18597,N_9249,N_5569);
nor U18598 (N_18598,N_7574,N_5682);
or U18599 (N_18599,N_4300,N_4900);
and U18600 (N_18600,N_6847,N_1481);
or U18601 (N_18601,N_5670,N_7559);
nand U18602 (N_18602,N_9465,N_8788);
or U18603 (N_18603,N_3406,N_547);
nor U18604 (N_18604,N_5227,N_697);
xor U18605 (N_18605,N_5754,N_1240);
or U18606 (N_18606,N_5008,N_3587);
and U18607 (N_18607,N_7085,N_3986);
and U18608 (N_18608,N_2988,N_6043);
and U18609 (N_18609,N_2969,N_9968);
or U18610 (N_18610,N_3299,N_858);
xor U18611 (N_18611,N_2933,N_7962);
nor U18612 (N_18612,N_8145,N_9497);
nor U18613 (N_18613,N_8036,N_5885);
nor U18614 (N_18614,N_2276,N_6859);
xnor U18615 (N_18615,N_3810,N_8189);
nor U18616 (N_18616,N_9398,N_9304);
nor U18617 (N_18617,N_1225,N_3489);
or U18618 (N_18618,N_6611,N_8262);
or U18619 (N_18619,N_7665,N_5019);
or U18620 (N_18620,N_5230,N_1655);
nor U18621 (N_18621,N_7852,N_444);
or U18622 (N_18622,N_8497,N_1559);
or U18623 (N_18623,N_2399,N_1787);
nor U18624 (N_18624,N_5761,N_5938);
nand U18625 (N_18625,N_2473,N_8879);
nor U18626 (N_18626,N_7402,N_3332);
nand U18627 (N_18627,N_6261,N_8431);
and U18628 (N_18628,N_2822,N_2131);
xnor U18629 (N_18629,N_5371,N_3872);
and U18630 (N_18630,N_4253,N_8796);
nor U18631 (N_18631,N_4450,N_592);
and U18632 (N_18632,N_4349,N_6870);
nor U18633 (N_18633,N_5670,N_1791);
xor U18634 (N_18634,N_6873,N_7086);
nor U18635 (N_18635,N_6488,N_6816);
nor U18636 (N_18636,N_1274,N_4032);
nand U18637 (N_18637,N_4131,N_6079);
nand U18638 (N_18638,N_6382,N_103);
xnor U18639 (N_18639,N_8287,N_2387);
xnor U18640 (N_18640,N_3876,N_150);
or U18641 (N_18641,N_2806,N_710);
nor U18642 (N_18642,N_4656,N_5618);
xor U18643 (N_18643,N_506,N_8475);
xor U18644 (N_18644,N_1159,N_8662);
nand U18645 (N_18645,N_6675,N_4394);
nand U18646 (N_18646,N_9750,N_8077);
and U18647 (N_18647,N_3143,N_236);
or U18648 (N_18648,N_1491,N_3663);
nor U18649 (N_18649,N_1331,N_4459);
nand U18650 (N_18650,N_9244,N_7279);
or U18651 (N_18651,N_313,N_8677);
nand U18652 (N_18652,N_8258,N_8869);
nor U18653 (N_18653,N_7753,N_8839);
and U18654 (N_18654,N_6152,N_7791);
nand U18655 (N_18655,N_1514,N_8825);
xor U18656 (N_18656,N_6809,N_2153);
and U18657 (N_18657,N_7748,N_2219);
nor U18658 (N_18658,N_7449,N_1562);
nand U18659 (N_18659,N_6601,N_8354);
and U18660 (N_18660,N_7585,N_525);
and U18661 (N_18661,N_7332,N_6792);
xnor U18662 (N_18662,N_8845,N_6477);
nor U18663 (N_18663,N_9729,N_9588);
nor U18664 (N_18664,N_3817,N_1498);
xnor U18665 (N_18665,N_6324,N_4753);
nand U18666 (N_18666,N_861,N_1049);
nor U18667 (N_18667,N_4852,N_6858);
nand U18668 (N_18668,N_2407,N_6673);
xnor U18669 (N_18669,N_4648,N_9757);
and U18670 (N_18670,N_8270,N_2165);
xor U18671 (N_18671,N_6724,N_1306);
and U18672 (N_18672,N_8480,N_7534);
nor U18673 (N_18673,N_756,N_1863);
nand U18674 (N_18674,N_7574,N_5030);
nand U18675 (N_18675,N_4114,N_8333);
xor U18676 (N_18676,N_8218,N_7482);
xnor U18677 (N_18677,N_8547,N_3667);
and U18678 (N_18678,N_4292,N_3333);
nor U18679 (N_18679,N_1826,N_9505);
nand U18680 (N_18680,N_3122,N_5455);
xnor U18681 (N_18681,N_7470,N_1982);
and U18682 (N_18682,N_5258,N_717);
and U18683 (N_18683,N_8990,N_2248);
nand U18684 (N_18684,N_4851,N_3451);
xor U18685 (N_18685,N_6570,N_7976);
nor U18686 (N_18686,N_5248,N_4040);
nor U18687 (N_18687,N_6353,N_536);
and U18688 (N_18688,N_6350,N_4259);
and U18689 (N_18689,N_4806,N_7567);
or U18690 (N_18690,N_8136,N_604);
and U18691 (N_18691,N_6156,N_4588);
or U18692 (N_18692,N_5506,N_525);
nand U18693 (N_18693,N_603,N_3802);
nand U18694 (N_18694,N_2556,N_4437);
nor U18695 (N_18695,N_2308,N_3746);
nand U18696 (N_18696,N_7802,N_8729);
or U18697 (N_18697,N_9947,N_2521);
or U18698 (N_18698,N_7810,N_3945);
nand U18699 (N_18699,N_9461,N_5368);
and U18700 (N_18700,N_3974,N_2662);
and U18701 (N_18701,N_6548,N_7872);
and U18702 (N_18702,N_2991,N_6410);
nand U18703 (N_18703,N_2939,N_1065);
nor U18704 (N_18704,N_8275,N_4723);
or U18705 (N_18705,N_961,N_2061);
and U18706 (N_18706,N_3044,N_3252);
nand U18707 (N_18707,N_985,N_6939);
or U18708 (N_18708,N_1586,N_1928);
and U18709 (N_18709,N_7963,N_3833);
xor U18710 (N_18710,N_2729,N_4290);
nor U18711 (N_18711,N_8933,N_4183);
or U18712 (N_18712,N_1563,N_5842);
and U18713 (N_18713,N_1590,N_4810);
nor U18714 (N_18714,N_1928,N_1378);
xnor U18715 (N_18715,N_1071,N_337);
or U18716 (N_18716,N_9299,N_2921);
nor U18717 (N_18717,N_6004,N_5638);
or U18718 (N_18718,N_9562,N_8161);
nor U18719 (N_18719,N_6129,N_2440);
xor U18720 (N_18720,N_9689,N_6956);
nand U18721 (N_18721,N_3111,N_7630);
or U18722 (N_18722,N_6638,N_9994);
xor U18723 (N_18723,N_3376,N_8781);
and U18724 (N_18724,N_1140,N_8341);
and U18725 (N_18725,N_4122,N_1259);
or U18726 (N_18726,N_5464,N_4215);
xor U18727 (N_18727,N_6027,N_9818);
nor U18728 (N_18728,N_5375,N_1404);
nor U18729 (N_18729,N_2805,N_5596);
nor U18730 (N_18730,N_9768,N_2390);
nor U18731 (N_18731,N_2968,N_3706);
nand U18732 (N_18732,N_2557,N_7180);
or U18733 (N_18733,N_5901,N_5131);
or U18734 (N_18734,N_8765,N_8149);
xnor U18735 (N_18735,N_9964,N_2140);
nand U18736 (N_18736,N_1034,N_8847);
xor U18737 (N_18737,N_487,N_7420);
nor U18738 (N_18738,N_8940,N_4897);
and U18739 (N_18739,N_8505,N_8355);
nor U18740 (N_18740,N_4620,N_2744);
nor U18741 (N_18741,N_6284,N_2569);
and U18742 (N_18742,N_2920,N_924);
xor U18743 (N_18743,N_4924,N_3231);
and U18744 (N_18744,N_2898,N_6527);
nand U18745 (N_18745,N_2540,N_1573);
or U18746 (N_18746,N_4725,N_689);
nand U18747 (N_18747,N_7960,N_1573);
xnor U18748 (N_18748,N_4010,N_9115);
xnor U18749 (N_18749,N_9884,N_701);
nand U18750 (N_18750,N_5724,N_9612);
xnor U18751 (N_18751,N_3758,N_8364);
nand U18752 (N_18752,N_8063,N_5291);
nand U18753 (N_18753,N_6078,N_5093);
nand U18754 (N_18754,N_338,N_4253);
nand U18755 (N_18755,N_9259,N_4273);
nand U18756 (N_18756,N_8252,N_9343);
xor U18757 (N_18757,N_9171,N_9338);
xnor U18758 (N_18758,N_9917,N_8187);
nor U18759 (N_18759,N_7316,N_1532);
nor U18760 (N_18760,N_5871,N_4353);
or U18761 (N_18761,N_1492,N_8391);
xnor U18762 (N_18762,N_2681,N_7792);
nand U18763 (N_18763,N_7872,N_7274);
or U18764 (N_18764,N_8552,N_186);
nand U18765 (N_18765,N_2225,N_8361);
or U18766 (N_18766,N_8807,N_5535);
nand U18767 (N_18767,N_4722,N_6970);
and U18768 (N_18768,N_787,N_8144);
or U18769 (N_18769,N_1861,N_7687);
nor U18770 (N_18770,N_6041,N_6005);
nand U18771 (N_18771,N_2844,N_8219);
xor U18772 (N_18772,N_4881,N_9349);
xor U18773 (N_18773,N_7859,N_7646);
nand U18774 (N_18774,N_2835,N_6595);
nand U18775 (N_18775,N_7547,N_3038);
and U18776 (N_18776,N_2312,N_800);
nor U18777 (N_18777,N_8233,N_2548);
and U18778 (N_18778,N_8085,N_3467);
nand U18779 (N_18779,N_1696,N_949);
nor U18780 (N_18780,N_3748,N_9174);
nand U18781 (N_18781,N_9702,N_217);
xnor U18782 (N_18782,N_23,N_1565);
or U18783 (N_18783,N_6310,N_7260);
and U18784 (N_18784,N_4119,N_9770);
or U18785 (N_18785,N_4189,N_1991);
nor U18786 (N_18786,N_5699,N_302);
xnor U18787 (N_18787,N_4174,N_1080);
xnor U18788 (N_18788,N_798,N_3875);
nand U18789 (N_18789,N_3868,N_1553);
xor U18790 (N_18790,N_4252,N_7045);
nor U18791 (N_18791,N_9696,N_5785);
nand U18792 (N_18792,N_3297,N_3009);
or U18793 (N_18793,N_9543,N_2708);
xnor U18794 (N_18794,N_4855,N_5243);
xor U18795 (N_18795,N_9436,N_7069);
nand U18796 (N_18796,N_5028,N_2151);
nor U18797 (N_18797,N_2886,N_4113);
xnor U18798 (N_18798,N_3346,N_4907);
or U18799 (N_18799,N_3139,N_7563);
or U18800 (N_18800,N_5651,N_2711);
xnor U18801 (N_18801,N_2125,N_3654);
nand U18802 (N_18802,N_8597,N_8515);
nand U18803 (N_18803,N_7574,N_3364);
or U18804 (N_18804,N_6332,N_4741);
nor U18805 (N_18805,N_2451,N_5642);
and U18806 (N_18806,N_731,N_6262);
and U18807 (N_18807,N_2633,N_1923);
and U18808 (N_18808,N_2657,N_1368);
xor U18809 (N_18809,N_1623,N_1867);
nand U18810 (N_18810,N_3777,N_2148);
or U18811 (N_18811,N_884,N_7507);
nand U18812 (N_18812,N_4525,N_5036);
and U18813 (N_18813,N_4103,N_5571);
or U18814 (N_18814,N_1206,N_3250);
nor U18815 (N_18815,N_8624,N_2755);
or U18816 (N_18816,N_5875,N_5720);
xnor U18817 (N_18817,N_8195,N_4694);
nor U18818 (N_18818,N_9481,N_284);
xnor U18819 (N_18819,N_5282,N_424);
or U18820 (N_18820,N_26,N_6969);
xnor U18821 (N_18821,N_4476,N_4638);
nand U18822 (N_18822,N_5390,N_2532);
or U18823 (N_18823,N_7273,N_9035);
nand U18824 (N_18824,N_6467,N_2382);
and U18825 (N_18825,N_9512,N_4743);
nand U18826 (N_18826,N_6556,N_133);
nand U18827 (N_18827,N_1628,N_5232);
and U18828 (N_18828,N_9072,N_1606);
nor U18829 (N_18829,N_6946,N_200);
and U18830 (N_18830,N_5738,N_4958);
nor U18831 (N_18831,N_1335,N_2061);
or U18832 (N_18832,N_1964,N_3045);
nand U18833 (N_18833,N_1987,N_8935);
and U18834 (N_18834,N_8870,N_5938);
xnor U18835 (N_18835,N_2636,N_1913);
xnor U18836 (N_18836,N_4060,N_4201);
xnor U18837 (N_18837,N_8782,N_3616);
nand U18838 (N_18838,N_1681,N_3070);
and U18839 (N_18839,N_3897,N_178);
or U18840 (N_18840,N_2560,N_9169);
nand U18841 (N_18841,N_8571,N_9484);
and U18842 (N_18842,N_3076,N_9042);
nand U18843 (N_18843,N_4152,N_1707);
nand U18844 (N_18844,N_1837,N_8707);
and U18845 (N_18845,N_6804,N_3085);
nor U18846 (N_18846,N_6537,N_6964);
nand U18847 (N_18847,N_6234,N_2993);
or U18848 (N_18848,N_5000,N_7691);
nor U18849 (N_18849,N_6678,N_3993);
or U18850 (N_18850,N_6369,N_4482);
nor U18851 (N_18851,N_2072,N_1463);
nand U18852 (N_18852,N_5182,N_6709);
or U18853 (N_18853,N_3417,N_1874);
nor U18854 (N_18854,N_2913,N_4238);
nor U18855 (N_18855,N_540,N_2417);
nand U18856 (N_18856,N_7732,N_9257);
xor U18857 (N_18857,N_1819,N_6638);
nand U18858 (N_18858,N_6475,N_1834);
nor U18859 (N_18859,N_1582,N_4139);
xor U18860 (N_18860,N_5488,N_7249);
or U18861 (N_18861,N_4354,N_9255);
nor U18862 (N_18862,N_3806,N_3550);
or U18863 (N_18863,N_2239,N_3333);
xnor U18864 (N_18864,N_6880,N_3493);
nor U18865 (N_18865,N_54,N_17);
nand U18866 (N_18866,N_6128,N_7925);
nand U18867 (N_18867,N_2917,N_6567);
xnor U18868 (N_18868,N_8161,N_1355);
nand U18869 (N_18869,N_9938,N_1332);
nand U18870 (N_18870,N_7904,N_7335);
nand U18871 (N_18871,N_4882,N_2640);
nor U18872 (N_18872,N_6885,N_8957);
nand U18873 (N_18873,N_4462,N_8085);
nor U18874 (N_18874,N_9247,N_7335);
or U18875 (N_18875,N_4992,N_5149);
and U18876 (N_18876,N_6842,N_468);
nand U18877 (N_18877,N_1117,N_8742);
or U18878 (N_18878,N_4999,N_6658);
and U18879 (N_18879,N_698,N_7402);
and U18880 (N_18880,N_5777,N_4096);
xnor U18881 (N_18881,N_5100,N_6514);
and U18882 (N_18882,N_6724,N_8512);
or U18883 (N_18883,N_8113,N_6987);
and U18884 (N_18884,N_8816,N_6576);
nand U18885 (N_18885,N_6709,N_1144);
nor U18886 (N_18886,N_5922,N_8944);
nor U18887 (N_18887,N_7563,N_7893);
nor U18888 (N_18888,N_7968,N_8632);
xor U18889 (N_18889,N_3544,N_2245);
and U18890 (N_18890,N_1206,N_1261);
and U18891 (N_18891,N_1577,N_3178);
nor U18892 (N_18892,N_5475,N_3733);
and U18893 (N_18893,N_6461,N_6364);
or U18894 (N_18894,N_7581,N_937);
and U18895 (N_18895,N_7974,N_9590);
nor U18896 (N_18896,N_7904,N_5040);
nand U18897 (N_18897,N_6648,N_6222);
nor U18898 (N_18898,N_2274,N_2091);
nand U18899 (N_18899,N_5116,N_5409);
and U18900 (N_18900,N_8675,N_5560);
xnor U18901 (N_18901,N_6839,N_3623);
or U18902 (N_18902,N_3122,N_9618);
xnor U18903 (N_18903,N_9447,N_715);
and U18904 (N_18904,N_5312,N_8341);
xor U18905 (N_18905,N_3480,N_3035);
nor U18906 (N_18906,N_4275,N_9946);
nand U18907 (N_18907,N_6293,N_8466);
xor U18908 (N_18908,N_9701,N_5550);
nand U18909 (N_18909,N_7394,N_2208);
nand U18910 (N_18910,N_5644,N_5472);
xnor U18911 (N_18911,N_6102,N_6735);
and U18912 (N_18912,N_2643,N_43);
nand U18913 (N_18913,N_9339,N_243);
xnor U18914 (N_18914,N_1415,N_680);
xnor U18915 (N_18915,N_4806,N_2676);
nor U18916 (N_18916,N_5711,N_8877);
and U18917 (N_18917,N_6465,N_8416);
nand U18918 (N_18918,N_6405,N_9511);
or U18919 (N_18919,N_3659,N_9637);
xor U18920 (N_18920,N_9981,N_6199);
nor U18921 (N_18921,N_4754,N_501);
nor U18922 (N_18922,N_191,N_3018);
nand U18923 (N_18923,N_3918,N_3988);
xnor U18924 (N_18924,N_5762,N_2145);
nand U18925 (N_18925,N_7501,N_9099);
and U18926 (N_18926,N_6938,N_3748);
xor U18927 (N_18927,N_8706,N_4619);
nor U18928 (N_18928,N_7096,N_4873);
nand U18929 (N_18929,N_6223,N_8027);
nand U18930 (N_18930,N_5908,N_9874);
and U18931 (N_18931,N_7141,N_7341);
xnor U18932 (N_18932,N_6931,N_8869);
and U18933 (N_18933,N_8017,N_3942);
xnor U18934 (N_18934,N_6503,N_693);
nand U18935 (N_18935,N_6195,N_1339);
xnor U18936 (N_18936,N_8081,N_6922);
nand U18937 (N_18937,N_7785,N_315);
nor U18938 (N_18938,N_5051,N_5036);
xor U18939 (N_18939,N_2385,N_2722);
nor U18940 (N_18940,N_7508,N_6784);
nor U18941 (N_18941,N_6819,N_8108);
and U18942 (N_18942,N_754,N_5806);
or U18943 (N_18943,N_7220,N_7895);
and U18944 (N_18944,N_6878,N_1497);
xnor U18945 (N_18945,N_6283,N_6316);
xor U18946 (N_18946,N_4825,N_4470);
nor U18947 (N_18947,N_7216,N_9450);
and U18948 (N_18948,N_9726,N_6476);
and U18949 (N_18949,N_5415,N_3433);
nor U18950 (N_18950,N_4157,N_7296);
xor U18951 (N_18951,N_799,N_875);
nor U18952 (N_18952,N_1117,N_4793);
and U18953 (N_18953,N_7169,N_3920);
nor U18954 (N_18954,N_999,N_3411);
xor U18955 (N_18955,N_9168,N_7568);
nor U18956 (N_18956,N_4046,N_5307);
nor U18957 (N_18957,N_1197,N_5202);
or U18958 (N_18958,N_6767,N_1728);
nand U18959 (N_18959,N_1635,N_1087);
and U18960 (N_18960,N_9386,N_8876);
nor U18961 (N_18961,N_236,N_4336);
nor U18962 (N_18962,N_1400,N_2259);
and U18963 (N_18963,N_9481,N_3698);
nor U18964 (N_18964,N_5256,N_3030);
or U18965 (N_18965,N_2190,N_9364);
nand U18966 (N_18966,N_2702,N_4861);
and U18967 (N_18967,N_5342,N_2576);
nor U18968 (N_18968,N_8584,N_623);
or U18969 (N_18969,N_9310,N_9184);
xor U18970 (N_18970,N_3466,N_6375);
xor U18971 (N_18971,N_2134,N_7327);
and U18972 (N_18972,N_9262,N_4738);
and U18973 (N_18973,N_9007,N_4460);
xor U18974 (N_18974,N_8600,N_7856);
xor U18975 (N_18975,N_8752,N_4748);
and U18976 (N_18976,N_748,N_4371);
or U18977 (N_18977,N_1989,N_9784);
xor U18978 (N_18978,N_2830,N_5750);
nand U18979 (N_18979,N_8099,N_7283);
and U18980 (N_18980,N_3616,N_4271);
xnor U18981 (N_18981,N_8253,N_2013);
xnor U18982 (N_18982,N_2573,N_3131);
nor U18983 (N_18983,N_6648,N_1295);
xnor U18984 (N_18984,N_1443,N_791);
nor U18985 (N_18985,N_7578,N_6816);
nor U18986 (N_18986,N_3154,N_874);
nor U18987 (N_18987,N_2809,N_8739);
nand U18988 (N_18988,N_6019,N_323);
nor U18989 (N_18989,N_8777,N_5594);
xnor U18990 (N_18990,N_1722,N_3736);
or U18991 (N_18991,N_1551,N_2032);
or U18992 (N_18992,N_9619,N_8534);
and U18993 (N_18993,N_6708,N_9821);
nor U18994 (N_18994,N_1470,N_515);
nand U18995 (N_18995,N_7756,N_1344);
or U18996 (N_18996,N_9996,N_287);
nand U18997 (N_18997,N_3490,N_7780);
nand U18998 (N_18998,N_343,N_3070);
or U18999 (N_18999,N_532,N_2731);
nand U19000 (N_19000,N_6575,N_9126);
xnor U19001 (N_19001,N_3188,N_866);
xor U19002 (N_19002,N_5310,N_1113);
or U19003 (N_19003,N_1652,N_1938);
xor U19004 (N_19004,N_1963,N_2044);
or U19005 (N_19005,N_4070,N_3727);
nor U19006 (N_19006,N_5735,N_534);
nand U19007 (N_19007,N_9842,N_3762);
and U19008 (N_19008,N_8953,N_1501);
nand U19009 (N_19009,N_7121,N_9547);
and U19010 (N_19010,N_2625,N_6517);
nor U19011 (N_19011,N_910,N_1980);
nor U19012 (N_19012,N_7735,N_2555);
nor U19013 (N_19013,N_3229,N_3045);
and U19014 (N_19014,N_3993,N_6313);
and U19015 (N_19015,N_6846,N_460);
xnor U19016 (N_19016,N_9157,N_2006);
or U19017 (N_19017,N_8433,N_4733);
nor U19018 (N_19018,N_8680,N_3597);
and U19019 (N_19019,N_6258,N_1272);
nor U19020 (N_19020,N_2724,N_7306);
or U19021 (N_19021,N_5242,N_8232);
xor U19022 (N_19022,N_5578,N_636);
or U19023 (N_19023,N_9335,N_1137);
or U19024 (N_19024,N_2573,N_9637);
and U19025 (N_19025,N_8425,N_2000);
nor U19026 (N_19026,N_9818,N_719);
or U19027 (N_19027,N_7237,N_8480);
or U19028 (N_19028,N_3666,N_1906);
xnor U19029 (N_19029,N_8674,N_4799);
xor U19030 (N_19030,N_7307,N_4975);
or U19031 (N_19031,N_5171,N_9654);
nor U19032 (N_19032,N_7913,N_8863);
or U19033 (N_19033,N_1207,N_6377);
nand U19034 (N_19034,N_9703,N_6146);
nor U19035 (N_19035,N_591,N_2430);
nand U19036 (N_19036,N_3319,N_7309);
nand U19037 (N_19037,N_1924,N_2493);
and U19038 (N_19038,N_8521,N_1998);
and U19039 (N_19039,N_8133,N_8237);
nand U19040 (N_19040,N_8929,N_386);
nand U19041 (N_19041,N_9455,N_5327);
or U19042 (N_19042,N_8729,N_2249);
nor U19043 (N_19043,N_3920,N_8491);
and U19044 (N_19044,N_8606,N_4403);
xor U19045 (N_19045,N_8625,N_3598);
or U19046 (N_19046,N_9505,N_3988);
or U19047 (N_19047,N_6607,N_9873);
nand U19048 (N_19048,N_6802,N_5699);
or U19049 (N_19049,N_9879,N_2090);
nor U19050 (N_19050,N_4128,N_3706);
and U19051 (N_19051,N_3365,N_5827);
or U19052 (N_19052,N_1463,N_3847);
nand U19053 (N_19053,N_2247,N_4638);
nor U19054 (N_19054,N_3222,N_9937);
nand U19055 (N_19055,N_3282,N_6423);
nor U19056 (N_19056,N_8382,N_4091);
and U19057 (N_19057,N_8479,N_2744);
and U19058 (N_19058,N_8908,N_6084);
nor U19059 (N_19059,N_7263,N_1068);
or U19060 (N_19060,N_288,N_6588);
or U19061 (N_19061,N_5371,N_1920);
and U19062 (N_19062,N_7369,N_8942);
nor U19063 (N_19063,N_2754,N_164);
and U19064 (N_19064,N_5532,N_8603);
and U19065 (N_19065,N_2628,N_3281);
nor U19066 (N_19066,N_3736,N_3767);
xnor U19067 (N_19067,N_8840,N_8739);
nor U19068 (N_19068,N_7395,N_4367);
or U19069 (N_19069,N_1161,N_4157);
nand U19070 (N_19070,N_1740,N_6914);
xor U19071 (N_19071,N_5927,N_7266);
nand U19072 (N_19072,N_6230,N_5988);
or U19073 (N_19073,N_6687,N_5786);
nor U19074 (N_19074,N_9103,N_5413);
nor U19075 (N_19075,N_4419,N_7509);
and U19076 (N_19076,N_4089,N_8980);
nor U19077 (N_19077,N_2743,N_2653);
nor U19078 (N_19078,N_3408,N_5222);
nor U19079 (N_19079,N_3196,N_803);
nand U19080 (N_19080,N_4251,N_4043);
or U19081 (N_19081,N_8747,N_9223);
xnor U19082 (N_19082,N_9472,N_113);
nor U19083 (N_19083,N_7648,N_5298);
or U19084 (N_19084,N_609,N_2279);
or U19085 (N_19085,N_1225,N_7685);
xnor U19086 (N_19086,N_7767,N_4342);
nand U19087 (N_19087,N_3487,N_792);
xor U19088 (N_19088,N_494,N_8512);
or U19089 (N_19089,N_3733,N_7500);
nand U19090 (N_19090,N_8106,N_5828);
nand U19091 (N_19091,N_3578,N_5206);
nand U19092 (N_19092,N_3991,N_2513);
and U19093 (N_19093,N_856,N_4684);
nor U19094 (N_19094,N_4757,N_1166);
xnor U19095 (N_19095,N_1021,N_3497);
or U19096 (N_19096,N_2306,N_1171);
or U19097 (N_19097,N_2162,N_3073);
and U19098 (N_19098,N_2435,N_2867);
or U19099 (N_19099,N_3549,N_7528);
xnor U19100 (N_19100,N_3453,N_4967);
nor U19101 (N_19101,N_1818,N_4899);
and U19102 (N_19102,N_9999,N_1086);
xnor U19103 (N_19103,N_9832,N_6108);
and U19104 (N_19104,N_6105,N_6849);
nor U19105 (N_19105,N_3942,N_3245);
nand U19106 (N_19106,N_1974,N_7970);
and U19107 (N_19107,N_5391,N_7013);
nand U19108 (N_19108,N_4007,N_7040);
xor U19109 (N_19109,N_7156,N_9936);
xor U19110 (N_19110,N_3738,N_1615);
or U19111 (N_19111,N_4864,N_2202);
and U19112 (N_19112,N_2210,N_8115);
nand U19113 (N_19113,N_1924,N_2415);
nor U19114 (N_19114,N_8063,N_2996);
and U19115 (N_19115,N_9386,N_957);
and U19116 (N_19116,N_6911,N_3989);
nand U19117 (N_19117,N_9962,N_9764);
and U19118 (N_19118,N_2159,N_240);
nor U19119 (N_19119,N_3794,N_2842);
xnor U19120 (N_19120,N_365,N_3773);
nand U19121 (N_19121,N_6717,N_8360);
or U19122 (N_19122,N_4573,N_5584);
nand U19123 (N_19123,N_9920,N_2875);
nand U19124 (N_19124,N_3496,N_9654);
and U19125 (N_19125,N_5972,N_346);
nor U19126 (N_19126,N_6628,N_6581);
or U19127 (N_19127,N_7774,N_1022);
nor U19128 (N_19128,N_8740,N_5838);
nand U19129 (N_19129,N_3917,N_7782);
xor U19130 (N_19130,N_3314,N_4116);
nor U19131 (N_19131,N_7768,N_8461);
or U19132 (N_19132,N_7321,N_7685);
xnor U19133 (N_19133,N_9290,N_7821);
or U19134 (N_19134,N_3127,N_4600);
xor U19135 (N_19135,N_4460,N_1988);
and U19136 (N_19136,N_7242,N_2629);
nand U19137 (N_19137,N_7881,N_4316);
nand U19138 (N_19138,N_2286,N_6622);
nor U19139 (N_19139,N_2281,N_1375);
and U19140 (N_19140,N_7394,N_6558);
nand U19141 (N_19141,N_1630,N_354);
nor U19142 (N_19142,N_1165,N_9347);
xor U19143 (N_19143,N_562,N_3983);
and U19144 (N_19144,N_9458,N_3778);
xor U19145 (N_19145,N_5392,N_4398);
nor U19146 (N_19146,N_8848,N_7556);
or U19147 (N_19147,N_6729,N_3471);
and U19148 (N_19148,N_8958,N_2322);
xor U19149 (N_19149,N_7302,N_2846);
nand U19150 (N_19150,N_9648,N_7141);
nor U19151 (N_19151,N_2598,N_2030);
and U19152 (N_19152,N_2844,N_9973);
xnor U19153 (N_19153,N_3081,N_3758);
or U19154 (N_19154,N_6305,N_5222);
nand U19155 (N_19155,N_3490,N_4548);
or U19156 (N_19156,N_5894,N_885);
or U19157 (N_19157,N_2002,N_1714);
nand U19158 (N_19158,N_9193,N_8003);
nand U19159 (N_19159,N_8975,N_7654);
or U19160 (N_19160,N_66,N_2067);
or U19161 (N_19161,N_6938,N_4518);
or U19162 (N_19162,N_9263,N_9528);
xnor U19163 (N_19163,N_100,N_1044);
and U19164 (N_19164,N_3970,N_9425);
nand U19165 (N_19165,N_6230,N_3944);
nor U19166 (N_19166,N_621,N_8323);
nand U19167 (N_19167,N_1534,N_2845);
nand U19168 (N_19168,N_5414,N_1453);
nor U19169 (N_19169,N_4801,N_472);
xnor U19170 (N_19170,N_9646,N_7655);
xor U19171 (N_19171,N_2213,N_4873);
nand U19172 (N_19172,N_4211,N_1492);
nand U19173 (N_19173,N_2625,N_7722);
nor U19174 (N_19174,N_7763,N_3561);
and U19175 (N_19175,N_8404,N_8360);
nor U19176 (N_19176,N_8011,N_4015);
xnor U19177 (N_19177,N_1632,N_9418);
nand U19178 (N_19178,N_8614,N_2657);
xnor U19179 (N_19179,N_3372,N_9277);
and U19180 (N_19180,N_365,N_1045);
nor U19181 (N_19181,N_6681,N_7535);
nand U19182 (N_19182,N_16,N_6356);
nand U19183 (N_19183,N_6034,N_4903);
nand U19184 (N_19184,N_8478,N_1343);
and U19185 (N_19185,N_2616,N_641);
nand U19186 (N_19186,N_4900,N_3831);
or U19187 (N_19187,N_8966,N_9265);
and U19188 (N_19188,N_2382,N_619);
xor U19189 (N_19189,N_6980,N_4855);
nor U19190 (N_19190,N_8550,N_2131);
nand U19191 (N_19191,N_5218,N_6528);
xnor U19192 (N_19192,N_2534,N_5160);
or U19193 (N_19193,N_9119,N_8962);
or U19194 (N_19194,N_3854,N_4777);
xnor U19195 (N_19195,N_9020,N_4894);
nand U19196 (N_19196,N_4185,N_3343);
nor U19197 (N_19197,N_7780,N_1703);
xor U19198 (N_19198,N_3383,N_5512);
or U19199 (N_19199,N_211,N_4560);
nor U19200 (N_19200,N_8551,N_346);
nor U19201 (N_19201,N_5887,N_8822);
nor U19202 (N_19202,N_9038,N_8943);
or U19203 (N_19203,N_7769,N_2801);
nand U19204 (N_19204,N_3163,N_804);
nor U19205 (N_19205,N_5775,N_9720);
nor U19206 (N_19206,N_9584,N_4798);
nor U19207 (N_19207,N_4943,N_3462);
and U19208 (N_19208,N_5612,N_6215);
nor U19209 (N_19209,N_9802,N_3499);
nand U19210 (N_19210,N_1697,N_1792);
nor U19211 (N_19211,N_2108,N_6895);
and U19212 (N_19212,N_7926,N_300);
nand U19213 (N_19213,N_3796,N_5988);
nand U19214 (N_19214,N_9090,N_1805);
or U19215 (N_19215,N_3571,N_1611);
or U19216 (N_19216,N_9783,N_8912);
nor U19217 (N_19217,N_215,N_9704);
xor U19218 (N_19218,N_2558,N_8811);
and U19219 (N_19219,N_242,N_3836);
xor U19220 (N_19220,N_1782,N_7544);
and U19221 (N_19221,N_1298,N_8497);
xor U19222 (N_19222,N_5716,N_2761);
and U19223 (N_19223,N_4817,N_8465);
nor U19224 (N_19224,N_5874,N_761);
nor U19225 (N_19225,N_8807,N_4751);
nand U19226 (N_19226,N_5010,N_8831);
and U19227 (N_19227,N_6567,N_3052);
or U19228 (N_19228,N_4467,N_4491);
and U19229 (N_19229,N_4457,N_6711);
nor U19230 (N_19230,N_4932,N_3215);
or U19231 (N_19231,N_6755,N_4520);
xor U19232 (N_19232,N_7774,N_9074);
xor U19233 (N_19233,N_5715,N_8514);
nor U19234 (N_19234,N_760,N_5755);
nor U19235 (N_19235,N_3764,N_8949);
or U19236 (N_19236,N_116,N_6950);
or U19237 (N_19237,N_7595,N_7593);
or U19238 (N_19238,N_3171,N_8556);
and U19239 (N_19239,N_7741,N_7487);
nor U19240 (N_19240,N_3139,N_7682);
or U19241 (N_19241,N_7267,N_1974);
or U19242 (N_19242,N_3906,N_8334);
or U19243 (N_19243,N_7454,N_6654);
nand U19244 (N_19244,N_3457,N_9398);
and U19245 (N_19245,N_4235,N_5478);
nand U19246 (N_19246,N_7536,N_1175);
or U19247 (N_19247,N_6893,N_9956);
nor U19248 (N_19248,N_1443,N_4766);
nand U19249 (N_19249,N_7381,N_6098);
xnor U19250 (N_19250,N_1690,N_8577);
nand U19251 (N_19251,N_4516,N_6706);
xnor U19252 (N_19252,N_4291,N_8694);
nor U19253 (N_19253,N_6118,N_7422);
nor U19254 (N_19254,N_4134,N_2818);
and U19255 (N_19255,N_1334,N_9516);
nand U19256 (N_19256,N_3267,N_4188);
nand U19257 (N_19257,N_8065,N_1269);
xnor U19258 (N_19258,N_7578,N_9411);
or U19259 (N_19259,N_2499,N_4467);
nand U19260 (N_19260,N_2414,N_9077);
xor U19261 (N_19261,N_3145,N_1165);
or U19262 (N_19262,N_4238,N_9837);
and U19263 (N_19263,N_2111,N_4493);
and U19264 (N_19264,N_3681,N_6298);
xor U19265 (N_19265,N_5019,N_6433);
nor U19266 (N_19266,N_2010,N_467);
nor U19267 (N_19267,N_3540,N_8818);
and U19268 (N_19268,N_9135,N_4439);
xor U19269 (N_19269,N_740,N_1738);
and U19270 (N_19270,N_9263,N_9106);
nand U19271 (N_19271,N_1768,N_7491);
and U19272 (N_19272,N_9789,N_5565);
xor U19273 (N_19273,N_5210,N_6234);
nor U19274 (N_19274,N_5213,N_469);
or U19275 (N_19275,N_4266,N_4496);
xnor U19276 (N_19276,N_1559,N_2971);
or U19277 (N_19277,N_3643,N_4659);
xor U19278 (N_19278,N_6908,N_1424);
nor U19279 (N_19279,N_8623,N_4738);
and U19280 (N_19280,N_430,N_8285);
or U19281 (N_19281,N_7795,N_1304);
and U19282 (N_19282,N_7008,N_1179);
nand U19283 (N_19283,N_9733,N_8974);
nor U19284 (N_19284,N_9140,N_7658);
nor U19285 (N_19285,N_7569,N_5278);
nand U19286 (N_19286,N_2668,N_3476);
nor U19287 (N_19287,N_2790,N_81);
and U19288 (N_19288,N_8577,N_6478);
xor U19289 (N_19289,N_1128,N_6760);
and U19290 (N_19290,N_593,N_1636);
xnor U19291 (N_19291,N_7530,N_2651);
nand U19292 (N_19292,N_3284,N_4180);
nor U19293 (N_19293,N_7855,N_8203);
or U19294 (N_19294,N_4194,N_270);
nand U19295 (N_19295,N_4283,N_6636);
nand U19296 (N_19296,N_2429,N_7588);
xor U19297 (N_19297,N_3586,N_2320);
nor U19298 (N_19298,N_5191,N_9017);
or U19299 (N_19299,N_3927,N_1377);
or U19300 (N_19300,N_4313,N_3211);
and U19301 (N_19301,N_1747,N_6976);
nand U19302 (N_19302,N_5979,N_8760);
xor U19303 (N_19303,N_6614,N_4925);
and U19304 (N_19304,N_6656,N_9704);
nor U19305 (N_19305,N_3557,N_4278);
and U19306 (N_19306,N_6162,N_1895);
or U19307 (N_19307,N_5550,N_9655);
nand U19308 (N_19308,N_8023,N_9169);
nand U19309 (N_19309,N_4801,N_8029);
or U19310 (N_19310,N_1582,N_6436);
or U19311 (N_19311,N_6072,N_8690);
and U19312 (N_19312,N_6602,N_7510);
xor U19313 (N_19313,N_2610,N_2800);
or U19314 (N_19314,N_2978,N_4415);
nand U19315 (N_19315,N_5229,N_7237);
and U19316 (N_19316,N_2788,N_6730);
or U19317 (N_19317,N_8777,N_7659);
or U19318 (N_19318,N_1738,N_7865);
or U19319 (N_19319,N_1139,N_874);
xnor U19320 (N_19320,N_300,N_8976);
nor U19321 (N_19321,N_5971,N_406);
nor U19322 (N_19322,N_9383,N_6798);
nand U19323 (N_19323,N_57,N_5024);
nand U19324 (N_19324,N_1273,N_3304);
nand U19325 (N_19325,N_2453,N_8558);
nor U19326 (N_19326,N_1929,N_9276);
nor U19327 (N_19327,N_1686,N_4511);
xor U19328 (N_19328,N_1996,N_6391);
and U19329 (N_19329,N_2258,N_3399);
or U19330 (N_19330,N_842,N_1804);
or U19331 (N_19331,N_3973,N_3260);
and U19332 (N_19332,N_879,N_8274);
or U19333 (N_19333,N_6245,N_449);
nor U19334 (N_19334,N_4958,N_176);
nor U19335 (N_19335,N_5963,N_722);
nand U19336 (N_19336,N_4187,N_8257);
xor U19337 (N_19337,N_7176,N_9007);
or U19338 (N_19338,N_7081,N_3635);
and U19339 (N_19339,N_9063,N_6576);
xnor U19340 (N_19340,N_7270,N_5344);
nor U19341 (N_19341,N_2648,N_9885);
xor U19342 (N_19342,N_3257,N_5305);
or U19343 (N_19343,N_853,N_4747);
nor U19344 (N_19344,N_6324,N_6985);
xor U19345 (N_19345,N_1000,N_1026);
or U19346 (N_19346,N_7591,N_5878);
nand U19347 (N_19347,N_823,N_6516);
or U19348 (N_19348,N_9705,N_399);
or U19349 (N_19349,N_9556,N_2912);
nand U19350 (N_19350,N_5854,N_4365);
or U19351 (N_19351,N_1733,N_4366);
and U19352 (N_19352,N_5383,N_1465);
nand U19353 (N_19353,N_3855,N_4118);
and U19354 (N_19354,N_3220,N_9503);
nand U19355 (N_19355,N_8055,N_239);
nor U19356 (N_19356,N_78,N_826);
xnor U19357 (N_19357,N_2551,N_5946);
and U19358 (N_19358,N_9562,N_8219);
nand U19359 (N_19359,N_6901,N_2309);
or U19360 (N_19360,N_9243,N_3898);
and U19361 (N_19361,N_9231,N_432);
nor U19362 (N_19362,N_7728,N_2473);
xnor U19363 (N_19363,N_3436,N_6982);
xnor U19364 (N_19364,N_6769,N_6416);
nand U19365 (N_19365,N_5718,N_9011);
xnor U19366 (N_19366,N_3444,N_6516);
nor U19367 (N_19367,N_8725,N_4423);
or U19368 (N_19368,N_215,N_1125);
nand U19369 (N_19369,N_1007,N_2827);
and U19370 (N_19370,N_8739,N_4355);
or U19371 (N_19371,N_7166,N_5294);
nand U19372 (N_19372,N_8836,N_9);
nor U19373 (N_19373,N_8080,N_8197);
nand U19374 (N_19374,N_8277,N_8853);
or U19375 (N_19375,N_5408,N_6862);
and U19376 (N_19376,N_6230,N_5709);
or U19377 (N_19377,N_2662,N_9118);
xnor U19378 (N_19378,N_7368,N_751);
xnor U19379 (N_19379,N_7203,N_1111);
and U19380 (N_19380,N_2806,N_2447);
or U19381 (N_19381,N_8189,N_7893);
nand U19382 (N_19382,N_9859,N_9002);
or U19383 (N_19383,N_254,N_4550);
nand U19384 (N_19384,N_8438,N_6528);
and U19385 (N_19385,N_9931,N_3896);
nor U19386 (N_19386,N_2894,N_4036);
nand U19387 (N_19387,N_2967,N_6401);
or U19388 (N_19388,N_6649,N_1580);
nor U19389 (N_19389,N_9553,N_3174);
or U19390 (N_19390,N_7653,N_8736);
nand U19391 (N_19391,N_6259,N_6120);
xor U19392 (N_19392,N_6835,N_5509);
nor U19393 (N_19393,N_1610,N_2080);
nor U19394 (N_19394,N_3115,N_9767);
nand U19395 (N_19395,N_6800,N_9963);
and U19396 (N_19396,N_4161,N_8693);
xnor U19397 (N_19397,N_244,N_7366);
and U19398 (N_19398,N_2950,N_2648);
nor U19399 (N_19399,N_3578,N_6468);
and U19400 (N_19400,N_3714,N_565);
or U19401 (N_19401,N_7905,N_2545);
xor U19402 (N_19402,N_9614,N_697);
nand U19403 (N_19403,N_265,N_7616);
or U19404 (N_19404,N_7655,N_136);
xnor U19405 (N_19405,N_8060,N_3340);
and U19406 (N_19406,N_5533,N_8171);
xor U19407 (N_19407,N_5059,N_2009);
and U19408 (N_19408,N_6664,N_7749);
nand U19409 (N_19409,N_6489,N_772);
and U19410 (N_19410,N_2002,N_7254);
nor U19411 (N_19411,N_9801,N_2008);
nand U19412 (N_19412,N_6558,N_7717);
or U19413 (N_19413,N_7558,N_4400);
xor U19414 (N_19414,N_2743,N_9078);
and U19415 (N_19415,N_7262,N_3441);
and U19416 (N_19416,N_2286,N_9264);
xnor U19417 (N_19417,N_6819,N_2051);
xor U19418 (N_19418,N_3156,N_2262);
or U19419 (N_19419,N_9439,N_7066);
or U19420 (N_19420,N_174,N_4234);
nand U19421 (N_19421,N_8582,N_9191);
xor U19422 (N_19422,N_3759,N_2865);
and U19423 (N_19423,N_6993,N_8984);
and U19424 (N_19424,N_9222,N_9967);
and U19425 (N_19425,N_388,N_9820);
or U19426 (N_19426,N_6117,N_9309);
xnor U19427 (N_19427,N_6267,N_2529);
and U19428 (N_19428,N_5121,N_7389);
and U19429 (N_19429,N_6209,N_863);
and U19430 (N_19430,N_6841,N_4721);
xor U19431 (N_19431,N_6123,N_7236);
nor U19432 (N_19432,N_1316,N_7588);
nor U19433 (N_19433,N_684,N_1586);
and U19434 (N_19434,N_3178,N_9332);
xor U19435 (N_19435,N_4185,N_7151);
nand U19436 (N_19436,N_2382,N_5434);
nor U19437 (N_19437,N_7637,N_4029);
nand U19438 (N_19438,N_5385,N_9192);
and U19439 (N_19439,N_9819,N_8627);
nor U19440 (N_19440,N_8645,N_8214);
and U19441 (N_19441,N_6176,N_7417);
nand U19442 (N_19442,N_5109,N_5048);
nor U19443 (N_19443,N_9895,N_6153);
nor U19444 (N_19444,N_9821,N_9610);
nand U19445 (N_19445,N_8740,N_4004);
nand U19446 (N_19446,N_5928,N_4202);
xnor U19447 (N_19447,N_6096,N_3222);
nand U19448 (N_19448,N_3006,N_9453);
nor U19449 (N_19449,N_1087,N_2261);
nor U19450 (N_19450,N_2189,N_4260);
and U19451 (N_19451,N_256,N_3746);
nor U19452 (N_19452,N_7698,N_6982);
xor U19453 (N_19453,N_6553,N_5651);
and U19454 (N_19454,N_1483,N_2981);
nor U19455 (N_19455,N_4284,N_6536);
and U19456 (N_19456,N_1653,N_237);
xnor U19457 (N_19457,N_2207,N_3574);
and U19458 (N_19458,N_6808,N_3559);
nand U19459 (N_19459,N_2300,N_2007);
nor U19460 (N_19460,N_9301,N_9246);
nand U19461 (N_19461,N_7267,N_8872);
xor U19462 (N_19462,N_5257,N_2318);
xor U19463 (N_19463,N_8785,N_2340);
xor U19464 (N_19464,N_3445,N_3952);
and U19465 (N_19465,N_9339,N_2729);
xnor U19466 (N_19466,N_9547,N_9584);
xnor U19467 (N_19467,N_8051,N_5367);
xnor U19468 (N_19468,N_9262,N_4406);
nor U19469 (N_19469,N_3134,N_2383);
nand U19470 (N_19470,N_205,N_2045);
and U19471 (N_19471,N_2405,N_756);
nor U19472 (N_19472,N_5272,N_8611);
or U19473 (N_19473,N_2500,N_9947);
and U19474 (N_19474,N_9283,N_3539);
xor U19475 (N_19475,N_4915,N_167);
or U19476 (N_19476,N_3674,N_2748);
xor U19477 (N_19477,N_4051,N_5722);
nand U19478 (N_19478,N_5045,N_4523);
nor U19479 (N_19479,N_5974,N_7576);
nand U19480 (N_19480,N_7624,N_4805);
nand U19481 (N_19481,N_8534,N_5557);
nand U19482 (N_19482,N_2716,N_8169);
and U19483 (N_19483,N_3286,N_2267);
xnor U19484 (N_19484,N_2691,N_1823);
nor U19485 (N_19485,N_7815,N_9504);
or U19486 (N_19486,N_3611,N_2628);
or U19487 (N_19487,N_267,N_8557);
xnor U19488 (N_19488,N_9589,N_7645);
or U19489 (N_19489,N_3756,N_1525);
nor U19490 (N_19490,N_3094,N_7391);
nor U19491 (N_19491,N_3924,N_8322);
nor U19492 (N_19492,N_3904,N_6711);
nand U19493 (N_19493,N_9847,N_3707);
nand U19494 (N_19494,N_2401,N_1043);
nor U19495 (N_19495,N_8382,N_7414);
or U19496 (N_19496,N_2929,N_733);
or U19497 (N_19497,N_7529,N_2298);
nor U19498 (N_19498,N_3813,N_260);
xnor U19499 (N_19499,N_202,N_9987);
nor U19500 (N_19500,N_4908,N_158);
nor U19501 (N_19501,N_3171,N_7493);
and U19502 (N_19502,N_6738,N_886);
or U19503 (N_19503,N_4253,N_8169);
nand U19504 (N_19504,N_9432,N_8613);
nor U19505 (N_19505,N_3693,N_6296);
or U19506 (N_19506,N_9620,N_4549);
or U19507 (N_19507,N_9937,N_2765);
xnor U19508 (N_19508,N_3541,N_6186);
nand U19509 (N_19509,N_5268,N_4689);
nor U19510 (N_19510,N_1755,N_3296);
nand U19511 (N_19511,N_183,N_135);
or U19512 (N_19512,N_6072,N_3369);
and U19513 (N_19513,N_4649,N_4612);
xnor U19514 (N_19514,N_3580,N_101);
xnor U19515 (N_19515,N_2603,N_6787);
nor U19516 (N_19516,N_5953,N_5758);
and U19517 (N_19517,N_737,N_4453);
and U19518 (N_19518,N_9027,N_3856);
xnor U19519 (N_19519,N_89,N_5002);
xnor U19520 (N_19520,N_1834,N_2258);
and U19521 (N_19521,N_4758,N_7251);
nand U19522 (N_19522,N_6252,N_7530);
and U19523 (N_19523,N_6376,N_793);
xor U19524 (N_19524,N_4614,N_1667);
nor U19525 (N_19525,N_6037,N_8900);
nand U19526 (N_19526,N_6590,N_2742);
nor U19527 (N_19527,N_1113,N_9615);
nand U19528 (N_19528,N_7289,N_3396);
and U19529 (N_19529,N_9292,N_4594);
and U19530 (N_19530,N_9620,N_8141);
nor U19531 (N_19531,N_5698,N_5459);
nand U19532 (N_19532,N_7001,N_9026);
xnor U19533 (N_19533,N_8403,N_731);
nand U19534 (N_19534,N_7257,N_6550);
nor U19535 (N_19535,N_4327,N_7782);
nand U19536 (N_19536,N_3159,N_2867);
nand U19537 (N_19537,N_8183,N_3780);
nor U19538 (N_19538,N_2159,N_5928);
or U19539 (N_19539,N_3289,N_4647);
nand U19540 (N_19540,N_4051,N_2371);
and U19541 (N_19541,N_9323,N_5899);
nor U19542 (N_19542,N_4308,N_7828);
nor U19543 (N_19543,N_9802,N_6913);
nand U19544 (N_19544,N_1827,N_8532);
and U19545 (N_19545,N_3368,N_3377);
nor U19546 (N_19546,N_5777,N_1946);
nand U19547 (N_19547,N_7252,N_1020);
nor U19548 (N_19548,N_4739,N_3826);
nor U19549 (N_19549,N_2223,N_7062);
and U19550 (N_19550,N_1511,N_8833);
nor U19551 (N_19551,N_3847,N_7871);
nand U19552 (N_19552,N_6067,N_3788);
or U19553 (N_19553,N_1680,N_5474);
nor U19554 (N_19554,N_3955,N_9601);
and U19555 (N_19555,N_1713,N_8450);
nor U19556 (N_19556,N_869,N_9480);
nor U19557 (N_19557,N_6809,N_7123);
and U19558 (N_19558,N_6445,N_4425);
nor U19559 (N_19559,N_3778,N_7300);
xor U19560 (N_19560,N_9975,N_4060);
and U19561 (N_19561,N_3973,N_8230);
nand U19562 (N_19562,N_2885,N_343);
or U19563 (N_19563,N_757,N_7371);
xor U19564 (N_19564,N_7312,N_3505);
or U19565 (N_19565,N_2058,N_6664);
nand U19566 (N_19566,N_4324,N_6187);
nor U19567 (N_19567,N_4,N_1994);
xor U19568 (N_19568,N_9505,N_528);
or U19569 (N_19569,N_5919,N_535);
nor U19570 (N_19570,N_1938,N_6655);
xnor U19571 (N_19571,N_2308,N_3936);
and U19572 (N_19572,N_636,N_1837);
nor U19573 (N_19573,N_7720,N_2911);
nor U19574 (N_19574,N_9006,N_4409);
or U19575 (N_19575,N_9349,N_7428);
nand U19576 (N_19576,N_9713,N_4930);
xnor U19577 (N_19577,N_585,N_4643);
xor U19578 (N_19578,N_7352,N_2987);
nor U19579 (N_19579,N_3309,N_473);
nor U19580 (N_19580,N_8484,N_7449);
xnor U19581 (N_19581,N_5383,N_1492);
nor U19582 (N_19582,N_2140,N_7042);
nand U19583 (N_19583,N_85,N_48);
and U19584 (N_19584,N_4931,N_8626);
nand U19585 (N_19585,N_5285,N_6551);
nand U19586 (N_19586,N_6276,N_6267);
xor U19587 (N_19587,N_8547,N_6209);
xnor U19588 (N_19588,N_2794,N_8198);
nor U19589 (N_19589,N_1095,N_3208);
xor U19590 (N_19590,N_5011,N_5009);
or U19591 (N_19591,N_9463,N_7695);
xnor U19592 (N_19592,N_1996,N_480);
and U19593 (N_19593,N_8912,N_2302);
nor U19594 (N_19594,N_4132,N_3358);
nor U19595 (N_19595,N_6004,N_7581);
xor U19596 (N_19596,N_2815,N_6577);
xnor U19597 (N_19597,N_8953,N_2279);
and U19598 (N_19598,N_43,N_9192);
or U19599 (N_19599,N_9199,N_8755);
nand U19600 (N_19600,N_7907,N_7654);
nor U19601 (N_19601,N_2533,N_8614);
and U19602 (N_19602,N_7505,N_7298);
or U19603 (N_19603,N_1135,N_4739);
xor U19604 (N_19604,N_9618,N_3712);
and U19605 (N_19605,N_5434,N_9872);
or U19606 (N_19606,N_7939,N_9693);
and U19607 (N_19607,N_9892,N_9443);
xor U19608 (N_19608,N_4710,N_1032);
nor U19609 (N_19609,N_2745,N_3640);
and U19610 (N_19610,N_3256,N_3006);
xnor U19611 (N_19611,N_3057,N_6135);
nor U19612 (N_19612,N_7067,N_4884);
nand U19613 (N_19613,N_1534,N_9263);
or U19614 (N_19614,N_7154,N_8834);
nor U19615 (N_19615,N_1345,N_3146);
or U19616 (N_19616,N_9395,N_1902);
nand U19617 (N_19617,N_9156,N_4190);
xor U19618 (N_19618,N_2444,N_4672);
or U19619 (N_19619,N_2455,N_655);
or U19620 (N_19620,N_5482,N_2544);
and U19621 (N_19621,N_6585,N_2849);
nor U19622 (N_19622,N_1817,N_1052);
or U19623 (N_19623,N_8319,N_104);
and U19624 (N_19624,N_6601,N_9397);
and U19625 (N_19625,N_795,N_2775);
xnor U19626 (N_19626,N_5869,N_6692);
xnor U19627 (N_19627,N_9489,N_837);
nor U19628 (N_19628,N_6983,N_3368);
xnor U19629 (N_19629,N_6472,N_7194);
nand U19630 (N_19630,N_7497,N_969);
and U19631 (N_19631,N_1164,N_4840);
xnor U19632 (N_19632,N_2789,N_5511);
and U19633 (N_19633,N_8551,N_9073);
nand U19634 (N_19634,N_2676,N_9921);
nor U19635 (N_19635,N_8273,N_1742);
or U19636 (N_19636,N_7478,N_5831);
or U19637 (N_19637,N_9226,N_6670);
xnor U19638 (N_19638,N_7351,N_9128);
nor U19639 (N_19639,N_9978,N_4371);
and U19640 (N_19640,N_3839,N_9944);
nand U19641 (N_19641,N_2258,N_8991);
xor U19642 (N_19642,N_5309,N_6161);
nor U19643 (N_19643,N_1154,N_5699);
xnor U19644 (N_19644,N_4701,N_5633);
xnor U19645 (N_19645,N_6022,N_2884);
nor U19646 (N_19646,N_5628,N_9812);
and U19647 (N_19647,N_2171,N_7426);
and U19648 (N_19648,N_2321,N_1166);
nor U19649 (N_19649,N_9304,N_7393);
xor U19650 (N_19650,N_8842,N_3442);
xnor U19651 (N_19651,N_5765,N_4972);
or U19652 (N_19652,N_1538,N_2181);
nand U19653 (N_19653,N_8719,N_8116);
nand U19654 (N_19654,N_4895,N_4413);
xnor U19655 (N_19655,N_2988,N_7346);
or U19656 (N_19656,N_2027,N_3493);
or U19657 (N_19657,N_4337,N_1287);
nand U19658 (N_19658,N_4568,N_2364);
or U19659 (N_19659,N_3529,N_2251);
xnor U19660 (N_19660,N_7788,N_9270);
nor U19661 (N_19661,N_8700,N_5419);
nand U19662 (N_19662,N_143,N_641);
nand U19663 (N_19663,N_6582,N_7301);
or U19664 (N_19664,N_5578,N_1112);
nor U19665 (N_19665,N_7737,N_3568);
nand U19666 (N_19666,N_2314,N_2890);
xnor U19667 (N_19667,N_7117,N_9311);
or U19668 (N_19668,N_1504,N_3603);
nor U19669 (N_19669,N_424,N_9560);
nand U19670 (N_19670,N_4826,N_8320);
or U19671 (N_19671,N_4739,N_6560);
or U19672 (N_19672,N_4890,N_1082);
xnor U19673 (N_19673,N_6469,N_5901);
or U19674 (N_19674,N_30,N_2413);
and U19675 (N_19675,N_5510,N_7710);
nor U19676 (N_19676,N_8341,N_6358);
xor U19677 (N_19677,N_8138,N_5098);
nand U19678 (N_19678,N_9791,N_8170);
or U19679 (N_19679,N_6370,N_1387);
and U19680 (N_19680,N_3063,N_1729);
nor U19681 (N_19681,N_4500,N_523);
nor U19682 (N_19682,N_2057,N_3062);
and U19683 (N_19683,N_7627,N_343);
nor U19684 (N_19684,N_7651,N_5424);
nand U19685 (N_19685,N_5157,N_9478);
xnor U19686 (N_19686,N_3666,N_2637);
nor U19687 (N_19687,N_6534,N_7713);
xnor U19688 (N_19688,N_8098,N_7624);
or U19689 (N_19689,N_7506,N_6930);
or U19690 (N_19690,N_5289,N_654);
xnor U19691 (N_19691,N_5687,N_4852);
nor U19692 (N_19692,N_8088,N_7658);
or U19693 (N_19693,N_2398,N_1772);
xor U19694 (N_19694,N_1911,N_8723);
nand U19695 (N_19695,N_1543,N_3277);
and U19696 (N_19696,N_4966,N_725);
nor U19697 (N_19697,N_5661,N_7438);
and U19698 (N_19698,N_3392,N_270);
nor U19699 (N_19699,N_5670,N_2773);
nor U19700 (N_19700,N_5630,N_9771);
nand U19701 (N_19701,N_274,N_5021);
nand U19702 (N_19702,N_5270,N_6964);
nand U19703 (N_19703,N_5898,N_7694);
nor U19704 (N_19704,N_7562,N_597);
or U19705 (N_19705,N_7966,N_6119);
nand U19706 (N_19706,N_1613,N_3372);
or U19707 (N_19707,N_1165,N_5758);
and U19708 (N_19708,N_7828,N_6728);
and U19709 (N_19709,N_1829,N_8130);
and U19710 (N_19710,N_5698,N_4608);
nand U19711 (N_19711,N_189,N_4647);
and U19712 (N_19712,N_414,N_9103);
nor U19713 (N_19713,N_8365,N_3218);
nor U19714 (N_19714,N_1177,N_4106);
or U19715 (N_19715,N_8279,N_2051);
nor U19716 (N_19716,N_9789,N_9409);
nor U19717 (N_19717,N_910,N_1467);
or U19718 (N_19718,N_7522,N_2205);
or U19719 (N_19719,N_3950,N_9609);
nand U19720 (N_19720,N_4491,N_1551);
xor U19721 (N_19721,N_1317,N_2771);
xor U19722 (N_19722,N_9359,N_2476);
and U19723 (N_19723,N_292,N_8936);
and U19724 (N_19724,N_1243,N_4657);
nand U19725 (N_19725,N_1183,N_4381);
or U19726 (N_19726,N_2904,N_7713);
or U19727 (N_19727,N_6052,N_6720);
or U19728 (N_19728,N_5852,N_2478);
xor U19729 (N_19729,N_4543,N_3442);
or U19730 (N_19730,N_767,N_9954);
nand U19731 (N_19731,N_8302,N_6455);
xor U19732 (N_19732,N_574,N_5864);
nor U19733 (N_19733,N_9558,N_9820);
or U19734 (N_19734,N_1525,N_2237);
and U19735 (N_19735,N_633,N_7460);
or U19736 (N_19736,N_6064,N_1989);
xor U19737 (N_19737,N_5794,N_3045);
nor U19738 (N_19738,N_1585,N_8088);
and U19739 (N_19739,N_2318,N_6681);
xnor U19740 (N_19740,N_1410,N_8070);
xor U19741 (N_19741,N_7881,N_2862);
and U19742 (N_19742,N_3095,N_7969);
and U19743 (N_19743,N_7858,N_1074);
xnor U19744 (N_19744,N_8804,N_9664);
and U19745 (N_19745,N_630,N_3283);
and U19746 (N_19746,N_1011,N_7356);
and U19747 (N_19747,N_5619,N_9097);
nor U19748 (N_19748,N_3554,N_5553);
nor U19749 (N_19749,N_6656,N_5860);
nand U19750 (N_19750,N_6474,N_2858);
and U19751 (N_19751,N_9511,N_4682);
nand U19752 (N_19752,N_607,N_7826);
xnor U19753 (N_19753,N_2072,N_3006);
nor U19754 (N_19754,N_7230,N_587);
and U19755 (N_19755,N_185,N_6952);
nor U19756 (N_19756,N_7099,N_3273);
or U19757 (N_19757,N_2280,N_2685);
and U19758 (N_19758,N_3650,N_7482);
or U19759 (N_19759,N_2672,N_3231);
xnor U19760 (N_19760,N_2993,N_9962);
and U19761 (N_19761,N_4485,N_2569);
or U19762 (N_19762,N_1961,N_8140);
and U19763 (N_19763,N_7093,N_2791);
and U19764 (N_19764,N_1690,N_8931);
xor U19765 (N_19765,N_2702,N_3013);
nor U19766 (N_19766,N_7310,N_5306);
nor U19767 (N_19767,N_4153,N_9829);
and U19768 (N_19768,N_982,N_4944);
and U19769 (N_19769,N_3474,N_4175);
nand U19770 (N_19770,N_5859,N_965);
xor U19771 (N_19771,N_298,N_2081);
or U19772 (N_19772,N_6014,N_7181);
or U19773 (N_19773,N_9720,N_7924);
nor U19774 (N_19774,N_3581,N_6793);
or U19775 (N_19775,N_1139,N_1416);
or U19776 (N_19776,N_4264,N_2499);
and U19777 (N_19777,N_2567,N_4105);
and U19778 (N_19778,N_7339,N_2482);
or U19779 (N_19779,N_7539,N_8144);
or U19780 (N_19780,N_4813,N_7767);
nand U19781 (N_19781,N_7822,N_7144);
nor U19782 (N_19782,N_7329,N_3264);
nand U19783 (N_19783,N_7592,N_1222);
nand U19784 (N_19784,N_2048,N_7793);
xor U19785 (N_19785,N_9963,N_2411);
or U19786 (N_19786,N_8384,N_8349);
xor U19787 (N_19787,N_498,N_612);
xnor U19788 (N_19788,N_4327,N_5571);
or U19789 (N_19789,N_8296,N_8233);
nor U19790 (N_19790,N_5824,N_9123);
xnor U19791 (N_19791,N_8887,N_1326);
nand U19792 (N_19792,N_1501,N_4539);
and U19793 (N_19793,N_4289,N_9727);
or U19794 (N_19794,N_9918,N_9293);
nor U19795 (N_19795,N_2293,N_4086);
or U19796 (N_19796,N_9375,N_3781);
nand U19797 (N_19797,N_3543,N_3032);
xor U19798 (N_19798,N_695,N_8026);
and U19799 (N_19799,N_8869,N_7994);
nand U19800 (N_19800,N_5424,N_6240);
xor U19801 (N_19801,N_7760,N_966);
and U19802 (N_19802,N_6458,N_1283);
or U19803 (N_19803,N_6403,N_8381);
xnor U19804 (N_19804,N_7790,N_2858);
and U19805 (N_19805,N_7120,N_2840);
or U19806 (N_19806,N_9064,N_6537);
and U19807 (N_19807,N_5041,N_3293);
nand U19808 (N_19808,N_860,N_2258);
nand U19809 (N_19809,N_6061,N_6155);
or U19810 (N_19810,N_3003,N_1581);
and U19811 (N_19811,N_1290,N_8090);
or U19812 (N_19812,N_8166,N_9260);
nand U19813 (N_19813,N_8755,N_6361);
or U19814 (N_19814,N_6621,N_4244);
xor U19815 (N_19815,N_8180,N_3037);
nor U19816 (N_19816,N_8733,N_8834);
nor U19817 (N_19817,N_4286,N_665);
and U19818 (N_19818,N_7942,N_1589);
nor U19819 (N_19819,N_1574,N_2552);
xnor U19820 (N_19820,N_489,N_5486);
nor U19821 (N_19821,N_5764,N_7904);
nor U19822 (N_19822,N_4039,N_6155);
nand U19823 (N_19823,N_3354,N_7372);
or U19824 (N_19824,N_3904,N_2883);
nand U19825 (N_19825,N_1634,N_8854);
or U19826 (N_19826,N_4533,N_1343);
nor U19827 (N_19827,N_101,N_8891);
nand U19828 (N_19828,N_2610,N_9245);
xnor U19829 (N_19829,N_6253,N_2398);
and U19830 (N_19830,N_277,N_3180);
nand U19831 (N_19831,N_5813,N_3080);
nor U19832 (N_19832,N_8589,N_6229);
and U19833 (N_19833,N_3562,N_317);
and U19834 (N_19834,N_4346,N_4000);
nand U19835 (N_19835,N_9361,N_7795);
xor U19836 (N_19836,N_8912,N_2111);
nor U19837 (N_19837,N_2118,N_2161);
or U19838 (N_19838,N_1672,N_4097);
nand U19839 (N_19839,N_9482,N_4297);
xnor U19840 (N_19840,N_6430,N_4492);
xor U19841 (N_19841,N_3369,N_5777);
and U19842 (N_19842,N_9518,N_6690);
and U19843 (N_19843,N_7056,N_3677);
xor U19844 (N_19844,N_5750,N_5457);
xor U19845 (N_19845,N_3006,N_657);
xnor U19846 (N_19846,N_158,N_345);
nor U19847 (N_19847,N_9287,N_1432);
or U19848 (N_19848,N_5683,N_429);
xor U19849 (N_19849,N_3053,N_1046);
or U19850 (N_19850,N_7950,N_2722);
xor U19851 (N_19851,N_9037,N_7204);
xor U19852 (N_19852,N_5455,N_1951);
and U19853 (N_19853,N_571,N_2385);
or U19854 (N_19854,N_923,N_6245);
and U19855 (N_19855,N_526,N_1893);
xor U19856 (N_19856,N_4786,N_469);
nor U19857 (N_19857,N_401,N_9474);
xor U19858 (N_19858,N_4966,N_7762);
or U19859 (N_19859,N_3214,N_395);
nor U19860 (N_19860,N_1414,N_3816);
nor U19861 (N_19861,N_7139,N_3269);
xnor U19862 (N_19862,N_2153,N_6441);
and U19863 (N_19863,N_1328,N_4651);
nand U19864 (N_19864,N_511,N_9335);
nand U19865 (N_19865,N_3153,N_6408);
nor U19866 (N_19866,N_2680,N_9579);
xnor U19867 (N_19867,N_8897,N_7096);
xor U19868 (N_19868,N_4591,N_4253);
nand U19869 (N_19869,N_1702,N_7090);
nand U19870 (N_19870,N_8418,N_6766);
and U19871 (N_19871,N_8487,N_813);
and U19872 (N_19872,N_1383,N_6826);
nand U19873 (N_19873,N_7341,N_130);
nand U19874 (N_19874,N_6420,N_705);
xnor U19875 (N_19875,N_1778,N_3233);
nor U19876 (N_19876,N_5545,N_989);
xnor U19877 (N_19877,N_1650,N_7971);
and U19878 (N_19878,N_788,N_8438);
and U19879 (N_19879,N_4339,N_1452);
xnor U19880 (N_19880,N_9824,N_5260);
and U19881 (N_19881,N_5993,N_5932);
or U19882 (N_19882,N_5312,N_7940);
xor U19883 (N_19883,N_7958,N_6179);
nand U19884 (N_19884,N_4002,N_524);
and U19885 (N_19885,N_7279,N_9874);
or U19886 (N_19886,N_9804,N_1052);
or U19887 (N_19887,N_6256,N_7870);
and U19888 (N_19888,N_2105,N_3798);
xor U19889 (N_19889,N_7822,N_7023);
or U19890 (N_19890,N_9779,N_2743);
nor U19891 (N_19891,N_6319,N_6288);
nand U19892 (N_19892,N_9348,N_9448);
nor U19893 (N_19893,N_4257,N_9947);
and U19894 (N_19894,N_3838,N_1538);
or U19895 (N_19895,N_9070,N_1880);
or U19896 (N_19896,N_1264,N_8212);
or U19897 (N_19897,N_1320,N_2609);
nand U19898 (N_19898,N_1483,N_1113);
and U19899 (N_19899,N_173,N_9373);
nor U19900 (N_19900,N_7370,N_5392);
and U19901 (N_19901,N_8622,N_1277);
nand U19902 (N_19902,N_5313,N_7929);
or U19903 (N_19903,N_9551,N_1854);
nor U19904 (N_19904,N_3042,N_6326);
xnor U19905 (N_19905,N_1249,N_3159);
nor U19906 (N_19906,N_6492,N_5005);
or U19907 (N_19907,N_2529,N_8914);
nand U19908 (N_19908,N_9561,N_7093);
and U19909 (N_19909,N_7915,N_448);
xor U19910 (N_19910,N_371,N_6352);
xnor U19911 (N_19911,N_8131,N_5928);
nor U19912 (N_19912,N_2735,N_5162);
xor U19913 (N_19913,N_2782,N_423);
nand U19914 (N_19914,N_836,N_7893);
xor U19915 (N_19915,N_2093,N_6633);
xnor U19916 (N_19916,N_2935,N_2697);
xor U19917 (N_19917,N_6618,N_7977);
and U19918 (N_19918,N_7378,N_8372);
or U19919 (N_19919,N_1345,N_4178);
xor U19920 (N_19920,N_8594,N_8083);
or U19921 (N_19921,N_2861,N_7588);
nand U19922 (N_19922,N_3287,N_978);
and U19923 (N_19923,N_4536,N_8684);
and U19924 (N_19924,N_5897,N_4538);
and U19925 (N_19925,N_1563,N_8014);
xor U19926 (N_19926,N_4761,N_8056);
xnor U19927 (N_19927,N_6937,N_1305);
xor U19928 (N_19928,N_4586,N_1341);
and U19929 (N_19929,N_3622,N_8977);
xnor U19930 (N_19930,N_5672,N_533);
or U19931 (N_19931,N_3945,N_4939);
nand U19932 (N_19932,N_9213,N_8310);
xnor U19933 (N_19933,N_9432,N_170);
or U19934 (N_19934,N_5796,N_6321);
or U19935 (N_19935,N_8252,N_7364);
xor U19936 (N_19936,N_2959,N_1843);
or U19937 (N_19937,N_3228,N_7758);
and U19938 (N_19938,N_7601,N_7704);
and U19939 (N_19939,N_9876,N_890);
xnor U19940 (N_19940,N_6028,N_8603);
xor U19941 (N_19941,N_3980,N_4252);
nand U19942 (N_19942,N_8205,N_5100);
and U19943 (N_19943,N_4023,N_7896);
nand U19944 (N_19944,N_8657,N_6791);
or U19945 (N_19945,N_6583,N_3811);
and U19946 (N_19946,N_416,N_3610);
or U19947 (N_19947,N_9951,N_7783);
nand U19948 (N_19948,N_4958,N_8384);
or U19949 (N_19949,N_6520,N_5101);
xnor U19950 (N_19950,N_3662,N_2150);
nor U19951 (N_19951,N_1926,N_9474);
nor U19952 (N_19952,N_6274,N_6140);
or U19953 (N_19953,N_2680,N_4584);
xnor U19954 (N_19954,N_9350,N_9391);
and U19955 (N_19955,N_5335,N_6950);
xor U19956 (N_19956,N_8304,N_3296);
or U19957 (N_19957,N_6120,N_5041);
nand U19958 (N_19958,N_9530,N_4036);
nand U19959 (N_19959,N_5375,N_2052);
nor U19960 (N_19960,N_1978,N_6068);
and U19961 (N_19961,N_6665,N_4753);
or U19962 (N_19962,N_1419,N_8013);
or U19963 (N_19963,N_8632,N_9325);
nor U19964 (N_19964,N_4664,N_9272);
or U19965 (N_19965,N_6587,N_496);
and U19966 (N_19966,N_8670,N_8023);
and U19967 (N_19967,N_7157,N_5333);
and U19968 (N_19968,N_3130,N_1448);
or U19969 (N_19969,N_9464,N_2460);
nor U19970 (N_19970,N_7681,N_67);
xor U19971 (N_19971,N_1129,N_8962);
or U19972 (N_19972,N_812,N_6566);
or U19973 (N_19973,N_8098,N_3406);
or U19974 (N_19974,N_4714,N_562);
nand U19975 (N_19975,N_709,N_5359);
and U19976 (N_19976,N_5462,N_6097);
nor U19977 (N_19977,N_5700,N_3619);
xor U19978 (N_19978,N_1111,N_3670);
or U19979 (N_19979,N_367,N_2278);
xnor U19980 (N_19980,N_4815,N_3979);
and U19981 (N_19981,N_5548,N_2732);
nand U19982 (N_19982,N_6753,N_8511);
and U19983 (N_19983,N_533,N_36);
and U19984 (N_19984,N_866,N_9071);
nor U19985 (N_19985,N_5031,N_7231);
or U19986 (N_19986,N_3190,N_9204);
and U19987 (N_19987,N_5948,N_6046);
xnor U19988 (N_19988,N_8118,N_6502);
and U19989 (N_19989,N_4018,N_7487);
nand U19990 (N_19990,N_5369,N_7121);
and U19991 (N_19991,N_6105,N_2919);
and U19992 (N_19992,N_3887,N_9821);
and U19993 (N_19993,N_2633,N_3460);
xor U19994 (N_19994,N_2111,N_2408);
nand U19995 (N_19995,N_639,N_647);
nor U19996 (N_19996,N_4337,N_2803);
nand U19997 (N_19997,N_9985,N_9643);
and U19998 (N_19998,N_1712,N_7187);
nand U19999 (N_19999,N_1326,N_443);
nor U20000 (N_20000,N_14817,N_11650);
and U20001 (N_20001,N_14876,N_11956);
nand U20002 (N_20002,N_15411,N_18164);
nand U20003 (N_20003,N_16340,N_15450);
or U20004 (N_20004,N_12388,N_10363);
and U20005 (N_20005,N_19249,N_15717);
xnor U20006 (N_20006,N_13355,N_18466);
xnor U20007 (N_20007,N_16993,N_14502);
xnor U20008 (N_20008,N_11097,N_15727);
xor U20009 (N_20009,N_19515,N_10633);
nand U20010 (N_20010,N_11130,N_14395);
nand U20011 (N_20011,N_13934,N_18861);
xor U20012 (N_20012,N_17262,N_12609);
xnor U20013 (N_20013,N_15360,N_14254);
xor U20014 (N_20014,N_10804,N_13496);
and U20015 (N_20015,N_16922,N_12879);
or U20016 (N_20016,N_14285,N_16857);
xor U20017 (N_20017,N_10632,N_10716);
and U20018 (N_20018,N_18988,N_16149);
xor U20019 (N_20019,N_12579,N_11174);
nand U20020 (N_20020,N_19913,N_14378);
or U20021 (N_20021,N_11727,N_10728);
xnor U20022 (N_20022,N_19564,N_17564);
or U20023 (N_20023,N_16834,N_19883);
or U20024 (N_20024,N_15183,N_10955);
xor U20025 (N_20025,N_18589,N_19219);
nor U20026 (N_20026,N_14077,N_10651);
and U20027 (N_20027,N_15057,N_11570);
nor U20028 (N_20028,N_15107,N_16514);
or U20029 (N_20029,N_10259,N_17311);
nor U20030 (N_20030,N_16425,N_18784);
or U20031 (N_20031,N_11039,N_16999);
or U20032 (N_20032,N_18142,N_10879);
xnor U20033 (N_20033,N_10807,N_17176);
nor U20034 (N_20034,N_18924,N_17475);
xnor U20035 (N_20035,N_19407,N_16729);
and U20036 (N_20036,N_17280,N_16003);
and U20037 (N_20037,N_17361,N_14619);
nor U20038 (N_20038,N_10614,N_10588);
xor U20039 (N_20039,N_13088,N_11886);
or U20040 (N_20040,N_10635,N_11361);
and U20041 (N_20041,N_13593,N_16883);
or U20042 (N_20042,N_17689,N_10886);
nor U20043 (N_20043,N_13878,N_11288);
nand U20044 (N_20044,N_15096,N_19496);
or U20045 (N_20045,N_11697,N_14074);
nand U20046 (N_20046,N_15045,N_10518);
or U20047 (N_20047,N_17547,N_16271);
nand U20048 (N_20048,N_18816,N_11232);
or U20049 (N_20049,N_15789,N_12433);
xor U20050 (N_20050,N_18324,N_16562);
xnor U20051 (N_20051,N_16748,N_11185);
xnor U20052 (N_20052,N_19850,N_10220);
xor U20053 (N_20053,N_16850,N_16973);
nor U20054 (N_20054,N_12686,N_10860);
and U20055 (N_20055,N_14553,N_14321);
xor U20056 (N_20056,N_12199,N_11731);
nand U20057 (N_20057,N_11090,N_16813);
and U20058 (N_20058,N_15810,N_15482);
nor U20059 (N_20059,N_12022,N_12976);
xnor U20060 (N_20060,N_12474,N_18225);
nor U20061 (N_20061,N_17667,N_12097);
xor U20062 (N_20062,N_11002,N_19930);
or U20063 (N_20063,N_19526,N_12325);
xnor U20064 (N_20064,N_11824,N_17650);
xnor U20065 (N_20065,N_16670,N_15580);
and U20066 (N_20066,N_14197,N_11675);
and U20067 (N_20067,N_15742,N_19052);
nand U20068 (N_20068,N_10231,N_18869);
nand U20069 (N_20069,N_14347,N_17157);
or U20070 (N_20070,N_18827,N_16653);
and U20071 (N_20071,N_15130,N_10668);
xnor U20072 (N_20072,N_16099,N_13200);
nor U20073 (N_20073,N_17010,N_19429);
or U20074 (N_20074,N_19678,N_11416);
nor U20075 (N_20075,N_16490,N_18104);
xor U20076 (N_20076,N_18519,N_19586);
nand U20077 (N_20077,N_11101,N_17495);
and U20078 (N_20078,N_18739,N_13480);
or U20079 (N_20079,N_19634,N_10704);
and U20080 (N_20080,N_11024,N_15716);
xnor U20081 (N_20081,N_17720,N_11709);
nand U20082 (N_20082,N_12883,N_12058);
nor U20083 (N_20083,N_18526,N_19375);
or U20084 (N_20084,N_18862,N_12154);
xor U20085 (N_20085,N_10270,N_18448);
or U20086 (N_20086,N_14009,N_12113);
and U20087 (N_20087,N_15233,N_13823);
and U20088 (N_20088,N_13807,N_12905);
xor U20089 (N_20089,N_10744,N_13845);
and U20090 (N_20090,N_18343,N_18981);
and U20091 (N_20091,N_13085,N_11925);
nand U20092 (N_20092,N_18282,N_11139);
and U20093 (N_20093,N_16566,N_11739);
and U20094 (N_20094,N_16202,N_14786);
xnor U20095 (N_20095,N_10180,N_13037);
nor U20096 (N_20096,N_12441,N_11620);
or U20097 (N_20097,N_18157,N_12994);
or U20098 (N_20098,N_12024,N_16779);
nor U20099 (N_20099,N_19792,N_12408);
or U20100 (N_20100,N_11729,N_10771);
and U20101 (N_20101,N_12251,N_13078);
xnor U20102 (N_20102,N_19800,N_19730);
nor U20103 (N_20103,N_15622,N_16780);
and U20104 (N_20104,N_18752,N_18396);
xor U20105 (N_20105,N_13343,N_12021);
xor U20106 (N_20106,N_13608,N_12849);
xor U20107 (N_20107,N_17437,N_10344);
nand U20108 (N_20108,N_16279,N_15744);
or U20109 (N_20109,N_18534,N_12076);
nand U20110 (N_20110,N_17096,N_12587);
and U20111 (N_20111,N_17609,N_10634);
nor U20112 (N_20112,N_17357,N_12871);
nor U20113 (N_20113,N_16840,N_17577);
and U20114 (N_20114,N_16184,N_18806);
or U20115 (N_20115,N_14204,N_17540);
or U20116 (N_20116,N_14274,N_16406);
nand U20117 (N_20117,N_19708,N_17462);
nand U20118 (N_20118,N_15026,N_18755);
and U20119 (N_20119,N_19262,N_19700);
nor U20120 (N_20120,N_10899,N_12847);
xnor U20121 (N_20121,N_12435,N_11161);
and U20122 (N_20122,N_19138,N_17319);
nand U20123 (N_20123,N_18801,N_12415);
nor U20124 (N_20124,N_10821,N_15150);
nor U20125 (N_20125,N_13021,N_16571);
or U20126 (N_20126,N_10020,N_11874);
nand U20127 (N_20127,N_13000,N_18707);
and U20128 (N_20128,N_18669,N_13975);
nand U20129 (N_20129,N_11515,N_10975);
and U20130 (N_20130,N_19383,N_12772);
nor U20131 (N_20131,N_13839,N_12747);
nand U20132 (N_20132,N_12735,N_19129);
nor U20133 (N_20133,N_15937,N_10688);
xnor U20134 (N_20134,N_12712,N_16310);
and U20135 (N_20135,N_10339,N_14960);
nor U20136 (N_20136,N_10534,N_17464);
nand U20137 (N_20137,N_13082,N_12594);
or U20138 (N_20138,N_12346,N_18386);
and U20139 (N_20139,N_19966,N_12283);
and U20140 (N_20140,N_10576,N_16606);
nand U20141 (N_20141,N_19333,N_18555);
nor U20142 (N_20142,N_16899,N_12581);
nand U20143 (N_20143,N_16258,N_16080);
nand U20144 (N_20144,N_14364,N_14911);
nor U20145 (N_20145,N_18670,N_13310);
nand U20146 (N_20146,N_16659,N_12722);
or U20147 (N_20147,N_19377,N_17915);
xnor U20148 (N_20148,N_12115,N_19231);
nor U20149 (N_20149,N_15466,N_19806);
or U20150 (N_20150,N_17429,N_13632);
xor U20151 (N_20151,N_10187,N_18231);
nor U20152 (N_20152,N_11088,N_10580);
xor U20153 (N_20153,N_19544,N_17446);
nor U20154 (N_20154,N_16020,N_17603);
nor U20155 (N_20155,N_14614,N_10065);
or U20156 (N_20156,N_11474,N_15986);
nand U20157 (N_20157,N_12632,N_10481);
or U20158 (N_20158,N_19728,N_13427);
nand U20159 (N_20159,N_11470,N_13063);
and U20160 (N_20160,N_17206,N_18043);
nor U20161 (N_20161,N_16257,N_18251);
nor U20162 (N_20162,N_10579,N_12571);
nand U20163 (N_20163,N_15079,N_19037);
xnor U20164 (N_20164,N_12019,N_13010);
or U20165 (N_20165,N_14383,N_11839);
or U20166 (N_20166,N_17648,N_19187);
or U20167 (N_20167,N_15811,N_16843);
or U20168 (N_20168,N_18754,N_12004);
nand U20169 (N_20169,N_11265,N_18724);
xnor U20170 (N_20170,N_14873,N_14213);
nand U20171 (N_20171,N_13393,N_18045);
xor U20172 (N_20172,N_14279,N_19317);
and U20173 (N_20173,N_19466,N_18905);
and U20174 (N_20174,N_19523,N_11046);
xnor U20175 (N_20175,N_19028,N_12495);
xnor U20176 (N_20176,N_11663,N_17708);
xor U20177 (N_20177,N_13905,N_13853);
and U20178 (N_20178,N_12913,N_12373);
nand U20179 (N_20179,N_15574,N_19175);
nand U20180 (N_20180,N_10949,N_14184);
xor U20181 (N_20181,N_15004,N_15205);
nand U20182 (N_20182,N_18475,N_11551);
and U20183 (N_20183,N_16868,N_16126);
xnor U20184 (N_20184,N_13906,N_19424);
xnor U20185 (N_20185,N_10723,N_11371);
or U20186 (N_20186,N_11141,N_15729);
or U20187 (N_20187,N_15316,N_12889);
and U20188 (N_20188,N_14935,N_18266);
and U20189 (N_20189,N_17693,N_19390);
nor U20190 (N_20190,N_11256,N_13354);
nand U20191 (N_20191,N_18411,N_13536);
nand U20192 (N_20192,N_15192,N_14768);
xnor U20193 (N_20193,N_19826,N_15780);
xor U20194 (N_20194,N_12316,N_11999);
or U20195 (N_20195,N_12887,N_10224);
xor U20196 (N_20196,N_13923,N_15244);
and U20197 (N_20197,N_12612,N_14672);
and U20198 (N_20198,N_15549,N_16837);
xor U20199 (N_20199,N_17387,N_19232);
nor U20200 (N_20200,N_11266,N_14419);
or U20201 (N_20201,N_11058,N_12267);
and U20202 (N_20202,N_13419,N_15544);
or U20203 (N_20203,N_11841,N_11573);
nor U20204 (N_20204,N_18623,N_16461);
nand U20205 (N_20205,N_13655,N_19550);
and U20206 (N_20206,N_13102,N_12549);
nand U20207 (N_20207,N_12836,N_13855);
or U20208 (N_20208,N_15319,N_19702);
nand U20209 (N_20209,N_11677,N_14248);
nor U20210 (N_20210,N_17065,N_18120);
nand U20211 (N_20211,N_10075,N_19787);
nand U20212 (N_20212,N_17961,N_14936);
nand U20213 (N_20213,N_14982,N_14549);
xor U20214 (N_20214,N_12635,N_17496);
and U20215 (N_20215,N_11557,N_11719);
and U20216 (N_20216,N_10725,N_12759);
and U20217 (N_20217,N_14246,N_17635);
nor U20218 (N_20218,N_12506,N_19460);
and U20219 (N_20219,N_18605,N_10206);
nor U20220 (N_20220,N_19528,N_18455);
xnor U20221 (N_20221,N_16361,N_12401);
nor U20222 (N_20222,N_19545,N_15946);
or U20223 (N_20223,N_14460,N_15975);
or U20224 (N_20224,N_15144,N_15296);
nor U20225 (N_20225,N_14979,N_16484);
and U20226 (N_20226,N_10885,N_12992);
xor U20227 (N_20227,N_19376,N_16422);
and U20228 (N_20228,N_12173,N_15342);
nor U20229 (N_20229,N_11222,N_11505);
nor U20230 (N_20230,N_14131,N_15623);
or U20231 (N_20231,N_10396,N_19404);
nand U20232 (N_20232,N_15028,N_11664);
xor U20233 (N_20233,N_14511,N_16692);
nor U20234 (N_20234,N_11264,N_12513);
xnor U20235 (N_20235,N_15215,N_13927);
nor U20236 (N_20236,N_16696,N_17951);
xor U20237 (N_20237,N_11699,N_19227);
and U20238 (N_20238,N_17155,N_15629);
nand U20239 (N_20239,N_16905,N_14703);
and U20240 (N_20240,N_14543,N_17131);
or U20241 (N_20241,N_19285,N_14828);
nor U20242 (N_20242,N_12987,N_19044);
nand U20243 (N_20243,N_10999,N_12191);
and U20244 (N_20244,N_14656,N_10529);
or U20245 (N_20245,N_14483,N_18288);
nand U20246 (N_20246,N_19856,N_12067);
xor U20247 (N_20247,N_15019,N_17247);
xor U20248 (N_20248,N_10742,N_18818);
nor U20249 (N_20249,N_18952,N_18689);
nor U20250 (N_20250,N_14886,N_17977);
and U20251 (N_20251,N_12105,N_11914);
and U20252 (N_20252,N_13737,N_13557);
and U20253 (N_20253,N_19222,N_14870);
xnor U20254 (N_20254,N_14406,N_13242);
nor U20255 (N_20255,N_11464,N_11536);
nor U20256 (N_20256,N_19611,N_19156);
xor U20257 (N_20257,N_11271,N_10465);
nand U20258 (N_20258,N_16529,N_14179);
nor U20259 (N_20259,N_13132,N_10567);
or U20260 (N_20260,N_16387,N_15899);
and U20261 (N_20261,N_19915,N_12087);
xor U20262 (N_20262,N_19463,N_12529);
nand U20263 (N_20263,N_11154,N_19047);
nor U20264 (N_20264,N_10875,N_16633);
nor U20265 (N_20265,N_14467,N_10629);
nand U20266 (N_20266,N_15765,N_14332);
nand U20267 (N_20267,N_19859,N_13746);
nor U20268 (N_20268,N_10160,N_14915);
nand U20269 (N_20269,N_10636,N_18347);
and U20270 (N_20270,N_12493,N_17967);
xnor U20271 (N_20271,N_16315,N_10972);
or U20272 (N_20272,N_18609,N_11627);
nor U20273 (N_20273,N_17188,N_18648);
xor U20274 (N_20274,N_11646,N_10559);
nor U20275 (N_20275,N_11875,N_10453);
nor U20276 (N_20276,N_18038,N_12073);
nor U20277 (N_20277,N_12121,N_19946);
nor U20278 (N_20278,N_18701,N_12095);
or U20279 (N_20279,N_10347,N_10754);
or U20280 (N_20280,N_13585,N_14806);
nand U20281 (N_20281,N_12174,N_13766);
nor U20282 (N_20282,N_16825,N_13789);
or U20283 (N_20283,N_17352,N_17578);
and U20284 (N_20284,N_10230,N_18645);
or U20285 (N_20285,N_18837,N_19416);
or U20286 (N_20286,N_18366,N_13328);
xor U20287 (N_20287,N_10805,N_11960);
and U20288 (N_20288,N_16062,N_16026);
nor U20289 (N_20289,N_17548,N_13980);
or U20290 (N_20290,N_11151,N_14740);
nand U20291 (N_20291,N_14844,N_18853);
or U20292 (N_20292,N_15171,N_16222);
xor U20293 (N_20293,N_18786,N_15879);
nand U20294 (N_20294,N_11425,N_16789);
and U20295 (N_20295,N_11817,N_17420);
or U20296 (N_20296,N_16821,N_10263);
or U20297 (N_20297,N_14331,N_19462);
xnor U20298 (N_20298,N_10929,N_18508);
or U20299 (N_20299,N_11947,N_14087);
nand U20300 (N_20300,N_18350,N_14894);
or U20301 (N_20301,N_17138,N_15615);
nand U20302 (N_20302,N_11964,N_15980);
nand U20303 (N_20303,N_13772,N_19905);
nor U20304 (N_20304,N_19816,N_15621);
nor U20305 (N_20305,N_10120,N_16122);
nor U20306 (N_20306,N_19842,N_15427);
nor U20307 (N_20307,N_13054,N_12803);
xor U20308 (N_20308,N_16097,N_11613);
nand U20309 (N_20309,N_14583,N_11418);
nor U20310 (N_20310,N_19226,N_19321);
nand U20311 (N_20311,N_16796,N_18616);
nor U20312 (N_20312,N_11867,N_10039);
nor U20313 (N_20313,N_19744,N_15317);
xnor U20314 (N_20314,N_16327,N_13898);
and U20315 (N_20315,N_14309,N_16684);
or U20316 (N_20316,N_18176,N_18427);
nor U20317 (N_20317,N_13559,N_16129);
or U20318 (N_20318,N_11420,N_17427);
nand U20319 (N_20319,N_13030,N_13040);
and U20320 (N_20320,N_10333,N_19395);
nand U20321 (N_20321,N_15039,N_14596);
or U20322 (N_20322,N_11050,N_18571);
xnor U20323 (N_20323,N_17422,N_12501);
nor U20324 (N_20324,N_19334,N_18575);
and U20325 (N_20325,N_15772,N_11370);
nor U20326 (N_20326,N_17143,N_11694);
or U20327 (N_20327,N_14375,N_17465);
or U20328 (N_20328,N_16345,N_11305);
and U20329 (N_20329,N_11652,N_12534);
nand U20330 (N_20330,N_17187,N_10294);
xor U20331 (N_20331,N_13587,N_17733);
nor U20332 (N_20332,N_11489,N_14963);
nor U20333 (N_20333,N_19260,N_16833);
and U20334 (N_20334,N_19996,N_19729);
and U20335 (N_20335,N_10587,N_11683);
xor U20336 (N_20336,N_15421,N_12952);
xor U20337 (N_20337,N_18492,N_11186);
and U20338 (N_20338,N_18116,N_12463);
nand U20339 (N_20339,N_19300,N_16826);
or U20340 (N_20340,N_14303,N_16169);
nand U20341 (N_20341,N_11228,N_14007);
xnor U20342 (N_20342,N_11527,N_13325);
or U20343 (N_20343,N_11029,N_14727);
xnor U20344 (N_20344,N_13398,N_10229);
nor U20345 (N_20345,N_12432,N_11865);
and U20346 (N_20346,N_13304,N_18733);
nor U20347 (N_20347,N_15209,N_12371);
and U20348 (N_20348,N_13064,N_11885);
or U20349 (N_20349,N_12820,N_19815);
xnor U20350 (N_20350,N_14194,N_15407);
or U20351 (N_20351,N_14252,N_13674);
xor U20352 (N_20352,N_18082,N_15981);
xnor U20353 (N_20353,N_18649,N_18208);
nand U20354 (N_20354,N_17287,N_10168);
and U20355 (N_20355,N_18388,N_17834);
and U20356 (N_20356,N_16346,N_18572);
xnor U20357 (N_20357,N_14122,N_10467);
xnor U20358 (N_20358,N_10447,N_12743);
and U20359 (N_20359,N_11635,N_16249);
and U20360 (N_20360,N_10652,N_14676);
xor U20361 (N_20361,N_16464,N_15161);
xnor U20362 (N_20362,N_15646,N_12297);
nand U20363 (N_20363,N_17724,N_13381);
nor U20364 (N_20364,N_15398,N_19503);
xor U20365 (N_20365,N_14250,N_14232);
nand U20366 (N_20366,N_17314,N_19801);
nand U20367 (N_20367,N_10987,N_14965);
xnor U20368 (N_20368,N_17736,N_14615);
xor U20369 (N_20369,N_19918,N_10193);
nand U20370 (N_20370,N_19870,N_17534);
or U20371 (N_20371,N_18783,N_13552);
nand U20372 (N_20372,N_10321,N_11533);
nor U20373 (N_20373,N_13192,N_14139);
or U20374 (N_20374,N_11014,N_10442);
nor U20375 (N_20375,N_10854,N_16352);
nor U20376 (N_20376,N_16435,N_19735);
and U20377 (N_20377,N_10441,N_14048);
nor U20378 (N_20378,N_16354,N_12578);
or U20379 (N_20379,N_11204,N_13486);
nor U20380 (N_20380,N_13420,N_19867);
and U20381 (N_20381,N_12968,N_11556);
nand U20382 (N_20382,N_10426,N_19438);
nand U20383 (N_20383,N_15196,N_18062);
xnor U20384 (N_20384,N_19516,N_12018);
nor U20385 (N_20385,N_13567,N_18437);
nand U20386 (N_20386,N_15149,N_18332);
xnor U20387 (N_20387,N_15769,N_17607);
nor U20388 (N_20388,N_16523,N_13092);
and U20389 (N_20389,N_10844,N_15782);
nor U20390 (N_20390,N_11409,N_12909);
xnor U20391 (N_20391,N_14721,N_19115);
and U20392 (N_20392,N_14925,N_19446);
or U20393 (N_20393,N_15074,N_11357);
and U20394 (N_20394,N_11250,N_14575);
xor U20395 (N_20395,N_18073,N_11172);
nor U20396 (N_20396,N_13313,N_15551);
xor U20397 (N_20397,N_12894,N_16316);
xnor U20398 (N_20398,N_12430,N_11106);
and U20399 (N_20399,N_10905,N_13209);
nor U20400 (N_20400,N_14295,N_18847);
and U20401 (N_20401,N_17747,N_18954);
xor U20402 (N_20402,N_13475,N_10539);
or U20403 (N_20403,N_17080,N_14036);
and U20404 (N_20404,N_19518,N_15325);
nor U20405 (N_20405,N_19218,N_16783);
nand U20406 (N_20406,N_11512,N_13399);
and U20407 (N_20407,N_11203,N_12178);
or U20408 (N_20408,N_18409,N_16641);
nand U20409 (N_20409,N_18564,N_16985);
and U20410 (N_20410,N_13193,N_15214);
or U20411 (N_20411,N_10026,N_12730);
nand U20412 (N_20412,N_17396,N_11594);
xor U20413 (N_20413,N_13276,N_19180);
nand U20414 (N_20414,N_16602,N_14433);
xnor U20415 (N_20415,N_19086,N_14078);
nor U20416 (N_20416,N_14944,N_11692);
nand U20417 (N_20417,N_18219,N_13890);
nor U20418 (N_20418,N_15538,N_19143);
nor U20419 (N_20419,N_10328,N_11803);
and U20420 (N_20420,N_14317,N_19844);
xnor U20421 (N_20421,N_18226,N_18740);
or U20422 (N_20422,N_15626,N_16074);
nand U20423 (N_20423,N_10416,N_10563);
or U20424 (N_20424,N_11157,N_15949);
xnor U20425 (N_20425,N_12785,N_19674);
or U20426 (N_20426,N_16071,N_14120);
nand U20427 (N_20427,N_13981,N_17779);
and U20428 (N_20428,N_10173,N_14092);
nand U20429 (N_20429,N_13631,N_16998);
or U20430 (N_20430,N_10264,N_14043);
or U20431 (N_20431,N_11661,N_16621);
or U20432 (N_20432,N_15955,N_14566);
nor U20433 (N_20433,N_17546,N_14461);
and U20434 (N_20434,N_13992,N_16479);
and U20435 (N_20435,N_10996,N_14186);
nand U20436 (N_20436,N_18684,N_15043);
or U20437 (N_20437,N_18734,N_19690);
nand U20438 (N_20438,N_10338,N_16819);
nor U20439 (N_20439,N_15996,N_11966);
nor U20440 (N_20440,N_13424,N_17434);
nand U20441 (N_20441,N_10455,N_15619);
or U20442 (N_20442,N_18741,N_15644);
xnor U20443 (N_20443,N_18108,N_10469);
and U20444 (N_20444,N_16113,N_16781);
xor U20445 (N_20445,N_17356,N_15088);
nand U20446 (N_20446,N_19743,N_13116);
xor U20447 (N_20447,N_13774,N_18635);
nand U20448 (N_20448,N_18843,N_13228);
or U20449 (N_20449,N_18556,N_12941);
and U20450 (N_20450,N_10681,N_16671);
nor U20451 (N_20451,N_18598,N_13595);
nor U20452 (N_20452,N_15997,N_18690);
and U20453 (N_20453,N_10181,N_15339);
or U20454 (N_20454,N_15486,N_16173);
nand U20455 (N_20455,N_17217,N_13635);
nand U20456 (N_20456,N_12709,N_10109);
and U20457 (N_20457,N_13361,N_10842);
xnor U20458 (N_20458,N_14634,N_18760);
nor U20459 (N_20459,N_12418,N_11226);
or U20460 (N_20460,N_11511,N_19447);
nor U20461 (N_20461,N_17112,N_19063);
xnor U20462 (N_20462,N_16193,N_11774);
xnor U20463 (N_20463,N_10155,N_14358);
nand U20464 (N_20464,N_10169,N_12036);
nor U20465 (N_20465,N_14127,N_10483);
xor U20466 (N_20466,N_11133,N_11870);
and U20467 (N_20467,N_12380,N_19234);
nor U20468 (N_20468,N_17618,N_17149);
nand U20469 (N_20469,N_14280,N_10242);
xor U20470 (N_20470,N_17412,N_19837);
nand U20471 (N_20471,N_19605,N_10279);
or U20472 (N_20472,N_11084,N_19271);
nor U20473 (N_20473,N_10492,N_10908);
or U20474 (N_20474,N_14520,N_11291);
or U20475 (N_20475,N_16775,N_17823);
or U20476 (N_20476,N_16564,N_13842);
nor U20477 (N_20477,N_16734,N_14525);
and U20478 (N_20478,N_17572,N_15932);
and U20479 (N_20479,N_13633,N_12782);
or U20480 (N_20480,N_10343,N_19750);
nor U20481 (N_20481,N_12449,N_16700);
or U20482 (N_20482,N_18200,N_17403);
and U20483 (N_20483,N_11765,N_11622);
nand U20484 (N_20484,N_17071,N_18979);
xor U20485 (N_20485,N_15651,N_10697);
nand U20486 (N_20486,N_15847,N_17294);
nand U20487 (N_20487,N_16599,N_18209);
and U20488 (N_20488,N_15610,N_12944);
nor U20489 (N_20489,N_10197,N_14753);
or U20490 (N_20490,N_15871,N_15963);
and U20491 (N_20491,N_11388,N_13533);
or U20492 (N_20492,N_17883,N_18547);
xnor U20493 (N_20493,N_13653,N_18285);
nand U20494 (N_20494,N_14144,N_13947);
nand U20495 (N_20495,N_10736,N_10045);
nand U20496 (N_20496,N_11566,N_17530);
or U20497 (N_20497,N_16655,N_18349);
nor U20498 (N_20498,N_10694,N_12478);
and U20499 (N_20499,N_10074,N_13479);
xor U20500 (N_20500,N_17838,N_19822);
or U20501 (N_20501,N_12809,N_13532);
nor U20502 (N_20502,N_19942,N_15535);
nand U20503 (N_20503,N_19060,N_18268);
xnor U20504 (N_20504,N_12570,N_12742);
nor U20505 (N_20505,N_18710,N_14244);
nand U20506 (N_20506,N_15563,N_11087);
or U20507 (N_20507,N_13275,N_11869);
nand U20508 (N_20508,N_13685,N_15102);
and U20509 (N_20509,N_12672,N_11366);
nor U20510 (N_20510,N_18368,N_17580);
or U20511 (N_20511,N_19208,N_14103);
nor U20512 (N_20512,N_19804,N_16563);
nand U20513 (N_20513,N_10918,N_16148);
nand U20514 (N_20514,N_13356,N_19761);
nand U20515 (N_20515,N_14411,N_11303);
xor U20516 (N_20516,N_17278,N_17404);
nor U20517 (N_20517,N_18533,N_10462);
and U20518 (N_20518,N_14187,N_19612);
nand U20519 (N_20519,N_18640,N_13779);
nor U20520 (N_20520,N_15724,N_11766);
or U20521 (N_20521,N_12741,N_11299);
nand U20522 (N_20522,N_13405,N_15483);
or U20523 (N_20523,N_13925,N_11877);
and U20524 (N_20524,N_11460,N_15204);
nor U20525 (N_20525,N_14760,N_11146);
or U20526 (N_20526,N_17115,N_10501);
or U20527 (N_20527,N_19981,N_15513);
and U20528 (N_20528,N_13344,N_17056);
nor U20529 (N_20529,N_11784,N_12293);
and U20530 (N_20530,N_19851,N_15854);
and U20531 (N_20531,N_17668,N_18187);
and U20532 (N_20532,N_19128,N_14064);
nand U20533 (N_20533,N_18221,N_17794);
nand U20534 (N_20534,N_15739,N_15384);
nor U20535 (N_20535,N_13696,N_17844);
and U20536 (N_20536,N_19877,N_18997);
nand U20537 (N_20537,N_19306,N_11534);
nor U20538 (N_20538,N_15506,N_12824);
nor U20539 (N_20539,N_17867,N_16908);
nand U20540 (N_20540,N_18838,N_17850);
nor U20541 (N_20541,N_17461,N_18066);
nand U20542 (N_20542,N_14695,N_12516);
xnor U20543 (N_20543,N_14329,N_14547);
xor U20544 (N_20544,N_19401,N_10618);
nor U20545 (N_20545,N_17591,N_18551);
nor U20546 (N_20546,N_11180,N_10097);
or U20547 (N_20547,N_10881,N_16224);
nand U20548 (N_20548,N_15243,N_17301);
and U20549 (N_20549,N_12298,N_15800);
nor U20550 (N_20550,N_14305,N_12713);
or U20551 (N_20551,N_11124,N_19847);
nand U20552 (N_20552,N_15691,N_18406);
or U20553 (N_20553,N_14555,N_17943);
or U20554 (N_20554,N_13022,N_10995);
xor U20555 (N_20555,N_13781,N_16530);
xor U20556 (N_20556,N_10115,N_11827);
nand U20557 (N_20557,N_19569,N_19547);
and U20558 (N_20558,N_16976,N_11140);
and U20559 (N_20559,N_19013,N_16007);
and U20560 (N_20560,N_15258,N_13333);
xor U20561 (N_20561,N_15680,N_16940);
and U20562 (N_20562,N_14455,N_16369);
or U20563 (N_20563,N_11778,N_16554);
xor U20564 (N_20564,N_13188,N_11412);
or U20565 (N_20565,N_17959,N_16644);
nand U20566 (N_20566,N_15848,N_12602);
or U20567 (N_20567,N_19449,N_15661);
nor U20568 (N_20568,N_10114,N_16194);
nand U20569 (N_20569,N_18614,N_17537);
nand U20570 (N_20570,N_12837,N_15953);
nand U20571 (N_20571,N_15386,N_10530);
nand U20572 (N_20572,N_11362,N_12303);
nor U20573 (N_20573,N_16572,N_11928);
nor U20574 (N_20574,N_17221,N_15597);
nor U20575 (N_20575,N_17421,N_19409);
and U20576 (N_20576,N_14840,N_18523);
and U20577 (N_20577,N_17478,N_15476);
nand U20578 (N_20578,N_12212,N_14464);
xor U20579 (N_20579,N_19912,N_16835);
nor U20580 (N_20580,N_16134,N_11033);
xnor U20581 (N_20581,N_16716,N_16017);
nor U20582 (N_20582,N_16521,N_19939);
nand U20583 (N_20583,N_19274,N_16704);
nand U20584 (N_20584,N_17013,N_19191);
xnor U20585 (N_20585,N_14417,N_10227);
and U20586 (N_20586,N_14326,N_14701);
xnor U20587 (N_20587,N_10682,N_13152);
or U20588 (N_20588,N_15272,N_15395);
nor U20589 (N_20589,N_19195,N_10233);
xnor U20590 (N_20590,N_19559,N_12063);
and U20591 (N_20591,N_12526,N_10841);
nand U20592 (N_20592,N_18936,N_15452);
nand U20593 (N_20593,N_11735,N_19752);
and U20594 (N_20594,N_15324,N_14865);
or U20595 (N_20595,N_11989,N_19623);
or U20596 (N_20596,N_17360,N_17453);
or U20597 (N_20597,N_19632,N_12826);
or U20598 (N_20598,N_15032,N_11597);
or U20599 (N_20599,N_13261,N_13113);
xnor U20600 (N_20600,N_14053,N_12843);
nor U20601 (N_20601,N_16947,N_16916);
nand U20602 (N_20602,N_17783,N_17510);
nand U20603 (N_20603,N_19765,N_10646);
nand U20604 (N_20604,N_12638,N_12814);
nand U20605 (N_20605,N_16895,N_10795);
or U20606 (N_20606,N_10719,N_17156);
nand U20607 (N_20607,N_14601,N_15676);
and U20608 (N_20608,N_15973,N_19980);
nor U20609 (N_20609,N_12096,N_19582);
or U20610 (N_20610,N_12204,N_18250);
and U20611 (N_20611,N_15945,N_15268);
and U20612 (N_20612,N_14730,N_14882);
xnor U20613 (N_20613,N_10400,N_14785);
nor U20614 (N_20614,N_17450,N_17432);
nor U20615 (N_20615,N_13935,N_13679);
xor U20616 (N_20616,N_13933,N_18013);
and U20617 (N_20617,N_19958,N_12522);
or U20618 (N_20618,N_11447,N_14738);
xor U20619 (N_20619,N_11293,N_19579);
or U20620 (N_20620,N_17821,N_10422);
nand U20621 (N_20621,N_13378,N_10393);
or U20622 (N_20622,N_16713,N_15014);
nand U20623 (N_20623,N_16355,N_19574);
and U20624 (N_20624,N_18770,N_19911);
and U20625 (N_20625,N_18213,N_14531);
nor U20626 (N_20626,N_10004,N_12728);
nand U20627 (N_20627,N_13126,N_17833);
xor U20628 (N_20628,N_16476,N_15058);
nand U20629 (N_20629,N_18577,N_10837);
nand U20630 (N_20630,N_16302,N_10599);
nand U20631 (N_20631,N_17334,N_11095);
nand U20632 (N_20632,N_18527,N_12437);
or U20633 (N_20633,N_15503,N_15669);
or U20634 (N_20634,N_13008,N_13880);
or U20635 (N_20635,N_14810,N_14401);
or U20636 (N_20636,N_13139,N_17180);
and U20637 (N_20637,N_14800,N_16373);
and U20638 (N_20638,N_10468,N_15967);
nor U20639 (N_20639,N_10228,N_12165);
nor U20640 (N_20640,N_10062,N_12315);
nor U20641 (N_20641,N_14051,N_12804);
and U20642 (N_20642,N_18242,N_12084);
nand U20643 (N_20643,N_12524,N_14998);
nand U20644 (N_20644,N_17817,N_15025);
nor U20645 (N_20645,N_14203,N_18891);
nand U20646 (N_20646,N_14076,N_18859);
and U20647 (N_20647,N_18620,N_10098);
nor U20648 (N_20648,N_16106,N_17505);
or U20649 (N_20649,N_18781,N_10348);
nand U20650 (N_20650,N_10390,N_17574);
and U20651 (N_20651,N_14230,N_16047);
xor U20652 (N_20652,N_14950,N_16274);
nor U20653 (N_20653,N_14170,N_14130);
xnor U20654 (N_20654,N_10198,N_18425);
nand U20655 (N_20655,N_12767,N_19637);
nand U20656 (N_20656,N_11003,N_11744);
nand U20657 (N_20657,N_18139,N_17225);
or U20658 (N_20658,N_13995,N_13720);
nor U20659 (N_20659,N_11082,N_18280);
and U20660 (N_20660,N_12170,N_10311);
nand U20661 (N_20661,N_12485,N_19099);
nand U20662 (N_20662,N_13406,N_11068);
and U20663 (N_20663,N_15712,N_11747);
nand U20664 (N_20664,N_16982,N_14106);
xor U20665 (N_20665,N_19075,N_17827);
nand U20666 (N_20666,N_19209,N_18898);
xor U20667 (N_20667,N_18910,N_15399);
nand U20668 (N_20668,N_13426,N_11499);
nand U20669 (N_20669,N_15711,N_17418);
or U20670 (N_20670,N_17238,N_19328);
or U20671 (N_20671,N_19600,N_11421);
nor U20672 (N_20672,N_14320,N_12758);
nor U20673 (N_20673,N_15966,N_17655);
xnor U20674 (N_20674,N_12841,N_13983);
nor U20675 (N_20675,N_13877,N_16002);
and U20676 (N_20676,N_11340,N_16427);
xor U20677 (N_20677,N_15954,N_19618);
nor U20678 (N_20678,N_11679,N_17805);
nand U20679 (N_20679,N_10676,N_12679);
nand U20680 (N_20680,N_13465,N_11601);
or U20681 (N_20681,N_13833,N_13960);
nand U20682 (N_20682,N_17235,N_14102);
nand U20683 (N_20683,N_19378,N_19303);
nand U20684 (N_20684,N_16350,N_13131);
or U20685 (N_20685,N_10094,N_15242);
or U20686 (N_20686,N_10461,N_10948);
nand U20687 (N_20687,N_10640,N_16496);
and U20688 (N_20688,N_19671,N_15897);
or U20689 (N_20689,N_10974,N_19428);
and U20690 (N_20690,N_13062,N_18109);
nor U20691 (N_20691,N_10748,N_19382);
and U20692 (N_20692,N_15874,N_13695);
or U20693 (N_20693,N_18041,N_11982);
nand U20694 (N_20694,N_13643,N_18585);
nor U20695 (N_20695,N_11589,N_12793);
and U20696 (N_20696,N_16028,N_19928);
and U20697 (N_20697,N_18035,N_12052);
xnor U20698 (N_20698,N_12808,N_13303);
or U20699 (N_20699,N_14431,N_18541);
or U20700 (N_20700,N_10305,N_17789);
and U20701 (N_20701,N_15902,N_14587);
or U20702 (N_20702,N_13622,N_15722);
nand U20703 (N_20703,N_10868,N_10023);
and U20704 (N_20704,N_10565,N_17560);
nor U20705 (N_20705,N_14752,N_16291);
nor U20706 (N_20706,N_12830,N_18730);
xnor U20707 (N_20707,N_13203,N_17614);
xor U20708 (N_20708,N_16096,N_16750);
xnor U20709 (N_20709,N_18792,N_19318);
nand U20710 (N_20710,N_16649,N_13210);
xnor U20711 (N_20711,N_15984,N_12796);
or U20712 (N_20712,N_11690,N_19581);
and U20713 (N_20713,N_18216,N_14257);
or U20714 (N_20714,N_17590,N_19532);
and U20715 (N_20715,N_13597,N_14990);
nand U20716 (N_20716,N_13598,N_15613);
and U20717 (N_20717,N_14192,N_17159);
nor U20718 (N_20718,N_13474,N_18940);
nor U20719 (N_20719,N_16233,N_14454);
xnor U20720 (N_20720,N_10527,N_18899);
or U20721 (N_20721,N_15307,N_19527);
or U20722 (N_20722,N_15723,N_15282);
nor U20723 (N_20723,N_15923,N_11121);
nand U20724 (N_20724,N_15794,N_17939);
or U20725 (N_20725,N_17712,N_17315);
and U20726 (N_20726,N_14576,N_12862);
nand U20727 (N_20727,N_16433,N_19812);
xor U20728 (N_20728,N_15745,N_11684);
nor U20729 (N_20729,N_18596,N_18115);
xor U20730 (N_20730,N_13752,N_14425);
nand U20731 (N_20731,N_14393,N_11304);
xnor U20732 (N_20732,N_12279,N_19412);
nor U20733 (N_20733,N_17739,N_14643);
nor U20734 (N_20734,N_19542,N_10760);
nor U20735 (N_20735,N_15821,N_11169);
and U20736 (N_20736,N_18472,N_14926);
nor U20737 (N_20737,N_10374,N_18672);
or U20738 (N_20738,N_12764,N_11815);
xor U20739 (N_20739,N_10572,N_15698);
nand U20740 (N_20740,N_14677,N_19890);
nand U20741 (N_20741,N_15101,N_19109);
or U20742 (N_20742,N_17317,N_14794);
nand U20743 (N_20743,N_16038,N_14249);
nand U20744 (N_20744,N_16838,N_17769);
nor U20745 (N_20745,N_16411,N_17531);
and U20746 (N_20746,N_17253,N_14405);
nor U20747 (N_20747,N_15013,N_15835);
and U20748 (N_20748,N_10940,N_13423);
and U20749 (N_20749,N_19495,N_18673);
xnor U20750 (N_20750,N_17364,N_11401);
nand U20751 (N_20751,N_16246,N_15468);
or U20752 (N_20752,N_11670,N_17521);
or U20753 (N_20753,N_14031,N_10508);
or U20754 (N_20754,N_18421,N_13942);
xnor U20755 (N_20755,N_17958,N_17318);
nand U20756 (N_20756,N_10324,N_19164);
and U20757 (N_20757,N_13083,N_10123);
nand U20758 (N_20758,N_15385,N_12186);
nor U20759 (N_20759,N_16478,N_11801);
and U20760 (N_20760,N_18093,N_10607);
xnor U20761 (N_20761,N_11653,N_14751);
or U20762 (N_20762,N_19188,N_15140);
and U20763 (N_20763,N_10159,N_14769);
xor U20764 (N_20764,N_13722,N_15248);
nor U20765 (N_20765,N_10548,N_18913);
and U20766 (N_20766,N_12817,N_16963);
nor U20767 (N_20767,N_13971,N_15683);
xor U20768 (N_20768,N_19386,N_16766);
xnor U20769 (N_20769,N_19727,N_15488);
nor U20770 (N_20770,N_10254,N_12075);
and U20771 (N_20771,N_15077,N_12625);
xor U20772 (N_20772,N_15689,N_16044);
nand U20773 (N_20773,N_14286,N_15852);
xor U20774 (N_20774,N_15693,N_13321);
nor U20775 (N_20775,N_16732,N_16925);
and U20776 (N_20776,N_19417,N_11704);
xor U20777 (N_20777,N_14958,N_15813);
or U20778 (N_20778,N_12781,N_15655);
nand U20779 (N_20779,N_13467,N_19149);
nand U20780 (N_20780,N_16235,N_14964);
xnor U20781 (N_20781,N_10484,N_18053);
or U20782 (N_20782,N_16549,N_10138);
xor U20783 (N_20783,N_10093,N_16970);
or U20784 (N_20784,N_19731,N_10490);
and U20785 (N_20785,N_15499,N_13862);
xnor U20786 (N_20786,N_11550,N_14193);
nand U20787 (N_20787,N_14835,N_19695);
nand U20788 (N_20788,N_17342,N_13135);
or U20789 (N_20789,N_11413,N_19916);
nand U20790 (N_20790,N_11972,N_16344);
nor U20791 (N_20791,N_14021,N_10990);
nand U20792 (N_20792,N_18369,N_12755);
nor U20793 (N_20793,N_16695,N_19964);
and U20794 (N_20794,N_12589,N_19502);
xnor U20795 (N_20795,N_13264,N_14899);
or U20796 (N_20796,N_10638,N_13736);
xnor U20797 (N_20797,N_16177,N_19694);
and U20798 (N_20798,N_11441,N_16376);
nand U20799 (N_20799,N_10673,N_12690);
nand U20800 (N_20800,N_15031,N_16162);
and U20801 (N_20801,N_19272,N_17727);
nor U20802 (N_20802,N_11623,N_10401);
xor U20803 (N_20803,N_13238,N_19920);
and U20804 (N_20804,N_12653,N_14188);
or U20805 (N_20805,N_16932,N_13520);
nand U20806 (N_20806,N_19173,N_16570);
or U20807 (N_20807,N_10806,N_15285);
or U20808 (N_20808,N_15659,N_18461);
xnor U20809 (N_20809,N_17663,N_12275);
and U20810 (N_20810,N_15362,N_14402);
xor U20811 (N_20811,N_16232,N_16923);
and U20812 (N_20812,N_17513,N_18091);
xor U20813 (N_20813,N_11100,N_17281);
xnor U20814 (N_20814,N_18301,N_18135);
xnor U20815 (N_20815,N_19114,N_12970);
or U20816 (N_20816,N_18151,N_19628);
and U20817 (N_20817,N_12511,N_19692);
nor U20818 (N_20818,N_16747,N_16705);
or U20819 (N_20819,N_14666,N_10965);
xor U20820 (N_20820,N_19161,N_16321);
xor U20821 (N_20821,N_14606,N_19038);
nand U20822 (N_20822,N_15873,N_14505);
xor U20823 (N_20823,N_13978,N_16992);
xor U20824 (N_20824,N_15909,N_12243);
nor U20825 (N_20825,N_15093,N_19740);
nor U20826 (N_20826,N_15938,N_12844);
nor U20827 (N_20827,N_13367,N_11590);
xnor U20828 (N_20828,N_16596,N_16170);
or U20829 (N_20829,N_15264,N_11122);
and U20830 (N_20830,N_19997,N_18911);
xor U20831 (N_20831,N_13036,N_10477);
nand U20832 (N_20832,N_11049,N_19033);
nand U20833 (N_20833,N_14149,N_12977);
or U20834 (N_20834,N_15990,N_16587);
nor U20835 (N_20835,N_18751,N_12588);
and U20836 (N_20836,N_17175,N_16200);
or U20837 (N_20837,N_13690,N_17785);
nor U20838 (N_20838,N_12715,N_17857);
xor U20839 (N_20839,N_13059,N_18168);
and U20840 (N_20840,N_15756,N_11569);
and U20841 (N_20841,N_11777,N_10134);
and U20842 (N_20842,N_11775,N_15797);
or U20843 (N_20843,N_13938,N_13076);
or U20844 (N_20844,N_11245,N_17597);
xnor U20845 (N_20845,N_13716,N_13527);
or U20846 (N_20846,N_18078,N_11878);
nand U20847 (N_20847,N_19948,N_17191);
or U20848 (N_20848,N_10738,N_11072);
xnor U20849 (N_20849,N_13436,N_15379);
or U20850 (N_20850,N_14611,N_14918);
and U20851 (N_20851,N_17001,N_11395);
xor U20852 (N_20852,N_15802,N_19923);
xor U20853 (N_20853,N_12788,N_13614);
xor U20854 (N_20854,N_16374,N_13699);
xnor U20855 (N_20855,N_11379,N_10286);
nor U20856 (N_20856,N_19216,N_16971);
and U20857 (N_20857,N_13339,N_18017);
or U20858 (N_20858,N_12027,N_11217);
or U20859 (N_20859,N_19960,N_10192);
nand U20860 (N_20860,N_12584,N_17452);
or U20861 (N_20861,N_19332,N_12056);
and U20862 (N_20862,N_12940,N_12031);
or U20863 (N_20863,N_14168,N_10510);
nand U20864 (N_20864,N_13128,N_14967);
or U20865 (N_20865,N_15633,N_10542);
xnor U20866 (N_20866,N_13412,N_18083);
or U20867 (N_20867,N_12870,N_12385);
xnor U20868 (N_20868,N_15352,N_13103);
and U20869 (N_20869,N_15176,N_19123);
nand U20870 (N_20870,N_18926,N_10302);
nor U20871 (N_20871,N_11609,N_18102);
nor U20872 (N_20872,N_10296,N_13484);
nor U20873 (N_20873,N_14376,N_12645);
and U20874 (N_20874,N_13299,N_16791);
xnor U20875 (N_20875,N_10261,N_13053);
nor U20876 (N_20876,N_19820,N_16590);
nand U20877 (N_20877,N_11821,N_18732);
xor U20878 (N_20878,N_18507,N_13060);
nor U20879 (N_20879,N_11493,N_14071);
nor U20880 (N_20880,N_11953,N_18536);
and U20881 (N_20881,N_16305,N_18810);
or U20882 (N_20882,N_12948,N_15453);
or U20883 (N_20883,N_19342,N_11000);
and U20884 (N_20884,N_17528,N_14707);
or U20885 (N_20885,N_10671,N_18074);
nor U20886 (N_20886,N_18064,N_14158);
or U20887 (N_20887,N_10058,N_17881);
nor U20888 (N_20888,N_16578,N_18126);
and U20889 (N_20889,N_11916,N_17353);
and U20890 (N_20890,N_18593,N_19103);
or U20891 (N_20891,N_16341,N_12288);
and U20892 (N_20892,N_16256,N_19999);
nor U20893 (N_20893,N_17900,N_10430);
xnor U20894 (N_20894,N_12416,N_14421);
nor U20895 (N_20895,N_10434,N_11247);
xor U20896 (N_20896,N_14782,N_11017);
or U20897 (N_20897,N_13286,N_16994);
or U20898 (N_20898,N_18775,N_19441);
and U20899 (N_20899,N_19287,N_11826);
or U20900 (N_20900,N_16396,N_11076);
xnor U20901 (N_20901,N_18866,N_18121);
and U20902 (N_20902,N_17643,N_17896);
and U20903 (N_20903,N_12226,N_13735);
or U20904 (N_20904,N_12885,N_12563);
nand U20905 (N_20905,N_19313,N_11595);
xnor U20906 (N_20906,N_17841,N_16016);
or U20907 (N_20907,N_15212,N_12402);
xor U20908 (N_20908,N_13899,N_11776);
xor U20909 (N_20909,N_12102,N_19588);
nor U20910 (N_20910,N_15709,N_13105);
nand U20911 (N_20911,N_11642,N_13762);
nand U20912 (N_20912,N_16746,N_14353);
nor U20913 (N_20913,N_10619,N_10749);
and U20914 (N_20914,N_13574,N_18569);
nand U20915 (N_20915,N_19500,N_18574);
nor U20916 (N_20916,N_14917,N_12656);
nand U20917 (N_20917,N_11144,N_19046);
xor U20918 (N_20918,N_19584,N_13672);
or U20919 (N_20919,N_15583,N_15173);
nor U20920 (N_20920,N_19650,N_12801);
xor U20921 (N_20921,N_17839,N_19293);
nor U20922 (N_20922,N_19641,N_16363);
nand U20923 (N_20923,N_11404,N_15527);
nor U20924 (N_20924,N_10133,N_18061);
nand U20925 (N_20925,N_11338,N_14942);
xor U20926 (N_20926,N_11298,N_19348);
or U20927 (N_20927,N_19202,N_17646);
nor U20928 (N_20928,N_11491,N_12129);
nor U20929 (N_20929,N_16853,N_12201);
nand U20930 (N_20930,N_13111,N_18283);
or U20931 (N_20931,N_13840,N_16794);
and U20932 (N_20932,N_17022,N_12482);
and U20933 (N_20933,N_18287,N_10297);
nand U20934 (N_20934,N_11189,N_11270);
or U20935 (N_20935,N_12140,N_18199);
nand U20936 (N_20936,N_10161,N_14371);
nand U20937 (N_20937,N_16269,N_14747);
xnor U20938 (N_20938,N_16088,N_18980);
xor U20939 (N_20939,N_18540,N_10925);
nor U20940 (N_20940,N_14567,N_17955);
nor U20941 (N_20941,N_13640,N_19855);
or U20942 (N_20942,N_14128,N_19602);
xnor U20943 (N_20943,N_17859,N_18478);
nor U20944 (N_20944,N_19477,N_17804);
xor U20945 (N_20945,N_18978,N_15936);
or U20946 (N_20946,N_13153,N_13662);
or U20947 (N_20947,N_13617,N_18608);
and U20948 (N_20948,N_17240,N_15255);
nor U20949 (N_20949,N_13137,N_13796);
nor U20950 (N_20950,N_14625,N_19739);
and U20951 (N_20951,N_15876,N_11733);
and U20952 (N_20952,N_17837,N_16618);
xor U20953 (N_20953,N_18180,N_13900);
nor U20954 (N_20954,N_14148,N_14245);
nor U20955 (N_20955,N_18680,N_12390);
nand U20956 (N_20956,N_12991,N_13792);
nand U20957 (N_20957,N_16755,N_17500);
and U20958 (N_20958,N_12010,N_14714);
and U20959 (N_20959,N_15682,N_13359);
nand U20960 (N_20960,N_14308,N_13347);
and U20961 (N_20961,N_11749,N_13363);
nor U20962 (N_20962,N_17331,N_19922);
and U20963 (N_20963,N_12189,N_16095);
nand U20964 (N_20964,N_16679,N_18103);
xnor U20965 (N_20965,N_14928,N_12357);
nand U20966 (N_20966,N_15658,N_17433);
xnor U20967 (N_20967,N_16174,N_19917);
xnor U20968 (N_20968,N_19746,N_10489);
nor U20969 (N_20969,N_19549,N_18028);
xor U20970 (N_20970,N_15241,N_14493);
or U20971 (N_20971,N_17889,N_18240);
or U20972 (N_20972,N_15358,N_12012);
nor U20973 (N_20973,N_12773,N_11004);
nand U20974 (N_20974,N_17263,N_17706);
nand U20975 (N_20975,N_15223,N_11907);
nor U20976 (N_20976,N_11754,N_10964);
and U20977 (N_20977,N_15987,N_13918);
nor U20978 (N_20978,N_18255,N_10361);
xnor U20979 (N_20979,N_14763,N_19145);
xor U20980 (N_20980,N_17172,N_18659);
nor U20981 (N_20981,N_19677,N_12134);
or U20982 (N_20982,N_16188,N_13387);
or U20983 (N_20983,N_15060,N_16543);
or U20984 (N_20984,N_15136,N_12467);
and U20985 (N_20985,N_13179,N_13777);
nand U20986 (N_20986,N_16845,N_14093);
and U20987 (N_20987,N_12364,N_11746);
nor U20988 (N_20988,N_10443,N_11853);
nand U20989 (N_20989,N_12945,N_10921);
nand U20990 (N_20990,N_11686,N_17299);
or U20991 (N_20991,N_17487,N_18671);
nor U20992 (N_20992,N_14352,N_14607);
nand U20993 (N_20993,N_13421,N_16820);
xor U20994 (N_20994,N_12377,N_12667);
nand U20995 (N_20995,N_17234,N_12210);
xnor U20996 (N_20996,N_13348,N_14579);
or U20997 (N_20997,N_12518,N_19071);
nor U20998 (N_20998,N_18674,N_12784);
xor U20999 (N_20999,N_12240,N_15558);
nand U21000 (N_21000,N_18341,N_10547);
nor U21001 (N_21001,N_15134,N_12412);
nor U21002 (N_21002,N_14744,N_17237);
nor U21003 (N_21003,N_12215,N_13294);
or U21004 (N_21004,N_12285,N_16103);
nand U21005 (N_21005,N_16446,N_12239);
nand U21006 (N_21006,N_18813,N_11123);
nand U21007 (N_21007,N_13052,N_16070);
or U21008 (N_21008,N_13289,N_17899);
nand U21009 (N_21009,N_14478,N_12453);
nor U21010 (N_21010,N_14126,N_18619);
or U21011 (N_21011,N_15947,N_15972);
xnor U21012 (N_21012,N_10290,N_12001);
and U21013 (N_21013,N_13851,N_12447);
nand U21014 (N_21014,N_13582,N_13642);
nand U21015 (N_21015,N_10113,N_15898);
or U21016 (N_21016,N_18844,N_19933);
or U21017 (N_21017,N_18736,N_17879);
nand U21018 (N_21018,N_16861,N_16712);
or U21019 (N_21019,N_10554,N_15041);
xnor U21020 (N_21020,N_18029,N_11958);
xnor U21021 (N_21021,N_16334,N_17529);
nand U21022 (N_21022,N_18727,N_17194);
nand U21023 (N_21023,N_15576,N_18263);
or U21024 (N_21024,N_19758,N_19938);
xnor U21025 (N_21025,N_14190,N_11211);
nor U21026 (N_21026,N_18446,N_10930);
nand U21027 (N_21027,N_12378,N_14866);
nor U21028 (N_21028,N_15286,N_19594);
nand U21029 (N_21029,N_14741,N_17582);
and U21030 (N_21030,N_13014,N_18165);
or U21031 (N_21031,N_17079,N_10141);
and U21032 (N_21032,N_18322,N_10185);
and U21033 (N_21033,N_11852,N_13508);
xnor U21034 (N_21034,N_14327,N_16195);
nor U21035 (N_21035,N_13926,N_10873);
nand U21036 (N_21036,N_10721,N_17953);
nand U21037 (N_21037,N_19255,N_12141);
and U21038 (N_21038,N_14808,N_16398);
xor U21039 (N_21039,N_12723,N_16342);
xor U21040 (N_21040,N_14242,N_11104);
nand U21041 (N_21041,N_12389,N_13554);
xnor U21042 (N_21042,N_18828,N_14724);
nor U21043 (N_21043,N_13491,N_11829);
nand U21044 (N_21044,N_15968,N_17158);
or U21045 (N_21045,N_16522,N_12703);
and U21046 (N_21046,N_11848,N_14243);
nor U21047 (N_21047,N_18581,N_10260);
or U21048 (N_21048,N_16332,N_15083);
and U21049 (N_21049,N_10622,N_17916);
nand U21050 (N_21050,N_13482,N_18016);
xnor U21051 (N_21051,N_11034,N_19048);
or U21052 (N_21052,N_16852,N_16225);
and U21053 (N_21053,N_19796,N_15710);
or U21054 (N_21054,N_12439,N_15569);
xnor U21055 (N_21055,N_19903,N_12644);
nand U21056 (N_21056,N_17973,N_15891);
or U21057 (N_21057,N_17891,N_19697);
nand U21058 (N_21058,N_14019,N_16260);
nand U21059 (N_21059,N_17726,N_15666);
nand U21060 (N_21060,N_16090,N_14535);
nand U21061 (N_21061,N_13442,N_13673);
xor U21062 (N_21062,N_11944,N_12417);
and U21063 (N_21063,N_17545,N_11814);
or U21064 (N_21064,N_16211,N_11541);
nand U21065 (N_21065,N_18092,N_18912);
or U21066 (N_21066,N_10306,N_15387);
nor U21067 (N_21067,N_13973,N_15786);
nand U21068 (N_21068,N_19458,N_11312);
or U21069 (N_21069,N_11745,N_18098);
nor U21070 (N_21070,N_13525,N_11896);
xor U21071 (N_21071,N_12908,N_17532);
nor U21072 (N_21072,N_13821,N_16555);
or U21073 (N_21073,N_17417,N_13984);
or U21074 (N_21074,N_16429,N_19657);
nand U21075 (N_21075,N_19535,N_16114);
nand U21076 (N_21076,N_16296,N_16141);
and U21077 (N_21077,N_19005,N_15290);
or U21078 (N_21078,N_19872,N_14811);
nor U21079 (N_21079,N_13318,N_19940);
xor U21080 (N_21080,N_10699,N_10158);
xnor U21081 (N_21081,N_16137,N_17980);
nand U21082 (N_21082,N_19442,N_16778);
nand U21083 (N_21083,N_14762,N_18915);
and U21084 (N_21084,N_18696,N_11194);
nand U21085 (N_21085,N_11109,N_19738);
and U21086 (N_21086,N_11846,N_10498);
nor U21087 (N_21087,N_11563,N_14355);
xnor U21088 (N_21088,N_16214,N_11147);
nor U21089 (N_21089,N_10938,N_13605);
nor U21090 (N_21090,N_14256,N_11518);
and U21091 (N_21091,N_12827,N_16380);
nand U21092 (N_21092,N_14039,N_18125);
or U21093 (N_21093,N_10631,N_18929);
nand U21094 (N_21094,N_19529,N_14546);
nand U21095 (N_21095,N_17057,N_14277);
nor U21096 (N_21096,N_10196,N_17623);
or U21097 (N_21097,N_12032,N_11094);
nor U21098 (N_21098,N_19077,N_15126);
and U21099 (N_21099,N_16737,N_16681);
xnor U21100 (N_21100,N_11725,N_11728);
xnor U21101 (N_21101,N_16418,N_12523);
or U21102 (N_21102,N_13832,N_14096);
nand U21103 (N_21103,N_15494,N_18317);
or U21104 (N_21104,N_13441,N_13531);
nor U21105 (N_21105,N_19004,N_17754);
or U21106 (N_21106,N_16836,N_12361);
or U21107 (N_21107,N_11884,N_14418);
and U21108 (N_21108,N_17994,N_12229);
xor U21109 (N_21109,N_14681,N_10040);
or U21110 (N_21110,N_12256,N_19045);
nand U21111 (N_21111,N_15071,N_11485);
and U21112 (N_21112,N_16912,N_10289);
xor U21113 (N_21113,N_13658,N_17681);
nand U21114 (N_21114,N_13308,N_18717);
or U21115 (N_21115,N_19142,N_17064);
nand U21116 (N_21116,N_10088,N_14282);
nand U21117 (N_21117,N_13012,N_15390);
nand U21118 (N_21118,N_18114,N_14105);
and U21119 (N_21119,N_16281,N_12359);
and U21120 (N_21120,N_18454,N_11374);
nand U21121 (N_21121,N_15159,N_14205);
nand U21122 (N_21122,N_14608,N_10878);
xor U21123 (N_21123,N_14972,N_18111);
nor U21124 (N_21124,N_18153,N_17744);
and U21125 (N_21125,N_10216,N_18858);
nand U21126 (N_21126,N_13186,N_12492);
nor U21127 (N_21127,N_17229,N_18808);
nand U21128 (N_21128,N_16085,N_17469);
nand U21129 (N_21129,N_18506,N_15749);
or U21130 (N_21130,N_13600,N_13217);
xnor U21131 (N_21131,N_16365,N_16581);
nand U21132 (N_21132,N_14491,N_17613);
and U21133 (N_21133,N_19998,N_18417);
nand U21134 (N_21134,N_12477,N_12494);
nor U21135 (N_21135,N_14504,N_19366);
nand U21136 (N_21136,N_11500,N_16728);
xor U21137 (N_21137,N_10586,N_18834);
or U21138 (N_21138,N_19818,N_11048);
or U21139 (N_21139,N_18884,N_16855);
xor U21140 (N_21140,N_13184,N_13464);
nor U21141 (N_21141,N_10457,N_17428);
nand U21142 (N_21142,N_19459,N_10322);
nor U21143 (N_21143,N_13703,N_19435);
xor U21144 (N_21144,N_18260,N_14569);
or U21145 (N_21145,N_13230,N_18630);
or U21146 (N_21146,N_12880,N_19054);
nor U21147 (N_21147,N_10561,N_19190);
nor U21148 (N_21148,N_13346,N_10377);
nand U21149 (N_21149,N_10695,N_10984);
nor U21150 (N_21150,N_16493,N_19268);
nor U21151 (N_21151,N_10402,N_17200);
nor U21152 (N_21152,N_17244,N_17209);
and U21153 (N_21153,N_17608,N_11923);
or U21154 (N_21154,N_12853,N_16961);
nand U21155 (N_21155,N_12925,N_16960);
and U21156 (N_21156,N_18840,N_11044);
nand U21157 (N_21157,N_15566,N_16920);
nand U21158 (N_21158,N_15461,N_13606);
or U21159 (N_21159,N_16412,N_19240);
and U21160 (N_21160,N_11530,N_16161);
or U21161 (N_21161,N_19001,N_10818);
and U21162 (N_21162,N_13477,N_18694);
xor U21163 (N_21163,N_15692,N_19244);
nor U21164 (N_21164,N_11564,N_14764);
xnor U21165 (N_21165,N_14152,N_12309);
and U21166 (N_21166,N_19610,N_12350);
and U21167 (N_21167,N_10178,N_18557);
nor U21168 (N_21168,N_17414,N_17134);
or U21169 (N_21169,N_15668,N_11372);
nor U21170 (N_21170,N_11224,N_12179);
nand U21171 (N_21171,N_12753,N_12555);
or U21172 (N_21172,N_15730,N_13417);
xnor U21173 (N_21173,N_18889,N_17483);
and U21174 (N_21174,N_16116,N_12372);
nand U21175 (N_21175,N_10284,N_15294);
nor U21176 (N_21176,N_10352,N_14877);
nand U21177 (N_21177,N_17691,N_15175);
nand U21178 (N_21178,N_14693,N_12544);
nor U21179 (N_21179,N_18431,N_19121);
nor U21180 (N_21180,N_15530,N_10832);
and U21181 (N_21181,N_10013,N_18814);
xor U21182 (N_21182,N_13196,N_12498);
xnor U21183 (N_21183,N_13856,N_19327);
and U21184 (N_21184,N_18426,N_13509);
nor U21185 (N_21185,N_15302,N_17142);
and U21186 (N_21186,N_19927,N_10456);
nor U21187 (N_21187,N_11117,N_19900);
and U21188 (N_21188,N_14821,N_17634);
nand U21189 (N_21189,N_16603,N_13743);
xor U21190 (N_21190,N_18590,N_16898);
xnor U21191 (N_21191,N_14020,N_10866);
or U21192 (N_21192,N_12185,N_15238);
or U21193 (N_21193,N_18928,N_13618);
or U21194 (N_21194,N_19414,N_15734);
or U21195 (N_21195,N_12558,N_15904);
nand U21196 (N_21196,N_14919,N_12454);
nor U21197 (N_21197,N_16459,N_11382);
nor U21198 (N_21198,N_14369,N_13243);
and U21199 (N_21199,N_12247,N_13562);
or U21200 (N_21200,N_11238,N_16849);
and U21201 (N_21201,N_17767,N_13678);
xnor U21202 (N_21202,N_10480,N_10643);
xnor U21203 (N_21203,N_17494,N_14174);
nand U21204 (N_21204,N_10856,N_19879);
xor U21205 (N_21205,N_17936,N_15271);
nor U21206 (N_21206,N_11150,N_10323);
xor U21207 (N_21207,N_15230,N_19755);
nor U21208 (N_21208,N_16050,N_10820);
and U21209 (N_21209,N_10451,N_17725);
nor U21210 (N_21210,N_15575,N_12980);
or U21211 (N_21211,N_15289,N_12697);
nor U21212 (N_21212,N_15091,N_14040);
nand U21213 (N_21213,N_17835,N_19921);
xor U21214 (N_21214,N_18352,N_17083);
nor U21215 (N_21215,N_19546,N_14586);
nand U21216 (N_21216,N_12659,N_10512);
xnor U21217 (N_21217,N_17593,N_13253);
or U21218 (N_21218,N_19525,N_10982);
and U21219 (N_21219,N_16472,N_17343);
nor U21220 (N_21220,N_13271,N_16494);
xor U21221 (N_21221,N_19955,N_13592);
nand U21222 (N_21222,N_15943,N_14268);
or U21223 (N_21223,N_14939,N_14100);
nor U21224 (N_21224,N_15526,N_13647);
nor U21225 (N_21225,N_11637,N_18147);
nor U21226 (N_21226,N_16788,N_13503);
nor U21227 (N_21227,N_12582,N_11807);
nor U21228 (N_21228,N_19615,N_14646);
xnor U21229 (N_21229,N_14976,N_15596);
and U21230 (N_21230,N_11419,N_19557);
nand U21231 (N_21231,N_12904,N_17460);
nor U21232 (N_21232,N_18832,N_13954);
or U21233 (N_21233,N_14498,N_11892);
and U21234 (N_21234,N_12397,N_13928);
nor U21235 (N_21235,N_13623,N_15141);
or U21236 (N_21236,N_11062,N_15525);
nand U21237 (N_21237,N_16157,N_17332);
nand U21238 (N_21238,N_14517,N_13967);
nand U21239 (N_21239,N_10432,N_11233);
and U21240 (N_21240,N_18949,N_17926);
nor U21241 (N_21241,N_14610,N_15762);
or U21242 (N_21242,N_16227,N_10340);
nand U21243 (N_21243,N_13513,N_12775);
nand U21244 (N_21244,N_17044,N_15701);
nand U21245 (N_21245,N_11319,N_13750);
and U21246 (N_21246,N_16120,N_19609);
and U21247 (N_21247,N_16743,N_14600);
or U21248 (N_21248,N_15773,N_15354);
nand U21249 (N_21249,N_16392,N_19355);
and U21250 (N_21250,N_19302,N_18974);
xor U21251 (N_21251,N_19865,N_14635);
or U21252 (N_21252,N_19176,N_16988);
nor U21253 (N_21253,N_15434,N_14901);
xnor U21254 (N_21254,N_13882,N_11339);
nor U21255 (N_21255,N_16431,N_12633);
nor U21256 (N_21256,N_12794,N_13047);
and U21257 (N_21257,N_10221,N_12816);
xnor U21258 (N_21258,N_14154,N_17711);
nand U21259 (N_21259,N_17869,N_12459);
nand U21260 (N_21260,N_12344,N_11423);
xor U21261 (N_21261,N_13998,N_15704);
or U21262 (N_21262,N_15970,N_13358);
xor U21263 (N_21263,N_18904,N_18955);
nand U21264 (N_21264,N_16102,N_10884);
and U21265 (N_21265,N_18223,N_12425);
nor U21266 (N_21266,N_10602,N_17113);
xnor U21267 (N_21267,N_14969,N_12542);
and U21268 (N_21268,N_14659,N_14577);
or U21269 (N_21269,N_10491,N_17685);
and U21270 (N_21270,N_19010,N_13376);
or U21271 (N_21271,N_12835,N_16203);
xor U21272 (N_21272,N_19166,N_11950);
xor U21273 (N_21273,N_13841,N_10421);
and U21274 (N_21274,N_10090,N_10048);
nand U21275 (N_21275,N_16772,N_13319);
nor U21276 (N_21276,N_13863,N_11605);
and U21277 (N_21277,N_13615,N_12332);
nor U21278 (N_21278,N_12281,N_18405);
or U21279 (N_21279,N_19693,N_13715);
xnor U21280 (N_21280,N_15455,N_10720);
and U21281 (N_21281,N_17753,N_10110);
or U21282 (N_21282,N_17519,N_18166);
and U21283 (N_21283,N_19887,N_16388);
nor U21284 (N_21284,N_11171,N_18591);
or U21285 (N_21285,N_12392,N_14824);
xnor U21286 (N_21286,N_10408,N_15763);
nand U21287 (N_21287,N_12238,N_10617);
nand U21288 (N_21288,N_11968,N_10840);
and U21289 (N_21289,N_17818,N_18921);
xor U21290 (N_21290,N_11804,N_10517);
xor U21291 (N_21291,N_10200,N_14847);
and U21292 (N_21292,N_10222,N_14773);
nand U21293 (N_21293,N_10520,N_18768);
nand U21294 (N_21294,N_13609,N_10499);
nor U21295 (N_21295,N_13669,N_14908);
nor U21296 (N_21296,N_14399,N_14859);
nor U21297 (N_21297,N_11443,N_19757);
and U21298 (N_21298,N_16645,N_10473);
nand U21299 (N_21299,N_19571,N_14397);
nor U21300 (N_21300,N_13603,N_19403);
nor U21301 (N_21301,N_12051,N_12138);
and U21302 (N_21302,N_17752,N_14337);
nor U21303 (N_21303,N_14632,N_10128);
nor U21304 (N_21304,N_18944,N_12146);
xnor U21305 (N_21305,N_10942,N_13776);
nand U21306 (N_21306,N_18878,N_11930);
nand U21307 (N_21307,N_10952,N_14795);
nand U21308 (N_21308,N_19347,N_14438);
and U21309 (N_21309,N_18748,N_14472);
nand U21310 (N_21310,N_18276,N_10726);
and U21311 (N_21311,N_13122,N_16415);
or U21312 (N_21312,N_13543,N_16597);
and U21313 (N_21313,N_14044,N_11555);
xnor U21314 (N_21314,N_15156,N_14480);
nor U21315 (N_21315,N_13537,N_13951);
nand U21316 (N_21316,N_16347,N_16301);
xor U21317 (N_21317,N_19654,N_16154);
and U21318 (N_21318,N_12646,N_11262);
nor U21319 (N_21319,N_13369,N_11207);
and U21320 (N_21320,N_16574,N_13240);
nand U21321 (N_21321,N_15977,N_18096);
nor U21322 (N_21322,N_15715,N_12479);
nor U21323 (N_21323,N_17036,N_15550);
or U21324 (N_21324,N_11648,N_11538);
and U21325 (N_21325,N_16553,N_12020);
xnor U21326 (N_21326,N_18316,N_16626);
xor U21327 (N_21327,N_19799,N_11389);
and U21328 (N_21328,N_11695,N_19672);
nor U21329 (N_21329,N_11316,N_16414);
or U21330 (N_21330,N_19021,N_14916);
nor U21331 (N_21331,N_11336,N_11086);
xor U21332 (N_21332,N_17511,N_15767);
nand U21333 (N_21333,N_19606,N_10907);
xnor U21334 (N_21334,N_19450,N_15118);
or U21335 (N_21335,N_12159,N_13414);
or U21336 (N_21336,N_15064,N_11501);
nand U21337 (N_21337,N_18613,N_10867);
nor U21338 (N_21338,N_13692,N_12443);
nand U21339 (N_21339,N_16469,N_17114);
and U21340 (N_21340,N_17369,N_19172);
nand U21341 (N_21341,N_10415,N_10735);
nor U21342 (N_21342,N_15922,N_15371);
or U21343 (N_21343,N_16014,N_16098);
xor U21344 (N_21344,N_18953,N_19684);
xor U21345 (N_21345,N_13011,N_11837);
and U21346 (N_21346,N_17335,N_15747);
nand U21347 (N_21347,N_14686,N_12762);
or U21348 (N_21348,N_12028,N_14373);
and U21349 (N_21349,N_15416,N_17674);
and U21350 (N_21350,N_17664,N_10085);
or U21351 (N_21351,N_15917,N_11038);
xor U21352 (N_21352,N_14896,N_12230);
or U21353 (N_21353,N_10199,N_16769);
nor U21354 (N_21354,N_11927,N_18222);
and U21355 (N_21355,N_13439,N_14216);
or U21356 (N_21356,N_16576,N_16600);
nand U21357 (N_21357,N_16701,N_17165);
nand U21358 (N_21358,N_12901,N_15768);
and U21359 (N_21359,N_16371,N_18065);
or U21360 (N_21360,N_15262,N_19029);
nor U21361 (N_21361,N_16913,N_16558);
nand U21362 (N_21362,N_17886,N_15085);
nand U21363 (N_21363,N_16420,N_19185);
xnor U21364 (N_21364,N_16312,N_16190);
or U21365 (N_21365,N_14793,N_18562);
and U21366 (N_21366,N_16209,N_10766);
nand U21367 (N_21367,N_11900,N_14292);
nor U21368 (N_21368,N_12903,N_10537);
and U21369 (N_21369,N_12184,N_13639);
xnor U21370 (N_21370,N_11047,N_14934);
or U21371 (N_21371,N_12535,N_13099);
nand U21372 (N_21372,N_17605,N_12777);
xnor U21373 (N_21373,N_13765,N_10139);
or U21374 (N_21374,N_10689,N_15170);
xnor U21375 (N_21375,N_10831,N_13619);
xor U21376 (N_21376,N_10372,N_19483);
xnor U21377 (N_21377,N_10170,N_17291);
xor U21378 (N_21378,N_19467,N_17447);
xnor U21379 (N_21379,N_16893,N_16632);
xor U21380 (N_21380,N_11797,N_14687);
or U21381 (N_21381,N_12374,N_11376);
xnor U21382 (N_21382,N_15795,N_17081);
and U21383 (N_21383,N_18467,N_18119);
nor U21384 (N_21384,N_18355,N_15200);
nor U21385 (N_21385,N_12974,N_12301);
xnor U21386 (N_21386,N_12321,N_16328);
nor U21387 (N_21387,N_10096,N_12916);
nor U21388 (N_21388,N_17672,N_18415);
and U21389 (N_21389,N_19733,N_18766);
xnor U21390 (N_21390,N_18232,N_16535);
or U21391 (N_21391,N_13389,N_18326);
nand U21392 (N_21392,N_11187,N_18943);
or U21393 (N_21393,N_17087,N_18118);
and U21394 (N_21394,N_14834,N_14118);
xor U21395 (N_21395,N_11149,N_13437);
or U21396 (N_21396,N_12831,N_17575);
or U21397 (N_21397,N_12130,N_19896);
and U21398 (N_21398,N_10095,N_16972);
and U21399 (N_21399,N_11796,N_19090);
xor U21400 (N_21400,N_19793,N_19660);
nor U21401 (N_21401,N_18380,N_14754);
or U21402 (N_21402,N_12317,N_17204);
or U21403 (N_21403,N_18253,N_16773);
nand U21404 (N_21404,N_10811,N_16635);
or U21405 (N_21405,N_18495,N_17745);
xor U21406 (N_21406,N_10630,N_18854);
xnor U21407 (N_21407,N_11201,N_12043);
nor U21408 (N_21408,N_11458,N_11857);
or U21409 (N_21409,N_16725,N_15599);
or U21410 (N_21410,N_16511,N_16041);
and U21411 (N_21411,N_16471,N_13039);
xor U21412 (N_21412,N_15228,N_10624);
or U21413 (N_21413,N_14335,N_15369);
xor U21414 (N_21414,N_18150,N_19863);
xnor U21415 (N_21415,N_15219,N_17588);
or U21416 (N_21416,N_16891,N_19479);
and U21417 (N_21417,N_11173,N_15495);
nor U21418 (N_21418,N_19215,N_14476);
nor U21419 (N_21419,N_10215,N_15868);
nor U21420 (N_21420,N_18975,N_10078);
xor U21421 (N_21421,N_17076,N_15487);
or U21422 (N_21422,N_13494,N_14722);
nand U21423 (N_21423,N_11552,N_15906);
or U21424 (N_21424,N_18418,N_15603);
nand U21425 (N_21425,N_10140,N_15882);
and U21426 (N_21426,N_18704,N_14143);
and U21427 (N_21427,N_10135,N_17266);
and U21428 (N_21428,N_17050,N_19595);
nand U21429 (N_21429,N_19714,N_15462);
and U21430 (N_21430,N_16946,N_17374);
nor U21431 (N_21431,N_12183,N_12422);
and U21432 (N_21432,N_10888,N_17179);
nand U21433 (N_21433,N_17697,N_10891);
nor U21434 (N_21434,N_19832,N_10751);
nor U21435 (N_21435,N_19335,N_10063);
nand U21436 (N_21436,N_14668,N_10887);
and U21437 (N_21437,N_17694,N_17947);
or U21438 (N_21438,N_18390,N_10598);
xnor U21439 (N_21439,N_18799,N_10712);
xor U21440 (N_21440,N_17275,N_14423);
xor U21441 (N_21441,N_17682,N_18503);
and U21442 (N_21442,N_19405,N_18214);
xor U21443 (N_21443,N_16817,N_15157);
xnor U21444 (N_21444,N_13191,N_16969);
xor U21445 (N_21445,N_10175,N_16266);
and U21446 (N_21446,N_14273,N_12559);
nor U21447 (N_21447,N_10507,N_12807);
nand U21448 (N_21448,N_15760,N_12424);
nand U21449 (N_21449,N_13248,N_14737);
nor U21450 (N_21450,N_13469,N_17219);
xor U21451 (N_21451,N_13208,N_12985);
xor U21452 (N_21452,N_14097,N_10277);
and U21453 (N_21453,N_16723,N_15915);
xnor U21454 (N_21454,N_15443,N_18484);
or U21455 (N_21455,N_11794,N_11722);
xnor U21456 (N_21456,N_14798,N_10367);
and U21457 (N_21457,N_16956,N_18015);
nor U21458 (N_21458,N_19194,N_17362);
nand U21459 (N_21459,N_10358,N_16462);
nand U21460 (N_21460,N_13522,N_16860);
and U21461 (N_21461,N_15903,N_16273);
and U21462 (N_21462,N_15591,N_14887);
nand U21463 (N_21463,N_17088,N_12268);
nand U21464 (N_21464,N_11575,N_16991);
nor U21465 (N_21465,N_14544,N_14088);
nand U21466 (N_21466,N_19621,N_11951);
nand U21467 (N_21467,N_14443,N_17388);
nand U21468 (N_21468,N_17983,N_19022);
nor U21469 (N_21469,N_17481,N_11917);
nor U21470 (N_21470,N_16492,N_10759);
or U21471 (N_21471,N_18387,N_17507);
nand U21472 (N_21472,N_12989,N_19280);
nor U21473 (N_21473,N_17012,N_17170);
nand U21474 (N_21474,N_19393,N_13686);
and U21475 (N_21475,N_16029,N_19399);
xor U21476 (N_21476,N_15778,N_13976);
xor U21477 (N_21477,N_19932,N_17193);
and U21478 (N_21478,N_11019,N_15764);
and U21479 (N_21479,N_13886,N_19759);
or U21480 (N_21480,N_16661,N_11941);
or U21481 (N_21481,N_18393,N_17909);
nor U21482 (N_21482,N_17380,N_10904);
xor U21483 (N_21483,N_13106,N_11738);
nor U21484 (N_21484,N_15180,N_13815);
or U21485 (N_21485,N_17557,N_11432);
and U21486 (N_21486,N_11651,N_17239);
xnor U21487 (N_21487,N_13222,N_18378);
nand U21488 (N_21488,N_15781,N_13107);
and U21489 (N_21489,N_16181,N_17642);
xnor U21490 (N_21490,N_12136,N_14211);
or U21491 (N_21491,N_10774,N_10317);
nor U21492 (N_21492,N_12023,N_13061);
and U21493 (N_21493,N_19620,N_13939);
nor U21494 (N_21494,N_19555,N_10176);
xnor U21495 (N_21495,N_14094,N_15869);
and U21496 (N_21496,N_17675,N_12047);
nor U21497 (N_21497,N_17327,N_19537);
nand U21498 (N_21498,N_19135,N_11678);
nand U21499 (N_21499,N_17908,N_19698);
nor U21500 (N_21500,N_18789,N_13921);
xnor U21501 (N_21501,N_10359,N_17459);
xor U21502 (N_21502,N_15792,N_12597);
nand U21503 (N_21503,N_14557,N_17740);
xor U21504 (N_21504,N_15638,N_16534);
nor U21505 (N_21505,N_16667,N_14265);
nor U21506 (N_21506,N_10703,N_15181);
xnor U21507 (N_21507,N_13371,N_11965);
or U21508 (N_21508,N_19036,N_16890);
or U21509 (N_21509,N_14949,N_15090);
nand U21510 (N_21510,N_16297,N_14713);
nor U21511 (N_21511,N_13773,N_14173);
xor U21512 (N_21512,N_13161,N_14494);
or U21513 (N_21513,N_14356,N_16485);
xnor U21514 (N_21514,N_10557,N_11079);
or U21515 (N_21515,N_16542,N_10024);
nor U21516 (N_21516,N_16643,N_10010);
nor U21517 (N_21517,N_18275,N_12358);
and U21518 (N_21518,N_11259,N_10288);
and U21519 (N_21519,N_19091,N_11492);
and U21520 (N_21520,N_17602,N_12041);
and U21521 (N_21521,N_15458,N_13146);
nand U21522 (N_21522,N_14997,N_16657);
xor U21523 (N_21523,N_12245,N_19397);
or U21524 (N_21524,N_14878,N_11579);
nor U21525 (N_21525,N_13901,N_10368);
xnor U21526 (N_21526,N_15276,N_15139);
nor U21527 (N_21527,N_12634,N_14767);
nor U21528 (N_21528,N_10979,N_18058);
nand U21529 (N_21529,N_18812,N_15519);
or U21530 (N_21530,N_14025,N_13656);
and U21531 (N_21531,N_12046,N_18342);
nand U21532 (N_21532,N_10172,N_18348);
xor U21533 (N_21533,N_11074,N_14006);
xor U21534 (N_21534,N_10855,N_14299);
nor U21535 (N_21535,N_17638,N_17624);
or U21536 (N_21536,N_17918,N_14902);
and U21537 (N_21537,N_13293,N_14906);
nand U21538 (N_21538,N_13066,N_19655);
nand U21539 (N_21539,N_11905,N_18072);
or U21540 (N_21540,N_14201,N_13048);
or U21541 (N_21541,N_17610,N_13638);
and U21542 (N_21542,N_13351,N_13911);
or U21543 (N_21543,N_10449,N_12086);
nor U21544 (N_21544,N_14674,N_11156);
or U21545 (N_21545,N_17104,N_15313);
nand U21546 (N_21546,N_12527,N_12623);
or U21547 (N_21547,N_16678,N_15153);
or U21548 (N_21548,N_16022,N_19908);
or U21549 (N_21549,N_18149,N_17105);
nand U21550 (N_21550,N_12823,N_18031);
and U21551 (N_21551,N_13025,N_15612);
or U21552 (N_21552,N_19858,N_16752);
and U21553 (N_21553,N_14209,N_16907);
nor U21554 (N_21554,N_18726,N_12249);
or U21555 (N_21555,N_19778,N_14237);
nor U21556 (N_21556,N_17224,N_17018);
and U21557 (N_21557,N_16797,N_18252);
xnor U21558 (N_21558,N_10765,N_10445);
nand U21559 (N_21559,N_10089,N_14787);
nand U21560 (N_21560,N_14671,N_16882);
xnor U21561 (N_21561,N_13768,N_18697);
nor U21562 (N_21562,N_17765,N_17737);
and U21563 (N_21563,N_12988,N_15460);
and U21564 (N_21564,N_11565,N_13804);
nand U21565 (N_21565,N_18246,N_18359);
and U21566 (N_21566,N_19995,N_19649);
or U21567 (N_21567,N_15783,N_18903);
and U21568 (N_21568,N_11089,N_19337);
or U21569 (N_21569,N_16611,N_17174);
xor U21570 (N_21570,N_11066,N_10406);
xor U21571 (N_21571,N_10091,N_17302);
or U21572 (N_21572,N_14561,N_18229);
and U21573 (N_21573,N_10664,N_14871);
or U21574 (N_21574,N_16816,N_17241);
xnor U21575 (N_21575,N_17061,N_14957);
or U21576 (N_21576,N_13616,N_18173);
nand U21577 (N_21577,N_14125,N_17907);
xnor U21578 (N_21578,N_17038,N_13296);
or U21579 (N_21579,N_16810,N_14429);
or U21580 (N_21580,N_10407,N_17276);
or U21581 (N_21581,N_17423,N_12754);
or U21582 (N_21582,N_16885,N_17488);
nor U21583 (N_21583,N_16848,N_17870);
nor U21584 (N_21584,N_12606,N_16012);
nor U21585 (N_21585,N_17903,N_18494);
xor U21586 (N_21586,N_11787,N_12643);
nor U21587 (N_21587,N_18195,N_14221);
nor U21588 (N_21588,N_18796,N_19298);
and U21589 (N_21589,N_10653,N_16045);
xor U21590 (N_21590,N_17391,N_10514);
and U21591 (N_21591,N_15069,N_12221);
nor U21592 (N_21592,N_16715,N_10156);
and U21593 (N_21593,N_10253,N_19914);
or U21594 (N_21594,N_13651,N_11192);
nor U21595 (N_21595,N_10051,N_18501);
and U21596 (N_21596,N_18688,N_16579);
or U21597 (N_21597,N_18592,N_17758);
and U21598 (N_21598,N_15738,N_15887);
xor U21599 (N_21599,N_17987,N_12965);
nor U21600 (N_21600,N_14952,N_17583);
nand U21601 (N_21601,N_10794,N_14857);
or U21602 (N_21602,N_16463,N_14488);
and U21603 (N_21603,N_19862,N_16247);
nor U21604 (N_21604,N_12616,N_17806);
and U21605 (N_21605,N_19603,N_16254);
nor U21606 (N_21606,N_13287,N_11582);
nand U21607 (N_21607,N_15410,N_10544);
nor U21608 (N_21608,N_15138,N_19150);
nand U21609 (N_21609,N_18566,N_16282);
or U21610 (N_21610,N_11510,N_19499);
or U21611 (N_21611,N_13056,N_15572);
or U21612 (N_21612,N_10268,N_16460);
xnor U21613 (N_21613,N_16945,N_14898);
nor U21614 (N_21614,N_16756,N_14593);
nand U21615 (N_21615,N_17686,N_14075);
and U21616 (N_21616,N_15528,N_10330);
and U21617 (N_21617,N_15958,N_11991);
xnor U21618 (N_21618,N_13702,N_14380);
xnor U21619 (N_21619,N_15158,N_12074);
xor U21620 (N_21620,N_10503,N_11384);
and U21621 (N_21621,N_13285,N_19782);
xnor U21622 (N_21622,N_17536,N_17949);
or U21623 (N_21623,N_13590,N_10926);
xnor U21624 (N_21624,N_15137,N_10310);
nor U21625 (N_21625,N_17449,N_19206);
and U21626 (N_21626,N_19374,N_19464);
nand U21627 (N_21627,N_12620,N_16864);
xnor U21628 (N_21628,N_18932,N_18856);
xnor U21629 (N_21629,N_10861,N_15927);
nand U21630 (N_21630,N_18227,N_15880);
and U21631 (N_21631,N_18374,N_14226);
nor U21632 (N_21632,N_14836,N_12756);
nand U21633 (N_21633,N_11134,N_17653);
xnor U21634 (N_21634,N_17151,N_18545);
and U21635 (N_21635,N_18248,N_13453);
xor U21636 (N_21636,N_16634,N_14109);
nor U21637 (N_21637,N_17304,N_17954);
and U21638 (N_21638,N_18749,N_19267);
nor U21639 (N_21639,N_17562,N_17535);
or U21640 (N_21640,N_16018,N_17004);
nor U21641 (N_21641,N_10079,N_15732);
nor U21642 (N_21642,N_19710,N_16025);
and U21643 (N_21643,N_11269,N_19889);
nand U21644 (N_21644,N_18525,N_19821);
nand U21645 (N_21645,N_19139,N_18968);
nand U21646 (N_21646,N_19919,N_19305);
nand U21647 (N_21647,N_19504,N_15334);
nor U21648 (N_21648,N_17722,N_11036);
nand U21649 (N_21649,N_11502,N_16482);
nand U21650 (N_21650,N_18795,N_18661);
nor U21651 (N_21651,N_14616,N_18408);
or U21652 (N_21652,N_16575,N_16518);
or U21653 (N_21653,N_16656,N_14099);
or U21654 (N_21654,N_17549,N_11871);
xnor U21655 (N_21655,N_10793,N_18893);
and U21656 (N_21656,N_19198,N_11213);
nor U21657 (N_21657,N_19986,N_13502);
nor U21658 (N_21658,N_14895,N_15600);
xor U21659 (N_21659,N_17375,N_11660);
nand U21660 (N_21660,N_12410,N_14313);
nor U21661 (N_21661,N_18033,N_10280);
xor U21662 (N_21662,N_16547,N_19089);
nor U21663 (N_21663,N_13162,N_11195);
and U21664 (N_21664,N_18377,N_12890);
nor U21665 (N_21665,N_14663,N_11358);
nor U21666 (N_21666,N_10162,N_12554);
xnor U21667 (N_21667,N_11724,N_11482);
nand U21668 (N_21668,N_11581,N_15812);
xnor U21669 (N_21669,N_14261,N_12481);
xor U21670 (N_21670,N_14509,N_16668);
and U21671 (N_21671,N_19420,N_13314);
or U21672 (N_21672,N_14123,N_19803);
nor U21673 (N_21673,N_13545,N_16801);
xnor U21674 (N_21674,N_10037,N_17359);
nor U21675 (N_21675,N_18465,N_18985);
nand U21676 (N_21676,N_10958,N_18325);
nand U21677 (N_21677,N_18785,N_12957);
nor U21678 (N_21678,N_16762,N_13711);
nand U21679 (N_21679,N_19182,N_11347);
nand U21680 (N_21680,N_15122,N_16262);
xnor U21681 (N_21681,N_15775,N_18872);
xor U21682 (N_21682,N_12490,N_17632);
or U21683 (N_21683,N_19653,N_10000);
or U21684 (N_21684,N_15397,N_12312);
or U21685 (N_21685,N_17596,N_11844);
nand U21686 (N_21686,N_18457,N_13090);
nand U21687 (N_21687,N_19019,N_10423);
xnor U21688 (N_21688,N_10755,N_12101);
xor U21689 (N_21689,N_18621,N_11808);
and U21690 (N_21690,N_11971,N_18647);
xnor U21691 (N_21691,N_12918,N_12103);
xor U21692 (N_21692,N_18665,N_14005);
nor U21693 (N_21693,N_17543,N_10770);
nand U21694 (N_21694,N_12175,N_11621);
and U21695 (N_21695,N_15785,N_10257);
nand U21696 (N_21696,N_13227,N_18638);
nor U21697 (N_21697,N_13985,N_12457);
nand U21698 (N_21698,N_10248,N_10371);
or U21699 (N_21699,N_13534,N_11616);
and U21700 (N_21700,N_15512,N_17363);
nand U21701 (N_21701,N_17408,N_18099);
or U21702 (N_21702,N_14907,N_14255);
nor U21703 (N_21703,N_11522,N_13350);
xnor U21704 (N_21704,N_10394,N_19824);
or U21705 (N_21705,N_16787,N_17456);
nand U21706 (N_21706,N_11850,N_12008);
or U21707 (N_21707,N_10146,N_17125);
and U21708 (N_21708,N_18990,N_19651);
xnor U21709 (N_21709,N_15529,N_16468);
nand U21710 (N_21710,N_14161,N_17964);
or U21711 (N_21711,N_18451,N_17702);
xor U21712 (N_21712,N_17289,N_15681);
or U21713 (N_21713,N_10122,N_14367);
nand U21714 (N_21714,N_14435,N_10714);
nor U21715 (N_21715,N_11255,N_17937);
and U21716 (N_21716,N_14334,N_17633);
nand U21717 (N_21717,N_13224,N_12618);
nor U21718 (N_21718,N_19247,N_16818);
and U21719 (N_21719,N_17355,N_10353);
or U21720 (N_21720,N_10417,N_18982);
xnor U21721 (N_21721,N_12335,N_17945);
nor U21722 (N_21722,N_14165,N_15776);
and U21723 (N_21723,N_11897,N_14013);
nor U21724 (N_21724,N_11126,N_13941);
nand U21725 (N_21725,N_18713,N_17377);
xor U21726 (N_21726,N_11355,N_18846);
xnor U21727 (N_21727,N_13786,N_12104);
nor U21728 (N_21728,N_11909,N_11790);
and U21729 (N_21729,N_14684,N_18186);
nor U21730 (N_21730,N_19361,N_16951);
nand U21731 (N_21731,N_13081,N_11647);
xnor U21732 (N_21732,N_12195,N_11393);
xor U21733 (N_21733,N_13993,N_17132);
nand U21734 (N_21734,N_10046,N_14104);
nor U21735 (N_21735,N_15378,N_18538);
nor U21736 (N_21736,N_10611,N_14340);
nor U21737 (N_21737,N_15799,N_10511);
nand U21738 (N_21738,N_12640,N_12322);
nor U21739 (N_21739,N_17486,N_18860);
nand U21740 (N_21740,N_12168,N_15746);
xnor U21741 (N_21741,N_11615,N_18714);
nand U21742 (N_21742,N_11445,N_13229);
xor U21743 (N_21743,N_14699,N_14302);
nand U21744 (N_21744,N_18825,N_16440);
xnor U21745 (N_21745,N_12787,N_17710);
and U21746 (N_21746,N_12233,N_10053);
and U21747 (N_21747,N_14937,N_12258);
and U21748 (N_21748,N_11755,N_17759);
and U21749 (N_21749,N_18100,N_15218);
nor U21750 (N_21750,N_13345,N_17842);
and U21751 (N_21751,N_14484,N_18906);
and U21752 (N_21752,N_15751,N_13338);
or U21753 (N_21753,N_12708,N_16207);
nor U21754 (N_21754,N_12469,N_12272);
and U21755 (N_21755,N_18063,N_14930);
or U21756 (N_21756,N_15962,N_16595);
or U21757 (N_21757,N_12912,N_13215);
or U21758 (N_21758,N_17196,N_13027);
xnor U21759 (N_21759,N_14238,N_11127);
or U21760 (N_21760,N_16901,N_19310);
xor U21761 (N_21761,N_14617,N_14003);
and U21762 (N_21762,N_18685,N_17011);
nand U21763 (N_21763,N_18138,N_14336);
xnor U21764 (N_21764,N_18463,N_14669);
nand U21765 (N_21765,N_18782,N_19237);
nand U21766 (N_21766,N_17671,N_16319);
and U21767 (N_21767,N_12166,N_12207);
xor U21768 (N_21768,N_17358,N_11976);
xnor U21769 (N_21769,N_16497,N_11524);
or U21770 (N_21770,N_19491,N_19885);
nand U21771 (N_21771,N_19481,N_19745);
xnor U21772 (N_21772,N_11349,N_17700);
or U21773 (N_21773,N_18156,N_14604);
or U21774 (N_21774,N_11181,N_17255);
xnor U21775 (N_21775,N_12461,N_11931);
nand U21776 (N_21776,N_17876,N_17144);
nand U21777 (N_21777,N_18951,N_10924);
nor U21778 (N_21778,N_17286,N_14177);
and U21779 (N_21779,N_13604,N_18003);
nor U21780 (N_21780,N_11643,N_18699);
and U21781 (N_21781,N_10513,N_10777);
nor U21782 (N_21782,N_15517,N_16944);
nor U21783 (N_21783,N_15011,N_11845);
xnor U21784 (N_21784,N_15587,N_11367);
or U21785 (N_21785,N_13808,N_11313);
xnor U21786 (N_21786,N_16933,N_14757);
or U21787 (N_21787,N_12975,N_11577);
xnor U21788 (N_21788,N_14850,N_17840);
xnor U21789 (N_21789,N_13586,N_18563);
xor U21790 (N_21790,N_16995,N_18021);
or U21791 (N_21791,N_18535,N_10817);
or U21792 (N_21792,N_11495,N_13664);
and U21793 (N_21793,N_11514,N_10890);
and U21794 (N_21794,N_14157,N_10897);
and U21795 (N_21795,N_10909,N_16516);
and U21796 (N_21796,N_17039,N_16910);
nand U21797 (N_21797,N_19652,N_19326);
or U21798 (N_21798,N_17348,N_18090);
nor U21799 (N_21799,N_10946,N_10889);
or U21800 (N_21800,N_19023,N_17215);
xnor U21801 (N_21801,N_13080,N_19626);
or U21802 (N_21802,N_14473,N_18583);
or U21803 (N_21803,N_16869,N_18385);
and U21804 (N_21804,N_11954,N_18737);
nand U21805 (N_21805,N_17378,N_16565);
xor U21806 (N_21806,N_11764,N_11403);
xor U21807 (N_21807,N_19967,N_12237);
nand U21808 (N_21808,N_13570,N_12203);
nand U21809 (N_21809,N_16448,N_16306);
nand U21810 (N_21810,N_19971,N_19886);
or U21811 (N_21811,N_19617,N_16902);
or U21812 (N_21812,N_17730,N_16583);
xnor U21813 (N_21813,N_14734,N_14000);
or U21814 (N_21814,N_12695,N_16759);
or U21815 (N_21815,N_16842,N_18992);
xnor U21816 (N_21816,N_17851,N_11341);
nor U21817 (N_21817,N_10436,N_18916);
and U21818 (N_21818,N_14755,N_12539);
or U21819 (N_21819,N_19869,N_13749);
nor U21820 (N_21820,N_16311,N_18389);
or U21821 (N_21821,N_15401,N_10150);
and U21822 (N_21822,N_11588,N_13018);
nor U21823 (N_21823,N_18067,N_11994);
xnor U21824 (N_21824,N_18277,N_15901);
and U21825 (N_21825,N_18935,N_18196);
xor U21826 (N_21826,N_10916,N_17749);
and U21827 (N_21827,N_18230,N_10983);
and U21828 (N_21828,N_17815,N_13675);
nand U21829 (N_21829,N_19102,N_17616);
and U21830 (N_21830,N_11277,N_14422);
and U21831 (N_21831,N_11065,N_11737);
and U21832 (N_21832,N_19852,N_17345);
or U21833 (N_21833,N_12935,N_18211);
nand U21834 (N_21834,N_10944,N_12930);
and U21835 (N_21835,N_17223,N_11561);
nor U21836 (N_21836,N_15308,N_15964);
nor U21837 (N_21837,N_15628,N_12811);
xnor U21838 (N_21838,N_11910,N_12954);
nor U21839 (N_21839,N_12668,N_15145);
nor U21840 (N_21840,N_11322,N_19391);
xor U21841 (N_21841,N_18500,N_12375);
nor U21842 (N_21842,N_19489,N_14492);
nor U21843 (N_21843,N_16954,N_16917);
nor U21844 (N_21844,N_13860,N_17902);
and U21845 (N_21845,N_15166,N_19476);
nor U21846 (N_21846,N_17407,N_19357);
nand U21847 (N_21847,N_11356,N_19193);
or U21848 (N_21848,N_15700,N_19130);
xor U21849 (N_21849,N_15279,N_10761);
nand U21850 (N_21850,N_12037,N_17892);
and U21851 (N_21851,N_17062,N_10970);
xnor U21852 (N_21852,N_15861,N_19154);
nor U21853 (N_21853,N_13225,N_12761);
xnor U21854 (N_21854,N_12961,N_14439);
xnor U21855 (N_21855,N_14271,N_15198);
and U21856 (N_21856,N_18473,N_18514);
or U21857 (N_21857,N_18141,N_17952);
or U21858 (N_21858,N_12628,N_14159);
or U21859 (N_21859,N_15284,N_10127);
xor U21860 (N_21860,N_17222,N_13826);
and U21861 (N_21861,N_10082,N_17124);
xor U21862 (N_21862,N_15338,N_18207);
xnor U21863 (N_21863,N_11943,N_15112);
nand U21864 (N_21864,N_14178,N_18983);
nand U21865 (N_21865,N_10201,N_10252);
and U21866 (N_21866,N_19353,N_18442);
nand U21867 (N_21867,N_12651,N_17069);
nand U21868 (N_21868,N_12356,N_12035);
nor U21869 (N_21869,N_17595,N_18416);
and U21870 (N_21870,N_10382,N_19372);
nor U21871 (N_21871,N_13372,N_17746);
and U21872 (N_21872,N_18743,N_15263);
and U21873 (N_21873,N_12464,N_11096);
nor U21874 (N_21874,N_14580,N_15344);
nand U21875 (N_21875,N_18382,N_17025);
and U21876 (N_21876,N_19985,N_17161);
and U21877 (N_21877,N_14098,N_13485);
nand U21878 (N_21878,N_10610,N_18880);
nand U21879 (N_21879,N_18757,N_16027);
or U21880 (N_21880,N_11937,N_10272);
xnor U21881 (N_21881,N_15148,N_12568);
nor U21882 (N_21882,N_11196,N_10116);
or U21883 (N_21883,N_17108,N_15894);
and U21884 (N_21884,N_12429,N_16379);
xnor U21885 (N_21885,N_17942,N_17874);
nor U21886 (N_21886,N_12034,N_13432);
nand U21887 (N_21887,N_16568,N_13870);
or U21888 (N_21888,N_14442,N_17541);
and U21889 (N_21889,N_10131,N_12960);
and U21890 (N_21890,N_16625,N_15501);
xor U21891 (N_21891,N_17316,N_11008);
nor U21892 (N_21892,N_12246,N_11220);
nand U21893 (N_21893,N_12426,N_11586);
xor U21894 (N_21894,N_18077,N_13883);
and U21895 (N_21895,N_10488,N_10910);
nand U21896 (N_21896,N_11307,N_19860);
nand U21897 (N_21897,N_19984,N_18131);
nand U21898 (N_21898,N_13729,N_12384);
nor U21899 (N_21899,N_18646,N_18691);
or U21900 (N_21900,N_12532,N_11060);
or U21901 (N_21901,N_16851,N_16776);
and U21902 (N_21902,N_11215,N_19263);
nand U21903 (N_21903,N_19101,N_18330);
nand U21904 (N_21904,N_17454,N_15346);
xnor U21905 (N_21905,N_11183,N_18769);
nor U21906 (N_21906,N_16243,N_11351);
xor U21907 (N_21907,N_19486,N_13902);
nor U21908 (N_21908,N_18587,N_14300);
and U21909 (N_21909,N_10001,N_13657);
nor U21910 (N_21910,N_11759,N_10600);
nor U21911 (N_21911,N_15306,N_10309);
nand U21912 (N_21912,N_12607,N_12194);
xnor U21913 (N_21913,N_13413,N_13301);
nor U21914 (N_21914,N_11431,N_14220);
nand U21915 (N_21915,N_10007,N_10105);
nand U21916 (N_21916,N_17052,N_16601);
nand U21917 (N_21917,N_12919,N_16741);
nor U21918 (N_21918,N_11862,N_18517);
xor U21919 (N_21919,N_19763,N_15007);
nor U21920 (N_21920,N_18019,N_17373);
or U21921 (N_21921,N_12124,N_17922);
nand U21922 (N_21922,N_17862,N_13390);
and U21923 (N_21923,N_19080,N_13006);
and U21924 (N_21924,N_18582,N_15706);
and U21925 (N_21925,N_10414,N_13997);
xnor U21926 (N_21926,N_11311,N_14287);
nor U21927 (N_21927,N_12874,N_19703);
and U21928 (N_21928,N_16795,N_11437);
or U21929 (N_21929,N_12066,N_12510);
and U21930 (N_21930,N_13178,N_18611);
nand U21931 (N_21931,N_15234,N_10460);
and U21932 (N_21932,N_14023,N_11542);
xnor U21933 (N_21933,N_13687,N_12419);
nand U21934 (N_21934,N_15133,N_10989);
and U21935 (N_21935,N_14012,N_19720);
nor U21936 (N_21936,N_17110,N_19178);
nand U21937 (N_21937,N_15128,N_13282);
nand U21938 (N_21938,N_10667,N_19116);
xnor U21939 (N_21939,N_17037,N_11767);
and U21940 (N_21940,N_11547,N_15860);
and U21941 (N_21941,N_12294,N_12351);
xnor U21942 (N_21942,N_17472,N_15095);
nand U21943 (N_21943,N_17893,N_13185);
or U21944 (N_21944,N_19880,N_14578);
or U21945 (N_21945,N_19256,N_17035);
and U21946 (N_21946,N_14240,N_11835);
nand U21947 (N_21947,N_19451,N_17371);
or U21948 (N_21948,N_15830,N_15920);
and U21949 (N_21949,N_16031,N_10153);
nor U21950 (N_21950,N_17802,N_12922);
or U21951 (N_21951,N_17539,N_19699);
nand U21952 (N_21952,N_17394,N_11598);
nand U21953 (N_21953,N_19320,N_15656);
nand U21954 (N_21954,N_16330,N_10103);
or U21955 (N_21955,N_10843,N_18037);
or U21956 (N_21956,N_13667,N_13016);
nand U21957 (N_21957,N_16451,N_19795);
nand U21958 (N_21958,N_12328,N_16569);
nand U21959 (N_21959,N_12639,N_13257);
and U21960 (N_21960,N_11306,N_18363);
xor U21961 (N_21961,N_16058,N_10019);
xnor U21962 (N_21962,N_19884,N_19840);
or U21963 (N_21963,N_19124,N_19057);
xor U21964 (N_21964,N_10291,N_10069);
or U21965 (N_21965,N_13307,N_19371);
xnor U21966 (N_21966,N_13147,N_16043);
nand U21967 (N_21967,N_18192,N_19514);
nand U21968 (N_21968,N_13150,N_15131);
xnor U21969 (N_21969,N_17182,N_19125);
nand U21970 (N_21970,N_13251,N_13397);
or U21971 (N_21971,N_17814,N_13914);
and U21972 (N_21972,N_16764,N_12655);
and U21973 (N_21973,N_19443,N_13676);
nand U21974 (N_21974,N_19636,N_11369);
nor U21975 (N_21975,N_15259,N_16140);
nor U21976 (N_21976,N_13199,N_17381);
nor U21977 (N_21977,N_16580,N_12143);
nor U21978 (N_21978,N_17913,N_12990);
xor U21979 (N_21979,N_13915,N_18201);
nor U21980 (N_21980,N_16087,N_15174);
or U21981 (N_21981,N_19539,N_11544);
or U21982 (N_21982,N_11410,N_14839);
xnor U21983 (N_21983,N_17026,N_16444);
and U21984 (N_21984,N_15021,N_15470);
nand U21985 (N_21985,N_11614,N_19379);
and U21986 (N_21986,N_11252,N_10137);
xor U21987 (N_21987,N_16336,N_11856);
nor U21988 (N_21988,N_17509,N_11760);
nand U21989 (N_21989,N_12360,N_10049);
nand U21990 (N_21990,N_12090,N_15624);
nand U21991 (N_21991,N_12984,N_19593);
nand U21992 (N_21992,N_16453,N_17111);
nor U21993 (N_21993,N_11053,N_12867);
and U21994 (N_21994,N_14137,N_12015);
nand U21995 (N_21995,N_19953,N_13682);
and U21996 (N_21996,N_15087,N_16034);
nand U21997 (N_21997,N_10083,N_16953);
nand U21998 (N_21998,N_10251,N_14776);
or U21999 (N_21999,N_15803,N_12859);
or U22000 (N_22000,N_11743,N_17666);
xnor U22001 (N_22001,N_14862,N_14387);
xor U22002 (N_22002,N_13500,N_19646);
nor U22003 (N_22003,N_16782,N_17625);
and U22004 (N_22004,N_18333,N_13785);
xor U22005 (N_22005,N_14059,N_19893);
nand U22006 (N_22006,N_18946,N_14670);
nand U22007 (N_22007,N_11708,N_17846);
and U22008 (N_22008,N_16751,N_17129);
or U22009 (N_22009,N_17709,N_15866);
and U22010 (N_22010,N_17041,N_18991);
and U22011 (N_22011,N_16708,N_10934);
xor U22012 (N_22012,N_18835,N_19607);
nand U22013 (N_22013,N_11730,N_11847);
nand U22014 (N_22014,N_10797,N_13493);
nor U22015 (N_22015,N_14113,N_17669);
nand U22016 (N_22016,N_14897,N_14207);
nor U22017 (N_22017,N_18907,N_19275);
nand U22018 (N_22018,N_15908,N_12860);
or U22019 (N_22019,N_12562,N_14033);
nand U22020 (N_22020,N_13236,N_19907);
or U22021 (N_22021,N_11855,N_17699);
and U22022 (N_22022,N_12866,N_11456);
xnor U22023 (N_22023,N_11486,N_16163);
nand U22024 (N_22024,N_11221,N_13070);
nand U22025 (N_22025,N_19601,N_15905);
xor U22026 (N_22026,N_18224,N_14377);
nor U22027 (N_22027,N_15929,N_13326);
and U22028 (N_22028,N_13385,N_11005);
nor U22029 (N_22029,N_19667,N_15940);
xor U22030 (N_22030,N_15757,N_14642);
xnor U22031 (N_22031,N_12779,N_14833);
nor U22032 (N_22032,N_17468,N_12304);
or U22033 (N_22033,N_10583,N_18189);
xor U22034 (N_22034,N_12216,N_17576);
and U22035 (N_22035,N_15976,N_17074);
xor U22036 (N_22036,N_11310,N_19522);
nor U22037 (N_22037,N_10351,N_14661);
and U22038 (N_22038,N_10645,N_19556);
nor U22039 (N_22039,N_18075,N_14169);
nor U22040 (N_22040,N_19235,N_11619);
nand U22041 (N_22041,N_17705,N_10858);
and U22042 (N_22042,N_10386,N_16986);
nor U22043 (N_22043,N_19817,N_13875);
nor U22044 (N_22044,N_16941,N_12329);
nor U22045 (N_22045,N_14655,N_15431);
xor U22046 (N_22046,N_11741,N_17781);
xor U22047 (N_22047,N_11015,N_10785);
nand U22048 (N_22048,N_17661,N_11782);
nor U22049 (N_22049,N_14436,N_18292);
xnor U22050 (N_22050,N_12865,N_10132);
nor U22051 (N_22051,N_14052,N_17594);
and U22052 (N_22052,N_10388,N_13723);
nor U22053 (N_22053,N_12595,N_19577);
or U22054 (N_22054,N_15253,N_14206);
nand U22055 (N_22055,N_12091,N_10313);
nand U22056 (N_22056,N_16339,N_13377);
xnor U22057 (N_22057,N_11105,N_16489);
or U22058 (N_22058,N_11970,N_17919);
and U22059 (N_22059,N_12366,N_18989);
nand U22060 (N_22060,N_13733,N_16894);
or U22061 (N_22061,N_18863,N_10177);
nand U22062 (N_22062,N_17470,N_15132);
xor U22063 (N_22063,N_11043,N_10894);
xnor U22064 (N_22064,N_17430,N_15327);
nor U22065 (N_22065,N_11710,N_14682);
or U22066 (N_22066,N_11895,N_16865);
nor U22067 (N_22067,N_19025,N_19485);
xnor U22068 (N_22068,N_16079,N_11521);
and U22069 (N_22069,N_13375,N_17213);
and U22070 (N_22070,N_16470,N_15948);
and U22071 (N_22071,N_16544,N_16727);
or U22072 (N_22072,N_10531,N_15645);
xnor U22073 (N_22073,N_15500,N_19713);
nor U22074 (N_22074,N_16689,N_19248);
or U22075 (N_22075,N_13444,N_16438);
nor U22076 (N_22076,N_17250,N_13212);
nor U22077 (N_22077,N_16121,N_19259);
xor U22078 (N_22078,N_17960,N_16888);
xor U22079 (N_22079,N_14140,N_14804);
nor U22080 (N_22080,N_17212,N_12197);
and U22081 (N_22081,N_18805,N_18049);
nor U22082 (N_22082,N_10399,N_16441);
nor U22083 (N_22083,N_10522,N_16844);
nor U22084 (N_22084,N_15520,N_13895);
nand U22085 (N_22085,N_17567,N_13948);
xor U22086 (N_22086,N_13127,N_14432);
nor U22087 (N_22087,N_19241,N_18468);
xor U22088 (N_22088,N_18496,N_12536);
nand U22089 (N_22089,N_19307,N_12799);
and U22090 (N_22090,N_14145,N_14381);
or U22091 (N_22091,N_16753,N_15818);
or U22092 (N_22092,N_18606,N_12394);
xor U22093 (N_22093,N_10623,N_15985);
or U22094 (N_22094,N_19567,N_18588);
xor U22095 (N_22095,N_16146,N_16086);
or U22096 (N_22096,N_17309,N_15598);
nor U22097 (N_22097,N_14452,N_18515);
xor U22098 (N_22098,N_17969,N_13353);
nor U22099 (N_22099,N_10551,N_13806);
nor U22100 (N_22100,N_14057,N_17203);
xnor U22101 (N_22101,N_13038,N_16828);
xnor U22102 (N_22102,N_14891,N_15754);
and U22103 (N_22103,N_10816,N_17887);
or U22104 (N_22104,N_10977,N_12423);
and U22105 (N_22105,N_10385,N_15896);
xnor U22106 (N_22106,N_13072,N_18948);
nand U22107 (N_22107,N_13576,N_18498);
nand U22108 (N_22108,N_16389,N_17910);
and U22109 (N_22109,N_18633,N_17063);
xnor U22110 (N_22110,N_15036,N_10519);
xnor U22111 (N_22111,N_14551,N_16997);
and U22112 (N_22112,N_10574,N_15436);
or U22113 (N_22113,N_12938,N_10691);
xnor U22114 (N_22114,N_12065,N_18938);
xor U22115 (N_22115,N_13741,N_12774);
nor U22116 (N_22116,N_14973,N_17256);
and U22117 (N_22117,N_11979,N_13380);
nor U22118 (N_22118,N_10739,N_11478);
or U22119 (N_22119,N_15770,N_17479);
and U22120 (N_22120,N_18169,N_10166);
nand U22121 (N_22121,N_13129,N_12530);
xor U22122 (N_22122,N_15864,N_17764);
nand U22123 (N_22123,N_12855,N_14732);
nand U22124 (N_22124,N_14927,N_14067);
nand U22125 (N_22125,N_18833,N_19257);
or U22126 (N_22126,N_18358,N_14657);
and U22127 (N_22127,N_12144,N_18594);
or U22128 (N_22128,N_14114,N_14150);
nor U22129 (N_22129,N_12142,N_14796);
xnor U22130 (N_22130,N_12731,N_15493);
nor U22131 (N_22131,N_18836,N_19126);
and U22132 (N_22132,N_17972,N_11833);
nand U22133 (N_22133,N_17150,N_14568);
nand U22134 (N_22134,N_12951,N_13297);
and U22135 (N_22135,N_14620,N_15660);
nor U22136 (N_22136,N_13891,N_14350);
nand U22137 (N_22137,N_19494,N_16735);
nor U22138 (N_22138,N_14664,N_14803);
xnor U22139 (N_22139,N_11092,N_19225);
nor U22140 (N_22140,N_12550,N_15546);
and U22141 (N_22141,N_13156,N_12152);
xor U22142 (N_22142,N_19501,N_15320);
and U22143 (N_22143,N_11509,N_13168);
nand U22144 (N_22144,N_14947,N_17137);
and U22145 (N_22145,N_15688,N_14880);
nor U22146 (N_22146,N_17935,N_18113);
nor U22147 (N_22147,N_19362,N_18552);
nor U22148 (N_22148,N_14136,N_17401);
and U22149 (N_22149,N_19945,N_11633);
nor U22150 (N_22150,N_10763,N_14658);
nor U22151 (N_22151,N_16930,N_12362);
and U22152 (N_22152,N_12227,N_11911);
nor U22153 (N_22153,N_12125,N_18000);
xor U22154 (N_22154,N_12600,N_11031);
and U22155 (N_22155,N_14379,N_10066);
and U22156 (N_22156,N_17778,N_14284);
and U22157 (N_22157,N_17492,N_15957);
nor U22158 (N_22158,N_15855,N_16488);
xor U22159 (N_22159,N_15926,N_10616);
xor U22160 (N_22160,N_15412,N_12119);
and U22161 (N_22161,N_14058,N_14026);
or U22162 (N_22162,N_17095,N_18060);
xor U22163 (N_22163,N_15254,N_19032);
or U22164 (N_22164,N_17875,N_13663);
and U22165 (N_22165,N_11452,N_14115);
xnor U22166 (N_22166,N_11294,N_18305);
nor U22167 (N_22167,N_16760,N_13148);
or U22168 (N_22168,N_17858,N_14749);
nor U22169 (N_22169,N_10571,N_18993);
and U22170 (N_22170,N_10124,N_10954);
xnor U22171 (N_22171,N_11603,N_14061);
xor U22172 (N_22172,N_13519,N_17031);
or U22173 (N_22173,N_14913,N_11975);
or U22174 (N_22174,N_16814,N_14542);
nor U22175 (N_22175,N_11182,N_14717);
and U22176 (N_22176,N_18579,N_16639);
and U22177 (N_22177,N_13884,N_12694);
nand U22178 (N_22178,N_16006,N_14362);
nor U22179 (N_22179,N_17871,N_17554);
or U22180 (N_22180,N_12802,N_14970);
and U22181 (N_22181,N_15187,N_11654);
xnor U22182 (N_22182,N_18450,N_19163);
and U22183 (N_22183,N_14107,N_17641);
nand U22184 (N_22184,N_10225,N_14293);
or U22185 (N_22185,N_12337,N_13448);
or U22186 (N_22186,N_13283,N_12271);
nand U22187 (N_22187,N_17911,N_14171);
nand U22188 (N_22188,N_18321,N_12192);
xnor U22189 (N_22189,N_11430,N_11325);
nor U22190 (N_22190,N_16183,N_16937);
or U22191 (N_22191,N_10356,N_14069);
xor U22192 (N_22192,N_11696,N_14872);
or U22193 (N_22193,N_12924,N_12026);
xnor U22194 (N_22194,N_18269,N_10217);
nor U22195 (N_22195,N_19214,N_17341);
or U22196 (N_22196,N_14940,N_12475);
or U22197 (N_22197,N_17245,N_17102);
xor U22198 (N_22198,N_17934,N_13709);
nand U22199 (N_22199,N_15420,N_10308);
and U22200 (N_22200,N_14932,N_18423);
nand U22201 (N_22201,N_17502,N_12622);
xnor U22202 (N_22202,N_14060,N_18742);
and U22203 (N_22203,N_15396,N_13751);
and U22204 (N_22204,N_18429,N_16237);
nand U22205 (N_22205,N_15003,N_11434);
and U22206 (N_22206,N_11290,N_11006);
nand U22207 (N_22207,N_14585,N_19105);
xnor U22208 (N_22208,N_10061,N_18976);
and U22209 (N_22209,N_11417,N_13388);
or U22210 (N_22210,N_13336,N_11129);
nor U22211 (N_22211,N_12502,N_15828);
and U22212 (N_22212,N_16436,N_10895);
xor U22213 (N_22213,N_13220,N_12473);
nand U22214 (N_22214,N_11868,N_19848);
nand U22215 (N_22215,N_10234,N_13889);
and U22216 (N_22216,N_14832,N_17561);
or U22217 (N_22217,N_11740,N_13265);
xnor U22218 (N_22218,N_16567,N_14999);
nor U22219 (N_22219,N_11422,N_18152);
xnor U22220 (N_22220,N_13422,N_16278);
and U22221 (N_22221,N_10951,N_14291);
or U22222 (N_22222,N_10550,N_19113);
or U22223 (N_22223,N_19480,N_14175);
nor U22224 (N_22224,N_19704,N_15065);
xor U22225 (N_22225,N_13824,N_18677);
nand U22226 (N_22226,N_16064,N_19991);
nand U22227 (N_22227,N_17426,N_12950);
and U22228 (N_22228,N_18256,N_12289);
and U22229 (N_22229,N_10033,N_19712);
or U22230 (N_22230,N_10341,N_15592);
or U22231 (N_22231,N_12795,N_19825);
xnor U22232 (N_22232,N_16286,N_12480);
xor U22233 (N_22233,N_16931,N_17184);
or U22234 (N_22234,N_16964,N_15910);
xor U22235 (N_22235,N_13478,N_18570);
or U22236 (N_22236,N_12253,N_11517);
or U22237 (N_22237,N_19622,N_18022);
and U22238 (N_22238,N_14924,N_18908);
and U22239 (N_22239,N_10729,N_13044);
xor U22240 (N_22240,N_10535,N_19299);
nand U22241 (N_22241,N_10267,N_16255);
or U22242 (N_22242,N_13825,N_15435);
and U22243 (N_22243,N_15402,N_19661);
nand U22244 (N_22244,N_17094,N_14953);
xnor U22245 (N_22245,N_11391,N_15555);
nor U22246 (N_22246,N_14609,N_17640);
or U22247 (N_22247,N_16219,N_13175);
and U22248 (N_22248,N_13144,N_13697);
nor U22249 (N_22249,N_18778,N_13861);
nor U22250 (N_22250,N_16467,N_14883);
nand U22251 (N_22251,N_13051,N_12789);
or U22252 (N_22252,N_11471,N_10621);
and U22253 (N_22253,N_15609,N_17463);
nand U22254 (N_22254,N_18586,N_14962);
nor U22255 (N_22255,N_19314,N_11571);
xnor U22256 (N_22256,N_11054,N_13628);
nor U22257 (N_22257,N_15408,N_15838);
nor U22258 (N_22258,N_11111,N_17854);
nand U22259 (N_22259,N_17948,N_17878);
xor U22260 (N_22260,N_17514,N_17474);
nand U22261 (N_22261,N_16561,N_15643);
or U22262 (N_22262,N_15537,N_18345);
nor U22263 (N_22263,N_14311,N_16777);
nor U22264 (N_22264,N_18476,N_13972);
or U22265 (N_22265,N_12484,N_14995);
nand U22266 (N_22266,N_12072,N_12280);
nand U22267 (N_22267,N_15952,N_13214);
xnor U22268 (N_22268,N_15226,N_13130);
xor U22269 (N_22269,N_16673,N_17652);
nand U22270 (N_22270,N_16324,N_11618);
nor U22271 (N_22271,N_13530,N_17800);
nand U22272 (N_22272,N_10130,N_11926);
or U22273 (N_22273,N_10998,N_16690);
or U22274 (N_22274,N_17145,N_10015);
or U22275 (N_22275,N_15147,N_13197);
and U22276 (N_22276,N_13084,N_17782);
nor U22277 (N_22277,N_15496,N_15152);
and U22278 (N_22278,N_16531,N_12718);
nand U22279 (N_22279,N_19839,N_18177);
nor U22280 (N_22280,N_11059,N_15736);
nand U22281 (N_22281,N_12610,N_10828);
or U22282 (N_22282,N_18787,N_12468);
nand U22283 (N_22283,N_17673,N_15273);
xor U22284 (N_22284,N_18631,N_17506);
and U22285 (N_22285,N_14434,N_11216);
and U22286 (N_22286,N_18403,N_13155);
xnor U22287 (N_22287,N_18531,N_19944);
nand U22288 (N_22288,N_13305,N_11476);
and U22289 (N_22289,N_16720,N_11178);
nand U22290 (N_22290,N_17877,N_18984);
and U22291 (N_22291,N_10362,N_18247);
nand U22292 (N_22292,N_12800,N_13798);
nand U22293 (N_22293,N_17985,N_10568);
xor U22294 (N_22294,N_10506,N_14180);
xor U22295 (N_22295,N_10911,N_11468);
nand U22296 (N_22296,N_17473,N_14164);
or U22297 (N_22297,N_17991,N_14526);
nand U22298 (N_22298,N_14879,N_19950);
xnor U22299 (N_22299,N_10345,N_18470);
nor U22300 (N_22300,N_10440,N_18868);
nand U22301 (N_22301,N_16221,N_18144);
xor U22302 (N_22302,N_13221,N_18394);
nand U22303 (N_22303,N_17298,N_10418);
nand U22304 (N_22304,N_14955,N_13331);
nand U22305 (N_22305,N_15473,N_13584);
xor U22306 (N_22306,N_10758,N_11177);
nand U22307 (N_22307,N_14516,N_12428);
and U22308 (N_22308,N_13583,N_15515);
xnor U22309 (N_22309,N_11263,N_16556);
nand U22310 (N_22310,N_13255,N_13986);
xor U22311 (N_22311,N_16502,N_14054);
or U22312 (N_22312,N_11939,N_18025);
or U22313 (N_22313,N_17411,N_14288);
or U22314 (N_22314,N_17884,N_16308);
nor U22315 (N_22315,N_19419,N_10269);
or U22316 (N_22316,N_18774,N_11328);
and U22317 (N_22317,N_16879,N_14081);
nor U22318 (N_22318,N_14966,N_19861);
nand U22319 (N_22319,N_12982,N_17490);
and U22320 (N_22320,N_10274,N_12353);
xnor U22321 (N_22321,N_14644,N_18700);
nand U22322 (N_22322,N_16437,N_19079);
or U22323 (N_22323,N_12005,N_11973);
and U22324 (N_22324,N_11450,N_12497);
and U22325 (N_22325,N_18271,N_18407);
xnor U22326 (N_22326,N_16400,N_12451);
or U22327 (N_22327,N_11860,N_12434);
or U22328 (N_22328,N_15359,N_19034);
and U22329 (N_22329,N_13273,N_17515);
nor U22330 (N_22330,N_15304,N_11021);
or U22331 (N_22331,N_18106,N_13302);
nor U22332 (N_22332,N_19053,N_13514);
or U22333 (N_22333,N_10370,N_11592);
xnor U22334 (N_22334,N_18259,N_13001);
nor U22335 (N_22335,N_10606,N_12647);
xnor U22336 (N_22336,N_17233,N_14385);
nand U22337 (N_22337,N_15856,N_18183);
or U22338 (N_22338,N_15796,N_14772);
or U22339 (N_22339,N_15465,N_10285);
xnor U22340 (N_22340,N_15432,N_16377);
xnor U22341 (N_22341,N_10318,N_13843);
or U22342 (N_22342,N_13516,N_12311);
or U22343 (N_22343,N_14229,N_19076);
or U22344 (N_22344,N_15759,N_18831);
and U22345 (N_22345,N_10626,N_11209);
nand U22346 (N_22346,N_16557,N_11261);
or U22347 (N_22347,N_10707,N_13109);
nor U22348 (N_22348,N_13869,N_10678);
nand U22349 (N_22349,N_16914,N_19871);
nor U22350 (N_22350,N_16742,N_13594);
nand U22351 (N_22351,N_13896,N_18914);
nor U22352 (N_22352,N_16283,N_14384);
nand U22353 (N_22353,N_12117,N_18815);
nor U22354 (N_22354,N_11889,N_15119);
and U22355 (N_22355,N_14465,N_18372);
nor U22356 (N_22356,N_16802,N_13705);
or U22357 (N_22357,N_19431,N_18615);
or U22358 (N_22358,N_15790,N_13241);
and U22359 (N_22359,N_18731,N_17885);
and U22360 (N_22360,N_18617,N_18486);
xnor U22361 (N_22361,N_19456,N_12308);
and U22362 (N_22362,N_11921,N_14554);
nor U22363 (N_22363,N_17982,N_19440);
nand U22364 (N_22364,N_14354,N_11331);
nand U22365 (N_22365,N_16499,N_16432);
and U22366 (N_22366,N_12604,N_11600);
and U22367 (N_22367,N_12040,N_10696);
or U22368 (N_22368,N_14166,N_15374);
and U22369 (N_22369,N_16650,N_13920);
and U22370 (N_22370,N_15084,N_17703);
and U22371 (N_22371,N_19358,N_16217);
and U22372 (N_22372,N_19983,N_15252);
nand U22373 (N_22373,N_19478,N_13913);
and U22374 (N_22374,N_14022,N_16428);
nand U22375 (N_22375,N_17498,N_19956);
nor U22376 (N_22376,N_14636,N_15366);
xnor U22377 (N_22377,N_11283,N_12209);
nand U22378 (N_22378,N_11981,N_15035);
or U22379 (N_22379,N_14733,N_12232);
xnor U22380 (N_22380,N_17366,N_13634);
xor U22381 (N_22381,N_18530,N_13636);
nand U22382 (N_22382,N_12693,N_19613);
nand U22383 (N_22383,N_12448,N_15883);
or U22384 (N_22384,N_19572,N_16495);
and U22385 (N_22385,N_10593,N_19158);
and U22386 (N_22386,N_16139,N_14196);
nand U22387 (N_22387,N_15602,N_15221);
and U22388 (N_22388,N_17698,N_15441);
and U22389 (N_22389,N_11268,N_14297);
nor U22390 (N_22390,N_14451,N_13201);
or U22391 (N_22391,N_10815,N_18522);
and U22392 (N_22392,N_16630,N_19813);
xnor U22393 (N_22393,N_10871,N_15251);
or U22394 (N_22394,N_15179,N_15332);
or U22395 (N_22395,N_16800,N_17761);
nand U22396 (N_22396,N_13827,N_17436);
nor U22397 (N_22397,N_16540,N_11540);
or U22398 (N_22398,N_15961,N_18401);
nand U22399 (N_22399,N_16984,N_12631);
xor U22400 (N_22400,N_11713,N_15677);
and U22401 (N_22401,N_14739,N_13110);
and U22402 (N_22402,N_18129,N_10920);
xor U22403 (N_22403,N_13714,N_11831);
xor U22404 (N_22404,N_13364,N_13386);
xor U22405 (N_22405,N_12740,N_15092);
or U22406 (N_22406,N_18011,N_16589);
xnor U22407 (N_22407,N_16677,N_13822);
or U22408 (N_22408,N_13907,N_13924);
xor U22409 (N_22409,N_15347,N_16897);
or U22410 (N_22410,N_10556,N_16093);
nand U22411 (N_22411,N_14660,N_19308);
or U22412 (N_22412,N_19455,N_15082);
nor U22413 (N_22413,N_17612,N_14784);
nand U22414 (N_22414,N_11992,N_16052);
or U22415 (N_22415,N_13816,N_10118);
nand U22416 (N_22416,N_17995,N_17400);
nor U22417 (N_22417,N_18917,N_14545);
xnor U22418 (N_22418,N_13095,N_19789);
nor U22419 (N_22419,N_18361,N_17014);
nor U22420 (N_22420,N_12851,N_16128);
and U22421 (N_22421,N_18233,N_13055);
and U22422 (N_22422,N_19153,N_15005);
xor U22423 (N_22423,N_15559,N_18758);
and U22424 (N_22424,N_17795,N_17160);
nor U22425 (N_22425,N_15370,N_13916);
nand U22426 (N_22426,N_15562,N_11819);
nor U22427 (N_22427,N_13159,N_14223);
nand U22428 (N_22428,N_11711,N_11955);
nor U22429 (N_22429,N_13136,N_18883);
nand U22430 (N_22430,N_10205,N_13254);
nand U22431 (N_22431,N_15235,N_19838);
xnor U22432 (N_22432,N_13340,N_15437);
and U22433 (N_22433,N_17734,N_19351);
nor U22434 (N_22434,N_18300,N_19296);
nand U22435 (N_22435,N_15348,N_13190);
xnor U22436 (N_22436,N_10239,N_10446);
or U22437 (N_22437,N_12100,N_13125);
nand U22438 (N_22438,N_11985,N_10903);
and U22439 (N_22439,N_19066,N_16831);
or U22440 (N_22440,N_18170,N_10021);
nand U22441 (N_22441,N_16761,N_18206);
or U22442 (N_22442,N_10776,N_17721);
nor U22443 (N_22443,N_14814,N_10737);
xor U22444 (N_22444,N_18595,N_14552);
and U22445 (N_22445,N_16573,N_13151);
nor U22446 (N_22446,N_11681,N_10743);
nand U22447 (N_22447,N_17439,N_19474);
nand U22448 (N_22448,N_19561,N_17068);
nor U22449 (N_22449,N_11274,N_11780);
or U22450 (N_22450,N_19273,N_19780);
nor U22451 (N_22451,N_13394,N_17713);
xor U22452 (N_22452,N_18565,N_15274);
and U22453 (N_22453,N_10223,N_14588);
nand U22454 (N_22454,N_14697,N_13017);
xnor U22455 (N_22455,N_12120,N_19747);
or U22456 (N_22456,N_19233,N_10644);
and U22457 (N_22457,N_13258,N_18274);
nor U22458 (N_22458,N_16353,N_13032);
xor U22459 (N_22459,N_11532,N_19811);
xor U22460 (N_22460,N_18811,N_15062);
nor U22461 (N_22461,N_17825,N_15521);
and U22462 (N_22462,N_12818,N_15301);
nand U22463 (N_22463,N_17376,N_12160);
nor U22464 (N_22464,N_12094,N_19352);
or U22465 (N_22465,N_18245,N_11098);
xnor U22466 (N_22466,N_12878,N_17382);
and U22467 (N_22467,N_12214,N_18807);
xnor U22468 (N_22468,N_15194,N_11012);
nor U22469 (N_22469,N_18424,N_11866);
xor U22470 (N_22470,N_11300,N_15817);
nand U22471 (N_22471,N_14444,N_16223);
nand U22472 (N_22472,N_16153,N_19926);
and U22473 (N_22473,N_14499,N_13987);
nand U22474 (N_22474,N_19184,N_15056);
nor U22475 (N_22475,N_17264,N_11273);
and U22476 (N_22476,N_14008,N_12861);
and U22477 (N_22477,N_15925,N_10381);
and U22478 (N_22478,N_15571,N_12611);
nor U22479 (N_22479,N_16551,N_18162);
nor U22480 (N_22480,N_15815,N_19834);
nand U22481 (N_22481,N_11337,N_13955);
or U22482 (N_22482,N_19828,N_17741);
and U22483 (N_22483,N_16152,N_12547);
or U22484 (N_22484,N_16536,N_17471);
or U22485 (N_22485,N_11645,N_16929);
xnor U22486 (N_22486,N_15748,N_11011);
or U22487 (N_22487,N_11535,N_18356);
and U22488 (N_22488,N_15182,N_17385);
or U22489 (N_22489,N_11408,N_13988);
nor U22490 (N_22490,N_15210,N_18124);
xor U22491 (N_22491,N_14626,N_14801);
and U22492 (N_22492,N_19088,N_14041);
nand U22493 (N_22493,N_19630,N_11457);
nand U22494 (N_22494,N_10219,N_13828);
and U22495 (N_22495,N_14519,N_16620);
nor U22496 (N_22496,N_15750,N_11894);
and U22497 (N_22497,N_12669,N_17308);
or U22498 (N_22498,N_15935,N_10813);
nor U22499 (N_22499,N_11703,N_11454);
nand U22500 (N_22500,N_16458,N_18744);
nand U22501 (N_22501,N_16197,N_19396);
or U22502 (N_22502,N_14027,N_17895);
or U22503 (N_22503,N_10702,N_19295);
and U22504 (N_22504,N_12873,N_14662);
and U22505 (N_22505,N_14017,N_14613);
or U22506 (N_22506,N_14726,N_12856);
nor U22507 (N_22507,N_15606,N_15649);
and U22508 (N_22508,N_16100,N_19992);
xor U22509 (N_22509,N_18528,N_10502);
xnor U22510 (N_22510,N_16804,N_16165);
nor U22511 (N_22511,N_10787,N_19020);
or U22512 (N_22512,N_12685,N_14199);
nand U22513 (N_22513,N_14853,N_12383);
xnor U22514 (N_22514,N_16921,N_18436);
nand U22515 (N_22515,N_12869,N_15853);
or U22516 (N_22516,N_18502,N_14260);
xnor U22517 (N_22517,N_16455,N_18776);
or U22518 (N_22518,N_18048,N_11137);
and U22519 (N_22519,N_16322,N_18759);
nand U22520 (N_22520,N_17135,N_13524);
nand U22521 (N_22521,N_13249,N_13281);
and U22522 (N_22522,N_13181,N_18664);
or U22523 (N_22523,N_17657,N_13795);
or U22524 (N_22524,N_15539,N_10836);
nand U22525 (N_22525,N_19261,N_17847);
nor U22526 (N_22526,N_13266,N_11668);
nor U22527 (N_22527,N_15480,N_14599);
or U22528 (N_22528,N_14711,N_12112);
nor U22529 (N_22529,N_13931,N_12608);
nor U22530 (N_22530,N_10625,N_17152);
or U22531 (N_22531,N_13108,N_11963);
and U22532 (N_22532,N_12675,N_14258);
and U22533 (N_22533,N_15584,N_19619);
nor U22534 (N_22534,N_12603,N_18887);
or U22535 (N_22535,N_11078,N_15728);
nor U22536 (N_22536,N_18395,N_15100);
or U22537 (N_22537,N_12470,N_16081);
nand U22538 (N_22538,N_15870,N_13739);
xor U22539 (N_22539,N_10869,N_18790);
nor U22540 (N_22540,N_19266,N_12888);
and U22541 (N_22541,N_19788,N_14083);
nand U22542 (N_22542,N_14365,N_16048);
xor U22543 (N_22543,N_18262,N_10314);
or U22544 (N_22544,N_16714,N_12011);
nand U22545 (N_22545,N_16909,N_17027);
or U22546 (N_22546,N_13274,N_12716);
and U22547 (N_22547,N_13747,N_12398);
or U22548 (N_22548,N_16487,N_15992);
xor U22549 (N_22549,N_12711,N_16402);
and U22550 (N_22550,N_17409,N_11957);
nor U22551 (N_22551,N_13725,N_18117);
nand U22552 (N_22552,N_14678,N_13712);
or U22553 (N_22553,N_10893,N_10741);
and U22554 (N_22554,N_18052,N_18364);
or U22555 (N_22555,N_12440,N_14630);
or U22556 (N_22556,N_19312,N_13404);
or U22557 (N_22557,N_13846,N_10143);
and U22558 (N_22558,N_13831,N_15478);
xnor U22559 (N_22559,N_18384,N_15167);
and U22560 (N_22560,N_19144,N_10558);
or U22561 (N_22561,N_11191,N_10536);
xnor U22562 (N_22562,N_13403,N_16230);
nand U22563 (N_22563,N_18145,N_18329);
xor U22564 (N_22564,N_16975,N_10981);
nand U22565 (N_22565,N_10214,N_15579);
nand U22566 (N_22566,N_13204,N_12926);
nor U22567 (N_22567,N_10566,N_14062);
or U22568 (N_22568,N_10271,N_12572);
or U22569 (N_22569,N_18323,N_16948);
or U22570 (N_22570,N_19211,N_15561);
or U22571 (N_22571,N_16078,N_10404);
xnor U22572 (N_22572,N_13233,N_10802);
nand U22573 (N_22573,N_15418,N_18076);
nand U22574 (N_22574,N_15565,N_19741);
xnor U22575 (N_22575,N_13648,N_14262);
or U22576 (N_22576,N_13169,N_10336);
and U22577 (N_22577,N_14307,N_10872);
nor U22578 (N_22578,N_19316,N_11608);
xnor U22579 (N_22579,N_16107,N_12979);
nand U22580 (N_22580,N_15731,N_16386);
and U22581 (N_22581,N_17966,N_12171);
nand U22582 (N_22582,N_11903,N_15277);
and U22583 (N_22583,N_15740,N_16808);
xor U22584 (N_22584,N_18800,N_19599);
nor U22585 (N_22585,N_16295,N_13601);
xor U22586 (N_22586,N_12349,N_12663);
nand U22587 (N_22587,N_11170,N_10859);
nand U22588 (N_22588,N_14386,N_17389);
xor U22589 (N_22589,N_14529,N_12654);
xor U22590 (N_22590,N_19167,N_13719);
xnor U22591 (N_22591,N_15111,N_16586);
or U22592 (N_22592,N_17757,N_15073);
xnor U22593 (N_22593,N_12525,N_16552);
xor U22594 (N_22594,N_11938,N_18353);
nor U22595 (N_22595,N_17017,N_14398);
xnor U22596 (N_22596,N_17169,N_10439);
xnor U22597 (N_22597,N_10379,N_12884);
nand U22598 (N_22598,N_14761,N_18244);
and U22599 (N_22599,N_17743,N_19205);
or U22600 (N_22600,N_18404,N_10243);
nand U22601 (N_22601,N_12966,N_18918);
nor U22602 (N_22602,N_16313,N_12521);
nor U22603 (N_22603,N_18567,N_14072);
or U22604 (N_22604,N_12766,N_16443);
xnor U22605 (N_22605,N_16158,N_18842);
nand U22606 (N_22606,N_15052,N_18422);
nand U22607 (N_22607,N_12445,N_18132);
xnor U22608 (N_22608,N_12698,N_12274);
xor U22609 (N_22609,N_19924,N_16185);
nor U22610 (N_22610,N_10814,N_12822);
or U22611 (N_22611,N_12657,N_17208);
nor U22612 (N_22612,N_18599,N_11246);
nor U22613 (N_22613,N_16506,N_13368);
or U22614 (N_22614,N_17097,N_12089);
and U22615 (N_22615,N_13370,N_16507);
and U22616 (N_22616,N_15078,N_15834);
nor U22617 (N_22617,N_12915,N_17484);
or U22618 (N_22618,N_16528,N_14665);
nand U22619 (N_22619,N_19753,N_11851);
xnor U22620 (N_22620,N_14267,N_10655);
nand U22621 (N_22621,N_11020,N_19070);
and U22622 (N_22622,N_16417,N_14989);
nor U22623 (N_22623,N_14111,N_10862);
nor U22624 (N_22624,N_11279,N_13133);
nand U22625 (N_22625,N_16229,N_10994);
nand U22626 (N_22626,N_17898,N_17177);
or U22627 (N_22627,N_14153,N_14791);
nor U22628 (N_22628,N_19797,N_13277);
or U22629 (N_22629,N_13395,N_14980);
or U22630 (N_22630,N_12381,N_18110);
and U22631 (N_22631,N_10068,N_12333);
and U22632 (N_22632,N_11716,N_13124);
and U22633 (N_22633,N_11809,N_17904);
nor U22634 (N_22634,N_16046,N_16605);
or U22635 (N_22635,N_11873,N_11469);
xnor U22636 (N_22636,N_15373,N_15428);
nand U22637 (N_22637,N_16674,N_16664);
xor U22638 (N_22638,N_16509,N_10923);
xnor U22639 (N_22639,N_19170,N_10665);
or U22640 (N_22640,N_10500,N_17678);
xor U22641 (N_22641,N_10003,N_12003);
or U22642 (N_22642,N_12649,N_19565);
nor U22643 (N_22643,N_17270,N_17272);
or U22644 (N_22644,N_11488,N_12002);
or U22645 (N_22645,N_19137,N_12725);
nor U22646 (N_22646,N_14888,N_19049);
nor U22647 (N_22647,N_17790,N_18050);
xor U22648 (N_22648,N_14018,N_14372);
and U22649 (N_22649,N_18683,N_19786);
nor U22650 (N_22650,N_11438,N_17190);
or U22651 (N_22651,N_19898,N_10775);
nand U22652 (N_22652,N_12248,N_17251);
or U22653 (N_22653,N_12151,N_16423);
and U22654 (N_22654,N_11360,N_10538);
nand U22655 (N_22655,N_14032,N_19092);
and U22656 (N_22656,N_12340,N_14119);
and U22657 (N_22657,N_18490,N_12650);
nand U22658 (N_22658,N_17228,N_11442);
xnor U22659 (N_22659,N_11386,N_10218);
and U22660 (N_22660,N_17252,N_16919);
or U22661 (N_22661,N_19473,N_15361);
and U22662 (N_22662,N_18477,N_19279);
or U22663 (N_22663,N_18159,N_11260);
xor U22664 (N_22664,N_18963,N_17989);
or U22665 (N_22665,N_16672,N_12637);
nor U22666 (N_22666,N_10740,N_16651);
and U22667 (N_22667,N_11604,N_19365);
nand U22668 (N_22668,N_10287,N_14771);
nor U22669 (N_22669,N_10006,N_11983);
or U22670 (N_22670,N_17816,N_14612);
and U22671 (N_22671,N_16980,N_12326);
nor U22672 (N_22672,N_13443,N_15393);
and U22673 (N_22673,N_16758,N_18315);
xnor U22674 (N_22674,N_17917,N_16559);
and U22675 (N_22675,N_11995,N_18931);
nor U22676 (N_22676,N_19717,N_15720);
nand U22677 (N_22677,N_11210,N_18243);
nand U22678 (N_22678,N_15893,N_18027);
nor U22679 (N_22679,N_19783,N_19277);
nor U22680 (N_22680,N_15072,N_18009);
nand U22681 (N_22681,N_11219,N_15113);
and U22682 (N_22682,N_14712,N_17077);
xnor U22683 (N_22683,N_14725,N_17444);
or U22684 (N_22684,N_14910,N_16604);
nand U22685 (N_22685,N_19726,N_10902);
and U22686 (N_22686,N_14217,N_11108);
nand U22687 (N_22687,N_12254,N_16613);
and U22688 (N_22688,N_11658,N_14720);
nor U22689 (N_22689,N_11516,N_14921);
nand U22690 (N_22690,N_16272,N_12009);
xor U22691 (N_22691,N_10577,N_12720);
nand U22692 (N_22692,N_19590,N_12705);
nand U22693 (N_22693,N_14407,N_19679);
nor U22694 (N_22694,N_14323,N_13529);
or U22695 (N_22695,N_17259,N_11244);
nand U22696 (N_22696,N_14134,N_12936);
nor U22697 (N_22697,N_17873,N_13867);
nor U22698 (N_22698,N_11572,N_19833);
and U22699 (N_22699,N_10541,N_16617);
nand U22700 (N_22700,N_14705,N_18376);
xor U22701 (N_22701,N_17799,N_14141);
or U22702 (N_22702,N_14933,N_11676);
xor U22703 (N_22703,N_17274,N_13661);
nand U22704 (N_22704,N_16876,N_19691);
nand U22705 (N_22705,N_17719,N_14789);
and U22706 (N_22706,N_11225,N_10262);
and U22707 (N_22707,N_14342,N_16757);
nand U22708 (N_22708,N_16663,N_10194);
nand U22709 (N_22709,N_10701,N_14673);
or U22710 (N_22710,N_17831,N_16730);
and U22711 (N_22711,N_17819,N_11812);
xnor U22712 (N_22712,N_17848,N_11302);
nor U22713 (N_22713,N_11974,N_18537);
nor U22714 (N_22714,N_16019,N_10331);
or U22715 (N_22715,N_13771,N_11160);
or U22716 (N_22716,N_18894,N_17670);
or U22717 (N_22717,N_18584,N_15117);
nand U22718 (N_22718,N_13504,N_14183);
xnor U22719 (N_22719,N_12414,N_18462);
nand U22720 (N_22720,N_19645,N_17078);
and U22721 (N_22721,N_16480,N_18004);
xnor U22722 (N_22722,N_17231,N_15679);
or U22723 (N_22723,N_19289,N_15467);
nor U22724 (N_22724,N_19288,N_13958);
and U22725 (N_22725,N_17101,N_18650);
nand U22726 (N_22726,N_12081,N_17349);
xor U22727 (N_22727,N_11625,N_15708);
xor U22728 (N_22728,N_11484,N_16491);
or U22729 (N_22729,N_10204,N_19769);
nand U22730 (N_22730,N_11599,N_14172);
and U22731 (N_22731,N_18306,N_19465);
or U22732 (N_22732,N_12158,N_16688);
nand U22733 (N_22733,N_19192,N_11069);
xor U22734 (N_22734,N_19350,N_10055);
nand U22735 (N_22735,N_13292,N_19638);
nor U22736 (N_22736,N_13075,N_18006);
xor U22737 (N_22737,N_19017,N_11284);
nand U22738 (N_22738,N_11752,N_12017);
nor U22739 (N_22739,N_11188,N_14729);
or U22740 (N_22740,N_17518,N_11475);
or U22741 (N_22741,N_14458,N_11762);
nand U22742 (N_22742,N_18444,N_14945);
xor U22743 (N_22743,N_10329,N_12234);
xnor U22744 (N_22744,N_17265,N_18485);
xnor U22745 (N_22745,N_16935,N_11295);
or U22746 (N_22746,N_17099,N_11052);
nor U22747 (N_22747,N_10853,N_10378);
or U22748 (N_22748,N_19841,N_15814);
nand U22749 (N_22749,N_14468,N_15652);
xnor U22750 (N_22750,N_10419,N_11091);
and U22751 (N_22751,N_16304,N_18532);
and U22752 (N_22752,N_19059,N_12500);
or U22753 (N_22753,N_14314,N_15678);
and U22754 (N_22754,N_11113,N_15105);
and U22755 (N_22755,N_14413,N_11546);
nor U22756 (N_22756,N_16680,N_13505);
xor U22757 (N_22757,N_10968,N_15590);
xor U22758 (N_22758,N_14269,N_17598);
nand U22759 (N_22759,N_10241,N_16383);
xnor U22760 (N_22760,N_13455,N_18973);
xor U22761 (N_22761,N_15808,N_19243);
and U22762 (N_22762,N_16419,N_16874);
or U22763 (N_22763,N_10099,N_18392);
or U22764 (N_22764,N_19598,N_17023);
or U22765 (N_22765,N_19706,N_14219);
and U22766 (N_22766,N_10931,N_13550);
and U22767 (N_22767,N_18957,N_14868);
nor U22768 (N_22768,N_17627,N_10978);
or U22769 (N_22769,N_18481,N_11241);
or U22770 (N_22770,N_18871,N_19387);
and U22771 (N_22771,N_12131,N_17297);
xor U22772 (N_22772,N_16083,N_17173);
xor U22773 (N_22773,N_16863,N_15446);
nor U22774 (N_22774,N_18651,N_10847);
nor U22775 (N_22775,N_19338,N_19836);
and U22776 (N_22776,N_18459,N_19437);
xnor U22777 (N_22777,N_18822,N_17059);
xnor U22778 (N_22778,N_16738,N_12139);
or U22779 (N_22779,N_16609,N_10669);
xor U22780 (N_22780,N_13352,N_13065);
nand U22781 (N_22781,N_15330,N_16771);
or U22782 (N_22782,N_11997,N_14001);
nand U22783 (N_22783,N_16036,N_19183);
nand U22784 (N_22784,N_19155,N_11107);
and U22785 (N_22785,N_16192,N_16977);
xor U22786 (N_22786,N_16873,N_13330);
or U22787 (N_22787,N_14363,N_18471);
and U22788 (N_22788,N_19947,N_11258);
or U22789 (N_22789,N_10709,N_15115);
xor U22790 (N_22790,N_11035,N_19631);
and U22791 (N_22791,N_12007,N_11612);
nor U22792 (N_22792,N_17792,N_13817);
nand U22793 (N_22793,N_13374,N_12177);
nor U22794 (N_22794,N_15010,N_16481);
and U22795 (N_22795,N_12438,N_13588);
xnor U22796 (N_22796,N_15755,N_16792);
and U22797 (N_22797,N_18719,N_11007);
nand U22798 (N_22798,N_14683,N_19854);
nor U22799 (N_22799,N_15098,N_14528);
xor U22800 (N_22800,N_13429,N_14574);
and U22801 (N_22801,N_17974,N_18010);
nand U22802 (N_22802,N_18970,N_14162);
nand U22803 (N_22803,N_15685,N_11649);
nand U22804 (N_22804,N_18453,N_19282);
and U22805 (N_22805,N_11843,N_17284);
nor U22806 (N_22806,N_13506,N_14874);
nand U22807 (N_22807,N_18249,N_12576);
or U22808 (N_22808,N_17163,N_11980);
nor U22809 (N_22809,N_13288,N_15070);
nand U22810 (N_22810,N_16023,N_15380);
xor U22811 (N_22811,N_14770,N_13473);
nand U22812 (N_22812,N_13818,N_14522);
nor U22813 (N_22813,N_11373,N_18085);
nand U22814 (N_22814,N_12624,N_14068);
xnor U22815 (N_22815,N_18721,N_11041);
or U22816 (N_22816,N_10119,N_16824);
nand U22817 (N_22817,N_15400,N_11080);
xor U22818 (N_22818,N_18513,N_17254);
nand U22819 (N_22819,N_14948,N_13910);
xnor U22820 (N_22820,N_16798,N_12172);
or U22821 (N_22821,N_13820,N_19258);
xor U22822 (N_22822,N_19186,N_19324);
nor U22823 (N_22823,N_17921,N_17729);
or U22824 (N_22824,N_19107,N_18703);
or U22825 (N_22825,N_17714,N_17965);
nor U22826 (N_22826,N_14780,N_17139);
and U22827 (N_22827,N_14696,N_10608);
and U22828 (N_22828,N_10298,N_17520);
nand U22829 (N_22829,N_17956,N_14890);
and U22830 (N_22830,N_19675,N_15950);
and U22831 (N_22831,N_17199,N_10042);
nand U22832 (N_22832,N_14045,N_18663);
and U22833 (N_22833,N_13754,N_15846);
and U22834 (N_22834,N_11948,N_12514);
or U22835 (N_22835,N_15991,N_12013);
and U22836 (N_22836,N_10540,N_17277);
nand U22837 (N_22837,N_10685,N_19201);
and U22838 (N_22838,N_14855,N_19957);
or U22839 (N_22839,N_17756,N_19453);
nand U22840 (N_22840,N_16094,N_12934);
nand U22841 (N_22841,N_12503,N_16268);
nor U22842 (N_22842,N_11732,N_10526);
and U22843 (N_22843,N_13157,N_18197);
xor U22844 (N_22844,N_11315,N_16250);
nand U22845 (N_22845,N_19364,N_11789);
nand U22846 (N_22846,N_13459,N_17933);
nand U22847 (N_22847,N_19551,N_19210);
and U22848 (N_22848,N_17340,N_18383);
or U22849 (N_22849,N_17153,N_19777);
or U22850 (N_22850,N_18137,N_15220);
or U22851 (N_22851,N_11881,N_16037);
xor U22852 (N_22852,N_10967,N_11063);
and U22853 (N_22853,N_11118,N_10613);
and U22854 (N_22854,N_10164,N_15779);
nand U22855 (N_22855,N_19269,N_18185);
nand U22856 (N_22856,N_10706,N_12910);
or U22857 (N_22857,N_13564,N_13239);
and U22858 (N_22858,N_17092,N_13847);
nor U22859 (N_22859,N_14010,N_11636);
and U22860 (N_22860,N_15492,N_13724);
nand U22861 (N_22861,N_11858,N_13812);
nand U22862 (N_22862,N_16145,N_14756);
nor U22863 (N_22863,N_10059,N_19772);
or U22864 (N_22864,N_12348,N_14641);
and U22865 (N_22865,N_19432,N_18198);
xnor U22866 (N_22866,N_18489,N_13362);
and U22867 (N_22867,N_19497,N_19026);
or U22868 (N_22868,N_11168,N_11480);
xnor U22869 (N_22869,N_17326,N_15737);
and U22870 (N_22870,N_14316,N_12409);
nand U22871 (N_22871,N_19935,N_16408);
nor U22872 (N_22872,N_18643,N_18217);
nand U22873 (N_22873,N_16054,N_18302);
and U22874 (N_22874,N_18370,N_17383);
xnor U22875 (N_22875,N_13259,N_17927);
xor U22876 (N_22876,N_16939,N_15108);
nand U22877 (N_22877,N_11723,N_12444);
and U22878 (N_22878,N_17457,N_11487);
and U22879 (N_22879,N_18042,N_11272);
xnor U22880 (N_22880,N_10100,N_19891);
xor U22881 (N_22881,N_16508,N_18281);
and U22882 (N_22882,N_10642,N_15474);
or U22883 (N_22883,N_12971,N_13710);
and U22884 (N_22884,N_13323,N_19104);
nor U22885 (N_22885,N_18521,N_18319);
nand U22886 (N_22886,N_10240,N_12917);
and U22887 (N_22887,N_14816,N_16928);
nand U22888 (N_22888,N_16736,N_19536);
and U22889 (N_22889,N_13953,N_17901);
nor U22890 (N_22890,N_10398,N_13961);
and U22891 (N_22891,N_10071,N_11742);
xor U22892 (N_22892,N_15578,N_17431);
nand U22893 (N_22893,N_18493,N_19809);
xor U22894 (N_22894,N_16934,N_16739);
and U22895 (N_22895,N_15516,N_13613);
xor U22896 (N_22896,N_15914,N_18652);
nor U22897 (N_22897,N_14034,N_19064);
and U22898 (N_22898,N_17551,N_18094);
xnor U22899 (N_22899,N_19881,N_17216);
or U22900 (N_22900,N_15573,N_15405);
or U22901 (N_22901,N_11986,N_16399);
nand U22902 (N_22902,N_18312,N_17141);
and U22903 (N_22903,N_15129,N_12543);
nor U22904 (N_22904,N_15012,N_15654);
and U22905 (N_22905,N_13791,N_17556);
or U22906 (N_22906,N_16915,N_13778);
nor U22907 (N_22907,N_13940,N_16694);
nand U22908 (N_22908,N_19748,N_18203);
nand U22909 (N_22909,N_15994,N_15581);
nor U22910 (N_22910,N_11280,N_10947);
nor U22911 (N_22911,N_15548,N_14116);
xor U22912 (N_22912,N_17826,N_16887);
or U22913 (N_22913,N_11023,N_12487);
xnor U22914 (N_22914,N_19493,N_10746);
and U22915 (N_22915,N_12025,N_18625);
and U22916 (N_22916,N_19682,N_14572);
xor U22917 (N_22917,N_16785,N_18761);
xor U22918 (N_22918,N_19003,N_14992);
nand U22919 (N_22919,N_16682,N_10077);
nand U22920 (N_22920,N_11148,N_15009);
xnor U22921 (N_22921,N_19505,N_10319);
or U22922 (N_22922,N_19707,N_16119);
nor U22923 (N_22923,N_10195,N_12963);
and U22924 (N_22924,N_18550,N_12671);
nand U22925 (N_22925,N_14797,N_18888);
nor U22926 (N_22926,N_15713,N_11888);
or U22927 (N_22927,N_17086,N_12295);
and U22928 (N_22928,N_13568,N_14251);
or U22929 (N_22929,N_14869,N_18046);
and U22930 (N_22930,N_13269,N_17499);
nor U22931 (N_22931,N_18220,N_17220);
or U22932 (N_22932,N_12379,N_15831);
and U22933 (N_22933,N_17944,N_18122);
and U22934 (N_22934,N_18875,N_11639);
and U22935 (N_22935,N_17628,N_17856);
nand U22936 (N_22936,N_19751,N_18400);
nand U22937 (N_22937,N_19961,N_14675);
nor U22938 (N_22938,N_12132,N_16660);
nand U22939 (N_22939,N_16707,N_19830);
and U22940 (N_22940,N_18304,N_13160);
and U22941 (N_22941,N_15684,N_10392);
or U22942 (N_22942,N_15822,N_12684);
and U22943 (N_22943,N_14424,N_17116);
nor U22944 (N_22944,N_19575,N_11934);
or U22945 (N_22945,N_19734,N_14594);
nor U22946 (N_22946,N_12236,N_16870);
and U22947 (N_22947,N_17601,N_19868);
xnor U22948 (N_22948,N_12619,N_18134);
xor U22949 (N_22949,N_10211,N_13753);
or U22950 (N_22950,N_10654,N_19876);
nand U22951 (N_22951,N_10880,N_12060);
xor U22952 (N_22952,N_11176,N_11861);
or U22953 (N_22953,N_14748,N_10515);
nand U22954 (N_22954,N_19345,N_11251);
and U22955 (N_22955,N_12899,N_18558);
nor U22956 (N_22956,N_17684,N_14827);
xnor U22957 (N_22957,N_11365,N_13625);
and U22958 (N_22958,N_10493,N_16198);
nand U22959 (N_22959,N_19095,N_19670);
or U22960 (N_22960,N_16251,N_10823);
nand U22961 (N_22961,N_13235,N_17600);
nor U22962 (N_22962,N_18234,N_12680);
nand U22963 (N_22963,N_15593,N_19344);
nand U22964 (N_22964,N_19147,N_18497);
nand U22965 (N_22965,N_18178,N_12757);
and U22966 (N_22966,N_14807,N_15620);
and U22967 (N_22967,N_13431,N_18686);
xor U22968 (N_22968,N_11115,N_12996);
xnor U22969 (N_22969,N_14253,N_12085);
xnor U22970 (N_22970,N_13068,N_12706);
and U22971 (N_22971,N_17435,N_13457);
nand U22972 (N_22972,N_19200,N_17398);
nand U22973 (N_22973,N_14563,N_18964);
or U22974 (N_22974,N_17338,N_16593);
nor U22975 (N_22975,N_15449,N_11560);
or U22976 (N_22976,N_19875,N_13033);
or U22977 (N_22977,N_13232,N_17072);
or U22978 (N_22978,N_14370,N_19767);
and U22979 (N_22979,N_12155,N_19989);
xor U22980 (N_22980,N_16292,N_14345);
or U22981 (N_22981,N_14155,N_10101);
nor U22982 (N_22982,N_15419,N_10945);
or U22983 (N_22983,N_18821,N_17542);
nand U22984 (N_22984,N_10157,N_15995);
nand U22985 (N_22985,N_13834,N_17073);
nor U22986 (N_22986,N_19228,N_16807);
xnor U22987 (N_22987,N_12724,N_15825);
or U22988 (N_22988,N_10188,N_12324);
nand U22989 (N_22989,N_15104,N_11197);
xnor U22990 (N_22990,N_11585,N_16504);
nand U22991 (N_22991,N_16594,N_11688);
xnor U22992 (N_22992,N_19530,N_13572);
nor U22993 (N_22993,N_11022,N_17133);
and U22994 (N_22994,N_15109,N_10184);
xor U22995 (N_22995,N_11893,N_10913);
xnor U22996 (N_22996,N_16299,N_11001);
or U22997 (N_22997,N_15665,N_12533);
nor U22998 (N_22998,N_13718,N_16117);
and U22999 (N_22999,N_12399,N_19963);
nand U23000 (N_23000,N_15250,N_16110);
and U23001 (N_23001,N_13194,N_14415);
nor U23002 (N_23002,N_18191,N_15392);
nand U23003 (N_23003,N_14030,N_11184);
or U23004 (N_23004,N_15675,N_11498);
xor U23005 (N_23005,N_12284,N_17525);
and U23006 (N_23006,N_14487,N_15055);
xor U23007 (N_23007,N_10041,N_16719);
nand U23008 (N_23008,N_11849,N_16166);
and U23009 (N_23009,N_12242,N_11200);
or U23010 (N_23010,N_16275,N_12367);
nand U23011 (N_23011,N_16841,N_12277);
nor U23012 (N_23012,N_17415,N_17798);
and U23013 (N_23013,N_11175,N_18826);
or U23014 (N_23014,N_18360,N_17929);
and U23015 (N_23015,N_11701,N_16500);
nand U23016 (N_23016,N_17047,N_15376);
or U23017 (N_23017,N_16950,N_10029);
xor U23018 (N_23018,N_13004,N_11064);
and U23019 (N_23019,N_15806,N_16722);
nor U23020 (N_23020,N_18618,N_12955);
and U23021 (N_23021,N_19845,N_19199);
nor U23022 (N_23022,N_14986,N_15804);
and U23023 (N_23023,N_10838,N_19168);
or U23024 (N_23024,N_17810,N_13630);
nor U23025 (N_23025,N_10650,N_15771);
nand U23026 (N_23026,N_12813,N_14049);
and U23027 (N_23027,N_19970,N_14500);
nand U23028 (N_23028,N_17336,N_11377);
nor U23029 (N_23029,N_19540,N_11208);
xnor U23030 (N_23030,N_18667,N_19230);
nor U23031 (N_23031,N_10226,N_19659);
or U23032 (N_23032,N_19336,N_11816);
or U23033 (N_23033,N_11548,N_11352);
nor U23034 (N_23034,N_19367,N_11237);
or U23035 (N_23035,N_13745,N_11940);
nand U23036 (N_23036,N_18433,N_15662);
xor U23037 (N_23037,N_11626,N_15391);
nand U23038 (N_23038,N_13446,N_13888);
xnor U23039 (N_23039,N_19487,N_15068);
or U23040 (N_23040,N_16005,N_10546);
xor U23041 (N_23041,N_19647,N_17103);
nand U23042 (N_23042,N_11559,N_14382);
and U23043 (N_23043,N_18127,N_14688);
or U23044 (N_23044,N_11906,N_14366);
nand U23045 (N_23045,N_14290,N_19669);
nand U23046 (N_23046,N_11103,N_14079);
or U23047 (N_23047,N_18273,N_11143);
or U23048 (N_23048,N_12273,N_18559);
xnor U23049 (N_23049,N_11467,N_17066);
and U23050 (N_23050,N_12354,N_14147);
nand U23051 (N_23051,N_18849,N_10142);
nand U23052 (N_23052,N_11102,N_17055);
and U23053 (N_23053,N_11081,N_16669);
and U23054 (N_23054,N_11788,N_14485);
or U23055 (N_23055,N_15718,N_10573);
nor U23056 (N_23056,N_10939,N_10670);
xnor U23057 (N_23057,N_13919,N_10479);
xor U23058 (N_23058,N_14047,N_12907);
nor U23059 (N_23059,N_15582,N_15116);
or U23060 (N_23060,N_15552,N_19009);
or U23061 (N_23061,N_11593,N_16407);
xnor U23062 (N_23062,N_18026,N_12259);
xnor U23063 (N_23063,N_14198,N_17183);
or U23064 (N_23064,N_18254,N_16104);
or U23065 (N_23065,N_15588,N_19931);
xor U23066 (N_23066,N_10674,N_17273);
and U23067 (N_23067,N_15514,N_16290);
xor U23068 (N_23068,N_18272,N_11644);
nor U23069 (N_23069,N_11949,N_13045);
nor U23070 (N_23070,N_19701,N_10034);
or U23071 (N_23071,N_17198,N_13317);
nor U23072 (N_23072,N_18881,N_13873);
and U23073 (N_23073,N_16858,N_15353);
or U23074 (N_23074,N_13023,N_16477);
nand U23075 (N_23075,N_12771,N_10752);
xor U23076 (N_23076,N_11490,N_19866);
and U23077 (N_23077,N_10258,N_12393);
xor U23078 (N_23078,N_15375,N_17971);
and U23079 (N_23079,N_15850,N_18641);
and U23080 (N_23080,N_12196,N_13908);
and U23081 (N_23081,N_17822,N_15415);
nand U23082 (N_23082,N_14063,N_18711);
or U23083 (N_23083,N_13742,N_16754);
xnor U23084 (N_23084,N_15106,N_10798);
nor U23085 (N_23085,N_14310,N_14112);
xor U23086 (N_23086,N_17167,N_11444);
nand U23087 (N_23087,N_12504,N_11093);
or U23088 (N_23088,N_10383,N_18087);
nor U23089 (N_23089,N_13764,N_18950);
or U23090 (N_23090,N_18032,N_14631);
nand U23091 (N_23091,N_11793,N_10675);
xnor U23092 (N_23092,N_14943,N_17040);
and U23093 (N_23093,N_10050,N_18313);
or U23094 (N_23094,N_10835,N_16143);
xnor U23095 (N_23095,N_11922,N_15944);
nor U23096 (N_23096,N_13793,N_10300);
nand U23097 (N_23097,N_13312,N_16124);
and U23098 (N_23098,N_12896,N_18068);
xnor U23099 (N_23099,N_15540,N_14603);
nand U23100 (N_23100,N_12902,N_16039);
and U23101 (N_23101,N_11908,N_12745);
xor U23102 (N_23102,N_12627,N_11545);
and U23103 (N_23103,N_10898,N_12442);
nand U23104 (N_23104,N_17344,N_15867);
and U23105 (N_23105,N_12276,N_14086);
or U23106 (N_23106,N_11920,N_15511);
nor U23107 (N_23107,N_11714,N_14845);
and U23108 (N_23108,N_19781,N_18059);
xor U23109 (N_23109,N_12167,N_10255);
nand U23110 (N_23110,N_10397,N_18511);
xor U23111 (N_23111,N_14202,N_13049);
nand U23112 (N_23112,N_14181,N_10724);
nand U23113 (N_23113,N_12840,N_12707);
nor U23114 (N_23114,N_19711,N_16699);
nand U23115 (N_23115,N_13211,N_14508);
nor U23116 (N_23116,N_16168,N_14843);
and U23117 (N_23117,N_11348,N_19341);
xor U23118 (N_23118,N_10922,N_10136);
nand U23119 (N_23119,N_14533,N_13298);
or U23120 (N_23120,N_13177,N_18999);
nand U23121 (N_23121,N_12744,N_18666);
or U23122 (N_23122,N_18297,N_19229);
and U23123 (N_23123,N_18706,N_12998);
or U23124 (N_23124,N_13523,N_17704);
nor U23125 (N_23125,N_14985,N_10246);
xor U23126 (N_23126,N_14573,N_15865);
nand U23127 (N_23127,N_17976,N_17442);
and U23128 (N_23128,N_13783,N_17762);
nand U23129 (N_23129,N_12296,N_11611);
nand U23130 (N_23130,N_17015,N_13767);
nor U23131 (N_23131,N_18258,N_14408);
xnor U23132 (N_23132,N_12071,N_14792);
or U23133 (N_23133,N_17325,N_12181);
xor U23134 (N_23134,N_14550,N_16130);
xor U23135 (N_23135,N_10475,N_12228);
or U23136 (N_23136,N_18479,N_12460);
and U23137 (N_23137,N_11659,N_15341);
nor U23138 (N_23138,N_11296,N_15951);
nor U23139 (N_23139,N_14987,N_16847);
xor U23140 (N_23140,N_10900,N_15321);
xor U23141 (N_23141,N_11967,N_17797);
nand U23142 (N_23142,N_17946,N_14011);
nand U23143 (N_23143,N_10569,N_12327);
nor U23144 (N_23144,N_15240,N_17024);
nor U23145 (N_23145,N_19134,N_11656);
and U23146 (N_23146,N_12250,N_13949);
nand U23147 (N_23147,N_17121,N_12156);
nor U23148 (N_23148,N_10395,N_15928);
nand U23149 (N_23149,N_18278,N_15477);
nor U23150 (N_23150,N_16118,N_17202);
nand U23151 (N_23151,N_17622,N_11772);
xor U23152 (N_23152,N_19937,N_14430);
and U23153 (N_23153,N_19031,N_13801);
nand U23154 (N_23154,N_13089,N_10727);
xor U23155 (N_23155,N_18610,N_17117);
xor U23156 (N_23156,N_15912,N_13117);
xnor U23157 (N_23157,N_15067,N_13932);
nand U23158 (N_23158,N_13542,N_12307);
or U23159 (N_23159,N_19094,N_18314);
nand U23160 (N_23160,N_14710,N_14361);
nor U23161 (N_23161,N_16178,N_14294);
nand U23162 (N_23162,N_14503,N_17021);
nand U23163 (N_23163,N_14029,N_18107);
xnor U23164 (N_23164,N_11823,N_11641);
nand U23165 (N_23165,N_14189,N_12688);
and U23166 (N_23166,N_15998,N_16683);
xor U23167 (N_23167,N_14016,N_11193);
nand U23168 (N_23168,N_13909,N_18939);
xor U23169 (N_23169,N_16323,N_16637);
nand U23170 (N_23170,N_17090,N_13553);
nand U23171 (N_23171,N_10437,N_13874);
xor U23172 (N_23172,N_15930,N_11674);
nor U23173 (N_23173,N_10036,N_19290);
xor U23174 (N_23174,N_15832,N_18865);
and U23175 (N_23175,N_16151,N_13790);
and U23176 (N_23176,N_16298,N_19018);
or U23177 (N_23177,N_18720,N_17477);
nor U23178 (N_23178,N_11665,N_17438);
nor U23179 (N_23179,N_18708,N_18578);
nor U23180 (N_23180,N_17043,N_19369);
nor U23181 (N_23181,N_16610,N_11899);
or U23182 (N_23182,N_13320,N_13565);
nor U23183 (N_23183,N_12062,N_15635);
nor U23184 (N_23184,N_11671,N_13809);
or U23185 (N_23185,N_12805,N_13683);
nor U23186 (N_23186,N_10591,N_18848);
and U23187 (N_23187,N_19445,N_19773);
xnor U23188 (N_23188,N_17127,N_13761);
nor U23189 (N_23189,N_13970,N_12386);
or U23190 (N_23190,N_18793,N_18237);
and U23191 (N_23191,N_11292,N_19785);
nor U23192 (N_23192,N_13668,N_15292);
and U23193 (N_23193,N_10786,N_10038);
nand U23194 (N_23194,N_17292,N_14156);
and U23195 (N_23195,N_16623,N_14652);
nor U23196 (N_23196,N_13300,N_10266);
or U23197 (N_23197,N_13539,N_18722);
nand U23198 (N_23198,N_17106,N_14138);
and U23199 (N_23199,N_11190,N_11685);
and U23200 (N_23200,N_17351,N_19766);
and U23201 (N_23201,N_14650,N_19683);
nor U23202 (N_23202,N_12683,N_18161);
nor U23203 (N_23203,N_14182,N_10236);
and U23204 (N_23204,N_16900,N_17267);
and U23205 (N_23205,N_11448,N_17865);
nor U23206 (N_23206,N_16395,N_12334);
xnor U23207 (N_23207,N_13952,N_14315);
xnor U23208 (N_23208,N_18675,N_16474);
or U23209 (N_23209,N_10627,N_10190);
nand U23210 (N_23210,N_10060,N_18698);
or U23211 (N_23211,N_18299,N_15191);
and U23212 (N_23212,N_15451,N_10745);
xnor U23213 (N_23213,N_11042,N_14359);
and U23214 (N_23214,N_13015,N_11736);
or U23215 (N_23215,N_19169,N_14864);
nand U23216 (N_23216,N_12838,N_18432);
and U23217 (N_23217,N_10680,N_14649);
xnor U23218 (N_23218,N_13226,N_15295);
xor U23219 (N_23219,N_12736,N_14306);
nor U23220 (N_23220,N_14892,N_10474);
or U23221 (N_23221,N_15049,N_17249);
nor U23222 (N_23222,N_17084,N_19074);
or U23223 (N_23223,N_10025,N_16533);
nor U23224 (N_23224,N_13198,N_19111);
or U23225 (N_23225,N_13872,N_13759);
and U23226 (N_23226,N_19724,N_12299);
and U23227 (N_23227,N_11539,N_14849);
or U23228 (N_23228,N_17690,N_15303);
and U23229 (N_23229,N_10080,N_14728);
and U23230 (N_23230,N_14778,N_15336);
nor U23231 (N_23231,N_15356,N_18399);
or U23232 (N_23232,N_15278,N_18662);
nor U23233 (N_23233,N_13007,N_15305);
nand U23234 (N_23234,N_13694,N_19534);
xnor U23235 (N_23235,N_15989,N_14133);
nor U23236 (N_23236,N_14024,N_19254);
and U23237 (N_23237,N_14788,N_12613);
nor U23238 (N_23238,N_17424,N_15426);
and U23239 (N_23239,N_18682,N_12931);
nand U23240 (N_23240,N_10800,N_13758);
xor U23241 (N_23241,N_11687,N_10592);
xnor U23242 (N_23242,N_17863,N_14702);
nand U23243 (N_23243,N_10609,N_16717);
nor U23244 (N_23244,N_18636,N_16987);
or U23245 (N_23245,N_12590,N_15761);
and U23246 (N_23246,N_17760,N_11075);
nor U23247 (N_23247,N_12126,N_10628);
xor U23248 (N_23248,N_19629,N_11883);
nor U23249 (N_23249,N_18295,N_15567);
nand U23250 (N_23250,N_16314,N_19625);
nor U23251 (N_23251,N_14863,N_14621);
or U23252 (N_23252,N_12287,N_13391);
xnor U23253 (N_23253,N_13599,N_11700);
nand U23254 (N_23254,N_17384,N_19294);
nor U23255 (N_23255,N_13026,N_15862);
nor U23256 (N_23256,N_19043,N_10915);
nand U23257 (N_23257,N_10826,N_11016);
or U23258 (N_23258,N_16199,N_18014);
and U23259 (N_23259,N_11381,N_11584);
and U23260 (N_23260,N_10052,N_11726);
and U23261 (N_23261,N_13950,N_12083);
nor U23262 (N_23262,N_11010,N_10773);
xor U23263 (N_23263,N_17920,N_16526);
xor U23264 (N_23264,N_12875,N_10829);
xnor U23265 (N_23265,N_19084,N_14448);
nor U23266 (N_23266,N_17924,N_12601);
and U23267 (N_23267,N_10596,N_18668);
nand U23268 (N_23268,N_19488,N_15863);
xnor U23269 (N_23269,N_16241,N_16608);
nor U23270 (N_23270,N_10409,N_14975);
or U23271 (N_23271,N_13858,N_13830);
nand U23272 (N_23272,N_16505,N_10312);
xor U23273 (N_23273,N_11825,N_10683);
nand U23274 (N_23274,N_18130,N_13167);
or U23275 (N_23275,N_10189,N_15890);
nand U23276 (N_23276,N_18205,N_11842);
nand U23277 (N_23277,N_18088,N_19977);
and U23278 (N_23278,N_16416,N_18560);
xor U23279 (N_23279,N_16068,N_10901);
and U23280 (N_23280,N_13498,N_17195);
and U23281 (N_23281,N_16239,N_10486);
nor U23282 (N_23282,N_17586,N_12898);
and U23283 (N_23283,N_13418,N_11223);
and U23284 (N_23284,N_16264,N_15154);
nor U23285 (N_23285,N_13024,N_12864);
or U23286 (N_23286,N_10590,N_16878);
nand U23287 (N_23287,N_19421,N_18967);
nand U23288 (N_23288,N_18089,N_14231);
xnor U23289 (N_23289,N_11345,N_14084);
and U23290 (N_23290,N_10179,N_13665);
xnor U23291 (N_23291,N_12692,N_17020);
nor U23292 (N_23292,N_13521,N_15725);
nor U23293 (N_23293,N_19012,N_14035);
and U23294 (N_23294,N_12161,N_10768);
xnor U23295 (N_23295,N_13463,N_16056);
and U23296 (N_23296,N_15531,N_18171);
and U23297 (N_23297,N_18339,N_16384);
or U23298 (N_23298,N_11128,N_10992);
xor U23299 (N_23299,N_10524,N_11378);
nand U23300 (N_23300,N_14875,N_11864);
or U23301 (N_23301,N_12575,N_17307);
xnor U23302 (N_23302,N_16357,N_18772);
or U23303 (N_23303,N_19087,N_18520);
xor U23304 (N_23304,N_19097,N_15185);
and U23305 (N_23305,N_18447,N_11392);
and U23306 (N_23306,N_10834,N_16180);
and U23307 (N_23307,N_17489,N_13077);
or U23308 (N_23308,N_13341,N_17008);
and U23309 (N_23309,N_11218,N_13143);
and U23310 (N_23310,N_11285,N_12765);
nand U23311 (N_23311,N_14312,N_13223);
nand U23312 (N_23312,N_13365,N_16187);
and U23313 (N_23313,N_12760,N_12548);
and U23314 (N_23314,N_16252,N_16598);
and U23315 (N_23315,N_17637,N_18681);
and U23316 (N_23316,N_16242,N_19624);
and U23317 (N_23317,N_13366,N_11350);
xnor U23318 (N_23318,N_19968,N_16248);
nand U23319 (N_23319,N_14420,N_18568);
or U23320 (N_23320,N_18410,N_13706);
xnor U23321 (N_23321,N_18311,N_17002);
and U23322 (N_23322,N_12352,N_13666);
nand U23323 (N_23323,N_15022,N_12400);
xnor U23324 (N_23324,N_15099,N_19507);
and U23325 (N_23325,N_19385,N_18823);
nor U23326 (N_23326,N_17197,N_16284);
or U23327 (N_23327,N_16358,N_11477);
xor U23328 (N_23328,N_12404,N_10991);
or U23329 (N_23329,N_15367,N_12517);
nor U23330 (N_23330,N_13237,N_19252);
xor U23331 (N_23331,N_19475,N_17950);
or U23332 (N_23332,N_19030,N_12512);
nand U23333 (N_23333,N_12093,N_19709);
and U23334 (N_23334,N_16585,N_17707);
xor U23335 (N_23335,N_11406,N_18851);
and U23336 (N_23336,N_13794,N_18966);
or U23337 (N_23337,N_19805,N_15907);
and U23338 (N_23338,N_14463,N_16799);
nand U23339 (N_23339,N_18054,N_12064);
and U23340 (N_23340,N_17801,N_18678);
nand U23341 (N_23341,N_12580,N_19784);
nand U23342 (N_23342,N_13805,N_14819);
and U23343 (N_23343,N_18257,N_13476);
nand U23344 (N_23344,N_16142,N_18624);
nand U23345 (N_23345,N_15061,N_10708);
xor U23346 (N_23346,N_10256,N_16368);
nor U23347 (N_23347,N_13788,N_11506);
or U23348 (N_23348,N_13430,N_18639);
and U23349 (N_23349,N_19554,N_14333);
nand U23350 (N_23350,N_19543,N_16726);
nand U23351 (N_23351,N_13267,N_16156);
and U23352 (N_23352,N_13681,N_18039);
or U23353 (N_23353,N_15721,N_15667);
or U23354 (N_23354,N_13892,N_10067);
or U23355 (N_23355,N_15351,N_18241);
and U23356 (N_23356,N_12702,N_19857);
nand U23357 (N_23357,N_12109,N_16175);
nor U23358 (N_23358,N_12198,N_18705);
nand U23359 (N_23359,N_17555,N_13332);
or U23360 (N_23360,N_10647,N_10906);
nand U23361 (N_23361,N_17784,N_18008);
xnor U23362 (N_23362,N_15674,N_16024);
and U23363 (N_23363,N_10064,N_12565);
nor U23364 (N_23364,N_16978,N_14038);
nand U23365 (N_23365,N_16244,N_14357);
or U23366 (N_23366,N_16133,N_11459);
nor U23367 (N_23367,N_12446,N_19426);
xor U23368 (N_23368,N_19242,N_12292);
xor U23369 (N_23369,N_15249,N_11838);
and U23370 (N_23370,N_13732,N_16936);
nor U23371 (N_23371,N_12790,N_11297);
nand U23372 (N_23372,N_10429,N_10801);
or U23373 (N_23373,N_18518,N_17051);
and U23374 (N_23374,N_11289,N_19756);
and U23375 (N_23375,N_19360,N_11429);
xor U23376 (N_23376,N_10073,N_12489);
and U23377 (N_23377,N_17210,N_15464);
nor U23378 (N_23378,N_11610,N_13311);
nor U23379 (N_23379,N_18179,N_16676);
nor U23380 (N_23380,N_12614,N_16303);
nand U23381 (N_23381,N_10487,N_10555);
nand U23382 (N_23382,N_19814,N_10730);
xor U23383 (N_23383,N_10485,N_13316);
and U23384 (N_23384,N_19895,N_10963);
and U23385 (N_23385,N_10163,N_10104);
xnor U23386 (N_23386,N_13727,N_18351);
and U23387 (N_23387,N_11286,N_11887);
nand U23388 (N_23388,N_19941,N_12157);
nand U23389 (N_23389,N_18235,N_18128);
nand U23390 (N_23390,N_10011,N_19081);
and U23391 (N_23391,N_18874,N_13134);
xnor U23392 (N_23392,N_17559,N_19969);
nand U23393 (N_23393,N_19011,N_19909);
xor U23394 (N_23394,N_12162,N_19433);
xor U23395 (N_23395,N_19596,N_13483);
nor U23396 (N_23396,N_14746,N_19949);
nor U23397 (N_23397,N_13810,N_19212);
nand U23398 (N_23398,N_17282,N_16513);
and U23399 (N_23399,N_14854,N_16253);
xor U23400 (N_23400,N_13688,N_12054);
or U23401 (N_23401,N_18279,N_11483);
xor U23402 (N_23402,N_15237,N_15663);
nor U23403 (N_23403,N_12546,N_18765);
nand U23404 (N_23404,N_11424,N_18890);
nor U23405 (N_23405,N_12269,N_13470);
and U23406 (N_23406,N_17395,N_19533);
nor U23407 (N_23407,N_14135,N_10971);
nor U23408 (N_23408,N_14818,N_19566);
and U23409 (N_23409,N_16806,N_10375);
and U23410 (N_23410,N_16008,N_13627);
or U23411 (N_23411,N_15605,N_12986);
nand U23412 (N_23412,N_19008,N_14391);
nor U23413 (N_23413,N_11329,N_15919);
xnor U23414 (N_23414,N_13836,N_10425);
or U23415 (N_23415,N_12220,N_10943);
nand U23416 (N_23416,N_12726,N_17130);
or U23417 (N_23417,N_19040,N_19112);
and U23418 (N_23418,N_15568,N_18971);
nand U23419 (N_23419,N_18402,N_10986);
nor U23420 (N_23420,N_12556,N_16456);
nand U23421 (N_23421,N_16483,N_12382);
nand U23422 (N_23422,N_15687,N_14996);
or U23423 (N_23423,N_10543,N_16872);
nand U23424 (N_23424,N_14654,N_10649);
nand U23425 (N_23425,N_17290,N_11969);
xor U23426 (N_23426,N_12881,N_17337);
and U23427 (N_23427,N_13848,N_14510);
nor U23428 (N_23428,N_13646,N_14264);
xor U23429 (N_23429,N_15216,N_13329);
xor U23430 (N_23430,N_15438,N_10276);
nand U23431 (N_23431,N_13819,N_19597);
nor U23432 (N_23432,N_13850,N_14718);
nor U23433 (N_23433,N_15983,N_14471);
xnor U23434 (N_23434,N_10747,N_18839);
nand U23435 (N_23435,N_14743,N_15146);
nor U23436 (N_23436,N_11479,N_15886);
and U23437 (N_23437,N_19760,N_18210);
xnor U23438 (N_23438,N_17123,N_16631);
and U23439 (N_23439,N_18105,N_11606);
and U23440 (N_23440,N_16300,N_18456);
xnor U23441 (N_23441,N_11346,N_12123);
nor U23442 (N_23442,N_13964,N_17226);
nor U23443 (N_23443,N_11206,N_10293);
and U23444 (N_23444,N_17313,N_17527);
and U23445 (N_23445,N_14716,N_16830);
and U23446 (N_23446,N_14597,N_14993);
nor U23447 (N_23447,N_11682,N_14618);
or U23448 (N_23448,N_16063,N_16135);
xor U23449 (N_23449,N_19823,N_19131);
xor U23450 (N_23450,N_12039,N_10993);
xnor U23451 (N_23451,N_13207,N_13865);
xor U23452 (N_23452,N_10384,N_15836);
nor U23453 (N_23453,N_12069,N_18958);
xnor U23454 (N_23454,N_18290,N_15027);
or U23455 (N_23455,N_12617,N_18873);
and U23456 (N_23456,N_13814,N_11799);
nand U23457 (N_23457,N_13123,N_14537);
or U23458 (N_23458,N_18972,N_11083);
nor U23459 (N_23459,N_12376,N_10235);
xnor U23460 (N_23460,N_17773,N_12200);
xor U23461 (N_23461,N_13142,N_14167);
xor U23462 (N_23462,N_14884,N_18756);
and U23463 (N_23463,N_15639,N_16226);
or U23464 (N_23464,N_10433,N_13671);
nor U23465 (N_23465,N_17367,N_18504);
nor U23466 (N_23466,N_11077,N_16965);
and U23467 (N_23467,N_18777,N_17573);
nor U23468 (N_23468,N_12538,N_10275);
or U23469 (N_23469,N_14266,N_17553);
and U23470 (N_23470,N_14449,N_18338);
xor U23471 (N_23471,N_18745,N_18642);
xor U23472 (N_23472,N_19027,N_16403);
nand U23473 (N_23473,N_16309,N_11634);
nand U23474 (N_23474,N_16421,N_13726);
and U23475 (N_23475,N_18855,N_17645);
nand U23476 (N_23476,N_12541,N_13803);
nand U23477 (N_23477,N_10427,N_18897);
xnor U23478 (N_23478,N_15015,N_11961);
nor U23479 (N_23479,N_12964,N_10792);
nor U23480 (N_23480,N_14700,N_14805);
xor U23481 (N_23481,N_10171,N_17968);
nand U23482 (N_23482,N_13965,N_10304);
and U23483 (N_23483,N_10661,N_18289);
and U23484 (N_23484,N_13091,N_18296);
or U23485 (N_23485,N_19972,N_16654);
nor U23486 (N_23486,N_18900,N_14276);
nor U23487 (N_23487,N_16906,N_11959);
nand U23488 (N_23488,N_14994,N_17370);
xor U23489 (N_23489,N_16228,N_13641);
xnor U23490 (N_23490,N_15777,N_16057);
and U23491 (N_23491,N_19794,N_19236);
xor U23492 (N_23492,N_13471,N_14466);
xor U23493 (N_23493,N_16267,N_13043);
nand U23494 (N_23494,N_11342,N_11707);
or U23495 (N_23495,N_12673,N_12110);
or U23496 (N_23496,N_19829,N_16548);
and U23497 (N_23497,N_18412,N_13262);
and U23498 (N_23498,N_14951,N_15631);
nor U23499 (N_23499,N_17458,N_18933);
and U23500 (N_23500,N_12658,N_14416);
nand U23501 (N_23501,N_18001,N_16942);
nor U23502 (N_23502,N_15497,N_15924);
xor U23503 (N_23503,N_14831,N_16206);
nand U23504 (N_23504,N_17843,N_15533);
nor U23505 (N_23505,N_11231,N_11820);
nand U23506 (N_23506,N_10687,N_10497);
nand U23507 (N_23507,N_18561,N_15518);
and U23508 (N_23508,N_13760,N_10969);
nand U23509 (N_23509,N_16541,N_18604);
and U23510 (N_23510,N_15409,N_12848);
nor U23511 (N_23511,N_12225,N_16370);
xnor U23512 (N_23512,N_17046,N_15315);
and U23513 (N_23513,N_12182,N_17166);
or U23514 (N_23514,N_15318,N_14428);
nor U23515 (N_23515,N_13748,N_19165);
or U23516 (N_23516,N_19973,N_16702);
nor U23517 (N_23517,N_13797,N_17524);
xnor U23518 (N_23518,N_17552,N_12967);
and U23519 (N_23519,N_10282,N_17493);
and U23520 (N_23520,N_15020,N_18987);
or U23521 (N_23521,N_15601,N_15827);
xnor U23522 (N_23522,N_16333,N_11834);
or U23523 (N_23523,N_10209,N_13041);
xnor U23524 (N_23524,N_10366,N_16884);
and U23525 (N_23525,N_12850,N_17189);
nand U23526 (N_23526,N_13428,N_10017);
nor U23527 (N_23527,N_15000,N_10018);
nand U23528 (N_23528,N_15993,N_14560);
nand U23529 (N_23529,N_14820,N_13903);
nand U23530 (N_23530,N_17410,N_14541);
nor U23531 (N_23531,N_10845,N_10912);
xnor U23532 (N_23532,N_19681,N_18723);
or U23533 (N_23533,N_19434,N_10035);
xnor U23534 (N_23534,N_12300,N_17809);
and U23535 (N_23535,N_12734,N_10810);
or U23536 (N_23536,N_17738,N_18460);
and U23537 (N_23537,N_12149,N_19736);
nand U23538 (N_23538,N_10830,N_18886);
and U23539 (N_23539,N_13140,N_14903);
xor U23540 (N_23540,N_17538,N_19315);
xnor U23541 (N_23541,N_15881,N_12959);
nand U23542 (N_23542,N_17715,N_11785);
or U23543 (N_23543,N_14073,N_19265);
or U23544 (N_23544,N_12355,N_16216);
nand U23545 (N_23545,N_17932,N_16082);
nand U23546 (N_23546,N_16749,N_11549);
nor U23547 (N_23547,N_11354,N_11114);
nor U23548 (N_23548,N_13894,N_10756);
xor U23549 (N_23549,N_16968,N_16326);
nand U23550 (N_23550,N_11904,N_15630);
xor U23551 (N_23551,N_12202,N_10935);
nor U23552 (N_23552,N_17154,N_17748);
and U23553 (N_23553,N_15135,N_17093);
and U23554 (N_23554,N_19987,N_16662);
xnor U23555 (N_23555,N_15231,N_18160);
xnor U23556 (N_23556,N_19015,N_11308);
nand U23557 (N_23557,N_10464,N_17075);
nor U23558 (N_23558,N_11125,N_19373);
or U23559 (N_23559,N_16519,N_10528);
xnor U23560 (N_23560,N_17323,N_15377);
or U23561 (N_23561,N_10956,N_13571);
nand U23562 (N_23562,N_18002,N_17211);
nor U23563 (N_23563,N_13263,N_16077);
or U23564 (N_23564,N_10597,N_10656);
or U23565 (N_23565,N_17868,N_14691);
nand U23566 (N_23566,N_14736,N_16832);
xor U23567 (N_23567,N_16866,N_12190);
and U23568 (N_23568,N_12947,N_18941);
nand U23569 (N_23569,N_10027,N_18034);
or U23570 (N_23570,N_12678,N_10022);
nand U23571 (N_23571,N_16616,N_17030);
xnor U23572 (N_23572,N_17849,N_10595);
or U23573 (N_23573,N_17813,N_10360);
or U23574 (N_23574,N_14984,N_19284);
nor U23575 (N_23575,N_18291,N_16473);
nand U23576 (N_23576,N_17503,N_18482);
xor U23577 (N_23577,N_10478,N_13458);
and U23578 (N_23578,N_12488,N_18857);
nor U23579 (N_23579,N_12211,N_16231);
or U23580 (N_23580,N_19410,N_15543);
and U23581 (N_23581,N_17808,N_11773);
xor U23582 (N_23582,N_19643,N_13416);
nand U23583 (N_23583,N_16066,N_14046);
nand U23584 (N_23584,N_15498,N_10937);
or U23585 (N_23585,N_17261,N_15017);
nand U23586 (N_23586,N_13730,N_16060);
xor U23587 (N_23587,N_14388,N_11446);
nor U23588 (N_23588,N_19281,N_10016);
and U23589 (N_23589,N_12465,N_15086);
or U23590 (N_23590,N_11854,N_16382);
and U23591 (N_23591,N_14799,N_10959);
nor U23592 (N_23592,N_13626,N_10988);
nor U23593 (N_23593,N_18870,N_19608);
xnor U23594 (N_23594,N_19264,N_14565);
nand U23595 (N_23595,N_17322,N_15350);
or U23596 (N_23596,N_18430,N_15889);
and U23597 (N_23597,N_16592,N_17930);
nor U23598 (N_23598,N_17497,N_18794);
and U23599 (N_23599,N_16740,N_18654);
nor U23600 (N_23600,N_15246,N_10874);
xor U23601 (N_23601,N_10827,N_12699);
and U23602 (N_23602,N_13541,N_13691);
and U23603 (N_23603,N_19159,N_19484);
or U23604 (N_23604,N_12270,N_18969);
and U23605 (N_23605,N_18375,N_15172);
nor U23606 (N_23606,N_19902,N_18709);
nor U23607 (N_23607,N_16812,N_10292);
and U23608 (N_23608,N_18542,N_12088);
or U23609 (N_23609,N_13507,N_15018);
nor U23610 (N_23610,N_11380,N_15697);
or U23611 (N_23611,N_15809,N_15169);
nand U23612 (N_23612,N_10494,N_15608);
nor U23613 (N_23613,N_12318,N_14624);
xnor U23614 (N_23614,N_14938,N_18335);
and U23615 (N_23615,N_18715,N_18687);
or U23616 (N_23616,N_18172,N_13434);
nand U23617 (N_23617,N_12845,N_18212);
and U23618 (N_23618,N_14360,N_16745);
or U23619 (N_23619,N_10941,N_15934);
xnor U23620 (N_23620,N_10850,N_13528);
nand U23621 (N_23621,N_19448,N_18852);
xnor U23622 (N_23622,N_12257,N_19152);
and U23623 (N_23623,N_14605,N_10129);
nor U23624 (N_23624,N_16001,N_17140);
nor U23625 (N_23625,N_14709,N_15389);
nor U23626 (N_23626,N_15207,N_14920);
and U23627 (N_23627,N_16337,N_18428);
or U23628 (N_23628,N_10031,N_11554);
and U23629 (N_23629,N_19952,N_19635);
nor U23630 (N_23630,N_15075,N_17218);
or U23631 (N_23631,N_11040,N_10796);
or U23632 (N_23632,N_15536,N_15557);
xor U23633 (N_23633,N_14988,N_17791);
xor U23634 (N_23634,N_19197,N_12670);
nand U23635 (N_23635,N_17570,N_11630);
nor U23636 (N_23636,N_11915,N_17750);
nand U23637 (N_23637,N_19427,N_16445);
nor U23638 (N_23638,N_18845,N_12057);
or U23639 (N_23639,N_10207,N_11783);
nor U23640 (N_23640,N_13558,N_18603);
xor U23641 (N_23641,N_19827,N_12431);
xor U23642 (N_23642,N_14639,N_16263);
nand U23643 (N_23643,N_17656,N_19552);
xnor U23644 (N_23644,N_12053,N_18184);
or U23645 (N_23645,N_19181,N_13707);
xor U23646 (N_23646,N_16127,N_19162);
nand U23647 (N_23647,N_13216,N_16881);
xnor U23648 (N_23648,N_17236,N_18044);
nand U23649 (N_23649,N_15164,N_15824);
xor U23650 (N_23650,N_14781,N_15314);
xnor U23651 (N_23651,N_17988,N_19517);
nand U23652 (N_23652,N_14495,N_16076);
nor U23653 (N_23653,N_14954,N_12540);
nor U23654 (N_23654,N_11935,N_14281);
xnor U23655 (N_23655,N_17328,N_13577);
nand U23656 (N_23656,N_17058,N_18509);
nand U23657 (N_23657,N_18379,N_18174);
xor U23658 (N_23658,N_19370,N_15444);
or U23659 (N_23659,N_12892,N_12180);
nand U23660 (N_23660,N_15851,N_15094);
xnor U23661 (N_23661,N_19050,N_17181);
or U23662 (N_23662,N_13990,N_14121);
nor U23663 (N_23663,N_18909,N_13982);
or U23664 (N_23664,N_19389,N_19402);
xnor U23665 (N_23665,N_13684,N_12626);
xnor U23666 (N_23666,N_17890,N_13708);
nor U23667 (N_23667,N_11912,N_17098);
or U23668 (N_23668,N_13701,N_11988);
and U23669 (N_23669,N_15703,N_17906);
nand U23670 (N_23670,N_13173,N_18204);
and U23671 (N_23671,N_14837,N_11673);
and U23672 (N_23672,N_19239,N_16051);
and U23673 (N_23673,N_10147,N_14325);
or U23674 (N_23674,N_17501,N_15719);
nor U23675 (N_23675,N_18902,N_19925);
and U23676 (N_23676,N_12729,N_14318);
nand U23677 (N_23677,N_15978,N_14538);
or U23678 (N_23678,N_19663,N_14218);
nand U23679 (N_23679,N_14042,N_17386);
nor U23680 (N_23680,N_19148,N_13922);
xnor U23681 (N_23681,N_14474,N_12491);
nor U23682 (N_23682,N_14330,N_17485);
and U23683 (N_23683,N_16981,N_17285);
or U23684 (N_23684,N_12369,N_11131);
nor U23685 (N_23685,N_10812,N_12858);
and U23686 (N_23686,N_11461,N_16405);
or U23687 (N_23687,N_16875,N_19553);
and U23688 (N_23688,N_14056,N_10620);
nor U23689 (N_23689,N_18773,N_17649);
nor U23690 (N_23690,N_10183,N_12029);
xnor U23691 (N_23691,N_10789,N_15322);
xor U23692 (N_23692,N_11013,N_17413);
nand U23693 (N_23693,N_17611,N_19892);
and U23694 (N_23694,N_15791,N_14571);
xor U23695 (N_23695,N_11326,N_11428);
nor U23696 (N_23696,N_14912,N_10822);
nand U23697 (N_23697,N_14591,N_19658);
or U23698 (N_23698,N_10043,N_17941);
xnor U23699 (N_23699,N_17701,N_13989);
or U23700 (N_23700,N_16089,N_13544);
nand U23701 (N_23701,N_16167,N_16718);
and U23702 (N_23702,N_12700,N_14506);
or U23703 (N_23703,N_10772,N_13857);
or U23704 (N_23704,N_16294,N_15859);
or U23705 (N_23705,N_18634,N_19133);
and U23706 (N_23706,N_12560,N_15034);
nor U23707 (N_23707,N_12666,N_17085);
nand U23708 (N_23708,N_11800,N_10782);
nand U23709 (N_23709,N_17000,N_16287);
or U23710 (N_23710,N_13517,N_17508);
or U23711 (N_23711,N_11791,N_16591);
nor U23712 (N_23712,N_13879,N_17246);
or U23713 (N_23713,N_18095,N_15326);
xnor U23714 (N_23714,N_17970,N_15577);
or U23715 (N_23715,N_10523,N_19680);
or U23716 (N_23716,N_17476,N_10552);
nor U23717 (N_23717,N_10917,N_14512);
nor U23718 (N_23718,N_14750,N_10342);
nand U23719 (N_23719,N_14055,N_12721);
and U23720 (N_23720,N_11818,N_16924);
and U23721 (N_23721,N_12828,N_14129);
or U23722 (N_23722,N_18294,N_13440);
xor U23723 (N_23723,N_13611,N_19644);
xnor U23724 (N_23724,N_16201,N_13050);
nand U23725 (N_23725,N_14527,N_15425);
xor U23726 (N_23726,N_14842,N_17550);
or U23727 (N_23727,N_16245,N_15484);
nand U23728 (N_23728,N_19771,N_11977);
or U23729 (N_23729,N_13963,N_18877);
nor U23730 (N_23730,N_11402,N_17882);
and U23731 (N_23731,N_19368,N_15634);
or U23732 (N_23732,N_10603,N_12265);
xor U23733 (N_23733,N_12471,N_10693);
nor U23734 (N_23734,N_16839,N_11717);
or U23735 (N_23735,N_19511,N_18788);
nand U23736 (N_23736,N_11385,N_19688);
nand U23737 (N_23737,N_13620,N_14812);
or U23738 (N_23738,N_11323,N_10238);
nor U23739 (N_23739,N_18959,N_11607);
nand U23740 (N_23740,N_19472,N_14403);
nand U23741 (N_23741,N_12897,N_11158);
xor U23742 (N_23742,N_15672,N_16004);
nor U23743 (N_23743,N_15839,N_17441);
and U23744 (N_23744,N_15114,N_16539);
nand U23745 (N_23745,N_16176,N_15942);
xor U23746 (N_23746,N_18441,N_13180);
or U23747 (N_23747,N_10953,N_11344);
nor U23748 (N_23748,N_16270,N_17512);
and U23749 (N_23749,N_19873,N_15471);
or U23750 (N_23750,N_16204,N_11119);
xor U23751 (N_23751,N_12660,N_15288);
or U23752 (N_23752,N_11276,N_14977);
xor U23753 (N_23753,N_14822,N_19253);
nand U23754 (N_23754,N_15186,N_10927);
nand U23755 (N_23755,N_15103,N_18112);
and U23756 (N_23756,N_12016,N_15042);
and U23757 (N_23757,N_12403,N_18998);
nand U23758 (N_23758,N_18005,N_18779);
nor U23759 (N_23759,N_13569,N_18101);
and U23760 (N_23760,N_18543,N_15229);
nor U23761 (N_23761,N_16624,N_13996);
or U23762 (N_23762,N_12006,N_13930);
xor U23763 (N_23763,N_12456,N_16010);
xor U23764 (N_23764,N_15840,N_19329);
or U23765 (N_23765,N_13497,N_19072);
nand U23766 (N_23766,N_14766,N_13268);
or U23767 (N_23767,N_15508,N_19725);
nand U23768 (N_23768,N_14893,N_17772);
nor U23769 (N_23769,N_18239,N_16768);
or U23770 (N_23770,N_16640,N_13165);
or U23771 (N_23771,N_16763,N_16577);
and U23772 (N_23772,N_15479,N_19359);
nor U23773 (N_23773,N_16059,N_10525);
nor U23774 (N_23774,N_17629,N_10985);
nor U23775 (N_23775,N_12806,N_19411);
xnor U23776 (N_23776,N_13596,N_15858);
or U23777 (N_23777,N_18163,N_11453);
nor U23778 (N_23778,N_19749,N_10245);
nor U23779 (N_23779,N_14685,N_14066);
or U23780 (N_23780,N_13466,N_11387);
nand U23781 (N_23781,N_19888,N_15224);
and U23782 (N_23782,N_12345,N_16709);
nand U23783 (N_23783,N_14328,N_16092);
xnor U23784 (N_23784,N_13700,N_17855);
nand U23785 (N_23785,N_11165,N_13334);
xor U23786 (N_23786,N_13740,N_14775);
xnor U23787 (N_23787,N_18820,N_10152);
nor U23788 (N_23788,N_17091,N_14595);
and U23789 (N_23789,N_10106,N_11519);
xnor U23790 (N_23790,N_12436,N_15971);
and U23791 (N_23791,N_18626,N_12128);
or U23792 (N_23792,N_16394,N_14176);
or U23793 (N_23793,N_14829,N_16636);
xnor U23794 (N_23794,N_16871,N_18876);
nand U23795 (N_23795,N_15029,N_16084);
or U23796 (N_23796,N_12033,N_12770);
and U23797 (N_23797,N_11913,N_11155);
nor U23798 (N_23798,N_15664,N_17082);
xor U23799 (N_23799,N_14437,N_16967);
xor U23800 (N_23800,N_18167,N_14301);
or U23801 (N_23801,N_15690,N_10482);
nand U23802 (N_23802,N_11112,N_13392);
and U23803 (N_23803,N_11712,N_15921);
and U23804 (N_23804,N_19189,N_19384);
xor U23805 (N_23805,N_16238,N_14427);
xor U23806 (N_23806,N_15752,N_19042);
nor U23807 (N_23807,N_12509,N_12972);
nor U23808 (N_23808,N_13563,N_10008);
or U23809 (N_23809,N_19906,N_12561);
nor U23810 (N_23810,N_15023,N_18367);
nand U23811 (N_23811,N_18397,N_12137);
nor U23812 (N_23812,N_18007,N_19509);
or U23813 (N_23813,N_17354,N_16182);
nor U23814 (N_23814,N_15030,N_14215);
and U23815 (N_23815,N_11748,N_18546);
or U23816 (N_23816,N_11574,N_16686);
xor U23817 (N_23817,N_13046,N_14470);
and U23818 (N_23818,N_19120,N_18867);
xnor U23819 (N_23819,N_14410,N_10532);
and U23820 (N_23820,N_12163,N_10562);
nand U23821 (N_23821,N_11275,N_11364);
nand U23822 (N_23822,N_13252,N_11987);
or U23823 (N_23823,N_17771,N_14708);
or U23824 (N_23824,N_14774,N_17516);
and U23825 (N_23825,N_19422,N_16996);
or U23826 (N_23826,N_12780,N_17830);
xnor U23827 (N_23827,N_14263,N_10056);
or U23828 (N_23828,N_15406,N_11465);
nor U23829 (N_23829,N_13548,N_19722);
xnor U23830 (N_23830,N_16903,N_14765);
xnor U23831 (N_23831,N_10686,N_17146);
and U23832 (N_23832,N_11531,N_12978);
xnor U23833 (N_23833,N_14941,N_11720);
or U23834 (N_23834,N_14004,N_17787);
nand U23835 (N_23835,N_18753,N_17122);
and U23836 (N_23836,N_16049,N_17732);
or U23837 (N_23837,N_15329,N_19132);
xnor U23838 (N_23838,N_12452,N_17606);
xor U23839 (N_23839,N_13835,N_19309);
nand U23840 (N_23840,N_14050,N_10764);
nor U23841 (N_23841,N_18133,N_13250);
or U23842 (N_23842,N_15213,N_16731);
and U23843 (N_23843,N_11427,N_10659);
and U23844 (N_23844,N_18308,N_18791);
and U23845 (N_23845,N_18804,N_13573);
nand U23846 (N_23846,N_14974,N_15245);
or U23847 (N_23847,N_14322,N_12605);
xor U23848 (N_23848,N_12147,N_17780);
nand U23849 (N_23849,N_19951,N_12320);
xor U23850 (N_23850,N_17820,N_14490);
or U23851 (N_23851,N_10851,N_15884);
nor U23852 (N_23852,N_14856,N_18175);
xnor U23853 (N_23853,N_16710,N_16733);
and U23854 (N_23854,N_12187,N_18267);
nor U23855 (N_23855,N_15472,N_16867);
nand U23856 (N_23856,N_19548,N_15647);
nand U23857 (N_23857,N_14885,N_11990);
nand U23858 (N_23858,N_16378,N_12483);
xnor U23859 (N_23859,N_16189,N_16329);
or U23860 (N_23860,N_14070,N_12266);
nor U23861 (N_23861,N_15463,N_19591);
nor U23862 (N_23862,N_10182,N_15270);
xnor U23863 (N_23863,N_14536,N_13009);
xor U23864 (N_23864,N_10791,N_19665);
and U23865 (N_23865,N_16390,N_14779);
and U23866 (N_23866,N_18892,N_17019);
nand U23867 (N_23867,N_15269,N_19418);
xnor U23868 (N_23868,N_14002,N_18780);
nand U23869 (N_23869,N_16560,N_12507);
and U23870 (N_23870,N_11198,N_15637);
and U23871 (N_23871,N_17119,N_13460);
and U23872 (N_23872,N_14539,N_16208);
and U23873 (N_23873,N_11602,N_14858);
nand U23874 (N_23874,N_19878,N_18487);
nor U23875 (N_23875,N_18628,N_18440);
xnor U23876 (N_23876,N_17894,N_17201);
nor U23877 (N_23877,N_11596,N_11229);
nor U23878 (N_23878,N_16648,N_16550);
nand U23879 (N_23879,N_12466,N_15632);
nor U23880 (N_23880,N_15280,N_13489);
nand U23881 (N_23881,N_12306,N_11891);
nand U23882 (N_23882,N_11898,N_19633);
xnor U23883 (N_23883,N_17584,N_10711);
nand U23884 (N_23884,N_14110,N_19585);
xor U23885 (N_23885,N_13526,N_11984);
nor U23886 (N_23886,N_10458,N_15368);
nand U23887 (N_23887,N_17990,N_13621);
xor U23888 (N_23888,N_11558,N_11116);
xnor U23889 (N_23889,N_18930,N_16803);
or U23890 (N_23890,N_10553,N_15265);
nor U23891 (N_23891,N_12391,N_15143);
xor U23892 (N_23892,N_15008,N_12077);
or U23893 (N_23893,N_15312,N_12900);
xnor U23894 (N_23894,N_19673,N_18188);
xnor U23895 (N_23895,N_11568,N_11830);
or U23896 (N_23896,N_13035,N_15805);
or U23897 (N_23897,N_11721,N_17751);
nor U23898 (N_23898,N_17054,N_12665);
and U23899 (N_23899,N_14426,N_10444);
xnor U23900 (N_23900,N_13670,N_17296);
and U23901 (N_23901,N_10369,N_13864);
or U23902 (N_23902,N_14338,N_18612);
or U23903 (N_23903,N_11394,N_12652);
nor U23904 (N_23904,N_14296,N_11832);
nor U23905 (N_23905,N_11018,N_16105);
xnor U23906 (N_23906,N_17448,N_16033);
xnor U23907 (N_23907,N_15872,N_12252);
nand U23908 (N_23908,N_15509,N_11396);
or U23909 (N_23909,N_15217,N_18414);
and U23910 (N_23910,N_15913,N_11496);
or U23911 (N_23911,N_17619,N_15454);
and U23912 (N_23912,N_13994,N_13580);
or U23913 (N_23913,N_15266,N_15829);
and U23914 (N_23914,N_14648,N_18081);
xnor U23915 (N_23915,N_13280,N_16424);
and U23916 (N_23916,N_16240,N_19381);
nor U23917 (N_23917,N_18622,N_13408);
xor U23918 (N_23918,N_15260,N_16220);
or U23919 (N_23919,N_19276,N_13579);
and U23920 (N_23920,N_11513,N_19512);
nand U23921 (N_23921,N_17864,N_16259);
and U23922 (N_23922,N_13452,N_14348);
or U23923 (N_23923,N_10357,N_11798);
nand U23924 (N_23924,N_11248,N_15016);
nand U23925 (N_23925,N_19065,N_17683);
nand U23926 (N_23926,N_17288,N_15247);
nor U23927 (N_23927,N_15585,N_17005);
or U23928 (N_23928,N_14848,N_16652);
and U23929 (N_23929,N_18354,N_15650);
nor U23930 (N_23930,N_14559,N_16101);
and U23931 (N_23931,N_19319,N_10332);
or U23932 (N_23932,N_16959,N_19664);
nand U23933 (N_23933,N_16317,N_12395);
nor U23934 (N_23934,N_17676,N_19108);
xnor U23935 (N_23935,N_15283,N_14704);
nor U23936 (N_23936,N_15900,N_11199);
nor U23937 (N_23937,N_15766,N_17728);
nand U23938 (N_23938,N_14978,N_11153);
nor U23939 (N_23939,N_18660,N_15695);
and U23940 (N_23940,N_16335,N_15447);
nor U23941 (N_23941,N_19278,N_14540);
nor U23942 (N_23942,N_17320,N_19962);
xnor U23943 (N_23943,N_18193,N_14815);
xnor U23944 (N_23944,N_10032,N_16515);
and U23945 (N_23945,N_16612,N_18265);
nand U23946 (N_23946,N_16409,N_16658);
or U23947 (N_23947,N_18996,N_12133);
xnor U23948 (N_23948,N_10014,N_19380);
nand U23949 (N_23949,N_18158,N_12911);
or U23950 (N_23950,N_11880,N_15469);
xnor U23951 (N_23951,N_10783,N_10165);
nand U23952 (N_23952,N_15445,N_15372);
nand U23953 (N_23953,N_16338,N_14813);
xnor U23954 (N_23954,N_10210,N_13189);
xnor U23955 (N_23955,N_19754,N_16989);
xor U23956 (N_23956,N_18012,N_10121);
or U23957 (N_23957,N_19568,N_11166);
nor U23958 (N_23958,N_19853,N_17480);
nor U23959 (N_23959,N_13704,N_12079);
and U23960 (N_23960,N_16949,N_13349);
nand U23961 (N_23961,N_13119,N_17089);
and U23962 (N_23962,N_18829,N_10072);
or U23963 (N_23963,N_11235,N_17397);
and U23964 (N_23964,N_16366,N_19394);
and U23965 (N_23965,N_16974,N_17853);
xor U23966 (N_23966,N_12586,N_17029);
nor U23967 (N_23967,N_11333,N_12710);
or U23968 (N_23968,N_17232,N_10232);
nand U23969 (N_23969,N_19490,N_10505);
nor U23970 (N_23970,N_11706,N_15733);
nand U23971 (N_23971,N_11085,N_17763);
or U23972 (N_23972,N_11667,N_19576);
or U23973 (N_23973,N_13315,N_17445);
nand U23974 (N_23974,N_10454,N_10424);
xor U23975 (N_23975,N_14777,N_10594);
and U23976 (N_23976,N_15044,N_15309);
xnor U23977 (N_23977,N_12286,N_13538);
xnor U23978 (N_23978,N_10316,N_18819);
nor U23979 (N_23979,N_16629,N_13763);
xor U23980 (N_23980,N_12783,N_15640);
nand U23981 (N_23981,N_16426,N_18154);
and U23982 (N_23982,N_19614,N_17565);
or U23983 (N_23983,N_16040,N_10549);
xnor U23984 (N_23984,N_12821,N_15911);
or U23985 (N_23985,N_16693,N_10799);
and U23986 (N_23986,N_14991,N_11440);
xor U23987 (N_23987,N_12596,N_16069);
and U23988 (N_23988,N_10283,N_11163);
nand U23989 (N_23989,N_14852,N_13402);
and U23990 (N_23990,N_10054,N_12557);
xnor U23991 (N_23991,N_14014,N_17033);
or U23992 (N_23992,N_10273,N_11132);
and U23993 (N_23993,N_10769,N_15300);
nor U23994 (N_23994,N_14224,N_12933);
nand U23995 (N_23995,N_14404,N_14374);
or U23996 (N_23996,N_11055,N_19770);
nor U23997 (N_23997,N_12347,N_12462);
xor U23998 (N_23998,N_14037,N_11666);
and U23999 (N_23999,N_15916,N_11472);
nor U24000 (N_24000,N_17998,N_10846);
nor U24001 (N_24001,N_16475,N_11243);
nor U24002 (N_24002,N_11435,N_12815);
xnor U24003 (N_24003,N_19082,N_16442);
nor U24004 (N_24004,N_12208,N_12048);
xor U24005 (N_24005,N_16854,N_16503);
xor U24006 (N_24006,N_15189,N_18071);
and U24007 (N_24007,N_11301,N_19994);
and U24008 (N_24008,N_14637,N_15735);
or U24009 (N_24009,N_10692,N_15299);
xor U24010 (N_24010,N_15648,N_19519);
xnor U24011 (N_24011,N_19238,N_15388);
or U24012 (N_24012,N_12145,N_13866);
xor U24013 (N_24013,N_14584,N_19513);
nor U24014 (N_24014,N_19221,N_18391);
or U24015 (N_24015,N_19468,N_11936);
and U24016 (N_24016,N_16774,N_13578);
nand U24017 (N_24017,N_14653,N_19006);
and U24018 (N_24018,N_16215,N_18057);
nand U24019 (N_24019,N_17126,N_17579);
xnor U24020 (N_24020,N_10112,N_12973);
and U24021 (N_24021,N_12798,N_12127);
xnor U24022 (N_24022,N_19988,N_18763);
xnor U24023 (N_24023,N_19764,N_16911);
or U24024 (N_24024,N_11998,N_13176);
and U24025 (N_24025,N_10803,N_12852);
or U24026 (N_24026,N_19041,N_10863);
nor U24027 (N_24027,N_14825,N_10778);
nor U24028 (N_24028,N_13449,N_13206);
or U24029 (N_24029,N_13897,N_18632);
xnor U24030 (N_24030,N_16030,N_16765);
nand U24031 (N_24031,N_12278,N_11638);
and U24032 (N_24032,N_13382,N_10380);
and U24033 (N_24033,N_19331,N_15048);
nor U24034 (N_24034,N_17803,N_11278);
and U24035 (N_24035,N_16155,N_14324);
nand U24036 (N_24036,N_18994,N_13121);
xnor U24037 (N_24037,N_18194,N_19506);
or U24038 (N_24038,N_14200,N_14089);
or U24039 (N_24039,N_16009,N_12049);
or U24040 (N_24040,N_11494,N_13689);
nor U24041 (N_24041,N_17723,N_12962);
xor U24042 (N_24042,N_12585,N_12981);
nand U24043 (N_24043,N_12458,N_17028);
nand U24044 (N_24044,N_14548,N_16822);
or U24045 (N_24045,N_15429,N_16711);
nand U24046 (N_24046,N_13929,N_14914);
xnor U24047 (N_24047,N_19580,N_18458);
xor U24048 (N_24048,N_17533,N_18413);
and U24049 (N_24049,N_14227,N_12687);
nor U24050 (N_24050,N_15618,N_19223);
or U24051 (N_24051,N_19174,N_10757);
and U24052 (N_24052,N_18143,N_15979);
nand U24053 (N_24053,N_10410,N_17329);
nand U24054 (N_24054,N_10883,N_12070);
or U24055 (N_24055,N_13728,N_18344);
and U24056 (N_24056,N_19790,N_10637);
xnor U24057 (N_24057,N_18307,N_15236);
xnor U24058 (N_24058,N_16360,N_12662);
and U24059 (N_24059,N_16829,N_17776);
or U24060 (N_24060,N_15168,N_19798);
and U24061 (N_24061,N_10734,N_11411);
nand U24062 (N_24062,N_11978,N_11503);
nand U24063 (N_24063,N_14225,N_17350);
nand U24064 (N_24064,N_10767,N_17295);
and U24065 (N_24065,N_18656,N_13409);
xor U24066 (N_24066,N_13962,N_10870);
nor U24067 (N_24067,N_19471,N_11946);
nand U24068 (N_24068,N_17243,N_19068);
and U24069 (N_24069,N_14581,N_15625);
xor U24070 (N_24070,N_10962,N_18505);
and U24071 (N_24071,N_15261,N_14400);
nor U24072 (N_24072,N_18961,N_10876);
and U24073 (N_24073,N_12330,N_12205);
or U24074 (N_24074,N_10346,N_13195);
or U24075 (N_24075,N_18850,N_19073);
xor U24076 (N_24076,N_14396,N_14514);
nand U24077 (N_24077,N_16697,N_16465);
xor U24078 (N_24078,N_19356,N_18750);
or U24079 (N_24079,N_11317,N_19096);
xnor U24080 (N_24080,N_17258,N_15553);
or U24081 (N_24081,N_15965,N_16035);
nor U24082 (N_24082,N_18264,N_15694);
and U24083 (N_24083,N_13115,N_12107);
and U24084 (N_24084,N_19083,N_13234);
nand U24085 (N_24085,N_19531,N_16348);
and U24086 (N_24086,N_11032,N_12677);
nor U24087 (N_24087,N_15816,N_15211);
or U24088 (N_24088,N_16147,N_15670);
nor U24089 (N_24089,N_10575,N_18925);
xor U24090 (N_24090,N_10722,N_15547);
nand U24091 (N_24091,N_19122,N_17770);
nor U24092 (N_24092,N_19291,N_17070);
nor U24093 (N_24093,N_14679,N_14698);
or U24094 (N_24094,N_12092,N_10005);
or U24095 (N_24095,N_15642,N_18320);
xor U24096 (N_24096,N_19100,N_13163);
xor U24097 (N_24097,N_18947,N_13447);
nor U24098 (N_24098,N_14117,N_19676);
xor U24099 (N_24099,N_15491,N_12876);
and U24100 (N_24100,N_13028,N_16288);
nand U24101 (N_24101,N_17996,N_13094);
xnor U24102 (N_24102,N_11715,N_11567);
nor U24103 (N_24103,N_13112,N_15297);
nor U24104 (N_24104,N_10961,N_19589);
or U24105 (N_24105,N_16053,N_16397);
or U24106 (N_24106,N_12681,N_17888);
nor U24107 (N_24107,N_13396,N_12342);
nor U24108 (N_24108,N_13245,N_16013);
and U24109 (N_24109,N_15381,N_13946);
or U24110 (N_24110,N_11779,N_14841);
and U24111 (N_24111,N_10896,N_12893);
nand U24112 (N_24112,N_12932,N_17718);
nor U24113 (N_24113,N_18202,N_10684);
and U24114 (N_24114,N_18762,N_13999);
xnor U24115 (N_24115,N_16191,N_15123);
and U24116 (N_24116,N_15047,N_12106);
xnor U24117 (N_24117,N_18334,N_16990);
and U24118 (N_24118,N_10028,N_10320);
nor U24119 (N_24119,N_11996,N_18018);
nor U24120 (N_24120,N_11368,N_12956);
nor U24121 (N_24121,N_10249,N_19061);
nor U24122 (N_24122,N_11343,N_14298);
or U24123 (N_24123,N_17768,N_16261);
nand U24124 (N_24124,N_15037,N_18381);
nand U24125 (N_24125,N_15960,N_15707);
or U24126 (N_24126,N_17491,N_16356);
nand U24127 (N_24127,N_12080,N_11758);
nand U24128 (N_24128,N_17828,N_12455);
nor U24129 (N_24129,N_12751,N_17128);
xor U24130 (N_24130,N_10578,N_16896);
nand U24131 (N_24131,N_11702,N_10914);
and U24132 (N_24132,N_19775,N_14241);
xnor U24133 (N_24133,N_10389,N_10732);
nand U24134 (N_24134,N_16582,N_19078);
nor U24135 (N_24135,N_16265,N_17581);
nand U24136 (N_24136,N_12921,N_17171);
xor U24137 (N_24137,N_12648,N_13813);
or U24138 (N_24138,N_18439,N_15433);
nor U24139 (N_24139,N_13561,N_11037);
nor U24140 (N_24140,N_14289,N_12515);
nor U24141 (N_24141,N_15671,N_15178);
nor U24142 (N_24142,N_15343,N_16393);
or U24143 (N_24143,N_18362,N_15956);
xor U24144 (N_24144,N_11359,N_18070);
and U24145 (N_24145,N_13738,N_13461);
or U24146 (N_24146,N_13769,N_18553);
xnor U24147 (N_24147,N_17617,N_18919);
or U24148 (N_24148,N_15758,N_17242);
and U24149 (N_24149,N_19413,N_18030);
or U24150 (N_24150,N_19454,N_13802);
or U24151 (N_24151,N_16160,N_15328);
nor U24152 (N_24152,N_13003,N_16375);
nor U24153 (N_24153,N_19346,N_17214);
and U24154 (N_24154,N_16957,N_12545);
or U24155 (N_24155,N_17365,N_12224);
nor U24156 (N_24156,N_13698,N_17993);
xnor U24157 (N_24157,N_10081,N_10809);
or U24158 (N_24158,N_14961,N_15287);
xor U24159 (N_24159,N_15232,N_13244);
nor U24160 (N_24160,N_12778,N_16622);
or U24161 (N_24161,N_11239,N_11466);
nor U24162 (N_24162,N_18601,N_19085);
nand U24163 (N_24163,N_19975,N_10825);
or U24164 (N_24164,N_14409,N_17402);
xor U24165 (N_24165,N_18637,N_13324);
nor U24166 (N_24166,N_12310,N_13337);
xor U24167 (N_24167,N_16212,N_13087);
or U24168 (N_24168,N_10365,N_18927);
xor U24169 (N_24169,N_11504,N_16061);
nand U24170 (N_24170,N_16109,N_10111);
and U24171 (N_24171,N_11802,N_11253);
xor U24172 (N_24172,N_10107,N_12363);
xnor U24173 (N_24173,N_12231,N_13187);
xnor U24174 (N_24174,N_19521,N_11537);
nand U24175 (N_24175,N_19978,N_18597);
xnor U24176 (N_24176,N_14830,N_12696);
xnor U24177 (N_24177,N_16525,N_12496);
xor U24178 (N_24178,N_10605,N_18310);
nand U24179 (N_24179,N_14534,N_15931);
nand U24180 (N_24180,N_13400,N_11840);
or U24181 (N_24181,N_18340,N_18728);
xor U24182 (N_24182,N_17774,N_19835);
or U24183 (N_24183,N_16691,N_19196);
nor U24184 (N_24184,N_15051,N_17777);
nor U24185 (N_24185,N_18148,N_12319);
xor U24186 (N_24186,N_13322,N_16958);
nor U24187 (N_24187,N_13309,N_16385);
xnor U24188 (N_24188,N_13490,N_16293);
nand U24189 (N_24189,N_16687,N_18488);
or U24190 (N_24190,N_16856,N_19398);
nand U24191 (N_24191,N_19899,N_19846);
xnor U24192 (N_24192,N_14523,N_15335);
nand U24193 (N_24193,N_10733,N_17677);
and U24194 (N_24194,N_19119,N_17660);
or U24195 (N_24195,N_15267,N_10533);
nand U24196 (N_24196,N_13959,N_15841);
or U24197 (N_24197,N_14680,N_13164);
xor U24198 (N_24198,N_11309,N_17324);
or U24199 (N_24199,N_11768,N_18474);
and U24200 (N_24200,N_18236,N_10612);
nor U24201 (N_24201,N_14667,N_12566);
or U24202 (N_24202,N_18024,N_10012);
xor U24203 (N_24203,N_17293,N_11587);
nand U24204 (N_24204,N_10960,N_11591);
or U24205 (N_24205,N_14790,N_12739);
or U24206 (N_24206,N_15293,N_10509);
nor U24207 (N_24207,N_14341,N_15510);
or U24208 (N_24208,N_18055,N_15636);
or U24209 (N_24209,N_14867,N_19791);
nor U24210 (N_24210,N_17793,N_10824);
nor U24211 (N_24211,N_18644,N_14622);
nand U24212 (N_24212,N_12593,N_11070);
or U24213 (N_24213,N_11433,N_17654);
or U24214 (N_24214,N_12574,N_11770);
and U24215 (N_24215,N_17984,N_19106);
and U24216 (N_24216,N_17905,N_18328);
and U24217 (N_24217,N_16927,N_14809);
nor U24218 (N_24218,N_19127,N_11901);
xor U24219 (N_24219,N_13734,N_11669);
or U24220 (N_24220,N_14556,N_14745);
nand U24221 (N_24221,N_19035,N_12099);
nor U24222 (N_24222,N_13488,N_10648);
and U24223 (N_24223,N_14719,N_12336);
xor U24224 (N_24224,N_14931,N_12061);
xnor U24225 (N_24225,N_13481,N_16614);
and U24226 (N_24226,N_15594,N_14339);
xor U24227 (N_24227,N_11750,N_14518);
xnor U24228 (N_24228,N_18797,N_10657);
and U24229 (N_24229,N_16767,N_13540);
nor U24230 (N_24230,N_15490,N_10672);
nor U24231 (N_24231,N_16926,N_19943);
xnor U24232 (N_24232,N_12906,N_12599);
or U24233 (N_24233,N_17568,N_16527);
nor U24234 (N_24234,N_11945,N_17451);
xnor U24235 (N_24235,N_19807,N_19339);
and U24236 (N_24236,N_11481,N_19024);
xor U24237 (N_24237,N_16171,N_12055);
nand U24238 (N_24238,N_14645,N_12476);
nor U24239 (N_24239,N_19689,N_18510);
nor U24240 (N_24240,N_18182,N_14900);
nand U24241 (N_24241,N_11628,N_16011);
nor U24242 (N_24242,N_11507,N_15197);
xnor U24243 (N_24243,N_13591,N_14304);
xor U24244 (N_24244,N_10936,N_11254);
xor U24245 (N_24245,N_15257,N_16706);
nor U24246 (N_24246,N_13383,N_15357);
and U24247 (N_24247,N_19965,N_16607);
nor U24248 (N_24248,N_14028,N_11240);
and U24249 (N_24249,N_12953,N_14091);
nor U24250 (N_24250,N_16073,N_18735);
nand U24251 (N_24251,N_17279,N_10438);
nand U24252 (N_24252,N_13885,N_11335);
nand U24253 (N_24253,N_18986,N_14694);
nand U24254 (N_24254,N_19270,N_15160);
or U24255 (N_24255,N_10731,N_12176);
nand U24256 (N_24256,N_19058,N_10452);
xnor U24257 (N_24257,N_14623,N_13438);
xor U24258 (N_24258,N_12958,N_12038);
nor U24259 (N_24259,N_14851,N_18539);
and U24260 (N_24260,N_13231,N_10658);
or U24261 (N_24261,N_11451,N_16276);
nor U24262 (N_24262,N_13787,N_13270);
or U24263 (N_24263,N_11529,N_15439);
nor U24264 (N_24264,N_10864,N_19323);
and U24265 (N_24265,N_19719,N_13213);
nor U24266 (N_24266,N_17981,N_14486);
and U24267 (N_24267,N_13290,N_12116);
or U24268 (N_24268,N_18373,N_17563);
nand U24269 (N_24269,N_19934,N_12219);
or U24270 (N_24270,N_14971,N_16186);
xor U24271 (N_24271,N_10057,N_11414);
nor U24272 (N_24272,N_16131,N_11693);
and U24273 (N_24273,N_18491,N_10303);
nand U24274 (N_24274,N_17330,N_12000);
nand U24275 (N_24275,N_14085,N_16619);
nand U24276 (N_24276,N_10788,N_14447);
and U24277 (N_24277,N_15798,N_19171);
xor U24278 (N_24278,N_10471,N_15657);
nor U24279 (N_24279,N_12863,N_10350);
nand U24280 (N_24280,N_17587,N_11761);
nor U24281 (N_24281,N_17120,N_11281);
nand U24282 (N_24282,N_17912,N_10117);
xor U24283 (N_24283,N_11028,N_17268);
nor U24284 (N_24284,N_10334,N_16164);
and U24285 (N_24285,N_10504,N_16532);
nor U24286 (N_24286,N_16015,N_16685);
and U24287 (N_24287,N_17957,N_10327);
and U24288 (N_24288,N_16042,N_14846);
xnor U24289 (N_24289,N_19016,N_16067);
and U24290 (N_24290,N_11242,N_10087);
or U24291 (N_24291,N_12797,N_17860);
nor U24292 (N_24292,N_15311,N_19640);
nor U24293 (N_24293,N_11397,N_16537);
and U24294 (N_24294,N_17665,N_17978);
nand U24295 (N_24295,N_12691,N_18443);
nand U24296 (N_24296,N_10496,N_12732);
and U24297 (N_24297,N_10070,N_16952);
xnor U24298 (N_24298,N_12832,N_10470);
and U24299 (N_24299,N_11449,N_14922);
and U24300 (N_24300,N_19774,N_17048);
nor U24301 (N_24301,N_10700,N_17406);
or U24302 (N_24302,N_15554,N_14640);
or U24303 (N_24303,N_10203,N_19461);
xor U24304 (N_24304,N_11918,N_10002);
nor U24305 (N_24305,N_11924,N_15225);
xnor U24306 (N_24306,N_15142,N_14860);
xor U24307 (N_24307,N_12188,N_14101);
xor U24308 (N_24308,N_12263,N_16918);
or U24309 (N_24309,N_16943,N_17880);
and U24310 (N_24310,N_16545,N_14344);
nand U24311 (N_24311,N_15837,N_13624);
or U24312 (N_24312,N_10784,N_12674);
xnor U24313 (N_24313,N_13757,N_10435);
or U24314 (N_24314,N_16627,N_19098);
or U24315 (N_24315,N_18764,N_16805);
nor U24316 (N_24316,N_14283,N_17393);
nand U24317 (N_24317,N_15121,N_19292);
xor U24318 (N_24318,N_19406,N_11919);
nor U24319 (N_24319,N_17742,N_11631);
xor U24320 (N_24320,N_18934,N_15275);
xnor U24321 (N_24321,N_11071,N_14015);
nand U24322 (N_24322,N_13652,N_15239);
nand U24323 (N_24323,N_15504,N_17526);
xor U24324 (N_24324,N_14259,N_15195);
and U24325 (N_24325,N_18023,N_14689);
nor U24326 (N_24326,N_17979,N_17067);
nor U24327 (N_24327,N_14651,N_12769);
or U24328 (N_24328,N_18452,N_19583);
xnor U24329 (N_24329,N_17992,N_19959);
or U24330 (N_24330,N_16823,N_10335);
or U24331 (N_24331,N_12078,N_14723);
or U24332 (N_24332,N_10472,N_19220);
or U24333 (N_24333,N_15403,N_14132);
nand U24334 (N_24334,N_18238,N_15310);
and U24335 (N_24335,N_13731,N_12114);
nor U24336 (N_24336,N_12206,N_12891);
or U24337 (N_24337,N_19014,N_18607);
or U24338 (N_24338,N_15459,N_14233);
nor U24339 (N_24339,N_14080,N_18676);
and U24340 (N_24340,N_16091,N_15199);
nor U24341 (N_24341,N_14065,N_12928);
nor U24342 (N_24342,N_17679,N_12895);
nand U24343 (N_24343,N_19204,N_15363);
or U24344 (N_24344,N_13775,N_14236);
or U24345 (N_24345,N_11405,N_14706);
nor U24346 (N_24346,N_15502,N_18573);
or U24347 (N_24347,N_13384,N_18036);
and U24348 (N_24348,N_11655,N_17347);
nand U24349 (N_24349,N_10564,N_14210);
or U24350 (N_24350,N_12737,N_12450);
xor U24351 (N_24351,N_15413,N_10584);
and U24352 (N_24352,N_19388,N_16115);
or U24353 (N_24353,N_16517,N_11415);
nor U24354 (N_24354,N_18693,N_19843);
or U24355 (N_24355,N_17986,N_11890);
nand U24356 (N_24356,N_16289,N_13589);
and U24357 (N_24357,N_16032,N_10715);
and U24358 (N_24358,N_15383,N_15481);
xnor U24359 (N_24359,N_14390,N_12244);
nand U24360 (N_24360,N_10047,N_11751);
xnor U24361 (N_24361,N_10753,N_19666);
and U24362 (N_24362,N_10030,N_18896);
xnor U24363 (N_24363,N_13451,N_19558);
nor U24364 (N_24364,N_15877,N_19560);
nor U24365 (N_24365,N_15616,N_14570);
nor U24366 (N_24366,N_13612,N_19213);
xnor U24367 (N_24367,N_19639,N_15895);
xor U24368 (N_24368,N_13966,N_13171);
and U24369 (N_24369,N_11523,N_18261);
nand U24370 (N_24370,N_19894,N_14082);
nor U24371 (N_24371,N_12717,N_11473);
or U24372 (N_24372,N_12314,N_12537);
xor U24373 (N_24373,N_19904,N_14142);
nand U24374 (N_24374,N_16889,N_17269);
and U24375 (N_24375,N_11162,N_17443);
nand U24376 (N_24376,N_17589,N_15457);
nand U24377 (N_24377,N_16827,N_17832);
and U24378 (N_24378,N_19570,N_14450);
nor U24379 (N_24379,N_18702,N_14923);
and U24380 (N_24380,N_12714,N_13575);
nor U24381 (N_24381,N_15331,N_17788);
and U24382 (N_24382,N_13020,N_17872);
xnor U24383 (N_24383,N_18445,N_19301);
nor U24384 (N_24384,N_16318,N_18480);
nor U24385 (N_24385,N_10250,N_15298);
or U24386 (N_24386,N_13256,N_17615);
or U24387 (N_24387,N_14234,N_11863);
nand U24388 (N_24388,N_15337,N_13407);
xor U24389 (N_24389,N_19203,N_10337);
xor U24390 (N_24390,N_19439,N_11009);
or U24391 (N_24391,N_10265,N_10448);
or U24392 (N_24392,N_18365,N_15345);
and U24393 (N_24393,N_11462,N_15857);
and U24394 (N_24394,N_11828,N_10679);
xor U24395 (N_24395,N_15422,N_10570);
nor U24396 (N_24396,N_10149,N_11025);
xor U24397 (N_24397,N_11030,N_19093);
nand U24398 (N_24398,N_16277,N_12630);
or U24399 (N_24399,N_12750,N_14627);
nor U24400 (N_24400,N_13182,N_17440);
and U24401 (N_24401,N_13945,N_16021);
or U24402 (N_24402,N_11135,N_19304);
or U24403 (N_24403,N_17716,N_15653);
nand U24404 (N_24404,N_13100,N_15542);
or U24405 (N_24405,N_13637,N_14589);
and U24406 (N_24406,N_11771,N_14124);
and U24407 (N_24407,N_19055,N_13141);
and U24408 (N_24408,N_14239,N_13097);
xor U24409 (N_24409,N_11455,N_13511);
and U24410 (N_24410,N_18679,N_13360);
or U24411 (N_24411,N_18695,N_17651);
nand U24412 (N_24412,N_14956,N_19715);
nand U24413 (N_24413,N_18945,N_15999);
and U24414 (N_24414,N_11952,N_11136);
xnor U24415 (N_24415,N_12164,N_12748);
xnor U24416 (N_24416,N_10307,N_12636);
xor U24417 (N_24417,N_14195,N_12942);
xnor U24418 (N_24418,N_15523,N_17032);
and U24419 (N_24419,N_17007,N_16325);
xor U24420 (N_24420,N_13379,N_17271);
or U24421 (N_24421,N_11056,N_15939);
nor U24422 (N_24422,N_12264,N_18438);
or U24423 (N_24423,N_10405,N_11705);
and U24424 (N_24424,N_12569,N_12877);
nor U24425 (N_24425,N_15059,N_10084);
nor U24426 (N_24426,N_15050,N_18738);
xnor U24427 (N_24427,N_13154,N_19656);
nand U24428 (N_24428,N_12829,N_14459);
and U24429 (N_24429,N_19286,N_14469);
and U24430 (N_24430,N_18419,N_12857);
xnor U24431 (N_24431,N_14530,N_17585);
xor U24432 (N_24432,N_10808,N_15823);
nand U24433 (N_24433,N_18653,N_19436);
or U24434 (N_24434,N_13979,N_15190);
nor U24435 (N_24435,N_16498,N_13005);
xnor U24436 (N_24436,N_11756,N_18284);
and U24437 (N_24437,N_18920,N_14349);
and U24438 (N_24438,N_11099,N_14445);
nor U24439 (N_24439,N_11932,N_12042);
xnor U24440 (N_24440,N_17053,N_18937);
nand U24441 (N_24441,N_14270,N_17164);
and U24442 (N_24442,N_13854,N_13450);
xnor U24443 (N_24443,N_11324,N_14638);
or U24444 (N_24444,N_19810,N_13073);
xor U24445 (N_24445,N_13546,N_13838);
or U24446 (N_24446,N_12260,N_11138);
xor U24447 (N_24447,N_18718,N_17866);
or U24448 (N_24448,N_19979,N_13644);
nor U24449 (N_24449,N_10710,N_14146);
xnor U24450 (N_24450,N_13074,N_18270);
xnor U24451 (N_24451,N_19245,N_14582);
or U24452 (N_24452,N_12014,N_13650);
nor U24453 (N_24453,N_12396,N_10780);
xnor U24454 (N_24454,N_18449,N_11617);
xor U24455 (N_24455,N_16372,N_18286);
nor U24456 (N_24456,N_12937,N_15545);
nand U24457 (N_24457,N_15833,N_15524);
nor U24458 (N_24458,N_15959,N_12059);
xnor U24459 (N_24459,N_18658,N_11314);
and U24460 (N_24460,N_15586,N_19250);
or U24461 (N_24461,N_18051,N_18922);
xor U24462 (N_24462,N_13799,N_12792);
nand U24463 (N_24463,N_13002,N_10690);
and U24464 (N_24464,N_15206,N_17931);
or U24465 (N_24465,N_15686,N_15820);
xor U24466 (N_24466,N_11320,N_15714);
and U24467 (N_24467,N_16770,N_17392);
xor U24468 (N_24468,N_18512,N_13800);
nand U24469 (N_24469,N_18977,N_10476);
xnor U24470 (N_24470,N_12290,N_19742);
xor U24471 (N_24471,N_16351,N_16859);
xnor U24472 (N_24472,N_12169,N_19297);
nor U24473 (N_24473,N_18746,N_17569);
and U24474 (N_24474,N_10877,N_12505);
nor U24475 (N_24475,N_19520,N_15595);
nand U24476 (N_24476,N_16938,N_16786);
and U24477 (N_24477,N_11543,N_13912);
nand U24478 (N_24478,N_10677,N_19160);
nor U24479 (N_24479,N_11334,N_18123);
nor U24480 (N_24480,N_13069,N_12834);
xor U24481 (N_24481,N_19069,N_16665);
nand U24482 (N_24482,N_15024,N_15741);
and U24483 (N_24483,N_13556,N_15888);
and U24484 (N_24484,N_11152,N_19897);
or U24485 (N_24485,N_11792,N_19662);
xor U24486 (N_24486,N_17626,N_15323);
and U24487 (N_24487,N_17346,N_19864);
or U24488 (N_24488,N_18725,N_13067);
nand U24489 (N_24489,N_13071,N_17136);
and U24490 (N_24490,N_15982,N_12553);
nor U24491 (N_24491,N_13295,N_18464);
or U24492 (N_24492,N_15038,N_12768);
and U24493 (N_24493,N_14881,N_16809);
nor U24494 (N_24494,N_17861,N_16877);
and U24495 (N_24495,N_12486,N_17522);
xnor U24496 (N_24496,N_17558,N_19110);
nor U24497 (N_24497,N_12872,N_13943);
nand U24498 (N_24498,N_10354,N_11249);
xor U24499 (N_24499,N_12573,N_13031);
xor U24500 (N_24500,N_14497,N_17300);
xor U24501 (N_24501,N_19768,N_13629);
or U24502 (N_24502,N_12531,N_18327);
and U24503 (N_24503,N_10373,N_11067);
or U24504 (N_24504,N_15743,N_14453);
nor U24505 (N_24505,N_16132,N_14394);
or U24506 (N_24506,N_18942,N_17419);
or U24507 (N_24507,N_12704,N_10315);
nand U24508 (N_24508,N_16359,N_18346);
xor U24509 (N_24509,N_17812,N_17999);
nor U24510 (N_24510,N_10144,N_11929);
nand U24511 (N_24511,N_14392,N_11691);
or U24512 (N_24512,N_17755,N_12577);
nand U24513 (N_24513,N_15705,N_15124);
or U24514 (N_24514,N_12995,N_16410);
xnor U24515 (N_24515,N_17100,N_19136);
or U24516 (N_24516,N_16520,N_18803);
nand U24517 (N_24517,N_17975,N_19616);
xnor U24518 (N_24518,N_16584,N_13868);
or U24519 (N_24519,N_13977,N_19587);
nand U24520 (N_24520,N_16538,N_13373);
nand U24521 (N_24521,N_16285,N_10463);
nand U24522 (N_24522,N_10295,N_12969);
nand U24523 (N_24523,N_19541,N_13445);
and U24524 (N_24524,N_17766,N_10355);
and U24525 (N_24525,N_17312,N_15203);
or U24526 (N_24526,N_12776,N_16055);
nand U24527 (N_24527,N_18885,N_19311);
or U24528 (N_24528,N_17786,N_18097);
or U24529 (N_24529,N_11680,N_11520);
xnor U24530 (N_24530,N_14160,N_12222);
nor U24531 (N_24531,N_14212,N_19062);
nand U24532 (N_24532,N_11497,N_19067);
nor U24533 (N_24533,N_14247,N_10247);
and U24534 (N_24534,N_14521,N_16546);
xor U24535 (N_24535,N_16430,N_18140);
or U24536 (N_24536,N_19990,N_12387);
and U24537 (N_24537,N_15151,N_15974);
nor U24538 (N_24538,N_13202,N_19423);
or U24539 (N_24539,N_12098,N_13086);
nand U24540 (N_24540,N_13342,N_17807);
nor U24541 (N_24541,N_19954,N_16698);
nor U24542 (N_24542,N_19737,N_13247);
and U24543 (N_24543,N_11580,N_13019);
and U24544 (N_24544,N_15033,N_18544);
nor U24545 (N_24545,N_17925,N_16196);
nor U24546 (N_24546,N_18817,N_14351);
nand U24547 (N_24547,N_14319,N_13956);
or U24548 (N_24548,N_11632,N_14742);
nand U24549 (N_24549,N_12946,N_11230);
nor U24550 (N_24550,N_14090,N_16159);
nor U24551 (N_24551,N_13279,N_15291);
and U24552 (N_24552,N_14783,N_15807);
and U24553 (N_24553,N_12564,N_16979);
and U24554 (N_24554,N_15193,N_17658);
xnor U24555 (N_24555,N_17405,N_15475);
or U24556 (N_24556,N_11332,N_12405);
nand U24557 (N_24557,N_17009,N_17639);
nand U24558 (N_24558,N_12949,N_19510);
nand U24559 (N_24559,N_15541,N_13246);
nand U24560 (N_24560,N_16454,N_19425);
and U24561 (N_24561,N_11813,N_18146);
xnor U24562 (N_24562,N_17644,N_17257);
and U24563 (N_24563,N_11781,N_12508);
nor U24564 (N_24564,N_17680,N_18879);
xnor U24565 (N_24565,N_16452,N_16179);
and U24566 (N_24566,N_12939,N_18181);
and U24567 (N_24567,N_16466,N_19415);
nand U24568 (N_24568,N_16962,N_16966);
xor U24569 (N_24569,N_18729,N_14477);
nor U24570 (N_24570,N_19430,N_13581);
or U24571 (N_24571,N_19874,N_12235);
nand U24572 (N_24572,N_18882,N_19246);
xnor U24573 (N_24573,N_12993,N_13492);
nand U24574 (N_24574,N_19482,N_12153);
nand U24575 (N_24575,N_16213,N_17260);
xor U24576 (N_24576,N_13093,N_18190);
or U24577 (N_24577,N_16072,N_15507);
or U24578 (N_24578,N_18336,N_14208);
and U24579 (N_24579,N_12520,N_17504);
or U24580 (N_24580,N_14690,N_10865);
or U24581 (N_24581,N_10108,N_15522);
xnor U24582 (N_24582,N_18629,N_11576);
nand U24583 (N_24583,N_11057,N_11027);
and U24584 (N_24584,N_19524,N_19642);
nor U24585 (N_24585,N_19762,N_10639);
nand U24586 (N_24586,N_11436,N_11689);
or U24587 (N_24587,N_15184,N_13936);
xor U24588 (N_24588,N_10604,N_16343);
nor U24589 (N_24589,N_14151,N_16075);
nor U24590 (N_24590,N_12082,N_10717);
xnor U24591 (N_24591,N_15165,N_11167);
nor U24592 (N_24592,N_12223,N_13096);
or U24593 (N_24593,N_16413,N_13649);
and U24594 (N_24594,N_15892,N_19538);
or U24595 (N_24595,N_10848,N_16524);
nand U24596 (N_24596,N_12122,N_19007);
or U24597 (N_24597,N_10145,N_16486);
xnor U24598 (N_24598,N_17006,N_12499);
nand U24599 (N_24599,N_10167,N_10450);
xnor U24600 (N_24600,N_15063,N_14909);
nor U24601 (N_24601,N_11110,N_17192);
or U24602 (N_24602,N_18398,N_12413);
xor U24603 (N_24603,N_17060,N_10244);
or U24604 (N_24604,N_11234,N_17963);
xnor U24605 (N_24605,N_10980,N_18549);
and U24606 (N_24606,N_15784,N_16349);
or U24607 (N_24607,N_17207,N_10076);
or U24608 (N_24608,N_16123,N_16983);
and U24609 (N_24609,N_15006,N_15485);
and U24610 (N_24610,N_15414,N_12839);
nand U24611 (N_24611,N_12567,N_18331);
and U24612 (N_24612,N_13893,N_19039);
nand U24613 (N_24613,N_19349,N_17695);
xnor U24614 (N_24614,N_16512,N_10364);
xnor U24615 (N_24615,N_19469,N_19330);
nor U24616 (N_24616,N_10126,N_17118);
nor U24617 (N_24617,N_11205,N_12341);
nor U24618 (N_24618,N_12812,N_14214);
nand U24619 (N_24619,N_14564,N_10762);
xor U24620 (N_24620,N_13876,N_17148);
and U24621 (N_24621,N_19470,N_10466);
and U24622 (N_24622,N_12217,N_12282);
xnor U24623 (N_24623,N_16125,N_18056);
nor U24624 (N_24624,N_13957,N_13357);
nand U24625 (N_24625,N_15127,N_10092);
nand U24626 (N_24626,N_12886,N_15155);
and U24627 (N_24627,N_18080,N_11399);
or U24628 (N_24628,N_18420,N_10125);
nor U24629 (N_24629,N_13272,N_17205);
nand U24630 (N_24630,N_13138,N_11120);
xnor U24631 (N_24631,N_17482,N_19444);
xor U24632 (N_24632,N_15611,N_10973);
xnor U24633 (N_24633,N_16811,N_12676);
or U24634 (N_24634,N_13401,N_11795);
nand U24635 (N_24635,N_16362,N_13852);
and U24636 (N_24636,N_14513,N_10403);
nor U24637 (N_24637,N_14602,N_15349);
or U24638 (N_24638,N_14823,N_14968);
or U24639 (N_24639,N_18747,N_19141);
nand U24640 (N_24640,N_19457,N_10428);
nand U24641 (N_24641,N_15340,N_13887);
and U24642 (N_24642,N_17455,N_17248);
nand U24643 (N_24643,N_12365,N_18155);
nor U24644 (N_24644,N_12810,N_13680);
or U24645 (N_24645,N_17416,N_11508);
and U24646 (N_24646,N_14562,N_14981);
xor U24647 (N_24647,N_13218,N_14524);
nand U24648 (N_24648,N_15556,N_18960);
nand U24649 (N_24649,N_15844,N_18554);
or U24650 (N_24650,N_15702,N_16144);
nor U24651 (N_24651,N_12111,N_17168);
xor U24652 (N_24652,N_15564,N_11882);
nand U24653 (N_24653,N_14462,N_13104);
or U24654 (N_24654,N_12343,N_16331);
xnor U24655 (N_24655,N_10391,N_17379);
nor U24656 (N_24656,N_10387,N_16108);
nor U24657 (N_24657,N_17321,N_11526);
xor U24658 (N_24658,N_16628,N_14532);
nor U24659 (N_24659,N_17599,N_17852);
nand U24660 (N_24660,N_15054,N_11327);
nand U24661 (N_24661,N_18580,N_12615);
or U24662 (N_24662,N_16638,N_16501);
and U24663 (N_24663,N_17305,N_13607);
nand U24664 (N_24664,N_16434,N_13013);
or U24665 (N_24665,N_17016,N_13677);
nor U24666 (N_24666,N_16449,N_14735);
nand U24667 (N_24667,N_16320,N_17230);
or U24668 (N_24668,N_12882,N_19668);
nand U24669 (N_24669,N_11257,N_13721);
nor U24670 (N_24670,N_17368,N_11822);
and U24671 (N_24671,N_15560,N_18040);
and U24672 (N_24672,N_15788,N_11061);
or U24673 (N_24673,N_18576,N_19779);
or U24674 (N_24674,N_15448,N_11142);
or U24675 (N_24675,N_15404,N_17109);
nor U24676 (N_24676,N_19976,N_10174);
nor U24677 (N_24677,N_18309,N_16136);
or U24678 (N_24678,N_19117,N_14441);
or U24679 (N_24679,N_17466,N_10237);
nand U24680 (N_24680,N_16510,N_16234);
and U24681 (N_24681,N_12719,N_19408);
xor U24682 (N_24682,N_10349,N_13456);
xnor U24683 (N_24683,N_11051,N_19974);
and U24684 (N_24684,N_14731,N_16724);
and U24685 (N_24685,N_14389,N_19721);
nor U24686 (N_24686,N_10932,N_19685);
or U24687 (N_24687,N_11876,N_13101);
nand U24688 (N_24688,N_11026,N_17829);
and U24689 (N_24689,N_15696,N_15002);
xor U24690 (N_24690,N_13645,N_13278);
xor U24691 (N_24691,N_13487,N_12833);
nand U24692 (N_24692,N_11407,N_10976);
nor U24693 (N_24693,N_18371,N_10560);
or U24694 (N_24694,N_15878,N_12338);
xor U24695 (N_24695,N_18136,N_10713);
or U24696 (N_24696,N_10882,N_15440);
or U24697 (N_24697,N_19207,N_13174);
and U24698 (N_24698,N_11400,N_17162);
xor U24699 (N_24699,N_10516,N_17735);
xnor U24700 (N_24700,N_18771,N_15364);
and U24701 (N_24701,N_14457,N_17659);
nor U24702 (N_24702,N_16815,N_11179);
and U24703 (N_24703,N_11439,N_15423);
or U24704 (N_24704,N_11879,N_12218);
nor U24705 (N_24705,N_12421,N_17467);
or U24706 (N_24706,N_15589,N_15046);
nor U24707 (N_24707,N_12983,N_13472);
or U24708 (N_24708,N_17796,N_11753);
and U24709 (N_24709,N_11363,N_14235);
nand U24710 (N_24710,N_12923,N_16210);
or U24711 (N_24711,N_12135,N_14108);
nand U24712 (N_24712,N_19718,N_19000);
or U24713 (N_24713,N_10202,N_17897);
nand U24714 (N_24714,N_16450,N_15417);
or U24715 (N_24715,N_10151,N_14412);
xnor U24716 (N_24716,N_11734,N_17775);
and U24717 (N_24717,N_18228,N_13260);
or U24718 (N_24718,N_17604,N_13744);
or U24719 (N_24719,N_10779,N_16236);
nor U24720 (N_24720,N_16904,N_16280);
xor U24721 (N_24721,N_18864,N_14507);
and U24722 (N_24722,N_11662,N_13327);
xnor U24723 (N_24723,N_19251,N_13969);
nand U24724 (N_24724,N_18655,N_13659);
nand U24725 (N_24725,N_15188,N_10933);
nand U24726 (N_24726,N_10459,N_11145);
nand U24727 (N_24727,N_13837,N_18293);
xnor U24728 (N_24728,N_12331,N_19151);
xor U24729 (N_24729,N_13512,N_13551);
nand U24730 (N_24730,N_15875,N_19687);
or U24731 (N_24731,N_10376,N_19776);
and U24732 (N_24732,N_10641,N_13415);
and U24733 (N_24733,N_11267,N_11227);
xnor U24734 (N_24734,N_19627,N_12519);
and U24735 (N_24735,N_12323,N_15097);
and U24736 (N_24736,N_14929,N_17592);
nor U24737 (N_24737,N_17692,N_15281);
nand U24738 (N_24738,N_13904,N_15843);
or U24739 (N_24739,N_11214,N_14489);
and U24740 (N_24740,N_18047,N_15627);
nand U24741 (N_24741,N_12241,N_17571);
or U24742 (N_24742,N_14629,N_17940);
xnor U24743 (N_24743,N_17621,N_15570);
and U24744 (N_24744,N_16642,N_19723);
nor U24745 (N_24745,N_15849,N_18548);
nand U24746 (N_24746,N_10589,N_17938);
xor U24747 (N_24747,N_10325,N_12997);
or U24748 (N_24748,N_19217,N_12791);
and U24749 (N_24749,N_14228,N_19686);
xor U24750 (N_24750,N_14905,N_17042);
or U24751 (N_24751,N_12846,N_10790);
and U24752 (N_24752,N_18830,N_11769);
nor U24753 (N_24753,N_18318,N_12621);
or U24754 (N_24754,N_19592,N_19901);
nand U24755 (N_24755,N_18469,N_11786);
nor U24756 (N_24756,N_11624,N_10615);
and U24757 (N_24757,N_14482,N_17824);
nand U24758 (N_24758,N_14838,N_19648);
or U24759 (N_24759,N_10957,N_13660);
nor U24760 (N_24760,N_13284,N_10705);
xor U24761 (N_24761,N_15673,N_12629);
and U24762 (N_24762,N_15489,N_10698);
xor U24763 (N_24763,N_12664,N_13610);
xnor U24764 (N_24764,N_13120,N_18956);
nor U24765 (N_24765,N_15208,N_19177);
nor U24766 (N_24766,N_19882,N_19056);
nand U24767 (N_24767,N_17333,N_13859);
nand U24768 (N_24768,N_14185,N_13306);
xor U24769 (N_24769,N_18692,N_10495);
nor U24770 (N_24770,N_12999,N_13219);
nand U24771 (N_24771,N_17631,N_12370);
xor U24772 (N_24772,N_17636,N_10186);
xnor U24773 (N_24773,N_10833,N_15333);
nor U24774 (N_24774,N_10966,N_16646);
and U24775 (N_24775,N_10928,N_11562);
nor U24776 (N_24776,N_17845,N_14759);
nor U24777 (N_24777,N_19146,N_18084);
nor U24778 (N_24778,N_16846,N_18627);
xnor U24779 (N_24779,N_13042,N_13881);
nand U24780 (N_24780,N_18524,N_14475);
and U24781 (N_24781,N_13170,N_15641);
and U24782 (N_24782,N_14479,N_14440);
or U24783 (N_24783,N_11318,N_11657);
nor U24784 (N_24784,N_16862,N_12150);
or U24785 (N_24785,N_17962,N_15826);
nor U24786 (N_24786,N_18337,N_11553);
or U24787 (N_24787,N_12305,N_14758);
nor U24788 (N_24788,N_19732,N_18602);
and U24789 (N_24789,N_19051,N_14275);
nor U24790 (N_24790,N_13435,N_13495);
nand U24791 (N_24791,N_15918,N_13433);
nor U24792 (N_24792,N_17283,N_12763);
xnor U24793 (N_24793,N_13172,N_18798);
nor U24794 (N_24794,N_18483,N_12914);
nand U24795 (N_24795,N_19910,N_11757);
or U24796 (N_24796,N_13499,N_10582);
nand U24797 (N_24797,N_12733,N_19118);
xnor U24798 (N_24798,N_12752,N_13547);
xor U24799 (N_24799,N_15202,N_12738);
and U24800 (N_24800,N_18516,N_11353);
xor U24801 (N_24801,N_17399,N_11321);
xnor U24802 (N_24802,N_11375,N_19831);
or U24803 (N_24803,N_12045,N_17647);
and U24804 (N_24804,N_15845,N_18298);
nor U24805 (N_24805,N_16065,N_18901);
nand U24806 (N_24806,N_16307,N_14272);
nor U24807 (N_24807,N_13468,N_18218);
nor U24808 (N_24808,N_17731,N_15382);
nand U24809 (N_24809,N_19400,N_11698);
nand U24810 (N_24810,N_13158,N_13784);
or U24811 (N_24811,N_19002,N_15505);
nor U24812 (N_24812,N_19179,N_18434);
nand U24813 (N_24813,N_15774,N_17544);
nor U24814 (N_24814,N_19224,N_17147);
xnor U24815 (N_24815,N_16955,N_14959);
nor U24816 (N_24816,N_17185,N_10662);
nand U24817 (N_24817,N_14889,N_14095);
nand U24818 (N_24818,N_10750,N_10857);
nor U24819 (N_24819,N_13057,N_16205);
and U24820 (N_24820,N_17566,N_17928);
and U24821 (N_24821,N_11806,N_14558);
xor U24822 (N_24822,N_16401,N_14802);
and U24823 (N_24823,N_17914,N_12068);
nor U24824 (N_24824,N_12030,N_12854);
and U24825 (N_24825,N_14633,N_19452);
or U24826 (N_24826,N_12598,N_17186);
nor U24827 (N_24827,N_12427,N_13717);
and U24828 (N_24828,N_14598,N_14826);
or U24829 (N_24829,N_12868,N_15066);
nand U24830 (N_24830,N_16391,N_10213);
or U24831 (N_24831,N_11836,N_14278);
or U24832 (N_24832,N_13755,N_15534);
nand U24833 (N_24833,N_14592,N_15988);
or U24834 (N_24834,N_16150,N_13535);
or U24835 (N_24835,N_15227,N_13149);
and U24836 (N_24836,N_18923,N_14946);
nor U24837 (N_24837,N_11164,N_14481);
xnor U24838 (N_24838,N_10009,N_19140);
xnor U24839 (N_24839,N_15941,N_19936);
nand U24840 (N_24840,N_11383,N_14647);
nand U24841 (N_24841,N_15256,N_11202);
nand U24842 (N_24842,N_14346,N_12302);
xor U24843 (N_24843,N_14222,N_10044);
or U24844 (N_24844,N_12420,N_17687);
or U24845 (N_24845,N_11426,N_15699);
nor U24846 (N_24846,N_12148,N_13871);
and U24847 (N_24847,N_15885,N_19498);
and U24848 (N_24848,N_19705,N_15001);
xor U24849 (N_24849,N_10581,N_12339);
xor U24850 (N_24850,N_14414,N_16703);
and U24851 (N_24851,N_12193,N_13166);
nand U24852 (N_24852,N_10413,N_18895);
nor U24853 (N_24853,N_17178,N_19508);
xor U24854 (N_24854,N_10278,N_18841);
and U24855 (N_24855,N_15969,N_13844);
nor U24856 (N_24856,N_11993,N_11212);
or U24857 (N_24857,N_10852,N_15753);
xnor U24858 (N_24858,N_14692,N_13098);
nand U24859 (N_24859,N_19340,N_13501);
and U24860 (N_24860,N_13944,N_14628);
nand U24861 (N_24861,N_11810,N_15726);
nor U24862 (N_24862,N_12929,N_15787);
nor U24863 (N_24863,N_16000,N_13756);
xnor U24864 (N_24864,N_14496,N_16457);
or U24865 (N_24865,N_15430,N_16784);
or U24866 (N_24866,N_10086,N_13654);
nand U24867 (N_24867,N_12825,N_14861);
nor U24868 (N_24868,N_10412,N_18069);
xor U24869 (N_24869,N_11672,N_19604);
and U24870 (N_24870,N_13029,N_16615);
xor U24871 (N_24871,N_10718,N_17696);
nor U24872 (N_24872,N_18962,N_16793);
nor U24873 (N_24873,N_13991,N_17662);
and U24874 (N_24874,N_14191,N_11525);
and U24875 (N_24875,N_19363,N_10208);
and U24876 (N_24876,N_12313,N_15801);
nand U24877 (N_24877,N_13515,N_15842);
and U24878 (N_24878,N_16744,N_18995);
and U24879 (N_24879,N_13425,N_11073);
and U24880 (N_24880,N_12261,N_11805);
nand U24881 (N_24881,N_10411,N_13602);
and U24882 (N_24882,N_17717,N_11287);
and U24883 (N_24883,N_15163,N_10212);
xor U24884 (N_24884,N_10950,N_19283);
or U24885 (N_24885,N_11578,N_12407);
xnor U24886 (N_24886,N_11718,N_11398);
nor U24887 (N_24887,N_13118,N_16790);
nand U24888 (N_24888,N_15456,N_15532);
and U24889 (N_24889,N_10326,N_14515);
and U24890 (N_24890,N_11640,N_14368);
nand U24891 (N_24891,N_10102,N_15120);
nand U24892 (N_24892,N_17107,N_11962);
xnor U24893 (N_24893,N_17372,N_17003);
or U24894 (N_24894,N_10585,N_12819);
nand U24895 (N_24895,N_14983,N_15394);
nand U24896 (N_24896,N_13518,N_19325);
nand U24897 (N_24897,N_13811,N_10281);
or U24898 (N_24898,N_16381,N_13974);
nor U24899 (N_24899,N_12411,N_17523);
or U24900 (N_24900,N_16112,N_12746);
xnor U24901 (N_24901,N_10299,N_13555);
and U24902 (N_24902,N_11282,N_10660);
or U24903 (N_24903,N_16675,N_17425);
and U24904 (N_24904,N_10431,N_14715);
nor U24905 (N_24905,N_15081,N_18809);
nand U24906 (N_24906,N_12255,N_14456);
or U24907 (N_24907,N_13937,N_16886);
xnor U24908 (N_24908,N_11528,N_13560);
nor U24909 (N_24909,N_15793,N_13462);
or U24910 (N_24910,N_19982,N_13205);
nand U24911 (N_24911,N_19993,N_12701);
nor U24912 (N_24912,N_12108,N_17997);
nor U24913 (N_24913,N_15076,N_12406);
xnor U24914 (N_24914,N_17303,N_19563);
nand U24915 (N_24915,N_12528,N_16647);
nand U24916 (N_24916,N_18215,N_10663);
and U24917 (N_24917,N_17620,N_15933);
and U24918 (N_24918,N_15201,N_12749);
nand U24919 (N_24919,N_11872,N_19929);
nand U24920 (N_24920,N_15819,N_11583);
nand U24921 (N_24921,N_13183,N_12291);
nand U24922 (N_24922,N_13079,N_17034);
nor U24923 (N_24923,N_16439,N_19696);
xnor U24924 (N_24924,N_10148,N_12689);
nor U24925 (N_24925,N_10781,N_13917);
xnor U24926 (N_24926,N_16367,N_19802);
nor U24927 (N_24927,N_15053,N_12591);
nor U24928 (N_24928,N_17923,N_13034);
or U24929 (N_24929,N_10666,N_11236);
or U24930 (N_24930,N_12118,N_12583);
and U24931 (N_24931,N_15614,N_15424);
nand U24932 (N_24932,N_19573,N_13780);
or U24933 (N_24933,N_13829,N_18716);
xnor U24934 (N_24934,N_12727,N_19492);
and U24935 (N_24935,N_13510,N_13770);
xnor U24936 (N_24936,N_16588,N_15040);
and U24937 (N_24937,N_11159,N_10420);
or U24938 (N_24938,N_16218,N_13411);
nor U24939 (N_24939,N_15177,N_12592);
nand U24940 (N_24940,N_19157,N_13549);
nor U24941 (N_24941,N_15222,N_13410);
nor U24942 (N_24942,N_19322,N_13849);
nand U24943 (N_24943,N_10892,N_13114);
xor U24944 (N_24944,N_17630,N_19562);
and U24945 (N_24945,N_14904,N_16111);
nor U24946 (N_24946,N_11942,N_18965);
xor U24947 (N_24947,N_18086,N_19849);
nor U24948 (N_24948,N_11902,N_16892);
and U24949 (N_24949,N_17339,N_12927);
nand U24950 (N_24950,N_10819,N_14446);
nor U24951 (N_24951,N_13454,N_19354);
nor U24952 (N_24952,N_18802,N_17811);
or U24953 (N_24953,N_13058,N_15607);
and U24954 (N_24954,N_19808,N_13782);
and U24955 (N_24955,N_12368,N_14163);
xnor U24956 (N_24956,N_16666,N_11463);
or U24957 (N_24957,N_14343,N_16364);
or U24958 (N_24958,N_15089,N_10545);
xnor U24959 (N_24959,N_19819,N_15080);
nand U24960 (N_24960,N_10997,N_18499);
nor U24961 (N_24961,N_19392,N_15162);
or U24962 (N_24962,N_12786,N_15604);
or U24963 (N_24963,N_12642,N_12682);
or U24964 (N_24964,N_17390,N_17517);
or U24965 (N_24965,N_10601,N_11933);
nand U24966 (N_24966,N_12661,N_18600);
and U24967 (N_24967,N_10849,N_18712);
nand U24968 (N_24968,N_13693,N_13566);
nor U24969 (N_24969,N_12213,N_14590);
and U24970 (N_24970,N_18657,N_17688);
nor U24971 (N_24971,N_16880,N_13145);
and U24972 (N_24972,N_15355,N_16172);
and U24973 (N_24973,N_15125,N_11390);
or U24974 (N_24974,N_12943,N_11045);
or U24975 (N_24975,N_19578,N_11330);
xnor U24976 (N_24976,N_10839,N_13335);
xnor U24977 (N_24977,N_11859,N_12551);
nand U24978 (N_24978,N_12920,N_10919);
nor U24979 (N_24979,N_16138,N_17306);
xnor U24980 (N_24980,N_16721,N_11763);
xnor U24981 (N_24981,N_18767,N_10521);
and U24982 (N_24982,N_18824,N_18529);
nand U24983 (N_24983,N_18079,N_16447);
nor U24984 (N_24984,N_15110,N_13968);
or U24985 (N_24985,N_12044,N_12472);
xnor U24986 (N_24986,N_12552,N_10301);
xor U24987 (N_24987,N_12262,N_11811);
and U24988 (N_24988,N_17310,N_18303);
nor U24989 (N_24989,N_17227,N_12842);
or U24990 (N_24990,N_15442,N_16404);
or U24991 (N_24991,N_15365,N_12641);
or U24992 (N_24992,N_15617,N_13291);
nand U24993 (N_24993,N_18435,N_18020);
nor U24994 (N_24994,N_17836,N_17045);
nor U24995 (N_24995,N_13713,N_12050);
nand U24996 (N_24996,N_14501,N_17049);
nand U24997 (N_24997,N_19716,N_19343);
nand U24998 (N_24998,N_10154,N_10191);
and U24999 (N_24999,N_11629,N_18357);
nor U25000 (N_25000,N_19022,N_18065);
xnor U25001 (N_25001,N_11874,N_17241);
nor U25002 (N_25002,N_15368,N_11766);
and U25003 (N_25003,N_12767,N_13034);
or U25004 (N_25004,N_14025,N_12730);
or U25005 (N_25005,N_17180,N_10149);
and U25006 (N_25006,N_19467,N_14423);
or U25007 (N_25007,N_14988,N_15990);
and U25008 (N_25008,N_16945,N_13104);
nand U25009 (N_25009,N_10920,N_17335);
and U25010 (N_25010,N_16949,N_18464);
xnor U25011 (N_25011,N_10923,N_10471);
or U25012 (N_25012,N_18239,N_17618);
xor U25013 (N_25013,N_13354,N_13103);
nor U25014 (N_25014,N_10036,N_11618);
nand U25015 (N_25015,N_18355,N_17909);
nor U25016 (N_25016,N_14337,N_18233);
nor U25017 (N_25017,N_16590,N_11506);
nand U25018 (N_25018,N_17866,N_14362);
or U25019 (N_25019,N_12403,N_13040);
nand U25020 (N_25020,N_15465,N_19595);
or U25021 (N_25021,N_15419,N_16697);
or U25022 (N_25022,N_10463,N_12924);
or U25023 (N_25023,N_18161,N_16823);
or U25024 (N_25024,N_11276,N_14665);
and U25025 (N_25025,N_18469,N_13779);
nand U25026 (N_25026,N_16276,N_11999);
xnor U25027 (N_25027,N_18292,N_12157);
nor U25028 (N_25028,N_13902,N_17081);
and U25029 (N_25029,N_12994,N_16204);
nor U25030 (N_25030,N_17254,N_19786);
and U25031 (N_25031,N_18305,N_18914);
nor U25032 (N_25032,N_11895,N_16222);
nand U25033 (N_25033,N_19207,N_11849);
xnor U25034 (N_25034,N_18893,N_11367);
and U25035 (N_25035,N_15223,N_16490);
or U25036 (N_25036,N_10997,N_12749);
and U25037 (N_25037,N_12197,N_12906);
or U25038 (N_25038,N_10340,N_13066);
or U25039 (N_25039,N_15843,N_12910);
nor U25040 (N_25040,N_17081,N_14787);
nand U25041 (N_25041,N_12274,N_19875);
nor U25042 (N_25042,N_17659,N_16440);
nor U25043 (N_25043,N_14727,N_18671);
or U25044 (N_25044,N_12488,N_13749);
nor U25045 (N_25045,N_17354,N_12975);
or U25046 (N_25046,N_19289,N_18870);
and U25047 (N_25047,N_15622,N_11265);
xor U25048 (N_25048,N_11118,N_17134);
nand U25049 (N_25049,N_19956,N_16507);
nor U25050 (N_25050,N_17100,N_18641);
and U25051 (N_25051,N_18966,N_14011);
and U25052 (N_25052,N_14785,N_14957);
xnor U25053 (N_25053,N_13427,N_14092);
or U25054 (N_25054,N_14774,N_12032);
and U25055 (N_25055,N_12325,N_14508);
and U25056 (N_25056,N_13102,N_13645);
xor U25057 (N_25057,N_11942,N_11915);
or U25058 (N_25058,N_18607,N_10637);
and U25059 (N_25059,N_18835,N_17590);
or U25060 (N_25060,N_15475,N_19008);
nor U25061 (N_25061,N_16456,N_18594);
and U25062 (N_25062,N_19054,N_18915);
and U25063 (N_25063,N_18303,N_12741);
nand U25064 (N_25064,N_11781,N_19651);
or U25065 (N_25065,N_16195,N_13075);
and U25066 (N_25066,N_15969,N_10983);
or U25067 (N_25067,N_19309,N_15314);
xor U25068 (N_25068,N_15138,N_10760);
nor U25069 (N_25069,N_12055,N_15913);
nor U25070 (N_25070,N_12023,N_11008);
or U25071 (N_25071,N_15140,N_15132);
nor U25072 (N_25072,N_19615,N_17551);
nor U25073 (N_25073,N_13766,N_18147);
and U25074 (N_25074,N_16931,N_15965);
or U25075 (N_25075,N_14603,N_17478);
nor U25076 (N_25076,N_17226,N_11077);
xor U25077 (N_25077,N_15477,N_15027);
and U25078 (N_25078,N_12174,N_10727);
and U25079 (N_25079,N_14401,N_16091);
nor U25080 (N_25080,N_17246,N_18429);
xor U25081 (N_25081,N_12617,N_11326);
or U25082 (N_25082,N_13317,N_10808);
nor U25083 (N_25083,N_11785,N_18727);
xnor U25084 (N_25084,N_18710,N_14579);
and U25085 (N_25085,N_14873,N_12459);
or U25086 (N_25086,N_19969,N_15639);
nand U25087 (N_25087,N_12201,N_18951);
nor U25088 (N_25088,N_10374,N_14990);
nand U25089 (N_25089,N_14817,N_11561);
or U25090 (N_25090,N_18005,N_11947);
and U25091 (N_25091,N_10439,N_15973);
xor U25092 (N_25092,N_17458,N_13841);
xor U25093 (N_25093,N_15388,N_15752);
and U25094 (N_25094,N_18634,N_16358);
nand U25095 (N_25095,N_18582,N_14923);
xnor U25096 (N_25096,N_14323,N_18734);
or U25097 (N_25097,N_12243,N_16410);
nand U25098 (N_25098,N_15552,N_18053);
and U25099 (N_25099,N_14612,N_14854);
xor U25100 (N_25100,N_16223,N_13008);
nor U25101 (N_25101,N_16145,N_13340);
or U25102 (N_25102,N_13569,N_11676);
nor U25103 (N_25103,N_10172,N_15344);
nor U25104 (N_25104,N_12898,N_12423);
and U25105 (N_25105,N_14522,N_11960);
xnor U25106 (N_25106,N_10096,N_14558);
xor U25107 (N_25107,N_16257,N_10913);
xor U25108 (N_25108,N_16884,N_17266);
xor U25109 (N_25109,N_19690,N_11284);
xor U25110 (N_25110,N_19696,N_19178);
nor U25111 (N_25111,N_18038,N_19769);
and U25112 (N_25112,N_19084,N_10517);
nand U25113 (N_25113,N_19463,N_14766);
nor U25114 (N_25114,N_11246,N_10027);
xor U25115 (N_25115,N_13150,N_19325);
nor U25116 (N_25116,N_16851,N_15525);
and U25117 (N_25117,N_12875,N_11297);
nand U25118 (N_25118,N_18186,N_17542);
nand U25119 (N_25119,N_19547,N_18145);
and U25120 (N_25120,N_11595,N_16074);
nand U25121 (N_25121,N_11644,N_17727);
nor U25122 (N_25122,N_19174,N_10574);
nor U25123 (N_25123,N_18291,N_12394);
nor U25124 (N_25124,N_15422,N_11723);
or U25125 (N_25125,N_16974,N_19972);
and U25126 (N_25126,N_15735,N_18243);
xor U25127 (N_25127,N_19389,N_18705);
xor U25128 (N_25128,N_15103,N_18883);
and U25129 (N_25129,N_14385,N_15203);
and U25130 (N_25130,N_18943,N_16170);
or U25131 (N_25131,N_14296,N_16088);
and U25132 (N_25132,N_16748,N_10919);
and U25133 (N_25133,N_19354,N_10445);
xnor U25134 (N_25134,N_11746,N_10876);
xnor U25135 (N_25135,N_11584,N_11653);
xnor U25136 (N_25136,N_18826,N_10208);
xor U25137 (N_25137,N_11874,N_10544);
or U25138 (N_25138,N_19403,N_18350);
nand U25139 (N_25139,N_14974,N_11686);
nor U25140 (N_25140,N_14093,N_10305);
nand U25141 (N_25141,N_19092,N_19523);
and U25142 (N_25142,N_11720,N_18357);
and U25143 (N_25143,N_19779,N_18480);
and U25144 (N_25144,N_15450,N_16255);
nor U25145 (N_25145,N_16279,N_13830);
nor U25146 (N_25146,N_10620,N_10680);
nor U25147 (N_25147,N_13618,N_15201);
or U25148 (N_25148,N_17812,N_11291);
nor U25149 (N_25149,N_13857,N_14679);
xnor U25150 (N_25150,N_11426,N_15840);
nand U25151 (N_25151,N_15821,N_17157);
nor U25152 (N_25152,N_10063,N_19915);
nor U25153 (N_25153,N_17177,N_11789);
nor U25154 (N_25154,N_15028,N_16022);
nor U25155 (N_25155,N_14841,N_10823);
nand U25156 (N_25156,N_10716,N_14951);
or U25157 (N_25157,N_19437,N_17402);
nand U25158 (N_25158,N_14403,N_13523);
and U25159 (N_25159,N_12843,N_15276);
nor U25160 (N_25160,N_15589,N_10319);
or U25161 (N_25161,N_15512,N_12969);
xor U25162 (N_25162,N_18318,N_13077);
nand U25163 (N_25163,N_19483,N_15372);
or U25164 (N_25164,N_11970,N_15980);
nand U25165 (N_25165,N_18542,N_19083);
xor U25166 (N_25166,N_15853,N_19046);
nor U25167 (N_25167,N_14881,N_19548);
nand U25168 (N_25168,N_18858,N_16536);
and U25169 (N_25169,N_13626,N_19952);
xor U25170 (N_25170,N_16658,N_16273);
and U25171 (N_25171,N_13423,N_15759);
and U25172 (N_25172,N_17777,N_18554);
or U25173 (N_25173,N_11211,N_10999);
and U25174 (N_25174,N_12915,N_17021);
nand U25175 (N_25175,N_12005,N_15372);
xor U25176 (N_25176,N_17708,N_14757);
nand U25177 (N_25177,N_10804,N_12557);
nand U25178 (N_25178,N_18662,N_19879);
xor U25179 (N_25179,N_18344,N_18881);
xor U25180 (N_25180,N_11265,N_17885);
xor U25181 (N_25181,N_10921,N_16374);
or U25182 (N_25182,N_13775,N_12629);
nor U25183 (N_25183,N_16325,N_11675);
and U25184 (N_25184,N_18600,N_15866);
nand U25185 (N_25185,N_15437,N_19593);
nand U25186 (N_25186,N_16116,N_16803);
or U25187 (N_25187,N_15510,N_12631);
nor U25188 (N_25188,N_10348,N_17579);
or U25189 (N_25189,N_18651,N_14475);
or U25190 (N_25190,N_10124,N_16266);
nand U25191 (N_25191,N_10749,N_10858);
nor U25192 (N_25192,N_11213,N_16466);
or U25193 (N_25193,N_10292,N_18799);
and U25194 (N_25194,N_16949,N_14436);
nand U25195 (N_25195,N_17652,N_17006);
xor U25196 (N_25196,N_18530,N_11285);
nand U25197 (N_25197,N_14113,N_16360);
nand U25198 (N_25198,N_11638,N_14748);
or U25199 (N_25199,N_13064,N_12489);
nor U25200 (N_25200,N_11528,N_11925);
or U25201 (N_25201,N_19667,N_12561);
nor U25202 (N_25202,N_18042,N_11380);
xor U25203 (N_25203,N_10237,N_13608);
xor U25204 (N_25204,N_12583,N_14696);
nor U25205 (N_25205,N_14584,N_12575);
and U25206 (N_25206,N_10565,N_18098);
nor U25207 (N_25207,N_10387,N_19440);
or U25208 (N_25208,N_14537,N_12848);
or U25209 (N_25209,N_10272,N_16862);
nor U25210 (N_25210,N_16602,N_11015);
or U25211 (N_25211,N_12445,N_13338);
xor U25212 (N_25212,N_15543,N_18304);
nand U25213 (N_25213,N_14639,N_14743);
xnor U25214 (N_25214,N_18132,N_14957);
or U25215 (N_25215,N_17753,N_12209);
xor U25216 (N_25216,N_11104,N_12943);
or U25217 (N_25217,N_19109,N_18505);
or U25218 (N_25218,N_14674,N_16840);
and U25219 (N_25219,N_10363,N_15111);
nand U25220 (N_25220,N_10827,N_13951);
and U25221 (N_25221,N_11831,N_14654);
nand U25222 (N_25222,N_18325,N_10661);
or U25223 (N_25223,N_11462,N_10445);
xor U25224 (N_25224,N_10009,N_19083);
or U25225 (N_25225,N_19734,N_16863);
nor U25226 (N_25226,N_15643,N_18152);
and U25227 (N_25227,N_18024,N_14173);
and U25228 (N_25228,N_10599,N_16796);
and U25229 (N_25229,N_14641,N_18927);
or U25230 (N_25230,N_17277,N_17416);
and U25231 (N_25231,N_16204,N_16168);
and U25232 (N_25232,N_12816,N_16610);
nor U25233 (N_25233,N_18721,N_17719);
xnor U25234 (N_25234,N_10515,N_17491);
nand U25235 (N_25235,N_11969,N_12851);
or U25236 (N_25236,N_10408,N_18071);
xnor U25237 (N_25237,N_14644,N_16417);
nor U25238 (N_25238,N_16966,N_14532);
or U25239 (N_25239,N_14017,N_15283);
nor U25240 (N_25240,N_16106,N_15100);
nor U25241 (N_25241,N_19563,N_12464);
xor U25242 (N_25242,N_16916,N_11847);
nand U25243 (N_25243,N_12621,N_14232);
xnor U25244 (N_25244,N_11573,N_19791);
or U25245 (N_25245,N_15235,N_17667);
and U25246 (N_25246,N_18137,N_17545);
or U25247 (N_25247,N_18142,N_14267);
and U25248 (N_25248,N_15746,N_16178);
and U25249 (N_25249,N_13350,N_11228);
and U25250 (N_25250,N_11145,N_17252);
xor U25251 (N_25251,N_18052,N_18664);
nand U25252 (N_25252,N_10078,N_16701);
and U25253 (N_25253,N_15909,N_10465);
xnor U25254 (N_25254,N_11451,N_16126);
xor U25255 (N_25255,N_16201,N_12152);
nand U25256 (N_25256,N_13170,N_18505);
or U25257 (N_25257,N_16885,N_16272);
xor U25258 (N_25258,N_14190,N_11458);
xnor U25259 (N_25259,N_12443,N_14745);
nor U25260 (N_25260,N_16116,N_19417);
xnor U25261 (N_25261,N_11147,N_14244);
or U25262 (N_25262,N_14954,N_14195);
and U25263 (N_25263,N_15470,N_14352);
xor U25264 (N_25264,N_12700,N_13571);
nand U25265 (N_25265,N_14929,N_12320);
nand U25266 (N_25266,N_11741,N_11165);
or U25267 (N_25267,N_18061,N_16380);
xnor U25268 (N_25268,N_18330,N_13923);
or U25269 (N_25269,N_10616,N_17916);
nor U25270 (N_25270,N_15396,N_15783);
xor U25271 (N_25271,N_14879,N_19177);
or U25272 (N_25272,N_10580,N_14386);
and U25273 (N_25273,N_18150,N_15705);
nor U25274 (N_25274,N_17289,N_10877);
or U25275 (N_25275,N_12412,N_15587);
or U25276 (N_25276,N_17098,N_11394);
nand U25277 (N_25277,N_19769,N_13082);
xnor U25278 (N_25278,N_14830,N_11163);
nand U25279 (N_25279,N_11105,N_19305);
and U25280 (N_25280,N_16871,N_19747);
or U25281 (N_25281,N_16917,N_16247);
xor U25282 (N_25282,N_13069,N_14893);
xnor U25283 (N_25283,N_14197,N_15352);
nand U25284 (N_25284,N_18954,N_16041);
nor U25285 (N_25285,N_16123,N_16184);
nand U25286 (N_25286,N_19872,N_17856);
and U25287 (N_25287,N_10091,N_10187);
nor U25288 (N_25288,N_17185,N_17212);
xor U25289 (N_25289,N_11585,N_15071);
or U25290 (N_25290,N_16073,N_16042);
or U25291 (N_25291,N_16037,N_12532);
and U25292 (N_25292,N_17209,N_14679);
nor U25293 (N_25293,N_10576,N_19714);
and U25294 (N_25294,N_17468,N_14758);
nor U25295 (N_25295,N_11115,N_12597);
or U25296 (N_25296,N_16956,N_18420);
or U25297 (N_25297,N_10702,N_15750);
xor U25298 (N_25298,N_13439,N_19488);
and U25299 (N_25299,N_16585,N_16956);
and U25300 (N_25300,N_18284,N_14367);
nand U25301 (N_25301,N_17343,N_15774);
or U25302 (N_25302,N_17509,N_15613);
and U25303 (N_25303,N_17466,N_10852);
and U25304 (N_25304,N_13134,N_12832);
xnor U25305 (N_25305,N_11104,N_10286);
nor U25306 (N_25306,N_12938,N_18732);
nand U25307 (N_25307,N_16390,N_11961);
and U25308 (N_25308,N_13425,N_14479);
and U25309 (N_25309,N_11515,N_12725);
nor U25310 (N_25310,N_18430,N_14109);
nand U25311 (N_25311,N_14116,N_10501);
and U25312 (N_25312,N_15292,N_13757);
nor U25313 (N_25313,N_14002,N_11770);
nor U25314 (N_25314,N_16713,N_16002);
or U25315 (N_25315,N_18860,N_14852);
nand U25316 (N_25316,N_12103,N_17755);
or U25317 (N_25317,N_11935,N_12301);
and U25318 (N_25318,N_12035,N_11224);
or U25319 (N_25319,N_15101,N_14860);
xnor U25320 (N_25320,N_17367,N_15973);
nand U25321 (N_25321,N_15014,N_16957);
nand U25322 (N_25322,N_10322,N_13752);
nand U25323 (N_25323,N_18122,N_19082);
xnor U25324 (N_25324,N_17395,N_17755);
or U25325 (N_25325,N_12016,N_19047);
or U25326 (N_25326,N_11934,N_10298);
and U25327 (N_25327,N_17380,N_14081);
and U25328 (N_25328,N_13452,N_16339);
xnor U25329 (N_25329,N_13429,N_16283);
xnor U25330 (N_25330,N_19384,N_14681);
nor U25331 (N_25331,N_14081,N_18017);
and U25332 (N_25332,N_17736,N_17514);
xnor U25333 (N_25333,N_19090,N_15683);
nor U25334 (N_25334,N_18204,N_14806);
nor U25335 (N_25335,N_19265,N_15652);
and U25336 (N_25336,N_17776,N_10590);
and U25337 (N_25337,N_17174,N_11513);
xor U25338 (N_25338,N_15147,N_13980);
nand U25339 (N_25339,N_14519,N_13995);
nand U25340 (N_25340,N_15748,N_19604);
or U25341 (N_25341,N_15758,N_13032);
or U25342 (N_25342,N_17011,N_19617);
xnor U25343 (N_25343,N_18187,N_16869);
and U25344 (N_25344,N_11499,N_10771);
and U25345 (N_25345,N_17894,N_17423);
and U25346 (N_25346,N_13806,N_10282);
or U25347 (N_25347,N_16348,N_10521);
nand U25348 (N_25348,N_11221,N_12513);
nand U25349 (N_25349,N_17555,N_19450);
nor U25350 (N_25350,N_16972,N_11005);
or U25351 (N_25351,N_12671,N_13490);
nor U25352 (N_25352,N_17605,N_19875);
xnor U25353 (N_25353,N_18478,N_19039);
nor U25354 (N_25354,N_14735,N_16456);
and U25355 (N_25355,N_17248,N_14393);
xor U25356 (N_25356,N_18822,N_14231);
xnor U25357 (N_25357,N_15405,N_13686);
nand U25358 (N_25358,N_12903,N_15738);
xor U25359 (N_25359,N_18905,N_12072);
and U25360 (N_25360,N_18512,N_10845);
or U25361 (N_25361,N_12188,N_10278);
or U25362 (N_25362,N_15632,N_18629);
xor U25363 (N_25363,N_18148,N_13102);
nor U25364 (N_25364,N_17903,N_16583);
xor U25365 (N_25365,N_11239,N_19239);
nand U25366 (N_25366,N_17905,N_16739);
and U25367 (N_25367,N_13326,N_10379);
xnor U25368 (N_25368,N_14848,N_12906);
and U25369 (N_25369,N_10758,N_11958);
and U25370 (N_25370,N_14070,N_14687);
xnor U25371 (N_25371,N_10159,N_17503);
or U25372 (N_25372,N_10244,N_16383);
nand U25373 (N_25373,N_19892,N_16899);
nor U25374 (N_25374,N_10394,N_19631);
nor U25375 (N_25375,N_19972,N_12858);
and U25376 (N_25376,N_19218,N_18914);
xnor U25377 (N_25377,N_15676,N_10821);
or U25378 (N_25378,N_17541,N_15436);
or U25379 (N_25379,N_16690,N_10733);
or U25380 (N_25380,N_17531,N_16268);
nand U25381 (N_25381,N_15746,N_18342);
nor U25382 (N_25382,N_18678,N_14528);
and U25383 (N_25383,N_19609,N_11618);
and U25384 (N_25384,N_17664,N_14931);
nand U25385 (N_25385,N_15016,N_19132);
nand U25386 (N_25386,N_17754,N_12060);
xnor U25387 (N_25387,N_19279,N_16011);
nand U25388 (N_25388,N_12064,N_19273);
and U25389 (N_25389,N_11360,N_10941);
nand U25390 (N_25390,N_14587,N_15730);
or U25391 (N_25391,N_19431,N_11015);
xor U25392 (N_25392,N_12188,N_14971);
and U25393 (N_25393,N_11513,N_13555);
and U25394 (N_25394,N_12374,N_10864);
xnor U25395 (N_25395,N_10357,N_12475);
and U25396 (N_25396,N_10980,N_10440);
nand U25397 (N_25397,N_18320,N_16044);
or U25398 (N_25398,N_18837,N_13095);
or U25399 (N_25399,N_19785,N_17415);
nor U25400 (N_25400,N_16509,N_12367);
nand U25401 (N_25401,N_17131,N_19258);
nor U25402 (N_25402,N_16737,N_14255);
and U25403 (N_25403,N_18077,N_16996);
nand U25404 (N_25404,N_16870,N_11515);
nor U25405 (N_25405,N_10932,N_19058);
and U25406 (N_25406,N_17753,N_11674);
or U25407 (N_25407,N_16327,N_14796);
and U25408 (N_25408,N_10492,N_19394);
nor U25409 (N_25409,N_15182,N_14012);
nand U25410 (N_25410,N_14663,N_16823);
nand U25411 (N_25411,N_10776,N_11764);
nor U25412 (N_25412,N_12303,N_16648);
nor U25413 (N_25413,N_12660,N_16025);
nand U25414 (N_25414,N_17912,N_15207);
nand U25415 (N_25415,N_17983,N_12222);
xor U25416 (N_25416,N_12665,N_18996);
nor U25417 (N_25417,N_16638,N_13662);
nand U25418 (N_25418,N_13447,N_12531);
nand U25419 (N_25419,N_12414,N_11888);
nor U25420 (N_25420,N_19799,N_14071);
or U25421 (N_25421,N_17617,N_14188);
nand U25422 (N_25422,N_18338,N_11000);
nand U25423 (N_25423,N_12221,N_16801);
or U25424 (N_25424,N_10903,N_16208);
nor U25425 (N_25425,N_16577,N_18241);
xor U25426 (N_25426,N_17369,N_17088);
nand U25427 (N_25427,N_17655,N_12799);
and U25428 (N_25428,N_15662,N_15305);
or U25429 (N_25429,N_12223,N_17069);
nand U25430 (N_25430,N_12017,N_13672);
or U25431 (N_25431,N_16207,N_11333);
and U25432 (N_25432,N_19014,N_16949);
nand U25433 (N_25433,N_19863,N_16676);
and U25434 (N_25434,N_12911,N_17223);
and U25435 (N_25435,N_19516,N_17616);
and U25436 (N_25436,N_12575,N_10638);
nor U25437 (N_25437,N_14463,N_16968);
nor U25438 (N_25438,N_19547,N_13824);
or U25439 (N_25439,N_12156,N_15961);
nand U25440 (N_25440,N_12698,N_18953);
nor U25441 (N_25441,N_10299,N_11368);
or U25442 (N_25442,N_13805,N_10804);
nor U25443 (N_25443,N_13295,N_14018);
nand U25444 (N_25444,N_15833,N_11808);
and U25445 (N_25445,N_14494,N_13897);
or U25446 (N_25446,N_18958,N_13628);
xnor U25447 (N_25447,N_17679,N_19617);
xor U25448 (N_25448,N_13832,N_17770);
nand U25449 (N_25449,N_10313,N_12981);
or U25450 (N_25450,N_18969,N_15319);
xnor U25451 (N_25451,N_16866,N_19902);
nor U25452 (N_25452,N_12250,N_16509);
or U25453 (N_25453,N_14303,N_15470);
nand U25454 (N_25454,N_18735,N_15184);
nor U25455 (N_25455,N_16414,N_19060);
xnor U25456 (N_25456,N_19706,N_14400);
nor U25457 (N_25457,N_15358,N_15197);
or U25458 (N_25458,N_13206,N_13002);
and U25459 (N_25459,N_17103,N_12102);
xor U25460 (N_25460,N_11220,N_15208);
or U25461 (N_25461,N_13630,N_19110);
xor U25462 (N_25462,N_16350,N_18785);
or U25463 (N_25463,N_18195,N_11278);
or U25464 (N_25464,N_11453,N_17862);
and U25465 (N_25465,N_15300,N_11621);
nand U25466 (N_25466,N_11247,N_10885);
xnor U25467 (N_25467,N_15870,N_11722);
and U25468 (N_25468,N_16577,N_10524);
nand U25469 (N_25469,N_10325,N_16736);
nor U25470 (N_25470,N_10109,N_13819);
or U25471 (N_25471,N_16166,N_12682);
and U25472 (N_25472,N_10669,N_14593);
xnor U25473 (N_25473,N_15207,N_13673);
nor U25474 (N_25474,N_17159,N_14721);
and U25475 (N_25475,N_14802,N_15350);
nand U25476 (N_25476,N_13806,N_16957);
and U25477 (N_25477,N_16471,N_15923);
and U25478 (N_25478,N_15827,N_16401);
nor U25479 (N_25479,N_16285,N_10943);
and U25480 (N_25480,N_10220,N_18849);
nor U25481 (N_25481,N_17959,N_18693);
xor U25482 (N_25482,N_11844,N_16881);
or U25483 (N_25483,N_14009,N_14431);
xnor U25484 (N_25484,N_11826,N_14112);
nor U25485 (N_25485,N_16823,N_11533);
nand U25486 (N_25486,N_11478,N_15251);
xnor U25487 (N_25487,N_12477,N_16357);
and U25488 (N_25488,N_18966,N_14345);
xnor U25489 (N_25489,N_14383,N_18504);
nor U25490 (N_25490,N_11251,N_16537);
or U25491 (N_25491,N_15489,N_16946);
and U25492 (N_25492,N_16725,N_14117);
or U25493 (N_25493,N_15822,N_18600);
xnor U25494 (N_25494,N_11861,N_15693);
and U25495 (N_25495,N_11387,N_13939);
nor U25496 (N_25496,N_14903,N_19106);
nor U25497 (N_25497,N_13226,N_15057);
nand U25498 (N_25498,N_17167,N_13514);
xnor U25499 (N_25499,N_14923,N_16829);
xnor U25500 (N_25500,N_14274,N_11862);
nand U25501 (N_25501,N_18054,N_18943);
or U25502 (N_25502,N_16387,N_12412);
xnor U25503 (N_25503,N_17844,N_16734);
or U25504 (N_25504,N_17913,N_13437);
nor U25505 (N_25505,N_15272,N_17169);
and U25506 (N_25506,N_19877,N_14367);
xnor U25507 (N_25507,N_11195,N_17665);
xnor U25508 (N_25508,N_11365,N_12534);
nor U25509 (N_25509,N_16959,N_10826);
xor U25510 (N_25510,N_10464,N_17517);
or U25511 (N_25511,N_11070,N_15015);
or U25512 (N_25512,N_19405,N_16154);
and U25513 (N_25513,N_15342,N_16532);
xor U25514 (N_25514,N_16616,N_12593);
nand U25515 (N_25515,N_12369,N_17105);
nor U25516 (N_25516,N_11740,N_15901);
xor U25517 (N_25517,N_10458,N_14336);
and U25518 (N_25518,N_10916,N_19038);
and U25519 (N_25519,N_15494,N_13905);
nor U25520 (N_25520,N_13459,N_13753);
xnor U25521 (N_25521,N_15217,N_17985);
nand U25522 (N_25522,N_11626,N_14198);
or U25523 (N_25523,N_11635,N_13531);
or U25524 (N_25524,N_14696,N_12273);
or U25525 (N_25525,N_18884,N_15007);
or U25526 (N_25526,N_10994,N_12588);
nor U25527 (N_25527,N_15355,N_19039);
and U25528 (N_25528,N_11578,N_16944);
and U25529 (N_25529,N_12649,N_15448);
nand U25530 (N_25530,N_14093,N_15973);
nand U25531 (N_25531,N_18387,N_19483);
nor U25532 (N_25532,N_10175,N_10370);
nor U25533 (N_25533,N_10090,N_15779);
and U25534 (N_25534,N_19497,N_10759);
nor U25535 (N_25535,N_15387,N_11398);
nor U25536 (N_25536,N_13138,N_12661);
xnor U25537 (N_25537,N_14289,N_14108);
nand U25538 (N_25538,N_12909,N_18915);
or U25539 (N_25539,N_13024,N_18801);
or U25540 (N_25540,N_11223,N_17594);
or U25541 (N_25541,N_18937,N_17921);
or U25542 (N_25542,N_15852,N_18465);
and U25543 (N_25543,N_13399,N_12871);
and U25544 (N_25544,N_11082,N_14846);
xor U25545 (N_25545,N_14482,N_11776);
nand U25546 (N_25546,N_11536,N_10687);
and U25547 (N_25547,N_16823,N_11231);
nor U25548 (N_25548,N_19807,N_12605);
or U25549 (N_25549,N_14115,N_10576);
and U25550 (N_25550,N_14915,N_15985);
nand U25551 (N_25551,N_11791,N_16900);
nand U25552 (N_25552,N_15527,N_13006);
nor U25553 (N_25553,N_12145,N_13054);
and U25554 (N_25554,N_11273,N_15943);
or U25555 (N_25555,N_17652,N_16729);
nand U25556 (N_25556,N_13316,N_14147);
nor U25557 (N_25557,N_13473,N_10083);
and U25558 (N_25558,N_17019,N_11803);
or U25559 (N_25559,N_10262,N_12916);
and U25560 (N_25560,N_19200,N_19824);
and U25561 (N_25561,N_16704,N_10893);
and U25562 (N_25562,N_19435,N_13022);
nand U25563 (N_25563,N_10383,N_14922);
xor U25564 (N_25564,N_13759,N_13023);
xor U25565 (N_25565,N_19882,N_17853);
xor U25566 (N_25566,N_17983,N_19041);
and U25567 (N_25567,N_12040,N_15866);
xor U25568 (N_25568,N_17321,N_12945);
nor U25569 (N_25569,N_11292,N_17336);
or U25570 (N_25570,N_15676,N_18817);
nor U25571 (N_25571,N_10390,N_10745);
and U25572 (N_25572,N_18946,N_15596);
nor U25573 (N_25573,N_18928,N_14777);
xor U25574 (N_25574,N_15764,N_19995);
xor U25575 (N_25575,N_17178,N_16618);
or U25576 (N_25576,N_15031,N_19625);
or U25577 (N_25577,N_13579,N_18487);
nor U25578 (N_25578,N_16266,N_17840);
nand U25579 (N_25579,N_18010,N_12992);
nand U25580 (N_25580,N_18748,N_17547);
nor U25581 (N_25581,N_19002,N_15347);
xnor U25582 (N_25582,N_14437,N_15703);
xnor U25583 (N_25583,N_12664,N_12424);
or U25584 (N_25584,N_13395,N_11399);
xnor U25585 (N_25585,N_14666,N_12593);
and U25586 (N_25586,N_13323,N_14771);
or U25587 (N_25587,N_14451,N_11342);
nor U25588 (N_25588,N_11895,N_11495);
xnor U25589 (N_25589,N_12748,N_17778);
nor U25590 (N_25590,N_19765,N_14316);
nor U25591 (N_25591,N_10424,N_17156);
nand U25592 (N_25592,N_11355,N_16166);
and U25593 (N_25593,N_10156,N_11038);
and U25594 (N_25594,N_17621,N_11134);
or U25595 (N_25595,N_15065,N_17352);
xnor U25596 (N_25596,N_12412,N_10934);
xnor U25597 (N_25597,N_15573,N_11418);
and U25598 (N_25598,N_18867,N_16855);
xnor U25599 (N_25599,N_15168,N_18051);
nor U25600 (N_25600,N_17158,N_15320);
xnor U25601 (N_25601,N_19946,N_13416);
and U25602 (N_25602,N_13084,N_12507);
nand U25603 (N_25603,N_15275,N_17664);
nor U25604 (N_25604,N_14262,N_10554);
nand U25605 (N_25605,N_15373,N_16418);
nand U25606 (N_25606,N_16408,N_12097);
nand U25607 (N_25607,N_18354,N_19039);
or U25608 (N_25608,N_14559,N_10149);
xnor U25609 (N_25609,N_18971,N_17395);
xor U25610 (N_25610,N_11711,N_14332);
nand U25611 (N_25611,N_19660,N_15675);
and U25612 (N_25612,N_13322,N_17988);
or U25613 (N_25613,N_11877,N_17837);
nand U25614 (N_25614,N_12108,N_13059);
nor U25615 (N_25615,N_19176,N_17299);
or U25616 (N_25616,N_19859,N_16653);
nor U25617 (N_25617,N_16211,N_11471);
nor U25618 (N_25618,N_11335,N_14405);
nand U25619 (N_25619,N_17835,N_12399);
xor U25620 (N_25620,N_13259,N_10456);
and U25621 (N_25621,N_17291,N_13257);
and U25622 (N_25622,N_13042,N_14344);
and U25623 (N_25623,N_12756,N_10865);
nand U25624 (N_25624,N_19782,N_16218);
nor U25625 (N_25625,N_18733,N_10096);
nor U25626 (N_25626,N_16898,N_14280);
nor U25627 (N_25627,N_18387,N_19901);
nor U25628 (N_25628,N_18811,N_12933);
nor U25629 (N_25629,N_17805,N_16730);
or U25630 (N_25630,N_17907,N_11202);
nand U25631 (N_25631,N_13787,N_15781);
nor U25632 (N_25632,N_11682,N_10386);
xor U25633 (N_25633,N_17599,N_13180);
nor U25634 (N_25634,N_16949,N_18642);
or U25635 (N_25635,N_16487,N_19429);
nand U25636 (N_25636,N_18532,N_10877);
nor U25637 (N_25637,N_18472,N_18817);
and U25638 (N_25638,N_10101,N_11278);
xnor U25639 (N_25639,N_16805,N_11338);
and U25640 (N_25640,N_13830,N_12738);
and U25641 (N_25641,N_15003,N_18123);
nor U25642 (N_25642,N_12358,N_14151);
nand U25643 (N_25643,N_10603,N_13227);
or U25644 (N_25644,N_10406,N_18120);
xor U25645 (N_25645,N_10697,N_11926);
xnor U25646 (N_25646,N_16121,N_14493);
xnor U25647 (N_25647,N_17221,N_14031);
nand U25648 (N_25648,N_16499,N_13836);
and U25649 (N_25649,N_18895,N_18317);
nor U25650 (N_25650,N_10295,N_18036);
and U25651 (N_25651,N_12357,N_11979);
nand U25652 (N_25652,N_10997,N_10750);
nand U25653 (N_25653,N_15964,N_16660);
and U25654 (N_25654,N_15972,N_16613);
nand U25655 (N_25655,N_13453,N_18284);
and U25656 (N_25656,N_19072,N_16705);
or U25657 (N_25657,N_13798,N_13453);
and U25658 (N_25658,N_11717,N_15323);
nor U25659 (N_25659,N_14567,N_11187);
and U25660 (N_25660,N_14202,N_16834);
or U25661 (N_25661,N_12722,N_19851);
or U25662 (N_25662,N_19185,N_11605);
xnor U25663 (N_25663,N_16469,N_11191);
nand U25664 (N_25664,N_14501,N_19519);
and U25665 (N_25665,N_12663,N_15481);
xor U25666 (N_25666,N_10847,N_16259);
or U25667 (N_25667,N_16173,N_19583);
or U25668 (N_25668,N_15519,N_11539);
nand U25669 (N_25669,N_10007,N_17073);
or U25670 (N_25670,N_17411,N_12965);
nor U25671 (N_25671,N_16992,N_15280);
nor U25672 (N_25672,N_17581,N_14084);
and U25673 (N_25673,N_15997,N_18476);
and U25674 (N_25674,N_19613,N_12060);
and U25675 (N_25675,N_19988,N_19793);
or U25676 (N_25676,N_15823,N_15278);
nand U25677 (N_25677,N_11713,N_10686);
nand U25678 (N_25678,N_14603,N_17030);
nor U25679 (N_25679,N_16312,N_13369);
nor U25680 (N_25680,N_10103,N_19615);
nor U25681 (N_25681,N_13178,N_11348);
nand U25682 (N_25682,N_11007,N_12015);
and U25683 (N_25683,N_15302,N_17712);
and U25684 (N_25684,N_18419,N_14346);
or U25685 (N_25685,N_15331,N_13202);
and U25686 (N_25686,N_16967,N_11651);
and U25687 (N_25687,N_14720,N_10395);
nor U25688 (N_25688,N_10061,N_14284);
and U25689 (N_25689,N_11829,N_10953);
nand U25690 (N_25690,N_15705,N_16513);
nand U25691 (N_25691,N_19521,N_11930);
xnor U25692 (N_25692,N_11441,N_10376);
nand U25693 (N_25693,N_19533,N_12586);
or U25694 (N_25694,N_18287,N_18101);
nor U25695 (N_25695,N_16950,N_10415);
nor U25696 (N_25696,N_17167,N_13546);
and U25697 (N_25697,N_16183,N_15907);
xnor U25698 (N_25698,N_15381,N_12778);
nor U25699 (N_25699,N_19776,N_16772);
or U25700 (N_25700,N_12620,N_19493);
nor U25701 (N_25701,N_12217,N_19466);
nand U25702 (N_25702,N_19934,N_15961);
nand U25703 (N_25703,N_16332,N_18449);
nand U25704 (N_25704,N_18901,N_14801);
nand U25705 (N_25705,N_13091,N_19327);
nand U25706 (N_25706,N_12974,N_11922);
or U25707 (N_25707,N_18750,N_15464);
nor U25708 (N_25708,N_14702,N_10983);
and U25709 (N_25709,N_17327,N_13527);
and U25710 (N_25710,N_16763,N_16643);
and U25711 (N_25711,N_10689,N_19614);
and U25712 (N_25712,N_13964,N_16696);
and U25713 (N_25713,N_16941,N_16674);
xnor U25714 (N_25714,N_10616,N_15239);
nor U25715 (N_25715,N_17933,N_17783);
and U25716 (N_25716,N_19018,N_12158);
or U25717 (N_25717,N_16010,N_14338);
xnor U25718 (N_25718,N_11317,N_11780);
xor U25719 (N_25719,N_16877,N_13712);
or U25720 (N_25720,N_14001,N_14636);
or U25721 (N_25721,N_17083,N_18691);
nor U25722 (N_25722,N_19748,N_15275);
and U25723 (N_25723,N_19240,N_11819);
or U25724 (N_25724,N_15696,N_17848);
and U25725 (N_25725,N_13141,N_15732);
or U25726 (N_25726,N_19931,N_14184);
nand U25727 (N_25727,N_14300,N_12120);
nand U25728 (N_25728,N_13464,N_13008);
nand U25729 (N_25729,N_16756,N_13205);
nor U25730 (N_25730,N_15227,N_16150);
and U25731 (N_25731,N_10615,N_14136);
xor U25732 (N_25732,N_12857,N_17377);
and U25733 (N_25733,N_16065,N_19833);
or U25734 (N_25734,N_14415,N_18230);
and U25735 (N_25735,N_12150,N_13710);
or U25736 (N_25736,N_10739,N_11722);
and U25737 (N_25737,N_14457,N_13885);
nor U25738 (N_25738,N_14521,N_13040);
nor U25739 (N_25739,N_16632,N_13563);
nand U25740 (N_25740,N_11699,N_19591);
nand U25741 (N_25741,N_14329,N_10256);
xnor U25742 (N_25742,N_19278,N_18608);
xor U25743 (N_25743,N_11549,N_11846);
or U25744 (N_25744,N_11108,N_19214);
nor U25745 (N_25745,N_16304,N_19634);
and U25746 (N_25746,N_14844,N_16344);
nand U25747 (N_25747,N_10215,N_19781);
or U25748 (N_25748,N_19615,N_14144);
nor U25749 (N_25749,N_13647,N_14997);
nand U25750 (N_25750,N_15523,N_15412);
nand U25751 (N_25751,N_13795,N_13939);
xnor U25752 (N_25752,N_13109,N_16090);
and U25753 (N_25753,N_12459,N_16627);
nor U25754 (N_25754,N_12568,N_10957);
or U25755 (N_25755,N_16561,N_10572);
nor U25756 (N_25756,N_19024,N_10352);
and U25757 (N_25757,N_10308,N_13905);
and U25758 (N_25758,N_19128,N_19305);
or U25759 (N_25759,N_16089,N_13350);
and U25760 (N_25760,N_13337,N_18169);
xor U25761 (N_25761,N_12486,N_16379);
and U25762 (N_25762,N_10068,N_18622);
nand U25763 (N_25763,N_16705,N_14241);
nand U25764 (N_25764,N_10148,N_14905);
xor U25765 (N_25765,N_17541,N_19010);
xnor U25766 (N_25766,N_18828,N_12677);
nor U25767 (N_25767,N_19954,N_17660);
nand U25768 (N_25768,N_13687,N_19748);
nor U25769 (N_25769,N_19613,N_15845);
nand U25770 (N_25770,N_15412,N_14432);
xnor U25771 (N_25771,N_17447,N_17510);
nand U25772 (N_25772,N_16243,N_11483);
or U25773 (N_25773,N_10666,N_15904);
nand U25774 (N_25774,N_10310,N_12087);
or U25775 (N_25775,N_15767,N_18658);
xnor U25776 (N_25776,N_14879,N_16628);
and U25777 (N_25777,N_12233,N_10558);
and U25778 (N_25778,N_14792,N_15895);
xor U25779 (N_25779,N_12824,N_10735);
nand U25780 (N_25780,N_11121,N_16783);
and U25781 (N_25781,N_19134,N_11259);
nand U25782 (N_25782,N_17469,N_14559);
or U25783 (N_25783,N_17515,N_14373);
nor U25784 (N_25784,N_12202,N_11897);
and U25785 (N_25785,N_10002,N_19237);
or U25786 (N_25786,N_13860,N_15000);
or U25787 (N_25787,N_19673,N_11943);
and U25788 (N_25788,N_19987,N_16963);
nor U25789 (N_25789,N_12077,N_14655);
and U25790 (N_25790,N_11614,N_13538);
xnor U25791 (N_25791,N_10315,N_17951);
or U25792 (N_25792,N_19514,N_18780);
nand U25793 (N_25793,N_17833,N_10362);
nand U25794 (N_25794,N_15317,N_16959);
or U25795 (N_25795,N_14033,N_14837);
and U25796 (N_25796,N_12627,N_11914);
nor U25797 (N_25797,N_19241,N_18628);
and U25798 (N_25798,N_15041,N_19465);
and U25799 (N_25799,N_14391,N_15665);
or U25800 (N_25800,N_15363,N_17093);
and U25801 (N_25801,N_13863,N_17304);
nor U25802 (N_25802,N_16267,N_18535);
and U25803 (N_25803,N_14901,N_15093);
or U25804 (N_25804,N_17551,N_12620);
nor U25805 (N_25805,N_17440,N_17866);
and U25806 (N_25806,N_13046,N_17474);
xnor U25807 (N_25807,N_10041,N_16146);
and U25808 (N_25808,N_10647,N_10533);
xnor U25809 (N_25809,N_10688,N_11071);
or U25810 (N_25810,N_19872,N_13650);
nand U25811 (N_25811,N_15766,N_11433);
nand U25812 (N_25812,N_19511,N_14101);
and U25813 (N_25813,N_19283,N_11913);
xor U25814 (N_25814,N_17936,N_14490);
nor U25815 (N_25815,N_13894,N_11285);
nand U25816 (N_25816,N_13444,N_10984);
nand U25817 (N_25817,N_16562,N_10154);
xnor U25818 (N_25818,N_19884,N_15680);
and U25819 (N_25819,N_18138,N_11638);
or U25820 (N_25820,N_18509,N_10548);
nor U25821 (N_25821,N_17842,N_16259);
xnor U25822 (N_25822,N_16601,N_16914);
xor U25823 (N_25823,N_17758,N_18932);
and U25824 (N_25824,N_15035,N_16219);
and U25825 (N_25825,N_13410,N_17739);
and U25826 (N_25826,N_14722,N_18489);
and U25827 (N_25827,N_18653,N_10497);
xnor U25828 (N_25828,N_10599,N_16384);
or U25829 (N_25829,N_19780,N_16481);
xor U25830 (N_25830,N_10562,N_15263);
or U25831 (N_25831,N_16028,N_18505);
nor U25832 (N_25832,N_12863,N_15630);
or U25833 (N_25833,N_18803,N_19242);
xnor U25834 (N_25834,N_11112,N_11732);
or U25835 (N_25835,N_16182,N_16593);
nor U25836 (N_25836,N_15299,N_17004);
or U25837 (N_25837,N_18819,N_18132);
and U25838 (N_25838,N_18983,N_14744);
xor U25839 (N_25839,N_16226,N_14175);
nand U25840 (N_25840,N_12327,N_19100);
or U25841 (N_25841,N_13489,N_10936);
nand U25842 (N_25842,N_11822,N_14590);
nor U25843 (N_25843,N_19263,N_13745);
and U25844 (N_25844,N_11383,N_15464);
nand U25845 (N_25845,N_17302,N_11338);
nor U25846 (N_25846,N_19109,N_17513);
nand U25847 (N_25847,N_13177,N_19256);
or U25848 (N_25848,N_19501,N_11483);
and U25849 (N_25849,N_15150,N_13414);
or U25850 (N_25850,N_16990,N_10096);
and U25851 (N_25851,N_13006,N_18666);
or U25852 (N_25852,N_14045,N_13316);
or U25853 (N_25853,N_13316,N_18933);
nand U25854 (N_25854,N_12624,N_19959);
nor U25855 (N_25855,N_12068,N_18019);
and U25856 (N_25856,N_17381,N_16371);
xor U25857 (N_25857,N_19178,N_17655);
or U25858 (N_25858,N_13536,N_10804);
xor U25859 (N_25859,N_12111,N_11208);
nand U25860 (N_25860,N_16614,N_13713);
or U25861 (N_25861,N_18517,N_15436);
nor U25862 (N_25862,N_19489,N_18425);
nand U25863 (N_25863,N_18603,N_13541);
xnor U25864 (N_25864,N_17412,N_15081);
xor U25865 (N_25865,N_18033,N_17663);
and U25866 (N_25866,N_11137,N_13877);
nor U25867 (N_25867,N_17302,N_14252);
xor U25868 (N_25868,N_14266,N_18132);
and U25869 (N_25869,N_13299,N_10130);
nor U25870 (N_25870,N_10955,N_15064);
nand U25871 (N_25871,N_15872,N_13687);
and U25872 (N_25872,N_11374,N_17396);
nor U25873 (N_25873,N_10825,N_16536);
nor U25874 (N_25874,N_18622,N_18247);
nand U25875 (N_25875,N_12264,N_15071);
and U25876 (N_25876,N_15304,N_10117);
and U25877 (N_25877,N_19053,N_10980);
nand U25878 (N_25878,N_18459,N_19372);
nor U25879 (N_25879,N_13951,N_11391);
and U25880 (N_25880,N_19467,N_16129);
xor U25881 (N_25881,N_11005,N_19727);
xnor U25882 (N_25882,N_18125,N_12402);
nand U25883 (N_25883,N_14206,N_11650);
xor U25884 (N_25884,N_16016,N_19168);
nand U25885 (N_25885,N_10523,N_11490);
xnor U25886 (N_25886,N_17914,N_17058);
xor U25887 (N_25887,N_19530,N_12326);
nand U25888 (N_25888,N_11454,N_14736);
or U25889 (N_25889,N_18782,N_10865);
nand U25890 (N_25890,N_10946,N_14385);
xor U25891 (N_25891,N_19681,N_18790);
nand U25892 (N_25892,N_13650,N_11843);
nand U25893 (N_25893,N_13620,N_19702);
nor U25894 (N_25894,N_14316,N_14135);
or U25895 (N_25895,N_11747,N_14433);
and U25896 (N_25896,N_16707,N_16003);
nor U25897 (N_25897,N_14421,N_18087);
nor U25898 (N_25898,N_10744,N_17799);
xnor U25899 (N_25899,N_18087,N_12890);
and U25900 (N_25900,N_16327,N_10549);
nand U25901 (N_25901,N_10137,N_18979);
nor U25902 (N_25902,N_19230,N_16061);
nand U25903 (N_25903,N_19865,N_16158);
xor U25904 (N_25904,N_18779,N_10738);
xor U25905 (N_25905,N_13422,N_18949);
and U25906 (N_25906,N_11963,N_12212);
nand U25907 (N_25907,N_19005,N_18928);
and U25908 (N_25908,N_16397,N_10849);
nand U25909 (N_25909,N_19046,N_11921);
and U25910 (N_25910,N_15324,N_11515);
nand U25911 (N_25911,N_13063,N_10489);
and U25912 (N_25912,N_19352,N_10470);
xnor U25913 (N_25913,N_11442,N_18940);
and U25914 (N_25914,N_13614,N_13611);
and U25915 (N_25915,N_15552,N_14193);
and U25916 (N_25916,N_13876,N_17609);
or U25917 (N_25917,N_13396,N_10162);
nand U25918 (N_25918,N_10724,N_11771);
or U25919 (N_25919,N_18690,N_12266);
xor U25920 (N_25920,N_13015,N_10547);
or U25921 (N_25921,N_17823,N_15650);
nand U25922 (N_25922,N_17004,N_16737);
nor U25923 (N_25923,N_12164,N_16707);
and U25924 (N_25924,N_18533,N_10115);
nor U25925 (N_25925,N_15996,N_15216);
xnor U25926 (N_25926,N_12105,N_14182);
nor U25927 (N_25927,N_10050,N_19650);
nand U25928 (N_25928,N_10539,N_14922);
xor U25929 (N_25929,N_16837,N_10641);
and U25930 (N_25930,N_10876,N_16105);
nor U25931 (N_25931,N_11062,N_13422);
or U25932 (N_25932,N_11333,N_11993);
or U25933 (N_25933,N_19018,N_16097);
nand U25934 (N_25934,N_10308,N_16070);
or U25935 (N_25935,N_10310,N_13016);
nand U25936 (N_25936,N_13488,N_16913);
or U25937 (N_25937,N_19338,N_12527);
and U25938 (N_25938,N_16841,N_11019);
xnor U25939 (N_25939,N_16695,N_14281);
and U25940 (N_25940,N_14548,N_18886);
nor U25941 (N_25941,N_13047,N_10550);
xor U25942 (N_25942,N_16968,N_14590);
nor U25943 (N_25943,N_16586,N_19803);
nor U25944 (N_25944,N_12071,N_10176);
and U25945 (N_25945,N_10548,N_16161);
and U25946 (N_25946,N_16873,N_19620);
nor U25947 (N_25947,N_11739,N_15583);
and U25948 (N_25948,N_13296,N_12300);
and U25949 (N_25949,N_18704,N_15796);
nor U25950 (N_25950,N_15194,N_18596);
nand U25951 (N_25951,N_13504,N_16565);
and U25952 (N_25952,N_19084,N_13643);
nand U25953 (N_25953,N_16961,N_13664);
and U25954 (N_25954,N_19840,N_11020);
xnor U25955 (N_25955,N_13139,N_13726);
and U25956 (N_25956,N_10471,N_19040);
and U25957 (N_25957,N_15069,N_16610);
nand U25958 (N_25958,N_11117,N_19678);
or U25959 (N_25959,N_12950,N_16001);
nand U25960 (N_25960,N_12274,N_10686);
nor U25961 (N_25961,N_15327,N_19688);
nand U25962 (N_25962,N_12461,N_11923);
nand U25963 (N_25963,N_16748,N_15392);
nand U25964 (N_25964,N_19859,N_14935);
and U25965 (N_25965,N_19656,N_12003);
and U25966 (N_25966,N_10271,N_13404);
xor U25967 (N_25967,N_19733,N_13082);
nor U25968 (N_25968,N_13391,N_17506);
nand U25969 (N_25969,N_17457,N_16647);
nor U25970 (N_25970,N_15032,N_15953);
and U25971 (N_25971,N_17571,N_13434);
or U25972 (N_25972,N_10559,N_10418);
nand U25973 (N_25973,N_12340,N_11152);
xor U25974 (N_25974,N_12298,N_10842);
and U25975 (N_25975,N_10402,N_16010);
xor U25976 (N_25976,N_10179,N_12596);
and U25977 (N_25977,N_11167,N_17243);
nor U25978 (N_25978,N_19881,N_12719);
and U25979 (N_25979,N_10549,N_13453);
or U25980 (N_25980,N_14032,N_19843);
nor U25981 (N_25981,N_12615,N_19816);
or U25982 (N_25982,N_11371,N_18676);
xor U25983 (N_25983,N_16311,N_18103);
nand U25984 (N_25984,N_14263,N_16187);
and U25985 (N_25985,N_14294,N_12816);
nor U25986 (N_25986,N_14982,N_10803);
xnor U25987 (N_25987,N_19502,N_10167);
xnor U25988 (N_25988,N_17186,N_14240);
and U25989 (N_25989,N_18884,N_12566);
nor U25990 (N_25990,N_10867,N_18885);
or U25991 (N_25991,N_13640,N_10227);
nand U25992 (N_25992,N_12922,N_17135);
nand U25993 (N_25993,N_10471,N_13640);
xnor U25994 (N_25994,N_15965,N_15035);
nand U25995 (N_25995,N_15150,N_18174);
and U25996 (N_25996,N_17183,N_14954);
or U25997 (N_25997,N_16006,N_17731);
xnor U25998 (N_25998,N_15784,N_16088);
xor U25999 (N_25999,N_11271,N_13409);
or U26000 (N_26000,N_14843,N_18597);
or U26001 (N_26001,N_15431,N_13254);
nand U26002 (N_26002,N_16831,N_10309);
xor U26003 (N_26003,N_16971,N_14694);
xnor U26004 (N_26004,N_15777,N_13549);
nand U26005 (N_26005,N_17629,N_14216);
nor U26006 (N_26006,N_18783,N_16131);
nand U26007 (N_26007,N_18759,N_14690);
nor U26008 (N_26008,N_15590,N_15625);
nand U26009 (N_26009,N_10433,N_12821);
nor U26010 (N_26010,N_19027,N_10717);
nor U26011 (N_26011,N_12094,N_14964);
and U26012 (N_26012,N_19240,N_16379);
xor U26013 (N_26013,N_15891,N_15866);
xnor U26014 (N_26014,N_16333,N_18861);
nor U26015 (N_26015,N_17201,N_11539);
and U26016 (N_26016,N_10231,N_16443);
nor U26017 (N_26017,N_13050,N_17288);
xor U26018 (N_26018,N_12556,N_15758);
nor U26019 (N_26019,N_15616,N_19495);
nor U26020 (N_26020,N_17796,N_12218);
nand U26021 (N_26021,N_18544,N_14923);
nor U26022 (N_26022,N_11489,N_10617);
xor U26023 (N_26023,N_14300,N_19926);
or U26024 (N_26024,N_19383,N_16559);
or U26025 (N_26025,N_13799,N_18535);
or U26026 (N_26026,N_17699,N_12134);
or U26027 (N_26027,N_16642,N_11929);
and U26028 (N_26028,N_19903,N_11902);
nand U26029 (N_26029,N_17902,N_15275);
nor U26030 (N_26030,N_10390,N_18306);
nor U26031 (N_26031,N_15335,N_10755);
and U26032 (N_26032,N_14780,N_19399);
and U26033 (N_26033,N_15601,N_11508);
and U26034 (N_26034,N_19470,N_13316);
xnor U26035 (N_26035,N_18347,N_14694);
or U26036 (N_26036,N_15624,N_15797);
nand U26037 (N_26037,N_18252,N_13090);
or U26038 (N_26038,N_18858,N_10483);
nand U26039 (N_26039,N_15386,N_12992);
nor U26040 (N_26040,N_15623,N_18215);
or U26041 (N_26041,N_11008,N_18849);
xnor U26042 (N_26042,N_12192,N_15151);
xnor U26043 (N_26043,N_11301,N_11336);
nor U26044 (N_26044,N_18622,N_17516);
and U26045 (N_26045,N_17268,N_15091);
or U26046 (N_26046,N_10443,N_16823);
or U26047 (N_26047,N_10113,N_12756);
or U26048 (N_26048,N_13563,N_18041);
xnor U26049 (N_26049,N_10319,N_16691);
and U26050 (N_26050,N_18638,N_10712);
or U26051 (N_26051,N_15155,N_15531);
and U26052 (N_26052,N_18948,N_19523);
and U26053 (N_26053,N_15010,N_18182);
and U26054 (N_26054,N_15037,N_18418);
nor U26055 (N_26055,N_17800,N_18625);
and U26056 (N_26056,N_16690,N_13788);
xnor U26057 (N_26057,N_14677,N_10343);
xnor U26058 (N_26058,N_16104,N_14967);
and U26059 (N_26059,N_19036,N_12867);
and U26060 (N_26060,N_11357,N_16016);
xnor U26061 (N_26061,N_18148,N_12559);
nor U26062 (N_26062,N_18216,N_19618);
or U26063 (N_26063,N_19423,N_17394);
or U26064 (N_26064,N_19516,N_17791);
and U26065 (N_26065,N_10591,N_16703);
nand U26066 (N_26066,N_10371,N_14290);
xnor U26067 (N_26067,N_13997,N_14439);
and U26068 (N_26068,N_17702,N_18068);
or U26069 (N_26069,N_19948,N_15464);
nand U26070 (N_26070,N_19066,N_12220);
nand U26071 (N_26071,N_11854,N_10278);
nor U26072 (N_26072,N_13528,N_13941);
or U26073 (N_26073,N_19094,N_12903);
nor U26074 (N_26074,N_11708,N_14318);
or U26075 (N_26075,N_11674,N_13591);
nor U26076 (N_26076,N_19965,N_10921);
nor U26077 (N_26077,N_11713,N_19963);
xor U26078 (N_26078,N_11411,N_12007);
xnor U26079 (N_26079,N_13661,N_14996);
nand U26080 (N_26080,N_16089,N_18311);
nand U26081 (N_26081,N_14656,N_14098);
xnor U26082 (N_26082,N_13701,N_18543);
nor U26083 (N_26083,N_15888,N_18540);
and U26084 (N_26084,N_18903,N_19239);
nand U26085 (N_26085,N_18258,N_12903);
xor U26086 (N_26086,N_12103,N_14452);
nor U26087 (N_26087,N_13116,N_17418);
nand U26088 (N_26088,N_13251,N_18007);
or U26089 (N_26089,N_17207,N_15492);
or U26090 (N_26090,N_10037,N_15867);
nand U26091 (N_26091,N_19637,N_16102);
xnor U26092 (N_26092,N_17173,N_11187);
or U26093 (N_26093,N_11814,N_10142);
xor U26094 (N_26094,N_14037,N_15053);
or U26095 (N_26095,N_10694,N_11456);
nand U26096 (N_26096,N_17796,N_19775);
and U26097 (N_26097,N_16990,N_17992);
and U26098 (N_26098,N_18817,N_11000);
nand U26099 (N_26099,N_17472,N_11785);
nor U26100 (N_26100,N_19787,N_16221);
nor U26101 (N_26101,N_15721,N_16998);
nand U26102 (N_26102,N_12941,N_15780);
and U26103 (N_26103,N_11188,N_17816);
nor U26104 (N_26104,N_18640,N_15399);
nand U26105 (N_26105,N_16711,N_11794);
xnor U26106 (N_26106,N_14346,N_13092);
or U26107 (N_26107,N_18623,N_18863);
nand U26108 (N_26108,N_10227,N_17749);
nor U26109 (N_26109,N_16313,N_16432);
or U26110 (N_26110,N_14460,N_18486);
nand U26111 (N_26111,N_17754,N_17064);
nor U26112 (N_26112,N_17074,N_17374);
nor U26113 (N_26113,N_11027,N_18237);
nor U26114 (N_26114,N_10424,N_10713);
and U26115 (N_26115,N_10930,N_17853);
nand U26116 (N_26116,N_10689,N_10356);
and U26117 (N_26117,N_15898,N_19076);
xnor U26118 (N_26118,N_18822,N_18248);
nand U26119 (N_26119,N_12254,N_16132);
nand U26120 (N_26120,N_12085,N_18121);
xnor U26121 (N_26121,N_11728,N_14902);
and U26122 (N_26122,N_18872,N_15112);
xor U26123 (N_26123,N_16152,N_11289);
nand U26124 (N_26124,N_19182,N_15479);
xor U26125 (N_26125,N_10863,N_12609);
nor U26126 (N_26126,N_17649,N_15560);
or U26127 (N_26127,N_11331,N_19217);
nand U26128 (N_26128,N_19184,N_11158);
or U26129 (N_26129,N_12706,N_13574);
nor U26130 (N_26130,N_14899,N_15136);
nand U26131 (N_26131,N_16650,N_11293);
or U26132 (N_26132,N_16853,N_13586);
or U26133 (N_26133,N_17329,N_11480);
and U26134 (N_26134,N_10635,N_16859);
nand U26135 (N_26135,N_11071,N_10595);
nand U26136 (N_26136,N_16366,N_13049);
nand U26137 (N_26137,N_16596,N_12351);
and U26138 (N_26138,N_18242,N_19099);
nor U26139 (N_26139,N_13300,N_15454);
or U26140 (N_26140,N_15668,N_15044);
or U26141 (N_26141,N_11389,N_15537);
nor U26142 (N_26142,N_18406,N_15469);
nor U26143 (N_26143,N_13277,N_10547);
nand U26144 (N_26144,N_13509,N_16011);
nor U26145 (N_26145,N_13151,N_13817);
nor U26146 (N_26146,N_16480,N_18061);
nand U26147 (N_26147,N_18976,N_16710);
and U26148 (N_26148,N_19970,N_17170);
nand U26149 (N_26149,N_19158,N_14977);
nor U26150 (N_26150,N_16232,N_10211);
and U26151 (N_26151,N_19779,N_19670);
nand U26152 (N_26152,N_13861,N_19912);
or U26153 (N_26153,N_11678,N_17616);
nand U26154 (N_26154,N_16604,N_13846);
and U26155 (N_26155,N_17283,N_17992);
nor U26156 (N_26156,N_16724,N_15205);
or U26157 (N_26157,N_14053,N_15716);
nand U26158 (N_26158,N_15466,N_16111);
xor U26159 (N_26159,N_17588,N_16735);
or U26160 (N_26160,N_16850,N_16929);
nor U26161 (N_26161,N_14611,N_15193);
and U26162 (N_26162,N_11659,N_15993);
or U26163 (N_26163,N_16109,N_16373);
nor U26164 (N_26164,N_15867,N_18821);
xor U26165 (N_26165,N_15213,N_16680);
nor U26166 (N_26166,N_19162,N_12527);
nor U26167 (N_26167,N_15179,N_10481);
xnor U26168 (N_26168,N_18447,N_19449);
nor U26169 (N_26169,N_17731,N_11177);
nand U26170 (N_26170,N_14884,N_17608);
or U26171 (N_26171,N_10280,N_17234);
or U26172 (N_26172,N_17916,N_11621);
and U26173 (N_26173,N_16837,N_12168);
or U26174 (N_26174,N_10873,N_13669);
xor U26175 (N_26175,N_10497,N_10122);
and U26176 (N_26176,N_19461,N_15460);
xor U26177 (N_26177,N_15795,N_18647);
nand U26178 (N_26178,N_18040,N_15235);
and U26179 (N_26179,N_19190,N_12821);
or U26180 (N_26180,N_19999,N_16631);
nor U26181 (N_26181,N_14945,N_12971);
and U26182 (N_26182,N_18354,N_12624);
nor U26183 (N_26183,N_17199,N_18092);
xnor U26184 (N_26184,N_10247,N_12279);
and U26185 (N_26185,N_13753,N_19541);
nand U26186 (N_26186,N_12501,N_13003);
and U26187 (N_26187,N_11122,N_15850);
nor U26188 (N_26188,N_15479,N_10615);
nor U26189 (N_26189,N_12503,N_12723);
xnor U26190 (N_26190,N_12348,N_18732);
or U26191 (N_26191,N_18367,N_12659);
or U26192 (N_26192,N_13955,N_16363);
xnor U26193 (N_26193,N_16620,N_13042);
and U26194 (N_26194,N_10761,N_18771);
nor U26195 (N_26195,N_14516,N_15863);
and U26196 (N_26196,N_10839,N_18777);
xnor U26197 (N_26197,N_15588,N_17459);
and U26198 (N_26198,N_14177,N_11531);
nand U26199 (N_26199,N_18584,N_14453);
nand U26200 (N_26200,N_18612,N_12081);
or U26201 (N_26201,N_15523,N_15126);
nor U26202 (N_26202,N_11167,N_12785);
xor U26203 (N_26203,N_11246,N_11867);
nand U26204 (N_26204,N_12724,N_17099);
and U26205 (N_26205,N_17189,N_11971);
nand U26206 (N_26206,N_17763,N_10377);
nor U26207 (N_26207,N_10154,N_16717);
xnor U26208 (N_26208,N_14403,N_18910);
xor U26209 (N_26209,N_16959,N_11607);
and U26210 (N_26210,N_19142,N_19407);
nand U26211 (N_26211,N_16431,N_15919);
and U26212 (N_26212,N_13563,N_14069);
nor U26213 (N_26213,N_19728,N_19362);
nand U26214 (N_26214,N_18396,N_16186);
nor U26215 (N_26215,N_12604,N_13916);
xnor U26216 (N_26216,N_14579,N_17955);
and U26217 (N_26217,N_18192,N_18803);
or U26218 (N_26218,N_10239,N_12612);
xor U26219 (N_26219,N_14293,N_10614);
xnor U26220 (N_26220,N_19766,N_13025);
or U26221 (N_26221,N_15513,N_12645);
or U26222 (N_26222,N_13531,N_11875);
and U26223 (N_26223,N_18243,N_16490);
and U26224 (N_26224,N_10520,N_12359);
or U26225 (N_26225,N_17468,N_11917);
or U26226 (N_26226,N_15936,N_18186);
nor U26227 (N_26227,N_16830,N_10691);
nor U26228 (N_26228,N_10005,N_17300);
xnor U26229 (N_26229,N_19732,N_17443);
nor U26230 (N_26230,N_15061,N_16341);
or U26231 (N_26231,N_10834,N_12905);
xnor U26232 (N_26232,N_13989,N_13766);
and U26233 (N_26233,N_11975,N_11798);
xor U26234 (N_26234,N_18651,N_17156);
xor U26235 (N_26235,N_16364,N_17191);
nand U26236 (N_26236,N_12308,N_17160);
and U26237 (N_26237,N_13621,N_11277);
nor U26238 (N_26238,N_19075,N_10790);
or U26239 (N_26239,N_18493,N_16508);
and U26240 (N_26240,N_19588,N_14945);
and U26241 (N_26241,N_14634,N_12049);
nor U26242 (N_26242,N_12772,N_11072);
or U26243 (N_26243,N_16893,N_11800);
nor U26244 (N_26244,N_13905,N_13937);
nor U26245 (N_26245,N_14787,N_14119);
or U26246 (N_26246,N_11986,N_13602);
xnor U26247 (N_26247,N_14296,N_17336);
nor U26248 (N_26248,N_19961,N_11502);
xor U26249 (N_26249,N_17225,N_10241);
or U26250 (N_26250,N_15644,N_17641);
nand U26251 (N_26251,N_10461,N_16911);
or U26252 (N_26252,N_13279,N_14322);
or U26253 (N_26253,N_11429,N_18135);
nor U26254 (N_26254,N_18044,N_14405);
nand U26255 (N_26255,N_11083,N_11543);
and U26256 (N_26256,N_14171,N_18129);
or U26257 (N_26257,N_14703,N_12448);
and U26258 (N_26258,N_15536,N_13457);
xnor U26259 (N_26259,N_10415,N_10492);
and U26260 (N_26260,N_17429,N_10778);
or U26261 (N_26261,N_19981,N_18979);
xnor U26262 (N_26262,N_13394,N_19245);
nand U26263 (N_26263,N_19856,N_13903);
nand U26264 (N_26264,N_11780,N_14102);
nand U26265 (N_26265,N_16637,N_14330);
or U26266 (N_26266,N_15854,N_17710);
or U26267 (N_26267,N_13673,N_16809);
nor U26268 (N_26268,N_15413,N_14901);
nand U26269 (N_26269,N_13458,N_16163);
nand U26270 (N_26270,N_18172,N_17499);
and U26271 (N_26271,N_16753,N_13758);
nand U26272 (N_26272,N_12962,N_19547);
nor U26273 (N_26273,N_15393,N_11394);
and U26274 (N_26274,N_16139,N_15682);
and U26275 (N_26275,N_11555,N_16602);
xor U26276 (N_26276,N_10200,N_11131);
nand U26277 (N_26277,N_17068,N_18967);
and U26278 (N_26278,N_15883,N_10192);
nand U26279 (N_26279,N_11807,N_19854);
nand U26280 (N_26280,N_13900,N_13455);
and U26281 (N_26281,N_11096,N_10470);
and U26282 (N_26282,N_10025,N_13965);
nor U26283 (N_26283,N_14181,N_14804);
nor U26284 (N_26284,N_13630,N_15390);
or U26285 (N_26285,N_19948,N_16554);
nor U26286 (N_26286,N_19708,N_14746);
nor U26287 (N_26287,N_10998,N_18406);
nand U26288 (N_26288,N_19688,N_16752);
nand U26289 (N_26289,N_13082,N_16682);
nand U26290 (N_26290,N_10920,N_15915);
and U26291 (N_26291,N_17379,N_16403);
nor U26292 (N_26292,N_18280,N_17447);
or U26293 (N_26293,N_17306,N_10154);
or U26294 (N_26294,N_18096,N_15936);
or U26295 (N_26295,N_16633,N_17603);
nand U26296 (N_26296,N_18339,N_15903);
xnor U26297 (N_26297,N_17227,N_17023);
nand U26298 (N_26298,N_18159,N_15036);
xor U26299 (N_26299,N_18384,N_14417);
or U26300 (N_26300,N_10930,N_11521);
nand U26301 (N_26301,N_13000,N_17660);
nor U26302 (N_26302,N_11877,N_19327);
xor U26303 (N_26303,N_13664,N_17231);
nor U26304 (N_26304,N_17194,N_12581);
nand U26305 (N_26305,N_17358,N_15693);
nor U26306 (N_26306,N_15289,N_14125);
nor U26307 (N_26307,N_17649,N_12783);
nand U26308 (N_26308,N_11667,N_14626);
or U26309 (N_26309,N_14406,N_10939);
xnor U26310 (N_26310,N_17822,N_13101);
and U26311 (N_26311,N_16049,N_14142);
xor U26312 (N_26312,N_11438,N_17162);
xor U26313 (N_26313,N_13529,N_12453);
nor U26314 (N_26314,N_12278,N_16265);
nor U26315 (N_26315,N_12260,N_16856);
nor U26316 (N_26316,N_17075,N_13005);
nand U26317 (N_26317,N_11315,N_17734);
or U26318 (N_26318,N_11081,N_12159);
and U26319 (N_26319,N_16015,N_19673);
nand U26320 (N_26320,N_14040,N_10092);
or U26321 (N_26321,N_12516,N_14644);
nor U26322 (N_26322,N_13876,N_19165);
or U26323 (N_26323,N_15718,N_11406);
or U26324 (N_26324,N_16412,N_18926);
xnor U26325 (N_26325,N_18637,N_10927);
nand U26326 (N_26326,N_12870,N_17381);
nor U26327 (N_26327,N_19748,N_15662);
and U26328 (N_26328,N_10681,N_16137);
nand U26329 (N_26329,N_15993,N_19732);
or U26330 (N_26330,N_10139,N_19176);
and U26331 (N_26331,N_17643,N_11326);
or U26332 (N_26332,N_15420,N_16408);
nor U26333 (N_26333,N_17513,N_13445);
and U26334 (N_26334,N_15630,N_18744);
or U26335 (N_26335,N_18989,N_12755);
or U26336 (N_26336,N_12058,N_15790);
nor U26337 (N_26337,N_14936,N_14925);
xnor U26338 (N_26338,N_18504,N_11434);
nand U26339 (N_26339,N_11324,N_18786);
nor U26340 (N_26340,N_12903,N_15757);
or U26341 (N_26341,N_10204,N_10821);
nor U26342 (N_26342,N_14746,N_10101);
nor U26343 (N_26343,N_19587,N_17740);
and U26344 (N_26344,N_19998,N_12136);
or U26345 (N_26345,N_14267,N_13565);
nor U26346 (N_26346,N_19537,N_14742);
xnor U26347 (N_26347,N_10950,N_19606);
xnor U26348 (N_26348,N_19089,N_17793);
xor U26349 (N_26349,N_10249,N_12114);
and U26350 (N_26350,N_15779,N_19788);
and U26351 (N_26351,N_19986,N_12362);
xnor U26352 (N_26352,N_12910,N_16599);
xnor U26353 (N_26353,N_12710,N_10326);
or U26354 (N_26354,N_17236,N_17581);
nand U26355 (N_26355,N_14396,N_14230);
nor U26356 (N_26356,N_16969,N_10820);
and U26357 (N_26357,N_13808,N_15296);
nor U26358 (N_26358,N_16395,N_13378);
and U26359 (N_26359,N_10491,N_15460);
and U26360 (N_26360,N_18840,N_19301);
xor U26361 (N_26361,N_16376,N_12980);
or U26362 (N_26362,N_10861,N_12681);
nand U26363 (N_26363,N_12279,N_12078);
nand U26364 (N_26364,N_18529,N_17457);
xnor U26365 (N_26365,N_12787,N_12817);
nor U26366 (N_26366,N_14162,N_12552);
nor U26367 (N_26367,N_14207,N_12168);
nand U26368 (N_26368,N_18139,N_15386);
or U26369 (N_26369,N_19585,N_10223);
nor U26370 (N_26370,N_11996,N_11835);
xor U26371 (N_26371,N_13610,N_15116);
and U26372 (N_26372,N_13121,N_19953);
and U26373 (N_26373,N_11063,N_15143);
nor U26374 (N_26374,N_12654,N_19714);
nand U26375 (N_26375,N_19188,N_14067);
nand U26376 (N_26376,N_11269,N_17774);
or U26377 (N_26377,N_14214,N_13946);
and U26378 (N_26378,N_15293,N_12627);
or U26379 (N_26379,N_12915,N_10658);
or U26380 (N_26380,N_16185,N_13588);
xnor U26381 (N_26381,N_19701,N_11672);
or U26382 (N_26382,N_13227,N_18892);
xnor U26383 (N_26383,N_13807,N_19593);
nand U26384 (N_26384,N_13200,N_17216);
or U26385 (N_26385,N_15080,N_15639);
nor U26386 (N_26386,N_11769,N_16434);
and U26387 (N_26387,N_15987,N_17431);
or U26388 (N_26388,N_13502,N_13001);
or U26389 (N_26389,N_14004,N_12577);
nor U26390 (N_26390,N_12496,N_17194);
and U26391 (N_26391,N_15335,N_13753);
and U26392 (N_26392,N_12710,N_11127);
nand U26393 (N_26393,N_19497,N_11564);
and U26394 (N_26394,N_13066,N_13657);
and U26395 (N_26395,N_10591,N_11259);
and U26396 (N_26396,N_11288,N_11104);
nor U26397 (N_26397,N_16428,N_17811);
xnor U26398 (N_26398,N_18978,N_10713);
nor U26399 (N_26399,N_12885,N_11730);
and U26400 (N_26400,N_13778,N_17743);
nor U26401 (N_26401,N_10799,N_10830);
or U26402 (N_26402,N_11669,N_19319);
or U26403 (N_26403,N_15142,N_19203);
or U26404 (N_26404,N_16793,N_10117);
or U26405 (N_26405,N_10209,N_15260);
nor U26406 (N_26406,N_16303,N_17959);
nand U26407 (N_26407,N_18297,N_19102);
or U26408 (N_26408,N_12017,N_14056);
or U26409 (N_26409,N_13127,N_17198);
nand U26410 (N_26410,N_10059,N_16638);
or U26411 (N_26411,N_11473,N_12104);
or U26412 (N_26412,N_13165,N_19385);
and U26413 (N_26413,N_17415,N_12420);
xnor U26414 (N_26414,N_16370,N_14401);
nand U26415 (N_26415,N_11308,N_11881);
or U26416 (N_26416,N_19675,N_13164);
and U26417 (N_26417,N_16273,N_10930);
xor U26418 (N_26418,N_10185,N_10387);
and U26419 (N_26419,N_11425,N_19734);
and U26420 (N_26420,N_13539,N_16077);
nand U26421 (N_26421,N_16948,N_13434);
nor U26422 (N_26422,N_11644,N_15317);
nand U26423 (N_26423,N_18403,N_18694);
and U26424 (N_26424,N_16325,N_19155);
xor U26425 (N_26425,N_14092,N_10681);
nor U26426 (N_26426,N_17876,N_11068);
xor U26427 (N_26427,N_15547,N_17489);
nor U26428 (N_26428,N_10700,N_16697);
or U26429 (N_26429,N_10216,N_17838);
or U26430 (N_26430,N_13182,N_12320);
nand U26431 (N_26431,N_14466,N_13247);
and U26432 (N_26432,N_15260,N_12123);
nor U26433 (N_26433,N_13452,N_13607);
nor U26434 (N_26434,N_10595,N_11682);
xnor U26435 (N_26435,N_13487,N_17245);
xnor U26436 (N_26436,N_17980,N_19521);
nand U26437 (N_26437,N_14010,N_18170);
and U26438 (N_26438,N_19045,N_19515);
or U26439 (N_26439,N_19538,N_16356);
and U26440 (N_26440,N_16558,N_12986);
xnor U26441 (N_26441,N_15986,N_17549);
nand U26442 (N_26442,N_16868,N_19325);
and U26443 (N_26443,N_16939,N_17874);
nor U26444 (N_26444,N_17640,N_18741);
xnor U26445 (N_26445,N_13513,N_18634);
nand U26446 (N_26446,N_10980,N_19293);
xnor U26447 (N_26447,N_15486,N_11763);
xnor U26448 (N_26448,N_15975,N_17732);
nor U26449 (N_26449,N_14384,N_15829);
and U26450 (N_26450,N_14044,N_11644);
or U26451 (N_26451,N_17671,N_19755);
and U26452 (N_26452,N_19897,N_16308);
or U26453 (N_26453,N_16904,N_12662);
nand U26454 (N_26454,N_18165,N_17533);
and U26455 (N_26455,N_19988,N_10451);
xor U26456 (N_26456,N_12773,N_12163);
or U26457 (N_26457,N_17335,N_13644);
xnor U26458 (N_26458,N_12843,N_19687);
or U26459 (N_26459,N_13760,N_16356);
nand U26460 (N_26460,N_10554,N_12761);
nand U26461 (N_26461,N_13078,N_17355);
or U26462 (N_26462,N_18818,N_16193);
or U26463 (N_26463,N_14541,N_12908);
or U26464 (N_26464,N_15499,N_18286);
xor U26465 (N_26465,N_19149,N_10714);
xnor U26466 (N_26466,N_16564,N_15242);
xnor U26467 (N_26467,N_10403,N_19932);
nor U26468 (N_26468,N_16588,N_14661);
xor U26469 (N_26469,N_15140,N_13869);
nor U26470 (N_26470,N_13652,N_10330);
or U26471 (N_26471,N_14420,N_17434);
xnor U26472 (N_26472,N_15786,N_17463);
nand U26473 (N_26473,N_16946,N_19603);
or U26474 (N_26474,N_19803,N_16496);
xnor U26475 (N_26475,N_17662,N_14219);
xnor U26476 (N_26476,N_13259,N_15709);
and U26477 (N_26477,N_15630,N_10043);
nor U26478 (N_26478,N_15809,N_19413);
nor U26479 (N_26479,N_12843,N_15666);
nor U26480 (N_26480,N_12357,N_16039);
nor U26481 (N_26481,N_18381,N_17400);
nor U26482 (N_26482,N_17083,N_10599);
xor U26483 (N_26483,N_14866,N_15808);
nand U26484 (N_26484,N_19078,N_12279);
nand U26485 (N_26485,N_17864,N_12485);
and U26486 (N_26486,N_18062,N_12196);
xor U26487 (N_26487,N_17454,N_10389);
xnor U26488 (N_26488,N_15860,N_13804);
xor U26489 (N_26489,N_16089,N_13567);
and U26490 (N_26490,N_17691,N_19802);
nand U26491 (N_26491,N_16896,N_12577);
or U26492 (N_26492,N_11016,N_15457);
or U26493 (N_26493,N_15784,N_15762);
xnor U26494 (N_26494,N_12997,N_10278);
nor U26495 (N_26495,N_17600,N_12034);
xnor U26496 (N_26496,N_13767,N_10703);
and U26497 (N_26497,N_12302,N_15949);
and U26498 (N_26498,N_17386,N_11178);
xnor U26499 (N_26499,N_16546,N_12985);
nor U26500 (N_26500,N_11612,N_15160);
nand U26501 (N_26501,N_15618,N_15644);
nor U26502 (N_26502,N_15375,N_15945);
xnor U26503 (N_26503,N_18874,N_13989);
and U26504 (N_26504,N_12283,N_10976);
and U26505 (N_26505,N_16365,N_10879);
nor U26506 (N_26506,N_14766,N_12272);
and U26507 (N_26507,N_15819,N_11767);
nor U26508 (N_26508,N_10742,N_17451);
xor U26509 (N_26509,N_13094,N_14721);
or U26510 (N_26510,N_11800,N_12152);
nor U26511 (N_26511,N_16456,N_10217);
and U26512 (N_26512,N_17848,N_15136);
nand U26513 (N_26513,N_18087,N_10307);
and U26514 (N_26514,N_13014,N_15449);
and U26515 (N_26515,N_18607,N_19373);
and U26516 (N_26516,N_14098,N_16374);
nor U26517 (N_26517,N_11208,N_19713);
xnor U26518 (N_26518,N_14773,N_11512);
xnor U26519 (N_26519,N_13304,N_19133);
or U26520 (N_26520,N_17750,N_17093);
or U26521 (N_26521,N_10845,N_19529);
or U26522 (N_26522,N_19730,N_11236);
or U26523 (N_26523,N_16541,N_16570);
nand U26524 (N_26524,N_19362,N_13188);
and U26525 (N_26525,N_18336,N_16716);
nand U26526 (N_26526,N_18582,N_19911);
or U26527 (N_26527,N_13784,N_12139);
or U26528 (N_26528,N_15565,N_11410);
and U26529 (N_26529,N_12079,N_12502);
nor U26530 (N_26530,N_10976,N_19168);
nand U26531 (N_26531,N_10121,N_14231);
nand U26532 (N_26532,N_16056,N_13920);
or U26533 (N_26533,N_17835,N_18369);
or U26534 (N_26534,N_11347,N_17063);
nand U26535 (N_26535,N_19995,N_12879);
xor U26536 (N_26536,N_10645,N_17320);
xnor U26537 (N_26537,N_19360,N_14129);
or U26538 (N_26538,N_14358,N_18518);
nor U26539 (N_26539,N_12153,N_19072);
or U26540 (N_26540,N_11870,N_13534);
xor U26541 (N_26541,N_19003,N_13529);
nand U26542 (N_26542,N_19370,N_11069);
and U26543 (N_26543,N_11961,N_15249);
and U26544 (N_26544,N_16266,N_15359);
and U26545 (N_26545,N_18327,N_17754);
xor U26546 (N_26546,N_12967,N_19965);
nor U26547 (N_26547,N_15602,N_13125);
nand U26548 (N_26548,N_16852,N_16167);
nand U26549 (N_26549,N_12625,N_15309);
and U26550 (N_26550,N_17942,N_14709);
or U26551 (N_26551,N_12326,N_17186);
nand U26552 (N_26552,N_17304,N_14289);
xor U26553 (N_26553,N_13469,N_13336);
and U26554 (N_26554,N_17972,N_10451);
nand U26555 (N_26555,N_16384,N_16961);
and U26556 (N_26556,N_11070,N_13382);
nor U26557 (N_26557,N_11090,N_11668);
and U26558 (N_26558,N_19274,N_17448);
xnor U26559 (N_26559,N_11554,N_18802);
nand U26560 (N_26560,N_10782,N_14805);
or U26561 (N_26561,N_10628,N_12943);
nand U26562 (N_26562,N_19535,N_11788);
nand U26563 (N_26563,N_13249,N_16901);
or U26564 (N_26564,N_13373,N_14646);
or U26565 (N_26565,N_12336,N_17733);
and U26566 (N_26566,N_16553,N_13814);
or U26567 (N_26567,N_16307,N_17861);
and U26568 (N_26568,N_19361,N_14981);
and U26569 (N_26569,N_16004,N_15243);
or U26570 (N_26570,N_18386,N_17591);
nand U26571 (N_26571,N_11545,N_16960);
nand U26572 (N_26572,N_14074,N_17380);
and U26573 (N_26573,N_16499,N_14876);
and U26574 (N_26574,N_12958,N_17485);
nand U26575 (N_26575,N_19134,N_12925);
or U26576 (N_26576,N_14880,N_11090);
and U26577 (N_26577,N_19621,N_18042);
xnor U26578 (N_26578,N_12145,N_14789);
or U26579 (N_26579,N_19303,N_13410);
and U26580 (N_26580,N_10123,N_10009);
and U26581 (N_26581,N_17621,N_14253);
nand U26582 (N_26582,N_12220,N_17445);
nor U26583 (N_26583,N_14137,N_12677);
nand U26584 (N_26584,N_15647,N_15245);
nand U26585 (N_26585,N_15947,N_19081);
nor U26586 (N_26586,N_11085,N_12744);
nor U26587 (N_26587,N_17831,N_10560);
nand U26588 (N_26588,N_18053,N_16832);
nor U26589 (N_26589,N_19817,N_13137);
and U26590 (N_26590,N_14449,N_16537);
nor U26591 (N_26591,N_18804,N_17884);
nand U26592 (N_26592,N_14752,N_15154);
xnor U26593 (N_26593,N_17634,N_12788);
nor U26594 (N_26594,N_11027,N_10372);
nor U26595 (N_26595,N_13067,N_10271);
nor U26596 (N_26596,N_16174,N_17551);
nor U26597 (N_26597,N_16009,N_17717);
xnor U26598 (N_26598,N_17098,N_16049);
nor U26599 (N_26599,N_13411,N_16669);
nor U26600 (N_26600,N_11148,N_17973);
nor U26601 (N_26601,N_10387,N_15492);
nor U26602 (N_26602,N_11233,N_13500);
nand U26603 (N_26603,N_12655,N_19247);
xnor U26604 (N_26604,N_10461,N_16361);
nand U26605 (N_26605,N_19107,N_14288);
nor U26606 (N_26606,N_11723,N_15890);
xor U26607 (N_26607,N_11814,N_14315);
or U26608 (N_26608,N_16045,N_18159);
xor U26609 (N_26609,N_15234,N_11945);
nand U26610 (N_26610,N_17002,N_13046);
nand U26611 (N_26611,N_14256,N_14793);
or U26612 (N_26612,N_16010,N_11091);
nor U26613 (N_26613,N_18949,N_18874);
and U26614 (N_26614,N_18553,N_17769);
and U26615 (N_26615,N_11980,N_19698);
or U26616 (N_26616,N_13103,N_13242);
and U26617 (N_26617,N_13356,N_19692);
or U26618 (N_26618,N_15393,N_16977);
xor U26619 (N_26619,N_12778,N_12498);
xnor U26620 (N_26620,N_12140,N_11398);
xnor U26621 (N_26621,N_11078,N_15866);
nor U26622 (N_26622,N_13453,N_14497);
xor U26623 (N_26623,N_10101,N_18072);
xor U26624 (N_26624,N_15457,N_19827);
and U26625 (N_26625,N_14065,N_14494);
nor U26626 (N_26626,N_17790,N_12985);
and U26627 (N_26627,N_11732,N_10119);
xnor U26628 (N_26628,N_13501,N_12979);
nand U26629 (N_26629,N_11697,N_16601);
nor U26630 (N_26630,N_14855,N_10571);
or U26631 (N_26631,N_19207,N_10032);
nand U26632 (N_26632,N_12927,N_19017);
xnor U26633 (N_26633,N_11293,N_16836);
nand U26634 (N_26634,N_18966,N_18666);
xnor U26635 (N_26635,N_13519,N_10232);
xor U26636 (N_26636,N_14494,N_18974);
and U26637 (N_26637,N_12424,N_14258);
nor U26638 (N_26638,N_16218,N_13412);
nor U26639 (N_26639,N_15656,N_19415);
xnor U26640 (N_26640,N_17784,N_14131);
nor U26641 (N_26641,N_18979,N_16260);
nand U26642 (N_26642,N_18161,N_14485);
nand U26643 (N_26643,N_12081,N_16029);
and U26644 (N_26644,N_19834,N_16627);
nand U26645 (N_26645,N_12903,N_16797);
or U26646 (N_26646,N_19112,N_16740);
nand U26647 (N_26647,N_18704,N_13543);
xor U26648 (N_26648,N_15616,N_11214);
or U26649 (N_26649,N_12646,N_19940);
nand U26650 (N_26650,N_16805,N_11462);
xnor U26651 (N_26651,N_10523,N_13927);
xnor U26652 (N_26652,N_13756,N_12561);
nor U26653 (N_26653,N_11704,N_10385);
nand U26654 (N_26654,N_11460,N_12705);
nand U26655 (N_26655,N_17367,N_18404);
xnor U26656 (N_26656,N_13106,N_16589);
or U26657 (N_26657,N_11557,N_11167);
and U26658 (N_26658,N_19398,N_16203);
nand U26659 (N_26659,N_18216,N_16851);
or U26660 (N_26660,N_13674,N_15794);
or U26661 (N_26661,N_19268,N_14859);
xnor U26662 (N_26662,N_14321,N_16614);
or U26663 (N_26663,N_17212,N_11154);
and U26664 (N_26664,N_19574,N_13467);
nor U26665 (N_26665,N_11922,N_19501);
nor U26666 (N_26666,N_17890,N_15683);
xor U26667 (N_26667,N_17576,N_17533);
and U26668 (N_26668,N_18749,N_10698);
xnor U26669 (N_26669,N_17197,N_18500);
and U26670 (N_26670,N_10882,N_13861);
nand U26671 (N_26671,N_12788,N_13999);
or U26672 (N_26672,N_14730,N_12199);
nor U26673 (N_26673,N_14451,N_10781);
and U26674 (N_26674,N_15311,N_12424);
nor U26675 (N_26675,N_19820,N_18585);
xnor U26676 (N_26676,N_16305,N_17313);
nand U26677 (N_26677,N_16718,N_14508);
and U26678 (N_26678,N_17635,N_16894);
nor U26679 (N_26679,N_19043,N_11257);
and U26680 (N_26680,N_10660,N_13563);
nor U26681 (N_26681,N_19657,N_18049);
xor U26682 (N_26682,N_15078,N_10012);
and U26683 (N_26683,N_17257,N_12830);
nand U26684 (N_26684,N_11112,N_13038);
nor U26685 (N_26685,N_11949,N_15033);
and U26686 (N_26686,N_16372,N_18565);
or U26687 (N_26687,N_12029,N_12354);
nor U26688 (N_26688,N_19434,N_15764);
nand U26689 (N_26689,N_13049,N_12414);
and U26690 (N_26690,N_19554,N_17025);
nand U26691 (N_26691,N_14677,N_11315);
nor U26692 (N_26692,N_14477,N_15955);
nand U26693 (N_26693,N_18693,N_16939);
nand U26694 (N_26694,N_17547,N_12410);
xnor U26695 (N_26695,N_12798,N_10998);
nand U26696 (N_26696,N_18983,N_14272);
nand U26697 (N_26697,N_13750,N_15427);
nor U26698 (N_26698,N_10582,N_19593);
and U26699 (N_26699,N_16315,N_10179);
xor U26700 (N_26700,N_10679,N_19469);
or U26701 (N_26701,N_15581,N_11299);
or U26702 (N_26702,N_13863,N_14644);
or U26703 (N_26703,N_19990,N_18874);
nor U26704 (N_26704,N_15038,N_18236);
nand U26705 (N_26705,N_12743,N_16734);
or U26706 (N_26706,N_11980,N_12284);
and U26707 (N_26707,N_18696,N_15143);
nor U26708 (N_26708,N_11406,N_13638);
nand U26709 (N_26709,N_14675,N_10950);
xor U26710 (N_26710,N_19646,N_17441);
and U26711 (N_26711,N_10935,N_19859);
xnor U26712 (N_26712,N_19123,N_18194);
and U26713 (N_26713,N_16602,N_11308);
nor U26714 (N_26714,N_13866,N_10436);
nand U26715 (N_26715,N_17332,N_11414);
xor U26716 (N_26716,N_18380,N_14173);
nor U26717 (N_26717,N_14533,N_18678);
nand U26718 (N_26718,N_12145,N_11699);
and U26719 (N_26719,N_13338,N_11248);
nor U26720 (N_26720,N_17467,N_11641);
nand U26721 (N_26721,N_11133,N_18497);
nor U26722 (N_26722,N_12908,N_10221);
nor U26723 (N_26723,N_11772,N_16955);
nand U26724 (N_26724,N_12490,N_10229);
and U26725 (N_26725,N_13859,N_11053);
and U26726 (N_26726,N_17891,N_17553);
nor U26727 (N_26727,N_14266,N_14410);
xor U26728 (N_26728,N_14761,N_12815);
and U26729 (N_26729,N_11698,N_13172);
and U26730 (N_26730,N_14549,N_18514);
xnor U26731 (N_26731,N_16551,N_10425);
xnor U26732 (N_26732,N_15389,N_11389);
or U26733 (N_26733,N_15739,N_14919);
nand U26734 (N_26734,N_19217,N_11170);
or U26735 (N_26735,N_12597,N_15767);
and U26736 (N_26736,N_18851,N_11451);
nor U26737 (N_26737,N_10330,N_13845);
nand U26738 (N_26738,N_10232,N_10955);
xor U26739 (N_26739,N_19933,N_19464);
xnor U26740 (N_26740,N_15924,N_19037);
or U26741 (N_26741,N_10088,N_18731);
nor U26742 (N_26742,N_19316,N_18470);
nand U26743 (N_26743,N_13185,N_13418);
nor U26744 (N_26744,N_18048,N_15263);
nor U26745 (N_26745,N_13354,N_19641);
or U26746 (N_26746,N_13789,N_14227);
nor U26747 (N_26747,N_18042,N_14933);
and U26748 (N_26748,N_12738,N_13600);
or U26749 (N_26749,N_11426,N_16587);
nand U26750 (N_26750,N_19993,N_12549);
xor U26751 (N_26751,N_18653,N_19784);
or U26752 (N_26752,N_10825,N_15587);
xor U26753 (N_26753,N_12017,N_12244);
and U26754 (N_26754,N_12317,N_18110);
nor U26755 (N_26755,N_11577,N_16234);
nor U26756 (N_26756,N_13200,N_13168);
nand U26757 (N_26757,N_11726,N_17298);
and U26758 (N_26758,N_16678,N_16813);
xnor U26759 (N_26759,N_13629,N_15563);
xnor U26760 (N_26760,N_16692,N_15452);
nor U26761 (N_26761,N_13791,N_13895);
nor U26762 (N_26762,N_16811,N_18323);
xor U26763 (N_26763,N_14982,N_13995);
nor U26764 (N_26764,N_19019,N_14325);
nand U26765 (N_26765,N_10285,N_18184);
nand U26766 (N_26766,N_10661,N_15060);
and U26767 (N_26767,N_15667,N_14666);
and U26768 (N_26768,N_15324,N_17772);
xnor U26769 (N_26769,N_12296,N_17625);
nand U26770 (N_26770,N_18509,N_18566);
nand U26771 (N_26771,N_18972,N_19456);
nor U26772 (N_26772,N_16755,N_13732);
xnor U26773 (N_26773,N_10756,N_16397);
or U26774 (N_26774,N_18633,N_17210);
nand U26775 (N_26775,N_17434,N_16500);
or U26776 (N_26776,N_19404,N_19783);
xor U26777 (N_26777,N_10087,N_18703);
nor U26778 (N_26778,N_17913,N_12478);
nor U26779 (N_26779,N_16658,N_14874);
xnor U26780 (N_26780,N_15631,N_14420);
and U26781 (N_26781,N_13054,N_11674);
nand U26782 (N_26782,N_17020,N_10798);
nor U26783 (N_26783,N_15690,N_18822);
or U26784 (N_26784,N_11883,N_11410);
and U26785 (N_26785,N_18150,N_17353);
or U26786 (N_26786,N_18334,N_10759);
xnor U26787 (N_26787,N_11362,N_15387);
or U26788 (N_26788,N_18329,N_11417);
nand U26789 (N_26789,N_17713,N_16160);
or U26790 (N_26790,N_10443,N_14644);
nor U26791 (N_26791,N_17852,N_17844);
and U26792 (N_26792,N_10105,N_11560);
nand U26793 (N_26793,N_17677,N_16081);
or U26794 (N_26794,N_16059,N_11588);
and U26795 (N_26795,N_13683,N_14500);
or U26796 (N_26796,N_12817,N_13045);
xnor U26797 (N_26797,N_13685,N_10891);
xor U26798 (N_26798,N_11666,N_15177);
nand U26799 (N_26799,N_17115,N_11628);
or U26800 (N_26800,N_19455,N_11019);
or U26801 (N_26801,N_15825,N_14107);
nand U26802 (N_26802,N_11171,N_13144);
nand U26803 (N_26803,N_13012,N_16390);
nor U26804 (N_26804,N_11393,N_17200);
and U26805 (N_26805,N_15608,N_18237);
xnor U26806 (N_26806,N_15998,N_13459);
and U26807 (N_26807,N_16825,N_15586);
nand U26808 (N_26808,N_10723,N_18776);
nor U26809 (N_26809,N_15405,N_15829);
xor U26810 (N_26810,N_10000,N_15128);
nor U26811 (N_26811,N_18264,N_10009);
nand U26812 (N_26812,N_10553,N_14193);
nand U26813 (N_26813,N_15450,N_17073);
and U26814 (N_26814,N_18147,N_16213);
or U26815 (N_26815,N_19168,N_19868);
nand U26816 (N_26816,N_17488,N_19649);
nor U26817 (N_26817,N_18159,N_14942);
xnor U26818 (N_26818,N_16910,N_10135);
xor U26819 (N_26819,N_14053,N_19008);
nor U26820 (N_26820,N_13726,N_11553);
nor U26821 (N_26821,N_16976,N_10772);
or U26822 (N_26822,N_11167,N_10159);
and U26823 (N_26823,N_16843,N_15920);
nand U26824 (N_26824,N_10177,N_11919);
nor U26825 (N_26825,N_17157,N_17459);
or U26826 (N_26826,N_11113,N_13573);
xor U26827 (N_26827,N_15728,N_18058);
or U26828 (N_26828,N_16305,N_19264);
nand U26829 (N_26829,N_10723,N_13166);
or U26830 (N_26830,N_12490,N_11551);
xnor U26831 (N_26831,N_18141,N_11539);
or U26832 (N_26832,N_16465,N_17478);
and U26833 (N_26833,N_18317,N_19706);
and U26834 (N_26834,N_11401,N_12961);
nor U26835 (N_26835,N_10479,N_13894);
xnor U26836 (N_26836,N_15091,N_16918);
nor U26837 (N_26837,N_13385,N_12706);
nand U26838 (N_26838,N_17002,N_19013);
nor U26839 (N_26839,N_19593,N_15329);
and U26840 (N_26840,N_15047,N_12613);
xor U26841 (N_26841,N_10416,N_14617);
nor U26842 (N_26842,N_12397,N_11130);
nand U26843 (N_26843,N_11456,N_12581);
nor U26844 (N_26844,N_17651,N_10001);
nand U26845 (N_26845,N_17794,N_11564);
nor U26846 (N_26846,N_17324,N_17735);
or U26847 (N_26847,N_13106,N_16263);
xnor U26848 (N_26848,N_11454,N_11455);
nor U26849 (N_26849,N_14116,N_14576);
and U26850 (N_26850,N_12699,N_11288);
and U26851 (N_26851,N_14989,N_17524);
or U26852 (N_26852,N_19773,N_18084);
nor U26853 (N_26853,N_16958,N_11311);
nand U26854 (N_26854,N_13996,N_16517);
nand U26855 (N_26855,N_13004,N_16797);
nand U26856 (N_26856,N_17740,N_17484);
or U26857 (N_26857,N_11526,N_15587);
or U26858 (N_26858,N_13269,N_17856);
and U26859 (N_26859,N_17296,N_14202);
nand U26860 (N_26860,N_10807,N_12409);
and U26861 (N_26861,N_15576,N_13408);
xnor U26862 (N_26862,N_16572,N_11994);
and U26863 (N_26863,N_11343,N_17715);
and U26864 (N_26864,N_14213,N_16394);
xnor U26865 (N_26865,N_15185,N_15750);
nand U26866 (N_26866,N_12952,N_19110);
nand U26867 (N_26867,N_12677,N_14084);
nor U26868 (N_26868,N_16632,N_19400);
nand U26869 (N_26869,N_14825,N_14123);
xnor U26870 (N_26870,N_11708,N_17617);
xnor U26871 (N_26871,N_16587,N_18942);
xnor U26872 (N_26872,N_14972,N_10398);
and U26873 (N_26873,N_11023,N_18554);
or U26874 (N_26874,N_14235,N_15027);
or U26875 (N_26875,N_16436,N_17995);
or U26876 (N_26876,N_18831,N_17658);
and U26877 (N_26877,N_16927,N_19972);
or U26878 (N_26878,N_10424,N_13646);
nand U26879 (N_26879,N_14780,N_15326);
xnor U26880 (N_26880,N_19123,N_12558);
or U26881 (N_26881,N_11327,N_17739);
nand U26882 (N_26882,N_11131,N_15201);
and U26883 (N_26883,N_18104,N_12084);
nor U26884 (N_26884,N_17998,N_19501);
or U26885 (N_26885,N_17677,N_18491);
or U26886 (N_26886,N_14597,N_19478);
nor U26887 (N_26887,N_11939,N_19537);
and U26888 (N_26888,N_14139,N_10776);
nor U26889 (N_26889,N_11120,N_14141);
nand U26890 (N_26890,N_13094,N_13654);
and U26891 (N_26891,N_15647,N_15641);
nor U26892 (N_26892,N_18847,N_14946);
and U26893 (N_26893,N_13947,N_13885);
and U26894 (N_26894,N_11166,N_18150);
nand U26895 (N_26895,N_10579,N_17060);
xor U26896 (N_26896,N_16771,N_19521);
nor U26897 (N_26897,N_10577,N_18963);
nand U26898 (N_26898,N_10287,N_14434);
xnor U26899 (N_26899,N_18298,N_17458);
xnor U26900 (N_26900,N_15213,N_16546);
and U26901 (N_26901,N_14179,N_19453);
xor U26902 (N_26902,N_14513,N_19730);
or U26903 (N_26903,N_19183,N_11524);
nor U26904 (N_26904,N_14871,N_15542);
or U26905 (N_26905,N_15771,N_13711);
xnor U26906 (N_26906,N_12414,N_14290);
nor U26907 (N_26907,N_12037,N_15157);
and U26908 (N_26908,N_19636,N_16344);
nor U26909 (N_26909,N_11386,N_10959);
and U26910 (N_26910,N_17538,N_16251);
and U26911 (N_26911,N_15405,N_17241);
nand U26912 (N_26912,N_13297,N_13021);
xnor U26913 (N_26913,N_11467,N_12194);
nor U26914 (N_26914,N_18610,N_15442);
nor U26915 (N_26915,N_18292,N_13077);
and U26916 (N_26916,N_17231,N_16548);
xor U26917 (N_26917,N_13023,N_19249);
xnor U26918 (N_26918,N_13874,N_17549);
and U26919 (N_26919,N_11181,N_17080);
nor U26920 (N_26920,N_12398,N_11040);
nor U26921 (N_26921,N_17771,N_13357);
nand U26922 (N_26922,N_10470,N_16832);
nand U26923 (N_26923,N_12487,N_14379);
or U26924 (N_26924,N_10878,N_10009);
nor U26925 (N_26925,N_10271,N_16663);
xor U26926 (N_26926,N_15052,N_11391);
nand U26927 (N_26927,N_14421,N_15281);
and U26928 (N_26928,N_14401,N_14498);
or U26929 (N_26929,N_10196,N_15989);
xor U26930 (N_26930,N_13483,N_11675);
nand U26931 (N_26931,N_15531,N_11374);
xnor U26932 (N_26932,N_17485,N_18109);
or U26933 (N_26933,N_11939,N_13352);
nor U26934 (N_26934,N_17821,N_15720);
or U26935 (N_26935,N_11938,N_16500);
nand U26936 (N_26936,N_16130,N_19241);
xnor U26937 (N_26937,N_14103,N_10882);
nor U26938 (N_26938,N_19450,N_19820);
or U26939 (N_26939,N_15874,N_10181);
nand U26940 (N_26940,N_19942,N_17621);
and U26941 (N_26941,N_10976,N_11332);
nand U26942 (N_26942,N_16015,N_18084);
nand U26943 (N_26943,N_17325,N_10113);
xor U26944 (N_26944,N_18864,N_18071);
and U26945 (N_26945,N_17642,N_18853);
and U26946 (N_26946,N_12149,N_17203);
and U26947 (N_26947,N_16237,N_17122);
nor U26948 (N_26948,N_12813,N_14277);
nor U26949 (N_26949,N_16421,N_10654);
xor U26950 (N_26950,N_19596,N_14684);
and U26951 (N_26951,N_16972,N_13157);
nand U26952 (N_26952,N_19047,N_19995);
xnor U26953 (N_26953,N_14563,N_14570);
nand U26954 (N_26954,N_11029,N_19014);
and U26955 (N_26955,N_18655,N_18353);
nor U26956 (N_26956,N_11258,N_19583);
and U26957 (N_26957,N_16529,N_14669);
or U26958 (N_26958,N_17666,N_15284);
nand U26959 (N_26959,N_11803,N_18437);
nor U26960 (N_26960,N_18284,N_17986);
or U26961 (N_26961,N_12159,N_13349);
xor U26962 (N_26962,N_19799,N_16084);
nor U26963 (N_26963,N_16086,N_10482);
nand U26964 (N_26964,N_17252,N_16114);
xor U26965 (N_26965,N_14880,N_14777);
nand U26966 (N_26966,N_14433,N_14340);
nand U26967 (N_26967,N_13824,N_16111);
or U26968 (N_26968,N_12728,N_11664);
nand U26969 (N_26969,N_17886,N_15951);
and U26970 (N_26970,N_18382,N_15358);
and U26971 (N_26971,N_16522,N_16462);
xnor U26972 (N_26972,N_17919,N_15680);
nor U26973 (N_26973,N_13517,N_16090);
xnor U26974 (N_26974,N_14681,N_10692);
xor U26975 (N_26975,N_15908,N_10343);
or U26976 (N_26976,N_12062,N_12173);
nand U26977 (N_26977,N_19580,N_10083);
nor U26978 (N_26978,N_15424,N_18640);
xnor U26979 (N_26979,N_14791,N_18753);
nand U26980 (N_26980,N_15040,N_19044);
and U26981 (N_26981,N_16473,N_17796);
xor U26982 (N_26982,N_18541,N_18248);
nand U26983 (N_26983,N_18199,N_12074);
nor U26984 (N_26984,N_12634,N_11449);
nor U26985 (N_26985,N_17408,N_14706);
and U26986 (N_26986,N_15822,N_15096);
nand U26987 (N_26987,N_15907,N_15810);
xnor U26988 (N_26988,N_13771,N_14345);
nor U26989 (N_26989,N_12964,N_18117);
nand U26990 (N_26990,N_16522,N_19490);
nand U26991 (N_26991,N_11551,N_11738);
xnor U26992 (N_26992,N_13123,N_12497);
xnor U26993 (N_26993,N_17158,N_11665);
or U26994 (N_26994,N_12413,N_16503);
nand U26995 (N_26995,N_10173,N_13904);
nand U26996 (N_26996,N_14507,N_19131);
and U26997 (N_26997,N_18639,N_19482);
and U26998 (N_26998,N_16334,N_11710);
or U26999 (N_26999,N_14849,N_17035);
or U27000 (N_27000,N_19860,N_12571);
nand U27001 (N_27001,N_17858,N_11153);
xnor U27002 (N_27002,N_15966,N_11261);
xor U27003 (N_27003,N_17602,N_18141);
xnor U27004 (N_27004,N_11083,N_16060);
xnor U27005 (N_27005,N_16327,N_11080);
nand U27006 (N_27006,N_18580,N_17783);
xor U27007 (N_27007,N_17390,N_14006);
and U27008 (N_27008,N_15200,N_18666);
nand U27009 (N_27009,N_13145,N_12537);
nand U27010 (N_27010,N_16406,N_17543);
nor U27011 (N_27011,N_18221,N_16622);
nor U27012 (N_27012,N_12536,N_12057);
or U27013 (N_27013,N_12582,N_19483);
and U27014 (N_27014,N_13145,N_10663);
nand U27015 (N_27015,N_10503,N_11440);
nand U27016 (N_27016,N_11698,N_10122);
or U27017 (N_27017,N_19471,N_14218);
and U27018 (N_27018,N_17697,N_17439);
nor U27019 (N_27019,N_15313,N_13775);
nand U27020 (N_27020,N_17220,N_16894);
nand U27021 (N_27021,N_18986,N_19299);
and U27022 (N_27022,N_18443,N_10577);
or U27023 (N_27023,N_11416,N_12465);
nand U27024 (N_27024,N_11796,N_10559);
and U27025 (N_27025,N_16388,N_19834);
and U27026 (N_27026,N_11938,N_13283);
xnor U27027 (N_27027,N_13189,N_19947);
or U27028 (N_27028,N_15057,N_12965);
nand U27029 (N_27029,N_15032,N_16897);
nor U27030 (N_27030,N_18764,N_19258);
xor U27031 (N_27031,N_10833,N_12780);
xor U27032 (N_27032,N_12446,N_13759);
nor U27033 (N_27033,N_12369,N_12180);
nand U27034 (N_27034,N_17197,N_17116);
nor U27035 (N_27035,N_16529,N_16756);
xor U27036 (N_27036,N_18581,N_13036);
xor U27037 (N_27037,N_11273,N_12600);
nand U27038 (N_27038,N_13353,N_18790);
xor U27039 (N_27039,N_11887,N_12924);
or U27040 (N_27040,N_17132,N_14866);
nand U27041 (N_27041,N_16627,N_15834);
or U27042 (N_27042,N_19010,N_16537);
xnor U27043 (N_27043,N_16218,N_19387);
nor U27044 (N_27044,N_19614,N_11722);
or U27045 (N_27045,N_15431,N_13267);
nand U27046 (N_27046,N_10393,N_15742);
or U27047 (N_27047,N_17949,N_17389);
nor U27048 (N_27048,N_18819,N_19583);
nor U27049 (N_27049,N_12305,N_17515);
xor U27050 (N_27050,N_19105,N_19586);
xnor U27051 (N_27051,N_18224,N_18809);
xnor U27052 (N_27052,N_18583,N_16825);
nand U27053 (N_27053,N_12697,N_19789);
nand U27054 (N_27054,N_14036,N_12542);
and U27055 (N_27055,N_19844,N_15548);
and U27056 (N_27056,N_19572,N_17610);
nand U27057 (N_27057,N_12237,N_14806);
xnor U27058 (N_27058,N_17134,N_15201);
nor U27059 (N_27059,N_10097,N_12793);
xor U27060 (N_27060,N_11221,N_12220);
or U27061 (N_27061,N_17405,N_15370);
and U27062 (N_27062,N_19228,N_15216);
and U27063 (N_27063,N_13840,N_12230);
nand U27064 (N_27064,N_10240,N_11432);
nand U27065 (N_27065,N_18679,N_13848);
or U27066 (N_27066,N_18381,N_13709);
nor U27067 (N_27067,N_12667,N_18305);
nand U27068 (N_27068,N_18306,N_19112);
xnor U27069 (N_27069,N_15588,N_18380);
and U27070 (N_27070,N_11692,N_16736);
nor U27071 (N_27071,N_14701,N_10629);
and U27072 (N_27072,N_18661,N_10422);
nand U27073 (N_27073,N_14973,N_13549);
nor U27074 (N_27074,N_17652,N_17309);
nor U27075 (N_27075,N_19537,N_16906);
nor U27076 (N_27076,N_16029,N_17336);
and U27077 (N_27077,N_16155,N_19411);
xnor U27078 (N_27078,N_12847,N_13434);
and U27079 (N_27079,N_19885,N_14905);
and U27080 (N_27080,N_19678,N_17121);
or U27081 (N_27081,N_10303,N_15136);
and U27082 (N_27082,N_16362,N_19851);
nand U27083 (N_27083,N_18315,N_12529);
xor U27084 (N_27084,N_13653,N_13669);
and U27085 (N_27085,N_15174,N_17200);
or U27086 (N_27086,N_11080,N_16038);
and U27087 (N_27087,N_17682,N_14735);
xor U27088 (N_27088,N_15835,N_18040);
nor U27089 (N_27089,N_16856,N_15491);
nor U27090 (N_27090,N_19995,N_15853);
nor U27091 (N_27091,N_19574,N_17189);
and U27092 (N_27092,N_10232,N_18914);
and U27093 (N_27093,N_15666,N_16178);
nor U27094 (N_27094,N_15413,N_12591);
xor U27095 (N_27095,N_15729,N_13075);
or U27096 (N_27096,N_16985,N_14541);
nand U27097 (N_27097,N_18450,N_16746);
nand U27098 (N_27098,N_12907,N_13690);
nand U27099 (N_27099,N_15825,N_10320);
or U27100 (N_27100,N_12028,N_12282);
or U27101 (N_27101,N_11944,N_10304);
xnor U27102 (N_27102,N_14171,N_10173);
nor U27103 (N_27103,N_11347,N_15386);
nor U27104 (N_27104,N_16313,N_18063);
nand U27105 (N_27105,N_10627,N_19715);
or U27106 (N_27106,N_10505,N_10361);
or U27107 (N_27107,N_16906,N_17668);
xnor U27108 (N_27108,N_12911,N_11833);
xor U27109 (N_27109,N_14499,N_16640);
nor U27110 (N_27110,N_19026,N_17017);
nand U27111 (N_27111,N_14542,N_11503);
nor U27112 (N_27112,N_17912,N_19372);
and U27113 (N_27113,N_13602,N_11779);
and U27114 (N_27114,N_16694,N_16410);
xnor U27115 (N_27115,N_19484,N_12595);
nand U27116 (N_27116,N_18298,N_11962);
nor U27117 (N_27117,N_11514,N_10030);
and U27118 (N_27118,N_13048,N_10678);
nand U27119 (N_27119,N_15164,N_15063);
nor U27120 (N_27120,N_13414,N_18383);
and U27121 (N_27121,N_19796,N_15559);
and U27122 (N_27122,N_14838,N_17352);
nor U27123 (N_27123,N_11636,N_10346);
nand U27124 (N_27124,N_16013,N_11311);
or U27125 (N_27125,N_14851,N_17242);
nand U27126 (N_27126,N_12455,N_10156);
xnor U27127 (N_27127,N_15803,N_10756);
nor U27128 (N_27128,N_15163,N_17597);
and U27129 (N_27129,N_17467,N_12437);
and U27130 (N_27130,N_13680,N_15290);
or U27131 (N_27131,N_19900,N_13820);
nor U27132 (N_27132,N_17132,N_17551);
or U27133 (N_27133,N_15415,N_16255);
xnor U27134 (N_27134,N_14520,N_18871);
nor U27135 (N_27135,N_19478,N_11527);
nand U27136 (N_27136,N_12730,N_12930);
or U27137 (N_27137,N_10769,N_18070);
nor U27138 (N_27138,N_19373,N_12356);
nand U27139 (N_27139,N_19412,N_13826);
xor U27140 (N_27140,N_11109,N_19521);
xnor U27141 (N_27141,N_19165,N_10737);
xor U27142 (N_27142,N_13282,N_11857);
nor U27143 (N_27143,N_13475,N_17794);
nand U27144 (N_27144,N_11446,N_17504);
and U27145 (N_27145,N_12600,N_16924);
or U27146 (N_27146,N_18547,N_19298);
xnor U27147 (N_27147,N_12830,N_13942);
nand U27148 (N_27148,N_16483,N_16309);
nand U27149 (N_27149,N_10851,N_13331);
nand U27150 (N_27150,N_10858,N_15369);
xor U27151 (N_27151,N_17641,N_14946);
or U27152 (N_27152,N_14965,N_19174);
xor U27153 (N_27153,N_15469,N_13715);
or U27154 (N_27154,N_18699,N_14959);
or U27155 (N_27155,N_19417,N_19882);
nand U27156 (N_27156,N_14680,N_13070);
and U27157 (N_27157,N_19014,N_17650);
nor U27158 (N_27158,N_15288,N_17656);
and U27159 (N_27159,N_14845,N_17142);
xor U27160 (N_27160,N_16149,N_19450);
xnor U27161 (N_27161,N_13141,N_13049);
and U27162 (N_27162,N_16820,N_16510);
or U27163 (N_27163,N_15210,N_18115);
nand U27164 (N_27164,N_13641,N_15066);
nand U27165 (N_27165,N_13120,N_12503);
nand U27166 (N_27166,N_10213,N_11519);
nor U27167 (N_27167,N_11056,N_12756);
or U27168 (N_27168,N_19739,N_11543);
nor U27169 (N_27169,N_14519,N_12460);
or U27170 (N_27170,N_15243,N_18346);
nor U27171 (N_27171,N_13626,N_16063);
and U27172 (N_27172,N_10508,N_13585);
nor U27173 (N_27173,N_16479,N_12204);
nor U27174 (N_27174,N_16681,N_19757);
nor U27175 (N_27175,N_12424,N_17140);
nor U27176 (N_27176,N_11453,N_13749);
nor U27177 (N_27177,N_13704,N_15239);
and U27178 (N_27178,N_18803,N_15869);
or U27179 (N_27179,N_11070,N_11939);
or U27180 (N_27180,N_15314,N_15523);
xnor U27181 (N_27181,N_17591,N_14274);
nand U27182 (N_27182,N_17824,N_10769);
nor U27183 (N_27183,N_19836,N_10854);
nand U27184 (N_27184,N_13100,N_10350);
nor U27185 (N_27185,N_10095,N_11332);
and U27186 (N_27186,N_17106,N_16507);
xnor U27187 (N_27187,N_10404,N_17112);
or U27188 (N_27188,N_19641,N_18696);
and U27189 (N_27189,N_14647,N_11310);
nor U27190 (N_27190,N_19144,N_17475);
nand U27191 (N_27191,N_18386,N_13389);
or U27192 (N_27192,N_17585,N_17232);
nand U27193 (N_27193,N_12230,N_10196);
nor U27194 (N_27194,N_10828,N_15219);
nor U27195 (N_27195,N_15134,N_16279);
and U27196 (N_27196,N_10686,N_11418);
or U27197 (N_27197,N_11741,N_15812);
and U27198 (N_27198,N_12609,N_14188);
and U27199 (N_27199,N_18153,N_16766);
xor U27200 (N_27200,N_18902,N_19162);
and U27201 (N_27201,N_11060,N_17991);
and U27202 (N_27202,N_17013,N_10587);
nor U27203 (N_27203,N_16529,N_13213);
nor U27204 (N_27204,N_19595,N_16762);
nand U27205 (N_27205,N_12007,N_17576);
and U27206 (N_27206,N_17340,N_14749);
xor U27207 (N_27207,N_17358,N_18439);
and U27208 (N_27208,N_16698,N_18084);
nand U27209 (N_27209,N_17152,N_11714);
nor U27210 (N_27210,N_17882,N_15719);
nor U27211 (N_27211,N_11705,N_10327);
nand U27212 (N_27212,N_10740,N_13978);
nand U27213 (N_27213,N_12723,N_14927);
or U27214 (N_27214,N_15776,N_11774);
or U27215 (N_27215,N_16069,N_18103);
nor U27216 (N_27216,N_11882,N_15560);
and U27217 (N_27217,N_17060,N_19790);
or U27218 (N_27218,N_11276,N_11348);
or U27219 (N_27219,N_17880,N_17137);
nor U27220 (N_27220,N_13983,N_14751);
and U27221 (N_27221,N_19751,N_13668);
and U27222 (N_27222,N_13136,N_11291);
xor U27223 (N_27223,N_16146,N_10558);
nor U27224 (N_27224,N_13208,N_13241);
xor U27225 (N_27225,N_16674,N_14490);
xor U27226 (N_27226,N_19041,N_18573);
and U27227 (N_27227,N_18987,N_15703);
xnor U27228 (N_27228,N_13281,N_12504);
nand U27229 (N_27229,N_15385,N_18548);
xor U27230 (N_27230,N_13827,N_11750);
nand U27231 (N_27231,N_10952,N_10055);
and U27232 (N_27232,N_10613,N_16045);
nor U27233 (N_27233,N_11777,N_11333);
and U27234 (N_27234,N_12930,N_10840);
nand U27235 (N_27235,N_12389,N_18036);
or U27236 (N_27236,N_17191,N_14703);
nor U27237 (N_27237,N_13241,N_14197);
nand U27238 (N_27238,N_16239,N_11093);
or U27239 (N_27239,N_15568,N_18256);
nand U27240 (N_27240,N_17010,N_17480);
xnor U27241 (N_27241,N_15474,N_11703);
xor U27242 (N_27242,N_14182,N_17321);
nor U27243 (N_27243,N_13031,N_13427);
and U27244 (N_27244,N_18151,N_17069);
nand U27245 (N_27245,N_18510,N_16957);
nand U27246 (N_27246,N_12293,N_17631);
or U27247 (N_27247,N_19255,N_10213);
and U27248 (N_27248,N_17726,N_13344);
nor U27249 (N_27249,N_19209,N_16222);
and U27250 (N_27250,N_16571,N_14171);
xor U27251 (N_27251,N_10168,N_10465);
and U27252 (N_27252,N_14285,N_16838);
nor U27253 (N_27253,N_15412,N_12617);
xor U27254 (N_27254,N_17784,N_14316);
nor U27255 (N_27255,N_14345,N_17176);
and U27256 (N_27256,N_12030,N_17090);
or U27257 (N_27257,N_10761,N_17038);
xnor U27258 (N_27258,N_12027,N_15327);
nand U27259 (N_27259,N_17084,N_14020);
nor U27260 (N_27260,N_14577,N_14413);
and U27261 (N_27261,N_19265,N_14139);
xnor U27262 (N_27262,N_12267,N_15290);
nor U27263 (N_27263,N_16407,N_16721);
nand U27264 (N_27264,N_10114,N_16204);
xnor U27265 (N_27265,N_11929,N_13829);
and U27266 (N_27266,N_14537,N_19775);
and U27267 (N_27267,N_12254,N_17436);
or U27268 (N_27268,N_16065,N_18945);
and U27269 (N_27269,N_10632,N_16486);
xnor U27270 (N_27270,N_12563,N_10313);
nand U27271 (N_27271,N_16696,N_14833);
and U27272 (N_27272,N_19393,N_11018);
and U27273 (N_27273,N_15165,N_11418);
xnor U27274 (N_27274,N_19507,N_18833);
and U27275 (N_27275,N_17346,N_17442);
nor U27276 (N_27276,N_14177,N_12724);
xnor U27277 (N_27277,N_11771,N_15721);
nand U27278 (N_27278,N_16992,N_17038);
nor U27279 (N_27279,N_18144,N_12247);
and U27280 (N_27280,N_12158,N_11477);
and U27281 (N_27281,N_10962,N_15234);
nor U27282 (N_27282,N_18020,N_15925);
xor U27283 (N_27283,N_16518,N_19357);
or U27284 (N_27284,N_15389,N_10980);
and U27285 (N_27285,N_19479,N_16305);
nor U27286 (N_27286,N_15471,N_13273);
and U27287 (N_27287,N_18921,N_17938);
and U27288 (N_27288,N_10341,N_13778);
and U27289 (N_27289,N_16430,N_19662);
xnor U27290 (N_27290,N_10434,N_13072);
nor U27291 (N_27291,N_19921,N_19146);
and U27292 (N_27292,N_18507,N_16727);
nor U27293 (N_27293,N_18379,N_13087);
or U27294 (N_27294,N_13841,N_11226);
and U27295 (N_27295,N_16659,N_14008);
nor U27296 (N_27296,N_10424,N_11093);
nand U27297 (N_27297,N_15177,N_16054);
or U27298 (N_27298,N_10226,N_12136);
and U27299 (N_27299,N_19141,N_17965);
xnor U27300 (N_27300,N_13297,N_19262);
nor U27301 (N_27301,N_10538,N_17420);
or U27302 (N_27302,N_16604,N_14340);
xor U27303 (N_27303,N_18954,N_12643);
xnor U27304 (N_27304,N_11804,N_18627);
or U27305 (N_27305,N_12162,N_19351);
nor U27306 (N_27306,N_11039,N_12182);
and U27307 (N_27307,N_13841,N_16998);
xor U27308 (N_27308,N_11989,N_10192);
xnor U27309 (N_27309,N_15151,N_10674);
and U27310 (N_27310,N_16251,N_13279);
or U27311 (N_27311,N_18481,N_16152);
xor U27312 (N_27312,N_18141,N_14806);
nor U27313 (N_27313,N_11558,N_16825);
and U27314 (N_27314,N_19548,N_17934);
xnor U27315 (N_27315,N_14823,N_15614);
nor U27316 (N_27316,N_17905,N_19947);
and U27317 (N_27317,N_11461,N_11289);
nor U27318 (N_27318,N_13485,N_16257);
xnor U27319 (N_27319,N_18578,N_17442);
nor U27320 (N_27320,N_14330,N_14110);
xor U27321 (N_27321,N_11158,N_11103);
nor U27322 (N_27322,N_16496,N_14313);
and U27323 (N_27323,N_12431,N_13101);
and U27324 (N_27324,N_17911,N_14336);
and U27325 (N_27325,N_16619,N_19889);
xor U27326 (N_27326,N_18988,N_14491);
or U27327 (N_27327,N_19562,N_12857);
or U27328 (N_27328,N_13003,N_14807);
and U27329 (N_27329,N_12330,N_14186);
nor U27330 (N_27330,N_15024,N_18022);
nor U27331 (N_27331,N_13572,N_14485);
xor U27332 (N_27332,N_19780,N_18540);
nor U27333 (N_27333,N_11877,N_17906);
and U27334 (N_27334,N_10091,N_18301);
nor U27335 (N_27335,N_10191,N_19794);
nor U27336 (N_27336,N_15504,N_14282);
nor U27337 (N_27337,N_14460,N_15087);
or U27338 (N_27338,N_17570,N_15792);
xor U27339 (N_27339,N_19587,N_12895);
nand U27340 (N_27340,N_12239,N_14621);
xor U27341 (N_27341,N_18275,N_12673);
and U27342 (N_27342,N_14899,N_19363);
nand U27343 (N_27343,N_14797,N_19208);
or U27344 (N_27344,N_18791,N_10305);
nor U27345 (N_27345,N_12787,N_19248);
and U27346 (N_27346,N_14571,N_16785);
or U27347 (N_27347,N_12218,N_12882);
or U27348 (N_27348,N_10378,N_13089);
or U27349 (N_27349,N_15545,N_19769);
nor U27350 (N_27350,N_18725,N_10021);
xor U27351 (N_27351,N_19959,N_10358);
or U27352 (N_27352,N_19940,N_19197);
nor U27353 (N_27353,N_16947,N_17148);
and U27354 (N_27354,N_15129,N_14078);
or U27355 (N_27355,N_12175,N_14718);
nand U27356 (N_27356,N_18636,N_16795);
and U27357 (N_27357,N_12615,N_11845);
nor U27358 (N_27358,N_19337,N_12696);
xor U27359 (N_27359,N_14871,N_10238);
and U27360 (N_27360,N_13674,N_15254);
or U27361 (N_27361,N_10155,N_15996);
nand U27362 (N_27362,N_15176,N_19461);
nand U27363 (N_27363,N_17297,N_13332);
or U27364 (N_27364,N_14271,N_18931);
nand U27365 (N_27365,N_14204,N_10939);
nor U27366 (N_27366,N_10087,N_18377);
and U27367 (N_27367,N_15071,N_15634);
and U27368 (N_27368,N_15915,N_11462);
nand U27369 (N_27369,N_13159,N_15929);
xnor U27370 (N_27370,N_12759,N_16366);
nor U27371 (N_27371,N_16832,N_19059);
nand U27372 (N_27372,N_10060,N_12164);
or U27373 (N_27373,N_17254,N_15750);
and U27374 (N_27374,N_17537,N_19680);
xnor U27375 (N_27375,N_15917,N_14238);
nand U27376 (N_27376,N_15388,N_14130);
or U27377 (N_27377,N_19878,N_19269);
nor U27378 (N_27378,N_19507,N_10285);
nand U27379 (N_27379,N_10123,N_15771);
and U27380 (N_27380,N_18503,N_17144);
or U27381 (N_27381,N_10677,N_13390);
and U27382 (N_27382,N_18142,N_19764);
nand U27383 (N_27383,N_18672,N_10535);
nand U27384 (N_27384,N_18215,N_13848);
nor U27385 (N_27385,N_16585,N_14060);
and U27386 (N_27386,N_17072,N_16585);
nor U27387 (N_27387,N_19317,N_12958);
nand U27388 (N_27388,N_11176,N_15811);
and U27389 (N_27389,N_11643,N_12464);
nor U27390 (N_27390,N_14097,N_13430);
and U27391 (N_27391,N_16171,N_19317);
xor U27392 (N_27392,N_16516,N_17436);
nor U27393 (N_27393,N_10883,N_12643);
nor U27394 (N_27394,N_17784,N_14618);
and U27395 (N_27395,N_12191,N_18598);
nand U27396 (N_27396,N_14989,N_17237);
xnor U27397 (N_27397,N_13055,N_19104);
or U27398 (N_27398,N_13632,N_14492);
nand U27399 (N_27399,N_16995,N_19082);
nand U27400 (N_27400,N_16130,N_15420);
nand U27401 (N_27401,N_12220,N_19997);
nor U27402 (N_27402,N_14253,N_14379);
nand U27403 (N_27403,N_17353,N_16727);
or U27404 (N_27404,N_18750,N_17806);
xor U27405 (N_27405,N_11384,N_10898);
or U27406 (N_27406,N_17278,N_12392);
xor U27407 (N_27407,N_10087,N_11954);
and U27408 (N_27408,N_11559,N_16591);
nor U27409 (N_27409,N_10299,N_11023);
nand U27410 (N_27410,N_15732,N_18666);
nand U27411 (N_27411,N_10212,N_14972);
nand U27412 (N_27412,N_16905,N_10360);
xnor U27413 (N_27413,N_10997,N_14062);
xnor U27414 (N_27414,N_13398,N_14565);
xnor U27415 (N_27415,N_13278,N_12975);
or U27416 (N_27416,N_12441,N_18388);
xor U27417 (N_27417,N_11447,N_18228);
or U27418 (N_27418,N_10679,N_10304);
nand U27419 (N_27419,N_10348,N_19905);
and U27420 (N_27420,N_12295,N_16814);
xnor U27421 (N_27421,N_15017,N_16426);
and U27422 (N_27422,N_15356,N_13567);
and U27423 (N_27423,N_15633,N_19739);
xnor U27424 (N_27424,N_10093,N_10258);
and U27425 (N_27425,N_19649,N_19717);
or U27426 (N_27426,N_15035,N_18324);
or U27427 (N_27427,N_14626,N_10519);
nand U27428 (N_27428,N_16658,N_18459);
nor U27429 (N_27429,N_14066,N_11459);
nand U27430 (N_27430,N_18420,N_14566);
or U27431 (N_27431,N_12314,N_19827);
nor U27432 (N_27432,N_14201,N_15977);
nand U27433 (N_27433,N_12285,N_10498);
and U27434 (N_27434,N_14361,N_10239);
nor U27435 (N_27435,N_14883,N_11344);
xnor U27436 (N_27436,N_11116,N_13769);
nand U27437 (N_27437,N_10354,N_10925);
and U27438 (N_27438,N_13448,N_10713);
and U27439 (N_27439,N_13162,N_15022);
nor U27440 (N_27440,N_16291,N_13153);
and U27441 (N_27441,N_17309,N_10931);
nand U27442 (N_27442,N_10453,N_12450);
or U27443 (N_27443,N_13542,N_18322);
xnor U27444 (N_27444,N_15503,N_13926);
nand U27445 (N_27445,N_18025,N_12346);
or U27446 (N_27446,N_17716,N_14011);
nand U27447 (N_27447,N_10664,N_11218);
nor U27448 (N_27448,N_18966,N_12250);
nor U27449 (N_27449,N_11753,N_16486);
nor U27450 (N_27450,N_11678,N_11607);
or U27451 (N_27451,N_19326,N_15936);
and U27452 (N_27452,N_10557,N_10848);
nand U27453 (N_27453,N_12684,N_15762);
nand U27454 (N_27454,N_19375,N_15184);
nor U27455 (N_27455,N_12979,N_11349);
or U27456 (N_27456,N_15791,N_10359);
xnor U27457 (N_27457,N_13129,N_17035);
and U27458 (N_27458,N_17679,N_19509);
or U27459 (N_27459,N_18796,N_14398);
nor U27460 (N_27460,N_11918,N_11079);
or U27461 (N_27461,N_13886,N_10994);
nor U27462 (N_27462,N_14557,N_15665);
nor U27463 (N_27463,N_16090,N_18139);
nand U27464 (N_27464,N_11473,N_12484);
nand U27465 (N_27465,N_15222,N_19320);
or U27466 (N_27466,N_14655,N_10320);
or U27467 (N_27467,N_19108,N_19504);
nand U27468 (N_27468,N_19845,N_10974);
nand U27469 (N_27469,N_18726,N_14203);
and U27470 (N_27470,N_19817,N_11418);
xnor U27471 (N_27471,N_16293,N_13463);
nor U27472 (N_27472,N_17266,N_14546);
or U27473 (N_27473,N_17219,N_16352);
or U27474 (N_27474,N_18958,N_15358);
nand U27475 (N_27475,N_19234,N_16411);
and U27476 (N_27476,N_11681,N_19998);
or U27477 (N_27477,N_13593,N_10215);
nand U27478 (N_27478,N_16856,N_19211);
nor U27479 (N_27479,N_19747,N_10635);
or U27480 (N_27480,N_10389,N_13641);
nand U27481 (N_27481,N_11873,N_12052);
nand U27482 (N_27482,N_10219,N_19000);
nand U27483 (N_27483,N_14251,N_11891);
nand U27484 (N_27484,N_13984,N_19095);
nand U27485 (N_27485,N_11172,N_11497);
nor U27486 (N_27486,N_14592,N_15126);
or U27487 (N_27487,N_10619,N_19325);
and U27488 (N_27488,N_19369,N_19718);
xor U27489 (N_27489,N_18337,N_12208);
xor U27490 (N_27490,N_12405,N_10586);
nor U27491 (N_27491,N_16265,N_12685);
and U27492 (N_27492,N_11176,N_18926);
nand U27493 (N_27493,N_17296,N_19290);
xnor U27494 (N_27494,N_11881,N_11343);
nor U27495 (N_27495,N_18971,N_13139);
nand U27496 (N_27496,N_11328,N_19229);
nand U27497 (N_27497,N_11913,N_10335);
and U27498 (N_27498,N_19545,N_18205);
xnor U27499 (N_27499,N_11401,N_14076);
nor U27500 (N_27500,N_10263,N_15099);
or U27501 (N_27501,N_16069,N_17337);
xnor U27502 (N_27502,N_12619,N_14280);
and U27503 (N_27503,N_17449,N_14190);
xor U27504 (N_27504,N_15925,N_14457);
xnor U27505 (N_27505,N_18517,N_19987);
nor U27506 (N_27506,N_17172,N_17348);
nand U27507 (N_27507,N_13347,N_16270);
nor U27508 (N_27508,N_11601,N_13376);
nor U27509 (N_27509,N_11132,N_14291);
xor U27510 (N_27510,N_11528,N_17239);
and U27511 (N_27511,N_12392,N_15692);
and U27512 (N_27512,N_14136,N_14021);
and U27513 (N_27513,N_19082,N_13847);
and U27514 (N_27514,N_15194,N_10066);
nor U27515 (N_27515,N_11690,N_17067);
and U27516 (N_27516,N_13931,N_19746);
and U27517 (N_27517,N_16959,N_19068);
xnor U27518 (N_27518,N_15453,N_19159);
xor U27519 (N_27519,N_19487,N_19199);
or U27520 (N_27520,N_14793,N_14779);
xnor U27521 (N_27521,N_19858,N_17184);
nand U27522 (N_27522,N_15039,N_18959);
nand U27523 (N_27523,N_11706,N_11300);
xnor U27524 (N_27524,N_15849,N_10035);
and U27525 (N_27525,N_17042,N_12780);
or U27526 (N_27526,N_12414,N_10926);
and U27527 (N_27527,N_16936,N_11069);
or U27528 (N_27528,N_12396,N_14165);
nand U27529 (N_27529,N_16417,N_15328);
xor U27530 (N_27530,N_12488,N_15115);
xor U27531 (N_27531,N_10489,N_15902);
and U27532 (N_27532,N_12591,N_11179);
and U27533 (N_27533,N_16112,N_10027);
or U27534 (N_27534,N_14495,N_15122);
xnor U27535 (N_27535,N_11858,N_13372);
and U27536 (N_27536,N_17958,N_18425);
nand U27537 (N_27537,N_17001,N_10602);
or U27538 (N_27538,N_17448,N_18668);
and U27539 (N_27539,N_14451,N_12210);
xor U27540 (N_27540,N_12132,N_15432);
xor U27541 (N_27541,N_19602,N_10602);
and U27542 (N_27542,N_15461,N_19202);
or U27543 (N_27543,N_14480,N_13447);
nor U27544 (N_27544,N_12831,N_15134);
nand U27545 (N_27545,N_16498,N_13138);
nand U27546 (N_27546,N_10542,N_14581);
nand U27547 (N_27547,N_11202,N_19431);
or U27548 (N_27548,N_15857,N_17282);
or U27549 (N_27549,N_14554,N_11116);
and U27550 (N_27550,N_10789,N_14734);
nand U27551 (N_27551,N_14105,N_16834);
xor U27552 (N_27552,N_16818,N_15363);
nand U27553 (N_27553,N_10950,N_11935);
nor U27554 (N_27554,N_11643,N_16544);
or U27555 (N_27555,N_19292,N_18931);
nand U27556 (N_27556,N_17707,N_16674);
and U27557 (N_27557,N_19127,N_11581);
nand U27558 (N_27558,N_15259,N_12482);
xnor U27559 (N_27559,N_11654,N_12725);
or U27560 (N_27560,N_12921,N_15911);
or U27561 (N_27561,N_10343,N_13910);
or U27562 (N_27562,N_14594,N_19559);
xnor U27563 (N_27563,N_10029,N_10721);
or U27564 (N_27564,N_15477,N_18238);
and U27565 (N_27565,N_11837,N_15287);
xnor U27566 (N_27566,N_13936,N_10026);
nand U27567 (N_27567,N_13923,N_14515);
or U27568 (N_27568,N_10340,N_13628);
xnor U27569 (N_27569,N_19069,N_13274);
nand U27570 (N_27570,N_11181,N_11711);
nor U27571 (N_27571,N_18760,N_14369);
nor U27572 (N_27572,N_12839,N_15844);
xnor U27573 (N_27573,N_10609,N_12183);
xor U27574 (N_27574,N_10488,N_15684);
or U27575 (N_27575,N_13564,N_16239);
xor U27576 (N_27576,N_18217,N_13337);
or U27577 (N_27577,N_16291,N_12183);
xnor U27578 (N_27578,N_19027,N_18349);
nor U27579 (N_27579,N_16482,N_18217);
nor U27580 (N_27580,N_18319,N_12600);
nand U27581 (N_27581,N_10419,N_19372);
xnor U27582 (N_27582,N_13171,N_18577);
and U27583 (N_27583,N_16821,N_17698);
nand U27584 (N_27584,N_11721,N_19780);
or U27585 (N_27585,N_11534,N_15830);
and U27586 (N_27586,N_19481,N_11155);
nor U27587 (N_27587,N_13149,N_17411);
nand U27588 (N_27588,N_10896,N_16053);
nand U27589 (N_27589,N_10724,N_15565);
nor U27590 (N_27590,N_18249,N_11914);
nand U27591 (N_27591,N_18758,N_19514);
or U27592 (N_27592,N_17136,N_16497);
or U27593 (N_27593,N_10949,N_10384);
nand U27594 (N_27594,N_12671,N_10422);
and U27595 (N_27595,N_11861,N_12241);
xor U27596 (N_27596,N_14334,N_16928);
nor U27597 (N_27597,N_10683,N_12180);
or U27598 (N_27598,N_16911,N_12869);
or U27599 (N_27599,N_18212,N_10957);
or U27600 (N_27600,N_11766,N_15968);
or U27601 (N_27601,N_18812,N_17913);
and U27602 (N_27602,N_16778,N_19841);
xnor U27603 (N_27603,N_14411,N_14892);
nand U27604 (N_27604,N_13971,N_15486);
nand U27605 (N_27605,N_13765,N_11740);
xnor U27606 (N_27606,N_18588,N_12943);
or U27607 (N_27607,N_15391,N_14643);
or U27608 (N_27608,N_16553,N_11349);
xor U27609 (N_27609,N_14297,N_15167);
or U27610 (N_27610,N_13031,N_19798);
and U27611 (N_27611,N_19193,N_12141);
nor U27612 (N_27612,N_18962,N_14596);
xnor U27613 (N_27613,N_12040,N_16645);
xnor U27614 (N_27614,N_15100,N_16978);
or U27615 (N_27615,N_15778,N_12928);
nor U27616 (N_27616,N_12632,N_10150);
xnor U27617 (N_27617,N_10151,N_16228);
nand U27618 (N_27618,N_11416,N_15447);
nand U27619 (N_27619,N_19959,N_13829);
or U27620 (N_27620,N_16943,N_11442);
nor U27621 (N_27621,N_11054,N_16064);
nand U27622 (N_27622,N_18521,N_11634);
or U27623 (N_27623,N_13524,N_14599);
nor U27624 (N_27624,N_16331,N_11150);
nor U27625 (N_27625,N_14999,N_17195);
nand U27626 (N_27626,N_12072,N_18099);
or U27627 (N_27627,N_13596,N_17655);
nand U27628 (N_27628,N_17328,N_18814);
or U27629 (N_27629,N_14676,N_12052);
and U27630 (N_27630,N_16421,N_14212);
nand U27631 (N_27631,N_10221,N_11593);
nand U27632 (N_27632,N_14656,N_17778);
nor U27633 (N_27633,N_14680,N_19933);
nor U27634 (N_27634,N_17448,N_11998);
xor U27635 (N_27635,N_19955,N_14296);
xnor U27636 (N_27636,N_12052,N_17321);
and U27637 (N_27637,N_18359,N_18423);
and U27638 (N_27638,N_14746,N_15612);
xor U27639 (N_27639,N_13330,N_12576);
and U27640 (N_27640,N_13491,N_14494);
and U27641 (N_27641,N_14474,N_10398);
xnor U27642 (N_27642,N_11739,N_14409);
or U27643 (N_27643,N_14760,N_11355);
xnor U27644 (N_27644,N_14616,N_16740);
and U27645 (N_27645,N_11811,N_11729);
nor U27646 (N_27646,N_19386,N_10384);
xor U27647 (N_27647,N_16811,N_10678);
and U27648 (N_27648,N_18218,N_17935);
or U27649 (N_27649,N_11350,N_15904);
nor U27650 (N_27650,N_15068,N_18418);
or U27651 (N_27651,N_11301,N_18233);
and U27652 (N_27652,N_18967,N_14313);
and U27653 (N_27653,N_10598,N_15956);
and U27654 (N_27654,N_10964,N_14174);
nor U27655 (N_27655,N_18459,N_18357);
xnor U27656 (N_27656,N_11057,N_12078);
nor U27657 (N_27657,N_11949,N_10600);
nor U27658 (N_27658,N_18618,N_18897);
or U27659 (N_27659,N_12558,N_14743);
xnor U27660 (N_27660,N_10177,N_16438);
and U27661 (N_27661,N_17088,N_10141);
or U27662 (N_27662,N_12694,N_11234);
xnor U27663 (N_27663,N_19619,N_12134);
xnor U27664 (N_27664,N_14839,N_11850);
nand U27665 (N_27665,N_10238,N_16306);
or U27666 (N_27666,N_11461,N_15115);
nand U27667 (N_27667,N_18196,N_18326);
nor U27668 (N_27668,N_16715,N_11316);
xnor U27669 (N_27669,N_12920,N_11910);
and U27670 (N_27670,N_10085,N_12478);
xor U27671 (N_27671,N_10234,N_18942);
and U27672 (N_27672,N_14973,N_19600);
nor U27673 (N_27673,N_14862,N_19766);
and U27674 (N_27674,N_16223,N_13242);
xnor U27675 (N_27675,N_15943,N_15250);
nand U27676 (N_27676,N_13273,N_16414);
and U27677 (N_27677,N_15808,N_19360);
nor U27678 (N_27678,N_10002,N_18329);
xnor U27679 (N_27679,N_15692,N_14512);
nand U27680 (N_27680,N_18628,N_14098);
or U27681 (N_27681,N_15653,N_17788);
nor U27682 (N_27682,N_13656,N_10856);
xor U27683 (N_27683,N_16766,N_14590);
xnor U27684 (N_27684,N_19510,N_15154);
nor U27685 (N_27685,N_10217,N_18666);
nand U27686 (N_27686,N_16305,N_15210);
nand U27687 (N_27687,N_16931,N_13906);
xnor U27688 (N_27688,N_16902,N_13631);
nand U27689 (N_27689,N_10954,N_15199);
and U27690 (N_27690,N_15757,N_10734);
xnor U27691 (N_27691,N_14978,N_15032);
and U27692 (N_27692,N_18876,N_16888);
and U27693 (N_27693,N_12122,N_11298);
nand U27694 (N_27694,N_11261,N_10632);
xor U27695 (N_27695,N_16288,N_13356);
and U27696 (N_27696,N_14313,N_18200);
xor U27697 (N_27697,N_18434,N_17281);
xnor U27698 (N_27698,N_11501,N_16108);
and U27699 (N_27699,N_17263,N_16142);
xnor U27700 (N_27700,N_13219,N_18216);
xor U27701 (N_27701,N_16414,N_12489);
or U27702 (N_27702,N_11068,N_10683);
nor U27703 (N_27703,N_11982,N_14970);
and U27704 (N_27704,N_19623,N_11525);
nand U27705 (N_27705,N_12928,N_15332);
nor U27706 (N_27706,N_13892,N_14855);
and U27707 (N_27707,N_12026,N_11404);
or U27708 (N_27708,N_17425,N_14152);
nor U27709 (N_27709,N_12351,N_18713);
nand U27710 (N_27710,N_10871,N_12526);
and U27711 (N_27711,N_15714,N_19256);
xnor U27712 (N_27712,N_16935,N_14890);
xor U27713 (N_27713,N_18071,N_18452);
or U27714 (N_27714,N_18723,N_12341);
xor U27715 (N_27715,N_13982,N_10152);
nand U27716 (N_27716,N_19885,N_18934);
nand U27717 (N_27717,N_12880,N_17064);
xnor U27718 (N_27718,N_12797,N_11979);
xor U27719 (N_27719,N_13572,N_15779);
nor U27720 (N_27720,N_10474,N_14461);
nand U27721 (N_27721,N_10645,N_17220);
nand U27722 (N_27722,N_12574,N_18472);
nand U27723 (N_27723,N_15691,N_13746);
nand U27724 (N_27724,N_13366,N_18665);
and U27725 (N_27725,N_12735,N_18353);
xor U27726 (N_27726,N_16096,N_10406);
nor U27727 (N_27727,N_15920,N_17094);
or U27728 (N_27728,N_15114,N_12621);
nor U27729 (N_27729,N_15507,N_11535);
and U27730 (N_27730,N_11695,N_18883);
xor U27731 (N_27731,N_13197,N_19248);
xnor U27732 (N_27732,N_16841,N_18007);
or U27733 (N_27733,N_18798,N_15902);
and U27734 (N_27734,N_19268,N_13577);
and U27735 (N_27735,N_11280,N_15426);
or U27736 (N_27736,N_13423,N_16922);
nand U27737 (N_27737,N_12728,N_13973);
or U27738 (N_27738,N_11790,N_18925);
xor U27739 (N_27739,N_16708,N_14188);
or U27740 (N_27740,N_17116,N_13273);
and U27741 (N_27741,N_13123,N_16330);
nand U27742 (N_27742,N_15617,N_18455);
xnor U27743 (N_27743,N_12226,N_17099);
xnor U27744 (N_27744,N_11344,N_17291);
xor U27745 (N_27745,N_15917,N_11674);
nand U27746 (N_27746,N_10935,N_19870);
or U27747 (N_27747,N_18814,N_19986);
and U27748 (N_27748,N_16293,N_11554);
xnor U27749 (N_27749,N_19931,N_16938);
and U27750 (N_27750,N_19167,N_10832);
nor U27751 (N_27751,N_13994,N_11843);
nor U27752 (N_27752,N_15968,N_17629);
xor U27753 (N_27753,N_10644,N_18376);
or U27754 (N_27754,N_11941,N_10157);
or U27755 (N_27755,N_11067,N_17389);
or U27756 (N_27756,N_18416,N_19518);
or U27757 (N_27757,N_19395,N_10224);
nand U27758 (N_27758,N_16769,N_17310);
nand U27759 (N_27759,N_10853,N_11655);
xnor U27760 (N_27760,N_11365,N_19205);
nand U27761 (N_27761,N_11313,N_16818);
nand U27762 (N_27762,N_17511,N_11039);
nand U27763 (N_27763,N_18113,N_13563);
nor U27764 (N_27764,N_14411,N_15319);
or U27765 (N_27765,N_13878,N_13275);
or U27766 (N_27766,N_11332,N_13873);
or U27767 (N_27767,N_13357,N_12378);
nor U27768 (N_27768,N_11530,N_19183);
and U27769 (N_27769,N_15398,N_16635);
xnor U27770 (N_27770,N_15532,N_13550);
nor U27771 (N_27771,N_19993,N_19689);
nor U27772 (N_27772,N_16435,N_13364);
or U27773 (N_27773,N_10017,N_10671);
or U27774 (N_27774,N_11269,N_18373);
or U27775 (N_27775,N_18274,N_12608);
and U27776 (N_27776,N_14219,N_17590);
xnor U27777 (N_27777,N_19223,N_18012);
xnor U27778 (N_27778,N_14888,N_12835);
nand U27779 (N_27779,N_10423,N_12546);
nand U27780 (N_27780,N_15086,N_11832);
xor U27781 (N_27781,N_12993,N_13534);
nor U27782 (N_27782,N_12938,N_15827);
xor U27783 (N_27783,N_14390,N_10168);
xor U27784 (N_27784,N_15716,N_18821);
nand U27785 (N_27785,N_19536,N_19148);
xnor U27786 (N_27786,N_16924,N_18939);
xnor U27787 (N_27787,N_17196,N_18042);
and U27788 (N_27788,N_15217,N_10793);
nand U27789 (N_27789,N_12681,N_14486);
xor U27790 (N_27790,N_14192,N_19453);
xnor U27791 (N_27791,N_10473,N_16435);
or U27792 (N_27792,N_15882,N_13931);
nand U27793 (N_27793,N_19588,N_13812);
and U27794 (N_27794,N_13380,N_17612);
or U27795 (N_27795,N_10301,N_17316);
xnor U27796 (N_27796,N_15400,N_11945);
xor U27797 (N_27797,N_19204,N_19716);
and U27798 (N_27798,N_11227,N_11141);
xnor U27799 (N_27799,N_18742,N_18895);
nand U27800 (N_27800,N_14593,N_14627);
xor U27801 (N_27801,N_19694,N_15383);
xnor U27802 (N_27802,N_15413,N_10344);
or U27803 (N_27803,N_18328,N_12459);
or U27804 (N_27804,N_16006,N_13639);
nor U27805 (N_27805,N_12770,N_15880);
or U27806 (N_27806,N_11115,N_17740);
nor U27807 (N_27807,N_15935,N_10190);
xor U27808 (N_27808,N_13620,N_10103);
nand U27809 (N_27809,N_11068,N_13902);
nor U27810 (N_27810,N_15884,N_11709);
nand U27811 (N_27811,N_17195,N_11466);
or U27812 (N_27812,N_11162,N_10752);
nor U27813 (N_27813,N_13554,N_10609);
nand U27814 (N_27814,N_13612,N_16881);
nand U27815 (N_27815,N_10601,N_15438);
xor U27816 (N_27816,N_19795,N_11578);
nor U27817 (N_27817,N_12611,N_17283);
nand U27818 (N_27818,N_16296,N_15575);
xor U27819 (N_27819,N_13073,N_19161);
and U27820 (N_27820,N_16120,N_16915);
nor U27821 (N_27821,N_12085,N_19505);
nor U27822 (N_27822,N_13425,N_12064);
nor U27823 (N_27823,N_17299,N_16201);
xnor U27824 (N_27824,N_10815,N_18329);
or U27825 (N_27825,N_17123,N_19521);
xor U27826 (N_27826,N_16063,N_18803);
or U27827 (N_27827,N_12084,N_16193);
nand U27828 (N_27828,N_12902,N_18276);
nand U27829 (N_27829,N_15892,N_14826);
and U27830 (N_27830,N_16102,N_13496);
xor U27831 (N_27831,N_11324,N_19497);
or U27832 (N_27832,N_16094,N_13857);
xor U27833 (N_27833,N_10173,N_10125);
xnor U27834 (N_27834,N_16111,N_13082);
or U27835 (N_27835,N_11474,N_13310);
nand U27836 (N_27836,N_10160,N_15689);
nor U27837 (N_27837,N_18444,N_15616);
nand U27838 (N_27838,N_14729,N_11123);
nand U27839 (N_27839,N_15202,N_19091);
nor U27840 (N_27840,N_16638,N_10274);
nand U27841 (N_27841,N_14066,N_11369);
or U27842 (N_27842,N_13202,N_18301);
nor U27843 (N_27843,N_12632,N_15873);
nor U27844 (N_27844,N_12859,N_15915);
and U27845 (N_27845,N_10882,N_12323);
or U27846 (N_27846,N_19567,N_14449);
nand U27847 (N_27847,N_12166,N_12556);
and U27848 (N_27848,N_16238,N_14918);
nand U27849 (N_27849,N_14933,N_13619);
or U27850 (N_27850,N_12379,N_12081);
and U27851 (N_27851,N_13119,N_13767);
xor U27852 (N_27852,N_11094,N_11502);
nand U27853 (N_27853,N_19173,N_15109);
nor U27854 (N_27854,N_13904,N_10082);
or U27855 (N_27855,N_15660,N_16730);
xnor U27856 (N_27856,N_19799,N_17706);
nand U27857 (N_27857,N_18381,N_16171);
or U27858 (N_27858,N_10006,N_17029);
nor U27859 (N_27859,N_17607,N_16047);
nand U27860 (N_27860,N_11725,N_19184);
xnor U27861 (N_27861,N_14810,N_19250);
or U27862 (N_27862,N_19819,N_19903);
and U27863 (N_27863,N_14078,N_17879);
and U27864 (N_27864,N_15100,N_13156);
xnor U27865 (N_27865,N_11036,N_19066);
nand U27866 (N_27866,N_17754,N_13252);
nor U27867 (N_27867,N_19147,N_11970);
nand U27868 (N_27868,N_12070,N_17940);
and U27869 (N_27869,N_19251,N_19243);
xor U27870 (N_27870,N_10450,N_12833);
nor U27871 (N_27871,N_11582,N_17762);
nand U27872 (N_27872,N_14142,N_17477);
nor U27873 (N_27873,N_10909,N_15781);
xor U27874 (N_27874,N_19902,N_18025);
or U27875 (N_27875,N_12471,N_15680);
nor U27876 (N_27876,N_10613,N_10996);
nand U27877 (N_27877,N_13864,N_14102);
xor U27878 (N_27878,N_15371,N_13071);
xor U27879 (N_27879,N_15308,N_14970);
nor U27880 (N_27880,N_19543,N_11083);
xor U27881 (N_27881,N_15769,N_19386);
nand U27882 (N_27882,N_13812,N_12082);
or U27883 (N_27883,N_15805,N_14267);
or U27884 (N_27884,N_18501,N_17431);
or U27885 (N_27885,N_19546,N_18006);
xnor U27886 (N_27886,N_14013,N_10057);
nand U27887 (N_27887,N_19225,N_19932);
xor U27888 (N_27888,N_14686,N_10718);
nand U27889 (N_27889,N_12655,N_18305);
and U27890 (N_27890,N_17593,N_10748);
nand U27891 (N_27891,N_18064,N_16612);
and U27892 (N_27892,N_17717,N_14130);
or U27893 (N_27893,N_17346,N_13251);
nand U27894 (N_27894,N_15347,N_12192);
xnor U27895 (N_27895,N_15195,N_16041);
xnor U27896 (N_27896,N_19608,N_12340);
and U27897 (N_27897,N_18812,N_19333);
nor U27898 (N_27898,N_11986,N_13550);
nand U27899 (N_27899,N_13688,N_13766);
xnor U27900 (N_27900,N_18659,N_10919);
nand U27901 (N_27901,N_15916,N_14680);
nor U27902 (N_27902,N_14580,N_15686);
nor U27903 (N_27903,N_15549,N_13879);
xor U27904 (N_27904,N_19436,N_17967);
nor U27905 (N_27905,N_18094,N_19338);
and U27906 (N_27906,N_19114,N_15539);
and U27907 (N_27907,N_10369,N_13072);
or U27908 (N_27908,N_14521,N_18044);
or U27909 (N_27909,N_14837,N_10720);
nand U27910 (N_27910,N_18771,N_17495);
and U27911 (N_27911,N_11742,N_11205);
and U27912 (N_27912,N_11480,N_12337);
xor U27913 (N_27913,N_13625,N_13360);
nand U27914 (N_27914,N_18006,N_15278);
xnor U27915 (N_27915,N_18473,N_15032);
nor U27916 (N_27916,N_19066,N_15695);
nor U27917 (N_27917,N_17508,N_10392);
xor U27918 (N_27918,N_10696,N_13789);
nand U27919 (N_27919,N_19923,N_12060);
nor U27920 (N_27920,N_19355,N_12558);
and U27921 (N_27921,N_12004,N_17136);
and U27922 (N_27922,N_18677,N_17617);
nand U27923 (N_27923,N_13881,N_12300);
or U27924 (N_27924,N_19779,N_15697);
nor U27925 (N_27925,N_13226,N_13338);
nor U27926 (N_27926,N_14626,N_19999);
or U27927 (N_27927,N_13495,N_10928);
nand U27928 (N_27928,N_17012,N_15158);
xnor U27929 (N_27929,N_11869,N_11614);
xnor U27930 (N_27930,N_10770,N_19822);
and U27931 (N_27931,N_15740,N_12800);
and U27932 (N_27932,N_14918,N_12436);
or U27933 (N_27933,N_18953,N_18802);
nor U27934 (N_27934,N_18696,N_18641);
nand U27935 (N_27935,N_15630,N_18222);
or U27936 (N_27936,N_10969,N_19923);
and U27937 (N_27937,N_14591,N_10496);
or U27938 (N_27938,N_17213,N_12673);
nand U27939 (N_27939,N_17589,N_14638);
or U27940 (N_27940,N_16348,N_15643);
nor U27941 (N_27941,N_14207,N_10452);
nand U27942 (N_27942,N_15190,N_14956);
nor U27943 (N_27943,N_14230,N_19858);
and U27944 (N_27944,N_18152,N_11365);
xor U27945 (N_27945,N_11866,N_12013);
xnor U27946 (N_27946,N_19260,N_19379);
and U27947 (N_27947,N_14085,N_15434);
or U27948 (N_27948,N_10517,N_15907);
xor U27949 (N_27949,N_11275,N_12134);
nand U27950 (N_27950,N_13433,N_19195);
nor U27951 (N_27951,N_11051,N_17883);
nand U27952 (N_27952,N_13243,N_15618);
and U27953 (N_27953,N_11397,N_14682);
or U27954 (N_27954,N_14904,N_16551);
nor U27955 (N_27955,N_11535,N_18122);
nor U27956 (N_27956,N_13348,N_12882);
and U27957 (N_27957,N_14725,N_12094);
nand U27958 (N_27958,N_11898,N_10885);
and U27959 (N_27959,N_17608,N_10320);
xnor U27960 (N_27960,N_19488,N_15446);
or U27961 (N_27961,N_12737,N_17952);
nand U27962 (N_27962,N_16511,N_12032);
or U27963 (N_27963,N_16365,N_18159);
nor U27964 (N_27964,N_13817,N_11150);
and U27965 (N_27965,N_12925,N_10843);
xnor U27966 (N_27966,N_13984,N_16500);
and U27967 (N_27967,N_14255,N_15633);
nor U27968 (N_27968,N_10054,N_15833);
nand U27969 (N_27969,N_10407,N_17909);
nor U27970 (N_27970,N_16598,N_11671);
or U27971 (N_27971,N_18599,N_17715);
nand U27972 (N_27972,N_15930,N_10836);
and U27973 (N_27973,N_17659,N_12837);
and U27974 (N_27974,N_12010,N_10729);
or U27975 (N_27975,N_15623,N_19665);
xor U27976 (N_27976,N_16659,N_14347);
and U27977 (N_27977,N_10517,N_13652);
or U27978 (N_27978,N_11328,N_12262);
nand U27979 (N_27979,N_19134,N_18925);
xor U27980 (N_27980,N_10839,N_18595);
xnor U27981 (N_27981,N_11014,N_17905);
nand U27982 (N_27982,N_10811,N_19484);
nand U27983 (N_27983,N_15797,N_13090);
and U27984 (N_27984,N_18134,N_11674);
nor U27985 (N_27985,N_19979,N_16941);
or U27986 (N_27986,N_17713,N_18204);
nor U27987 (N_27987,N_18901,N_11476);
nand U27988 (N_27988,N_17462,N_10834);
nand U27989 (N_27989,N_17824,N_12500);
nor U27990 (N_27990,N_19913,N_17205);
nand U27991 (N_27991,N_12662,N_16977);
or U27992 (N_27992,N_16756,N_12062);
and U27993 (N_27993,N_10509,N_14110);
nor U27994 (N_27994,N_12336,N_14049);
xnor U27995 (N_27995,N_11803,N_19744);
nand U27996 (N_27996,N_16445,N_11138);
nor U27997 (N_27997,N_11280,N_19930);
nand U27998 (N_27998,N_10724,N_19521);
xor U27999 (N_27999,N_12117,N_10829);
nand U28000 (N_28000,N_10499,N_17839);
nand U28001 (N_28001,N_11616,N_11933);
and U28002 (N_28002,N_16181,N_11499);
or U28003 (N_28003,N_19831,N_14656);
xor U28004 (N_28004,N_12350,N_14694);
or U28005 (N_28005,N_19458,N_12250);
nand U28006 (N_28006,N_15388,N_12822);
and U28007 (N_28007,N_14894,N_17346);
or U28008 (N_28008,N_12312,N_18984);
or U28009 (N_28009,N_13296,N_12816);
and U28010 (N_28010,N_18449,N_16047);
nor U28011 (N_28011,N_16915,N_18506);
or U28012 (N_28012,N_16044,N_12415);
xor U28013 (N_28013,N_13133,N_14614);
xnor U28014 (N_28014,N_18674,N_13950);
or U28015 (N_28015,N_10412,N_12537);
nor U28016 (N_28016,N_16465,N_16248);
nor U28017 (N_28017,N_17625,N_14885);
xnor U28018 (N_28018,N_11812,N_12881);
nor U28019 (N_28019,N_10354,N_18196);
xor U28020 (N_28020,N_15488,N_13935);
nor U28021 (N_28021,N_17547,N_19318);
nor U28022 (N_28022,N_17707,N_18715);
xnor U28023 (N_28023,N_13954,N_18777);
nand U28024 (N_28024,N_15157,N_16348);
or U28025 (N_28025,N_11348,N_10326);
or U28026 (N_28026,N_17192,N_18534);
nor U28027 (N_28027,N_12215,N_12222);
nand U28028 (N_28028,N_18709,N_11927);
nand U28029 (N_28029,N_15389,N_16859);
and U28030 (N_28030,N_10717,N_15489);
xor U28031 (N_28031,N_17762,N_15223);
xor U28032 (N_28032,N_13624,N_10725);
nor U28033 (N_28033,N_18820,N_16536);
xnor U28034 (N_28034,N_11953,N_17019);
nand U28035 (N_28035,N_10690,N_18396);
and U28036 (N_28036,N_12912,N_16164);
xnor U28037 (N_28037,N_12133,N_12971);
nand U28038 (N_28038,N_11098,N_12236);
nand U28039 (N_28039,N_17075,N_16137);
nor U28040 (N_28040,N_15107,N_12253);
and U28041 (N_28041,N_14362,N_18850);
or U28042 (N_28042,N_11039,N_12258);
xor U28043 (N_28043,N_18939,N_18485);
or U28044 (N_28044,N_13123,N_17011);
nand U28045 (N_28045,N_19096,N_11840);
and U28046 (N_28046,N_19390,N_10171);
nand U28047 (N_28047,N_18925,N_12503);
xor U28048 (N_28048,N_11652,N_13853);
nor U28049 (N_28049,N_12676,N_16843);
or U28050 (N_28050,N_15157,N_14206);
or U28051 (N_28051,N_10198,N_11668);
or U28052 (N_28052,N_11026,N_19368);
nand U28053 (N_28053,N_19778,N_11839);
nand U28054 (N_28054,N_16679,N_17891);
and U28055 (N_28055,N_14225,N_11230);
nand U28056 (N_28056,N_15128,N_16803);
xnor U28057 (N_28057,N_16362,N_11862);
nand U28058 (N_28058,N_10537,N_16435);
or U28059 (N_28059,N_11312,N_13753);
and U28060 (N_28060,N_11218,N_19633);
nor U28061 (N_28061,N_12530,N_18061);
nand U28062 (N_28062,N_19977,N_10310);
nand U28063 (N_28063,N_17610,N_15928);
nor U28064 (N_28064,N_19098,N_15473);
nor U28065 (N_28065,N_13902,N_13570);
or U28066 (N_28066,N_13523,N_18656);
or U28067 (N_28067,N_17250,N_19151);
or U28068 (N_28068,N_16111,N_12102);
xor U28069 (N_28069,N_16243,N_12455);
or U28070 (N_28070,N_17924,N_10556);
nor U28071 (N_28071,N_18888,N_17550);
or U28072 (N_28072,N_17810,N_19209);
and U28073 (N_28073,N_15552,N_18661);
xnor U28074 (N_28074,N_13254,N_17198);
nand U28075 (N_28075,N_19812,N_16499);
or U28076 (N_28076,N_13848,N_13703);
xor U28077 (N_28077,N_14319,N_14284);
and U28078 (N_28078,N_13159,N_14031);
and U28079 (N_28079,N_18322,N_12724);
and U28080 (N_28080,N_11759,N_10432);
and U28081 (N_28081,N_15279,N_14242);
xnor U28082 (N_28082,N_13501,N_17746);
nand U28083 (N_28083,N_10886,N_19604);
xor U28084 (N_28084,N_10601,N_19569);
xnor U28085 (N_28085,N_16590,N_18605);
xor U28086 (N_28086,N_13078,N_14899);
xor U28087 (N_28087,N_11569,N_13454);
and U28088 (N_28088,N_18887,N_12586);
nand U28089 (N_28089,N_13099,N_12403);
or U28090 (N_28090,N_15504,N_16375);
and U28091 (N_28091,N_11664,N_19595);
nand U28092 (N_28092,N_18061,N_18641);
xnor U28093 (N_28093,N_10962,N_19648);
and U28094 (N_28094,N_13954,N_14056);
xnor U28095 (N_28095,N_16989,N_10138);
nor U28096 (N_28096,N_11193,N_13068);
nand U28097 (N_28097,N_14752,N_14476);
nand U28098 (N_28098,N_14530,N_14268);
nor U28099 (N_28099,N_15813,N_19922);
xor U28100 (N_28100,N_10462,N_10147);
nor U28101 (N_28101,N_10281,N_11421);
nor U28102 (N_28102,N_12328,N_10353);
nand U28103 (N_28103,N_12054,N_15996);
nor U28104 (N_28104,N_19804,N_12590);
and U28105 (N_28105,N_14454,N_18174);
nor U28106 (N_28106,N_13597,N_14422);
nor U28107 (N_28107,N_14647,N_17012);
nor U28108 (N_28108,N_14708,N_13700);
and U28109 (N_28109,N_12310,N_17936);
and U28110 (N_28110,N_16197,N_13820);
xor U28111 (N_28111,N_11743,N_10576);
and U28112 (N_28112,N_16054,N_19443);
nand U28113 (N_28113,N_15033,N_12187);
nand U28114 (N_28114,N_12866,N_14801);
nor U28115 (N_28115,N_13021,N_13248);
nor U28116 (N_28116,N_16387,N_12499);
xor U28117 (N_28117,N_17428,N_19907);
or U28118 (N_28118,N_17640,N_14531);
xor U28119 (N_28119,N_18871,N_14474);
xor U28120 (N_28120,N_11636,N_14272);
nand U28121 (N_28121,N_10003,N_11184);
and U28122 (N_28122,N_13256,N_13415);
or U28123 (N_28123,N_12213,N_14307);
xor U28124 (N_28124,N_14359,N_17366);
xor U28125 (N_28125,N_11202,N_19166);
or U28126 (N_28126,N_10637,N_13516);
nand U28127 (N_28127,N_11847,N_17015);
xnor U28128 (N_28128,N_14118,N_19660);
or U28129 (N_28129,N_16058,N_18767);
or U28130 (N_28130,N_11271,N_14672);
and U28131 (N_28131,N_10828,N_17263);
and U28132 (N_28132,N_18070,N_14514);
xor U28133 (N_28133,N_10011,N_13447);
and U28134 (N_28134,N_18789,N_13765);
and U28135 (N_28135,N_11130,N_18753);
nand U28136 (N_28136,N_19415,N_11920);
or U28137 (N_28137,N_18955,N_11677);
nand U28138 (N_28138,N_10377,N_14224);
or U28139 (N_28139,N_15478,N_11123);
xor U28140 (N_28140,N_14167,N_19595);
and U28141 (N_28141,N_15660,N_12873);
and U28142 (N_28142,N_13120,N_11163);
xor U28143 (N_28143,N_16730,N_10731);
and U28144 (N_28144,N_12885,N_14874);
or U28145 (N_28145,N_12757,N_18591);
and U28146 (N_28146,N_13353,N_14050);
nor U28147 (N_28147,N_17089,N_15275);
nor U28148 (N_28148,N_11405,N_16221);
nand U28149 (N_28149,N_11608,N_13568);
and U28150 (N_28150,N_10347,N_13979);
nor U28151 (N_28151,N_17669,N_19281);
and U28152 (N_28152,N_17306,N_16492);
nand U28153 (N_28153,N_13650,N_12982);
nor U28154 (N_28154,N_14228,N_12404);
xor U28155 (N_28155,N_16196,N_17860);
nand U28156 (N_28156,N_11899,N_14041);
nand U28157 (N_28157,N_19006,N_12558);
xor U28158 (N_28158,N_12452,N_17851);
nand U28159 (N_28159,N_19386,N_18593);
or U28160 (N_28160,N_15577,N_11565);
xor U28161 (N_28161,N_18841,N_16310);
and U28162 (N_28162,N_10805,N_10354);
xnor U28163 (N_28163,N_18951,N_14672);
and U28164 (N_28164,N_12804,N_14424);
xnor U28165 (N_28165,N_10182,N_10264);
or U28166 (N_28166,N_15469,N_11890);
and U28167 (N_28167,N_13274,N_17856);
and U28168 (N_28168,N_19164,N_10491);
nor U28169 (N_28169,N_12619,N_13441);
nor U28170 (N_28170,N_10504,N_10212);
or U28171 (N_28171,N_12941,N_19130);
nor U28172 (N_28172,N_17883,N_13600);
xnor U28173 (N_28173,N_19494,N_14283);
nor U28174 (N_28174,N_11635,N_17654);
nand U28175 (N_28175,N_12532,N_10815);
nor U28176 (N_28176,N_10218,N_16975);
nor U28177 (N_28177,N_10287,N_18013);
and U28178 (N_28178,N_15950,N_16937);
xnor U28179 (N_28179,N_10226,N_18239);
xor U28180 (N_28180,N_18612,N_19822);
nand U28181 (N_28181,N_10194,N_15558);
nand U28182 (N_28182,N_14921,N_14908);
and U28183 (N_28183,N_13458,N_11499);
and U28184 (N_28184,N_16363,N_15046);
nand U28185 (N_28185,N_12266,N_15001);
nor U28186 (N_28186,N_13611,N_19054);
xor U28187 (N_28187,N_14417,N_14879);
nand U28188 (N_28188,N_13691,N_11959);
or U28189 (N_28189,N_10073,N_16760);
nor U28190 (N_28190,N_14538,N_17149);
or U28191 (N_28191,N_11133,N_15015);
nor U28192 (N_28192,N_17875,N_15388);
nor U28193 (N_28193,N_13501,N_10530);
nand U28194 (N_28194,N_17092,N_12881);
nand U28195 (N_28195,N_13584,N_10192);
nand U28196 (N_28196,N_19809,N_13365);
or U28197 (N_28197,N_19437,N_15891);
nand U28198 (N_28198,N_13080,N_18620);
nand U28199 (N_28199,N_10401,N_13265);
nor U28200 (N_28200,N_12184,N_14089);
or U28201 (N_28201,N_15371,N_15970);
or U28202 (N_28202,N_13588,N_13143);
nand U28203 (N_28203,N_14065,N_17456);
nor U28204 (N_28204,N_14409,N_10771);
nor U28205 (N_28205,N_12199,N_17147);
or U28206 (N_28206,N_17921,N_17740);
or U28207 (N_28207,N_16795,N_15181);
nor U28208 (N_28208,N_14554,N_14842);
nor U28209 (N_28209,N_19147,N_17915);
xnor U28210 (N_28210,N_12333,N_11074);
and U28211 (N_28211,N_18759,N_12369);
and U28212 (N_28212,N_10626,N_18323);
nor U28213 (N_28213,N_14528,N_10086);
nor U28214 (N_28214,N_15435,N_13527);
xor U28215 (N_28215,N_11971,N_11347);
and U28216 (N_28216,N_17869,N_13655);
or U28217 (N_28217,N_14859,N_19143);
nand U28218 (N_28218,N_14711,N_12528);
and U28219 (N_28219,N_19597,N_13103);
nor U28220 (N_28220,N_15011,N_12498);
nor U28221 (N_28221,N_12152,N_13006);
nand U28222 (N_28222,N_15886,N_12682);
or U28223 (N_28223,N_13349,N_18408);
or U28224 (N_28224,N_13874,N_19566);
and U28225 (N_28225,N_17992,N_14461);
or U28226 (N_28226,N_13741,N_14409);
nand U28227 (N_28227,N_13624,N_18670);
or U28228 (N_28228,N_14595,N_17184);
and U28229 (N_28229,N_11232,N_19349);
nor U28230 (N_28230,N_14926,N_14910);
and U28231 (N_28231,N_16539,N_12830);
and U28232 (N_28232,N_11546,N_11231);
or U28233 (N_28233,N_18121,N_15084);
xor U28234 (N_28234,N_12597,N_13927);
nand U28235 (N_28235,N_17446,N_18210);
nor U28236 (N_28236,N_17966,N_13328);
and U28237 (N_28237,N_15677,N_15097);
or U28238 (N_28238,N_16133,N_10737);
and U28239 (N_28239,N_17802,N_12018);
xor U28240 (N_28240,N_13941,N_10425);
nor U28241 (N_28241,N_19278,N_17066);
nand U28242 (N_28242,N_16071,N_14265);
xnor U28243 (N_28243,N_11694,N_12243);
xor U28244 (N_28244,N_13113,N_19252);
and U28245 (N_28245,N_11272,N_18243);
and U28246 (N_28246,N_14525,N_17341);
nor U28247 (N_28247,N_16227,N_10767);
or U28248 (N_28248,N_19623,N_16125);
or U28249 (N_28249,N_16224,N_13650);
and U28250 (N_28250,N_15553,N_12996);
nand U28251 (N_28251,N_18963,N_14190);
and U28252 (N_28252,N_16850,N_19493);
nand U28253 (N_28253,N_14627,N_13643);
nand U28254 (N_28254,N_11036,N_17301);
nand U28255 (N_28255,N_12938,N_16891);
or U28256 (N_28256,N_17788,N_16346);
nand U28257 (N_28257,N_11775,N_19552);
nand U28258 (N_28258,N_15638,N_17892);
or U28259 (N_28259,N_17824,N_18224);
and U28260 (N_28260,N_11884,N_11423);
or U28261 (N_28261,N_19846,N_11523);
nor U28262 (N_28262,N_17023,N_10356);
and U28263 (N_28263,N_11012,N_11736);
nor U28264 (N_28264,N_18193,N_19625);
and U28265 (N_28265,N_12544,N_15242);
nor U28266 (N_28266,N_18007,N_13785);
or U28267 (N_28267,N_17389,N_15212);
and U28268 (N_28268,N_15297,N_18588);
nand U28269 (N_28269,N_19379,N_17243);
nand U28270 (N_28270,N_15120,N_18262);
nand U28271 (N_28271,N_16213,N_13104);
nor U28272 (N_28272,N_10589,N_13291);
or U28273 (N_28273,N_11312,N_12051);
and U28274 (N_28274,N_15724,N_13771);
nor U28275 (N_28275,N_10908,N_13599);
xor U28276 (N_28276,N_14609,N_19021);
and U28277 (N_28277,N_10028,N_15199);
or U28278 (N_28278,N_11703,N_18059);
nand U28279 (N_28279,N_10331,N_14972);
nor U28280 (N_28280,N_16083,N_19978);
and U28281 (N_28281,N_11784,N_11800);
nor U28282 (N_28282,N_17815,N_17937);
nand U28283 (N_28283,N_13916,N_14268);
and U28284 (N_28284,N_17867,N_16810);
and U28285 (N_28285,N_17990,N_18054);
and U28286 (N_28286,N_19243,N_12428);
and U28287 (N_28287,N_15841,N_18837);
xnor U28288 (N_28288,N_18870,N_17318);
nor U28289 (N_28289,N_14445,N_11794);
or U28290 (N_28290,N_11161,N_14123);
xor U28291 (N_28291,N_12462,N_10083);
nand U28292 (N_28292,N_15954,N_12101);
and U28293 (N_28293,N_13524,N_12210);
xnor U28294 (N_28294,N_17597,N_17038);
or U28295 (N_28295,N_16915,N_10571);
nor U28296 (N_28296,N_16691,N_19123);
xor U28297 (N_28297,N_12830,N_14476);
nand U28298 (N_28298,N_11225,N_10989);
nand U28299 (N_28299,N_15322,N_16595);
and U28300 (N_28300,N_11107,N_15226);
nor U28301 (N_28301,N_12578,N_10407);
nand U28302 (N_28302,N_11884,N_13846);
or U28303 (N_28303,N_16621,N_18993);
nand U28304 (N_28304,N_18004,N_10679);
nand U28305 (N_28305,N_17302,N_16642);
nor U28306 (N_28306,N_10086,N_13360);
nor U28307 (N_28307,N_11679,N_18611);
nand U28308 (N_28308,N_10054,N_17935);
nor U28309 (N_28309,N_16955,N_11486);
nor U28310 (N_28310,N_19730,N_13347);
and U28311 (N_28311,N_17680,N_14132);
and U28312 (N_28312,N_14158,N_12044);
or U28313 (N_28313,N_11766,N_16369);
nand U28314 (N_28314,N_14755,N_17018);
nand U28315 (N_28315,N_12509,N_11047);
or U28316 (N_28316,N_12677,N_18991);
nand U28317 (N_28317,N_12438,N_15557);
nor U28318 (N_28318,N_11861,N_16697);
xnor U28319 (N_28319,N_14425,N_19350);
nor U28320 (N_28320,N_12761,N_10540);
nand U28321 (N_28321,N_18055,N_10288);
nand U28322 (N_28322,N_13739,N_15420);
xnor U28323 (N_28323,N_15659,N_17515);
or U28324 (N_28324,N_19925,N_18855);
nand U28325 (N_28325,N_11116,N_17051);
and U28326 (N_28326,N_14098,N_19263);
or U28327 (N_28327,N_18421,N_13812);
xnor U28328 (N_28328,N_12763,N_15655);
and U28329 (N_28329,N_17036,N_11727);
and U28330 (N_28330,N_12244,N_18934);
and U28331 (N_28331,N_17033,N_10723);
nand U28332 (N_28332,N_11944,N_14346);
xor U28333 (N_28333,N_12478,N_12369);
nand U28334 (N_28334,N_10759,N_14574);
nor U28335 (N_28335,N_19055,N_17121);
nor U28336 (N_28336,N_14503,N_15231);
xnor U28337 (N_28337,N_12403,N_12794);
or U28338 (N_28338,N_11651,N_19556);
nand U28339 (N_28339,N_17880,N_15490);
nor U28340 (N_28340,N_16066,N_19151);
and U28341 (N_28341,N_19929,N_15177);
or U28342 (N_28342,N_15351,N_14554);
nand U28343 (N_28343,N_11628,N_14966);
and U28344 (N_28344,N_11477,N_12295);
nor U28345 (N_28345,N_13527,N_10082);
nor U28346 (N_28346,N_19990,N_10334);
and U28347 (N_28347,N_19315,N_15659);
nor U28348 (N_28348,N_12622,N_11808);
and U28349 (N_28349,N_15263,N_12735);
nor U28350 (N_28350,N_11990,N_18196);
nand U28351 (N_28351,N_11674,N_18404);
xnor U28352 (N_28352,N_13259,N_17771);
nand U28353 (N_28353,N_11962,N_11292);
and U28354 (N_28354,N_13632,N_15791);
and U28355 (N_28355,N_11993,N_10222);
or U28356 (N_28356,N_17210,N_18836);
or U28357 (N_28357,N_13154,N_12524);
xor U28358 (N_28358,N_13148,N_14361);
xnor U28359 (N_28359,N_10800,N_17805);
nand U28360 (N_28360,N_19859,N_13472);
and U28361 (N_28361,N_12711,N_11476);
nor U28362 (N_28362,N_17577,N_19222);
and U28363 (N_28363,N_18711,N_13647);
nand U28364 (N_28364,N_15145,N_15680);
or U28365 (N_28365,N_11940,N_17624);
and U28366 (N_28366,N_15050,N_16934);
xor U28367 (N_28367,N_11544,N_12845);
nand U28368 (N_28368,N_15145,N_14844);
xor U28369 (N_28369,N_13640,N_18635);
or U28370 (N_28370,N_10672,N_19413);
or U28371 (N_28371,N_16176,N_14743);
or U28372 (N_28372,N_12981,N_18915);
nor U28373 (N_28373,N_15935,N_13246);
and U28374 (N_28374,N_17829,N_12261);
or U28375 (N_28375,N_18625,N_12373);
xor U28376 (N_28376,N_19808,N_15250);
nand U28377 (N_28377,N_16355,N_19679);
nor U28378 (N_28378,N_19373,N_16806);
xnor U28379 (N_28379,N_10813,N_16473);
and U28380 (N_28380,N_15693,N_15270);
or U28381 (N_28381,N_15371,N_16491);
or U28382 (N_28382,N_17845,N_11138);
nand U28383 (N_28383,N_14541,N_11745);
xnor U28384 (N_28384,N_15063,N_10081);
and U28385 (N_28385,N_16551,N_12234);
and U28386 (N_28386,N_15820,N_19801);
or U28387 (N_28387,N_14341,N_17396);
or U28388 (N_28388,N_13670,N_16992);
or U28389 (N_28389,N_12223,N_18030);
nor U28390 (N_28390,N_12227,N_12440);
nand U28391 (N_28391,N_15200,N_10671);
and U28392 (N_28392,N_16201,N_19542);
nand U28393 (N_28393,N_11443,N_18345);
nor U28394 (N_28394,N_16369,N_16045);
nor U28395 (N_28395,N_13544,N_13738);
or U28396 (N_28396,N_14678,N_18010);
or U28397 (N_28397,N_15079,N_15652);
and U28398 (N_28398,N_16589,N_11190);
nand U28399 (N_28399,N_12614,N_11795);
and U28400 (N_28400,N_13283,N_13514);
and U28401 (N_28401,N_16990,N_11150);
and U28402 (N_28402,N_15560,N_12280);
nand U28403 (N_28403,N_14596,N_12719);
nand U28404 (N_28404,N_17014,N_15011);
nand U28405 (N_28405,N_11687,N_10975);
nor U28406 (N_28406,N_10994,N_18891);
xnor U28407 (N_28407,N_13253,N_11744);
nor U28408 (N_28408,N_17196,N_15679);
nor U28409 (N_28409,N_11873,N_14158);
nand U28410 (N_28410,N_10568,N_10067);
nand U28411 (N_28411,N_10362,N_14446);
nor U28412 (N_28412,N_18566,N_14791);
and U28413 (N_28413,N_18238,N_15539);
xnor U28414 (N_28414,N_13620,N_14891);
or U28415 (N_28415,N_14033,N_19667);
and U28416 (N_28416,N_19492,N_18739);
and U28417 (N_28417,N_16818,N_15176);
nor U28418 (N_28418,N_19142,N_17410);
nand U28419 (N_28419,N_19281,N_19930);
or U28420 (N_28420,N_18061,N_12316);
and U28421 (N_28421,N_11689,N_14341);
and U28422 (N_28422,N_10207,N_11141);
and U28423 (N_28423,N_16044,N_13876);
or U28424 (N_28424,N_15890,N_11994);
and U28425 (N_28425,N_13988,N_10847);
nor U28426 (N_28426,N_15822,N_18243);
or U28427 (N_28427,N_13364,N_11582);
xnor U28428 (N_28428,N_13428,N_15082);
and U28429 (N_28429,N_18426,N_13610);
nor U28430 (N_28430,N_17990,N_10287);
xnor U28431 (N_28431,N_18011,N_19305);
xor U28432 (N_28432,N_11671,N_19621);
xor U28433 (N_28433,N_10218,N_12040);
and U28434 (N_28434,N_13398,N_19304);
xnor U28435 (N_28435,N_19401,N_13486);
and U28436 (N_28436,N_11885,N_12858);
nand U28437 (N_28437,N_14193,N_18255);
xor U28438 (N_28438,N_15232,N_18432);
or U28439 (N_28439,N_14085,N_16605);
nor U28440 (N_28440,N_16595,N_18311);
or U28441 (N_28441,N_18338,N_14907);
xnor U28442 (N_28442,N_13763,N_13789);
nor U28443 (N_28443,N_13924,N_12332);
nor U28444 (N_28444,N_19864,N_15157);
nor U28445 (N_28445,N_16115,N_19642);
or U28446 (N_28446,N_18750,N_12831);
or U28447 (N_28447,N_13825,N_15198);
and U28448 (N_28448,N_12156,N_15221);
and U28449 (N_28449,N_14419,N_11058);
or U28450 (N_28450,N_11861,N_18692);
xor U28451 (N_28451,N_19465,N_11935);
xnor U28452 (N_28452,N_10008,N_11620);
or U28453 (N_28453,N_13187,N_12764);
xor U28454 (N_28454,N_17620,N_17003);
or U28455 (N_28455,N_11110,N_12274);
nor U28456 (N_28456,N_18901,N_18455);
nor U28457 (N_28457,N_10668,N_19822);
or U28458 (N_28458,N_14579,N_13989);
and U28459 (N_28459,N_14475,N_12209);
xnor U28460 (N_28460,N_15837,N_15162);
xor U28461 (N_28461,N_14270,N_18367);
nand U28462 (N_28462,N_15247,N_11793);
nand U28463 (N_28463,N_19804,N_18614);
nand U28464 (N_28464,N_12417,N_16207);
nand U28465 (N_28465,N_18076,N_14964);
or U28466 (N_28466,N_16155,N_12695);
xor U28467 (N_28467,N_14781,N_14423);
nand U28468 (N_28468,N_16649,N_11923);
nand U28469 (N_28469,N_17660,N_19499);
nor U28470 (N_28470,N_17169,N_15629);
nand U28471 (N_28471,N_16661,N_19860);
and U28472 (N_28472,N_10750,N_19785);
and U28473 (N_28473,N_16784,N_17932);
xor U28474 (N_28474,N_16505,N_10124);
and U28475 (N_28475,N_18682,N_13782);
xnor U28476 (N_28476,N_12274,N_14421);
nor U28477 (N_28477,N_15784,N_14215);
xor U28478 (N_28478,N_11068,N_15223);
nor U28479 (N_28479,N_11889,N_18242);
nand U28480 (N_28480,N_10031,N_16348);
nand U28481 (N_28481,N_17425,N_16365);
and U28482 (N_28482,N_13567,N_13852);
xor U28483 (N_28483,N_16790,N_19299);
nand U28484 (N_28484,N_18398,N_10157);
or U28485 (N_28485,N_17744,N_11761);
or U28486 (N_28486,N_17844,N_17601);
or U28487 (N_28487,N_11505,N_14746);
nor U28488 (N_28488,N_15658,N_18537);
and U28489 (N_28489,N_17287,N_10006);
and U28490 (N_28490,N_17691,N_12251);
or U28491 (N_28491,N_11017,N_14822);
xnor U28492 (N_28492,N_14729,N_10029);
xnor U28493 (N_28493,N_19484,N_14134);
and U28494 (N_28494,N_16400,N_18666);
nand U28495 (N_28495,N_18653,N_12602);
nand U28496 (N_28496,N_11927,N_13180);
xnor U28497 (N_28497,N_10145,N_13475);
or U28498 (N_28498,N_17927,N_18639);
and U28499 (N_28499,N_11419,N_12037);
nor U28500 (N_28500,N_11770,N_14055);
nand U28501 (N_28501,N_19313,N_16658);
or U28502 (N_28502,N_13664,N_16325);
or U28503 (N_28503,N_17878,N_12743);
and U28504 (N_28504,N_12976,N_12140);
xor U28505 (N_28505,N_11940,N_16897);
nand U28506 (N_28506,N_14798,N_12381);
xor U28507 (N_28507,N_10952,N_19251);
nor U28508 (N_28508,N_10764,N_14871);
or U28509 (N_28509,N_14178,N_17579);
nor U28510 (N_28510,N_10549,N_16296);
or U28511 (N_28511,N_19857,N_19091);
and U28512 (N_28512,N_14764,N_19502);
xor U28513 (N_28513,N_16972,N_15949);
nand U28514 (N_28514,N_17324,N_19890);
or U28515 (N_28515,N_12648,N_10977);
and U28516 (N_28516,N_15606,N_11054);
xor U28517 (N_28517,N_10289,N_11877);
and U28518 (N_28518,N_19760,N_18541);
nand U28519 (N_28519,N_17639,N_18211);
xor U28520 (N_28520,N_15362,N_17422);
and U28521 (N_28521,N_10839,N_10135);
xnor U28522 (N_28522,N_19093,N_18320);
nand U28523 (N_28523,N_13586,N_13848);
or U28524 (N_28524,N_14952,N_12615);
nand U28525 (N_28525,N_13133,N_17810);
xnor U28526 (N_28526,N_15388,N_13327);
nand U28527 (N_28527,N_14147,N_17139);
nand U28528 (N_28528,N_11297,N_18616);
nor U28529 (N_28529,N_13106,N_19738);
nor U28530 (N_28530,N_16993,N_10843);
nor U28531 (N_28531,N_17636,N_14482);
xor U28532 (N_28532,N_15349,N_11640);
and U28533 (N_28533,N_16242,N_19253);
nand U28534 (N_28534,N_13831,N_18873);
or U28535 (N_28535,N_14644,N_13864);
nor U28536 (N_28536,N_14846,N_17549);
or U28537 (N_28537,N_17445,N_12928);
nor U28538 (N_28538,N_16067,N_12097);
or U28539 (N_28539,N_16930,N_19817);
nor U28540 (N_28540,N_11032,N_19058);
nand U28541 (N_28541,N_11116,N_14402);
and U28542 (N_28542,N_13000,N_11363);
nor U28543 (N_28543,N_14071,N_14443);
xor U28544 (N_28544,N_13735,N_11096);
or U28545 (N_28545,N_18537,N_11809);
nand U28546 (N_28546,N_18860,N_16517);
or U28547 (N_28547,N_12402,N_12592);
nor U28548 (N_28548,N_16757,N_11209);
and U28549 (N_28549,N_17934,N_14700);
or U28550 (N_28550,N_13093,N_13613);
and U28551 (N_28551,N_12514,N_16586);
and U28552 (N_28552,N_12145,N_12031);
nor U28553 (N_28553,N_12166,N_13682);
nor U28554 (N_28554,N_11512,N_19260);
nand U28555 (N_28555,N_17808,N_19876);
nand U28556 (N_28556,N_19315,N_18508);
xor U28557 (N_28557,N_19688,N_18107);
xor U28558 (N_28558,N_14896,N_18410);
nand U28559 (N_28559,N_15504,N_16020);
or U28560 (N_28560,N_16397,N_15870);
nor U28561 (N_28561,N_10653,N_15275);
xor U28562 (N_28562,N_10983,N_18381);
or U28563 (N_28563,N_14316,N_13936);
nor U28564 (N_28564,N_17102,N_11299);
nor U28565 (N_28565,N_18522,N_17217);
nor U28566 (N_28566,N_17552,N_12597);
nand U28567 (N_28567,N_12417,N_19944);
nand U28568 (N_28568,N_11351,N_18100);
xor U28569 (N_28569,N_14837,N_17158);
and U28570 (N_28570,N_10482,N_14527);
or U28571 (N_28571,N_10838,N_10069);
xor U28572 (N_28572,N_12792,N_19818);
xor U28573 (N_28573,N_16466,N_19579);
or U28574 (N_28574,N_18324,N_18918);
xnor U28575 (N_28575,N_12338,N_17344);
nand U28576 (N_28576,N_12339,N_12187);
nor U28577 (N_28577,N_10355,N_12633);
and U28578 (N_28578,N_17324,N_15769);
nand U28579 (N_28579,N_13985,N_16999);
or U28580 (N_28580,N_15828,N_15862);
or U28581 (N_28581,N_17367,N_10689);
nand U28582 (N_28582,N_15661,N_17791);
xnor U28583 (N_28583,N_15433,N_10823);
nand U28584 (N_28584,N_14246,N_19628);
or U28585 (N_28585,N_12149,N_14722);
and U28586 (N_28586,N_14647,N_19650);
xnor U28587 (N_28587,N_18847,N_15031);
xor U28588 (N_28588,N_10466,N_15307);
nand U28589 (N_28589,N_18305,N_12077);
nand U28590 (N_28590,N_16345,N_12700);
nor U28591 (N_28591,N_11806,N_10208);
and U28592 (N_28592,N_15349,N_14156);
nand U28593 (N_28593,N_19453,N_17295);
nor U28594 (N_28594,N_10962,N_13006);
nor U28595 (N_28595,N_13602,N_12627);
nor U28596 (N_28596,N_11323,N_15833);
nand U28597 (N_28597,N_15977,N_18684);
nand U28598 (N_28598,N_14006,N_11011);
nor U28599 (N_28599,N_17034,N_19282);
and U28600 (N_28600,N_12195,N_17434);
nand U28601 (N_28601,N_10279,N_15249);
xnor U28602 (N_28602,N_16379,N_18695);
and U28603 (N_28603,N_11345,N_10360);
and U28604 (N_28604,N_13104,N_18037);
nand U28605 (N_28605,N_12851,N_15902);
nor U28606 (N_28606,N_18136,N_11120);
and U28607 (N_28607,N_12718,N_15471);
or U28608 (N_28608,N_15533,N_13711);
nand U28609 (N_28609,N_14302,N_16350);
xnor U28610 (N_28610,N_15677,N_11241);
or U28611 (N_28611,N_16171,N_18405);
or U28612 (N_28612,N_11322,N_10491);
or U28613 (N_28613,N_19854,N_12341);
nor U28614 (N_28614,N_16977,N_17680);
and U28615 (N_28615,N_18936,N_16365);
nand U28616 (N_28616,N_13429,N_14296);
or U28617 (N_28617,N_10790,N_14407);
and U28618 (N_28618,N_18499,N_11496);
xnor U28619 (N_28619,N_15237,N_11798);
or U28620 (N_28620,N_12137,N_16523);
xnor U28621 (N_28621,N_17750,N_11862);
and U28622 (N_28622,N_15281,N_14068);
nand U28623 (N_28623,N_16778,N_13726);
and U28624 (N_28624,N_19867,N_14055);
nor U28625 (N_28625,N_17467,N_16391);
nand U28626 (N_28626,N_13553,N_13021);
and U28627 (N_28627,N_12661,N_14575);
nand U28628 (N_28628,N_12875,N_15902);
or U28629 (N_28629,N_13061,N_14319);
nor U28630 (N_28630,N_11030,N_13268);
and U28631 (N_28631,N_12183,N_10438);
or U28632 (N_28632,N_11818,N_15258);
or U28633 (N_28633,N_19602,N_17907);
nand U28634 (N_28634,N_18373,N_18032);
xor U28635 (N_28635,N_17865,N_13964);
nand U28636 (N_28636,N_15736,N_12167);
nor U28637 (N_28637,N_17315,N_12817);
and U28638 (N_28638,N_15859,N_17108);
and U28639 (N_28639,N_18721,N_11670);
or U28640 (N_28640,N_17297,N_11500);
or U28641 (N_28641,N_14791,N_18980);
xnor U28642 (N_28642,N_18849,N_18970);
and U28643 (N_28643,N_19488,N_13358);
and U28644 (N_28644,N_13622,N_17458);
and U28645 (N_28645,N_10824,N_12433);
nor U28646 (N_28646,N_19588,N_16134);
nor U28647 (N_28647,N_12394,N_12163);
nand U28648 (N_28648,N_15630,N_11670);
nor U28649 (N_28649,N_14883,N_18565);
nor U28650 (N_28650,N_14571,N_10705);
xor U28651 (N_28651,N_17228,N_11331);
nand U28652 (N_28652,N_14104,N_13715);
or U28653 (N_28653,N_16540,N_11038);
xor U28654 (N_28654,N_18090,N_16516);
nor U28655 (N_28655,N_11235,N_11686);
nor U28656 (N_28656,N_12785,N_18138);
or U28657 (N_28657,N_17448,N_12831);
and U28658 (N_28658,N_16678,N_19294);
nand U28659 (N_28659,N_14342,N_16016);
nor U28660 (N_28660,N_14185,N_13618);
or U28661 (N_28661,N_10872,N_14091);
and U28662 (N_28662,N_12534,N_15560);
nand U28663 (N_28663,N_12061,N_19741);
nor U28664 (N_28664,N_16638,N_17230);
nor U28665 (N_28665,N_12905,N_13490);
xor U28666 (N_28666,N_12894,N_16353);
nand U28667 (N_28667,N_15877,N_18809);
nand U28668 (N_28668,N_10861,N_19788);
nor U28669 (N_28669,N_13660,N_10073);
or U28670 (N_28670,N_14919,N_19831);
nor U28671 (N_28671,N_10322,N_14746);
xnor U28672 (N_28672,N_15475,N_13437);
nor U28673 (N_28673,N_13207,N_15350);
nor U28674 (N_28674,N_17621,N_14692);
nand U28675 (N_28675,N_12780,N_15726);
nor U28676 (N_28676,N_18924,N_16309);
nor U28677 (N_28677,N_16393,N_12258);
and U28678 (N_28678,N_17004,N_16265);
or U28679 (N_28679,N_14047,N_16714);
or U28680 (N_28680,N_16625,N_12762);
xor U28681 (N_28681,N_13665,N_10678);
xnor U28682 (N_28682,N_12488,N_15026);
nor U28683 (N_28683,N_11560,N_17248);
or U28684 (N_28684,N_19672,N_14216);
or U28685 (N_28685,N_17928,N_10746);
nand U28686 (N_28686,N_11201,N_15244);
nand U28687 (N_28687,N_11560,N_19203);
and U28688 (N_28688,N_11741,N_11046);
or U28689 (N_28689,N_14674,N_11127);
nand U28690 (N_28690,N_14812,N_14784);
xnor U28691 (N_28691,N_12664,N_19379);
xnor U28692 (N_28692,N_12223,N_17154);
nand U28693 (N_28693,N_12288,N_10027);
or U28694 (N_28694,N_17611,N_14421);
nand U28695 (N_28695,N_12631,N_18473);
xnor U28696 (N_28696,N_11970,N_16618);
nor U28697 (N_28697,N_11261,N_16305);
xor U28698 (N_28698,N_17629,N_15628);
nand U28699 (N_28699,N_18455,N_17045);
nand U28700 (N_28700,N_19966,N_12759);
or U28701 (N_28701,N_10722,N_14069);
or U28702 (N_28702,N_14175,N_10343);
xnor U28703 (N_28703,N_12711,N_19852);
xnor U28704 (N_28704,N_19444,N_14292);
nand U28705 (N_28705,N_18133,N_16267);
or U28706 (N_28706,N_17025,N_11103);
nand U28707 (N_28707,N_10973,N_12066);
nor U28708 (N_28708,N_19989,N_12943);
nand U28709 (N_28709,N_17211,N_12319);
and U28710 (N_28710,N_14287,N_18564);
nor U28711 (N_28711,N_19839,N_13401);
and U28712 (N_28712,N_14516,N_18598);
nand U28713 (N_28713,N_15156,N_19100);
nand U28714 (N_28714,N_14042,N_11821);
or U28715 (N_28715,N_11726,N_16235);
and U28716 (N_28716,N_19065,N_11220);
xnor U28717 (N_28717,N_15619,N_15806);
xor U28718 (N_28718,N_19217,N_15263);
and U28719 (N_28719,N_13636,N_11025);
or U28720 (N_28720,N_14441,N_10905);
and U28721 (N_28721,N_15084,N_19466);
nor U28722 (N_28722,N_19814,N_13735);
nand U28723 (N_28723,N_18761,N_11962);
nand U28724 (N_28724,N_14400,N_10178);
nand U28725 (N_28725,N_10171,N_11789);
nor U28726 (N_28726,N_15578,N_15369);
xnor U28727 (N_28727,N_19541,N_12676);
nor U28728 (N_28728,N_11763,N_15136);
and U28729 (N_28729,N_15800,N_13658);
nand U28730 (N_28730,N_11986,N_12716);
and U28731 (N_28731,N_19246,N_11938);
nor U28732 (N_28732,N_17590,N_13923);
nor U28733 (N_28733,N_13388,N_18551);
xor U28734 (N_28734,N_10101,N_10290);
xor U28735 (N_28735,N_15787,N_14032);
and U28736 (N_28736,N_15630,N_17545);
xor U28737 (N_28737,N_14992,N_13440);
and U28738 (N_28738,N_15691,N_17577);
nand U28739 (N_28739,N_16226,N_13041);
nor U28740 (N_28740,N_18469,N_16334);
or U28741 (N_28741,N_17106,N_12977);
and U28742 (N_28742,N_10131,N_12356);
xnor U28743 (N_28743,N_16040,N_11929);
nand U28744 (N_28744,N_16089,N_17056);
and U28745 (N_28745,N_16419,N_15209);
and U28746 (N_28746,N_17879,N_15364);
and U28747 (N_28747,N_11827,N_11165);
or U28748 (N_28748,N_10722,N_18773);
or U28749 (N_28749,N_17747,N_15348);
or U28750 (N_28750,N_12863,N_12900);
and U28751 (N_28751,N_18867,N_18431);
or U28752 (N_28752,N_10602,N_14666);
xor U28753 (N_28753,N_11372,N_17415);
or U28754 (N_28754,N_13677,N_11868);
nand U28755 (N_28755,N_15305,N_17801);
nor U28756 (N_28756,N_12736,N_16501);
nor U28757 (N_28757,N_16481,N_18722);
nand U28758 (N_28758,N_17320,N_11997);
and U28759 (N_28759,N_11498,N_11599);
and U28760 (N_28760,N_18107,N_10118);
xor U28761 (N_28761,N_15171,N_13796);
and U28762 (N_28762,N_19457,N_16053);
xor U28763 (N_28763,N_12726,N_16218);
or U28764 (N_28764,N_11049,N_19751);
nand U28765 (N_28765,N_10184,N_19090);
xnor U28766 (N_28766,N_10988,N_16384);
or U28767 (N_28767,N_12979,N_10219);
nor U28768 (N_28768,N_12746,N_14473);
nor U28769 (N_28769,N_10036,N_16753);
nor U28770 (N_28770,N_17736,N_15282);
nor U28771 (N_28771,N_13845,N_17634);
and U28772 (N_28772,N_10217,N_13947);
and U28773 (N_28773,N_13343,N_18183);
and U28774 (N_28774,N_12123,N_16644);
nand U28775 (N_28775,N_10567,N_17137);
nand U28776 (N_28776,N_11760,N_19610);
or U28777 (N_28777,N_18471,N_16180);
xnor U28778 (N_28778,N_11864,N_11580);
or U28779 (N_28779,N_16036,N_19545);
or U28780 (N_28780,N_13958,N_15829);
or U28781 (N_28781,N_16311,N_16690);
nand U28782 (N_28782,N_11663,N_18615);
or U28783 (N_28783,N_14298,N_14623);
or U28784 (N_28784,N_17521,N_14979);
xnor U28785 (N_28785,N_18506,N_18389);
and U28786 (N_28786,N_18890,N_14579);
nor U28787 (N_28787,N_11306,N_18088);
nand U28788 (N_28788,N_18093,N_11004);
xor U28789 (N_28789,N_19203,N_18402);
nand U28790 (N_28790,N_17225,N_18826);
nand U28791 (N_28791,N_19462,N_18620);
nor U28792 (N_28792,N_11941,N_12318);
xnor U28793 (N_28793,N_10851,N_14363);
and U28794 (N_28794,N_16950,N_14582);
and U28795 (N_28795,N_16801,N_16945);
or U28796 (N_28796,N_17996,N_12058);
xor U28797 (N_28797,N_13120,N_19583);
xor U28798 (N_28798,N_17252,N_11773);
or U28799 (N_28799,N_18272,N_12936);
and U28800 (N_28800,N_11073,N_10824);
xnor U28801 (N_28801,N_12370,N_13351);
nand U28802 (N_28802,N_10820,N_13049);
nor U28803 (N_28803,N_10876,N_15381);
nor U28804 (N_28804,N_15167,N_15265);
nand U28805 (N_28805,N_14483,N_18449);
nor U28806 (N_28806,N_16895,N_10478);
or U28807 (N_28807,N_18081,N_16200);
and U28808 (N_28808,N_10769,N_10411);
or U28809 (N_28809,N_19722,N_19584);
xnor U28810 (N_28810,N_13545,N_18948);
or U28811 (N_28811,N_14147,N_12486);
and U28812 (N_28812,N_19857,N_14263);
or U28813 (N_28813,N_19709,N_15925);
xnor U28814 (N_28814,N_12496,N_10708);
nand U28815 (N_28815,N_17737,N_17226);
or U28816 (N_28816,N_12022,N_14382);
nand U28817 (N_28817,N_19583,N_15977);
and U28818 (N_28818,N_19710,N_13983);
xnor U28819 (N_28819,N_16834,N_15237);
nand U28820 (N_28820,N_10159,N_19997);
nor U28821 (N_28821,N_16605,N_14655);
or U28822 (N_28822,N_12872,N_16627);
or U28823 (N_28823,N_16073,N_14004);
or U28824 (N_28824,N_17986,N_15589);
xnor U28825 (N_28825,N_16142,N_12168);
nand U28826 (N_28826,N_12708,N_19110);
or U28827 (N_28827,N_15295,N_19388);
nand U28828 (N_28828,N_18802,N_13032);
nor U28829 (N_28829,N_12152,N_14467);
or U28830 (N_28830,N_16894,N_18742);
nand U28831 (N_28831,N_19187,N_13418);
nor U28832 (N_28832,N_11386,N_15239);
and U28833 (N_28833,N_17030,N_16558);
and U28834 (N_28834,N_16924,N_10511);
and U28835 (N_28835,N_19774,N_15215);
and U28836 (N_28836,N_16085,N_13626);
and U28837 (N_28837,N_18476,N_14345);
xor U28838 (N_28838,N_17687,N_17782);
xnor U28839 (N_28839,N_14119,N_14343);
nor U28840 (N_28840,N_17081,N_11565);
nand U28841 (N_28841,N_15111,N_18671);
and U28842 (N_28842,N_16085,N_13885);
or U28843 (N_28843,N_10294,N_13856);
nand U28844 (N_28844,N_13392,N_18399);
and U28845 (N_28845,N_17532,N_12283);
or U28846 (N_28846,N_18740,N_10808);
nand U28847 (N_28847,N_11291,N_18749);
nand U28848 (N_28848,N_18713,N_14186);
nor U28849 (N_28849,N_11041,N_10722);
and U28850 (N_28850,N_16272,N_17007);
xnor U28851 (N_28851,N_15692,N_13373);
or U28852 (N_28852,N_17303,N_14632);
and U28853 (N_28853,N_16980,N_16237);
nor U28854 (N_28854,N_19243,N_14982);
nor U28855 (N_28855,N_19201,N_11395);
xnor U28856 (N_28856,N_15250,N_16941);
nand U28857 (N_28857,N_14147,N_18533);
and U28858 (N_28858,N_10063,N_11025);
and U28859 (N_28859,N_13000,N_17471);
and U28860 (N_28860,N_11166,N_16597);
nor U28861 (N_28861,N_14870,N_13785);
nand U28862 (N_28862,N_14452,N_12617);
or U28863 (N_28863,N_19886,N_17574);
or U28864 (N_28864,N_14888,N_15514);
nand U28865 (N_28865,N_15222,N_15265);
or U28866 (N_28866,N_11697,N_19454);
nor U28867 (N_28867,N_14216,N_18607);
or U28868 (N_28868,N_13756,N_18877);
xnor U28869 (N_28869,N_11303,N_10697);
nand U28870 (N_28870,N_17168,N_10515);
xor U28871 (N_28871,N_18042,N_16225);
nand U28872 (N_28872,N_19483,N_18983);
or U28873 (N_28873,N_14330,N_16878);
nand U28874 (N_28874,N_18564,N_12122);
xnor U28875 (N_28875,N_17287,N_11795);
nand U28876 (N_28876,N_11492,N_16111);
or U28877 (N_28877,N_15115,N_16212);
xor U28878 (N_28878,N_18207,N_12745);
xnor U28879 (N_28879,N_11888,N_18743);
nand U28880 (N_28880,N_19189,N_11190);
nor U28881 (N_28881,N_11898,N_13924);
nor U28882 (N_28882,N_14607,N_16674);
nand U28883 (N_28883,N_19475,N_15594);
and U28884 (N_28884,N_11723,N_19275);
nor U28885 (N_28885,N_17491,N_15887);
or U28886 (N_28886,N_17470,N_18395);
or U28887 (N_28887,N_14940,N_11265);
xor U28888 (N_28888,N_19747,N_11971);
or U28889 (N_28889,N_17266,N_18547);
and U28890 (N_28890,N_17671,N_12102);
nor U28891 (N_28891,N_15790,N_11474);
nor U28892 (N_28892,N_11451,N_19634);
and U28893 (N_28893,N_13251,N_13620);
and U28894 (N_28894,N_15596,N_16975);
xnor U28895 (N_28895,N_14633,N_17538);
or U28896 (N_28896,N_17938,N_10821);
or U28897 (N_28897,N_14000,N_11110);
and U28898 (N_28898,N_19362,N_11806);
nand U28899 (N_28899,N_15325,N_17576);
xnor U28900 (N_28900,N_18176,N_11169);
xor U28901 (N_28901,N_11017,N_14943);
xor U28902 (N_28902,N_11604,N_19771);
nor U28903 (N_28903,N_10741,N_13864);
nor U28904 (N_28904,N_15294,N_16713);
nor U28905 (N_28905,N_10574,N_18437);
nand U28906 (N_28906,N_14915,N_12623);
xnor U28907 (N_28907,N_11296,N_16098);
or U28908 (N_28908,N_15091,N_18341);
and U28909 (N_28909,N_17521,N_17424);
nand U28910 (N_28910,N_12626,N_16968);
nor U28911 (N_28911,N_19721,N_16525);
or U28912 (N_28912,N_12047,N_13617);
xnor U28913 (N_28913,N_19854,N_12040);
nand U28914 (N_28914,N_10551,N_15915);
nor U28915 (N_28915,N_13104,N_10050);
xor U28916 (N_28916,N_14759,N_10504);
nand U28917 (N_28917,N_11879,N_17898);
nor U28918 (N_28918,N_11668,N_10356);
nand U28919 (N_28919,N_19153,N_11194);
or U28920 (N_28920,N_12230,N_17775);
xnor U28921 (N_28921,N_13183,N_18769);
xor U28922 (N_28922,N_18024,N_11528);
and U28923 (N_28923,N_14712,N_19425);
and U28924 (N_28924,N_16646,N_12658);
or U28925 (N_28925,N_16140,N_13230);
and U28926 (N_28926,N_15847,N_17650);
nor U28927 (N_28927,N_17038,N_10420);
and U28928 (N_28928,N_18182,N_11094);
nor U28929 (N_28929,N_10690,N_15393);
nand U28930 (N_28930,N_14380,N_13767);
and U28931 (N_28931,N_15903,N_13706);
nor U28932 (N_28932,N_13809,N_18514);
nand U28933 (N_28933,N_13610,N_14699);
nor U28934 (N_28934,N_15637,N_11883);
and U28935 (N_28935,N_16397,N_12041);
and U28936 (N_28936,N_11412,N_14179);
nand U28937 (N_28937,N_17891,N_10304);
or U28938 (N_28938,N_14478,N_14733);
or U28939 (N_28939,N_15292,N_16802);
nand U28940 (N_28940,N_10109,N_18891);
nand U28941 (N_28941,N_19974,N_18042);
xnor U28942 (N_28942,N_16254,N_12845);
nand U28943 (N_28943,N_15239,N_12107);
xor U28944 (N_28944,N_10156,N_11217);
nor U28945 (N_28945,N_17404,N_16519);
nor U28946 (N_28946,N_18341,N_14588);
nor U28947 (N_28947,N_10067,N_14008);
xor U28948 (N_28948,N_10291,N_16027);
nand U28949 (N_28949,N_14125,N_10311);
or U28950 (N_28950,N_10106,N_13584);
nor U28951 (N_28951,N_12414,N_10672);
xor U28952 (N_28952,N_10856,N_11695);
and U28953 (N_28953,N_13841,N_14214);
and U28954 (N_28954,N_17606,N_13966);
nand U28955 (N_28955,N_15408,N_11670);
xor U28956 (N_28956,N_11839,N_15463);
nor U28957 (N_28957,N_13789,N_10627);
or U28958 (N_28958,N_12579,N_17816);
nor U28959 (N_28959,N_12020,N_11798);
xnor U28960 (N_28960,N_15796,N_11772);
and U28961 (N_28961,N_12421,N_19609);
nand U28962 (N_28962,N_11671,N_16791);
and U28963 (N_28963,N_16036,N_12307);
or U28964 (N_28964,N_13218,N_16920);
nor U28965 (N_28965,N_15391,N_10571);
nand U28966 (N_28966,N_18317,N_18432);
xor U28967 (N_28967,N_14526,N_18919);
and U28968 (N_28968,N_14260,N_11514);
or U28969 (N_28969,N_14299,N_10170);
and U28970 (N_28970,N_11668,N_12274);
xor U28971 (N_28971,N_11015,N_15609);
and U28972 (N_28972,N_18840,N_19030);
nor U28973 (N_28973,N_12839,N_10001);
xor U28974 (N_28974,N_14800,N_11024);
and U28975 (N_28975,N_18900,N_19173);
and U28976 (N_28976,N_18515,N_15374);
nor U28977 (N_28977,N_15723,N_19510);
and U28978 (N_28978,N_12434,N_11207);
nand U28979 (N_28979,N_12218,N_11580);
nand U28980 (N_28980,N_10629,N_15485);
and U28981 (N_28981,N_16736,N_10077);
xor U28982 (N_28982,N_17093,N_16177);
or U28983 (N_28983,N_12893,N_18433);
nand U28984 (N_28984,N_12449,N_17689);
nand U28985 (N_28985,N_17377,N_15304);
xnor U28986 (N_28986,N_13558,N_18912);
and U28987 (N_28987,N_12832,N_15862);
and U28988 (N_28988,N_11819,N_14462);
xnor U28989 (N_28989,N_14428,N_18966);
or U28990 (N_28990,N_15666,N_16165);
and U28991 (N_28991,N_13515,N_18079);
nor U28992 (N_28992,N_18291,N_18847);
xnor U28993 (N_28993,N_10733,N_12550);
xnor U28994 (N_28994,N_11672,N_16009);
nand U28995 (N_28995,N_14541,N_19218);
nor U28996 (N_28996,N_13083,N_10912);
nand U28997 (N_28997,N_18724,N_10772);
and U28998 (N_28998,N_18223,N_10631);
or U28999 (N_28999,N_10758,N_12106);
nand U29000 (N_29000,N_14165,N_11296);
or U29001 (N_29001,N_18093,N_13089);
nor U29002 (N_29002,N_18510,N_10091);
and U29003 (N_29003,N_11489,N_13177);
or U29004 (N_29004,N_11339,N_16233);
or U29005 (N_29005,N_19964,N_19276);
nor U29006 (N_29006,N_14589,N_16003);
nor U29007 (N_29007,N_17315,N_10294);
or U29008 (N_29008,N_19483,N_19096);
nor U29009 (N_29009,N_18263,N_14150);
or U29010 (N_29010,N_12593,N_18213);
xnor U29011 (N_29011,N_12091,N_17396);
and U29012 (N_29012,N_12885,N_17179);
nor U29013 (N_29013,N_11499,N_13017);
xnor U29014 (N_29014,N_11203,N_11464);
nor U29015 (N_29015,N_10020,N_11259);
nand U29016 (N_29016,N_17400,N_16821);
nand U29017 (N_29017,N_16345,N_12417);
and U29018 (N_29018,N_15113,N_16398);
nand U29019 (N_29019,N_11309,N_10755);
or U29020 (N_29020,N_17844,N_17187);
nor U29021 (N_29021,N_18252,N_19528);
nand U29022 (N_29022,N_18935,N_10952);
and U29023 (N_29023,N_17108,N_19590);
nand U29024 (N_29024,N_12816,N_12264);
or U29025 (N_29025,N_19810,N_15430);
and U29026 (N_29026,N_10721,N_10728);
and U29027 (N_29027,N_10774,N_18714);
nor U29028 (N_29028,N_12727,N_15389);
and U29029 (N_29029,N_17125,N_17881);
and U29030 (N_29030,N_13352,N_12665);
xor U29031 (N_29031,N_17803,N_19064);
or U29032 (N_29032,N_10859,N_18908);
or U29033 (N_29033,N_15432,N_14751);
and U29034 (N_29034,N_18724,N_16722);
and U29035 (N_29035,N_17468,N_17358);
xor U29036 (N_29036,N_19662,N_19997);
and U29037 (N_29037,N_10862,N_14037);
nand U29038 (N_29038,N_15315,N_11788);
and U29039 (N_29039,N_19037,N_11818);
nor U29040 (N_29040,N_16823,N_19049);
nor U29041 (N_29041,N_11518,N_17032);
or U29042 (N_29042,N_19138,N_10451);
or U29043 (N_29043,N_11816,N_18330);
or U29044 (N_29044,N_19212,N_18651);
nand U29045 (N_29045,N_15212,N_13810);
nand U29046 (N_29046,N_10889,N_14690);
nor U29047 (N_29047,N_19286,N_15042);
nand U29048 (N_29048,N_19094,N_10930);
xor U29049 (N_29049,N_14414,N_13242);
nand U29050 (N_29050,N_16904,N_18585);
or U29051 (N_29051,N_11570,N_19716);
nand U29052 (N_29052,N_18030,N_15714);
nor U29053 (N_29053,N_14631,N_10364);
nor U29054 (N_29054,N_17910,N_13288);
nand U29055 (N_29055,N_15680,N_10830);
nand U29056 (N_29056,N_15769,N_12145);
xnor U29057 (N_29057,N_16676,N_16176);
nor U29058 (N_29058,N_11542,N_13032);
xor U29059 (N_29059,N_18525,N_18744);
nor U29060 (N_29060,N_14695,N_16303);
and U29061 (N_29061,N_17420,N_15267);
and U29062 (N_29062,N_11633,N_15466);
nor U29063 (N_29063,N_16826,N_15396);
or U29064 (N_29064,N_14247,N_19812);
and U29065 (N_29065,N_16009,N_19925);
xor U29066 (N_29066,N_16800,N_14864);
or U29067 (N_29067,N_12212,N_15735);
nor U29068 (N_29068,N_15943,N_16783);
xor U29069 (N_29069,N_19220,N_15484);
nor U29070 (N_29070,N_17519,N_10847);
or U29071 (N_29071,N_10271,N_18107);
nand U29072 (N_29072,N_13381,N_19078);
and U29073 (N_29073,N_17889,N_16966);
and U29074 (N_29074,N_18260,N_11924);
nor U29075 (N_29075,N_19470,N_19707);
and U29076 (N_29076,N_13391,N_16312);
or U29077 (N_29077,N_15263,N_13785);
xor U29078 (N_29078,N_12811,N_15552);
and U29079 (N_29079,N_16672,N_15980);
nand U29080 (N_29080,N_16885,N_15296);
nand U29081 (N_29081,N_11514,N_12873);
xnor U29082 (N_29082,N_14950,N_18404);
and U29083 (N_29083,N_16149,N_15581);
nor U29084 (N_29084,N_12117,N_12090);
or U29085 (N_29085,N_10021,N_16362);
or U29086 (N_29086,N_17521,N_19227);
and U29087 (N_29087,N_12350,N_12253);
xor U29088 (N_29088,N_18102,N_10451);
nor U29089 (N_29089,N_15399,N_14485);
nor U29090 (N_29090,N_17523,N_13641);
or U29091 (N_29091,N_12346,N_18786);
nand U29092 (N_29092,N_18678,N_10172);
nor U29093 (N_29093,N_16778,N_15335);
and U29094 (N_29094,N_15522,N_13746);
nor U29095 (N_29095,N_17250,N_15464);
nand U29096 (N_29096,N_12284,N_18685);
xor U29097 (N_29097,N_19280,N_14027);
xor U29098 (N_29098,N_11513,N_15920);
nor U29099 (N_29099,N_14202,N_15560);
or U29100 (N_29100,N_10187,N_18626);
or U29101 (N_29101,N_17209,N_15524);
xnor U29102 (N_29102,N_18690,N_15113);
or U29103 (N_29103,N_18557,N_17115);
or U29104 (N_29104,N_10296,N_16796);
nor U29105 (N_29105,N_14088,N_10804);
and U29106 (N_29106,N_18465,N_11262);
nand U29107 (N_29107,N_18846,N_15807);
or U29108 (N_29108,N_15938,N_12608);
and U29109 (N_29109,N_13260,N_18897);
nand U29110 (N_29110,N_10579,N_10451);
xor U29111 (N_29111,N_14821,N_15820);
nand U29112 (N_29112,N_11107,N_15504);
nor U29113 (N_29113,N_19615,N_17036);
and U29114 (N_29114,N_11464,N_10840);
or U29115 (N_29115,N_15317,N_10915);
and U29116 (N_29116,N_12480,N_19113);
nand U29117 (N_29117,N_14427,N_16927);
nor U29118 (N_29118,N_11196,N_18858);
nand U29119 (N_29119,N_10079,N_16622);
nor U29120 (N_29120,N_12965,N_10800);
or U29121 (N_29121,N_11488,N_16145);
xnor U29122 (N_29122,N_17837,N_11561);
and U29123 (N_29123,N_15888,N_16704);
and U29124 (N_29124,N_18491,N_17261);
nand U29125 (N_29125,N_16761,N_17636);
nand U29126 (N_29126,N_12234,N_13065);
or U29127 (N_29127,N_10140,N_16960);
and U29128 (N_29128,N_17804,N_15652);
or U29129 (N_29129,N_17797,N_18348);
nand U29130 (N_29130,N_17259,N_15501);
and U29131 (N_29131,N_16453,N_18484);
nor U29132 (N_29132,N_14021,N_19475);
nor U29133 (N_29133,N_13656,N_14565);
nand U29134 (N_29134,N_16072,N_19663);
xor U29135 (N_29135,N_12812,N_17745);
xnor U29136 (N_29136,N_11036,N_17902);
and U29137 (N_29137,N_15493,N_12603);
xor U29138 (N_29138,N_10227,N_14333);
nor U29139 (N_29139,N_19804,N_14178);
and U29140 (N_29140,N_11378,N_13108);
or U29141 (N_29141,N_14321,N_19449);
nor U29142 (N_29142,N_14753,N_14002);
nand U29143 (N_29143,N_18884,N_16838);
xnor U29144 (N_29144,N_14578,N_18453);
nand U29145 (N_29145,N_19799,N_10596);
nand U29146 (N_29146,N_19639,N_10545);
and U29147 (N_29147,N_14426,N_18771);
nor U29148 (N_29148,N_10613,N_10418);
and U29149 (N_29149,N_17222,N_11551);
nand U29150 (N_29150,N_13061,N_14425);
xnor U29151 (N_29151,N_18508,N_19351);
or U29152 (N_29152,N_18135,N_18788);
xor U29153 (N_29153,N_12096,N_16232);
xnor U29154 (N_29154,N_10562,N_11719);
xnor U29155 (N_29155,N_12585,N_19681);
and U29156 (N_29156,N_12412,N_13579);
nor U29157 (N_29157,N_19936,N_17104);
nor U29158 (N_29158,N_11534,N_15590);
nor U29159 (N_29159,N_10985,N_19635);
and U29160 (N_29160,N_11823,N_17086);
nand U29161 (N_29161,N_14160,N_16891);
and U29162 (N_29162,N_10530,N_19735);
nor U29163 (N_29163,N_12511,N_13198);
or U29164 (N_29164,N_13883,N_19841);
nand U29165 (N_29165,N_17721,N_12049);
xnor U29166 (N_29166,N_13624,N_14640);
nand U29167 (N_29167,N_16574,N_11700);
xor U29168 (N_29168,N_12447,N_16922);
xnor U29169 (N_29169,N_15303,N_12944);
nor U29170 (N_29170,N_13349,N_11856);
xor U29171 (N_29171,N_15007,N_16897);
nand U29172 (N_29172,N_14851,N_11086);
nor U29173 (N_29173,N_10494,N_13010);
nor U29174 (N_29174,N_13547,N_16046);
or U29175 (N_29175,N_11336,N_19954);
xor U29176 (N_29176,N_19816,N_18167);
nor U29177 (N_29177,N_12048,N_19245);
xnor U29178 (N_29178,N_14612,N_14161);
nor U29179 (N_29179,N_15837,N_19603);
and U29180 (N_29180,N_13030,N_15564);
and U29181 (N_29181,N_16030,N_15075);
xnor U29182 (N_29182,N_14598,N_10705);
and U29183 (N_29183,N_18215,N_18751);
and U29184 (N_29184,N_15555,N_14585);
nand U29185 (N_29185,N_19277,N_13213);
and U29186 (N_29186,N_15787,N_14660);
xnor U29187 (N_29187,N_13415,N_13509);
or U29188 (N_29188,N_16155,N_15571);
xor U29189 (N_29189,N_15227,N_11138);
xor U29190 (N_29190,N_12001,N_10246);
xnor U29191 (N_29191,N_19596,N_14730);
and U29192 (N_29192,N_18344,N_13048);
nor U29193 (N_29193,N_19481,N_17060);
or U29194 (N_29194,N_13704,N_13426);
nand U29195 (N_29195,N_10072,N_12630);
nor U29196 (N_29196,N_16282,N_18025);
nand U29197 (N_29197,N_16571,N_15660);
nor U29198 (N_29198,N_18026,N_19302);
nor U29199 (N_29199,N_13220,N_16941);
nand U29200 (N_29200,N_17886,N_13669);
and U29201 (N_29201,N_19135,N_16856);
xnor U29202 (N_29202,N_17662,N_16147);
and U29203 (N_29203,N_17957,N_18849);
and U29204 (N_29204,N_16986,N_16048);
and U29205 (N_29205,N_15318,N_18368);
or U29206 (N_29206,N_18537,N_13142);
nand U29207 (N_29207,N_11126,N_17843);
and U29208 (N_29208,N_12350,N_12078);
xor U29209 (N_29209,N_10401,N_13918);
and U29210 (N_29210,N_13517,N_18814);
and U29211 (N_29211,N_13305,N_18680);
xor U29212 (N_29212,N_14941,N_15191);
nor U29213 (N_29213,N_12359,N_15832);
nor U29214 (N_29214,N_13842,N_10756);
and U29215 (N_29215,N_18484,N_15778);
and U29216 (N_29216,N_16894,N_11639);
or U29217 (N_29217,N_19759,N_14625);
nand U29218 (N_29218,N_17464,N_10801);
nand U29219 (N_29219,N_10539,N_13399);
or U29220 (N_29220,N_12523,N_16662);
and U29221 (N_29221,N_16345,N_16878);
nand U29222 (N_29222,N_17971,N_12420);
nand U29223 (N_29223,N_16272,N_11537);
and U29224 (N_29224,N_13218,N_14064);
xnor U29225 (N_29225,N_19204,N_16352);
or U29226 (N_29226,N_15522,N_14081);
xor U29227 (N_29227,N_16466,N_11122);
xor U29228 (N_29228,N_16289,N_11754);
nor U29229 (N_29229,N_11726,N_17526);
xnor U29230 (N_29230,N_15600,N_11998);
and U29231 (N_29231,N_19932,N_17030);
or U29232 (N_29232,N_12158,N_18109);
nand U29233 (N_29233,N_14517,N_11394);
and U29234 (N_29234,N_12819,N_16930);
xnor U29235 (N_29235,N_13535,N_10826);
nor U29236 (N_29236,N_19948,N_14378);
or U29237 (N_29237,N_19879,N_10790);
or U29238 (N_29238,N_13012,N_14741);
xor U29239 (N_29239,N_13940,N_17164);
nor U29240 (N_29240,N_12506,N_16952);
nand U29241 (N_29241,N_12138,N_19190);
nor U29242 (N_29242,N_19780,N_16424);
nor U29243 (N_29243,N_12477,N_13624);
nor U29244 (N_29244,N_17755,N_14489);
xnor U29245 (N_29245,N_16870,N_10973);
nor U29246 (N_29246,N_19552,N_12059);
and U29247 (N_29247,N_15209,N_14294);
or U29248 (N_29248,N_13516,N_18633);
nand U29249 (N_29249,N_11875,N_16858);
and U29250 (N_29250,N_16559,N_18435);
nor U29251 (N_29251,N_13128,N_19577);
or U29252 (N_29252,N_19473,N_10415);
nor U29253 (N_29253,N_16125,N_11011);
nor U29254 (N_29254,N_14812,N_14146);
xor U29255 (N_29255,N_12723,N_16781);
and U29256 (N_29256,N_16555,N_13134);
or U29257 (N_29257,N_13978,N_16637);
nand U29258 (N_29258,N_17667,N_11111);
or U29259 (N_29259,N_10679,N_14994);
nand U29260 (N_29260,N_10964,N_19076);
xor U29261 (N_29261,N_18400,N_12091);
or U29262 (N_29262,N_15321,N_13523);
nor U29263 (N_29263,N_14919,N_14666);
or U29264 (N_29264,N_19084,N_15755);
or U29265 (N_29265,N_19338,N_15645);
nand U29266 (N_29266,N_16255,N_17855);
or U29267 (N_29267,N_18676,N_18022);
nor U29268 (N_29268,N_10446,N_12135);
and U29269 (N_29269,N_18157,N_12936);
xnor U29270 (N_29270,N_12873,N_18698);
nor U29271 (N_29271,N_13285,N_10196);
nand U29272 (N_29272,N_19209,N_11857);
xnor U29273 (N_29273,N_11632,N_11038);
and U29274 (N_29274,N_16651,N_12389);
nand U29275 (N_29275,N_12514,N_18956);
xor U29276 (N_29276,N_19941,N_16461);
xnor U29277 (N_29277,N_14716,N_12250);
nor U29278 (N_29278,N_17024,N_17287);
and U29279 (N_29279,N_11243,N_13476);
or U29280 (N_29280,N_17708,N_13675);
or U29281 (N_29281,N_15488,N_15044);
and U29282 (N_29282,N_13026,N_14832);
nor U29283 (N_29283,N_14022,N_12819);
nor U29284 (N_29284,N_13991,N_18920);
or U29285 (N_29285,N_17827,N_18442);
nand U29286 (N_29286,N_14671,N_13089);
xor U29287 (N_29287,N_10737,N_10114);
nor U29288 (N_29288,N_13635,N_19952);
or U29289 (N_29289,N_15556,N_19988);
nand U29290 (N_29290,N_11278,N_19381);
nor U29291 (N_29291,N_12516,N_13488);
and U29292 (N_29292,N_10968,N_18334);
and U29293 (N_29293,N_18745,N_14106);
nor U29294 (N_29294,N_16791,N_14805);
or U29295 (N_29295,N_11078,N_10966);
nand U29296 (N_29296,N_18029,N_11279);
nand U29297 (N_29297,N_19649,N_12560);
and U29298 (N_29298,N_13673,N_10183);
xnor U29299 (N_29299,N_16314,N_16579);
or U29300 (N_29300,N_19502,N_15213);
xnor U29301 (N_29301,N_16356,N_11162);
xor U29302 (N_29302,N_18497,N_18420);
and U29303 (N_29303,N_12577,N_14091);
nor U29304 (N_29304,N_12125,N_12269);
nand U29305 (N_29305,N_10007,N_13378);
xnor U29306 (N_29306,N_18519,N_15679);
or U29307 (N_29307,N_13909,N_19393);
nand U29308 (N_29308,N_16532,N_17771);
and U29309 (N_29309,N_15046,N_11413);
xor U29310 (N_29310,N_11162,N_16918);
and U29311 (N_29311,N_16687,N_11510);
and U29312 (N_29312,N_11745,N_18618);
nand U29313 (N_29313,N_10279,N_18628);
or U29314 (N_29314,N_14976,N_11084);
nand U29315 (N_29315,N_17961,N_12161);
nor U29316 (N_29316,N_18783,N_11335);
or U29317 (N_29317,N_16983,N_16159);
nor U29318 (N_29318,N_11297,N_15141);
nand U29319 (N_29319,N_14377,N_19537);
and U29320 (N_29320,N_15744,N_18667);
nor U29321 (N_29321,N_15444,N_18813);
xnor U29322 (N_29322,N_17145,N_11647);
and U29323 (N_29323,N_18762,N_14701);
nor U29324 (N_29324,N_13302,N_18802);
and U29325 (N_29325,N_16694,N_19460);
nand U29326 (N_29326,N_16924,N_19532);
or U29327 (N_29327,N_18141,N_11415);
and U29328 (N_29328,N_15382,N_18914);
nand U29329 (N_29329,N_17842,N_19485);
xor U29330 (N_29330,N_15036,N_12789);
or U29331 (N_29331,N_18745,N_16381);
or U29332 (N_29332,N_19383,N_17706);
or U29333 (N_29333,N_10175,N_17808);
nor U29334 (N_29334,N_17484,N_19952);
or U29335 (N_29335,N_15553,N_12774);
nor U29336 (N_29336,N_12848,N_18665);
or U29337 (N_29337,N_14603,N_12970);
and U29338 (N_29338,N_18185,N_11230);
and U29339 (N_29339,N_16008,N_13458);
and U29340 (N_29340,N_16673,N_19043);
nor U29341 (N_29341,N_12033,N_12483);
nand U29342 (N_29342,N_10101,N_16360);
nor U29343 (N_29343,N_17127,N_17354);
nand U29344 (N_29344,N_12594,N_13271);
and U29345 (N_29345,N_19343,N_12838);
nor U29346 (N_29346,N_14197,N_16067);
or U29347 (N_29347,N_10809,N_11923);
nor U29348 (N_29348,N_14312,N_13777);
nand U29349 (N_29349,N_12956,N_13942);
nand U29350 (N_29350,N_18519,N_13350);
nand U29351 (N_29351,N_17898,N_18844);
nor U29352 (N_29352,N_10744,N_17925);
nand U29353 (N_29353,N_14003,N_19055);
xor U29354 (N_29354,N_12866,N_10406);
or U29355 (N_29355,N_18232,N_19671);
nor U29356 (N_29356,N_18267,N_10437);
or U29357 (N_29357,N_19353,N_10030);
xnor U29358 (N_29358,N_16714,N_14831);
nor U29359 (N_29359,N_11183,N_10182);
xnor U29360 (N_29360,N_12861,N_17460);
nand U29361 (N_29361,N_14879,N_11623);
and U29362 (N_29362,N_13773,N_17081);
xor U29363 (N_29363,N_12492,N_17599);
nor U29364 (N_29364,N_19593,N_15605);
nand U29365 (N_29365,N_15170,N_14216);
or U29366 (N_29366,N_10473,N_10380);
xnor U29367 (N_29367,N_13017,N_15899);
or U29368 (N_29368,N_13248,N_16619);
xor U29369 (N_29369,N_14359,N_13240);
xnor U29370 (N_29370,N_13914,N_14495);
xnor U29371 (N_29371,N_17634,N_19712);
or U29372 (N_29372,N_12794,N_18122);
and U29373 (N_29373,N_15490,N_12954);
nor U29374 (N_29374,N_18723,N_10474);
nor U29375 (N_29375,N_11601,N_19166);
or U29376 (N_29376,N_15325,N_19788);
nor U29377 (N_29377,N_17125,N_12727);
nor U29378 (N_29378,N_19965,N_14389);
and U29379 (N_29379,N_19707,N_14761);
nand U29380 (N_29380,N_17756,N_10199);
nor U29381 (N_29381,N_15241,N_18086);
and U29382 (N_29382,N_13992,N_17218);
or U29383 (N_29383,N_10567,N_17915);
or U29384 (N_29384,N_11665,N_16866);
and U29385 (N_29385,N_12125,N_16270);
nor U29386 (N_29386,N_16921,N_10783);
or U29387 (N_29387,N_18184,N_17345);
nor U29388 (N_29388,N_19785,N_11297);
or U29389 (N_29389,N_14448,N_10317);
nand U29390 (N_29390,N_16525,N_19659);
or U29391 (N_29391,N_15096,N_16158);
nand U29392 (N_29392,N_13263,N_15163);
nand U29393 (N_29393,N_15137,N_15228);
nand U29394 (N_29394,N_11752,N_17626);
or U29395 (N_29395,N_10004,N_13855);
nand U29396 (N_29396,N_18666,N_10428);
and U29397 (N_29397,N_10680,N_11426);
xor U29398 (N_29398,N_17870,N_19746);
or U29399 (N_29399,N_16554,N_17411);
nand U29400 (N_29400,N_12424,N_18231);
nand U29401 (N_29401,N_17243,N_12875);
nand U29402 (N_29402,N_13448,N_13768);
or U29403 (N_29403,N_14846,N_14814);
or U29404 (N_29404,N_13496,N_17082);
and U29405 (N_29405,N_10382,N_16664);
nor U29406 (N_29406,N_13230,N_19181);
nor U29407 (N_29407,N_13420,N_17757);
or U29408 (N_29408,N_18561,N_14251);
nand U29409 (N_29409,N_17714,N_11386);
and U29410 (N_29410,N_10951,N_19365);
or U29411 (N_29411,N_14824,N_14672);
and U29412 (N_29412,N_19665,N_13108);
nand U29413 (N_29413,N_16622,N_11182);
or U29414 (N_29414,N_17852,N_12218);
nor U29415 (N_29415,N_14551,N_16126);
and U29416 (N_29416,N_11652,N_17212);
and U29417 (N_29417,N_14288,N_10963);
or U29418 (N_29418,N_18026,N_12485);
or U29419 (N_29419,N_10889,N_14282);
and U29420 (N_29420,N_12819,N_13388);
nand U29421 (N_29421,N_17319,N_17245);
nand U29422 (N_29422,N_11439,N_12907);
xnor U29423 (N_29423,N_10970,N_14080);
xor U29424 (N_29424,N_11461,N_19103);
xnor U29425 (N_29425,N_18715,N_11051);
nor U29426 (N_29426,N_11104,N_15449);
xor U29427 (N_29427,N_17574,N_12749);
nor U29428 (N_29428,N_19440,N_11054);
xnor U29429 (N_29429,N_11575,N_17867);
and U29430 (N_29430,N_16856,N_10554);
xnor U29431 (N_29431,N_12725,N_12865);
or U29432 (N_29432,N_19130,N_17733);
and U29433 (N_29433,N_10300,N_13258);
or U29434 (N_29434,N_17530,N_12653);
xor U29435 (N_29435,N_10888,N_16803);
xor U29436 (N_29436,N_16163,N_19119);
nor U29437 (N_29437,N_15556,N_18124);
or U29438 (N_29438,N_11765,N_14408);
and U29439 (N_29439,N_19682,N_11736);
and U29440 (N_29440,N_14813,N_13939);
xnor U29441 (N_29441,N_13891,N_16770);
nor U29442 (N_29442,N_18978,N_19143);
nand U29443 (N_29443,N_12617,N_14513);
nand U29444 (N_29444,N_16222,N_10793);
and U29445 (N_29445,N_12667,N_15042);
or U29446 (N_29446,N_11072,N_16622);
or U29447 (N_29447,N_19936,N_15283);
nor U29448 (N_29448,N_14150,N_14840);
or U29449 (N_29449,N_16153,N_12899);
xnor U29450 (N_29450,N_12827,N_17856);
xnor U29451 (N_29451,N_13652,N_16036);
nor U29452 (N_29452,N_12168,N_10503);
nor U29453 (N_29453,N_11565,N_16621);
xor U29454 (N_29454,N_18576,N_18433);
or U29455 (N_29455,N_19882,N_12607);
and U29456 (N_29456,N_17084,N_14915);
or U29457 (N_29457,N_17766,N_16783);
xnor U29458 (N_29458,N_19162,N_18968);
xor U29459 (N_29459,N_13687,N_10307);
xor U29460 (N_29460,N_17171,N_12897);
or U29461 (N_29461,N_13375,N_14986);
nand U29462 (N_29462,N_14266,N_11180);
xor U29463 (N_29463,N_16100,N_14598);
and U29464 (N_29464,N_19916,N_10793);
nand U29465 (N_29465,N_14762,N_14806);
nand U29466 (N_29466,N_15355,N_12101);
nor U29467 (N_29467,N_17983,N_15560);
nand U29468 (N_29468,N_16447,N_14911);
or U29469 (N_29469,N_16498,N_11003);
nand U29470 (N_29470,N_18746,N_19982);
nand U29471 (N_29471,N_12153,N_15624);
nand U29472 (N_29472,N_16431,N_11390);
xor U29473 (N_29473,N_13178,N_13226);
xnor U29474 (N_29474,N_13729,N_12125);
nor U29475 (N_29475,N_18665,N_16798);
nand U29476 (N_29476,N_13276,N_10561);
or U29477 (N_29477,N_17969,N_10298);
xor U29478 (N_29478,N_12818,N_17090);
nand U29479 (N_29479,N_19893,N_12766);
or U29480 (N_29480,N_11431,N_11781);
nand U29481 (N_29481,N_15742,N_13524);
nand U29482 (N_29482,N_16173,N_10420);
and U29483 (N_29483,N_13925,N_11975);
and U29484 (N_29484,N_15702,N_19229);
and U29485 (N_29485,N_11186,N_13270);
and U29486 (N_29486,N_13346,N_19418);
nand U29487 (N_29487,N_14302,N_13940);
nand U29488 (N_29488,N_13505,N_16940);
nand U29489 (N_29489,N_17120,N_14251);
and U29490 (N_29490,N_17049,N_11412);
or U29491 (N_29491,N_17345,N_19227);
or U29492 (N_29492,N_17075,N_11910);
xor U29493 (N_29493,N_16912,N_12634);
or U29494 (N_29494,N_19774,N_15942);
nor U29495 (N_29495,N_18637,N_11859);
or U29496 (N_29496,N_11133,N_12734);
and U29497 (N_29497,N_15226,N_17194);
and U29498 (N_29498,N_18899,N_12248);
or U29499 (N_29499,N_11652,N_14519);
or U29500 (N_29500,N_12772,N_13425);
nor U29501 (N_29501,N_12079,N_19464);
nand U29502 (N_29502,N_18223,N_16703);
xor U29503 (N_29503,N_10963,N_12741);
and U29504 (N_29504,N_16169,N_10847);
nor U29505 (N_29505,N_14534,N_10006);
nor U29506 (N_29506,N_12255,N_10382);
xnor U29507 (N_29507,N_15391,N_14742);
nand U29508 (N_29508,N_11774,N_19588);
xor U29509 (N_29509,N_10924,N_10732);
and U29510 (N_29510,N_12419,N_10148);
nand U29511 (N_29511,N_19968,N_14371);
nand U29512 (N_29512,N_15666,N_11422);
or U29513 (N_29513,N_14105,N_19959);
xnor U29514 (N_29514,N_16034,N_13586);
nor U29515 (N_29515,N_15851,N_17257);
and U29516 (N_29516,N_12078,N_14679);
nor U29517 (N_29517,N_19245,N_14680);
nor U29518 (N_29518,N_11831,N_12336);
or U29519 (N_29519,N_14079,N_16685);
and U29520 (N_29520,N_16776,N_12048);
or U29521 (N_29521,N_19973,N_15957);
nor U29522 (N_29522,N_13591,N_13157);
or U29523 (N_29523,N_18571,N_17380);
nor U29524 (N_29524,N_14432,N_17535);
xnor U29525 (N_29525,N_14470,N_18909);
xor U29526 (N_29526,N_13670,N_16786);
and U29527 (N_29527,N_11422,N_15865);
and U29528 (N_29528,N_11416,N_14776);
xor U29529 (N_29529,N_15275,N_15322);
nor U29530 (N_29530,N_19787,N_16458);
xnor U29531 (N_29531,N_10885,N_12675);
or U29532 (N_29532,N_10384,N_10719);
or U29533 (N_29533,N_11125,N_14740);
xnor U29534 (N_29534,N_13144,N_19943);
or U29535 (N_29535,N_19742,N_12680);
nand U29536 (N_29536,N_16399,N_18592);
nor U29537 (N_29537,N_15716,N_15563);
and U29538 (N_29538,N_14874,N_11391);
xnor U29539 (N_29539,N_11023,N_14969);
or U29540 (N_29540,N_10556,N_15980);
and U29541 (N_29541,N_18741,N_18274);
xnor U29542 (N_29542,N_16613,N_16587);
and U29543 (N_29543,N_10916,N_11003);
and U29544 (N_29544,N_16516,N_11486);
or U29545 (N_29545,N_14382,N_12338);
and U29546 (N_29546,N_13753,N_17516);
nor U29547 (N_29547,N_13545,N_17777);
nand U29548 (N_29548,N_19383,N_11503);
and U29549 (N_29549,N_12046,N_14827);
and U29550 (N_29550,N_13782,N_12637);
nand U29551 (N_29551,N_15606,N_16012);
nand U29552 (N_29552,N_14567,N_15438);
nand U29553 (N_29553,N_10700,N_13329);
xnor U29554 (N_29554,N_12054,N_14113);
xor U29555 (N_29555,N_17876,N_14891);
nor U29556 (N_29556,N_12081,N_12204);
xnor U29557 (N_29557,N_14371,N_15312);
nor U29558 (N_29558,N_16945,N_10044);
nor U29559 (N_29559,N_10666,N_17132);
nor U29560 (N_29560,N_19251,N_11927);
nor U29561 (N_29561,N_15955,N_12877);
and U29562 (N_29562,N_18432,N_11479);
xor U29563 (N_29563,N_17341,N_11206);
or U29564 (N_29564,N_15148,N_10762);
nor U29565 (N_29565,N_19645,N_12377);
xor U29566 (N_29566,N_18989,N_10376);
xor U29567 (N_29567,N_15317,N_19005);
nor U29568 (N_29568,N_11158,N_13515);
or U29569 (N_29569,N_18154,N_13758);
nor U29570 (N_29570,N_12836,N_18793);
or U29571 (N_29571,N_10275,N_12243);
nand U29572 (N_29572,N_15098,N_19873);
xor U29573 (N_29573,N_12204,N_11697);
xnor U29574 (N_29574,N_11240,N_18339);
xor U29575 (N_29575,N_13554,N_10805);
nand U29576 (N_29576,N_14458,N_13454);
and U29577 (N_29577,N_15930,N_12987);
xor U29578 (N_29578,N_18317,N_18855);
or U29579 (N_29579,N_14106,N_19125);
nand U29580 (N_29580,N_12966,N_18639);
nor U29581 (N_29581,N_19314,N_19919);
nor U29582 (N_29582,N_11185,N_17789);
nand U29583 (N_29583,N_13063,N_16243);
nor U29584 (N_29584,N_16729,N_19375);
xor U29585 (N_29585,N_18767,N_10895);
or U29586 (N_29586,N_15298,N_14963);
or U29587 (N_29587,N_14300,N_11694);
nor U29588 (N_29588,N_16735,N_17280);
and U29589 (N_29589,N_19866,N_15237);
nor U29590 (N_29590,N_18624,N_12442);
nor U29591 (N_29591,N_18336,N_18148);
and U29592 (N_29592,N_16255,N_10266);
and U29593 (N_29593,N_10129,N_17053);
or U29594 (N_29594,N_15289,N_12278);
or U29595 (N_29595,N_15222,N_14245);
nor U29596 (N_29596,N_13934,N_17196);
nor U29597 (N_29597,N_19146,N_13521);
xor U29598 (N_29598,N_12611,N_10779);
xnor U29599 (N_29599,N_11604,N_12196);
and U29600 (N_29600,N_12298,N_10874);
and U29601 (N_29601,N_19023,N_11466);
and U29602 (N_29602,N_16205,N_13543);
or U29603 (N_29603,N_15473,N_14087);
nand U29604 (N_29604,N_15937,N_15840);
nor U29605 (N_29605,N_19665,N_19570);
or U29606 (N_29606,N_13476,N_15790);
and U29607 (N_29607,N_17212,N_15348);
xnor U29608 (N_29608,N_14246,N_19140);
or U29609 (N_29609,N_18135,N_17997);
nor U29610 (N_29610,N_14241,N_17345);
nand U29611 (N_29611,N_19727,N_17977);
and U29612 (N_29612,N_18151,N_17650);
or U29613 (N_29613,N_15815,N_11699);
or U29614 (N_29614,N_13875,N_13998);
xor U29615 (N_29615,N_18565,N_11821);
nor U29616 (N_29616,N_12300,N_18737);
xnor U29617 (N_29617,N_14313,N_13038);
nor U29618 (N_29618,N_13338,N_11513);
xnor U29619 (N_29619,N_13493,N_11307);
and U29620 (N_29620,N_16719,N_19127);
xor U29621 (N_29621,N_13529,N_14486);
xor U29622 (N_29622,N_16348,N_17838);
and U29623 (N_29623,N_17695,N_11300);
nand U29624 (N_29624,N_15531,N_15408);
nand U29625 (N_29625,N_16508,N_11508);
and U29626 (N_29626,N_15905,N_10383);
nand U29627 (N_29627,N_15642,N_18329);
xor U29628 (N_29628,N_19698,N_16865);
or U29629 (N_29629,N_10732,N_14664);
nand U29630 (N_29630,N_16309,N_14221);
nand U29631 (N_29631,N_15487,N_11449);
nand U29632 (N_29632,N_14324,N_16769);
xor U29633 (N_29633,N_17661,N_15952);
nor U29634 (N_29634,N_15375,N_17753);
and U29635 (N_29635,N_15274,N_11251);
nand U29636 (N_29636,N_16733,N_13601);
or U29637 (N_29637,N_11514,N_15623);
xnor U29638 (N_29638,N_17762,N_13367);
nor U29639 (N_29639,N_17927,N_13751);
nor U29640 (N_29640,N_13004,N_17307);
nand U29641 (N_29641,N_10105,N_11733);
nand U29642 (N_29642,N_12753,N_17555);
xnor U29643 (N_29643,N_11648,N_16358);
nor U29644 (N_29644,N_15893,N_16848);
nor U29645 (N_29645,N_17194,N_16330);
nand U29646 (N_29646,N_17226,N_14514);
and U29647 (N_29647,N_14720,N_19902);
and U29648 (N_29648,N_10887,N_11037);
nor U29649 (N_29649,N_12734,N_16370);
and U29650 (N_29650,N_17275,N_11425);
xor U29651 (N_29651,N_13444,N_13195);
nand U29652 (N_29652,N_14601,N_10290);
xnor U29653 (N_29653,N_12959,N_10085);
nand U29654 (N_29654,N_10938,N_16436);
nand U29655 (N_29655,N_11796,N_18945);
nor U29656 (N_29656,N_17310,N_14803);
nor U29657 (N_29657,N_11029,N_13554);
nand U29658 (N_29658,N_18709,N_17635);
nor U29659 (N_29659,N_18401,N_17091);
and U29660 (N_29660,N_11134,N_18314);
nor U29661 (N_29661,N_13625,N_17167);
nor U29662 (N_29662,N_14313,N_16955);
xor U29663 (N_29663,N_14718,N_11621);
xnor U29664 (N_29664,N_17060,N_11735);
or U29665 (N_29665,N_16510,N_16875);
or U29666 (N_29666,N_11494,N_11227);
nor U29667 (N_29667,N_15275,N_15886);
nor U29668 (N_29668,N_14201,N_13064);
nand U29669 (N_29669,N_12515,N_16676);
xor U29670 (N_29670,N_13079,N_17698);
xor U29671 (N_29671,N_19549,N_13602);
xnor U29672 (N_29672,N_12635,N_16294);
nand U29673 (N_29673,N_19561,N_16031);
and U29674 (N_29674,N_17504,N_18152);
xnor U29675 (N_29675,N_14722,N_15358);
nand U29676 (N_29676,N_16185,N_16005);
and U29677 (N_29677,N_19941,N_14605);
and U29678 (N_29678,N_11392,N_17751);
or U29679 (N_29679,N_11693,N_15408);
or U29680 (N_29680,N_16078,N_19095);
xor U29681 (N_29681,N_17933,N_14599);
xor U29682 (N_29682,N_18167,N_11270);
or U29683 (N_29683,N_17130,N_12213);
nand U29684 (N_29684,N_11779,N_18395);
and U29685 (N_29685,N_18797,N_10923);
nand U29686 (N_29686,N_13192,N_17376);
xnor U29687 (N_29687,N_18782,N_16274);
or U29688 (N_29688,N_16679,N_10073);
nand U29689 (N_29689,N_14658,N_15494);
xor U29690 (N_29690,N_14036,N_18189);
nor U29691 (N_29691,N_14642,N_17356);
nor U29692 (N_29692,N_17907,N_14663);
or U29693 (N_29693,N_14281,N_11966);
nor U29694 (N_29694,N_18209,N_11243);
nand U29695 (N_29695,N_17317,N_10633);
or U29696 (N_29696,N_11748,N_12588);
nand U29697 (N_29697,N_10707,N_12474);
or U29698 (N_29698,N_19936,N_16047);
and U29699 (N_29699,N_15234,N_18511);
and U29700 (N_29700,N_16463,N_19985);
nand U29701 (N_29701,N_13285,N_17037);
and U29702 (N_29702,N_10259,N_12588);
nor U29703 (N_29703,N_17089,N_10819);
and U29704 (N_29704,N_11016,N_10303);
nor U29705 (N_29705,N_19810,N_17408);
nor U29706 (N_29706,N_13851,N_12206);
nand U29707 (N_29707,N_14552,N_13534);
or U29708 (N_29708,N_16781,N_15306);
nand U29709 (N_29709,N_11954,N_17104);
and U29710 (N_29710,N_13274,N_12129);
nand U29711 (N_29711,N_10029,N_16697);
xor U29712 (N_29712,N_14407,N_12040);
and U29713 (N_29713,N_11369,N_18543);
xor U29714 (N_29714,N_18914,N_14360);
and U29715 (N_29715,N_19263,N_17707);
xnor U29716 (N_29716,N_13687,N_18715);
nor U29717 (N_29717,N_13877,N_13250);
and U29718 (N_29718,N_19534,N_13077);
and U29719 (N_29719,N_15941,N_12314);
nand U29720 (N_29720,N_16296,N_10227);
nor U29721 (N_29721,N_19931,N_12190);
nor U29722 (N_29722,N_12350,N_18386);
xor U29723 (N_29723,N_10930,N_14667);
nand U29724 (N_29724,N_14865,N_18327);
nor U29725 (N_29725,N_18834,N_12898);
nand U29726 (N_29726,N_11984,N_17215);
or U29727 (N_29727,N_10917,N_11333);
or U29728 (N_29728,N_12143,N_12500);
or U29729 (N_29729,N_11572,N_19962);
and U29730 (N_29730,N_16791,N_17954);
or U29731 (N_29731,N_15646,N_19322);
nand U29732 (N_29732,N_18283,N_15705);
nor U29733 (N_29733,N_10427,N_18896);
or U29734 (N_29734,N_11694,N_12648);
and U29735 (N_29735,N_16548,N_10510);
and U29736 (N_29736,N_14310,N_18677);
or U29737 (N_29737,N_12609,N_12493);
and U29738 (N_29738,N_15458,N_10352);
or U29739 (N_29739,N_14205,N_14216);
xor U29740 (N_29740,N_12948,N_11352);
nor U29741 (N_29741,N_19167,N_12289);
and U29742 (N_29742,N_19205,N_13391);
and U29743 (N_29743,N_10895,N_12688);
and U29744 (N_29744,N_12445,N_19080);
xnor U29745 (N_29745,N_19312,N_17499);
xnor U29746 (N_29746,N_13637,N_10162);
xor U29747 (N_29747,N_13922,N_18470);
nor U29748 (N_29748,N_15984,N_14630);
or U29749 (N_29749,N_12216,N_12146);
xnor U29750 (N_29750,N_10911,N_18362);
nand U29751 (N_29751,N_14112,N_18281);
nand U29752 (N_29752,N_17231,N_15296);
xnor U29753 (N_29753,N_10361,N_12110);
and U29754 (N_29754,N_14849,N_12344);
nand U29755 (N_29755,N_14102,N_10760);
nand U29756 (N_29756,N_14560,N_15545);
and U29757 (N_29757,N_15364,N_11503);
nand U29758 (N_29758,N_12728,N_12499);
nand U29759 (N_29759,N_18003,N_12922);
or U29760 (N_29760,N_17715,N_15615);
xnor U29761 (N_29761,N_15530,N_17929);
nor U29762 (N_29762,N_19963,N_15308);
or U29763 (N_29763,N_17669,N_16847);
and U29764 (N_29764,N_14476,N_11382);
or U29765 (N_29765,N_19078,N_11407);
xor U29766 (N_29766,N_11288,N_16585);
or U29767 (N_29767,N_11429,N_16697);
and U29768 (N_29768,N_19018,N_19522);
nor U29769 (N_29769,N_15502,N_12860);
nand U29770 (N_29770,N_17832,N_12502);
and U29771 (N_29771,N_16078,N_17472);
nor U29772 (N_29772,N_17301,N_12175);
nand U29773 (N_29773,N_17028,N_10114);
xor U29774 (N_29774,N_19475,N_16087);
and U29775 (N_29775,N_16539,N_11679);
xnor U29776 (N_29776,N_17264,N_12124);
nand U29777 (N_29777,N_11604,N_12937);
xor U29778 (N_29778,N_14128,N_19182);
nor U29779 (N_29779,N_19250,N_10873);
xnor U29780 (N_29780,N_15807,N_17670);
xor U29781 (N_29781,N_12156,N_17781);
or U29782 (N_29782,N_12653,N_17146);
nand U29783 (N_29783,N_17733,N_17092);
nor U29784 (N_29784,N_19382,N_12374);
nor U29785 (N_29785,N_13907,N_17752);
nand U29786 (N_29786,N_18594,N_19169);
and U29787 (N_29787,N_16514,N_16106);
xnor U29788 (N_29788,N_18000,N_12811);
and U29789 (N_29789,N_16356,N_12440);
nor U29790 (N_29790,N_13667,N_12311);
and U29791 (N_29791,N_17362,N_16637);
xnor U29792 (N_29792,N_17514,N_15432);
or U29793 (N_29793,N_10266,N_18893);
or U29794 (N_29794,N_10768,N_17035);
xor U29795 (N_29795,N_12985,N_19670);
or U29796 (N_29796,N_10218,N_19542);
or U29797 (N_29797,N_18453,N_16216);
or U29798 (N_29798,N_12915,N_11638);
nor U29799 (N_29799,N_12009,N_14302);
nor U29800 (N_29800,N_11666,N_15956);
nand U29801 (N_29801,N_13276,N_10705);
nor U29802 (N_29802,N_18851,N_14187);
xnor U29803 (N_29803,N_13549,N_17756);
or U29804 (N_29804,N_11661,N_13656);
nand U29805 (N_29805,N_15128,N_14817);
nor U29806 (N_29806,N_19759,N_13728);
or U29807 (N_29807,N_10074,N_19753);
and U29808 (N_29808,N_12239,N_19778);
or U29809 (N_29809,N_16097,N_19710);
xnor U29810 (N_29810,N_12058,N_17382);
nor U29811 (N_29811,N_10373,N_14194);
or U29812 (N_29812,N_10174,N_11904);
and U29813 (N_29813,N_15821,N_18215);
and U29814 (N_29814,N_18456,N_13595);
or U29815 (N_29815,N_12726,N_15851);
xnor U29816 (N_29816,N_18331,N_11392);
xnor U29817 (N_29817,N_18323,N_19420);
or U29818 (N_29818,N_13558,N_14421);
or U29819 (N_29819,N_13451,N_11500);
or U29820 (N_29820,N_11208,N_13537);
xor U29821 (N_29821,N_19944,N_10033);
xnor U29822 (N_29822,N_11577,N_10902);
nand U29823 (N_29823,N_12129,N_18157);
and U29824 (N_29824,N_17902,N_13086);
and U29825 (N_29825,N_10446,N_11419);
nor U29826 (N_29826,N_11908,N_16290);
xor U29827 (N_29827,N_17481,N_12612);
nor U29828 (N_29828,N_10216,N_11830);
nor U29829 (N_29829,N_17581,N_17849);
xor U29830 (N_29830,N_16012,N_14627);
and U29831 (N_29831,N_13937,N_16446);
xnor U29832 (N_29832,N_18945,N_10700);
or U29833 (N_29833,N_19654,N_13805);
xnor U29834 (N_29834,N_11157,N_18223);
nand U29835 (N_29835,N_10062,N_12150);
nand U29836 (N_29836,N_12606,N_19174);
xor U29837 (N_29837,N_10128,N_13570);
or U29838 (N_29838,N_10715,N_16561);
or U29839 (N_29839,N_18326,N_16999);
xor U29840 (N_29840,N_12340,N_12344);
or U29841 (N_29841,N_11801,N_15937);
nor U29842 (N_29842,N_15292,N_15977);
or U29843 (N_29843,N_15639,N_17749);
or U29844 (N_29844,N_10878,N_16875);
or U29845 (N_29845,N_11529,N_19546);
nand U29846 (N_29846,N_15901,N_11021);
or U29847 (N_29847,N_18863,N_14421);
xnor U29848 (N_29848,N_15578,N_12671);
or U29849 (N_29849,N_10276,N_10385);
and U29850 (N_29850,N_17043,N_18115);
nor U29851 (N_29851,N_17408,N_16944);
nor U29852 (N_29852,N_12832,N_14298);
xnor U29853 (N_29853,N_19157,N_10271);
nand U29854 (N_29854,N_19331,N_15839);
and U29855 (N_29855,N_16004,N_17860);
nor U29856 (N_29856,N_11131,N_16301);
nor U29857 (N_29857,N_12081,N_10657);
nor U29858 (N_29858,N_15529,N_11467);
nand U29859 (N_29859,N_14562,N_14567);
xor U29860 (N_29860,N_19604,N_17448);
nor U29861 (N_29861,N_11601,N_10687);
xnor U29862 (N_29862,N_15226,N_19770);
or U29863 (N_29863,N_11109,N_18592);
nor U29864 (N_29864,N_13357,N_17339);
nand U29865 (N_29865,N_10244,N_11303);
nand U29866 (N_29866,N_18098,N_15401);
xor U29867 (N_29867,N_16418,N_16604);
or U29868 (N_29868,N_10399,N_16141);
nand U29869 (N_29869,N_18908,N_14971);
or U29870 (N_29870,N_18404,N_11363);
and U29871 (N_29871,N_13485,N_18947);
or U29872 (N_29872,N_15710,N_17340);
nand U29873 (N_29873,N_14374,N_12516);
nand U29874 (N_29874,N_11231,N_15223);
nor U29875 (N_29875,N_13915,N_17499);
nand U29876 (N_29876,N_19885,N_17165);
nor U29877 (N_29877,N_11256,N_18882);
nor U29878 (N_29878,N_19536,N_11047);
xor U29879 (N_29879,N_14056,N_11394);
nand U29880 (N_29880,N_13049,N_15012);
xnor U29881 (N_29881,N_17975,N_19728);
nor U29882 (N_29882,N_12286,N_17400);
nor U29883 (N_29883,N_18808,N_10794);
nand U29884 (N_29884,N_13008,N_19116);
nor U29885 (N_29885,N_18976,N_18633);
and U29886 (N_29886,N_11675,N_10095);
xnor U29887 (N_29887,N_10959,N_14866);
or U29888 (N_29888,N_12687,N_13785);
and U29889 (N_29889,N_19999,N_15246);
nor U29890 (N_29890,N_16187,N_15357);
nor U29891 (N_29891,N_16584,N_12713);
or U29892 (N_29892,N_19998,N_18783);
or U29893 (N_29893,N_13075,N_15437);
nand U29894 (N_29894,N_13474,N_17813);
nand U29895 (N_29895,N_14452,N_13529);
nor U29896 (N_29896,N_14585,N_18374);
xnor U29897 (N_29897,N_18682,N_19014);
nor U29898 (N_29898,N_14329,N_15722);
nor U29899 (N_29899,N_10118,N_17279);
xor U29900 (N_29900,N_17838,N_12576);
and U29901 (N_29901,N_19629,N_10765);
and U29902 (N_29902,N_14080,N_18493);
nand U29903 (N_29903,N_12909,N_13125);
xor U29904 (N_29904,N_19060,N_11260);
and U29905 (N_29905,N_16877,N_16415);
xnor U29906 (N_29906,N_19466,N_19067);
nand U29907 (N_29907,N_14001,N_18696);
or U29908 (N_29908,N_10781,N_10791);
nor U29909 (N_29909,N_11080,N_14936);
xnor U29910 (N_29910,N_14882,N_12658);
nor U29911 (N_29911,N_15951,N_17817);
or U29912 (N_29912,N_14591,N_13441);
and U29913 (N_29913,N_13366,N_14560);
and U29914 (N_29914,N_19822,N_19179);
or U29915 (N_29915,N_18601,N_18772);
or U29916 (N_29916,N_19104,N_17197);
nor U29917 (N_29917,N_11719,N_11912);
or U29918 (N_29918,N_10113,N_18323);
and U29919 (N_29919,N_16111,N_11851);
xnor U29920 (N_29920,N_15062,N_15617);
and U29921 (N_29921,N_13475,N_18501);
xnor U29922 (N_29922,N_14045,N_13162);
or U29923 (N_29923,N_10390,N_12871);
and U29924 (N_29924,N_11457,N_19864);
and U29925 (N_29925,N_15538,N_16896);
or U29926 (N_29926,N_10046,N_14207);
xor U29927 (N_29927,N_13800,N_10319);
or U29928 (N_29928,N_12561,N_18797);
or U29929 (N_29929,N_17521,N_10847);
xor U29930 (N_29930,N_10410,N_17842);
nand U29931 (N_29931,N_12480,N_16104);
nand U29932 (N_29932,N_18760,N_19774);
and U29933 (N_29933,N_17252,N_10613);
nor U29934 (N_29934,N_12798,N_11733);
or U29935 (N_29935,N_18544,N_14309);
or U29936 (N_29936,N_12412,N_14942);
nand U29937 (N_29937,N_11413,N_19602);
or U29938 (N_29938,N_18043,N_14632);
nand U29939 (N_29939,N_19681,N_19576);
or U29940 (N_29940,N_12373,N_19351);
nor U29941 (N_29941,N_12194,N_11842);
nand U29942 (N_29942,N_13202,N_15576);
and U29943 (N_29943,N_19647,N_15304);
nor U29944 (N_29944,N_12038,N_19358);
or U29945 (N_29945,N_18399,N_11334);
and U29946 (N_29946,N_18979,N_12382);
nor U29947 (N_29947,N_18300,N_18686);
nand U29948 (N_29948,N_13394,N_14275);
and U29949 (N_29949,N_12450,N_15292);
and U29950 (N_29950,N_10737,N_11581);
or U29951 (N_29951,N_15371,N_16789);
xnor U29952 (N_29952,N_14085,N_17899);
and U29953 (N_29953,N_15842,N_16616);
and U29954 (N_29954,N_11178,N_14559);
or U29955 (N_29955,N_16230,N_14491);
and U29956 (N_29956,N_17071,N_10315);
and U29957 (N_29957,N_13121,N_15569);
nor U29958 (N_29958,N_12644,N_19303);
nor U29959 (N_29959,N_18003,N_19094);
nand U29960 (N_29960,N_11562,N_10874);
nor U29961 (N_29961,N_19737,N_15978);
and U29962 (N_29962,N_11360,N_10292);
nor U29963 (N_29963,N_17181,N_16142);
and U29964 (N_29964,N_14955,N_18381);
or U29965 (N_29965,N_14415,N_18866);
nor U29966 (N_29966,N_17028,N_19015);
nor U29967 (N_29967,N_14633,N_12410);
nor U29968 (N_29968,N_11613,N_11063);
nand U29969 (N_29969,N_16367,N_16784);
or U29970 (N_29970,N_16283,N_17976);
nand U29971 (N_29971,N_15365,N_15661);
nand U29972 (N_29972,N_19162,N_11455);
and U29973 (N_29973,N_16489,N_10660);
nand U29974 (N_29974,N_11549,N_10498);
nor U29975 (N_29975,N_13380,N_13106);
or U29976 (N_29976,N_17242,N_16064);
nand U29977 (N_29977,N_14738,N_13233);
and U29978 (N_29978,N_17654,N_12400);
or U29979 (N_29979,N_10115,N_15292);
xor U29980 (N_29980,N_14923,N_16384);
xor U29981 (N_29981,N_17568,N_13069);
xor U29982 (N_29982,N_16451,N_10841);
or U29983 (N_29983,N_11399,N_15772);
xor U29984 (N_29984,N_10917,N_13329);
nand U29985 (N_29985,N_14217,N_19384);
nand U29986 (N_29986,N_14618,N_14985);
or U29987 (N_29987,N_12071,N_12567);
or U29988 (N_29988,N_18392,N_13775);
nand U29989 (N_29989,N_12729,N_16879);
nor U29990 (N_29990,N_13936,N_18211);
nor U29991 (N_29991,N_19344,N_11524);
nand U29992 (N_29992,N_16648,N_18023);
xnor U29993 (N_29993,N_17583,N_12341);
nor U29994 (N_29994,N_11117,N_12434);
and U29995 (N_29995,N_12337,N_16766);
xnor U29996 (N_29996,N_18760,N_13330);
or U29997 (N_29997,N_17607,N_11283);
or U29998 (N_29998,N_16146,N_11928);
nor U29999 (N_29999,N_13951,N_16770);
and U30000 (N_30000,N_20325,N_26132);
xnor U30001 (N_30001,N_21000,N_29168);
or U30002 (N_30002,N_25438,N_27079);
xnor U30003 (N_30003,N_23249,N_25659);
nand U30004 (N_30004,N_27131,N_23709);
xnor U30005 (N_30005,N_29956,N_24786);
nand U30006 (N_30006,N_27528,N_26640);
xnor U30007 (N_30007,N_28693,N_20068);
and U30008 (N_30008,N_25016,N_28463);
nand U30009 (N_30009,N_21134,N_24302);
xor U30010 (N_30010,N_28496,N_27115);
nor U30011 (N_30011,N_22763,N_26272);
nand U30012 (N_30012,N_25324,N_20035);
xnor U30013 (N_30013,N_29548,N_23055);
xnor U30014 (N_30014,N_21467,N_23441);
and U30015 (N_30015,N_25884,N_25109);
nand U30016 (N_30016,N_25425,N_21223);
nand U30017 (N_30017,N_27826,N_29719);
xnor U30018 (N_30018,N_29231,N_21849);
and U30019 (N_30019,N_29922,N_20894);
or U30020 (N_30020,N_21718,N_27363);
nor U30021 (N_30021,N_23303,N_21272);
and U30022 (N_30022,N_29770,N_24863);
and U30023 (N_30023,N_20016,N_27739);
and U30024 (N_30024,N_27856,N_25603);
and U30025 (N_30025,N_21571,N_22001);
nor U30026 (N_30026,N_27706,N_28561);
nor U30027 (N_30027,N_25913,N_27198);
or U30028 (N_30028,N_24548,N_29673);
xnor U30029 (N_30029,N_27109,N_21631);
or U30030 (N_30030,N_24536,N_25865);
or U30031 (N_30031,N_24840,N_22016);
and U30032 (N_30032,N_21900,N_26635);
or U30033 (N_30033,N_25175,N_27558);
and U30034 (N_30034,N_21182,N_21511);
xor U30035 (N_30035,N_28247,N_25390);
xor U30036 (N_30036,N_29759,N_23101);
and U30037 (N_30037,N_27974,N_29711);
xnor U30038 (N_30038,N_21181,N_28907);
or U30039 (N_30039,N_23814,N_21575);
and U30040 (N_30040,N_21988,N_25836);
and U30041 (N_30041,N_27124,N_29612);
nand U30042 (N_30042,N_26375,N_20339);
nor U30043 (N_30043,N_20455,N_23765);
xnor U30044 (N_30044,N_23328,N_28807);
or U30045 (N_30045,N_25440,N_20095);
nand U30046 (N_30046,N_21288,N_28574);
xnor U30047 (N_30047,N_28539,N_24526);
nand U30048 (N_30048,N_28350,N_21757);
or U30049 (N_30049,N_21381,N_27361);
nand U30050 (N_30050,N_24031,N_22384);
or U30051 (N_30051,N_27684,N_21123);
or U30052 (N_30052,N_25667,N_22441);
or U30053 (N_30053,N_20492,N_26795);
nor U30054 (N_30054,N_29876,N_20049);
xnor U30055 (N_30055,N_27880,N_28512);
nor U30056 (N_30056,N_29116,N_29000);
nor U30057 (N_30057,N_26893,N_20482);
and U30058 (N_30058,N_25012,N_25442);
nor U30059 (N_30059,N_26602,N_21504);
or U30060 (N_30060,N_27405,N_26203);
or U30061 (N_30061,N_22470,N_29024);
and U30062 (N_30062,N_21090,N_28251);
or U30063 (N_30063,N_29640,N_29855);
nor U30064 (N_30064,N_27063,N_22131);
or U30065 (N_30065,N_23953,N_24218);
and U30066 (N_30066,N_23531,N_20113);
nand U30067 (N_30067,N_24650,N_21772);
or U30068 (N_30068,N_26976,N_26346);
xnor U30069 (N_30069,N_26028,N_27537);
nand U30070 (N_30070,N_23439,N_25188);
xor U30071 (N_30071,N_23198,N_21336);
xor U30072 (N_30072,N_26589,N_21366);
nor U30073 (N_30073,N_26331,N_22654);
nand U30074 (N_30074,N_25228,N_21137);
nor U30075 (N_30075,N_28006,N_24534);
or U30076 (N_30076,N_27332,N_27799);
nor U30077 (N_30077,N_21488,N_28376);
or U30078 (N_30078,N_20926,N_27947);
or U30079 (N_30079,N_29887,N_27687);
nor U30080 (N_30080,N_21946,N_24472);
nand U30081 (N_30081,N_28983,N_29473);
xor U30082 (N_30082,N_22159,N_25156);
nand U30083 (N_30083,N_29300,N_25378);
and U30084 (N_30084,N_24149,N_21099);
xor U30085 (N_30085,N_24423,N_29947);
and U30086 (N_30086,N_27302,N_24221);
or U30087 (N_30087,N_27979,N_22209);
or U30088 (N_30088,N_28716,N_26461);
or U30089 (N_30089,N_25819,N_20144);
and U30090 (N_30090,N_29725,N_25220);
or U30091 (N_30091,N_25297,N_21565);
and U30092 (N_30092,N_23586,N_21717);
nand U30093 (N_30093,N_29696,N_23174);
and U30094 (N_30094,N_25990,N_20983);
or U30095 (N_30095,N_21537,N_23888);
xor U30096 (N_30096,N_24699,N_22436);
nor U30097 (N_30097,N_23701,N_24879);
xnor U30098 (N_30098,N_28123,N_28974);
or U30099 (N_30099,N_20361,N_28062);
xor U30100 (N_30100,N_29668,N_24499);
nor U30101 (N_30101,N_28962,N_20648);
nand U30102 (N_30102,N_22888,N_21379);
xor U30103 (N_30103,N_21727,N_20042);
xor U30104 (N_30104,N_26089,N_21522);
nand U30105 (N_30105,N_28276,N_24080);
nor U30106 (N_30106,N_27464,N_22116);
nor U30107 (N_30107,N_27403,N_23553);
nand U30108 (N_30108,N_24481,N_23666);
nor U30109 (N_30109,N_26031,N_28960);
and U30110 (N_30110,N_29523,N_28842);
and U30111 (N_30111,N_23039,N_28707);
or U30112 (N_30112,N_27362,N_24244);
and U30113 (N_30113,N_29124,N_24238);
xnor U30114 (N_30114,N_28015,N_24184);
xor U30115 (N_30115,N_29364,N_25089);
or U30116 (N_30116,N_21682,N_22293);
and U30117 (N_30117,N_29138,N_25627);
or U30118 (N_30118,N_26469,N_29512);
or U30119 (N_30119,N_22633,N_25365);
nand U30120 (N_30120,N_22919,N_20893);
nand U30121 (N_30121,N_26159,N_25907);
or U30122 (N_30122,N_24187,N_26384);
xnor U30123 (N_30123,N_20053,N_20000);
and U30124 (N_30124,N_21232,N_25769);
xnor U30125 (N_30125,N_20093,N_25980);
or U30126 (N_30126,N_28585,N_20071);
nand U30127 (N_30127,N_24966,N_27892);
and U30128 (N_30128,N_27509,N_22081);
or U30129 (N_30129,N_22271,N_20913);
or U30130 (N_30130,N_23092,N_28820);
or U30131 (N_30131,N_24801,N_24920);
xor U30132 (N_30132,N_27450,N_25831);
or U30133 (N_30133,N_29718,N_26418);
nand U30134 (N_30134,N_22903,N_28022);
xor U30135 (N_30135,N_28466,N_29964);
xor U30136 (N_30136,N_20850,N_21354);
nand U30137 (N_30137,N_22482,N_20369);
nor U30138 (N_30138,N_27905,N_20137);
xnor U30139 (N_30139,N_26593,N_27018);
nor U30140 (N_30140,N_23018,N_23869);
xnor U30141 (N_30141,N_21022,N_29918);
xnor U30142 (N_30142,N_28887,N_21027);
nor U30143 (N_30143,N_21435,N_27713);
and U30144 (N_30144,N_27126,N_20588);
nand U30145 (N_30145,N_29829,N_21876);
nor U30146 (N_30146,N_26652,N_29498);
nor U30147 (N_30147,N_20796,N_27328);
nor U30148 (N_30148,N_20950,N_22376);
nor U30149 (N_30149,N_24556,N_21461);
and U30150 (N_30150,N_22180,N_23202);
nor U30151 (N_30151,N_23449,N_21630);
or U30152 (N_30152,N_20067,N_23589);
nor U30153 (N_30153,N_29821,N_28448);
nor U30154 (N_30154,N_26393,N_23115);
nand U30155 (N_30155,N_23343,N_26883);
or U30156 (N_30156,N_27549,N_29741);
nor U30157 (N_30157,N_24940,N_27698);
xor U30158 (N_30158,N_21172,N_23399);
xnor U30159 (N_30159,N_28738,N_27099);
or U30160 (N_30160,N_25209,N_22440);
nand U30161 (N_30161,N_21785,N_27801);
or U30162 (N_30162,N_27266,N_23472);
nor U30163 (N_30163,N_27635,N_22770);
or U30164 (N_30164,N_27555,N_24643);
or U30165 (N_30165,N_25063,N_29485);
nor U30166 (N_30166,N_20277,N_24630);
and U30167 (N_30167,N_20064,N_23958);
and U30168 (N_30168,N_26670,N_20965);
nor U30169 (N_30169,N_21980,N_25981);
nor U30170 (N_30170,N_28285,N_22748);
nor U30171 (N_30171,N_24850,N_20753);
nor U30172 (N_30172,N_23098,N_20839);
nand U30173 (N_30173,N_28952,N_22089);
nand U30174 (N_30174,N_21294,N_26386);
nor U30175 (N_30175,N_25079,N_21708);
nand U30176 (N_30176,N_27616,N_24435);
or U30177 (N_30177,N_20907,N_28538);
or U30178 (N_30178,N_25041,N_25577);
nand U30179 (N_30179,N_26389,N_23175);
nor U30180 (N_30180,N_23990,N_21916);
nand U30181 (N_30181,N_28883,N_26765);
xor U30182 (N_30182,N_23703,N_21407);
nor U30183 (N_30183,N_27092,N_28316);
or U30184 (N_30184,N_22285,N_28313);
and U30185 (N_30185,N_29915,N_26179);
nor U30186 (N_30186,N_22539,N_25481);
xor U30187 (N_30187,N_26769,N_21784);
nor U30188 (N_30188,N_25232,N_24621);
xor U30189 (N_30189,N_25714,N_29306);
nand U30190 (N_30190,N_21450,N_27718);
or U30191 (N_30191,N_23535,N_24724);
and U30192 (N_30192,N_21868,N_27936);
and U30193 (N_30193,N_21841,N_26597);
nand U30194 (N_30194,N_25578,N_20643);
and U30195 (N_30195,N_21879,N_22336);
nand U30196 (N_30196,N_25931,N_29826);
xnor U30197 (N_30197,N_25689,N_28554);
nor U30198 (N_30198,N_22216,N_25951);
and U30199 (N_30199,N_22583,N_21041);
or U30200 (N_30200,N_27357,N_29465);
xor U30201 (N_30201,N_25541,N_20097);
and U30202 (N_30202,N_22920,N_25364);
and U30203 (N_30203,N_24718,N_28624);
nor U30204 (N_30204,N_28798,N_20689);
xor U30205 (N_30205,N_28275,N_27026);
and U30206 (N_30206,N_26921,N_29686);
nand U30207 (N_30207,N_28205,N_27762);
nand U30208 (N_30208,N_26142,N_22864);
or U30209 (N_30209,N_28548,N_21852);
nor U30210 (N_30210,N_24053,N_22789);
nor U30211 (N_30211,N_28060,N_28174);
nand U30212 (N_30212,N_24427,N_24150);
nor U30213 (N_30213,N_23520,N_24041);
and U30214 (N_30214,N_23534,N_22022);
nand U30215 (N_30215,N_24119,N_26822);
xnor U30216 (N_30216,N_28299,N_28633);
or U30217 (N_30217,N_26284,N_29987);
nand U30218 (N_30218,N_25007,N_26804);
xor U30219 (N_30219,N_24524,N_29784);
and U30220 (N_30220,N_29564,N_27052);
and U30221 (N_30221,N_24952,N_28287);
xor U30222 (N_30222,N_22853,N_26918);
nor U30223 (N_30223,N_23504,N_27525);
or U30224 (N_30224,N_25483,N_22126);
nand U30225 (N_30225,N_24628,N_20609);
or U30226 (N_30226,N_27247,N_24349);
nand U30227 (N_30227,N_22784,N_20251);
xor U30228 (N_30228,N_27506,N_26091);
or U30229 (N_30229,N_20876,N_24716);
nand U30230 (N_30230,N_26083,N_27765);
xor U30231 (N_30231,N_22195,N_20014);
or U30232 (N_30232,N_24931,N_26261);
xor U30233 (N_30233,N_22706,N_26685);
or U30234 (N_30234,N_20048,N_29480);
nand U30235 (N_30235,N_29596,N_24077);
xnor U30236 (N_30236,N_25219,N_24996);
and U30237 (N_30237,N_27303,N_20915);
and U30238 (N_30238,N_26025,N_28722);
and U30239 (N_30239,N_20452,N_21131);
xor U30240 (N_30240,N_27061,N_22123);
or U30241 (N_30241,N_29228,N_24819);
nor U30242 (N_30242,N_22523,N_28164);
and U30243 (N_30243,N_26547,N_20192);
and U30244 (N_30244,N_28226,N_23354);
or U30245 (N_30245,N_21857,N_22495);
or U30246 (N_30246,N_28347,N_27173);
and U30247 (N_30247,N_29284,N_28419);
or U30248 (N_30248,N_21471,N_20574);
xnor U30249 (N_30249,N_29370,N_21551);
nor U30250 (N_30250,N_20226,N_29200);
xor U30251 (N_30251,N_20139,N_28603);
xor U30252 (N_30252,N_25361,N_22786);
nand U30253 (N_30253,N_20208,N_20867);
xor U30254 (N_30254,N_27355,N_23281);
nor U30255 (N_30255,N_21109,N_24384);
and U30256 (N_30256,N_21590,N_21117);
or U30257 (N_30257,N_25302,N_20128);
or U30258 (N_30258,N_22316,N_23356);
nor U30259 (N_30259,N_27662,N_25904);
and U30260 (N_30260,N_20816,N_23781);
or U30261 (N_30261,N_23274,N_25550);
and U30262 (N_30262,N_22282,N_22509);
nand U30263 (N_30263,N_22727,N_28249);
nand U30264 (N_30264,N_21224,N_21752);
xor U30265 (N_30265,N_28033,N_23542);
xnor U30266 (N_30266,N_20754,N_28104);
nand U30267 (N_30267,N_24660,N_26931);
and U30268 (N_30268,N_25976,N_28348);
or U30269 (N_30269,N_23764,N_29699);
nand U30270 (N_30270,N_22532,N_22624);
or U30271 (N_30271,N_26361,N_23643);
and U30272 (N_30272,N_25526,N_23886);
nor U30273 (N_30273,N_21855,N_24419);
or U30274 (N_30274,N_25818,N_25244);
and U30275 (N_30275,N_23350,N_21078);
or U30276 (N_30276,N_24251,N_23443);
xnor U30277 (N_30277,N_22047,N_21888);
and U30278 (N_30278,N_20763,N_20107);
nand U30279 (N_30279,N_26338,N_27960);
nand U30280 (N_30280,N_27280,N_26618);
nor U30281 (N_30281,N_20903,N_23731);
nor U30282 (N_30282,N_23577,N_21886);
nor U30283 (N_30283,N_23426,N_24646);
and U30284 (N_30284,N_22833,N_23430);
or U30285 (N_30285,N_25991,N_26371);
or U30286 (N_30286,N_24904,N_23172);
xor U30287 (N_30287,N_20929,N_23784);
xnor U30288 (N_30288,N_27149,N_20830);
or U30289 (N_30289,N_27320,N_25509);
or U30290 (N_30290,N_23218,N_22467);
and U30291 (N_30291,N_26900,N_27078);
xnor U30292 (N_30292,N_26406,N_24290);
nand U30293 (N_30293,N_23629,N_21072);
nand U30294 (N_30294,N_25174,N_22063);
nor U30295 (N_30295,N_21419,N_28381);
and U30296 (N_30296,N_25166,N_22054);
or U30297 (N_30297,N_22430,N_24138);
and U30298 (N_30298,N_20709,N_21115);
and U30299 (N_30299,N_28206,N_24297);
nand U30300 (N_30300,N_23960,N_25103);
nor U30301 (N_30301,N_24124,N_21060);
or U30302 (N_30302,N_26303,N_27597);
and U30303 (N_30303,N_28999,N_21164);
xor U30304 (N_30304,N_20382,N_25136);
or U30305 (N_30305,N_22752,N_25668);
nand U30306 (N_30306,N_21581,N_20822);
nand U30307 (N_30307,N_29410,N_22405);
and U30308 (N_30308,N_26770,N_27903);
nand U30309 (N_30309,N_29463,N_20090);
nand U30310 (N_30310,N_26981,N_28110);
or U30311 (N_30311,N_26614,N_26874);
xor U30312 (N_30312,N_26004,N_22454);
and U30313 (N_30313,N_29760,N_21543);
xnor U30314 (N_30314,N_21698,N_28391);
xor U30315 (N_30315,N_25746,N_22881);
nor U30316 (N_30316,N_28578,N_20309);
nor U30317 (N_30317,N_20567,N_20991);
nand U30318 (N_30318,N_26725,N_26225);
and U30319 (N_30319,N_28521,N_28866);
and U30320 (N_30320,N_29620,N_22252);
or U30321 (N_30321,N_22905,N_21321);
or U30322 (N_30322,N_27530,N_24042);
nand U30323 (N_30323,N_26527,N_27704);
nor U30324 (N_30324,N_29560,N_23276);
and U30325 (N_30325,N_20881,N_26392);
nand U30326 (N_30326,N_21663,N_22820);
nand U30327 (N_30327,N_23912,N_20065);
or U30328 (N_30328,N_20184,N_27412);
nor U30329 (N_30329,N_28151,N_20552);
or U30330 (N_30330,N_25602,N_28748);
or U30331 (N_30331,N_26724,N_25795);
nand U30332 (N_30332,N_28238,N_28394);
xnor U30333 (N_30333,N_26431,N_22254);
nor U30334 (N_30334,N_29873,N_25524);
nor U30335 (N_30335,N_21148,N_29661);
or U30336 (N_30336,N_25712,N_22807);
or U30337 (N_30337,N_28584,N_29728);
and U30338 (N_30338,N_23187,N_20296);
or U30339 (N_30339,N_21409,N_24778);
and U30340 (N_30340,N_23183,N_20591);
and U30341 (N_30341,N_29360,N_24064);
nand U30342 (N_30342,N_25310,N_25817);
xor U30343 (N_30343,N_29288,N_21051);
nor U30344 (N_30344,N_26485,N_28344);
and U30345 (N_30345,N_25374,N_24166);
and U30346 (N_30346,N_25465,N_21157);
xor U30347 (N_30347,N_23468,N_21094);
and U30348 (N_30348,N_20166,N_20077);
and U30349 (N_30349,N_29587,N_23301);
nor U30350 (N_30350,N_21125,N_24429);
xnor U30351 (N_30351,N_23816,N_20928);
or U30352 (N_30352,N_21844,N_29891);
or U30353 (N_30353,N_25187,N_22240);
nor U30354 (N_30354,N_22055,N_22971);
nand U30355 (N_30355,N_26062,N_24637);
nor U30356 (N_30356,N_21647,N_27688);
or U30357 (N_30357,N_26932,N_21486);
nand U30358 (N_30358,N_29132,N_26733);
nand U30359 (N_30359,N_29082,N_21263);
nand U30360 (N_30360,N_26903,N_26189);
or U30361 (N_30361,N_24274,N_21616);
xnor U30362 (N_30362,N_24210,N_26949);
and U30363 (N_30363,N_25389,N_20174);
xnor U30364 (N_30364,N_20921,N_29779);
and U30365 (N_30365,N_24136,N_27264);
xor U30366 (N_30366,N_28638,N_23829);
xnor U30367 (N_30367,N_24783,N_21587);
and U30368 (N_30368,N_20631,N_27615);
or U30369 (N_30369,N_23223,N_22700);
and U30370 (N_30370,N_29246,N_21311);
and U30371 (N_30371,N_20414,N_25299);
xnor U30372 (N_30372,N_21282,N_29837);
xor U30373 (N_30373,N_23236,N_28925);
nand U30374 (N_30374,N_27674,N_20545);
or U30375 (N_30375,N_26862,N_26754);
nand U30376 (N_30376,N_22944,N_23125);
or U30377 (N_30377,N_27250,N_22113);
and U30378 (N_30378,N_27339,N_25521);
xnor U30379 (N_30379,N_22065,N_28417);
xor U30380 (N_30380,N_24692,N_23418);
and U30381 (N_30381,N_21293,N_21092);
nand U30382 (N_30382,N_23461,N_29795);
nand U30383 (N_30383,N_24457,N_22018);
xnor U30384 (N_30384,N_21364,N_29048);
or U30385 (N_30385,N_28525,N_24750);
or U30386 (N_30386,N_25009,N_22353);
or U30387 (N_30387,N_25347,N_24568);
nor U30388 (N_30388,N_28517,N_23311);
or U30389 (N_30389,N_20509,N_20898);
or U30390 (N_30390,N_24527,N_28118);
nand U30391 (N_30391,N_29967,N_26638);
nand U30392 (N_30392,N_26501,N_21524);
or U30393 (N_30393,N_26505,N_22787);
nor U30394 (N_30394,N_26776,N_21799);
and U30395 (N_30395,N_24252,N_25152);
and U30396 (N_30396,N_26078,N_22869);
nand U30397 (N_30397,N_25281,N_29994);
and U30398 (N_30398,N_25507,N_20219);
nor U30399 (N_30399,N_20598,N_27554);
nor U30400 (N_30400,N_27402,N_24372);
xor U30401 (N_30401,N_29287,N_21623);
and U30402 (N_30402,N_20498,N_29044);
and U30403 (N_30403,N_29221,N_26723);
or U30404 (N_30404,N_22476,N_29454);
or U30405 (N_30405,N_25148,N_27489);
nand U30406 (N_30406,N_27374,N_26763);
nor U30407 (N_30407,N_27116,N_26118);
or U30408 (N_30408,N_27730,N_20338);
or U30409 (N_30409,N_21594,N_28810);
nand U30410 (N_30410,N_22302,N_28209);
and U30411 (N_30411,N_22519,N_22671);
and U30412 (N_30412,N_27437,N_26106);
nor U30413 (N_30413,N_25333,N_27467);
and U30414 (N_30414,N_28830,N_27881);
nor U30415 (N_30415,N_20027,N_24224);
and U30416 (N_30416,N_21891,N_23800);
or U30417 (N_30417,N_29269,N_27950);
nand U30418 (N_30418,N_29274,N_28957);
xnor U30419 (N_30419,N_25475,N_23481);
nand U30420 (N_30420,N_29089,N_22810);
xnor U30421 (N_30421,N_22582,N_22184);
xor U30422 (N_30422,N_27317,N_25637);
xnor U30423 (N_30423,N_25595,N_24896);
nor U30424 (N_30424,N_23596,N_22259);
nand U30425 (N_30425,N_22576,N_24307);
nor U30426 (N_30426,N_23554,N_27686);
and U30427 (N_30427,N_20601,N_20801);
nor U30428 (N_30428,N_29373,N_26139);
nor U30429 (N_30429,N_23931,N_25682);
xnor U30430 (N_30430,N_20283,N_27417);
nor U30431 (N_30431,N_25031,N_29464);
or U30432 (N_30432,N_20860,N_23321);
or U30433 (N_30433,N_26668,N_29800);
nand U30434 (N_30434,N_29659,N_28679);
and U30435 (N_30435,N_21006,N_24444);
and U30436 (N_30436,N_26695,N_25290);
or U30437 (N_30437,N_24174,N_21417);
nand U30438 (N_30438,N_25258,N_29794);
nor U30439 (N_30439,N_28520,N_28655);
nor U30440 (N_30440,N_22988,N_24116);
nand U30441 (N_30441,N_23826,N_24507);
xnor U30442 (N_30442,N_22912,N_20103);
or U30443 (N_30443,N_21736,N_23459);
and U30444 (N_30444,N_28637,N_22725);
and U30445 (N_30445,N_20365,N_29580);
nand U30446 (N_30446,N_28429,N_22957);
nand U30447 (N_30447,N_25693,N_23661);
and U30448 (N_30448,N_29933,N_20556);
or U30449 (N_30449,N_20059,N_25340);
or U30450 (N_30450,N_27038,N_29256);
xor U30451 (N_30451,N_20052,N_27538);
and U30452 (N_30452,N_21593,N_25699);
nand U30453 (N_30453,N_27927,N_20542);
nand U30454 (N_30454,N_29926,N_26989);
nor U30455 (N_30455,N_28852,N_25939);
nor U30456 (N_30456,N_25767,N_22325);
nor U30457 (N_30457,N_24955,N_28059);
and U30458 (N_30458,N_21053,N_20232);
and U30459 (N_30459,N_26544,N_22696);
xnor U30460 (N_30460,N_21156,N_20846);
or U30461 (N_30461,N_21987,N_27352);
nand U30462 (N_30462,N_27691,N_23798);
nor U30463 (N_30463,N_23308,N_25610);
xor U30464 (N_30464,N_29601,N_21746);
xnor U30465 (N_30465,N_28864,N_26063);
xnor U30466 (N_30466,N_21510,N_20249);
xor U30467 (N_30467,N_22946,N_24823);
nand U30468 (N_30468,N_25083,N_24102);
and U30469 (N_30469,N_29626,N_29538);
or U30470 (N_30470,N_29258,N_28234);
or U30471 (N_30471,N_27922,N_26871);
or U30472 (N_30472,N_28310,N_29479);
nor U30473 (N_30473,N_25072,N_20444);
and U30474 (N_30474,N_23806,N_22067);
nor U30475 (N_30475,N_29263,N_28576);
or U30476 (N_30476,N_26200,N_28320);
nor U30477 (N_30477,N_28047,N_28608);
nor U30478 (N_30478,N_22061,N_22819);
nand U30479 (N_30479,N_27685,N_20378);
nand U30480 (N_30480,N_22965,N_23945);
xnor U30481 (N_30481,N_20145,N_21056);
xnor U30482 (N_30482,N_24129,N_24434);
nor U30483 (N_30483,N_25912,N_20920);
xnor U30484 (N_30484,N_21383,N_22442);
nor U30485 (N_30485,N_29244,N_25665);
nand U30486 (N_30486,N_27385,N_25396);
xnor U30487 (N_30487,N_23873,N_23635);
and U30488 (N_30488,N_28498,N_23246);
and U30489 (N_30489,N_25503,N_22361);
nand U30490 (N_30490,N_20678,N_20441);
nand U30491 (N_30491,N_29721,N_21477);
xor U30492 (N_30492,N_27513,N_27454);
nand U30493 (N_30493,N_26321,N_25633);
or U30494 (N_30494,N_26065,N_22518);
nand U30495 (N_30495,N_26454,N_26726);
and U30496 (N_30496,N_25048,N_22533);
or U30497 (N_30497,N_22120,N_22117);
xnor U30498 (N_30498,N_22359,N_25202);
and U30499 (N_30499,N_28465,N_22373);
nand U30500 (N_30500,N_20539,N_28240);
nor U30501 (N_30501,N_29945,N_20904);
and U30502 (N_30502,N_28121,N_22964);
or U30503 (N_30503,N_29303,N_21496);
and U30504 (N_30504,N_25873,N_26571);
xnor U30505 (N_30505,N_23695,N_27533);
nor U30506 (N_30506,N_29092,N_28076);
nor U30507 (N_30507,N_25807,N_29356);
nand U30508 (N_30508,N_28430,N_24059);
or U30509 (N_30509,N_26683,N_29056);
and U30510 (N_30510,N_21914,N_23982);
nor U30511 (N_30511,N_24014,N_29554);
or U30512 (N_30512,N_29091,N_21542);
nand U30513 (N_30513,N_25845,N_24214);
nor U30514 (N_30514,N_25329,N_26201);
and U30515 (N_30515,N_20167,N_26370);
nor U30516 (N_30516,N_28428,N_27980);
nand U30517 (N_30517,N_29158,N_20535);
nor U30518 (N_30518,N_26248,N_28618);
or U30519 (N_30519,N_25565,N_28241);
xnor U30520 (N_30520,N_26433,N_28278);
and U30521 (N_30521,N_23427,N_24596);
and U30522 (N_30522,N_21097,N_27368);
or U30523 (N_30523,N_27194,N_27961);
or U30524 (N_30524,N_22664,N_27353);
xor U30525 (N_30525,N_27824,N_20963);
or U30526 (N_30526,N_22591,N_27295);
or U30527 (N_30527,N_21351,N_28274);
xnor U30528 (N_30528,N_21777,N_24097);
or U30529 (N_30529,N_25843,N_25522);
nor U30530 (N_30530,N_25914,N_23412);
xor U30531 (N_30531,N_27014,N_21028);
nand U30532 (N_30532,N_24799,N_24144);
or U30533 (N_30533,N_23483,N_21699);
nand U30534 (N_30534,N_29417,N_25806);
xnor U30535 (N_30535,N_25275,N_27644);
and U30536 (N_30536,N_28850,N_25599);
nand U30537 (N_30537,N_21003,N_24828);
or U30538 (N_30538,N_27934,N_21729);
nand U30539 (N_30539,N_22627,N_22560);
nand U30540 (N_30540,N_24231,N_27226);
nor U30541 (N_30541,N_20304,N_22074);
xnor U30542 (N_30542,N_28345,N_29327);
or U30543 (N_30543,N_27143,N_25584);
or U30544 (N_30544,N_20112,N_29610);
or U30545 (N_30545,N_29907,N_25349);
xnor U30546 (N_30546,N_22354,N_29405);
and U30547 (N_30547,N_23995,N_23122);
nand U30548 (N_30548,N_27410,N_28991);
xor U30549 (N_30549,N_24094,N_24869);
xnor U30550 (N_30550,N_23621,N_20925);
and U30551 (N_30551,N_27671,N_24583);
xor U30552 (N_30552,N_25028,N_26497);
and U30553 (N_30553,N_24991,N_23193);
nor U30554 (N_30554,N_22407,N_21230);
xor U30555 (N_30555,N_24638,N_20833);
nor U30556 (N_30556,N_29943,N_21098);
nor U30557 (N_30557,N_21780,N_26224);
and U30558 (N_30558,N_24808,N_24002);
or U30559 (N_30559,N_23603,N_28685);
nand U30560 (N_30560,N_28010,N_26450);
nor U30561 (N_30561,N_20198,N_27029);
or U30562 (N_30562,N_25036,N_26270);
and U30563 (N_30563,N_29169,N_27445);
and U30564 (N_30564,N_20685,N_21715);
and U30565 (N_30565,N_29197,N_25453);
nor U30566 (N_30566,N_22522,N_21358);
xor U30567 (N_30567,N_27292,N_27968);
xnor U30568 (N_30568,N_21414,N_26301);
xor U30569 (N_30569,N_25715,N_25942);
xor U30570 (N_30570,N_20351,N_29776);
nor U30571 (N_30571,N_23824,N_27996);
xor U30572 (N_30572,N_27890,N_24280);
and U30573 (N_30573,N_26212,N_23129);
nand U30574 (N_30574,N_25874,N_28183);
xor U30575 (N_30575,N_29543,N_22141);
nor U30576 (N_30576,N_20948,N_23064);
nor U30577 (N_30577,N_25841,N_20126);
nor U30578 (N_30578,N_24972,N_27468);
or U30579 (N_30579,N_26039,N_29425);
nor U30580 (N_30580,N_25269,N_24939);
and U30581 (N_30581,N_29162,N_25106);
and U30582 (N_30582,N_21033,N_22567);
and U30583 (N_30583,N_23977,N_21700);
and U30584 (N_30584,N_25634,N_27861);
nor U30585 (N_30585,N_26875,N_20701);
or U30586 (N_30586,N_21723,N_23203);
and U30587 (N_30587,N_22385,N_27269);
nor U30588 (N_30588,N_24719,N_23025);
or U30589 (N_30589,N_23437,N_26649);
and U30590 (N_30590,N_28393,N_22303);
and U30591 (N_30591,N_24203,N_27700);
xor U30592 (N_30592,N_24437,N_28565);
or U30593 (N_30593,N_23233,N_21634);
or U30594 (N_30594,N_25341,N_22676);
nor U30595 (N_30595,N_26752,N_24948);
nor U30596 (N_30596,N_20519,N_23058);
nand U30597 (N_30597,N_29537,N_20952);
or U30598 (N_30598,N_27294,N_20723);
nand U30599 (N_30599,N_24607,N_28242);
nor U30600 (N_30600,N_26229,N_24946);
nor U30601 (N_30601,N_26578,N_25055);
xnor U30602 (N_30602,N_28879,N_27648);
xnor U30603 (N_30603,N_23271,N_20650);
nor U30604 (N_30604,N_26457,N_27952);
and U30605 (N_30605,N_24001,N_28724);
or U30606 (N_30606,N_25110,N_20319);
nor U30607 (N_30607,N_25772,N_28680);
xor U30608 (N_30608,N_24910,N_28993);
xnor U30609 (N_30609,N_23578,N_28439);
nand U30610 (N_30610,N_22618,N_20100);
or U30611 (N_30611,N_21037,N_25988);
or U30612 (N_30612,N_21365,N_28617);
xor U30613 (N_30613,N_22536,N_25683);
nor U30614 (N_30614,N_26595,N_22334);
and U30615 (N_30615,N_26599,N_26474);
nand U30616 (N_30616,N_22949,N_26611);
nand U30617 (N_30617,N_27617,N_29368);
or U30618 (N_30618,N_21149,N_23698);
xnor U30619 (N_30619,N_27563,N_22754);
or U30620 (N_30620,N_22085,N_23943);
nand U30621 (N_30621,N_21977,N_24958);
nor U30622 (N_30622,N_27763,N_27944);
nand U30623 (N_30623,N_20888,N_24126);
xnor U30624 (N_30624,N_25804,N_27815);
or U30625 (N_30625,N_25968,N_21732);
nor U30626 (N_30626,N_27101,N_23510);
and U30627 (N_30627,N_23243,N_28331);
nand U30628 (N_30628,N_20294,N_23825);
xnor U30629 (N_30629,N_26946,N_23846);
nand U30630 (N_30630,N_24118,N_27878);
nand U30631 (N_30631,N_20835,N_20187);
and U30632 (N_30632,N_26511,N_28994);
nor U30633 (N_30633,N_25303,N_28169);
or U30634 (N_30634,N_22808,N_23462);
or U30635 (N_30635,N_28488,N_20849);
nand U30636 (N_30636,N_20511,N_21341);
and U30637 (N_30637,N_21650,N_20640);
nor U30638 (N_30638,N_26098,N_26877);
and U30639 (N_30639,N_29419,N_21420);
xnor U30640 (N_30640,N_27393,N_21329);
nand U30641 (N_30641,N_25791,N_26170);
and U30642 (N_30642,N_28001,N_29290);
nor U30643 (N_30643,N_22023,N_28868);
or U30644 (N_30644,N_28934,N_25413);
nand U30645 (N_30645,N_24859,N_24575);
xor U30646 (N_30646,N_22986,N_27414);
or U30647 (N_30647,N_23591,N_23387);
nand U30648 (N_30648,N_25245,N_24911);
and U30649 (N_30649,N_22973,N_21615);
and U30650 (N_30650,N_29489,N_20914);
nand U30651 (N_30651,N_20942,N_26858);
or U30652 (N_30652,N_28778,N_27354);
or U30653 (N_30653,N_26647,N_26986);
and U30654 (N_30654,N_29320,N_20795);
nand U30655 (N_30655,N_28457,N_21853);
nor U30656 (N_30656,N_24176,N_23364);
nand U30657 (N_30657,N_25552,N_23163);
or U30658 (N_30658,N_21046,N_23763);
and U30659 (N_30659,N_24337,N_23887);
nand U30660 (N_30660,N_24862,N_24100);
nor U30661 (N_30661,N_29839,N_25849);
and U30662 (N_30662,N_20047,N_22397);
nor U30663 (N_30663,N_26416,N_23242);
or U30664 (N_30664,N_25071,N_28988);
and U30665 (N_30665,N_27251,N_22323);
nand U30666 (N_30666,N_28704,N_29086);
nand U30667 (N_30667,N_27775,N_23295);
xor U30668 (N_30668,N_21279,N_27550);
nand U30669 (N_30669,N_21199,N_21476);
or U30670 (N_30670,N_25581,N_28699);
nand U30671 (N_30671,N_28967,N_20800);
xnor U30672 (N_30672,N_29917,N_26653);
or U30673 (N_30673,N_29434,N_26808);
nand U30674 (N_30674,N_22549,N_23140);
nand U30675 (N_30675,N_27516,N_29326);
nor U30676 (N_30676,N_20985,N_29542);
xor U30677 (N_30677,N_28773,N_22894);
xnor U30678 (N_30678,N_26126,N_22465);
nand U30679 (N_30679,N_23612,N_29027);
nor U30680 (N_30680,N_21261,N_25383);
nor U30681 (N_30681,N_26873,N_29665);
and U30682 (N_30682,N_21541,N_26377);
nor U30683 (N_30683,N_26872,N_24602);
xor U30684 (N_30684,N_24364,N_21301);
xor U30685 (N_30685,N_27034,N_27260);
or U30686 (N_30686,N_24535,N_22493);
nor U30687 (N_30687,N_24213,N_27746);
or U30688 (N_30688,N_29858,N_27822);
xor U30689 (N_30689,N_27185,N_29971);
xnor U30690 (N_30690,N_25916,N_29384);
and U30691 (N_30691,N_28626,N_26426);
xor U30692 (N_30692,N_27531,N_24334);
xor U30693 (N_30693,N_24700,N_26681);
nor U30694 (N_30694,N_26466,N_21244);
nand U30695 (N_30695,N_28774,N_23047);
nor U30696 (N_30696,N_20142,N_26790);
nand U30697 (N_30697,N_29216,N_25081);
nand U30698 (N_30698,N_20730,N_21934);
and U30699 (N_30699,N_20565,N_26033);
or U30700 (N_30700,N_25786,N_29978);
nor U30701 (N_30701,N_23985,N_21143);
nor U30702 (N_30702,N_20895,N_22035);
or U30703 (N_30703,N_24936,N_25501);
nor U30704 (N_30704,N_28921,N_20501);
xor U30705 (N_30705,N_29649,N_27515);
nor U30706 (N_30706,N_26503,N_21996);
or U30707 (N_30707,N_26096,N_27566);
nand U30708 (N_30708,N_20858,N_26072);
nor U30709 (N_30709,N_22502,N_27823);
and U30710 (N_30710,N_26294,N_28129);
and U30711 (N_30711,N_20703,N_21877);
and U30712 (N_30712,N_25757,N_27954);
xor U30713 (N_30713,N_24509,N_24836);
or U30714 (N_30714,N_25640,N_20999);
xor U30715 (N_30715,N_26492,N_27122);
nor U30716 (N_30716,N_21773,N_22244);
nor U30717 (N_30717,N_29884,N_26845);
or U30718 (N_30718,N_22115,N_23677);
nand U30719 (N_30719,N_29146,N_25711);
and U30720 (N_30720,N_21453,N_26496);
nor U30721 (N_30721,N_29472,N_25261);
nand U30722 (N_30722,N_26322,N_27594);
xnor U30723 (N_30723,N_24125,N_20078);
nand U30724 (N_30724,N_20193,N_20573);
or U30725 (N_30725,N_28739,N_24781);
xor U30726 (N_30726,N_24817,N_22773);
xnor U30727 (N_30727,N_24062,N_22653);
and U30728 (N_30728,N_29702,N_22178);
and U30729 (N_30729,N_21733,N_25561);
and U30730 (N_30730,N_23624,N_24732);
and U30731 (N_30731,N_21983,N_22241);
nor U30732 (N_30732,N_24525,N_22093);
nor U30733 (N_30733,N_29903,N_20584);
nand U30734 (N_30734,N_26720,N_21418);
or U30735 (N_30735,N_29302,N_24901);
and U30736 (N_30736,N_29403,N_23147);
xor U30737 (N_30737,N_24078,N_29561);
or U30738 (N_30738,N_25537,N_29202);
or U30739 (N_30739,N_21176,N_27774);
xnor U30740 (N_30740,N_29857,N_25771);
xor U30741 (N_30741,N_23951,N_24332);
nor U30742 (N_30742,N_25829,N_26166);
or U30743 (N_30743,N_26171,N_22595);
and U30744 (N_30744,N_29615,N_29328);
or U30745 (N_30745,N_26736,N_23845);
nor U30746 (N_30746,N_23501,N_21497);
nor U30747 (N_30747,N_24667,N_24049);
nor U30748 (N_30748,N_25621,N_23533);
xnor U30749 (N_30749,N_21940,N_20466);
or U30750 (N_30750,N_26487,N_24861);
nor U30751 (N_30751,N_26130,N_26995);
xor U30752 (N_30752,N_22037,N_23194);
or U30753 (N_30753,N_26101,N_24578);
and U30754 (N_30754,N_25556,N_28489);
xor U30755 (N_30755,N_26109,N_29517);
nor U30756 (N_30756,N_21574,N_22622);
xor U30757 (N_30757,N_23150,N_28256);
or U30758 (N_30758,N_24633,N_28756);
and U30759 (N_30759,N_22610,N_27680);
xnor U30760 (N_30760,N_28790,N_20690);
xnor U30761 (N_30761,N_26803,N_29993);
nand U30762 (N_30762,N_23604,N_24788);
xor U30763 (N_30763,N_26175,N_28916);
and U30764 (N_30764,N_24040,N_24159);
and U30765 (N_30765,N_25890,N_27787);
xor U30766 (N_30766,N_28592,N_29714);
or U30767 (N_30767,N_25352,N_28644);
or U30768 (N_30768,N_28474,N_27888);
nor U30769 (N_30769,N_25020,N_20470);
xor U30770 (N_30770,N_23518,N_27027);
nand U30771 (N_30771,N_23402,N_20105);
nand U30772 (N_30772,N_25280,N_26435);
or U30773 (N_30773,N_20222,N_23579);
nand U30774 (N_30774,N_21236,N_26174);
nand U30775 (N_30775,N_20880,N_27002);
nor U30776 (N_30776,N_21874,N_28042);
or U30777 (N_30777,N_28154,N_21248);
and U30778 (N_30778,N_21113,N_28120);
nor U30779 (N_30779,N_24538,N_24655);
and U30780 (N_30780,N_24253,N_26344);
nand U30781 (N_30781,N_20420,N_27471);
xor U30782 (N_30782,N_26374,N_25073);
nand U30783 (N_30783,N_22941,N_27653);
or U30784 (N_30784,N_23685,N_20120);
and U30785 (N_30785,N_21389,N_24333);
and U30786 (N_30786,N_25735,N_27517);
xor U30787 (N_30787,N_29894,N_20507);
or U30788 (N_30788,N_26880,N_29268);
xor U30789 (N_30789,N_23802,N_21254);
or U30790 (N_30790,N_26914,N_21462);
xor U30791 (N_30791,N_26217,N_23352);
and U30792 (N_30792,N_20399,N_21095);
or U30793 (N_30793,N_24965,N_27276);
nand U30794 (N_30794,N_25434,N_25534);
xnor U30795 (N_30795,N_23214,N_24611);
or U30796 (N_30796,N_24970,N_25710);
or U30797 (N_30797,N_27918,N_29950);
nor U30798 (N_30798,N_21976,N_29088);
or U30799 (N_30799,N_22350,N_29787);
or U30800 (N_30800,N_28915,N_24230);
or U30801 (N_30801,N_24550,N_22210);
and U30802 (N_30802,N_28371,N_25563);
xor U30803 (N_30803,N_23381,N_25902);
nor U30804 (N_30804,N_20819,N_28491);
xnor U30805 (N_30805,N_29266,N_29275);
nor U30806 (N_30806,N_23928,N_21827);
nand U30807 (N_30807,N_25591,N_25546);
and U30808 (N_30808,N_28178,N_26050);
and U30809 (N_30809,N_27311,N_20682);
nand U30810 (N_30810,N_24820,N_26339);
and U30811 (N_30811,N_27215,N_25078);
xnor U30812 (N_30812,N_20435,N_25941);
nor U30813 (N_30813,N_26187,N_26771);
nand U30814 (N_30814,N_20964,N_22993);
and U30815 (N_30815,N_20986,N_29979);
and U30816 (N_30816,N_24895,N_22987);
and U30817 (N_30817,N_28382,N_22640);
and U30818 (N_30818,N_22585,N_24257);
nand U30819 (N_30819,N_20877,N_25381);
nor U30820 (N_30820,N_29817,N_28339);
nor U30821 (N_30821,N_25144,N_23694);
and U30822 (N_30822,N_22799,N_25747);
nor U30823 (N_30823,N_26145,N_28787);
or U30824 (N_30824,N_29786,N_23813);
xor U30825 (N_30825,N_25213,N_21239);
nand U30826 (N_30826,N_25235,N_29072);
xnor U30827 (N_30827,N_22223,N_26773);
nand U30828 (N_30828,N_28004,N_22882);
nand U30829 (N_30829,N_28708,N_29183);
and U30830 (N_30830,N_21824,N_29112);
nor U30831 (N_30831,N_21348,N_27179);
nor U30832 (N_30832,N_20534,N_24314);
nor U30833 (N_30833,N_26432,N_29406);
nand U30834 (N_30834,N_28217,N_20676);
xnor U30835 (N_30835,N_23668,N_27051);
or U30836 (N_30836,N_25684,N_20873);
or U30837 (N_30837,N_25318,N_25309);
xnor U30838 (N_30838,N_28614,N_20684);
or U30839 (N_30839,N_28410,N_22187);
nor U30840 (N_30840,N_25822,N_29676);
and U30841 (N_30841,N_26750,N_27457);
or U30842 (N_30842,N_27240,N_25506);
nand U30843 (N_30843,N_21629,N_23550);
and U30844 (N_30844,N_23667,N_24011);
xnor U30845 (N_30845,N_24893,N_26662);
nand U30846 (N_30846,N_21672,N_21611);
or U30847 (N_30847,N_28322,N_22075);
xnor U30848 (N_30848,N_27153,N_26115);
xnor U30849 (N_30849,N_27073,N_24229);
or U30850 (N_30850,N_28806,N_22079);
or U30851 (N_30851,N_28451,N_24366);
and U30852 (N_30852,N_20468,N_25445);
or U30853 (N_30853,N_27816,N_21908);
nand U30854 (N_30854,N_22229,N_25727);
xor U30855 (N_30855,N_26290,N_25094);
nor U30856 (N_30856,N_27394,N_26323);
nor U30857 (N_30857,N_21132,N_24087);
nand U30858 (N_30858,N_28869,N_22553);
and U30859 (N_30859,N_28063,N_24851);
xnor U30860 (N_30860,N_27318,N_28020);
or U30861 (N_30861,N_21029,N_26107);
and U30862 (N_30862,N_25377,N_29458);
nor U30863 (N_30863,N_27176,N_21064);
xnor U30864 (N_30864,N_20081,N_20233);
xor U30865 (N_30865,N_21062,N_26092);
or U30866 (N_30866,N_23077,N_21305);
or U30867 (N_30867,N_20306,N_25686);
or U30868 (N_30868,N_20131,N_24325);
nand U30869 (N_30869,N_28013,N_25054);
xor U30870 (N_30870,N_29944,N_29367);
and U30871 (N_30871,N_28612,N_25810);
and U30872 (N_30872,N_24034,N_28395);
nor U30873 (N_30873,N_22705,N_26785);
or U30874 (N_30874,N_20886,N_24237);
nor U30875 (N_30875,N_26035,N_26934);
xnor U30876 (N_30876,N_27504,N_29685);
nor U30877 (N_30877,N_20652,N_21122);
nand U30878 (N_30878,N_25692,N_27810);
and U30879 (N_30879,N_26844,N_29195);
nand U30880 (N_30880,N_25933,N_25971);
xnor U30881 (N_30881,N_20718,N_23482);
or U30882 (N_30882,N_22914,N_21685);
nor U30883 (N_30883,N_20465,N_22034);
or U30884 (N_30884,N_20551,N_21550);
nand U30885 (N_30885,N_22702,N_29019);
xnor U30886 (N_30886,N_24941,N_28995);
and U30887 (N_30887,N_20058,N_26923);
nand U30888 (N_30888,N_29380,N_28341);
and U30889 (N_30889,N_28190,N_24491);
and U30890 (N_30890,N_21973,N_25620);
and U30891 (N_30891,N_25911,N_21171);
nand U30892 (N_30892,N_23237,N_23054);
or U30893 (N_30893,N_26644,N_28283);
and U30894 (N_30894,N_23026,N_25376);
nor U30895 (N_30895,N_28794,N_24365);
nor U30896 (N_30896,N_26493,N_22485);
nand U30897 (N_30897,N_21105,N_23594);
or U30898 (N_30898,N_21845,N_24447);
xnor U30899 (N_30899,N_28049,N_24871);
or U30900 (N_30900,N_21026,N_27391);
nor U30901 (N_30901,N_24240,N_24177);
nand U30902 (N_30902,N_25708,N_26818);
nor U30903 (N_30903,N_28808,N_27675);
or U30904 (N_30904,N_21793,N_27683);
or U30905 (N_30905,N_22163,N_26838);
nor U30906 (N_30906,N_27797,N_21972);
nor U30907 (N_30907,N_22305,N_24178);
and U30908 (N_30908,N_23840,N_22674);
nand U30909 (N_30909,N_22677,N_25040);
xor U30910 (N_30910,N_22364,N_25197);
nor U30911 (N_30911,N_22781,N_24392);
xor U30912 (N_30912,N_21536,N_25196);
xor U30913 (N_30913,N_20582,N_28225);
nor U30914 (N_30914,N_28082,N_26019);
and U30915 (N_30915,N_26912,N_28914);
nand U30916 (N_30916,N_29526,N_20954);
nor U30917 (N_30917,N_25998,N_23013);
nor U30918 (N_30918,N_20433,N_20355);
nor U30919 (N_30919,N_27505,N_20889);
nor U30920 (N_30920,N_26341,N_23640);
nor U30921 (N_30921,N_27771,N_26658);
and U30922 (N_30922,N_29611,N_20024);
nand U30923 (N_30923,N_23315,N_22457);
xor U30924 (N_30924,N_22637,N_28342);
or U30925 (N_30925,N_26246,N_21854);
or U30926 (N_30926,N_20707,N_21850);
nand U30927 (N_30927,N_20554,N_21455);
or U30928 (N_30928,N_22422,N_26560);
or U30929 (N_30929,N_25237,N_29071);
nor U30930 (N_30930,N_29455,N_20218);
and U30931 (N_30931,N_20245,N_24192);
or U30932 (N_30932,N_27601,N_23219);
nand U30933 (N_30933,N_26252,N_29272);
xnor U30934 (N_30934,N_29942,N_21691);
xnor U30935 (N_30935,N_27211,N_25409);
xor U30936 (N_30936,N_20957,N_25995);
and U30937 (N_30937,N_22125,N_28289);
nand U30938 (N_30938,N_23262,N_26343);
or U30939 (N_30939,N_28326,N_23691);
nor U30940 (N_30940,N_24774,N_25316);
and U30941 (N_30941,N_24167,N_25011);
nor U30942 (N_30942,N_23706,N_24391);
and U30943 (N_30943,N_27526,N_21878);
nor U30944 (N_30944,N_20512,N_25759);
xor U30945 (N_30945,N_24402,N_28441);
nor U30946 (N_30946,N_26707,N_28505);
and U30947 (N_30947,N_24415,N_29047);
nor U30948 (N_30948,N_28803,N_24985);
nor U30949 (N_30949,N_27647,N_20523);
and U30950 (N_30950,N_22256,N_26586);
or U30951 (N_30951,N_29546,N_25619);
xnor U30952 (N_30952,N_28452,N_20761);
and U30953 (N_30953,N_20447,N_22452);
xnor U30954 (N_30954,N_27976,N_23976);
xnor U30955 (N_30955,N_27624,N_20286);
or U30956 (N_30956,N_26446,N_24113);
and U30957 (N_30957,N_27059,N_27305);
and U30958 (N_30958,N_22142,N_28030);
or U30959 (N_30959,N_27652,N_27083);
nor U30960 (N_30960,N_23778,N_29467);
nand U30961 (N_30961,N_24858,N_26369);
or U30962 (N_30962,N_25814,N_21584);
nor U30963 (N_30963,N_26878,N_20503);
or U30964 (N_30964,N_26766,N_27603);
and U30965 (N_30965,N_25164,N_27838);
nor U30966 (N_30966,N_27757,N_23346);
nand U30967 (N_30967,N_27743,N_29098);
nand U30968 (N_30968,N_27223,N_24951);
xor U30969 (N_30969,N_25037,N_27872);
nand U30970 (N_30970,N_21432,N_21030);
xor U30971 (N_30971,N_21653,N_21484);
and U30972 (N_30972,N_22435,N_28619);
xnor U30973 (N_30973,N_23060,N_20679);
or U30974 (N_30974,N_22665,N_28473);
nor U30975 (N_30975,N_20513,N_21011);
xor U30976 (N_30976,N_29521,N_27441);
nand U30977 (N_30977,N_22528,N_27241);
nand U30978 (N_30978,N_27197,N_20348);
and U30979 (N_30979,N_28432,N_21837);
nand U30980 (N_30980,N_21251,N_22907);
or U30981 (N_30981,N_25420,N_25496);
or U30982 (N_30982,N_20171,N_26922);
and U30983 (N_30983,N_24200,N_29062);
nand U30984 (N_30984,N_23934,N_29540);
nand U30985 (N_30985,N_23713,N_20638);
nor U30986 (N_30986,N_23251,N_20206);
nand U30987 (N_30987,N_27596,N_28051);
nand U30988 (N_30988,N_26622,N_24921);
nand U30989 (N_30989,N_22872,N_21478);
or U30990 (N_30990,N_26291,N_20706);
nand U30991 (N_30991,N_25191,N_20635);
and U30992 (N_30992,N_21711,N_20724);
xor U30993 (N_30993,N_29281,N_22790);
or U30994 (N_30994,N_27009,N_26606);
and U30995 (N_30995,N_20771,N_29912);
nand U30996 (N_30996,N_27987,N_26856);
and U30997 (N_30997,N_23988,N_28301);
nor U30998 (N_30998,N_24691,N_22942);
xnor U30999 (N_30999,N_24008,N_26634);
or U31000 (N_31000,N_20863,N_24686);
nor U31001 (N_31001,N_25134,N_25828);
and U31002 (N_31002,N_28421,N_22803);
nand U31003 (N_31003,N_29559,N_21851);
nor U31004 (N_31004,N_27853,N_24625);
and U31005 (N_31005,N_22730,N_29315);
and U31006 (N_31006,N_28703,N_26727);
nor U31007 (N_31007,N_25096,N_26952);
xor U31008 (N_31008,N_28497,N_26842);
xor U31009 (N_31009,N_22950,N_20813);
nor U31010 (N_31010,N_23230,N_21626);
or U31011 (N_31011,N_28897,N_26970);
xnor U31012 (N_31012,N_28812,N_23946);
nand U31013 (N_31013,N_29323,N_25082);
and U31014 (N_31014,N_28840,N_25630);
nor U31015 (N_31015,N_23867,N_23981);
and U31016 (N_31016,N_20343,N_22269);
xnor U31017 (N_31017,N_27023,N_29341);
and U31018 (N_31018,N_28492,N_26287);
xnor U31019 (N_31019,N_21145,N_29110);
nor U31020 (N_31020,N_29330,N_21016);
or U31021 (N_31021,N_27378,N_20916);
or U31022 (N_31022,N_22521,N_27407);
nand U31023 (N_31023,N_27422,N_26310);
or U31024 (N_31024,N_24063,N_26049);
nor U31025 (N_31025,N_27633,N_21047);
or U31026 (N_31026,N_25262,N_20661);
and U31027 (N_31027,N_26898,N_25987);
or U31028 (N_31028,N_22841,N_23290);
or U31029 (N_31029,N_25218,N_21501);
nand U31030 (N_31030,N_23365,N_21817);
and U31031 (N_31031,N_24644,N_20555);
or U31032 (N_31032,N_20599,N_21721);
nand U31033 (N_31033,N_22340,N_22208);
or U31034 (N_31034,N_21950,N_27802);
and U31035 (N_31035,N_23733,N_29201);
xnor U31036 (N_31036,N_22992,N_20570);
xor U31037 (N_31037,N_21714,N_21324);
nand U31038 (N_31038,N_26538,N_20788);
or U31039 (N_31039,N_24727,N_20201);
nand U31040 (N_31040,N_23700,N_25424);
nor U31041 (N_31041,N_20945,N_28526);
nand U31042 (N_31042,N_26902,N_29369);
or U31043 (N_31043,N_24886,N_21445);
or U31044 (N_31044,N_21410,N_25853);
or U31045 (N_31045,N_20380,N_27174);
and U31046 (N_31046,N_29205,N_27923);
and U31047 (N_31047,N_20947,N_24072);
and U31048 (N_31048,N_25569,N_21200);
and U31049 (N_31049,N_27587,N_26890);
nand U31050 (N_31050,N_26930,N_23438);
or U31051 (N_31051,N_23647,N_25796);
and U31052 (N_31052,N_22048,N_27584);
and U31053 (N_31053,N_27282,N_24761);
or U31054 (N_31054,N_26621,N_28559);
nor U31055 (N_31055,N_29075,N_26165);
nand U31056 (N_31056,N_22077,N_26507);
nor U31057 (N_31057,N_27752,N_24899);
nand U31058 (N_31058,N_27134,N_23120);
nand U31059 (N_31059,N_21635,N_25304);
nor U31060 (N_31060,N_21676,N_24051);
and U31061 (N_31061,N_27590,N_24241);
nor U31062 (N_31062,N_23329,N_25639);
xnor U31063 (N_31063,N_20760,N_25691);
xnor U31064 (N_31064,N_21218,N_23130);
or U31065 (N_31065,N_20909,N_26430);
and U31066 (N_31066,N_20018,N_23842);
and U31067 (N_31067,N_29142,N_28138);
nand U31068 (N_31068,N_29309,N_23085);
or U31069 (N_31069,N_28872,N_23689);
nand U31070 (N_31070,N_20263,N_24617);
xnor U31071 (N_31071,N_25247,N_25184);
xnor U31072 (N_31072,N_25339,N_28797);
xor U31073 (N_31073,N_25512,N_24653);
or U31074 (N_31074,N_25085,N_20457);
nand U31075 (N_31075,N_29541,N_26604);
and U31076 (N_31076,N_27049,N_25937);
nor U31077 (N_31077,N_27969,N_27213);
or U31078 (N_31078,N_21919,N_21274);
and U31079 (N_31079,N_22202,N_29882);
and U31080 (N_31080,N_26158,N_26835);
and U31081 (N_31081,N_28853,N_26666);
nand U31082 (N_31082,N_27062,N_27306);
nand U31083 (N_31083,N_23834,N_21958);
or U31084 (N_31084,N_24393,N_20101);
and U31085 (N_31085,N_25313,N_23744);
nor U31086 (N_31086,N_22740,N_23505);
nand U31087 (N_31087,N_27415,N_26897);
nor U31088 (N_31088,N_26630,N_28906);
or U31089 (N_31089,N_25539,N_26265);
xnor U31090 (N_31090,N_27184,N_22578);
nand U31091 (N_31091,N_22614,N_24744);
and U31092 (N_31092,N_22481,N_26828);
and U31093 (N_31093,N_23433,N_29186);
and U31094 (N_31094,N_22604,N_20590);
nor U31095 (N_31095,N_22461,N_20798);
nand U31096 (N_31096,N_26561,N_24157);
and U31097 (N_31097,N_26071,N_21856);
nand U31098 (N_31098,N_23080,N_28735);
xnor U31099 (N_31099,N_27261,N_21869);
or U31100 (N_31100,N_23326,N_25240);
xor U31101 (N_31101,N_28222,N_28095);
nand U31102 (N_31102,N_25348,N_21707);
xnor U31103 (N_31103,N_22963,N_21822);
xor U31104 (N_31104,N_22406,N_27012);
nand U31105 (N_31105,N_21231,N_24669);
or U31106 (N_31106,N_26220,N_24141);
or U31107 (N_31107,N_23159,N_26676);
or U31108 (N_31108,N_22775,N_28728);
nor U31109 (N_31109,N_22962,N_22450);
nor U31110 (N_31110,N_29121,N_22017);
or U31111 (N_31111,N_27239,N_25785);
and U31112 (N_31112,N_27932,N_27400);
or U31113 (N_31113,N_26613,N_22657);
nand U31114 (N_31114,N_23021,N_24110);
or U31115 (N_31115,N_20756,N_22227);
or U31116 (N_31116,N_23278,N_28134);
or U31117 (N_31117,N_26479,N_26114);
nand U31118 (N_31118,N_21110,N_24343);
xor U31119 (N_31119,N_23962,N_20840);
and U31120 (N_31120,N_25138,N_24785);
and U31121 (N_31121,N_23457,N_20119);
or U31122 (N_31122,N_26144,N_27638);
and U31123 (N_31123,N_20606,N_28527);
xor U31124 (N_31124,N_26868,N_27019);
or U31125 (N_31125,N_29716,N_25385);
and U31126 (N_31126,N_23113,N_20875);
xnor U31127 (N_31127,N_22434,N_23177);
and U31128 (N_31128,N_21458,N_28689);
xor U31129 (N_31129,N_24735,N_21583);
or U31130 (N_31130,N_28604,N_25286);
xor U31131 (N_31131,N_28427,N_28665);
xnor U31132 (N_31132,N_23657,N_24464);
xnor U31133 (N_31133,N_22999,N_20874);
nor U31134 (N_31134,N_25222,N_23752);
nand U31135 (N_31135,N_20912,N_25935);
xor U31136 (N_31136,N_27351,N_20413);
nor U31137 (N_31137,N_25965,N_20426);
xnor U31138 (N_31138,N_24683,N_24137);
nand U31139 (N_31139,N_22921,N_21479);
and U31140 (N_31140,N_29017,N_22284);
xor U31141 (N_31141,N_28849,N_29713);
or U31142 (N_31142,N_21373,N_22492);
nand U31143 (N_31143,N_25189,N_24736);
nand U31144 (N_31144,N_22408,N_29575);
xnor U31145 (N_31145,N_20141,N_23644);
and U31146 (N_31146,N_20203,N_20393);
nor U31147 (N_31147,N_22330,N_21598);
nor U31148 (N_31148,N_20854,N_25909);
or U31149 (N_31149,N_25104,N_20353);
xnor U31150 (N_31150,N_23112,N_27453);
xor U31151 (N_31151,N_23409,N_24758);
or U31152 (N_31152,N_20831,N_21597);
nor U31153 (N_31153,N_28184,N_28117);
and U31154 (N_31154,N_29105,N_21569);
nand U31155 (N_31155,N_21179,N_29593);
xnor U31156 (N_31156,N_23492,N_25671);
or U31157 (N_31157,N_29700,N_21965);
or U31158 (N_31158,N_21013,N_21918);
nand U31159 (N_31159,N_22889,N_25010);
nor U31160 (N_31160,N_27387,N_24714);
and U31161 (N_31161,N_25967,N_23355);
nand U31162 (N_31162,N_22983,N_26629);
and U31163 (N_31163,N_28501,N_20320);
or U31164 (N_31164,N_22174,N_26251);
xnor U31165 (N_31165,N_21966,N_22021);
xnor U31166 (N_31166,N_25008,N_24021);
nor U31167 (N_31167,N_29793,N_22314);
nand U31168 (N_31168,N_22424,N_23989);
nor U31169 (N_31169,N_29119,N_25229);
nor U31170 (N_31170,N_29798,N_29198);
nor U31171 (N_31171,N_27761,N_20572);
xor U31172 (N_31172,N_25050,N_24215);
and U31173 (N_31173,N_24196,N_27060);
nor U31174 (N_31174,N_25360,N_21111);
and U31175 (N_31175,N_29494,N_24765);
and U31176 (N_31176,N_27906,N_22327);
nor U31177 (N_31177,N_28102,N_21091);
nor U31178 (N_31178,N_25283,N_27629);
and U31179 (N_31179,N_27728,N_25862);
nor U31180 (N_31180,N_26082,N_23282);
or U31181 (N_31181,N_24467,N_29850);
xnor U31182 (N_31182,N_22680,N_20804);
nand U31183 (N_31183,N_29777,N_22924);
or U31184 (N_31184,N_23532,N_28355);
and U31185 (N_31185,N_22542,N_23361);
nor U31186 (N_31186,N_28648,N_23405);
nand U31187 (N_31187,N_24386,N_25894);
or U31188 (N_31188,N_21310,N_25108);
xnor U31189 (N_31189,N_22218,N_23935);
and U31190 (N_31190,N_22645,N_28046);
nand U31191 (N_31191,N_23107,N_22057);
nor U31192 (N_31192,N_28839,N_26282);
xnor U31193 (N_31193,N_29670,N_27150);
and U31194 (N_31194,N_28727,N_20292);
or U31195 (N_31195,N_29579,N_25794);
or U31196 (N_31196,N_20409,N_27655);
nor U31197 (N_31197,N_21936,N_20235);
xor U31198 (N_31198,N_28636,N_23336);
or U31199 (N_31199,N_20221,N_21081);
xor U31200 (N_31200,N_27783,N_27591);
xor U31201 (N_31201,N_29357,N_28434);
nand U31202 (N_31202,N_23641,N_25737);
nor U31203 (N_31203,N_20397,N_29982);
nand U31204 (N_31204,N_23723,N_23673);
and U31205 (N_31205,N_27224,N_26267);
nor U31206 (N_31206,N_26292,N_28855);
or U31207 (N_31207,N_26436,N_24520);
nand U31208 (N_31208,N_29814,N_28440);
nand U31209 (N_31209,N_27475,N_22602);
nor U31210 (N_31210,N_25417,N_23793);
or U31211 (N_31211,N_22910,N_21843);
nand U31212 (N_31212,N_26944,N_25495);
or U31213 (N_31213,N_22660,N_23728);
nor U31214 (N_31214,N_26833,N_23741);
and U31215 (N_31215,N_22288,N_29113);
nor U31216 (N_31216,N_26068,N_26959);
nor U31217 (N_31217,N_23947,N_25075);
and U31218 (N_31218,N_27301,N_26385);
nand U31219 (N_31219,N_27216,N_25734);
xnor U31220 (N_31220,N_28271,N_27430);
nand U31221 (N_31221,N_21807,N_28965);
xor U31222 (N_31222,N_23419,N_23528);
or U31223 (N_31223,N_27409,N_28156);
xor U31224 (N_31224,N_20098,N_23584);
nor U31225 (N_31225,N_25722,N_28390);
or U31226 (N_31226,N_29037,N_24012);
nor U31227 (N_31227,N_20311,N_27519);
or U31228 (N_31228,N_22737,N_21863);
or U31229 (N_31229,N_28479,N_27462);
xnor U31230 (N_31230,N_28340,N_22648);
xnor U31231 (N_31231,N_26732,N_27814);
and U31232 (N_31232,N_26081,N_29415);
xor U31233 (N_31233,N_23141,N_25001);
nand U31234 (N_31234,N_26515,N_29641);
nand U31235 (N_31235,N_24755,N_24721);
nor U31236 (N_31236,N_27245,N_26117);
xor U31237 (N_31237,N_27267,N_21277);
xor U31238 (N_31238,N_25282,N_20714);
or U31239 (N_31239,N_29726,N_29624);
or U31240 (N_31240,N_24837,N_23567);
xor U31241 (N_31241,N_20417,N_28358);
nand U31242 (N_31242,N_20755,N_22547);
xnor U31243 (N_31243,N_29022,N_20087);
and U31244 (N_31244,N_25112,N_25598);
and U31245 (N_31245,N_26397,N_27600);
nor U31246 (N_31246,N_24950,N_24830);
nor U31247 (N_31247,N_28296,N_20751);
or U31248 (N_31248,N_24449,N_29030);
nor U31249 (N_31249,N_27619,N_28198);
or U31250 (N_31250,N_27809,N_27864);
or U31251 (N_31251,N_22890,N_23169);
or U31252 (N_31252,N_28740,N_28223);
nor U31253 (N_31253,N_21696,N_25437);
nand U31254 (N_31254,N_27113,N_29506);
xor U31255 (N_31255,N_28351,N_21170);
nor U31256 (N_31256,N_22374,N_21749);
nor U31257 (N_31257,N_23769,N_21661);
and U31258 (N_31258,N_22080,N_22556);
nor U31259 (N_31259,N_26053,N_25513);
xor U31260 (N_31260,N_23487,N_22791);
or U31261 (N_31261,N_21396,N_28946);
or U31262 (N_31262,N_27484,N_20737);
nand U31263 (N_31263,N_29754,N_27889);
and U31264 (N_31264,N_23359,N_25548);
nor U31265 (N_31265,N_25609,N_21588);
and U31266 (N_31266,N_22631,N_21762);
nor U31267 (N_31267,N_26472,N_20732);
nand U31268 (N_31268,N_25760,N_24606);
or U31269 (N_31269,N_29296,N_28701);
and U31270 (N_31270,N_29692,N_29930);
or U31271 (N_31271,N_22855,N_20884);
xnor U31272 (N_31272,N_29140,N_28607);
or U31273 (N_31273,N_24690,N_21249);
and U31274 (N_31274,N_27358,N_25553);
or U31275 (N_31275,N_21296,N_28239);
or U31276 (N_31276,N_26490,N_26849);
xor U31277 (N_31277,N_27020,N_29150);
nand U31278 (N_31278,N_25276,N_29254);
nand U31279 (N_31279,N_29291,N_29387);
and U31280 (N_31280,N_28595,N_28824);
nand U31281 (N_31281,N_29591,N_25427);
nand U31282 (N_31282,N_29637,N_21424);
xnor U31283 (N_31283,N_26809,N_24387);
xor U31284 (N_31284,N_29299,N_28369);
or U31285 (N_31285,N_26262,N_27719);
or U31286 (N_31286,N_26941,N_22634);
nor U31287 (N_31287,N_21270,N_20121);
or U31288 (N_31288,N_26813,N_21423);
or U31289 (N_31289,N_26543,N_29064);
or U31290 (N_31290,N_26755,N_29392);
xor U31291 (N_31291,N_22825,N_25322);
nor U31292 (N_31292,N_22182,N_25950);
xor U31293 (N_31293,N_26241,N_27386);
nand U31294 (N_31294,N_28593,N_25956);
xor U31295 (N_31295,N_25241,N_29428);
nor U31296 (N_31296,N_21872,N_25590);
and U31297 (N_31297,N_29783,N_23454);
nand U31298 (N_31298,N_27022,N_26173);
nand U31299 (N_31299,N_21832,N_28930);
and U31300 (N_31300,N_22590,N_28757);
and U31301 (N_31301,N_26953,N_28413);
or U31302 (N_31302,N_22978,N_20366);
and U31303 (N_31303,N_24056,N_22718);
nand U31304 (N_31304,N_21651,N_23630);
nand U31305 (N_31305,N_29823,N_25816);
or U31306 (N_31306,N_24791,N_29450);
nand U31307 (N_31307,N_24355,N_21315);
nor U31308 (N_31308,N_29530,N_24891);
nand U31309 (N_31309,N_25351,N_22173);
and U31310 (N_31310,N_21967,N_24140);
nor U31311 (N_31311,N_21306,N_20841);
and U31312 (N_31312,N_26699,N_24707);
xnor U31313 (N_31313,N_29799,N_24478);
or U31314 (N_31314,N_27527,N_20994);
xnor U31315 (N_31315,N_25960,N_23507);
and U31316 (N_31316,N_22526,N_28650);
nand U31317 (N_31317,N_24532,N_26737);
xnor U31318 (N_31318,N_26916,N_20136);
and U31319 (N_31319,N_27111,N_20395);
nor U31320 (N_31320,N_27836,N_27090);
nand U31321 (N_31321,N_24679,N_25606);
and U31322 (N_31322,N_27800,N_29588);
nand U31323 (N_31323,N_29689,N_23406);
and U31324 (N_31324,N_23467,N_24767);
nor U31325 (N_31325,N_21573,N_22832);
nand U31326 (N_31326,N_21437,N_26296);
or U31327 (N_31327,N_26579,N_24256);
nor U31328 (N_31328,N_23102,N_20239);
or U31329 (N_31329,N_22322,N_22995);
or U31330 (N_31330,N_23043,N_22226);
xor U31331 (N_31331,N_28170,N_25802);
and U31332 (N_31332,N_29067,N_21810);
or U31333 (N_31333,N_27493,N_25368);
or U31334 (N_31334,N_21620,N_21017);
or U31335 (N_31335,N_24296,N_23660);
and U31336 (N_31336,N_23415,N_24232);
nor U31337 (N_31337,N_24081,N_27699);
nor U31338 (N_31338,N_26832,N_24598);
nand U31339 (N_31339,N_24495,N_27646);
or U31340 (N_31340,N_22453,N_27636);
nor U31341 (N_31341,N_24376,N_29365);
nand U31342 (N_31342,N_22294,N_26411);
nand U31343 (N_31343,N_23748,N_20602);
nor U31344 (N_31344,N_21258,N_22478);
or U31345 (N_31345,N_27191,N_26116);
and U31346 (N_31346,N_27998,N_20025);
nand U31347 (N_31347,N_23450,N_26906);
nand U31348 (N_31348,N_20577,N_28480);
nor U31349 (N_31349,N_25043,N_29347);
and U31350 (N_31350,N_24797,N_28112);
or U31351 (N_31351,N_24696,N_24877);
nor U31352 (N_31352,N_23200,N_27030);
and U31353 (N_31353,N_22879,N_23992);
or U31354 (N_31354,N_24554,N_28148);
xor U31355 (N_31355,N_24329,N_28107);
xor U31356 (N_31356,N_20471,N_21173);
xor U31357 (N_31357,N_27753,N_20710);
nand U31358 (N_31358,N_21359,N_21382);
nor U31359 (N_31359,N_29122,N_29722);
or U31360 (N_31360,N_28815,N_24807);
xnor U31361 (N_31361,N_26920,N_29476);
nor U31362 (N_31362,N_23617,N_23637);
or U31363 (N_31363,N_24703,N_28718);
nor U31364 (N_31364,N_24833,N_22392);
nand U31365 (N_31365,N_25953,N_26148);
nand U31366 (N_31366,N_24574,N_26660);
xor U31367 (N_31367,N_29233,N_22709);
xor U31368 (N_31368,N_21681,N_20029);
nand U31369 (N_31369,N_28008,N_22005);
or U31370 (N_31370,N_23937,N_26278);
nand U31371 (N_31371,N_28064,N_29809);
nor U31372 (N_31372,N_23849,N_27908);
or U31373 (N_31373,N_29638,N_29123);
xor U31374 (N_31374,N_22989,N_23654);
or U31375 (N_31375,N_21990,N_23633);
nand U31376 (N_31376,N_21991,N_25740);
xnor U31377 (N_31377,N_26958,N_20497);
nor U31378 (N_31378,N_24371,N_27965);
xnor U31379 (N_31379,N_27845,N_21287);
and U31380 (N_31380,N_25575,N_23240);
or U31381 (N_31381,N_29584,N_28742);
nand U31382 (N_31382,N_24772,N_26715);
xor U31383 (N_31383,N_28972,N_27388);
xor U31384 (N_31384,N_24541,N_20564);
or U31385 (N_31385,N_28954,N_21136);
xnor U31386 (N_31386,N_20583,N_29354);
or U31387 (N_31387,N_25679,N_22880);
or U31388 (N_31388,N_28519,N_25643);
or U31389 (N_31389,N_21735,N_20810);
nand U31390 (N_31390,N_22923,N_25508);
or U31391 (N_31391,N_24570,N_22554);
nand U31392 (N_31392,N_25419,N_20321);
nor U31393 (N_31393,N_20814,N_20085);
nand U31394 (N_31394,N_28980,N_26157);
or U31395 (N_31395,N_21981,N_29469);
and U31396 (N_31396,N_28050,N_25917);
or U31397 (N_31397,N_25963,N_26888);
or U31398 (N_31398,N_29636,N_26978);
nand U31399 (N_31399,N_24728,N_22956);
nand U31400 (N_31400,N_20373,N_20135);
and U31401 (N_31401,N_26895,N_28173);
xor U31402 (N_31402,N_21102,N_20528);
xnor U31403 (N_31403,N_20496,N_27203);
nand U31404 (N_31404,N_20961,N_20146);
nand U31405 (N_31405,N_22064,N_20130);
nor U31406 (N_31406,N_22328,N_26594);
or U31407 (N_31407,N_28600,N_20458);
or U31408 (N_31408,N_20096,N_21813);
nand U31409 (N_31409,N_23546,N_27668);
or U31410 (N_31410,N_25962,N_24179);
or U31411 (N_31411,N_24944,N_27390);
or U31412 (N_31412,N_24024,N_28003);
nand U31413 (N_31413,N_26881,N_24428);
nand U31414 (N_31414,N_29060,N_21207);
or U31415 (N_31415,N_29381,N_21935);
nor U31416 (N_31416,N_26680,N_25632);
and U31417 (N_31417,N_24605,N_28255);
and U31418 (N_31418,N_23217,N_24713);
nand U31419 (N_31419,N_22011,N_25289);
nor U31420 (N_31420,N_24058,N_25153);
and U31421 (N_31421,N_29294,N_29273);
and U31422 (N_31422,N_21448,N_28437);
and U31423 (N_31423,N_27712,N_24265);
xor U31424 (N_31424,N_25460,N_22052);
xnor U31425 (N_31425,N_21084,N_21513);
nand U31426 (N_31426,N_20086,N_29271);
or U31427 (N_31427,N_27983,N_20123);
nand U31428 (N_31428,N_20878,N_20514);
nor U31429 (N_31429,N_26863,N_24770);
or U31430 (N_31430,N_20949,N_29875);
nor U31431 (N_31431,N_29295,N_21446);
and U31432 (N_31432,N_26521,N_25654);
nand U31433 (N_31433,N_25321,N_25656);
nor U31434 (N_31434,N_24271,N_29492);
and U31435 (N_31435,N_29093,N_22616);
or U31436 (N_31436,N_25657,N_24022);
xnor U31437 (N_31437,N_23734,N_27040);
xnor U31438 (N_31438,N_23048,N_23396);
nor U31439 (N_31439,N_25623,N_20302);
xnor U31440 (N_31440,N_20216,N_23952);
nand U31441 (N_31441,N_20892,N_26394);
nand U31442 (N_31442,N_28819,N_26364);
xnor U31443 (N_31443,N_28291,N_24276);
and U31444 (N_31444,N_28158,N_24567);
or U31445 (N_31445,N_29411,N_23678);
or U31446 (N_31446,N_25099,N_21875);
xnor U31447 (N_31447,N_28903,N_25879);
nand U31448 (N_31448,N_24135,N_28352);
or U31449 (N_31449,N_22788,N_22876);
or U31450 (N_31450,N_28389,N_28746);
nand U31451 (N_31451,N_27875,N_28656);
nand U31452 (N_31452,N_23717,N_23618);
xor U31453 (N_31453,N_28085,N_21871);
and U31454 (N_31454,N_21604,N_24490);
and U31455 (N_31455,N_21790,N_23915);
and U31456 (N_31456,N_25421,N_23007);
and U31457 (N_31457,N_21093,N_29066);
or U31458 (N_31458,N_23939,N_24254);
or U31459 (N_31459,N_29525,N_23390);
and U31460 (N_31460,N_27794,N_22313);
and U31461 (N_31461,N_29968,N_22399);
nand U31462 (N_31462,N_29715,N_29180);
or U31463 (N_31463,N_27234,N_25448);
and U31464 (N_31464,N_20866,N_26665);
and U31465 (N_31465,N_24248,N_27607);
or U31466 (N_31466,N_29892,N_29888);
xnor U31467 (N_31467,N_26080,N_21128);
nor U31468 (N_31468,N_24272,N_24892);
or U31469 (N_31469,N_21209,N_27188);
or U31470 (N_31470,N_23819,N_22688);
and U31471 (N_31471,N_24190,N_25642);
nand U31472 (N_31472,N_21377,N_21521);
and U31473 (N_31473,N_24340,N_27666);
nor U31474 (N_31474,N_25314,N_24885);
and U31475 (N_31475,N_23897,N_21743);
and U31476 (N_31476,N_23747,N_24582);
nand U31477 (N_31477,N_27421,N_29448);
and U31478 (N_31478,N_20334,N_28702);
and U31479 (N_31479,N_22623,N_27170);
xor U31480 (N_31480,N_28450,N_29400);
or U31481 (N_31481,N_25101,N_21401);
or U31482 (N_31482,N_20350,N_29389);
nor U31483 (N_31483,N_25366,N_29974);
nor U31484 (N_31484,N_28630,N_25724);
xor U31485 (N_31485,N_27427,N_21907);
and U31486 (N_31486,N_22237,N_24460);
or U31487 (N_31487,N_27623,N_26823);
xor U31488 (N_31488,N_26563,N_21978);
nor U31489 (N_31489,N_21909,N_26764);
nand U31490 (N_31490,N_27789,N_23568);
nand U31491 (N_31491,N_25211,N_27127);
and U31492 (N_31492,N_26318,N_24983);
or U31493 (N_31493,N_21921,N_21533);
nand U31494 (N_31494,N_23696,N_23488);
nand U31495 (N_31495,N_26348,N_29684);
nand U31496 (N_31496,N_25661,N_21689);
or U31497 (N_31497,N_28140,N_22445);
xor U31498 (N_31498,N_29557,N_20372);
and U31499 (N_31499,N_26298,N_20460);
nor U31500 (N_31500,N_22875,N_21867);
nor U31501 (N_31501,N_22667,N_21404);
and U31502 (N_31502,N_21210,N_23719);
nand U31503 (N_31503,N_29585,N_23716);
and U31504 (N_31504,N_25062,N_28032);
or U31505 (N_31505,N_24170,N_21433);
xor U31506 (N_31506,N_22378,N_27911);
nand U31507 (N_31507,N_25705,N_21920);
and U31508 (N_31508,N_22290,N_24264);
nor U31509 (N_31509,N_27472,N_29185);
or U31510 (N_31510,N_20940,N_28691);
and U31511 (N_31511,N_24759,N_23436);
xor U31512 (N_31512,N_28094,N_22831);
nand U31513 (N_31513,N_25033,N_21428);
nand U31514 (N_31514,N_22658,N_27748);
xnor U31515 (N_31515,N_21280,N_26797);
xnor U31516 (N_31516,N_24884,N_27580);
or U31517 (N_31517,N_28659,N_29422);
xor U31518 (N_31518,N_20832,N_23051);
xor U31519 (N_31519,N_27895,N_24270);
or U31520 (N_31520,N_28108,N_21809);
and U31521 (N_31521,N_25395,N_23089);
and U31522 (N_31522,N_29331,N_23949);
nor U31523 (N_31523,N_28989,N_25077);
and U31524 (N_31524,N_25596,N_26402);
or U31525 (N_31525,N_22231,N_25068);
xor U31526 (N_31526,N_22307,N_21442);
nand U31527 (N_31527,N_23151,N_29396);
xor U31528 (N_31528,N_28532,N_22076);
nand U31529 (N_31529,N_24148,N_28948);
nand U31530 (N_31530,N_27972,N_27121);
nand U31531 (N_31531,N_28979,N_20972);
nor U31532 (N_31532,N_20191,N_21079);
nand U31533 (N_31533,N_21797,N_22650);
nor U31534 (N_31534,N_24857,N_21357);
and U31535 (N_31535,N_23489,N_27106);
nor U31536 (N_31536,N_21592,N_27844);
and U31537 (N_31537,N_21399,N_22529);
or U31538 (N_31538,N_29785,N_27165);
and U31539 (N_31539,N_27360,N_22996);
nor U31540 (N_31540,N_26729,N_21465);
or U31541 (N_31541,N_22049,N_28396);
nor U31542 (N_31542,N_23519,N_26651);
nor U31543 (N_31543,N_27016,N_23693);
nor U31544 (N_31544,N_25477,N_20537);
and U31545 (N_31545,N_25013,N_29534);
nand U31546 (N_31546,N_27994,N_21730);
or U31547 (N_31547,N_20463,N_22870);
or U31548 (N_31548,N_29010,N_27433);
or U31549 (N_31549,N_25861,N_25478);
xor U31550 (N_31550,N_21624,N_24459);
or U31551 (N_31551,N_20656,N_29133);
nor U31552 (N_31552,N_25034,N_26403);
xor U31553 (N_31553,N_24935,N_25159);
or U31554 (N_31554,N_23117,N_27325);
nor U31555 (N_31555,N_23035,N_21347);
nand U31556 (N_31556,N_26141,N_24436);
and U31557 (N_31557,N_20170,N_28635);
xnor U31558 (N_31558,N_28784,N_20941);
nor U31559 (N_31559,N_24513,N_27081);
xnor U31560 (N_31560,N_25285,N_22062);
xnor U31561 (N_31561,N_23593,N_27167);
xor U31562 (N_31562,N_29806,N_28935);
or U31563 (N_31563,N_29573,N_25178);
or U31564 (N_31564,N_22137,N_26342);
nor U31565 (N_31565,N_27208,N_29148);
xor U31566 (N_31566,N_27595,N_24142);
xor U31567 (N_31567,N_21820,N_29536);
xnor U31568 (N_31568,N_20580,N_22836);
and U31569 (N_31569,N_24731,N_27807);
xnor U31570 (N_31570,N_28975,N_29755);
xnor U31571 (N_31571,N_21402,N_23431);
nor U31572 (N_31572,N_29339,N_29308);
nor U31573 (N_31573,N_22661,N_23817);
and U31574 (N_31574,N_20838,N_28628);
nor U31575 (N_31575,N_21776,N_24933);
nor U31576 (N_31576,N_27135,N_25200);
xor U31577 (N_31577,N_25450,N_21114);
or U31578 (N_31578,N_28577,N_29671);
and U31579 (N_31579,N_22904,N_29550);
xor U31580 (N_31580,N_25203,N_27095);
or U31581 (N_31581,N_27520,N_24093);
and U31582 (N_31582,N_27265,N_28221);
or U31583 (N_31583,N_20740,N_29570);
nor U31584 (N_31584,N_26362,N_24061);
and U31585 (N_31585,N_24986,N_29229);
or U31586 (N_31586,N_22296,N_27214);
nor U31587 (N_31587,N_26011,N_24663);
nor U31588 (N_31588,N_21034,N_21519);
xnor U31589 (N_31589,N_23797,N_23160);
nand U31590 (N_31590,N_26250,N_27831);
xnor U31591 (N_31591,N_22540,N_28412);
nand U31592 (N_31592,N_26734,N_22577);
nand U31593 (N_31593,N_24737,N_21129);
nor U31594 (N_31594,N_23006,N_29901);
xor U31595 (N_31595,N_26972,N_23679);
xnor U31596 (N_31596,N_20129,N_21568);
nor U31597 (N_31597,N_24060,N_29544);
and U31598 (N_31598,N_24489,N_25205);
xnor U31599 (N_31599,N_20997,N_24977);
and U31600 (N_31600,N_20204,N_21955);
and U31601 (N_31601,N_23338,N_26121);
xor U31602 (N_31602,N_23019,N_24715);
or U31603 (N_31603,N_28528,N_24043);
and U31604 (N_31604,N_29502,N_28690);
xor U31605 (N_31605,N_26689,N_29650);
nor U31606 (N_31606,N_20557,N_28550);
nor U31607 (N_31607,N_26215,N_24420);
xor U31608 (N_31608,N_28530,N_25004);
xor U31609 (N_31609,N_23075,N_24309);
xor U31610 (N_31610,N_25293,N_23127);
nand U31611 (N_31611,N_28325,N_20423);
nor U31612 (N_31612,N_22525,N_23543);
nand U31613 (N_31613,N_29937,N_29322);
and U31614 (N_31614,N_21146,N_21747);
nand U31615 (N_31615,N_23344,N_29705);
or U31616 (N_31616,N_28288,N_24741);
xnor U31617 (N_31617,N_20190,N_21931);
or U31618 (N_31618,N_21318,N_28281);
nand U31619 (N_31619,N_27114,N_23498);
nor U31620 (N_31620,N_29208,N_26939);
nor U31621 (N_31621,N_22488,N_28399);
or U31622 (N_31622,N_24311,N_23028);
nor U31623 (N_31623,N_27676,N_27423);
nand U31624 (N_31624,N_21184,N_20774);
or U31625 (N_31625,N_25291,N_23866);
nand U31626 (N_31626,N_25169,N_27949);
or U31627 (N_31627,N_28754,N_24657);
or U31628 (N_31628,N_26153,N_26610);
nor U31629 (N_31629,N_26359,N_26216);
nor U31630 (N_31630,N_25729,N_24813);
nor U31631 (N_31631,N_22421,N_22306);
nand U31632 (N_31632,N_26965,N_25906);
and U31633 (N_31633,N_23009,N_24601);
nand U31634 (N_31634,N_21345,N_20394);
nor U31635 (N_31635,N_28029,N_21255);
nand U31636 (N_31636,N_26751,N_29822);
nand U31637 (N_31637,N_22496,N_25499);
xnor U31638 (N_31638,N_29911,N_20155);
nor U31639 (N_31639,N_20261,N_26703);
xor U31640 (N_31640,N_25644,N_27252);
or U31641 (N_31641,N_27796,N_24523);
and U31642 (N_31642,N_26826,N_27189);
xor U31643 (N_31643,N_22967,N_20062);
and U31644 (N_31644,N_29232,N_26954);
and U31645 (N_31645,N_21834,N_25027);
xnor U31646 (N_31646,N_22917,N_23664);
nor U31647 (N_31647,N_25749,N_25685);
nand U31648 (N_31648,N_23832,N_28891);
xnor U31649 (N_31649,N_24559,N_25408);
and U31650 (N_31650,N_28672,N_26796);
nor U31651 (N_31651,N_24974,N_29220);
or U31652 (N_31652,N_23583,N_27448);
nand U31653 (N_31653,N_21307,N_20408);
or U31654 (N_31654,N_22317,N_28564);
or U31655 (N_31655,N_29084,N_20778);
xnor U31656 (N_31656,N_28055,N_28467);
and U31657 (N_31657,N_26793,N_23096);
and U31658 (N_31658,N_21449,N_27058);
or U31659 (N_31659,N_29240,N_27788);
nand U31660 (N_31660,N_23742,N_25343);
xnor U31661 (N_31661,N_28964,N_24147);
or U31662 (N_31662,N_28495,N_25750);
nor U31663 (N_31663,N_22132,N_22675);
nor U31664 (N_31664,N_26673,N_29015);
or U31665 (N_31665,N_27442,N_25629);
nor U31666 (N_31666,N_26040,N_26048);
or U31667 (N_31667,N_25982,N_26127);
and U31668 (N_31668,N_28711,N_22659);
nor U31669 (N_31669,N_21892,N_26892);
nand U31670 (N_31670,N_21750,N_27511);
nor U31671 (N_31671,N_28772,N_23395);
xor U31672 (N_31672,N_23830,N_20389);
nor U31673 (N_31673,N_21119,N_26721);
or U31674 (N_31674,N_21031,N_26884);
or U31675 (N_31675,N_21050,N_23484);
or U31676 (N_31676,N_23561,N_20158);
and U31677 (N_31677,N_26330,N_28073);
nand U31678 (N_31678,N_26520,N_20017);
nor U31679 (N_31679,N_20336,N_23880);
nand U31680 (N_31680,N_23913,N_25436);
and U31681 (N_31681,N_22584,N_25885);
or U31682 (N_31682,N_20859,N_23560);
and U31683 (N_31683,N_22318,N_26424);
nand U31684 (N_31684,N_28043,N_24959);
or U31685 (N_31685,N_22728,N_20792);
nor U31686 (N_31686,N_24914,N_25344);
nand U31687 (N_31687,N_20704,N_27627);
and U31688 (N_31688,N_20614,N_21233);
or U31689 (N_31689,N_25224,N_27225);
nor U31690 (N_31690,N_25946,N_20205);
or U31691 (N_31691,N_24544,N_23300);
nand U31692 (N_31692,N_29739,N_20473);
nand U31693 (N_31693,N_29744,N_25239);
xnor U31694 (N_31694,N_20177,N_25428);
nand U31695 (N_31695,N_28641,N_26850);
nor U31696 (N_31696,N_23061,N_24247);
nand U31697 (N_31697,N_29764,N_26309);
and U31698 (N_31698,N_25901,N_28012);
and U31699 (N_31699,N_24318,N_22431);
nor U31700 (N_31700,N_25331,N_23353);
and U31701 (N_31701,N_27010,N_25616);
and U31702 (N_31702,N_24870,N_24310);
xor U31703 (N_31703,N_23942,N_29174);
nor U31704 (N_31704,N_22224,N_22261);
xor U31705 (N_31705,N_28590,N_29925);
and U31706 (N_31706,N_22750,N_28359);
nand U31707 (N_31707,N_26570,N_24796);
nand U31708 (N_31708,N_29736,N_27343);
nand U31709 (N_31709,N_26889,N_29131);
and U31710 (N_31710,N_28453,N_24824);
nand U31711 (N_31711,N_26701,N_25485);
or U31712 (N_31712,N_26624,N_23607);
xnor U31713 (N_31713,N_21595,N_29963);
xor U31714 (N_31714,N_23993,N_23622);
or U31715 (N_31715,N_26554,N_23782);
xnor U31716 (N_31716,N_23227,N_28556);
and U31717 (N_31717,N_28168,N_29007);
nor U31718 (N_31718,N_22597,N_28324);
nand U31719 (N_31719,N_24517,N_23164);
nand U31720 (N_31720,N_23231,N_26453);
and U31721 (N_31721,N_23477,N_22783);
or U31722 (N_31722,N_26355,N_25266);
nand U31723 (N_31723,N_25702,N_29781);
xor U31724 (N_31724,N_22953,N_29372);
nor U31725 (N_31725,N_27480,N_25243);
or U31726 (N_31726,N_22196,N_23291);
nor U31727 (N_31727,N_28067,N_28127);
xnor U31728 (N_31728,N_22605,N_20657);
nand U31729 (N_31729,N_29577,N_22286);
xor U31730 (N_31730,N_24480,N_22570);
nor U31731 (N_31731,N_25558,N_29648);
nand U31732 (N_31732,N_28162,N_20307);
nand U31733 (N_31733,N_21703,N_21085);
and U31734 (N_31734,N_27641,N_20360);
or U31735 (N_31735,N_26760,N_26399);
and U31736 (N_31736,N_22177,N_26997);
nand U31737 (N_31737,N_26567,N_23114);
nor U31738 (N_31738,N_23368,N_28567);
and U31739 (N_31739,N_27166,N_21926);
or U31740 (N_31740,N_24312,N_27767);
and U31741 (N_31741,N_28014,N_26007);
nand U31742 (N_31742,N_29325,N_21057);
nand U31743 (N_31743,N_21495,N_24146);
or U31744 (N_31744,N_29214,N_24401);
nand U31745 (N_31745,N_28128,N_25466);
nor U31746 (N_31746,N_20973,N_22849);
xor U31747 (N_31747,N_21754,N_26005);
and U31748 (N_31748,N_28257,N_23610);
and U31749 (N_31749,N_28329,N_27832);
and U31750 (N_31750,N_21413,N_27651);
nand U31751 (N_31751,N_22959,N_26812);
or U31752 (N_31752,N_26854,N_27096);
xnor U31753 (N_31753,N_23948,N_28697);
xor U31754 (N_31754,N_29135,N_20722);
nor U31755 (N_31755,N_27164,N_26186);
xnor U31756 (N_31756,N_23513,N_22230);
nand U31757 (N_31757,N_24279,N_20346);
nand U31758 (N_31758,N_27628,N_28337);
nand U31759 (N_31759,N_26702,N_27319);
or U31760 (N_31760,N_21162,N_25859);
nor U31761 (N_31761,N_21204,N_21192);
xor U31762 (N_31762,N_26400,N_28034);
nor U31763 (N_31763,N_25809,N_22589);
xnor U31764 (N_31764,N_29866,N_23903);
or U31765 (N_31765,N_22338,N_20411);
xor U31766 (N_31766,N_26254,N_28177);
nor U31767 (N_31767,N_22499,N_26354);
or U31768 (N_31768,N_28838,N_27734);
xor U31769 (N_31769,N_24992,N_25125);
nand U31770 (N_31770,N_23792,N_25797);
or U31771 (N_31771,N_20438,N_27990);
xnor U31772 (N_31772,N_26334,N_20384);
nor U31773 (N_31773,N_25024,N_22381);
nand U31774 (N_31774,N_27659,N_23408);
nand U31775 (N_31775,N_26553,N_21118);
nor U31776 (N_31776,N_28582,N_25492);
nand U31777 (N_31777,N_23259,N_22531);
nand U31778 (N_31778,N_25948,N_28041);
xor U31779 (N_31779,N_22692,N_20546);
xor U31780 (N_31780,N_29438,N_22980);
xor U31781 (N_31781,N_25172,N_22863);
or U31782 (N_31782,N_20480,N_25721);
nand U31783 (N_31783,N_21960,N_24560);
nand U31784 (N_31784,N_29830,N_27913);
and U31785 (N_31785,N_23232,N_22697);
or U31786 (N_31786,N_27253,N_28484);
or U31787 (N_31787,N_24878,N_20587);
and U31788 (N_31788,N_21331,N_27672);
xnor U31789 (N_31789,N_22516,N_23736);
xnor U31790 (N_31790,N_20968,N_24397);
or U31791 (N_31791,N_28572,N_25334);
xor U31792 (N_31792,N_22928,N_29748);
and U31793 (N_31793,N_29707,N_21405);
and U31794 (N_31794,N_20667,N_26353);
or U31795 (N_31795,N_24303,N_20152);
nand U31796 (N_31796,N_24777,N_28943);
nor U31797 (N_31797,N_24223,N_20079);
nor U31798 (N_31798,N_20270,N_27384);
or U31799 (N_31799,N_26131,N_22816);
or U31800 (N_31800,N_20910,N_22587);
or U31801 (N_31801,N_27933,N_22663);
and U31802 (N_31802,N_22342,N_27654);
or U31803 (N_31803,N_24048,N_23076);
or U31804 (N_31804,N_22222,N_25730);
nor U31805 (N_31805,N_25462,N_27946);
xor U31806 (N_31806,N_23020,N_28827);
nor U31807 (N_31807,N_27293,N_22326);
and U31808 (N_31808,N_24800,N_26383);
nand U31809 (N_31809,N_20041,N_20315);
nand U31810 (N_31810,N_28661,N_24586);
xor U31811 (N_31811,N_24545,N_20303);
or U31812 (N_31812,N_20404,N_27420);
and U31813 (N_31813,N_26950,N_29953);
nand U31814 (N_31814,N_29960,N_29057);
nor U31815 (N_31815,N_23891,N_24872);
nor U31816 (N_31816,N_23388,N_29674);
nor U31817 (N_31817,N_28266,N_29576);
nand U31818 (N_31818,N_23289,N_24195);
xnor U31819 (N_31819,N_26663,N_24206);
or U31820 (N_31820,N_24722,N_22423);
nor U31821 (N_31821,N_28237,N_25074);
nand U31822 (N_31822,N_29460,N_23864);
nand U31823 (N_31823,N_20207,N_20265);
or U31824 (N_31824,N_25221,N_29104);
and U31825 (N_31825,N_22608,N_22249);
nor U31826 (N_31826,N_22468,N_23562);
nor U31827 (N_31827,N_21139,N_28904);
nor U31828 (N_31828,N_20636,N_21264);
xor U31829 (N_31829,N_25824,N_27155);
xor U31830 (N_31830,N_27938,N_26137);
and U31831 (N_31831,N_22283,N_21043);
xor U31832 (N_31832,N_21811,N_24537);
nand U31833 (N_31833,N_22292,N_25770);
or U31834 (N_31834,N_26467,N_29076);
nand U31835 (N_31835,N_25192,N_24250);
nand U31836 (N_31836,N_27879,N_22299);
or U31837 (N_31837,N_26259,N_22776);
xnor U31838 (N_31838,N_24695,N_27598);
or U31839 (N_31839,N_24566,N_27795);
nor U31840 (N_31840,N_26253,N_27939);
or U31841 (N_31841,N_26249,N_22860);
or U31842 (N_31842,N_23297,N_20011);
and U31843 (N_31843,N_22418,N_20529);
nand U31844 (N_31844,N_29642,N_24666);
or U31845 (N_31845,N_21576,N_27645);
nor U31846 (N_31846,N_24641,N_21814);
and U31847 (N_31847,N_27381,N_22981);
nand U31848 (N_31848,N_22735,N_29028);
nor U31849 (N_31849,N_23872,N_24205);
xor U31850 (N_31850,N_20469,N_26781);
xnor U31851 (N_31851,N_22679,N_24954);
or U31852 (N_31852,N_27784,N_26757);
xor U31853 (N_31853,N_22628,N_24866);
and U31854 (N_31854,N_27805,N_29966);
xor U31855 (N_31855,N_24909,N_24793);
or U31856 (N_31856,N_21457,N_29586);
or U31857 (N_31857,N_23839,N_21363);
xor U31858 (N_31858,N_21514,N_23655);
or U31859 (N_31859,N_21803,N_23909);
nand U31860 (N_31860,N_22114,N_26438);
nor U31861 (N_31861,N_26927,N_28493);
nand U31862 (N_31862,N_22512,N_23756);
and U31863 (N_31863,N_28616,N_28056);
nand U31864 (N_31864,N_21599,N_29189);
nor U31865 (N_31865,N_26295,N_21220);
or U31866 (N_31866,N_26513,N_24864);
xor U31867 (N_31867,N_20713,N_22156);
nand U31868 (N_31868,N_28229,N_21601);
or U31869 (N_31869,N_29792,N_23384);
or U31870 (N_31870,N_24818,N_29959);
xor U31871 (N_31871,N_28926,N_22459);
nor U31872 (N_31872,N_29842,N_23549);
nand U31873 (N_31873,N_28951,N_24622);
and U31874 (N_31874,N_22817,N_26583);
xor U31875 (N_31875,N_25555,N_24915);
or U31876 (N_31876,N_21552,N_24433);
or U31877 (N_31877,N_22854,N_21355);
nor U31878 (N_31878,N_26580,N_24924);
or U31879 (N_31879,N_28900,N_21642);
and U31880 (N_31880,N_25327,N_25353);
or U31881 (N_31881,N_22724,N_28928);
nor U31882 (N_31882,N_26209,N_28818);
and U31883 (N_31883,N_24065,N_21885);
nand U31884 (N_31884,N_25480,N_22071);
xor U31885 (N_31885,N_22394,N_29013);
nand U31886 (N_31886,N_28732,N_20984);
nor U31887 (N_31887,N_23997,N_26786);
and U31888 (N_31888,N_20039,N_20110);
or U31889 (N_31889,N_25572,N_22031);
nor U31890 (N_31890,N_20377,N_27986);
and U31891 (N_31891,N_22133,N_28705);
or U31892 (N_31892,N_25798,N_22321);
nand U31893 (N_31893,N_23123,N_28985);
or U31894 (N_31894,N_26073,N_22822);
or U31895 (N_31895,N_25069,N_27657);
nor U31896 (N_31896,N_22847,N_29034);
or U31897 (N_31897,N_29825,N_24151);
and U31898 (N_31898,N_21463,N_24600);
xor U31899 (N_31899,N_21188,N_29590);
nor U31900 (N_31900,N_20924,N_28545);
and U31901 (N_31901,N_25498,N_28678);
nand U31902 (N_31902,N_21761,N_26093);
and U31903 (N_31903,N_29474,N_26489);
nand U31904 (N_31904,N_23072,N_28569);
and U31905 (N_31905,N_24656,N_26794);
and U31906 (N_31906,N_24418,N_29080);
nand U31907 (N_31907,N_28814,N_20269);
or U31908 (N_31908,N_24458,N_21369);
and U31909 (N_31909,N_24403,N_21954);
and U31910 (N_31910,N_25418,N_26076);
and U31911 (N_31911,N_23284,N_22566);
nand U31912 (N_31912,N_29114,N_26831);
and U31913 (N_31913,N_20381,N_23363);
xor U31914 (N_31914,N_26533,N_22517);
and U31915 (N_31915,N_28816,N_26966);
nor U31916 (N_31916,N_20505,N_26556);
or U31917 (N_31917,N_21177,N_21933);
and U31918 (N_31918,N_22726,N_20425);
or U31919 (N_31919,N_22601,N_22099);
nor U31920 (N_31920,N_24288,N_21997);
nor U31921 (N_31921,N_23391,N_21106);
xor U31922 (N_31922,N_28899,N_21406);
or U31923 (N_31923,N_23676,N_22734);
and U31924 (N_31924,N_21044,N_21252);
nor U31925 (N_31925,N_29743,N_27758);
nor U31926 (N_31926,N_24585,N_29054);
nand U31927 (N_31927,N_26566,N_21452);
xor U31928 (N_31928,N_23956,N_26147);
nor U31929 (N_31929,N_29127,N_28270);
and U31930 (N_31930,N_29147,N_21600);
and U31931 (N_31931,N_23392,N_23926);
and U31932 (N_31932,N_29329,N_29081);
xor U31933 (N_31933,N_23173,N_28019);
and U31934 (N_31934,N_21074,N_22909);
nor U31935 (N_31935,N_26111,N_21899);
nand U31936 (N_31936,N_25118,N_26956);
or U31937 (N_31937,N_25713,N_23456);
or U31938 (N_31938,N_29314,N_29143);
nor U31939 (N_31939,N_24594,N_27711);
and U31940 (N_31940,N_28911,N_29316);
or U31941 (N_31941,N_27917,N_27043);
nand U31942 (N_31942,N_24754,N_26061);
xnor U31943 (N_31943,N_23572,N_26277);
and U31944 (N_31944,N_26167,N_24506);
xnor U31945 (N_31945,N_23739,N_24969);
nand U31946 (N_31946,N_20310,N_24614);
nand U31947 (N_31947,N_26434,N_23811);
nand U31948 (N_31948,N_28652,N_23253);
xor U31949 (N_31949,N_29161,N_20987);
nor U31950 (N_31950,N_26620,N_28136);
xor U31951 (N_31951,N_23215,N_21451);
xor U31952 (N_31952,N_24746,N_21839);
and U31953 (N_31953,N_22835,N_21725);
and U31954 (N_31954,N_28203,N_20484);
nor U31955 (N_31955,N_25160,N_24760);
nor U31956 (N_31956,N_27971,N_21614);
and U31957 (N_31957,N_23794,N_22751);
xor U31958 (N_31958,N_20383,N_25731);
nor U31959 (N_31959,N_20215,N_20454);
nor U31960 (N_31960,N_23239,N_20975);
xnor U31961 (N_31961,N_21222,N_22742);
or U31962 (N_31962,N_22109,N_28845);
or U31963 (N_31963,N_24369,N_26206);
and U31964 (N_31964,N_20009,N_25687);
or U31965 (N_31965,N_29298,N_27677);
nand U31966 (N_31966,N_22409,N_24521);
xor U31967 (N_31967,N_21080,N_20559);
xor U31968 (N_31968,N_25246,N_22319);
xor U31969 (N_31969,N_28511,N_24903);
and U31970 (N_31970,N_26584,N_27882);
nand U31971 (N_31971,N_22059,N_23808);
xor U31972 (N_31972,N_27036,N_29236);
and U31973 (N_31973,N_21596,N_27610);
or U31974 (N_31974,N_23898,N_29693);
nand U31975 (N_31975,N_22685,N_26943);
and U31976 (N_31976,N_27750,N_28113);
and U31977 (N_31977,N_29639,N_28475);
xor U31978 (N_31978,N_22086,N_20070);
and U31979 (N_31979,N_27125,N_29812);
xor U31980 (N_31980,N_26859,N_22289);
or U31981 (N_31981,N_25957,N_29643);
xnor U31982 (N_31982,N_21025,N_25936);
xor U31983 (N_31983,N_25447,N_21036);
and U31984 (N_31984,N_27502,N_21782);
nor U31985 (N_31985,N_26829,N_27222);
xnor U31986 (N_31986,N_27105,N_21262);
nand U31987 (N_31987,N_25038,N_20043);
nand U31988 (N_31988,N_24540,N_28654);
xnor U31989 (N_31989,N_26172,N_25272);
xor U31990 (N_31990,N_20781,N_20500);
nand U31991 (N_31991,N_26021,N_23279);
nor U31992 (N_31992,N_26926,N_21970);
nand U31993 (N_31993,N_20746,N_25467);
and U31994 (N_31994,N_26716,N_29444);
xor U31995 (N_31995,N_20407,N_22162);
nor U31996 (N_31996,N_28959,N_26387);
and U31997 (N_31997,N_29226,N_27183);
nand U31998 (N_31998,N_21243,N_23335);
nand U31999 (N_31999,N_27877,N_28295);
and U32000 (N_32000,N_23821,N_20478);
nand U32001 (N_32001,N_23302,N_29137);
nor U32002 (N_32002,N_25930,N_29695);
or U32003 (N_32003,N_22729,N_29789);
xnor U32004 (N_32004,N_21360,N_23458);
xor U32005 (N_32005,N_29484,N_21760);
nor U32006 (N_32006,N_22694,N_24787);
nor U32007 (N_32007,N_26617,N_20890);
nor U32008 (N_32008,N_21748,N_25399);
or U32009 (N_32009,N_21999,N_22083);
nor U32010 (N_32010,N_23967,N_24932);
nand U32011 (N_32011,N_24485,N_27100);
nand U32012 (N_32012,N_22291,N_29522);
xnor U32013 (N_32013,N_25147,N_21684);
xnor U32014 (N_32014,N_27136,N_24197);
or U32015 (N_32015,N_24558,N_27024);
xor U32016 (N_32016,N_23773,N_23861);
and U32017 (N_32017,N_28293,N_26120);
nor U32018 (N_32018,N_26962,N_25893);
nand U32019 (N_32019,N_23964,N_26929);
or U32020 (N_32020,N_29973,N_21260);
or U32021 (N_32021,N_22777,N_21742);
and U32022 (N_32022,N_26710,N_27931);
xnor U32023 (N_32023,N_23455,N_20357);
xor U32024 (N_32024,N_22020,N_22490);
nor U32025 (N_32025,N_27714,N_25091);
xor U32026 (N_32026,N_24993,N_23486);
nand U32027 (N_32027,N_20229,N_24389);
xor U32028 (N_32028,N_27037,N_22798);
and U32029 (N_32029,N_29318,N_22366);
nand U32030 (N_32030,N_27255,N_21422);
or U32031 (N_32031,N_27383,N_28968);
nand U32032 (N_32032,N_23167,N_29621);
or U32033 (N_32033,N_29102,N_20616);
nor U32034 (N_32034,N_23220,N_24450);
xor U32035 (N_32035,N_24461,N_23094);
or U32036 (N_32036,N_27846,N_21821);
or U32037 (N_32037,N_22851,N_26791);
nor U32038 (N_32038,N_20276,N_25958);
or U32039 (N_32039,N_20151,N_23890);
nand U32040 (N_32040,N_28444,N_28723);
or U32041 (N_32041,N_24356,N_22805);
nor U32042 (N_32042,N_29230,N_20262);
nand U32043 (N_32043,N_20699,N_23766);
xnor U32044 (N_32044,N_20716,N_29618);
nand U32045 (N_32045,N_20625,N_24390);
xnor U32046 (N_32046,N_28870,N_23404);
xor U32047 (N_32047,N_20624,N_20337);
and U32048 (N_32048,N_26514,N_23823);
nor U32049 (N_32049,N_29675,N_23041);
xnor U32050 (N_32050,N_22246,N_23925);
xor U32051 (N_32051,N_22433,N_26404);
and U32052 (N_32052,N_23932,N_26637);
or U32053 (N_32053,N_22537,N_26420);
xnor U32054 (N_32054,N_24114,N_28403);
nor U32055 (N_32055,N_28308,N_28776);
nand U32056 (N_32056,N_26798,N_27331);
nand U32057 (N_32057,N_25215,N_20083);
nor U32058 (N_32058,N_24898,N_24942);
xnor U32059 (N_32059,N_28260,N_28945);
xor U32060 (N_32060,N_27238,N_28074);
or U32061 (N_32061,N_25416,N_27050);
or U32062 (N_32062,N_20617,N_20217);
xnor U32063 (N_32063,N_26682,N_23100);
nor U32064 (N_32064,N_29008,N_21312);
and U32065 (N_32065,N_23207,N_23730);
or U32066 (N_32066,N_26029,N_28865);
and U32067 (N_32067,N_23229,N_26465);
and U32068 (N_32068,N_22768,N_26820);
and U32069 (N_32069,N_28375,N_24361);
and U32070 (N_32070,N_24028,N_28912);
nand U32071 (N_32071,N_26345,N_26464);
nand U32072 (N_32072,N_23540,N_27817);
and U32073 (N_32073,N_26836,N_24117);
xnor U32074 (N_32074,N_29654,N_28929);
xnor U32075 (N_32075,N_21692,N_22038);
xnor U32076 (N_32076,N_22278,N_21175);
or U32077 (N_32077,N_26960,N_27389);
nor U32078 (N_32078,N_22739,N_26281);
and U32079 (N_32079,N_28286,N_25076);
and U32080 (N_32080,N_26026,N_22668);
and U32081 (N_32081,N_23847,N_29280);
and U32082 (N_32082,N_21530,N_22630);
or U32083 (N_32083,N_27057,N_22626);
or U32084 (N_32084,N_25489,N_25844);
or U32085 (N_32085,N_24023,N_29451);
nand U32086 (N_32086,N_21637,N_20533);
and U32087 (N_32087,N_23152,N_29863);
and U32088 (N_32088,N_28378,N_28368);
nand U32089 (N_32089,N_24373,N_21894);
nand U32090 (N_32090,N_27943,N_29459);
nand U32091 (N_32091,N_25882,N_20540);
xor U32092 (N_32092,N_23137,N_27041);
xnor U32093 (N_32093,N_26573,N_28832);
nor U32094 (N_32094,N_24815,N_20998);
or U32095 (N_32095,N_26891,N_28338);
nand U32096 (N_32096,N_24088,N_26784);
nor U32097 (N_32097,N_20931,N_29869);
and U32098 (N_32098,N_25840,N_28817);
and U32099 (N_32099,N_24723,N_20266);
nand U32100 (N_32100,N_22954,N_20162);
nand U32101 (N_32101,N_26090,N_27346);
nand U32102 (N_32102,N_26983,N_21001);
nand U32103 (N_32103,N_29416,N_23662);
nand U32104 (N_32104,N_21838,N_24096);
xor U32105 (N_32105,N_25039,N_28290);
nand U32106 (N_32106,N_20645,N_24414);
xor U32107 (N_32107,N_28405,N_22524);
and U32108 (N_32108,N_22580,N_25928);
nand U32109 (N_32109,N_21731,N_28841);
nand U32110 (N_32110,N_28847,N_21273);
nand U32111 (N_32111,N_23292,N_24108);
and U32112 (N_32112,N_29527,N_21124);
nand U32113 (N_32113,N_25827,N_23495);
nor U32114 (N_32114,N_24664,N_20281);
and U32115 (N_32115,N_27729,N_20213);
and U32116 (N_32116,N_22635,N_21211);
and U32117 (N_32117,N_23704,N_23133);
or U32118 (N_32118,N_20416,N_20527);
nor U32119 (N_32119,N_22719,N_22779);
or U32120 (N_32120,N_27047,N_22004);
or U32121 (N_32121,N_24286,N_25015);
or U32122 (N_32122,N_29815,N_29553);
xor U32123 (N_32123,N_27398,N_21905);
nor U32124 (N_32124,N_25319,N_27546);
nor U32125 (N_32125,N_26896,N_27821);
and U32126 (N_32126,N_27338,N_27573);
and U32127 (N_32127,N_21073,N_27552);
and U32128 (N_32128,N_21633,N_26099);
xor U32129 (N_32129,N_21738,N_20220);
and U32130 (N_32130,N_24562,N_20403);
nand U32131 (N_32131,N_20782,N_27579);
xnor U32132 (N_32132,N_28402,N_24249);
nor U32133 (N_32133,N_23566,N_23179);
nand U32134 (N_32134,N_21326,N_28356);
nand U32135 (N_32135,N_21460,N_27168);
or U32136 (N_32136,N_24122,N_26968);
xor U32137 (N_32137,N_21798,N_28811);
and U32138 (N_32138,N_21769,N_25158);
and U32139 (N_32139,N_21083,N_25675);
and U32140 (N_32140,N_23772,N_23835);
xnor U32141 (N_32141,N_23529,N_23062);
and U32142 (N_32142,N_21625,N_29511);
nor U32143 (N_32143,N_21266,N_25386);
and U32144 (N_32144,N_26985,N_22621);
xnor U32145 (N_32145,N_24734,N_26909);
or U32146 (N_32146,N_24809,N_21185);
nor U32147 (N_32147,N_24378,N_20641);
xnor U32148 (N_32148,N_23349,N_25716);
or U32149 (N_32149,N_27847,N_29627);
xor U32150 (N_32150,N_24242,N_21120);
xor U32151 (N_32151,N_20388,N_26074);
or U32152 (N_32152,N_24009,N_20273);
xnor U32153 (N_32153,N_24745,N_29248);
and U32154 (N_32154,N_28057,N_22387);
and U32155 (N_32155,N_28502,N_28687);
and U32156 (N_32156,N_27731,N_28613);
xnor U32157 (N_32157,N_27137,N_27576);
and U32158 (N_32158,N_29846,N_25728);
nand U32159 (N_32159,N_24285,N_28531);
and U32160 (N_32160,N_21995,N_21520);
or U32161 (N_32161,N_27025,N_25753);
nand U32162 (N_32162,N_21880,N_27937);
and U32163 (N_32163,N_23277,N_20051);
nor U32164 (N_32164,N_25300,N_21012);
and U32165 (N_32165,N_29401,N_21812);
nor U32166 (N_32166,N_25520,N_25920);
xor U32167 (N_32167,N_27162,N_28152);
nor U32168 (N_32168,N_26226,N_23602);
nor U32169 (N_32169,N_23894,N_23093);
nand U32170 (N_32170,N_27271,N_29249);
nor U32171 (N_32171,N_22715,N_23170);
nor U32172 (N_32172,N_29694,N_29350);
and U32173 (N_32173,N_21020,N_29491);
and U32174 (N_32174,N_21668,N_21135);
nor U32175 (N_32175,N_24300,N_24287);
or U32176 (N_32176,N_27490,N_28789);
nand U32177 (N_32177,N_22380,N_23088);
or U32178 (N_32178,N_20115,N_27466);
and U32179 (N_32179,N_28137,N_27650);
nor U32180 (N_32180,N_24739,N_22707);
and U32181 (N_32181,N_22897,N_23991);
nand U32182 (N_32182,N_27867,N_28252);
nor U32183 (N_32183,N_28143,N_24409);
nor U32184 (N_32184,N_20431,N_21052);
nand U32185 (N_32185,N_26210,N_20677);
and U32186 (N_32186,N_28763,N_24961);
and U32187 (N_32187,N_24026,N_23447);
nand U32188 (N_32188,N_27487,N_25231);
nand U32189 (N_32189,N_23105,N_21667);
nand U32190 (N_32190,N_23638,N_22711);
nand U32191 (N_32191,N_23548,N_27202);
or U32192 (N_32192,N_21679,N_26558);
nor U32193 (N_32193,N_22906,N_26519);
or U32194 (N_32194,N_25350,N_26509);
nand U32195 (N_32195,N_20495,N_28384);
xor U32196 (N_32196,N_29849,N_21070);
nand U32197 (N_32197,N_23836,N_26102);
and U32198 (N_32198,N_23270,N_23998);
or U32199 (N_32199,N_23417,N_25137);
or U32200 (N_32200,N_20757,N_28159);
nand U32201 (N_32201,N_22744,N_22464);
nor U32202 (N_32202,N_29991,N_27660);
nor U32203 (N_32203,N_27228,N_26018);
and U32204 (N_32204,N_28254,N_29058);
or U32205 (N_32205,N_28881,N_23082);
and U32206 (N_32206,N_21281,N_22877);
and U32207 (N_32207,N_28692,N_21547);
xnor U32208 (N_32208,N_29424,N_25554);
and U32209 (N_32209,N_21285,N_29551);
nor U32210 (N_32210,N_23509,N_25511);
and U32211 (N_32211,N_26625,N_23652);
nor U32212 (N_32212,N_26940,N_21502);
nand U32213 (N_32213,N_27722,N_23333);
or U32214 (N_32214,N_29896,N_23375);
nand U32215 (N_32215,N_27129,N_26452);
xnor U32216 (N_32216,N_20901,N_23799);
nand U32217 (N_32217,N_26971,N_21130);
and U32218 (N_32218,N_20508,N_23440);
xor U32219 (N_32219,N_24794,N_27740);
xor U32220 (N_32220,N_27849,N_21054);
nand U32221 (N_32221,N_24381,N_25934);
nor U32222 (N_32222,N_23978,N_27819);
nor U32223 (N_32223,N_22274,N_24635);
xnor U32224 (N_32224,N_22379,N_23959);
nand U32225 (N_32225,N_29219,N_25681);
xor U32226 (N_32226,N_28583,N_26190);
nor U32227 (N_32227,N_24324,N_24282);
nand U32228 (N_32228,N_25932,N_22415);
xor U32229 (N_32229,N_29604,N_24701);
nor U32230 (N_32230,N_23226,N_25455);
or U32231 (N_32231,N_20905,N_21067);
xnor U32232 (N_32232,N_27955,N_28836);
xor U32233 (N_32233,N_25124,N_21720);
nor U32234 (N_32234,N_24339,N_22958);
nand U32235 (N_32235,N_29756,N_25777);
or U32236 (N_32236,N_24315,N_28570);
nor U32237 (N_32237,N_27701,N_22771);
or U32238 (N_32238,N_23110,N_21677);
xnor U32239 (N_32239,N_29446,N_29681);
or U32240 (N_32240,N_29780,N_21283);
or U32241 (N_32241,N_24494,N_27690);
or U32242 (N_32242,N_27157,N_21923);
or U32243 (N_32243,N_27272,N_29069);
or U32244 (N_32244,N_29203,N_26759);
or U32245 (N_32245,N_21545,N_27721);
and U32246 (N_32246,N_29178,N_29518);
and U32247 (N_32247,N_29012,N_20280);
xnor U32248 (N_32248,N_26719,N_24553);
or U32249 (N_32249,N_26152,N_24101);
or U32250 (N_32250,N_23628,N_28597);
nor U32251 (N_32251,N_20969,N_25504);
and U32252 (N_32252,N_25143,N_22506);
and U32253 (N_32253,N_28611,N_25986);
nor U32254 (N_32254,N_22356,N_29851);
xnor U32255 (N_32255,N_27492,N_23235);
xor U32256 (N_32256,N_24688,N_20974);
nor U32257 (N_32257,N_28089,N_23984);
and U32258 (N_32258,N_27461,N_25127);
or U32259 (N_32259,N_21059,N_27945);
and U32260 (N_32260,N_21548,N_29144);
nor U32261 (N_32261,N_26202,N_21563);
xnor U32262 (N_32262,N_25359,N_27299);
nand U32263 (N_32263,N_27281,N_23144);
nor U32264 (N_32264,N_21493,N_27177);
nand U32265 (N_32265,N_24612,N_20374);
xor U32266 (N_32266,N_20099,N_28464);
or U32267 (N_32267,N_20768,N_29355);
nand U32268 (N_32268,N_23002,N_29046);
and U32269 (N_32269,N_24462,N_28366);
nor U32270 (N_32270,N_25133,N_22014);
and U32271 (N_32271,N_28715,N_29861);
xor U32272 (N_32272,N_20693,N_29932);
or U32273 (N_32273,N_29029,N_29547);
and U32274 (N_32274,N_24802,N_29324);
nand U32275 (N_32275,N_28072,N_21412);
nand U32276 (N_32276,N_25733,N_20324);
and U32277 (N_32277,N_27541,N_25186);
or U32278 (N_32278,N_27270,N_20787);
or U32279 (N_32279,N_23327,N_24684);
nand U32280 (N_32280,N_25070,N_29878);
nand U32281 (N_32281,N_20194,N_29908);
nor U32282 (N_32282,N_21889,N_27959);
nor U32283 (N_32283,N_28023,N_21482);
nand U32284 (N_32284,N_29836,N_23138);
nand U32285 (N_32285,N_21183,N_22148);
nor U32286 (N_32286,N_23473,N_22749);
nand U32287 (N_32287,N_20317,N_26234);
xor U32288 (N_32288,N_20634,N_29916);
nor U32289 (N_32289,N_26428,N_24145);
nor U32290 (N_32290,N_29227,N_21276);
xnor U32291 (N_32291,N_25790,N_23272);
or U32292 (N_32292,N_27428,N_28155);
xor U32293 (N_32293,N_26998,N_21309);
nand U32294 (N_32294,N_20668,N_20853);
nor U32295 (N_32295,N_28734,N_25574);
xnor U32296 (N_32296,N_22401,N_28218);
nor U32297 (N_32297,N_21608,N_22355);
xor U32298 (N_32298,N_25703,N_25707);
nor U32299 (N_32299,N_21415,N_29153);
nor U32300 (N_32300,N_25540,N_24547);
and U32301 (N_32301,N_20032,N_23648);
xor U32302 (N_32302,N_24441,N_24925);
xor U32303 (N_32303,N_27431,N_22845);
and U32304 (N_32304,N_29107,N_26182);
nor U32305 (N_32305,N_20671,N_20450);
nor U32306 (N_32306,N_20486,N_25525);
nand U32307 (N_32307,N_28236,N_24881);
xnor U32308 (N_32308,N_27401,N_25375);
nand U32309 (N_32309,N_22687,N_21208);
xor U32310 (N_32310,N_23885,N_28442);
nand U32311 (N_32311,N_24165,N_24907);
or U32312 (N_32312,N_28269,N_21246);
nand U32313 (N_32313,N_22837,N_25903);
or U32314 (N_32314,N_28219,N_21245);
nor U32315 (N_32315,N_27806,N_23010);
or U32316 (N_32316,N_22127,N_25820);
and U32317 (N_32317,N_29691,N_28420);
nand U32318 (N_32318,N_24328,N_25210);
and U32319 (N_32319,N_27854,N_25067);
and U32320 (N_32320,N_28086,N_25897);
nand U32321 (N_32321,N_20459,N_22599);
or U32322 (N_32322,N_25060,N_21014);
xnor U32323 (N_32323,N_29096,N_27736);
xor U32324 (N_32324,N_28506,N_24047);
and U32325 (N_32325,N_23244,N_25878);
nor U32326 (N_32326,N_29768,N_23317);
xor U32327 (N_32327,N_24811,N_25426);
nor U32328 (N_32328,N_25422,N_25989);
and U32329 (N_32329,N_28658,N_21906);
or U32330 (N_32330,N_21560,N_26816);
nor U32331 (N_32331,N_26774,N_25362);
xnor U32332 (N_32332,N_28752,N_28478);
nor U32333 (N_32333,N_26778,N_28336);
xor U32334 (N_32334,N_23189,N_23796);
or U32335 (N_32335,N_27344,N_20669);
nand U32336 (N_32336,N_29613,N_24768);
nor U32337 (N_32337,N_28805,N_21666);
xor U32338 (N_32338,N_24188,N_20406);
or U32339 (N_32339,N_23975,N_22625);
nand U32340 (N_32340,N_26964,N_21454);
xnor U32341 (N_32341,N_25648,N_25253);
and U32342 (N_32342,N_21042,N_26510);
or U32343 (N_32343,N_28780,N_21226);
and U32344 (N_32344,N_22119,N_22138);
xor U32345 (N_32345,N_20589,N_28736);
and U32346 (N_32346,N_24453,N_25208);
xor U32347 (N_32347,N_29657,N_22985);
xnor U32348 (N_32348,N_21771,N_25717);
xor U32349 (N_32349,N_22095,N_22102);
xor U32350 (N_32350,N_23770,N_22636);
or U32351 (N_32351,N_25742,N_27395);
nand U32352 (N_32352,N_24608,N_24120);
nand U32353 (N_32353,N_20558,N_27901);
nor U32354 (N_32354,N_26060,N_27035);
nand U32355 (N_32355,N_29353,N_25752);
nand U32356 (N_32356,N_27277,N_27565);
and U32357 (N_32357,N_25415,N_26564);
xnor U32358 (N_32358,N_26550,N_23690);
or U32359 (N_32359,N_28333,N_21160);
nor U32360 (N_32360,N_26518,N_24642);
or U32361 (N_32361,N_20603,N_28783);
nor U32362 (N_32362,N_20900,N_28284);
xor U32363 (N_32363,N_24015,N_23434);
and U32364 (N_32364,N_26557,N_25543);
nand U32365 (N_32365,N_22483,N_26161);
xor U32366 (N_32366,N_27522,N_22026);
or U32367 (N_32367,N_25720,N_24930);
or U32368 (N_32368,N_26905,N_26064);
xnor U32369 (N_32369,N_23309,N_26445);
xnor U32370 (N_32370,N_23804,N_29172);
or U32371 (N_32371,N_29184,N_29745);
nand U32372 (N_32372,N_25392,N_29317);
and U32373 (N_32373,N_28969,N_26899);
xor U32374 (N_32374,N_21605,N_25532);
or U32375 (N_32375,N_21702,N_21096);
nor U32376 (N_32376,N_29095,N_20069);
nand U32377 (N_32377,N_24843,N_23725);
or U32378 (N_32378,N_27669,N_20228);
xnor U32379 (N_32379,N_29727,N_24887);
nand U32380 (N_32380,N_27112,N_23429);
nor U32381 (N_32381,N_24273,N_25194);
nor U32382 (N_32382,N_27172,N_24217);
or U32383 (N_32383,N_26530,N_24133);
xor U32384 (N_32384,N_23850,N_22764);
nand U32385 (N_32385,N_29193,N_25373);
nor U32386 (N_32386,N_24889,N_25589);
or U32387 (N_32387,N_23585,N_21859);
nand U32388 (N_32388,N_23261,N_24522);
or U32389 (N_32389,N_27828,N_29021);
nor U32390 (N_32390,N_20966,N_26223);
xor U32391 (N_32391,N_22762,N_29061);
nand U32392 (N_32392,N_22961,N_25292);
or U32393 (N_32393,N_21716,N_28262);
and U32394 (N_32394,N_27985,N_29879);
and U32395 (N_32395,N_24266,N_28328);
or U32396 (N_32396,N_24953,N_23442);
nor U32397 (N_32397,N_23876,N_27583);
or U32398 (N_32398,N_27044,N_22219);
xnor U32399 (N_32399,N_27544,N_20815);
nor U32400 (N_32400,N_24317,N_20076);
nand U32401 (N_32401,N_24198,N_29503);
or U32402 (N_32402,N_27085,N_29337);
nor U32403 (N_32403,N_22746,N_21517);
nand U32404 (N_32404,N_25382,N_29251);
xnor U32405 (N_32405,N_27843,N_28863);
or U32406 (N_32406,N_23669,N_25952);
nand U32407 (N_32407,N_28100,N_28631);
xor U32408 (N_32408,N_25042,N_24398);
and U32409 (N_32409,N_22507,N_21104);
or U32410 (N_32410,N_28215,N_28449);
or U32411 (N_32411,N_27133,N_21512);
nand U32412 (N_32412,N_23757,N_22655);
xnor U32413 (N_32413,N_23608,N_27494);
or U32414 (N_32414,N_22632,N_26692);
xnor U32415 (N_32415,N_26329,N_22165);
and U32416 (N_32416,N_27140,N_20825);
or U32417 (N_32417,N_26124,N_20104);
nand U32418 (N_32418,N_24945,N_20477);
and U32419 (N_32419,N_24487,N_25274);
and U32420 (N_32420,N_28856,N_22251);
and U32421 (N_32421,N_24579,N_25743);
nor U32422 (N_32422,N_24090,N_22613);
nand U32423 (N_32423,N_26802,N_28663);
nand U32424 (N_32424,N_24661,N_20790);
nor U32425 (N_32425,N_20680,N_29838);
nand U32426 (N_32426,N_29740,N_26499);
or U32427 (N_32427,N_25398,N_25955);
and U32428 (N_32428,N_22008,N_27324);
nand U32429 (N_32429,N_24473,N_26442);
and U32430 (N_32430,N_27120,N_21395);
xnor U32431 (N_32431,N_28354,N_29090);
and U32432 (N_32432,N_21289,N_24590);
nand U32433 (N_32433,N_20168,N_20596);
nand U32434 (N_32434,N_26834,N_23722);
or U32435 (N_32435,N_25562,N_23156);
and U32436 (N_32436,N_27107,N_22260);
and U32437 (N_32437,N_21724,N_29032);
xnor U32438 (N_32438,N_28640,N_28446);
or U32439 (N_32439,N_24610,N_24922);
or U32440 (N_32440,N_28558,N_26805);
nor U32441 (N_32441,N_22092,N_20359);
nor U32442 (N_32442,N_20748,N_28373);
and U32443 (N_32443,N_20127,N_26088);
or U32444 (N_32444,N_24841,N_25238);
nand U32445 (N_32445,N_20021,N_21153);
xor U32446 (N_32446,N_23204,N_20659);
nor U32447 (N_32447,N_29361,N_20979);
xnor U32448 (N_32448,N_23605,N_24301);
xnor U32449 (N_32449,N_26608,N_25401);
and U32450 (N_32450,N_25472,N_23351);
or U32451 (N_32451,N_22297,N_24451);
or U32452 (N_32452,N_25338,N_29841);
or U32453 (N_32453,N_25308,N_21674);
nand U32454 (N_32454,N_29439,N_26792);
or U32455 (N_32455,N_21912,N_23145);
and U32456 (N_32456,N_20780,N_23515);
xor U32457 (N_32457,N_25474,N_22369);
or U32458 (N_32458,N_29600,N_21138);
nor U32459 (N_32459,N_22568,N_26686);
nor U32460 (N_32460,N_28846,N_20400);
or U32461 (N_32461,N_24726,N_28179);
and U32462 (N_32462,N_20305,N_27884);
or U32463 (N_32463,N_28349,N_24984);
xnor U32464 (N_32464,N_24994,N_28854);
nor U32465 (N_32465,N_28018,N_24504);
nand U32466 (N_32466,N_26181,N_26478);
nor U32467 (N_32467,N_20696,N_23907);
nand U32468 (N_32468,N_27084,N_22938);
nand U32469 (N_32469,N_29758,N_22220);
nand U32470 (N_32470,N_26306,N_26024);
xnor U32471 (N_32471,N_20681,N_24766);
or U32472 (N_32472,N_25206,N_24511);
xor U32473 (N_32473,N_20697,N_22009);
nand U32474 (N_32474,N_25490,N_23008);
xor U32475 (N_32475,N_26177,N_20852);
nor U32476 (N_32476,N_23933,N_29311);
nor U32477 (N_32477,N_27724,N_21949);
nand U32478 (N_32478,N_25064,N_23490);
nand U32479 (N_32479,N_21165,N_21076);
nand U32480 (N_32480,N_26047,N_27367);
and U32481 (N_32481,N_29923,N_28844);
and U32482 (N_32482,N_22161,N_23877);
nand U32483 (N_32483,N_22673,N_22280);
or U32484 (N_32484,N_24091,N_21444);
xnor U32485 (N_32485,N_22743,N_26163);
and U32486 (N_32486,N_23132,N_29477);
nand U32487 (N_32487,N_20633,N_25658);
and U32488 (N_32488,N_29262,N_29589);
and U32489 (N_32489,N_21873,N_29630);
nand U32490 (N_32490,N_26336,N_24278);
or U32491 (N_32491,N_23293,N_23645);
or U32492 (N_32492,N_23046,N_29155);
nand U32493 (N_32493,N_22425,N_29049);
or U32494 (N_32494,N_24875,N_22477);
and U32495 (N_32495,N_27542,N_27811);
nor U32496 (N_32496,N_29117,N_21021);
or U32497 (N_32497,N_29631,N_22466);
nor U32498 (N_32498,N_23049,N_26288);
nand U32499 (N_32499,N_23065,N_22813);
and U32500 (N_32500,N_25631,N_22358);
xor U32501 (N_32501,N_25236,N_23688);
and U32502 (N_32502,N_22720,N_27745);
nor U32503 (N_32503,N_28377,N_24593);
nand U32504 (N_32504,N_28762,N_23936);
or U32505 (N_32505,N_23086,N_24304);
or U32506 (N_32506,N_29835,N_26910);
or U32507 (N_32507,N_25404,N_29599);
nand U32508 (N_32508,N_21235,N_24019);
nand U32509 (N_32509,N_20865,N_24529);
nand U32510 (N_32510,N_22243,N_26937);
xnor U32511 (N_32511,N_23574,N_23889);
or U32512 (N_32512,N_27055,N_26925);
and U32513 (N_32513,N_24842,N_29919);
or U32514 (N_32514,N_23954,N_28386);
xnor U32515 (N_32515,N_24618,N_22974);
xnor U32516 (N_32516,N_29558,N_24867);
nor U32517 (N_32517,N_27754,N_20421);
xnor U32518 (N_32518,N_27304,N_27345);
nand U32519 (N_32519,N_28745,N_20971);
nor U32520 (N_32520,N_28037,N_21088);
or U32521 (N_32521,N_22712,N_27426);
nor U32522 (N_32522,N_28319,N_25528);
or U32523 (N_32523,N_22107,N_27793);
or U32524 (N_32524,N_29708,N_27697);
or U32525 (N_32525,N_25611,N_24834);
xor U32526 (N_32526,N_28212,N_28888);
or U32527 (N_32527,N_22693,N_26500);
or U32528 (N_32528,N_23255,N_28454);
nor U32529 (N_32529,N_21710,N_22200);
xor U32530 (N_32530,N_23210,N_27273);
nor U32531 (N_32531,N_26372,N_29853);
nand U32532 (N_32532,N_21791,N_21507);
xor U32533 (N_32533,N_28187,N_23737);
and U32534 (N_32534,N_28801,N_29151);
and U32535 (N_32535,N_20358,N_23780);
and U32536 (N_32536,N_26449,N_22931);
nor U32537 (N_32537,N_20092,N_26709);
and U32538 (N_32538,N_23599,N_26646);
xnor U32539 (N_32539,N_21216,N_29420);
and U32540 (N_32540,N_23161,N_27205);
nand U32541 (N_32541,N_26365,N_24624);
or U32542 (N_32542,N_27156,N_27248);
nand U32543 (N_32543,N_29955,N_26300);
and U32544 (N_32544,N_20114,N_28268);
or U32545 (N_32545,N_23157,N_24106);
or U32546 (N_32546,N_27091,N_25441);
xnor U32547 (N_32547,N_21335,N_29310);
or U32548 (N_32548,N_25650,N_24749);
nor U32549 (N_32549,N_21416,N_22662);
or U32550 (N_32550,N_28009,N_25886);
and U32551 (N_32551,N_25592,N_24542);
or U32552 (N_32552,N_25614,N_20278);
nand U32553 (N_32553,N_20490,N_22420);
nand U32554 (N_32554,N_26440,N_20046);
nand U32555 (N_32555,N_22896,N_23022);
and U32556 (N_32556,N_27786,N_28950);
or U32557 (N_32557,N_28407,N_27011);
nand U32558 (N_32558,N_22629,N_29505);
or U32559 (N_32559,N_26235,N_24477);
xor U32560 (N_32560,N_29253,N_22968);
nor U32561 (N_32561,N_29818,N_25457);
xnor U32562 (N_32562,N_28346,N_24071);
nand U32563 (N_32563,N_24193,N_28956);
nand U32564 (N_32564,N_28093,N_25165);
and U32565 (N_32565,N_21436,N_26688);
xnor U32566 (N_32566,N_27599,N_22097);
and U32567 (N_32567,N_20826,N_28146);
or U32568 (N_32568,N_25406,N_23940);
and U32569 (N_32569,N_28884,N_27634);
or U32570 (N_32570,N_23720,N_24687);
nand U32571 (N_32571,N_20739,N_25672);
and U32572 (N_32572,N_29965,N_27178);
nor U32573 (N_32573,N_21975,N_22649);
xnor U32574 (N_32574,N_22447,N_29927);
and U32575 (N_32575,N_29386,N_20173);
nor U32576 (N_32576,N_24763,N_28105);
or U32577 (N_32577,N_27337,N_23269);
nor U32578 (N_32578,N_26945,N_27964);
or U32579 (N_32579,N_23551,N_21213);
nor U32580 (N_32580,N_20410,N_29808);
nand U32581 (N_32581,N_21391,N_27848);
xor U32582 (N_32582,N_23569,N_21828);
and U32583 (N_32583,N_23313,N_27274);
or U32584 (N_32584,N_24917,N_24680);
nor U32585 (N_32585,N_28227,N_22874);
nand U32586 (N_32586,N_20827,N_28312);
nor U32587 (N_32587,N_29529,N_25146);
or U32588 (N_32588,N_23619,N_24561);
or U32589 (N_32589,N_25267,N_26205);
or U32590 (N_32590,N_26010,N_21398);
or U32591 (N_32591,N_20725,N_20066);
xor U32592 (N_32592,N_23865,N_26307);
xor U32593 (N_32593,N_20362,N_25026);
or U32594 (N_32594,N_22211,N_24422);
or U32595 (N_32595,N_29270,N_22873);
nor U32596 (N_32596,N_27899,N_20869);
or U32597 (N_32597,N_23791,N_29018);
nand U32598 (N_32598,N_20312,N_29909);
xor U32599 (N_32599,N_29285,N_21426);
xnor U32600 (N_32600,N_21759,N_25900);
and U32601 (N_32601,N_25701,N_29509);
nor U32602 (N_32602,N_27290,N_27643);
nor U32603 (N_32603,N_28357,N_21618);
or U32604 (N_32604,N_26633,N_20613);
nor U32605 (N_32605,N_28230,N_22927);
nand U32606 (N_32606,N_22145,N_26504);
xnor U32607 (N_32607,N_29874,N_23306);
and U32608 (N_32608,N_28599,N_21858);
and U32609 (N_32609,N_27212,N_20010);
and U32610 (N_32610,N_20040,N_27604);
nand U32611 (N_32611,N_28411,N_21313);
nand U32612 (N_32612,N_27470,N_28621);
nor U32613 (N_32613,N_23631,N_20089);
nor U32614 (N_32614,N_25140,N_20349);
nand U32615 (N_32615,N_25949,N_25190);
nor U32616 (N_32616,N_25726,N_27322);
nor U32617 (N_32617,N_26730,N_23070);
xor U32618 (N_32618,N_28150,N_23464);
or U32619 (N_32619,N_29688,N_29609);
nand U32620 (N_32620,N_29078,N_23986);
or U32621 (N_32621,N_29486,N_25523);
and U32622 (N_32622,N_26548,N_21259);
nand U32623 (N_32623,N_23283,N_21655);
xnor U32624 (N_32624,N_24533,N_21963);
or U32625 (N_32625,N_27742,N_26425);
nor U32626 (N_32626,N_27237,N_28443);
nor U32627 (N_32627,N_24342,N_29970);
xor U32628 (N_32628,N_24139,N_23410);
and U32629 (N_32629,N_23248,N_20993);
xnor U32630 (N_32630,N_28211,N_20188);
nor U32631 (N_32631,N_28315,N_28542);
and U32632 (N_32632,N_26705,N_25023);
or U32633 (N_32633,N_29986,N_21763);
or U32634 (N_32634,N_28862,N_27419);
and U32635 (N_32635,N_25212,N_29118);
nand U32636 (N_32636,N_24876,N_21673);
or U32637 (N_32637,N_28253,N_28163);
nor U32638 (N_32638,N_26276,N_27046);
or U32639 (N_32639,N_27760,N_20285);
nor U32640 (N_32640,N_29065,N_22272);
and U32641 (N_32641,N_29063,N_22489);
xnor U32642 (N_32642,N_27738,N_24018);
nor U32643 (N_32643,N_28115,N_22225);
or U32644 (N_32644,N_25059,N_26642);
nand U32645 (N_32645,N_23968,N_26155);
nor U32646 (N_32646,N_23875,N_25576);
nor U32647 (N_32647,N_27910,N_29706);
or U32648 (N_32648,N_25516,N_26085);
xnor U32649 (N_32649,N_23347,N_28363);
xor U32650 (N_32650,N_28323,N_21658);
nand U32651 (N_32651,N_28075,N_21786);
nor U32652 (N_32652,N_26846,N_29513);
nand U32653 (N_32653,N_24740,N_22846);
or U32654 (N_32654,N_27443,N_25847);
nand U32655 (N_32655,N_24626,N_27291);
and U32656 (N_32656,N_22104,N_21061);
nor U32657 (N_32657,N_23625,N_29828);
and U32658 (N_32658,N_27458,N_28977);
and U32659 (N_32659,N_26051,N_20967);
and U32660 (N_32660,N_28011,N_20019);
and U32661 (N_32661,N_28553,N_22474);
nor U32662 (N_32662,N_23305,N_20439);
nand U32663 (N_32663,N_25856,N_21896);
xor U32664 (N_32664,N_23996,N_21352);
nor U32665 (N_32665,N_21745,N_21613);
nor U32666 (N_32666,N_24557,N_23104);
xnor U32667 (N_32667,N_26014,N_23377);
nor U32668 (N_32668,N_24069,N_24228);
nand U32669 (N_32669,N_22772,N_22899);
and U32670 (N_32670,N_25454,N_27589);
nor U32671 (N_32671,N_29333,N_28987);
or U32672 (N_32672,N_21606,N_25100);
or U32673 (N_32673,N_28601,N_28905);
or U32674 (N_32674,N_29701,N_29900);
and U32675 (N_32675,N_27725,N_26913);
or U32676 (N_32676,N_24838,N_24748);
or U32677 (N_32677,N_29662,N_27007);
nor U32678 (N_32678,N_23672,N_28997);
nor U32679 (N_32679,N_26349,N_22170);
nand U32680 (N_32680,N_28759,N_22098);
and U32681 (N_32681,N_29239,N_29077);
xor U32682 (N_32682,N_21253,N_21058);
and U32683 (N_32683,N_28119,N_29614);
nor U32684 (N_32684,N_21116,N_28720);
and U32685 (N_32685,N_25864,N_20008);
and U32686 (N_32686,N_22901,N_22975);
and U32687 (N_32687,N_22128,N_25613);
nor U32688 (N_32688,N_20828,N_28695);
or U32689 (N_32689,N_28188,N_24162);
nor U32690 (N_32690,N_21256,N_22110);
nor U32691 (N_32691,N_22362,N_21481);
nand U32692 (N_32692,N_27071,N_26135);
nand U32693 (N_32693,N_27130,N_20259);
nand U32694 (N_32694,N_25605,N_24243);
and U32695 (N_32695,N_29962,N_25959);
nand U32696 (N_32696,N_20749,N_22082);
xnor U32697 (N_32697,N_28507,N_20301);
xnor U32698 (N_32698,N_20148,N_24086);
or U32699 (N_32699,N_25615,N_29211);
nand U32700 (N_32700,N_24260,N_26271);
xnor U32701 (N_32701,N_26378,N_29441);
nor U32702 (N_32702,N_21619,N_23296);
or U32703 (N_32703,N_26448,N_29645);
xor U32704 (N_32704,N_24597,N_27840);
or U32705 (N_32705,N_20268,N_21783);
nand U32706 (N_32706,N_29436,N_27312);
xnor U32707 (N_32707,N_24539,N_27469);
or U32708 (N_32708,N_24130,N_22559);
and U32709 (N_32709,N_27681,N_25837);
nor U32710 (N_32710,N_24377,N_24306);
and U32711 (N_32711,N_28581,N_27171);
nor U32712 (N_32712,N_29902,N_27309);
and U32713 (N_32713,N_20434,N_24383);
and U32714 (N_32714,N_25706,N_25758);
nand U32715 (N_32715,N_29334,N_21664);
or U32716 (N_32716,N_26758,N_23547);
nor U32717 (N_32717,N_23320,N_23263);
nand U32718 (N_32718,N_29342,N_27254);
nand U32719 (N_32719,N_25803,N_26067);
nand U32720 (N_32720,N_21024,N_26684);
and U32721 (N_32721,N_28267,N_27380);
or U32722 (N_32722,N_20953,N_21202);
nor U32723 (N_32723,N_25869,N_21938);
xnor U32724 (N_32724,N_20061,N_23340);
nor U32725 (N_32725,N_27703,N_28813);
xnor U32726 (N_32726,N_28487,N_24016);
xor U32727 (N_32727,N_29644,N_28566);
or U32728 (N_32728,N_24411,N_28483);
xnor U32729 (N_32729,N_28534,N_29782);
xnor U32730 (N_32730,N_29717,N_26324);
nor U32731 (N_32731,N_29408,N_27833);
and U32732 (N_32732,N_23941,N_23843);
xor U32733 (N_32733,N_28978,N_24565);
or U32734 (N_32734,N_21376,N_23868);
xnor U32735 (N_32735,N_24609,N_23166);
nand U32736 (N_32736,N_25583,N_24829);
or U32737 (N_32737,N_23564,N_21319);
nor U32738 (N_32738,N_24338,N_29432);
or U32739 (N_32739,N_23966,N_20196);
xor U32740 (N_32740,N_26669,N_21968);
or U32741 (N_32741,N_23479,N_21937);
nor U32742 (N_32742,N_20576,N_25265);
or U32743 (N_32743,N_27192,N_25294);
and U32744 (N_32744,N_29820,N_29906);
and U32745 (N_32745,N_21302,N_24979);
xnor U32746 (N_32746,N_23893,N_21163);
or U32747 (N_32747,N_24963,N_20401);
xor U32748 (N_32748,N_20124,N_26413);
and U32749 (N_32749,N_27438,N_27717);
nor U32750 (N_32750,N_24551,N_23924);
xnor U32751 (N_32751,N_20773,N_21964);
or U32752 (N_32752,N_28504,N_21161);
or U32753 (N_32753,N_23423,N_26522);
or U32754 (N_32754,N_28795,N_24949);
xnor U32755 (N_32755,N_20415,N_26612);
nand U32756 (N_32756,N_23787,N_23453);
or U32757 (N_32757,N_22039,N_21756);
or U32758 (N_32758,N_23221,N_20132);
nor U32759 (N_32759,N_29101,N_27460);
and U32760 (N_32760,N_28781,N_26974);
nor U32761 (N_32761,N_27626,N_24738);
or U32762 (N_32762,N_23037,N_20639);
nor U32763 (N_32763,N_26572,N_20738);
and U32764 (N_32764,N_29170,N_21392);
and U32765 (N_32765,N_29043,N_28081);
or U32766 (N_32766,N_27500,N_29164);
or U32767 (N_32767,N_20578,N_23199);
xnor U32768 (N_32768,N_24488,N_27921);
xor U32769 (N_32769,N_20862,N_20298);
nand U32770 (N_32770,N_29870,N_29175);
nand U32771 (N_32771,N_25130,N_28132);
xor U32772 (N_32772,N_23859,N_22883);
nand U32773 (N_32773,N_25855,N_22652);
xnor U32774 (N_32774,N_26864,N_23165);
xnor U32775 (N_32775,N_29466,N_20236);
xor U32776 (N_32776,N_29864,N_27956);
nor U32777 (N_32777,N_24131,N_29737);
or U32778 (N_32778,N_25154,N_28823);
nand U32779 (N_32779,N_22402,N_24822);
or U32780 (N_32780,N_27940,N_23923);
xor U32781 (N_32781,N_23972,N_20670);
xor U32782 (N_32782,N_22298,N_28518);
or U32783 (N_32783,N_26806,N_24938);
or U32784 (N_32784,N_25529,N_27962);
xnor U32785 (N_32785,N_23627,N_28482);
nand U32786 (N_32786,N_27957,N_26462);
or U32787 (N_32787,N_26409,N_27907);
and U32788 (N_32788,N_20244,N_28770);
or U32789 (N_32789,N_26607,N_21712);
nor U32790 (N_32790,N_23257,N_25860);
and U32791 (N_32791,N_29395,N_20742);
nor U32792 (N_32792,N_25414,N_20481);
or U32793 (N_32793,N_22309,N_27397);
nor U32794 (N_32794,N_22155,N_25053);
nor U32795 (N_32795,N_27902,N_23708);
or U32796 (N_32796,N_23499,N_25451);
and U32797 (N_32797,N_20186,N_28090);
and U32798 (N_32798,N_27013,N_24044);
or U32799 (N_32799,N_21902,N_25047);
nand U32800 (N_32800,N_25369,N_29154);
xor U32801 (N_32801,N_22543,N_26022);
xor U32802 (N_32802,N_24573,N_20642);
nor U32803 (N_32803,N_27925,N_28370);
nor U32804 (N_32804,N_28653,N_22096);
nand U32805 (N_32805,N_23131,N_21815);
xnor U32806 (N_32806,N_23268,N_29394);
xor U32807 (N_32807,N_21675,N_28130);
nor U32808 (N_32808,N_24812,N_22717);
and U32809 (N_32809,N_27637,N_25183);
and U32810 (N_32810,N_26984,N_20644);
nor U32811 (N_32811,N_26947,N_27989);
nor U32812 (N_32812,N_20561,N_21603);
nor U32813 (N_32813,N_29213,N_27951);
and U32814 (N_32814,N_29840,N_26439);
and U32815 (N_32815,N_24054,N_29109);
or U32816 (N_32816,N_24452,N_21789);
nor U32817 (N_32817,N_22839,N_21705);
nor U32818 (N_32818,N_22520,N_25698);
or U32819 (N_32819,N_21561,N_28031);
and U32820 (N_32820,N_29379,N_26494);
nor U32821 (N_32821,N_27289,N_22753);
nor U32822 (N_32822,N_25387,N_27283);
or U32823 (N_32823,N_26841,N_28575);
and U32824 (N_32824,N_25330,N_23074);
nor U32825 (N_32825,N_22287,N_29929);
nor U32826 (N_32826,N_20044,N_27780);
nand U32827 (N_32827,N_25898,N_23732);
or U32828 (N_32828,N_29619,N_28471);
or U32829 (N_32829,N_23563,N_26184);
nor U32830 (N_32830,N_27160,N_25355);
nand U32831 (N_32831,N_28314,N_20902);
and U32832 (N_32832,N_27474,N_25407);
nor U32833 (N_32833,N_20134,N_24855);
or U32834 (N_32834,N_25547,N_26003);
nand U32835 (N_32835,N_27768,N_25468);
xor U32836 (N_32836,N_29871,N_26659);
or U32837 (N_32837,N_28438,N_29877);
nand U32838 (N_32838,N_26783,N_20474);
xnor U32839 (N_32839,N_28775,N_24479);
or U32840 (N_32840,N_27359,N_22678);
xor U32841 (N_32841,N_25519,N_27287);
and U32842 (N_32842,N_22814,N_20524);
nor U32843 (N_32843,N_20323,N_20247);
xor U32844 (N_32844,N_21227,N_29103);
nor U32845 (N_32845,N_28066,N_25586);
nand U32846 (N_32846,N_24589,N_27813);
xor U32847 (N_32847,N_28024,N_23522);
xnor U32848 (N_32848,N_24564,N_28080);
and U32849 (N_32849,N_26994,N_23033);
or U32850 (N_32850,N_25354,N_26195);
nand U32851 (N_32851,N_20655,N_22463);
and U32852 (N_32852,N_26305,N_27545);
and U32853 (N_32853,N_24208,N_26935);
or U32854 (N_32854,N_26239,N_28549);
xor U32855 (N_32855,N_27557,N_20692);
or U32856 (N_32856,N_23385,N_26847);
nor U32857 (N_32857,N_20977,N_26160);
nand U32858 (N_32858,N_22747,N_20581);
xnor U32859 (N_32859,N_23957,N_27262);
nand U32860 (N_32860,N_21944,N_20932);
or U32861 (N_32861,N_29723,N_21942);
and U32862 (N_32862,N_22811,N_28208);
nor U32863 (N_32863,N_28364,N_28729);
and U32864 (N_32864,N_22069,N_27139);
xnor U32865 (N_32865,N_24163,N_25704);
nand U32866 (N_32866,N_27182,N_21475);
and U32867 (N_32867,N_27376,N_26749);
xor U32868 (N_32868,N_25719,N_20802);
or U32869 (N_32869,N_22315,N_22382);
and U32870 (N_32870,N_23027,N_22593);
nor U32871 (N_32871,N_21823,N_28309);
xnor U32872 (N_32872,N_26687,N_27708);
nand U32873 (N_32873,N_25774,N_29321);
or U32874 (N_32874,N_27119,N_22136);
and U32875 (N_32875,N_21154,N_20658);
and U32876 (N_32876,N_28265,N_26395);
nor U32877 (N_32877,N_28562,N_26151);
xnor U32878 (N_32878,N_25176,N_27098);
xnor U32879 (N_32879,N_23858,N_23000);
xnor U32880 (N_32880,N_21558,N_20935);
or U32881 (N_32881,N_21456,N_29426);
nand U32882 (N_32882,N_22758,N_27190);
nand U32883 (N_32883,N_28404,N_23497);
nor U32884 (N_32884,N_21795,N_23182);
or U32885 (N_32885,N_25751,N_26316);
or U32886 (N_32886,N_29578,N_23180);
or U32887 (N_32887,N_24971,N_22972);
nand U32888 (N_32888,N_20623,N_22000);
nor U32889 (N_32889,N_29592,N_26477);
nand U32890 (N_32890,N_23576,N_28327);
or U32891 (N_32891,N_20797,N_26360);
and U32892 (N_32892,N_21819,N_25910);
nor U32893 (N_32893,N_21400,N_22780);
xor U32894 (N_32894,N_22341,N_22257);
or U32895 (N_32895,N_22144,N_22505);
nand U32896 (N_32896,N_21150,N_29996);
or U32897 (N_32897,N_22487,N_28435);
xnor U32898 (N_32898,N_28586,N_29359);
xor U32899 (N_32899,N_24514,N_27257);
or U32900 (N_32900,N_21180,N_21739);
nor U32901 (N_32901,N_29998,N_21265);
xor U32902 (N_32902,N_24846,N_22221);
and U32903 (N_32903,N_27572,N_23452);
or U32904 (N_32904,N_20943,N_29732);
or U32905 (N_32905,N_20516,N_25056);
nor U32906 (N_32906,N_20386,N_20532);
or U32907 (N_32907,N_26549,N_26739);
or U32908 (N_32908,N_25964,N_20238);
and U32909 (N_32909,N_25328,N_27999);
and U32910 (N_32910,N_20687,N_27476);
nand U32911 (N_32911,N_28809,N_20257);
or U32912 (N_32912,N_23181,N_23503);
nand U32913 (N_32913,N_22025,N_29704);
xnor U32914 (N_32914,N_29283,N_23216);
or U32915 (N_32915,N_25566,N_27569);
nand U32916 (N_32916,N_28401,N_20164);
nand U32917 (N_32917,N_28859,N_24404);
nand U32918 (N_32918,N_25117,N_26807);
nand U32919 (N_32919,N_27673,N_28568);
nand U32920 (N_32920,N_25142,N_28800);
nor U32921 (N_32921,N_23544,N_27707);
xnor U32922 (N_32922,N_23222,N_29672);
and U32923 (N_32923,N_27904,N_23103);
xor U32924 (N_32924,N_22479,N_20736);
or U32925 (N_32925,N_29552,N_27984);
or U32926 (N_32926,N_20437,N_21334);
nor U32927 (N_32927,N_23314,N_21695);
nor U32928 (N_32928,N_23042,N_26274);
xnor U32929 (N_32929,N_27308,N_27477);
xor U32930 (N_32930,N_25826,N_21045);
nand U32931 (N_32931,N_28753,N_28670);
or U32932 (N_32932,N_27102,N_29597);
or U32933 (N_32933,N_28397,N_23614);
or U32934 (N_32934,N_28071,N_29173);
and U32935 (N_32935,N_20660,N_28114);
xor U32936 (N_32936,N_20075,N_25732);
or U32937 (N_32937,N_26814,N_20030);
xor U32938 (N_32938,N_26782,N_24219);
or U32939 (N_32939,N_24773,N_28147);
xnor U32940 (N_32940,N_27452,N_28543);
xor U32941 (N_32941,N_20995,N_26857);
or U32942 (N_32942,N_22932,N_22815);
or U32943 (N_32943,N_26588,N_28353);
nand U32944 (N_32944,N_29031,N_27883);
xor U32945 (N_32945,N_20946,N_29735);
nor U32946 (N_32946,N_29363,N_28889);
xor U32947 (N_32947,N_29349,N_29041);
nor U32948 (N_32948,N_23754,N_24109);
xor U32949 (N_32949,N_22157,N_27054);
or U32950 (N_32950,N_23697,N_20368);
and U32951 (N_32951,N_23508,N_22050);
and U32952 (N_32952,N_27336,N_22508);
xnor U32953 (N_32953,N_28160,N_24456);
nor U32954 (N_32954,N_24294,N_27440);
xnor U32955 (N_32955,N_23372,N_28516);
nor U32956 (N_32956,N_29003,N_27581);
and U32957 (N_32957,N_25105,N_26419);
or U32958 (N_32958,N_29209,N_23186);
nand U32959 (N_32959,N_25830,N_24039);
or U32960 (N_32960,N_24571,N_28116);
nand U32961 (N_32961,N_21808,N_25926);
and U32962 (N_32962,N_26851,N_21861);
or U32963 (N_32963,N_23827,N_28589);
nand U32964 (N_32964,N_21515,N_29941);
and U32965 (N_32965,N_27232,N_24476);
nand U32966 (N_32966,N_24668,N_20784);
and U32967 (N_32967,N_20675,N_26328);
nor U32968 (N_32968,N_25459,N_24595);
nor U32969 (N_32969,N_28334,N_23234);
nand U32970 (N_32970,N_25107,N_26674);
or U32971 (N_32971,N_27839,N_23871);
nand U32972 (N_32972,N_20728,N_24702);
nand U32973 (N_32973,N_29001,N_25061);
nand U32974 (N_32974,N_21498,N_27778);
or U32975 (N_32975,N_26459,N_23961);
nor U32976 (N_32976,N_20237,N_26819);
nor U32977 (N_32977,N_20340,N_21638);
xor U32978 (N_32978,N_28101,N_22669);
nand U32979 (N_32979,N_22199,N_25379);
nor U32980 (N_32980,N_22643,N_23212);
or U32981 (N_32981,N_27486,N_20538);
or U32982 (N_32982,N_29632,N_21941);
nor U32983 (N_32983,N_25690,N_22205);
xnor U32984 (N_32984,N_28726,N_23556);
nand U32985 (N_32985,N_20485,N_26853);
or U32986 (N_32986,N_20897,N_21337);
nand U32987 (N_32987,N_24380,N_29025);
xnor U32988 (N_32988,N_28909,N_21189);
nor U32989 (N_32989,N_28016,N_20297);
xor U32990 (N_32990,N_23367,N_28027);
or U32991 (N_32991,N_22193,N_24164);
and U32992 (N_32992,N_26506,N_22844);
nand U32993 (N_32993,N_28731,N_27612);
and U32994 (N_32994,N_28272,N_22118);
and U32995 (N_32995,N_21278,N_21291);
nand U32996 (N_32996,N_22638,N_24882);
nor U32997 (N_32997,N_21709,N_29567);
and U32998 (N_32998,N_20896,N_20691);
nand U32999 (N_32999,N_28195,N_29440);
nand U33000 (N_33000,N_27953,N_22861);
nand U33001 (N_33001,N_25538,N_21728);
and U33002 (N_33002,N_21796,N_22446);
xor U33003 (N_33003,N_24410,N_25173);
and U33004 (N_33004,N_29265,N_25371);
nand U33005 (N_33005,N_26366,N_23511);
and U33006 (N_33006,N_26756,N_25551);
nor U33007 (N_33007,N_25688,N_28332);
or U33008 (N_33008,N_27885,N_29038);
xor U33009 (N_33009,N_27556,N_24305);
and U33010 (N_33010,N_24226,N_26297);
nor U33011 (N_33011,N_23400,N_23357);
and U33012 (N_33012,N_21787,N_24292);
and U33013 (N_33013,N_28649,N_21421);
nand U33014 (N_33014,N_24708,N_20214);
and U33015 (N_33015,N_25204,N_23040);
or U33016 (N_33016,N_22058,N_29803);
nor U33017 (N_33017,N_29343,N_28874);
nand U33018 (N_33018,N_25479,N_29139);
or U33019 (N_33019,N_28700,N_28513);
or U33020 (N_33020,N_24555,N_26356);
xor U33021 (N_33021,N_24751,N_27145);
and U33022 (N_33022,N_20702,N_26569);
and U33023 (N_33023,N_27749,N_29683);
or U33024 (N_33024,N_21648,N_26800);
nor U33025 (N_33025,N_29050,N_24883);
and U33026 (N_33026,N_20627,N_23095);
or U33027 (N_33027,N_22281,N_27138);
and U33028 (N_33028,N_24375,N_28749);
or U33029 (N_33029,N_24079,N_24412);
nor U33030 (N_33030,N_24000,N_27733);
xnor U33031 (N_33031,N_23154,N_29634);
xor U33032 (N_33032,N_21680,N_21836);
nor U33033 (N_33033,N_29669,N_27364);
nand U33034 (N_33034,N_26337,N_29747);
nand U33035 (N_33035,N_22410,N_24888);
or U33036 (N_33036,N_26555,N_25973);
or U33037 (N_33037,N_29129,N_24616);
and U33038 (N_33038,N_25531,N_25494);
nor U33039 (N_33039,N_22930,N_25641);
nand U33040 (N_33040,N_26066,N_26304);
or U33041 (N_33041,N_22448,N_20775);
xor U33042 (N_33042,N_28365,N_21168);
and U33043 (N_33043,N_24443,N_29720);
and U33044 (N_33044,N_27313,N_25323);
or U33045 (N_33045,N_29605,N_26924);
or U33046 (N_33046,N_29375,N_20805);
nor U33047 (N_33047,N_26352,N_20812);
nand U33048 (N_33048,N_25115,N_23724);
nor U33049 (N_33049,N_23469,N_28263);
xor U33050 (N_33050,N_25473,N_29097);
and U33051 (N_33051,N_24245,N_22710);
nand U33052 (N_33052,N_21472,N_25870);
nand U33053 (N_33053,N_23914,N_27382);
nand U33054 (N_33054,N_23815,N_22367);
nand U33055 (N_33055,N_29975,N_25597);
xor U33056 (N_33056,N_25315,N_26311);
nor U33057 (N_33057,N_24468,N_26907);
xor U33058 (N_33058,N_24123,N_29811);
and U33059 (N_33059,N_27042,N_25491);
nand U33060 (N_33060,N_28426,N_28895);
nand U33061 (N_33061,N_23032,N_24469);
xnor U33062 (N_33062,N_27439,N_20252);
nor U33063 (N_33063,N_25157,N_28038);
nand U33064 (N_33064,N_22765,N_25662);
nor U33065 (N_33065,N_23785,N_29042);
and U33066 (N_33066,N_27159,N_28766);
and U33067 (N_33067,N_27897,N_29724);
or U33068 (N_33068,N_29881,N_29094);
xnor U33069 (N_33069,N_23892,N_25257);
nor U33070 (N_33070,N_29765,N_22201);
nand U33071 (N_33071,N_25264,N_25306);
or U33072 (N_33072,N_23921,N_22139);
xor U33073 (N_33073,N_23749,N_23851);
nand U33074 (N_33074,N_22514,N_24316);
xor U33075 (N_33075,N_25919,N_21572);
xnor U33076 (N_33076,N_22916,N_20159);
xor U33077 (N_33077,N_21801,N_23480);
or U33078 (N_33078,N_23517,N_25505);
xnor U33079 (N_33079,N_20872,N_22774);
or U33080 (N_33080,N_24440,N_21362);
or U33081 (N_33081,N_23795,N_26717);
and U33082 (N_33082,N_22339,N_22045);
and U33083 (N_33083,N_21903,N_28185);
nor U33084 (N_33084,N_21268,N_28292);
xor U33085 (N_33085,N_20959,N_25087);
nor U33086 (N_33086,N_22925,N_22295);
and U33087 (N_33087,N_24045,N_21831);
nor U33088 (N_33088,N_25111,N_29478);
or U33089 (N_33089,N_23097,N_23857);
xor U33090 (N_33090,N_27618,N_28625);
xnor U33091 (N_33091,N_27284,N_22976);
xor U33092 (N_33092,N_26904,N_20195);
and U33093 (N_33093,N_22611,N_29961);
nand U33094 (N_33094,N_28387,N_28924);
and U33095 (N_33095,N_21018,N_23003);
or U33096 (N_33096,N_23034,N_28552);
nor U33097 (N_33097,N_23646,N_20117);
or U33098 (N_33098,N_29767,N_20637);
nand U33099 (N_33099,N_20456,N_25252);
nor U33100 (N_33100,N_24036,N_29738);
and U33101 (N_33101,N_21344,N_29617);
and U33102 (N_33102,N_21932,N_21842);
nor U33103 (N_33103,N_26043,N_23045);
nor U33104 (N_33104,N_29264,N_27928);
or U33105 (N_33105,N_28207,N_23927);
nand U33106 (N_33106,N_20937,N_21077);
or U33107 (N_33107,N_26286,N_22186);
or U33108 (N_33108,N_22460,N_26821);
nand U33109 (N_33109,N_21494,N_22346);
or U33110 (N_33110,N_21644,N_28627);
and U33111 (N_33111,N_27622,N_26455);
xor U33112 (N_33112,N_23718,N_27632);
nand U33113 (N_33113,N_22574,N_24658);
nand U33114 (N_33114,N_20560,N_20715);
xor U33115 (N_33115,N_20488,N_20611);
or U33116 (N_33116,N_26973,N_29678);
and U33117 (N_33117,N_24752,N_27209);
xor U33118 (N_33118,N_25123,N_26936);
nor U33119 (N_33119,N_26963,N_27982);
nand U33120 (N_33120,N_22651,N_26197);
nand U33121 (N_33121,N_25709,N_26347);
and U33122 (N_33122,N_24475,N_24076);
nand U33123 (N_33123,N_24107,N_21384);
nor U33124 (N_33124,N_20857,N_23188);
xor U33125 (N_33125,N_28681,N_29004);
nor U33126 (N_33126,N_21860,N_27087);
or U33127 (N_33127,N_29087,N_29852);
nor U33128 (N_33128,N_22124,N_26079);
and U33129 (N_33129,N_22270,N_26308);
nor U33130 (N_33130,N_22562,N_23683);
xor U33131 (N_33131,N_26911,N_25305);
xnor U33132 (N_33132,N_25430,N_27436);
or U33133 (N_33133,N_25391,N_26020);
nand U33134 (N_33134,N_23788,N_21127);
nand U33135 (N_33135,N_24510,N_27605);
nor U33136 (N_33136,N_24057,N_22188);
and U33137 (N_33137,N_27003,N_26475);
or U33138 (N_33138,N_23266,N_25978);
and U33139 (N_33139,N_22388,N_25493);
or U33140 (N_33140,N_25999,N_26738);
and U33141 (N_33141,N_29045,N_25256);
and U33142 (N_33142,N_28667,N_25510);
or U33143 (N_33143,N_28470,N_21741);
nor U33144 (N_33144,N_29487,N_22690);
or U33145 (N_33145,N_22371,N_24795);
or U33146 (N_33146,N_25604,N_21913);
and U33147 (N_33147,N_25854,N_25170);
or U33148 (N_33148,N_27334,N_21529);
xnor U33149 (N_33149,N_20436,N_28061);
nor U33150 (N_33150,N_26698,N_20295);
nand U33151 (N_33151,N_27075,N_27103);
nand U33152 (N_33152,N_26441,N_24615);
nand U33153 (N_33153,N_27920,N_25943);
nor U33154 (N_33154,N_29827,N_24268);
and U33155 (N_33155,N_27413,N_24454);
xnor U33156 (N_33156,N_20153,N_25045);
nand U33157 (N_33157,N_20504,N_21570);
or U33158 (N_33158,N_20515,N_25051);
or U33159 (N_33159,N_27941,N_21726);
nand U33160 (N_33160,N_24753,N_25635);
xor U33161 (N_33161,N_27547,N_27201);
nand U33162 (N_33162,N_22088,N_26568);
or U33163 (N_33163,N_28244,N_23738);
xor U33164 (N_33164,N_23136,N_21169);
and U33165 (N_33165,N_25823,N_29399);
or U33166 (N_33166,N_22760,N_26315);
nor U33167 (N_33167,N_22194,N_28645);
nand U33168 (N_33168,N_22214,N_24623);
or U33169 (N_33169,N_29555,N_27523);
nor U33170 (N_33170,N_25850,N_25996);
nand U33171 (N_33171,N_29418,N_28998);
nor U33172 (N_33172,N_25984,N_27369);
nand U33173 (N_33173,N_29500,N_29409);
xor U33174 (N_33174,N_26468,N_22821);
and U33175 (N_33175,N_22084,N_23801);
xor U33176 (N_33176,N_22895,N_29307);
nand U33177 (N_33177,N_28204,N_29801);
nand U33178 (N_33178,N_22672,N_29304);
xnor U33179 (N_33179,N_21325,N_27855);
nand U33180 (N_33180,N_25394,N_23979);
xnor U33181 (N_33181,N_27039,N_25029);
or U33182 (N_33182,N_25317,N_21607);
xor U33183 (N_33183,N_21142,N_27217);
xor U33184 (N_33184,N_23360,N_29074);
xor U33185 (N_33185,N_21755,N_25799);
and U33186 (N_33186,N_26517,N_23209);
nand U33187 (N_33187,N_22151,N_25600);
nand U33188 (N_33188,N_29165,N_22940);
xor U33189 (N_33189,N_28153,N_24046);
nand U33190 (N_33190,N_23067,N_21464);
and U33191 (N_33191,N_29223,N_24913);
nand U33192 (N_33192,N_23162,N_29976);
and U33193 (N_33193,N_26825,N_29238);
xnor U33194 (N_33194,N_20517,N_26587);
and U33195 (N_33195,N_25057,N_20091);
nand U33196 (N_33196,N_23478,N_23485);
nor U33197 (N_33197,N_24368,N_24975);
nand U33198 (N_33198,N_29390,N_26713);
or U33199 (N_33199,N_29497,N_20856);
nand U33200 (N_33200,N_20332,N_22867);
or U33201 (N_33201,N_23446,N_29734);
nand U33202 (N_33202,N_27868,N_26502);
nor U33203 (N_33203,N_22494,N_25628);
and U33204 (N_33204,N_23238,N_21322);
xor U33205 (N_33205,N_22236,N_20007);
nor U33206 (N_33206,N_26712,N_23118);
xnor U33207 (N_33207,N_26581,N_22757);
or U33208 (N_33208,N_23374,N_20272);
nand U33209 (N_33209,N_20493,N_24790);
xor U33210 (N_33210,N_24503,N_26495);
xor U33211 (N_33211,N_28668,N_29191);
or U33212 (N_33212,N_20109,N_25515);
nand U33213 (N_33213,N_22106,N_29260);
nand U33214 (N_33214,N_20809,N_29456);
xnor U33215 (N_33215,N_27682,N_20169);
nor U33216 (N_33216,N_22732,N_23746);
xnor U33217 (N_33217,N_21887,N_24659);
and U33218 (N_33218,N_27242,N_24025);
and U33219 (N_33219,N_24711,N_27689);
xor U33220 (N_33220,N_21071,N_25139);
nor U33221 (N_33221,N_20666,N_23143);
xor U33222 (N_33222,N_28955,N_28246);
xor U33223 (N_33223,N_24665,N_27015);
nand U33224 (N_33224,N_27365,N_24900);
xor U33225 (N_33225,N_22607,N_24363);
and U33226 (N_33226,N_26987,N_26350);
and U33227 (N_33227,N_26069,N_25163);
nand U33228 (N_33228,N_25518,N_28259);
nand U33229 (N_33229,N_27507,N_21338);
xor U33230 (N_33230,N_20250,N_23862);
nor U33231 (N_33231,N_20548,N_22266);
and U33232 (N_33232,N_24990,N_25444);
xnor U33233 (N_33233,N_27204,N_27562);
or U33234 (N_33234,N_25250,N_26138);
nor U33235 (N_33235,N_25018,N_28544);
nand U33236 (N_33236,N_21704,N_29989);
or U33237 (N_33237,N_24299,N_20230);
nand U33238 (N_33238,N_23011,N_27482);
nor U33239 (N_33239,N_29860,N_21805);
or U33240 (N_33240,N_22936,N_23874);
xor U33241 (N_33241,N_24320,N_28510);
xor U33242 (N_33242,N_20483,N_20847);
or U33243 (N_33243,N_20597,N_25832);
or U33244 (N_33244,N_28193,N_26824);
and U33245 (N_33245,N_21993,N_25411);
nor U33246 (N_33246,N_22898,N_27564);
nand U33247 (N_33247,N_22391,N_22329);
and U33248 (N_33248,N_27825,N_25718);
nor U33249 (N_33249,N_25899,N_23031);
or U33250 (N_33250,N_28213,N_26257);
xor U33251 (N_33251,N_23403,N_26156);
nand U33252 (N_33252,N_26722,N_28751);
and U33253 (N_33253,N_29872,N_23973);
or U33254 (N_33254,N_25805,N_27152);
and U33255 (N_33255,N_29488,N_28696);
nand U33256 (N_33256,N_24358,N_22893);
xor U33257 (N_33257,N_29698,N_22859);
nor U33258 (N_33258,N_25922,N_25863);
and U33259 (N_33259,N_22823,N_23090);
xnor U33260 (N_33260,N_24173,N_22934);
nor U33261 (N_33261,N_24677,N_22228);
and U33262 (N_33262,N_21767,N_22486);
or U33263 (N_33263,N_23465,N_29832);
xor U33264 (N_33264,N_27642,N_22473);
or U33265 (N_33265,N_20313,N_23818);
xnor U33266 (N_33266,N_21234,N_25560);
xnor U33267 (N_33267,N_28372,N_21167);
and U33268 (N_33268,N_25400,N_29305);
nor U33269 (N_33269,N_29388,N_27560);
xnor U33270 (N_33270,N_25270,N_23294);
xor U33271 (N_33271,N_24406,N_20427);
nor U33272 (N_33272,N_24331,N_25587);
or U33273 (N_33273,N_22885,N_22100);
nor U33274 (N_33274,N_28937,N_20882);
nand U33275 (N_33275,N_24512,N_23273);
or U33276 (N_33276,N_23775,N_22563);
or U33277 (N_33277,N_28878,N_21380);
and U33278 (N_33278,N_29026,N_21408);
or U33279 (N_33279,N_21151,N_23820);
nand U33280 (N_33280,N_22268,N_27161);
or U33281 (N_33281,N_25739,N_23650);
nand U33282 (N_33282,N_24816,N_20316);
and U33283 (N_33283,N_23267,N_26373);
nand U33284 (N_33284,N_25618,N_26219);
xnor U33285 (N_33285,N_26484,N_23626);
nand U33286 (N_33286,N_23149,N_22615);
nor U33287 (N_33287,N_25363,N_22101);
nor U33288 (N_33288,N_20870,N_25412);
nand U33289 (N_33289,N_27732,N_21087);
nand U33290 (N_33290,N_29981,N_25765);
nor U33291 (N_33291,N_20001,N_24854);
nand U33292 (N_33292,N_24845,N_28709);
or U33293 (N_33293,N_24689,N_21346);
or U33294 (N_33294,N_22066,N_21121);
nand U33295 (N_33295,N_20618,N_20845);
and U33296 (N_33296,N_27329,N_26740);
or U33297 (N_33297,N_23225,N_24293);
nand U33298 (N_33298,N_24156,N_28873);
or U33299 (N_33299,N_28261,N_23171);
nand U33300 (N_33300,N_23146,N_29931);
nor U33301 (N_33301,N_29159,N_27263);
and U33302 (N_33302,N_27141,N_24017);
nand U33303 (N_33303,N_23500,N_22267);
nand U33304 (N_33304,N_20264,N_23735);
nand U33305 (N_33305,N_23325,N_29234);
or U33306 (N_33306,N_29854,N_20621);
and U33307 (N_33307,N_23310,N_25336);
or U33308 (N_33308,N_27064,N_25872);
nand U33309 (N_33309,N_21737,N_25649);
nand U33310 (N_33310,N_21962,N_22400);
nand U33311 (N_33311,N_29068,N_24416);
nand U33312 (N_33312,N_25927,N_25993);
or U33313 (N_33313,N_28876,N_21228);
xor U33314 (N_33314,N_27835,N_29910);
nand U33315 (N_33315,N_29889,N_20864);
and U33316 (N_33316,N_24908,N_21438);
and U33317 (N_33317,N_20199,N_29733);
and U33318 (N_33318,N_21579,N_29507);
nor U33319 (N_33319,N_22105,N_28765);
nor U33320 (N_33320,N_23428,N_24873);
and U33321 (N_33321,N_27896,N_21678);
nor U33322 (N_33322,N_21665,N_23153);
or U33323 (N_33323,N_28294,N_24186);
nand U33324 (N_33324,N_27236,N_22534);
nor U33325 (N_33325,N_22469,N_28931);
or U33326 (N_33326,N_20183,N_23416);
nand U33327 (N_33327,N_22704,N_21372);
or U33328 (N_33328,N_29245,N_20711);
and U33329 (N_33329,N_29771,N_29166);
and U33330 (N_33330,N_27089,N_22140);
xor U33331 (N_33331,N_24132,N_22335);
xnor U33332 (N_33332,N_27924,N_22033);
nor U33333 (N_33333,N_28303,N_22545);
nor U33334 (N_33334,N_21557,N_23777);
nand U33335 (N_33335,N_26367,N_26562);
or U33336 (N_33336,N_22456,N_22036);
xor U33337 (N_33337,N_29898,N_24207);
or U33338 (N_33338,N_23366,N_28890);
and U33339 (N_33339,N_26421,N_25484);
xor U33340 (N_33340,N_25226,N_28233);
nor U33341 (N_33341,N_22794,N_20375);
or U33342 (N_33342,N_21217,N_21582);
and U33343 (N_33343,N_29128,N_21589);
xnor U33344 (N_33344,N_27948,N_22887);
and U33345 (N_33345,N_26961,N_26552);
and U33346 (N_33346,N_29210,N_27350);
or U33347 (N_33347,N_21214,N_23084);
nor U33348 (N_33348,N_21038,N_25678);
nor U33349 (N_33349,N_27275,N_26314);
and U33350 (N_33350,N_28579,N_21833);
xor U33351 (N_33351,N_23155,N_24649);
xor U33352 (N_33352,N_26711,N_20547);
nor U33353 (N_33353,N_22850,N_27973);
xnor U33354 (N_33354,N_28458,N_26537);
xor U33355 (N_33355,N_25514,N_25846);
nor U33356 (N_33356,N_22918,N_23726);
and U33357 (N_33357,N_24417,N_22535);
nand U33358 (N_33358,N_21339,N_20327);
or U33359 (N_33359,N_26299,N_24202);
or U33360 (N_33360,N_22797,N_23451);
nand U33361 (N_33361,N_22878,N_20868);
nand U33362 (N_33362,N_28125,N_26260);
or U33363 (N_33363,N_27008,N_29449);
and U33364 (N_33364,N_25680,N_28682);
and U33365 (N_33365,N_29106,N_29083);
and U33366 (N_33366,N_22263,N_22966);
or U33367 (N_33367,N_23929,N_25887);
nor U33368 (N_33368,N_22755,N_28536);
xor U33369 (N_33369,N_26761,N_29445);
xor U33370 (N_33370,N_20322,N_27625);
nor U33371 (N_33371,N_20794,N_23178);
and U33372 (N_33372,N_26045,N_24121);
and U33373 (N_33373,N_22357,N_29893);
or U33374 (N_33374,N_26482,N_25497);
or U33375 (N_33375,N_23908,N_23029);
and U33376 (N_33376,N_20248,N_29005);
or U33377 (N_33377,N_23386,N_24516);
or U33378 (N_33378,N_22417,N_21539);
xnor U33379 (N_33379,N_23905,N_21035);
or U33380 (N_33380,N_21304,N_27045);
xnor U33381 (N_33381,N_27852,N_21862);
nand U33382 (N_33382,N_29762,N_26258);
xor U33383 (N_33383,N_26887,N_26526);
nand U33384 (N_33384,N_21290,N_20726);
xnor U33385 (N_33385,N_21238,N_22769);
and U33386 (N_33386,N_27086,N_28145);
xnor U33387 (N_33387,N_22375,N_22548);
or U33388 (N_33388,N_25248,N_29471);
nor U33389 (N_33389,N_29562,N_21430);
nand U33390 (N_33390,N_22756,N_28469);
or U33391 (N_33391,N_20440,N_27942);
or U33392 (N_33392,N_21327,N_27755);
nand U33393 (N_33393,N_21578,N_23755);
and U33394 (N_33394,N_29992,N_21089);
xnor U33395 (N_33395,N_29252,N_27529);
and U33396 (N_33396,N_29663,N_25151);
nand U33397 (N_33397,N_27321,N_23623);
or U33398 (N_33398,N_27993,N_28712);
nor U33399 (N_33399,N_24717,N_24405);
nor U33400 (N_33400,N_25449,N_29805);
and U33401 (N_33401,N_27123,N_28826);
nand U33402 (N_33402,N_25161,N_26136);
xor U33403 (N_33403,N_21895,N_20620);
or U33404 (N_33404,N_20063,N_21555);
and U33405 (N_33405,N_26429,N_26855);
and U33406 (N_33406,N_26590,N_21242);
xor U33407 (N_33407,N_25058,N_21580);
and U33408 (N_33408,N_22091,N_29224);
nand U33409 (N_33409,N_25761,N_21350);
xnor U33410 (N_33410,N_26293,N_28131);
nor U33411 (N_33411,N_26320,N_26198);
nand U33412 (N_33412,N_20608,N_23611);
xor U33413 (N_33413,N_22012,N_29120);
or U33414 (N_33414,N_20927,N_29293);
xnor U33415 (N_33415,N_24160,N_27370);
nand U33416 (N_33416,N_22275,N_20225);
nand U33417 (N_33417,N_21480,N_24227);
nand U33418 (N_33418,N_21591,N_27455);
nand U33419 (N_33419,N_20549,N_21375);
or U33420 (N_33420,N_25049,N_22644);
and U33421 (N_33421,N_29633,N_20758);
or U33422 (N_33422,N_29680,N_28560);
nor U33423 (N_33423,N_20719,N_29791);
or U33424 (N_33424,N_27348,N_29006);
or U33425 (N_33425,N_22203,N_28737);
xor U33426 (N_33426,N_27449,N_24502);
xnor U33427 (N_33427,N_21800,N_23444);
nor U33428 (N_33428,N_23208,N_20632);
nand U33429 (N_33429,N_27256,N_26128);
and U33430 (N_33430,N_23016,N_21371);
nand U33431 (N_33431,N_25700,N_25866);
or U33432 (N_33432,N_29206,N_22403);
nand U33433 (N_33433,N_29532,N_24379);
or U33434 (N_33434,N_21948,N_27404);
and U33435 (N_33435,N_27478,N_27863);
xor U33436 (N_33436,N_20765,N_27577);
and U33437 (N_33437,N_28455,N_29073);
nand U33438 (N_33438,N_27142,N_27818);
nor U33439 (N_33439,N_20211,N_20102);
xnor U33440 (N_33440,N_20243,N_27349);
nor U33441 (N_33441,N_22390,N_23211);
nor U33442 (N_33442,N_26704,N_21994);
xnor U33443 (N_33443,N_28165,N_28300);
xor U33444 (N_33444,N_26427,N_23558);
nand U33445 (N_33445,N_28210,N_22171);
or U33446 (N_33446,N_20122,N_26576);
xnor U33447 (N_33447,N_29679,N_24613);
and U33448 (N_33448,N_23571,N_28084);
and U33449 (N_33449,N_23705,N_28557);
and U33450 (N_33450,N_27592,N_29279);
nand U33451 (N_33451,N_23176,N_26456);
and U33452 (N_33452,N_24685,N_28902);
xor U33453 (N_33453,N_24344,N_27929);
xor U33454 (N_33454,N_22233,N_29856);
and U33455 (N_33455,N_23036,N_21342);
and U33456 (N_33456,N_29914,N_28563);
or U33457 (N_33457,N_27841,N_23330);
nand U33458 (N_33458,N_22670,N_21826);
or U33459 (N_33459,N_27715,N_26363);
or U33460 (N_33460,N_26626,N_27001);
and U33461 (N_33461,N_27891,N_29510);
and U33462 (N_33462,N_25035,N_23831);
nor U33463 (N_33463,N_26810,N_21602);
nor U33464 (N_33464,N_28547,N_25588);
or U33465 (N_33465,N_28306,N_25778);
or U33466 (N_33466,N_20530,N_26015);
or U33467 (N_33467,N_21439,N_29393);
nor U33468 (N_33468,N_27914,N_29652);
and U33469 (N_33469,N_27759,N_23379);
or U33470 (N_33470,N_21075,N_21516);
nor U33471 (N_33471,N_26044,N_22383);
nor U33472 (N_33472,N_29278,N_21386);
and U33473 (N_33473,N_24500,N_29433);
or U33474 (N_33474,N_27341,N_27195);
nand U33475 (N_33475,N_29749,N_29163);
xor U33476 (N_33476,N_23116,N_23570);
xnor U33477 (N_33477,N_28258,N_26801);
and U33478 (N_33478,N_21349,N_27830);
or U33479 (N_33479,N_23776,N_28228);
or U33480 (N_33480,N_26645,N_24421);
xnor U33481 (N_33481,N_22573,N_20922);
xor U33482 (N_33482,N_28091,N_26357);
or U33483 (N_33483,N_23397,N_26745);
and U33484 (N_33484,N_20364,N_26046);
or U33485 (N_33485,N_26696,N_26319);
xnor U33486 (N_33486,N_26901,N_22840);
nor U33487 (N_33487,N_21103,N_24032);
nor U33488 (N_33488,N_25977,N_24919);
xor U33489 (N_33489,N_28508,N_29423);
and U33490 (N_33490,N_20279,N_29810);
nand U33491 (N_33491,N_26700,N_29660);
nand U33492 (N_33492,N_20379,N_25938);
or U33493 (N_33493,N_26437,N_23810);
or U33494 (N_33494,N_21503,N_20464);
xor U33495 (N_33495,N_24482,N_26627);
or U33496 (N_33496,N_26414,N_20333);
nand U33497 (N_33497,N_24134,N_21953);
or U33498 (N_33498,N_20287,N_20593);
nor U33499 (N_33499,N_23389,N_27004);
nor U33500 (N_33500,N_29108,N_23056);
nor U33501 (N_33501,N_29939,N_22575);
and U33502 (N_33502,N_26002,N_27812);
and U33503 (N_33503,N_22175,N_24089);
and U33504 (N_33504,N_22427,N_27074);
nand U33505 (N_33505,N_29160,N_24308);
nor U33506 (N_33506,N_21049,N_20686);
xnor U33507 (N_33507,N_29470,N_26473);
xor U33508 (N_33508,N_25150,N_20026);
and U33509 (N_33509,N_21701,N_25216);
xor U33510 (N_33510,N_28643,N_25119);
or U33511 (N_33511,N_26866,N_24075);
nand U33512 (N_33512,N_25185,N_26001);
xnor U33513 (N_33513,N_23883,N_22455);
and U33514 (N_33514,N_24906,N_21609);
nor U33515 (N_33515,N_25573,N_26815);
or U33516 (N_33516,N_29194,N_29651);
nand U33517 (N_33517,N_20209,N_27444);
and U33518 (N_33518,N_20116,N_20200);
and U33519 (N_33519,N_21299,N_29237);
nand U33520 (N_33520,N_29255,N_22714);
xor U33521 (N_33521,N_26675,N_24810);
nor U33522 (N_33522,N_21429,N_28893);
and U33523 (N_33523,N_21055,N_27606);
nor U33524 (N_33524,N_29055,N_25470);
or U33525 (N_33525,N_20982,N_25230);
xnor U33526 (N_33526,N_25645,N_25813);
xnor U33527 (N_33527,N_21974,N_24762);
nor U33528 (N_33528,N_20764,N_28725);
xor U33529 (N_33529,N_22581,N_22792);
xnor U33530 (N_33530,N_22929,N_22365);
and U33531 (N_33531,N_28232,N_28606);
xor U33532 (N_33532,N_26388,N_21353);
and U33533 (N_33533,N_26100,N_24803);
and U33534 (N_33534,N_21284,N_29556);
nand U33535 (N_33535,N_28476,N_25384);
and U33536 (N_33536,N_26817,N_27396);
and U33537 (N_33537,N_21901,N_20154);
and U33538 (N_33538,N_23707,N_22800);
or U33539 (N_33539,N_26196,N_23904);
and U33540 (N_33540,N_23971,N_26780);
or U33541 (N_33541,N_29462,N_21617);
nand U33542 (N_33542,N_26837,N_25097);
or U33543 (N_33543,N_23362,N_29549);
or U33544 (N_33544,N_24632,N_22181);
and U33545 (N_33545,N_25000,N_28917);
or U33546 (N_33546,N_27377,N_22969);
xor U33547 (N_33547,N_22998,N_23121);
xor U33548 (N_33548,N_26027,N_28472);
and U33549 (N_33549,N_21866,N_20683);
or U33550 (N_33550,N_27463,N_28961);
xor U33551 (N_33551,N_29565,N_25918);
nor U33552 (N_33552,N_28834,N_22538);
and U33553 (N_33553,N_29545,N_27665);
nand U33554 (N_33554,N_21846,N_24530);
or U33555 (N_33555,N_29352,N_23205);
xor U33556 (N_33556,N_24957,N_27696);
xor U33557 (N_33557,N_24182,N_28005);
xnor U33558 (N_33558,N_27323,N_22206);
or U33559 (N_33559,N_27080,N_25542);
nand U33560 (N_33560,N_28044,N_20231);
and U33561 (N_33561,N_29247,N_25052);
and U33562 (N_33562,N_20274,N_29371);
xnor U33563 (N_33563,N_20396,N_20930);
or U33564 (N_33564,N_26565,N_26697);
or U33565 (N_33565,N_20335,N_26743);
nand U33566 (N_33566,N_29859,N_29181);
xnor U33567 (N_33567,N_25775,N_20143);
nor U33568 (N_33568,N_21174,N_22189);
or U33569 (N_33569,N_25005,N_26551);
xor U33570 (N_33570,N_28317,N_27613);
xor U33571 (N_33571,N_28760,N_20586);
nor U33572 (N_33572,N_28133,N_27514);
nand U33573 (N_33573,N_25564,N_28886);
or U33574 (N_33574,N_20422,N_27551);
or U33575 (N_33575,N_21427,N_27408);
xnor U33576 (N_33576,N_26207,N_23882);
nor U33577 (N_33577,N_26084,N_24439);
or U33578 (N_33578,N_22824,N_22235);
and U33579 (N_33579,N_23422,N_25638);
or U33580 (N_33580,N_24466,N_22701);
nand U33581 (N_33581,N_22609,N_29936);
xor U33582 (N_33582,N_28447,N_21361);
nor U33583 (N_33583,N_27066,N_27649);
nor U33584 (N_33584,N_22073,N_27678);
nand U33585 (N_33585,N_22731,N_29595);
and U33586 (N_33586,N_23910,N_22349);
nor U33587 (N_33587,N_26238,N_22265);
and U33588 (N_33588,N_29999,N_29880);
xnor U33589 (N_33589,N_21534,N_25129);
nand U33590 (N_33590,N_24764,N_21066);
xor U33591 (N_33591,N_25839,N_23675);
or U33592 (N_33592,N_28052,N_24222);
and U33593 (N_33593,N_28674,N_22977);
and U33594 (N_33594,N_29531,N_28970);
xnor U33595 (N_33595,N_21567,N_27032);
xnor U33596 (N_33596,N_22796,N_23053);
or U33597 (N_33597,N_25167,N_21015);
and U33598 (N_33598,N_22147,N_20575);
nor U33599 (N_33599,N_20752,N_27909);
nand U33600 (N_33600,N_26536,N_26423);
xnor U33601 (N_33601,N_25342,N_26193);
nor U33602 (N_33602,N_24236,N_27744);
and U33603 (N_33603,N_25080,N_29020);
or U33604 (N_33604,N_21959,N_28894);
xor U33605 (N_33605,N_22642,N_26882);
and U33606 (N_33606,N_27416,N_26264);
or U33607 (N_33607,N_26213,N_28000);
nand U33608 (N_33608,N_20461,N_21298);
nor U33609 (N_33609,N_28282,N_25335);
and U33610 (N_33610,N_21215,N_22112);
nor U33611 (N_33611,N_24832,N_20479);
xnor U33612 (N_33612,N_24185,N_26036);
and U33613 (N_33613,N_24928,N_24947);
or U33614 (N_33614,N_20939,N_26980);
and U33615 (N_33615,N_26140,N_24003);
and U33616 (N_33616,N_25268,N_22277);
nand U33617 (N_33617,N_25997,N_27995);
xnor U33618 (N_33618,N_27548,N_22370);
xor U33619 (N_33619,N_28273,N_27221);
nor U33620 (N_33620,N_22351,N_24733);
nand U33621 (N_33621,N_27330,N_23128);
nor U33622 (N_33622,N_28201,N_20328);
nand U33623 (N_33623,N_27310,N_23860);
nor U33624 (N_33624,N_23729,N_23466);
nand U33625 (N_33625,N_21411,N_25877);
or U33626 (N_33626,N_29528,N_28981);
nand U33627 (N_33627,N_26728,N_25032);
and U33628 (N_33628,N_22134,N_24430);
nand U33629 (N_33629,N_20673,N_24619);
or U33630 (N_33630,N_29742,N_21893);
nor U33631 (N_33631,N_26481,N_28039);
nand U33632 (N_33632,N_22530,N_25446);
and U33633 (N_33633,N_21205,N_23930);
xnor U33634 (N_33634,N_26498,N_21654);
nor U33635 (N_33635,N_26273,N_29447);
nor U33636 (N_33636,N_27210,N_24395);
nand U33637 (N_33637,N_22982,N_21640);
and U33638 (N_33638,N_20735,N_28623);
and U33639 (N_33639,N_25488,N_23275);
or U33640 (N_33640,N_25517,N_22681);
and U33641 (N_33641,N_21039,N_20161);
xor U33642 (N_33642,N_26055,N_26788);
nor U33643 (N_33643,N_22172,N_24926);
xor U33644 (N_33644,N_26534,N_22708);
xnor U33645 (N_33645,N_20111,N_29190);
and U33646 (N_33646,N_28330,N_22501);
and U33647 (N_33647,N_25780,N_20911);
or U33648 (N_33648,N_27631,N_29868);
xnor U33649 (N_33649,N_28406,N_23066);
and U33650 (N_33650,N_29404,N_27777);
xnor U33651 (N_33651,N_24918,N_21830);
and U33652 (N_33652,N_21775,N_21195);
and U33653 (N_33653,N_22990,N_20432);
nor U33654 (N_33654,N_28767,N_28721);
nand U33655 (N_33655,N_24446,N_28764);
nand U33656 (N_33656,N_24004,N_20824);
xor U33657 (N_33657,N_29629,N_27874);
and U33658 (N_33658,N_29250,N_24640);
nor U33659 (N_33659,N_22242,N_23190);
nand U33660 (N_33660,N_24998,N_28779);
nor U33661 (N_33661,N_26967,N_28938);
or U33662 (N_33662,N_28777,N_22053);
and U33663 (N_33663,N_24348,N_26545);
nor U33664 (N_33664,N_25594,N_23142);
nor U33665 (N_33665,N_24654,N_28927);
and U33666 (N_33666,N_29677,N_24577);
nor U33667 (N_33667,N_27435,N_23530);
nor U33668 (N_33668,N_25214,N_25557);
nor U33669 (N_33669,N_24216,N_22262);
or U33670 (N_33670,N_22475,N_21804);
nor U33671 (N_33671,N_23108,N_28367);
nor U33672 (N_33672,N_23573,N_25793);
nand U33673 (N_33673,N_24006,N_22484);
nor U33674 (N_33674,N_22497,N_21506);
nor U33675 (N_33675,N_27670,N_24853);
nor U33676 (N_33676,N_21320,N_22046);
or U33677 (N_33677,N_26632,N_23582);
xnor U33678 (N_33678,N_20934,N_26951);
nand U33679 (N_33679,N_24362,N_22806);
and U33680 (N_33680,N_26577,N_27434);
nand U33681 (N_33681,N_22843,N_23805);
xnor U33682 (N_33682,N_26992,N_25312);
xnor U33683 (N_33683,N_23609,N_29816);
or U33684 (N_33684,N_26169,N_25021);
or U33685 (N_33685,N_21333,N_27862);
or U33686 (N_33686,N_21403,N_24322);
nand U33687 (N_33687,N_29775,N_22273);
nor U33688 (N_33688,N_20721,N_20314);
and U33689 (N_33689,N_24775,N_22279);
nor U33690 (N_33690,N_21922,N_22255);
or U33691 (N_33691,N_25255,N_20980);
nor U33692 (N_33692,N_21753,N_20799);
and U33693 (N_33693,N_20125,N_28224);
xor U33694 (N_33694,N_29904,N_21621);
or U33695 (N_33695,N_27326,N_20525);
nand U33696 (N_33696,N_29533,N_25464);
nand U33697 (N_33697,N_27978,N_25871);
nor U33698 (N_33698,N_29002,N_29997);
nand U33699 (N_33699,N_22348,N_24620);
nand U33700 (N_33700,N_24330,N_21884);
or U33701 (N_33701,N_20663,N_22935);
or U33702 (N_33702,N_22782,N_23371);
or U33703 (N_33703,N_29398,N_20842);
or U33704 (N_33704,N_24505,N_23470);
nor U33705 (N_33705,N_26185,N_28741);
nor U33706 (N_33706,N_22444,N_26531);
nand U33707 (N_33707,N_20227,N_28515);
nand U33708 (N_33708,N_28202,N_20371);
xnor U33709 (N_33709,N_29431,N_26741);
and U33710 (N_33710,N_27667,N_23702);
nor U33711 (N_33711,N_29730,N_24508);
and U33712 (N_33712,N_24997,N_27785);
and U33713 (N_33713,N_20271,N_26154);
or U33714 (N_33714,N_20202,N_26848);
nand U33715 (N_33715,N_28250,N_22801);
nand U33716 (N_33716,N_22332,N_28684);
nand U33717 (N_33717,N_28851,N_22555);
xnor U33718 (N_33718,N_26735,N_29653);
xnor U33719 (N_33719,N_24648,N_21998);
xor U33720 (N_33720,N_23642,N_26105);
nor U33721 (N_33721,N_24826,N_22682);
or U33722 (N_33722,N_23252,N_24674);
xnor U33723 (N_33723,N_28996,N_22848);
nor U33724 (N_33724,N_28588,N_21186);
nor U33725 (N_33725,N_24682,N_20700);
and U33726 (N_33726,N_22948,N_21005);
nor U33727 (N_33727,N_25388,N_20289);
nor U33728 (N_33728,N_26333,N_20181);
nor U33729 (N_33729,N_28311,N_26775);
nand U33730 (N_33730,N_23918,N_27640);
or U33731 (N_33731,N_29292,N_25545);
or U33732 (N_33732,N_28431,N_26289);
and U33733 (N_33733,N_20629,N_27850);
nand U33734 (N_33734,N_25006,N_25452);
and U33735 (N_33735,N_22736,N_22852);
xnor U33736 (N_33736,N_26325,N_27146);
nor U33737 (N_33737,N_29921,N_29407);
and U33738 (N_33738,N_21911,N_20210);
xnor U33739 (N_33739,N_27764,N_24546);
and U33740 (N_33740,N_20996,N_24212);
xnor U33741 (N_33741,N_27163,N_20708);
nor U33742 (N_33742,N_28918,N_20446);
nor U33743 (N_33743,N_23581,N_28949);
and U33744 (N_33744,N_24880,N_25766);
and U33745 (N_33745,N_24259,N_27726);
xnor U33746 (N_33746,N_26957,N_29833);
or U33747 (N_33747,N_26204,N_23124);
nor U33748 (N_33748,N_29647,N_24027);
or U33749 (N_33749,N_28196,N_28669);
xnor U33750 (N_33750,N_21269,N_27834);
nand U33751 (N_33751,N_29225,N_25482);
nand U33752 (N_33752,N_22207,N_25122);
xor U33753 (N_33753,N_26990,N_26592);
xor U33754 (N_33754,N_25431,N_29608);
and U33755 (N_33755,N_23369,N_27710);
and U33756 (N_33756,N_25975,N_24326);
and U33757 (N_33757,N_26641,N_20600);
xnor U33758 (N_33758,N_22197,N_21370);
nor U33759 (N_33759,N_29983,N_24856);
and U33760 (N_33760,N_24181,N_26811);
xor U33761 (N_33761,N_22043,N_27031);
or U33762 (N_33762,N_26227,N_26113);
nand U33763 (N_33763,N_23980,N_21956);
or U33764 (N_33764,N_24636,N_23634);
xor U33765 (N_33765,N_28017,N_21527);
nor U33766 (N_33766,N_24442,N_22213);
nor U33767 (N_33767,N_20106,N_27798);
nand U33768 (N_33768,N_27720,N_24277);
xor U33769 (N_33769,N_20747,N_22812);
nor U33770 (N_33770,N_24267,N_21197);
xnor U33771 (N_33771,N_20462,N_24448);
nand U33772 (N_33772,N_29831,N_28048);
nor U33773 (N_33773,N_28189,N_22217);
or U33774 (N_33774,N_21108,N_23005);
xor U33775 (N_33775,N_27900,N_29972);
xor U33776 (N_33776,N_25233,N_28642);
nand U33777 (N_33777,N_25279,N_26655);
nand U33778 (N_33778,N_29481,N_29690);
nor U33779 (N_33779,N_25921,N_20837);
and U33780 (N_33780,N_22866,N_27118);
nand U33781 (N_33781,N_22504,N_24652);
nor U33782 (N_33782,N_23071,N_21622);
and U33783 (N_33783,N_27723,N_22176);
nor U33784 (N_33784,N_22345,N_24604);
nor U33785 (N_33785,N_23592,N_29051);
and U33786 (N_33786,N_22324,N_27621);
nand U33787 (N_33787,N_27935,N_20820);
nor U33788 (N_33788,N_21947,N_25736);
and U33789 (N_33789,N_24470,N_25273);
or U33790 (N_33790,N_27429,N_27912);
nand U33791 (N_33791,N_20960,N_23900);
nor U33792 (N_33792,N_25811,N_28186);
nor U33793 (N_33793,N_27865,N_25889);
xnor U33794 (N_33794,N_21368,N_26870);
nand U33795 (N_33795,N_21768,N_23475);
nand U33796 (N_33796,N_23265,N_21758);
nor U33797 (N_33797,N_27069,N_27288);
nor U33798 (N_33798,N_28126,N_26006);
nor U33799 (N_33799,N_21788,N_29332);
nand U33800 (N_33800,N_22913,N_28175);
and U33801 (N_33801,N_26867,N_25741);
and U33802 (N_33802,N_27747,N_22721);
nand U33803 (N_33803,N_28481,N_25135);
and U33804 (N_33804,N_22438,N_26194);
nand U33805 (N_33805,N_20612,N_28867);
nand U33806 (N_33806,N_27110,N_26180);
xor U33807 (N_33807,N_22250,N_23833);
nand U33808 (N_33808,N_24671,N_24849);
or U33809 (N_33809,N_25622,N_24074);
xnor U33810 (N_33810,N_29731,N_25582);
or U33811 (N_33811,N_26008,N_21178);
or U33812 (N_33812,N_26879,N_21825);
and U33813 (N_33813,N_23699,N_23493);
nor U33814 (N_33814,N_24916,N_23052);
or U33815 (N_33815,N_27021,N_25970);
nor U33816 (N_33816,N_20628,N_24987);
xnor U33817 (N_33817,N_22557,N_20698);
or U33818 (N_33818,N_20299,N_23916);
nand U33819 (N_33819,N_21829,N_26600);
or U33820 (N_33820,N_21556,N_25748);
xor U33821 (N_33821,N_22276,N_22056);
or U33822 (N_33822,N_27199,N_29949);
nand U33823 (N_33823,N_20585,N_27373);
xnor U33824 (N_33824,N_27966,N_20022);
or U33825 (N_33825,N_22600,N_24347);
nand U33826 (N_33826,N_27575,N_24168);
nor U33827 (N_33827,N_22333,N_21237);
and U33828 (N_33828,N_26942,N_21112);
xor U33829 (N_33829,N_24519,N_20829);
and U33830 (N_33830,N_23491,N_20284);
nand U33831 (N_33831,N_23527,N_21549);
nand U33832 (N_33832,N_25263,N_20054);
nand U33833 (N_33833,N_26317,N_28028);
and U33834 (N_33834,N_27779,N_23983);
or U33835 (N_33835,N_25776,N_23496);
xnor U33836 (N_33836,N_24161,N_20178);
xor U33837 (N_33837,N_28036,N_28833);
nand U33838 (N_33838,N_27181,N_27898);
or U33839 (N_33839,N_24235,N_26222);
or U33840 (N_33840,N_22472,N_27756);
and U33841 (N_33841,N_28400,N_20919);
or U33842 (N_33842,N_24496,N_25626);
xor U33843 (N_33843,N_26390,N_25994);
or U33844 (N_33844,N_23555,N_28103);
and U33845 (N_33845,N_22733,N_22565);
xnor U33846 (N_33846,N_29382,N_24821);
xnor U33847 (N_33847,N_27258,N_25296);
xor U33848 (N_33848,N_20412,N_28477);
and U33849 (N_33849,N_23280,N_25301);
xor U33850 (N_33850,N_26095,N_28896);
xor U33851 (N_33851,N_25141,N_21155);
xnor U33852 (N_33852,N_22858,N_24465);
nand U33853 (N_33853,N_29099,N_21986);
nor U33854 (N_33854,N_21193,N_20917);
xor U33855 (N_33855,N_24158,N_28423);
nand U33856 (N_33856,N_22462,N_26214);
or U33857 (N_33857,N_26275,N_21470);
or U33858 (N_33858,N_21152,N_26023);
nand U33859 (N_33859,N_23536,N_21297);
xnor U33860 (N_33860,N_23126,N_24662);
xnor U33861 (N_33861,N_20182,N_23004);
and U33862 (N_33862,N_26667,N_29946);
nand U33863 (N_33863,N_23091,N_28744);
nand U33864 (N_33864,N_25881,N_25095);
nand U33865 (N_33865,N_26327,N_28551);
nor U33866 (N_33866,N_22087,N_20108);
nor U33867 (N_33867,N_25876,N_21219);
and U33868 (N_33868,N_28747,N_26546);
xor U33869 (N_33869,N_27483,N_28647);
nand U33870 (N_33870,N_20510,N_23692);
or U33871 (N_33871,N_29453,N_20568);
nand U33872 (N_33872,N_25088,N_27132);
and U33873 (N_33873,N_23671,N_27088);
nor U33874 (N_33874,N_24705,N_22647);
nand U33875 (N_33875,N_26747,N_28782);
nand U33876 (N_33876,N_20789,N_24572);
nor U33877 (N_33877,N_23598,N_23786);
or U33878 (N_33878,N_23192,N_25271);
or U33879 (N_33879,N_26529,N_29772);
nand U33880 (N_33880,N_29865,N_22666);
nor U33881 (N_33881,N_23878,N_24289);
xnor U33882 (N_33882,N_23974,N_22363);
nand U33883 (N_33883,N_23917,N_22550);
xnor U33884 (N_33884,N_28098,N_20918);
or U33885 (N_33885,N_24576,N_24484);
xnor U33886 (N_33886,N_22396,N_20695);
or U33887 (N_33887,N_24769,N_20766);
nor U33888 (N_33888,N_22856,N_27886);
or U33889 (N_33889,N_22070,N_28971);
or U33890 (N_33890,N_24172,N_27411);
and U33891 (N_33891,N_25030,N_21792);
or U33892 (N_33892,N_27028,N_28719);
and U33893 (N_33893,N_21930,N_22480);
nor U33894 (N_33894,N_23081,N_26077);
and U33895 (N_33895,N_24180,N_26013);
and U33896 (N_33896,N_29867,N_29111);
nand U33897 (N_33897,N_29179,N_24143);
xnor U33898 (N_33898,N_24367,N_26247);
and U33899 (N_33899,N_22451,N_25664);
and U33900 (N_33900,N_29035,N_20807);
or U33901 (N_33901,N_27180,N_22078);
xor U33902 (N_33902,N_25500,N_23099);
nand U33903 (N_33903,N_26661,N_28880);
xor U33904 (N_33904,N_20770,N_23822);
nand U33905 (N_33905,N_28973,N_27147);
xor U33906 (N_33906,N_24757,N_25287);
and U33907 (N_33907,N_26628,N_27790);
or U33908 (N_33908,N_23541,N_23474);
xor U33909 (N_33909,N_24779,N_25533);
nand U33910 (N_33910,N_29667,N_23828);
nand U33911 (N_33911,N_20352,N_28522);
nand U33912 (N_33912,N_24073,N_26401);
xnor U33913 (N_33913,N_28380,N_29899);
or U33914 (N_33914,N_23245,N_22943);
xnor U33915 (N_33915,N_22042,N_27776);
or U33916 (N_33916,N_25044,N_22179);
xnor U33917 (N_33917,N_23838,N_28666);
nor U33918 (N_33918,N_21317,N_23424);
nor U33919 (N_33919,N_20475,N_20818);
nor U33920 (N_33920,N_27842,N_21528);
nand U33921 (N_33921,N_25568,N_20785);
and U33922 (N_33922,N_20189,N_28264);
xnor U33923 (N_33923,N_21659,N_21459);
and U33924 (N_33924,N_26230,N_26168);
and U33925 (N_33925,N_29778,N_26268);
nand U33926 (N_33926,N_26332,N_23322);
nor U33927 (N_33927,N_20163,N_25325);
xor U33928 (N_33928,N_29658,N_22698);
nand U33929 (N_33929,N_21286,N_25046);
xor U33930 (N_33930,N_28786,N_28857);
nand U33931 (N_33931,N_23516,N_29362);
nand U33932 (N_33932,N_23106,N_21343);
xnor U33933 (N_33933,N_27769,N_22028);
nor U33934 (N_33934,N_29622,N_29376);
xnor U33935 (N_33935,N_20074,N_22991);
nand U33936 (N_33936,N_20622,N_21441);
nand U33937 (N_33937,N_24474,N_21330);
or U33938 (N_33938,N_26654,N_20883);
nand U33939 (N_33939,N_21473,N_29563);
or U33940 (N_33940,N_25908,N_22304);
and U33941 (N_33941,N_28958,N_29033);
nand U33942 (N_33942,N_24706,N_28415);
and U33943 (N_33943,N_20767,N_29569);
or U33944 (N_33944,N_22984,N_29482);
and U33945 (N_33945,N_26460,N_27033);
nand U33946 (N_33946,N_21643,N_22689);
and U33947 (N_33947,N_22198,N_22030);
nand U33948 (N_33948,N_23812,N_27970);
or U33949 (N_33949,N_25102,N_20300);
nand U33950 (N_33950,N_25945,N_27792);
nand U33951 (N_33951,N_27220,N_29763);
nor U33952 (N_33952,N_24432,N_20050);
nor U33953 (N_33953,N_23870,N_20489);
xnor U33954 (N_33954,N_26086,N_26657);
or U33955 (N_33955,N_25251,N_22620);
and U33956 (N_33956,N_21241,N_20013);
nand U33957 (N_33957,N_24894,N_24587);
nor U33958 (N_33958,N_20579,N_27695);
nor U33959 (N_33959,N_25145,N_28245);
nor U33960 (N_33960,N_24425,N_24115);
nor U33961 (N_33961,N_27447,N_21770);
or U33962 (N_33962,N_24396,N_20418);
xor U33963 (N_33963,N_25815,N_20150);
and U33964 (N_33964,N_24225,N_27766);
nand U33965 (N_33965,N_26415,N_25380);
nand U33966 (N_33966,N_20817,N_21881);
nand U33967 (N_33967,N_26779,N_26176);
nand U33968 (N_33968,N_29413,N_29009);
and U33969 (N_33969,N_22158,N_23213);
xor U33970 (N_33970,N_26523,N_28096);
or U33971 (N_33971,N_28077,N_26192);
and U33972 (N_33972,N_26243,N_27692);
or U33973 (N_33973,N_21323,N_22032);
and U33974 (N_33974,N_25432,N_27246);
nor U33975 (N_33975,N_28555,N_26412);
and U33976 (N_33976,N_24693,N_24580);
and U33977 (N_33977,N_23759,N_28901);
nand U33978 (N_33978,N_23057,N_24678);
and U33979 (N_33979,N_28920,N_29014);
nand U33980 (N_33980,N_25570,N_28657);
or U33981 (N_33981,N_23197,N_26134);
nor U33982 (N_33982,N_25969,N_22168);
and U33983 (N_33983,N_26280,N_21221);
and U33984 (N_33984,N_26508,N_28456);
nand U33985 (N_33985,N_23069,N_28877);
nor U33986 (N_33986,N_28524,N_24067);
xor U33987 (N_33987,N_23902,N_26269);
or U33988 (N_33988,N_27570,N_29141);
nor U33989 (N_33989,N_25544,N_20419);
xnor U33990 (N_33990,N_28591,N_24627);
xnor U33991 (N_33991,N_20180,N_25666);
nor U33992 (N_33992,N_28587,N_22437);
nor U33993 (N_33993,N_25842,N_25779);
and U33994 (N_33994,N_22572,N_20197);
nor U33995 (N_33995,N_28615,N_21957);
or U33996 (N_33996,N_24400,N_29085);
and U33997 (N_33997,N_28923,N_28546);
nand U33998 (N_33998,N_22169,N_21447);
nand U33999 (N_33999,N_21688,N_29774);
and U34000 (N_34000,N_20958,N_23521);
and U34001 (N_34001,N_28468,N_20989);
nand U34002 (N_34002,N_28686,N_24175);
nand U34003 (N_34003,N_20472,N_28963);
nor U34004 (N_34004,N_22594,N_20326);
and U34005 (N_34005,N_21367,N_26731);
nor U34006 (N_34006,N_25867,N_28953);
or U34007 (N_34007,N_26789,N_21816);
and U34008 (N_34008,N_23853,N_22738);
xor U34009 (N_34009,N_21308,N_27144);
nor U34010 (N_34010,N_21645,N_22426);
or U34011 (N_34011,N_26679,N_25066);
nor U34012 (N_34012,N_22414,N_23955);
nand U34013 (N_34013,N_26041,N_21385);
nand U34014 (N_34014,N_25017,N_20604);
and U34015 (N_34015,N_25768,N_29344);
nand U34016 (N_34016,N_21100,N_29207);
or U34017 (N_34017,N_25696,N_23649);
and U34018 (N_34018,N_29335,N_20976);
nor U34019 (N_34019,N_24976,N_25579);
or U34020 (N_34020,N_29259,N_22068);
xnor U34021 (N_34021,N_25979,N_28821);
and U34022 (N_34022,N_25458,N_26603);
nand U34023 (N_34023,N_26255,N_26648);
nor U34024 (N_34024,N_24382,N_23616);
and U34025 (N_34025,N_28706,N_23460);
and U34026 (N_34026,N_20405,N_23710);
or U34027 (N_34027,N_21559,N_20476);
nand U34028 (N_34028,N_29267,N_21492);
xor U34029 (N_34029,N_26042,N_27017);
xnor U34030 (N_34030,N_27488,N_21794);
or U34031 (N_34031,N_26244,N_21671);
and U34032 (N_34032,N_29052,N_26233);
and U34033 (N_34033,N_20834,N_23139);
or U34034 (N_34034,N_29712,N_28235);
nand U34035 (N_34035,N_21627,N_25171);
nand U34036 (N_34036,N_21431,N_24283);
nand U34037 (N_34037,N_20223,N_25402);
or U34038 (N_34038,N_25476,N_21610);
nor U34039 (N_34039,N_27582,N_27869);
nor U34040 (N_34040,N_27456,N_21509);
or U34041 (N_34041,N_29623,N_24070);
xnor U34042 (N_34042,N_29437,N_26693);
or U34043 (N_34043,N_25356,N_26486);
xnor U34044 (N_34044,N_29171,N_27279);
nor U34045 (N_34045,N_29241,N_22723);
nor U34046 (N_34046,N_23670,N_29414);
nand U34047 (N_34047,N_25181,N_26017);
and U34048 (N_34048,N_28793,N_24865);
and U34049 (N_34049,N_21531,N_25788);
nor U34050 (N_34050,N_22135,N_20038);
nor U34051 (N_34051,N_20851,N_27479);
xnor U34052 (N_34052,N_24284,N_25624);
xor U34053 (N_34053,N_26672,N_20258);
nand U34054 (N_34054,N_27694,N_24111);
xnor U34055 (N_34055,N_26894,N_24291);
nand U34056 (N_34056,N_24319,N_20012);
xor U34057 (N_34057,N_27804,N_29443);
or U34058 (N_34058,N_29427,N_21719);
nor U34059 (N_34059,N_23413,N_29167);
xor U34060 (N_34060,N_25695,N_26143);
and U34061 (N_34061,N_23686,N_20073);
nand U34062 (N_34062,N_20080,N_24007);
nor U34063 (N_34063,N_29935,N_26245);
xnor U34064 (N_34064,N_21882,N_24353);
nor U34065 (N_34065,N_21340,N_20212);
nand U34066 (N_34066,N_24852,N_26714);
nor U34067 (N_34067,N_23083,N_22130);
and U34068 (N_34068,N_24827,N_20672);
nand U34069 (N_34069,N_24710,N_23224);
and U34070 (N_34070,N_27524,N_27539);
and U34071 (N_34071,N_23288,N_20020);
nand U34072 (N_34072,N_21632,N_21526);
nor U34073 (N_34073,N_24438,N_29377);
xnor U34074 (N_34074,N_23963,N_24068);
nand U34075 (N_34075,N_29635,N_23855);
and U34076 (N_34076,N_21540,N_23852);
nor U34077 (N_34077,N_20342,N_27327);
and U34078 (N_34078,N_25179,N_29429);
xor U34079 (N_34079,N_23258,N_20720);
xor U34080 (N_34080,N_27333,N_20520);
nand U34081 (N_34081,N_29977,N_25227);
nand U34082 (N_34082,N_21697,N_28602);
nor U34083 (N_34083,N_22432,N_29616);
nor U34084 (N_34084,N_29646,N_24105);
xor U34085 (N_34085,N_26869,N_29984);
or U34086 (N_34086,N_22900,N_28933);
or U34087 (N_34087,N_21201,N_24720);
and U34088 (N_34088,N_22166,N_22939);
or U34089 (N_34089,N_27268,N_20449);
xor U34090 (N_34090,N_27620,N_22301);
nand U34091 (N_34091,N_24647,N_20387);
and U34092 (N_34092,N_29397,N_24455);
nand U34093 (N_34093,N_27741,N_22204);
or U34094 (N_34094,N_27335,N_26718);
and U34095 (N_34095,N_24037,N_24771);
nand U34096 (N_34096,N_25370,N_24681);
nor U34097 (N_34097,N_21082,N_20002);
nor U34098 (N_34098,N_21649,N_23345);
and U34099 (N_34099,N_28620,N_25195);
and U34100 (N_34100,N_21133,N_20951);
nand U34101 (N_34101,N_21212,N_22603);
nand U34102 (N_34102,N_20653,N_20005);
nor U34103 (N_34103,N_27536,N_29885);
nand U34104 (N_34104,N_25567,N_28025);
xor U34105 (N_34105,N_29508,N_20392);
xor U34106 (N_34106,N_22997,N_21641);
or U34107 (N_34107,N_25838,N_26746);
and U34108 (N_34108,N_22248,N_27347);
xor U34109 (N_34109,N_29277,N_25463);
and U34110 (N_34110,N_23537,N_20843);
nor U34111 (N_34111,N_26744,N_29059);
and U34112 (N_34112,N_21300,N_20445);
nand U34113 (N_34113,N_21203,N_23514);
and U34114 (N_34114,N_26860,N_20055);
or U34115 (N_34115,N_21961,N_26108);
xor U34116 (N_34116,N_22013,N_20769);
nand U34117 (N_34117,N_27997,N_24155);
xor U34118 (N_34118,N_27406,N_29338);
or U34119 (N_34119,N_23407,N_20936);
and U34120 (N_34120,N_27894,N_25789);
xor U34121 (N_34121,N_21500,N_22612);
and U34122 (N_34122,N_28861,N_22994);
and U34123 (N_34123,N_24563,N_29625);
and U34124 (N_34124,N_27540,N_22010);
and U34125 (N_34125,N_20531,N_28829);
xnor U34126 (N_34126,N_20004,N_24847);
or U34127 (N_34127,N_25974,N_28743);
xnor U34128 (N_34128,N_29948,N_22347);
nor U34129 (N_34129,N_25022,N_24697);
nand U34130 (N_34130,N_24776,N_29581);
or U34131 (N_34131,N_22072,N_21393);
nor U34132 (N_34132,N_24592,N_29834);
nor U34133 (N_34133,N_22386,N_26982);
and U34134 (N_34134,N_25201,N_29848);
and U34135 (N_34135,N_24298,N_22428);
nor U34136 (N_34136,N_22429,N_28248);
or U34137 (N_34137,N_25647,N_24255);
nor U34138 (N_34138,N_20544,N_21686);
nand U34139 (N_34139,N_29136,N_25527);
and U34140 (N_34140,N_20356,N_29773);
xnor U34141 (N_34141,N_24083,N_20254);
nor U34142 (N_34142,N_23613,N_22703);
xor U34143 (N_34143,N_27693,N_24639);
xnor U34144 (N_34144,N_25723,N_27108);
nand U34145 (N_34145,N_28503,N_24501);
and U34146 (N_34146,N_28936,N_22745);
xnor U34147 (N_34147,N_27379,N_27151);
xor U34148 (N_34148,N_21328,N_24424);
nand U34149 (N_34149,N_27491,N_22892);
xor U34150 (N_34150,N_21126,N_22044);
and U34151 (N_34151,N_28172,N_21107);
and U34152 (N_34152,N_27000,N_29282);
nor U34153 (N_34153,N_21490,N_21267);
and U34154 (N_34154,N_24973,N_20733);
nand U34155 (N_34155,N_20844,N_21945);
and U34156 (N_34156,N_22951,N_23790);
or U34157 (N_34157,N_23196,N_29934);
and U34158 (N_34158,N_24152,N_26601);
nor U34159 (N_34159,N_22393,N_21890);
xnor U34160 (N_34160,N_26123,N_28297);
nand U34161 (N_34161,N_26380,N_27218);
nor U34162 (N_34162,N_25182,N_24937);
and U34163 (N_34163,N_23059,N_28398);
and U34164 (N_34164,N_27296,N_21554);
nor U34165 (N_34165,N_21864,N_26231);
nand U34166 (N_34166,N_20282,N_22041);
nor U34167 (N_34167,N_20694,N_24327);
nand U34168 (N_34168,N_29217,N_24407);
nand U34169 (N_34169,N_25763,N_25601);
nor U34170 (N_34170,N_24789,N_21469);
xnor U34171 (N_34171,N_25857,N_22551);
or U34172 (N_34172,N_27518,N_20118);
xnor U34173 (N_34173,N_25835,N_29286);
nor U34174 (N_34174,N_21928,N_20354);
or U34175 (N_34175,N_23779,N_21897);
and U34176 (N_34176,N_24629,N_22842);
nand U34177 (N_34177,N_20288,N_28058);
nor U34178 (N_34178,N_28828,N_25858);
xor U34179 (N_34179,N_27851,N_25199);
or U34180 (N_34180,N_26408,N_28835);
nor U34181 (N_34181,N_22826,N_28106);
xnor U34182 (N_34182,N_22503,N_29351);
or U34183 (N_34183,N_26032,N_22129);
nor U34184 (N_34184,N_26678,N_24246);
xnor U34185 (N_34185,N_29115,N_27148);
or U34186 (N_34186,N_29218,N_28698);
xor U34187 (N_34187,N_26876,N_27578);
nor U34188 (N_34188,N_23342,N_23307);
xor U34189 (N_34189,N_27372,N_28040);
xnor U34190 (N_34190,N_27068,N_26996);
nand U34191 (N_34191,N_21434,N_22122);
nand U34192 (N_34192,N_25852,N_25093);
or U34193 (N_34193,N_27300,N_29952);
nor U34194 (N_34194,N_23287,N_28514);
nor U34195 (N_34195,N_23448,N_21971);
nand U34196 (N_34196,N_23324,N_22146);
xor U34197 (N_34197,N_21292,N_20981);
or U34198 (N_34198,N_27975,N_28231);
nand U34199 (N_34199,N_21706,N_28335);
nor U34200 (N_34200,N_29769,N_25944);
and U34201 (N_34201,N_28053,N_21247);
and U34202 (N_34202,N_24528,N_20717);
and U34203 (N_34203,N_23970,N_21806);
nand U34204 (N_34204,N_29336,N_28026);
xnor U34205 (N_34205,N_21141,N_25260);
nand U34206 (N_34206,N_20185,N_24153);
and U34207 (N_34207,N_29666,N_28191);
xor U34208 (N_34208,N_24234,N_25929);
xor U34209 (N_34209,N_27770,N_23687);
nor U34210 (N_34210,N_28109,N_23191);
nor U34211 (N_34211,N_23425,N_20654);
and U34212 (N_34212,N_26443,N_26768);
xnor U34213 (N_34213,N_23557,N_22500);
nand U34214 (N_34214,N_22592,N_28383);
nand U34215 (N_34215,N_29023,N_21032);
nand U34216 (N_34216,N_26178,N_20776);
nand U34217 (N_34217,N_28302,N_26528);
nor U34218 (N_34218,N_27534,N_21636);
or U34219 (N_34219,N_24982,N_20750);
or U34220 (N_34220,N_28436,N_22152);
nor U34221 (N_34221,N_29504,N_28499);
nor U34222 (N_34222,N_22060,N_23109);
and U34223 (N_34223,N_26351,N_25825);
or U34224 (N_34224,N_27094,N_29535);
and U34225 (N_34225,N_25784,N_28660);
nand U34226 (N_34226,N_28523,N_25307);
or U34227 (N_34227,N_27915,N_27977);
nand U34228 (N_34228,N_28409,N_24634);
or U34229 (N_34229,N_21870,N_24591);
and U34230 (N_34230,N_29182,N_29134);
nand U34231 (N_34231,N_20448,N_26787);
xnor U34232 (N_34232,N_27499,N_24463);
nor U34233 (N_34233,N_27829,N_27887);
nand U34234 (N_34234,N_25660,N_27593);
nand U34235 (N_34235,N_26470,N_24211);
nor U34236 (N_34236,N_27820,N_24599);
or U34237 (N_34237,N_28758,N_22606);
nor U34238 (N_34238,N_29980,N_21694);
nand U34239 (N_34239,N_20224,N_29606);
xnor U34240 (N_34240,N_22377,N_23195);
nor U34241 (N_34241,N_25397,N_25607);
or U34242 (N_34242,N_23445,N_22164);
nand U34243 (N_34243,N_28651,N_25259);
xor U34244 (N_34244,N_26242,N_26410);
nand U34245 (N_34245,N_27588,N_23298);
or U34246 (N_34246,N_23597,N_25090);
nand U34247 (N_34247,N_22527,N_25834);
xor U34248 (N_34248,N_23285,N_28629);
nor U34249 (N_34249,N_29519,N_20347);
xnor U34250 (N_34250,N_23463,N_20630);
xnor U34251 (N_34251,N_26975,N_29374);
and U34252 (N_34252,N_26417,N_21883);
xnor U34253 (N_34253,N_24844,N_23588);
xor U34254 (N_34254,N_20734,N_25113);
xor U34255 (N_34255,N_29421,N_28804);
xnor U34256 (N_34256,N_28529,N_25697);
and U34257 (N_34257,N_21985,N_24962);
and U34258 (N_34258,N_29524,N_27664);
nor U34259 (N_34259,N_23524,N_22579);
nor U34260 (N_34260,N_23659,N_23050);
xnor U34261 (N_34261,N_26358,N_28343);
nor U34262 (N_34262,N_24066,N_28771);
or U34263 (N_34263,N_29757,N_28677);
and U34264 (N_34264,N_29940,N_29886);
xnor U34265 (N_34265,N_28598,N_23727);
or U34266 (N_34266,N_27298,N_21982);
xnor U34267 (N_34267,N_22253,N_23398);
nand U34268 (N_34268,N_22761,N_20906);
xnor U34269 (N_34269,N_24675,N_28065);
nand U34270 (N_34270,N_22372,N_29157);
and U34271 (N_34271,N_23620,N_22778);
or U34272 (N_34272,N_26285,N_23740);
xnor U34273 (N_34273,N_21374,N_27705);
nand U34274 (N_34274,N_24860,N_28216);
xor U34275 (N_34275,N_24313,N_28083);
xnor U34276 (N_34276,N_26228,N_22245);
and U34277 (N_34277,N_25225,N_27981);
nand U34278 (N_34278,N_20175,N_22239);
xnor U34279 (N_34279,N_24912,N_29346);
nor U34280 (N_34280,N_25875,N_29582);
nand U34281 (N_34281,N_25536,N_29572);
and U34282 (N_34282,N_27568,N_28609);
and U34283 (N_34283,N_20056,N_26463);
and U34284 (N_34284,N_23376,N_29319);
xnor U34285 (N_34285,N_20848,N_26056);
nand U34286 (N_34286,N_20759,N_28573);
and U34287 (N_34287,N_22412,N_22094);
nand U34288 (N_34288,N_20453,N_23994);
nand U34289 (N_34289,N_24874,N_20566);
xor U34290 (N_34290,N_23863,N_26335);
or U34291 (N_34291,N_25571,N_25966);
xor U34292 (N_34292,N_27857,N_25669);
and U34293 (N_34293,N_24258,N_25895);
nand U34294 (N_34294,N_20594,N_26379);
nand U34295 (N_34295,N_20651,N_25954);
and U34296 (N_34296,N_24848,N_24239);
or U34297 (N_34297,N_28500,N_24413);
nor U34298 (N_34298,N_26382,N_21225);
xnor U34299 (N_34299,N_27432,N_23674);
xor U34300 (N_34300,N_20646,N_25065);
or U34301 (N_34301,N_24370,N_22684);
and U34302 (N_34302,N_23896,N_27876);
nand U34303 (N_34303,N_21734,N_21898);
nand U34304 (N_34304,N_28321,N_20255);
xor U34305 (N_34305,N_28634,N_23841);
nand U34306 (N_34306,N_22891,N_27709);
and U34307 (N_34307,N_29813,N_27356);
nor U34308 (N_34308,N_28161,N_28622);
nor U34309 (N_34309,N_29594,N_27418);
nand U34310 (N_34310,N_28135,N_25295);
nor U34311 (N_34311,N_27893,N_26302);
xor U34312 (N_34312,N_25625,N_25337);
xor U34313 (N_34313,N_26582,N_26458);
or U34314 (N_34314,N_29261,N_27512);
or U34315 (N_34315,N_27567,N_23063);
or U34316 (N_34316,N_28944,N_29796);
xnor U34317 (N_34317,N_22546,N_27485);
and U34318 (N_34318,N_23337,N_24374);
or U34319 (N_34319,N_20138,N_24868);
and U34320 (N_34320,N_28858,N_25801);
or U34321 (N_34321,N_24233,N_29366);
nor U34322 (N_34322,N_24408,N_23001);
nand U34323 (N_34323,N_23012,N_23595);
nor U34324 (N_34324,N_29520,N_23024);
nand U34325 (N_34325,N_24336,N_26110);
and U34326 (N_34326,N_20731,N_25126);
nor U34327 (N_34327,N_29539,N_24651);
or U34328 (N_34328,N_24262,N_27340);
nand U34329 (N_34329,N_23411,N_24189);
nand U34330 (N_34330,N_21865,N_22029);
xor U34331 (N_34331,N_26767,N_28054);
nor U34332 (N_34332,N_26256,N_27553);
xor U34333 (N_34333,N_28710,N_27782);
xor U34334 (N_34334,N_27065,N_24281);
or U34335 (N_34335,N_26993,N_27230);
nand U34336 (N_34336,N_23506,N_23073);
and U34337 (N_34337,N_24814,N_26919);
and U34338 (N_34338,N_26615,N_20256);
or U34339 (N_34339,N_28181,N_21425);
xnor U34340 (N_34340,N_29924,N_28694);
or U34341 (N_34341,N_24191,N_27473);
and U34342 (N_34342,N_25808,N_26955);
xnor U34343 (N_34343,N_21779,N_23264);
nand U34344 (N_34344,N_24709,N_24552);
xor U34345 (N_34345,N_23711,N_24013);
xnor U34346 (N_34346,N_22395,N_23420);
xor U34347 (N_34347,N_25155,N_29176);
xnor U34348 (N_34348,N_22809,N_29752);
xor U34349 (N_34349,N_28070,N_25888);
xor U34350 (N_34350,N_28639,N_20147);
nor U34351 (N_34351,N_29079,N_24835);
xnor U34352 (N_34352,N_27481,N_26396);
xnor U34353 (N_34353,N_20390,N_22884);
nand U34354 (N_34354,N_26656,N_24967);
xnor U34355 (N_34355,N_29687,N_24729);
nor U34356 (N_34356,N_27425,N_25892);
nand U34357 (N_34357,N_23331,N_24194);
or U34358 (N_34358,N_23789,N_22827);
nor U34359 (N_34359,N_21577,N_21378);
and U34360 (N_34360,N_20662,N_28860);
nand U34361 (N_34361,N_29797,N_23750);
nand U34362 (N_34362,N_21927,N_29235);
xnor U34363 (N_34363,N_20772,N_20887);
xor U34364 (N_34364,N_23919,N_26034);
or U34365 (N_34365,N_20094,N_23837);
and U34366 (N_34366,N_22552,N_22232);
xor U34367 (N_34367,N_23552,N_22741);
or U34368 (N_34368,N_22979,N_25694);
xnor U34369 (N_34369,N_22040,N_20743);
and U34370 (N_34370,N_26559,N_21023);
xnor U34371 (N_34371,N_28671,N_22002);
nand U34372 (N_34372,N_24261,N_25764);
or U34373 (N_34373,N_27097,N_26240);
and U34374 (N_34374,N_21904,N_29493);
nand U34375 (N_34375,N_23879,N_24354);
and U34376 (N_34376,N_28992,N_27056);
xnor U34377 (N_34377,N_25559,N_28099);
nor U34378 (N_34378,N_22716,N_24209);
nor U34379 (N_34379,N_24352,N_25535);
xnor U34380 (N_34380,N_24220,N_23651);
xor U34381 (N_34381,N_22902,N_20727);
and U34382 (N_34382,N_23401,N_29703);
xnor U34383 (N_34383,N_26012,N_24350);
or U34384 (N_34384,N_25972,N_24672);
or U34385 (N_34385,N_21553,N_26237);
nor U34386 (N_34386,N_28892,N_23087);
nor U34387 (N_34387,N_24804,N_24784);
and U34388 (N_34388,N_21925,N_25754);
or U34389 (N_34389,N_25821,N_20647);
or U34390 (N_34390,N_22343,N_20443);
or U34391 (N_34391,N_27661,N_21662);
xor U34392 (N_34392,N_27465,N_20451);
nand U34393 (N_34393,N_26691,N_28139);
xor U34394 (N_34394,N_23715,N_23965);
and U34395 (N_34395,N_28885,N_23380);
nor U34396 (N_34396,N_26476,N_28675);
xnor U34397 (N_34397,N_21487,N_20045);
or U34398 (N_34398,N_27803,N_24052);
nor U34399 (N_34399,N_27702,N_26104);
or U34400 (N_34400,N_22511,N_20318);
nand U34401 (N_34401,N_24084,N_23987);
nor U34402 (N_34402,N_26591,N_25019);
and U34403 (N_34403,N_24999,N_23783);
and U34404 (N_34404,N_26532,N_26054);
nor U34405 (N_34405,N_29011,N_26266);
nor U34406 (N_34406,N_21683,N_23950);
nor U34407 (N_34407,N_21206,N_23256);
and U34408 (N_34408,N_21740,N_26037);
xor U34409 (N_34409,N_21048,N_28837);
and U34410 (N_34410,N_22691,N_29199);
xor U34411 (N_34411,N_28280,N_26483);
nand U34412 (N_34412,N_24743,N_29345);
and U34413 (N_34413,N_28664,N_26491);
or U34414 (N_34414,N_20165,N_29152);
and U34415 (N_34415,N_20808,N_29340);
nand U34416 (N_34416,N_29435,N_25787);
nor U34417 (N_34417,N_27679,N_23525);
or U34418 (N_34418,N_29928,N_21847);
xor U34419 (N_34419,N_28940,N_26326);
and U34420 (N_34420,N_20712,N_23312);
or U34421 (N_34421,N_26585,N_27791);
and U34422 (N_34422,N_21943,N_28848);
xnor U34423 (N_34423,N_20526,N_23761);
and U34424 (N_34424,N_29628,N_20649);
and U34425 (N_34425,N_23414,N_23768);
and U34426 (N_34426,N_25086,N_22617);
xnor U34427 (N_34427,N_22238,N_21257);
or U34428 (N_34428,N_20786,N_20885);
or U34429 (N_34429,N_28374,N_27175);
and U34430 (N_34430,N_22926,N_28461);
and U34431 (N_34431,N_27219,N_26619);
nand U34432 (N_34432,N_28871,N_27206);
or U34433 (N_34433,N_24020,N_25002);
nor U34434 (N_34434,N_22160,N_25114);
or U34435 (N_34435,N_20430,N_24742);
xnor U34436 (N_34436,N_28882,N_22300);
or U34437 (N_34437,N_29824,N_23999);
nor U34438 (N_34438,N_22596,N_24128);
and U34439 (N_34439,N_29412,N_23523);
and U34440 (N_34440,N_24543,N_20156);
nor U34441 (N_34441,N_27543,N_25288);
and U34442 (N_34442,N_28362,N_28796);
or U34443 (N_34443,N_24964,N_27837);
xnor U34444 (N_34444,N_23600,N_23658);
and U34445 (N_34445,N_21187,N_23681);
or U34446 (N_34446,N_26038,N_23774);
nor U34447 (N_34447,N_22829,N_28673);
nand U34448 (N_34448,N_24968,N_23526);
nand U34449 (N_34449,N_22368,N_22212);
or U34450 (N_34450,N_21086,N_20741);
nand U34451 (N_34451,N_24204,N_20179);
xor U34452 (N_34452,N_29766,N_29890);
and U34453 (N_34453,N_28788,N_22471);
nand U34454 (N_34454,N_20779,N_25992);
xnor U34455 (N_34455,N_20729,N_26650);
xnor U34456 (N_34456,N_26059,N_27193);
and U34457 (N_34457,N_22541,N_25149);
nand U34458 (N_34458,N_26677,N_23111);
and U34459 (N_34459,N_20705,N_27067);
and U34460 (N_34460,N_27930,N_29039);
nand U34461 (N_34461,N_21388,N_29958);
xor U34462 (N_34462,N_27227,N_23682);
or U34463 (N_34463,N_25121,N_24704);
nor U34464 (N_34464,N_29276,N_28792);
and U34465 (N_34465,N_25738,N_26988);
nand U34466 (N_34466,N_24426,N_28171);
and U34467 (N_34467,N_28194,N_29402);
nor U34468 (N_34468,N_26119,N_23250);
nand U34469 (N_34469,N_21140,N_29100);
or U34470 (N_34470,N_20308,N_28459);
or U34471 (N_34471,N_27072,N_28822);
nand U34472 (N_34472,N_28596,N_27158);
nor U34473 (N_34473,N_21713,N_28200);
nor U34474 (N_34474,N_22344,N_25223);
nor U34475 (N_34475,N_21397,N_28192);
or U34476 (N_34476,N_26690,N_27169);
and U34477 (N_34477,N_28662,N_21485);
and U34478 (N_34478,N_24035,N_27117);
nand U34479 (N_34479,N_23378,N_29468);
xor U34480 (N_34480,N_25198,N_25367);
xnor U34481 (N_34481,N_22154,N_27278);
and U34482 (N_34482,N_22331,N_24645);
nor U34483 (N_34483,N_28425,N_20553);
or U34484 (N_34484,N_24431,N_21009);
or U34485 (N_34485,N_21040,N_24321);
or U34486 (N_34486,N_23134,N_23899);
nor U34487 (N_34487,N_25617,N_23044);
or U34488 (N_34488,N_20506,N_25128);
and U34489 (N_34489,N_24569,N_22639);
and U34490 (N_34490,N_22862,N_24445);
xor U34491 (N_34491,N_23844,N_20234);
nand U34492 (N_34492,N_26948,N_27006);
nand U34493 (N_34493,N_25357,N_28197);
and U34494 (N_34494,N_20806,N_22886);
nor U34495 (N_34495,N_27873,N_27611);
xor U34496 (N_34496,N_29016,N_22019);
nor U34497 (N_34497,N_26885,N_20329);
or U34498 (N_34498,N_24980,N_21915);
nor U34499 (N_34499,N_23632,N_28180);
nor U34500 (N_34500,N_21652,N_27510);
nor U34501 (N_34501,N_24825,N_20428);
xor U34502 (N_34502,N_28799,N_27187);
and U34503 (N_34503,N_23323,N_25278);
or U34504 (N_34504,N_29378,N_24085);
or U34505 (N_34505,N_24098,N_23068);
nand U34506 (N_34506,N_23332,N_20923);
xor U34507 (N_34507,N_29969,N_24385);
nand U34508 (N_34508,N_27663,N_27495);
nand U34509 (N_34509,N_23922,N_21657);
xnor U34510 (N_34510,N_20082,N_29289);
nand U34511 (N_34511,N_20962,N_23135);
xor U34512 (N_34512,N_22458,N_29312);
xnor U34513 (N_34513,N_21499,N_25429);
nor U34514 (N_34514,N_25084,N_26742);
nor U34515 (N_34515,N_24694,N_22320);
nor U34516 (N_34516,N_24471,N_26000);
xnor U34517 (N_34517,N_29897,N_23771);
xor U34518 (N_34518,N_28243,N_23969);
and U34519 (N_34519,N_27128,N_20398);
and U34520 (N_34520,N_29602,N_23639);
and U34521 (N_34521,N_20610,N_22759);
or U34522 (N_34522,N_23920,N_21390);
nand U34523 (N_34523,N_25646,N_25502);
or U34524 (N_34524,N_23341,N_23684);
nor U34525 (N_34525,N_25443,N_22767);
or U34526 (N_34526,N_25549,N_28966);
nand U34527 (N_34527,N_29988,N_27244);
nor U34528 (N_34528,N_21532,N_23906);
nor U34529 (N_34529,N_20605,N_24171);
or U34530 (N_34530,N_26313,N_28580);
nor U34531 (N_34531,N_24486,N_26208);
nor U34532 (N_34532,N_20956,N_26480);
or U34533 (N_34533,N_20762,N_21835);
nor U34534 (N_34534,N_29501,N_23185);
and U34535 (N_34535,N_25756,N_25585);
nand U34536 (N_34536,N_24673,N_21508);
nand U34537 (N_34537,N_24698,N_20990);
or U34538 (N_34538,N_22793,N_24010);
or U34539 (N_34539,N_21158,N_22588);
xnor U34540 (N_34540,N_23803,N_27005);
and U34541 (N_34541,N_20291,N_21564);
or U34542 (N_34542,N_29951,N_28092);
nor U34543 (N_34543,N_26221,N_26188);
xnor U34544 (N_34544,N_24388,N_21144);
nor U34545 (N_34545,N_20172,N_29938);
and U34546 (N_34546,N_20823,N_29954);
xor U34547 (N_34547,N_28304,N_29126);
nor U34548 (N_34548,N_26623,N_28141);
xor U34549 (N_34549,N_24890,N_23615);
xnor U34550 (N_34550,N_24357,N_22857);
nand U34551 (N_34551,N_20023,N_20385);
xnor U34552 (N_34552,N_25924,N_28990);
and U34553 (N_34553,N_29187,N_21303);
nor U34554 (N_34554,N_21979,N_26103);
xor U34555 (N_34555,N_29348,N_20543);
xor U34556 (N_34556,N_22795,N_22915);
or U34557 (N_34557,N_29753,N_26471);
xnor U34558 (N_34558,N_21474,N_23228);
nand U34559 (N_34559,N_26122,N_24902);
or U34560 (N_34560,N_26574,N_22439);
nor U34561 (N_34561,N_20293,N_20595);
or U34562 (N_34562,N_29215,N_28408);
and U34563 (N_34563,N_25242,N_25673);
xnor U34564 (N_34564,N_23809,N_26999);
nor U34565 (N_34565,N_26236,N_22513);
or U34566 (N_34566,N_24492,N_21010);
and U34567 (N_34567,N_28769,N_23884);
or U34568 (N_34568,N_25781,N_20036);
and U34569 (N_34569,N_21765,N_28385);
and U34570 (N_34570,N_28485,N_28730);
nand U34571 (N_34571,N_29496,N_23807);
nand U34572 (N_34572,N_26969,N_20331);
nand U34573 (N_34573,N_23168,N_23895);
nand U34574 (N_34574,N_21566,N_21992);
and U34575 (N_34575,N_23545,N_21744);
and U34576 (N_34576,N_25234,N_26112);
and U34577 (N_34577,N_24934,N_29130);
nand U34578 (N_34578,N_23751,N_21840);
nor U34579 (N_34579,N_22150,N_22828);
and U34580 (N_34580,N_26542,N_27967);
nand U34581 (N_34581,N_21628,N_21917);
or U34582 (N_34582,N_26191,N_26524);
xnor U34583 (N_34583,N_25745,N_24295);
nand U34584 (N_34584,N_28445,N_25332);
xnor U34585 (N_34585,N_29301,N_23663);
xor U34586 (N_34586,N_22443,N_29957);
xnor U34587 (N_34587,N_29192,N_27399);
or U34588 (N_34588,N_23030,N_28298);
nand U34589 (N_34589,N_28676,N_28540);
and U34590 (N_34590,N_22491,N_28279);
or U34591 (N_34591,N_22818,N_20793);
xnor U34592 (N_34592,N_22641,N_20607);
and U34593 (N_34593,N_28717,N_25985);
or U34594 (N_34594,N_22955,N_27991);
nand U34595 (N_34595,N_21544,N_20899);
or U34596 (N_34596,N_28632,N_20429);
nor U34597 (N_34597,N_28490,N_26908);
xnor U34598 (N_34598,N_25744,N_25983);
xnor U34599 (N_34599,N_28045,N_29196);
nand U34600 (N_34600,N_23636,N_24099);
nand U34601 (N_34601,N_20494,N_25800);
xor U34602 (N_34602,N_20363,N_22646);
or U34603 (N_34603,N_21147,N_28122);
nand U34604 (N_34604,N_27737,N_27297);
or U34605 (N_34605,N_28124,N_29862);
or U34606 (N_34606,N_26639,N_21069);
nand U34607 (N_34607,N_29905,N_29391);
and U34608 (N_34608,N_24323,N_23286);
xnor U34609 (N_34609,N_28494,N_25320);
or U34610 (N_34610,N_20571,N_21538);
nand U34611 (N_34611,N_28947,N_29990);
and U34612 (N_34612,N_22419,N_27249);
and U34613 (N_34613,N_24603,N_20241);
and U34614 (N_34614,N_21525,N_26598);
nand U34615 (N_34615,N_27371,N_26991);
xor U34616 (N_34616,N_20034,N_20015);
and U34617 (N_34617,N_24995,N_27772);
and U34618 (N_34618,N_23665,N_22183);
or U34619 (N_34619,N_25851,N_22111);
or U34620 (N_34620,N_29729,N_26070);
or U34621 (N_34621,N_21802,N_20499);
xor U34622 (N_34622,N_20344,N_25277);
xor U34623 (N_34623,N_27916,N_22167);
nand U34624 (N_34624,N_29603,N_23767);
nand U34625 (N_34625,N_20149,N_20944);
nand U34626 (N_34626,N_20674,N_27104);
nand U34627 (N_34627,N_22143,N_24154);
nor U34628 (N_34628,N_26340,N_22713);
xor U34629 (N_34629,N_22190,N_26263);
or U34630 (N_34630,N_25580,N_22911);
nor U34631 (N_34631,N_25116,N_21639);
nor U34632 (N_34632,N_29222,N_26830);
or U34633 (N_34633,N_21356,N_22834);
and U34634 (N_34634,N_21240,N_24831);
or U34635 (N_34635,N_21332,N_20615);
and U34636 (N_34636,N_25435,N_28755);
nor U34637 (N_34637,N_27314,N_21295);
nand U34638 (N_34638,N_27963,N_25651);
nor U34639 (N_34639,N_28142,N_29583);
or U34640 (N_34640,N_23656,N_23721);
or U34641 (N_34641,N_28305,N_25755);
nor U34642 (N_34642,N_27630,N_28361);
xor U34643 (N_34643,N_20072,N_23148);
nand U34644 (N_34644,N_23512,N_25530);
and U34645 (N_34645,N_21660,N_28733);
and U34646 (N_34646,N_21314,N_22360);
and U34647 (N_34647,N_20133,N_20345);
nand U34648 (N_34648,N_21159,N_27076);
nand U34649 (N_34649,N_20562,N_29847);
nor U34650 (N_34650,N_27781,N_27609);
nand U34651 (N_34651,N_24104,N_28750);
or U34652 (N_34652,N_27602,N_27285);
nor U34653 (N_34653,N_24351,N_28007);
xnor U34654 (N_34654,N_29156,N_23494);
and U34655 (N_34655,N_26444,N_21443);
or U34656 (N_34656,N_23247,N_23370);
nand U34657 (N_34657,N_28825,N_28875);
xor U34658 (N_34658,N_26541,N_29036);
and U34659 (N_34659,N_25003,N_24549);
or U34660 (N_34660,N_20275,N_25608);
and U34661 (N_34661,N_29697,N_28220);
xor U34662 (N_34662,N_27496,N_26150);
or U34663 (N_34663,N_24038,N_23304);
nand U34664 (N_34664,N_27958,N_20246);
nor U34665 (N_34665,N_20467,N_28486);
and U34666 (N_34666,N_26777,N_26839);
or U34667 (N_34667,N_22312,N_29457);
xor U34668 (N_34668,N_25410,N_26886);
nor U34669 (N_34669,N_21939,N_24518);
nand U34670 (N_34670,N_23590,N_21063);
xor U34671 (N_34671,N_22498,N_26636);
nand U34672 (N_34672,N_20140,N_22337);
and U34673 (N_34673,N_29358,N_28910);
and U34674 (N_34674,N_20157,N_23394);
nor U34675 (N_34675,N_28843,N_28768);
and U34676 (N_34676,N_23538,N_26799);
and U34677 (N_34677,N_24676,N_25207);
nor U34678 (N_34678,N_29313,N_23316);
nor U34679 (N_34679,N_21656,N_24359);
nor U34680 (N_34680,N_27508,N_29383);
nor U34681 (N_34681,N_25346,N_29682);
xor U34682 (N_34682,N_20033,N_22215);
xor U34683 (N_34683,N_21774,N_21687);
nor U34684 (N_34684,N_23299,N_24981);
nand U34685 (N_34685,N_21007,N_27614);
xor U34686 (N_34686,N_26748,N_28713);
nor U34687 (N_34687,N_24050,N_27926);
nor U34688 (N_34688,N_28144,N_27608);
or U34689 (N_34689,N_23017,N_20688);
or U34690 (N_34690,N_26097,N_21101);
or U34691 (N_34691,N_28761,N_28688);
or U34692 (N_34692,N_24780,N_24360);
or U34693 (N_34693,N_21848,N_23319);
and U34694 (N_34694,N_27093,N_23653);
nand U34695 (N_34695,N_21766,N_23015);
or U34696 (N_34696,N_20088,N_28913);
nor U34697 (N_34697,N_26915,N_23339);
xor U34698 (N_34698,N_23318,N_22247);
nand U34699 (N_34699,N_27233,N_20664);
xor U34700 (N_34700,N_22838,N_26199);
or U34701 (N_34701,N_23079,N_25120);
nor U34702 (N_34702,N_23944,N_26232);
nand U34703 (N_34703,N_27451,N_20803);
xor U34704 (N_34704,N_28908,N_20955);
and U34705 (N_34705,N_25725,N_23014);
xnor U34706 (N_34706,N_23587,N_29070);
nor U34707 (N_34707,N_23119,N_24493);
and U34708 (N_34708,N_21778,N_29145);
and U34709 (N_34709,N_28610,N_26852);
nand U34710 (N_34710,N_29188,N_22191);
nor U34711 (N_34711,N_24782,N_20260);
and U34712 (N_34712,N_24798,N_22766);
and U34713 (N_34713,N_24103,N_24082);
xor U34714 (N_34714,N_28537,N_25677);
xnor U34715 (N_34715,N_25403,N_29807);
nor U34716 (N_34716,N_25670,N_25782);
nor U34717 (N_34717,N_24805,N_27459);
or U34718 (N_34718,N_25249,N_26643);
xnor U34719 (N_34719,N_28068,N_23038);
xor U34720 (N_34720,N_26016,N_23938);
or U34721 (N_34721,N_28683,N_27773);
and U34722 (N_34722,N_26405,N_21394);
xor U34723 (N_34723,N_29571,N_25612);
nand U34724 (N_34724,N_27077,N_21275);
nor U34725 (N_34725,N_24169,N_24029);
xnor U34726 (N_34726,N_27521,N_20908);
or U34727 (N_34727,N_26211,N_28088);
or U34728 (N_34728,N_27585,N_29452);
nor U34729 (N_34729,N_26094,N_27498);
and U34730 (N_34730,N_27574,N_20821);
or U34731 (N_34731,N_24792,N_24201);
xor U34732 (N_34732,N_26368,N_24183);
xnor U34733 (N_34733,N_22149,N_27375);
nand U34734 (N_34734,N_28392,N_28942);
xnor U34735 (N_34735,N_26671,N_29804);
nand U34736 (N_34736,N_25217,N_21008);
nand U34737 (N_34737,N_22544,N_29656);
or U34738 (N_34738,N_22234,N_24588);
nand U34739 (N_34739,N_24030,N_26539);
and U34740 (N_34740,N_21065,N_29499);
xnor U34741 (N_34741,N_26381,N_28182);
xor U34742 (N_34742,N_26840,N_24978);
nand U34743 (N_34743,N_26843,N_27919);
nor U34744 (N_34744,N_24346,N_23743);
xnor U34745 (N_34745,N_29664,N_29385);
or U34746 (N_34746,N_23680,N_29516);
and U34747 (N_34747,N_24127,N_20521);
xnor U34748 (N_34748,N_26488,N_26977);
nor U34749 (N_34749,N_29802,N_26865);
nand U34750 (N_34750,N_24199,N_29598);
nor U34751 (N_34751,N_22192,N_21693);
or U34752 (N_34752,N_26708,N_27658);
nor U34753 (N_34753,N_26575,N_25180);
nand U34754 (N_34754,N_22108,N_22515);
nor U34755 (N_34755,N_20370,N_29490);
xnor U34756 (N_34756,N_26030,N_29790);
nand U34757 (N_34757,N_26664,N_25393);
and U34758 (N_34758,N_27503,N_26753);
xnor U34759 (N_34759,N_22006,N_28087);
nor U34760 (N_34760,N_25254,N_28791);
xnor U34761 (N_34761,N_22868,N_28831);
nor U34762 (N_34762,N_27316,N_20267);
xor U34763 (N_34763,N_28986,N_29053);
and U34764 (N_34764,N_27866,N_28021);
xnor U34765 (N_34765,N_22952,N_27392);
nand U34766 (N_34766,N_24335,N_29568);
nor U34767 (N_34767,N_25132,N_26762);
xnor U34768 (N_34768,N_26938,N_27871);
nor U34769 (N_34769,N_25652,N_21818);
xor U34770 (N_34770,N_22922,N_28424);
nor U34771 (N_34771,N_21722,N_25326);
nor U34772 (N_34772,N_20988,N_28919);
nand U34773 (N_34773,N_28984,N_21271);
nor U34774 (N_34774,N_21190,N_20855);
or U34775 (N_34775,N_20592,N_23078);
and U34776 (N_34776,N_26052,N_28785);
and U34777 (N_34777,N_26422,N_27870);
and U34778 (N_34778,N_25655,N_20330);
or U34779 (N_34779,N_24269,N_27307);
or U34780 (N_34780,N_22308,N_24747);
and U34781 (N_34781,N_25423,N_24956);
xor U34782 (N_34782,N_28307,N_28414);
xnor U34783 (N_34783,N_25162,N_20563);
xor U34784 (N_34784,N_23580,N_27207);
nand U34785 (N_34785,N_28898,N_25372);
and U34786 (N_34786,N_26861,N_25896);
nand U34787 (N_34787,N_25891,N_22656);
and U34788 (N_34788,N_28166,N_20391);
nand U34789 (N_34789,N_29788,N_23476);
nor U34790 (N_34790,N_22586,N_27200);
or U34791 (N_34791,N_24531,N_29475);
nand U34792 (N_34792,N_22722,N_22871);
nand U34793 (N_34793,N_23254,N_25925);
and U34794 (N_34794,N_29212,N_28418);
and U34795 (N_34795,N_22003,N_22933);
and U34796 (N_34796,N_23559,N_24581);
nor U34797 (N_34797,N_25773,N_28388);
or U34798 (N_34798,N_27727,N_24927);
and U34799 (N_34799,N_28214,N_29709);
or U34800 (N_34800,N_24263,N_21646);
and U34801 (N_34801,N_25905,N_27243);
xnor U34802 (N_34802,N_22699,N_20938);
nand U34803 (N_34803,N_29574,N_23393);
or U34804 (N_34804,N_21535,N_26979);
and U34805 (N_34805,N_21764,N_23881);
or U34806 (N_34806,N_22449,N_23714);
and U34807 (N_34807,N_28535,N_24756);
or U34808 (N_34808,N_28922,N_23712);
nor U34809 (N_34809,N_20253,N_27259);
and U34810 (N_34810,N_29750,N_28111);
nand U34811 (N_34811,N_27808,N_29257);
or U34812 (N_34812,N_23348,N_24839);
and U34813 (N_34813,N_24095,N_23206);
xor U34814 (N_34814,N_21669,N_22413);
nand U34815 (N_34815,N_29297,N_26058);
nand U34816 (N_34816,N_29761,N_26009);
xnor U34817 (N_34817,N_23201,N_24033);
nor U34818 (N_34818,N_25880,N_28571);
nor U34819 (N_34819,N_20978,N_22571);
nand U34820 (N_34820,N_26694,N_23606);
nor U34821 (N_34821,N_25940,N_25636);
nor U34822 (N_34822,N_21194,N_28069);
or U34823 (N_34823,N_27315,N_22153);
and U34824 (N_34824,N_27988,N_23383);
xnor U34825 (N_34825,N_21019,N_24584);
nor U34826 (N_34826,N_28605,N_25405);
nand U34827 (N_34827,N_21585,N_22564);
or U34828 (N_34828,N_24960,N_20871);
nor U34829 (N_34829,N_22311,N_20745);
and U34830 (N_34830,N_23856,N_21781);
and U34831 (N_34831,N_21068,N_23753);
nand U34832 (N_34832,N_24989,N_22785);
and U34833 (N_34833,N_20240,N_22398);
xnor U34834 (N_34834,N_25284,N_24112);
or U34835 (N_34835,N_29843,N_20626);
or U34836 (N_34836,N_20442,N_20992);
nor U34837 (N_34837,N_26605,N_26146);
nand U34838 (N_34838,N_26917,N_27716);
or U34839 (N_34839,N_27186,N_24275);
nand U34840 (N_34840,N_26087,N_20522);
and U34841 (N_34841,N_27082,N_21198);
nand U34842 (N_34842,N_29920,N_27154);
nand U34843 (N_34843,N_23745,N_22389);
xor U34844 (N_34844,N_26407,N_29751);
nor U34845 (N_34845,N_20518,N_22830);
xor U34846 (N_34846,N_26525,N_27446);
nand U34847 (N_34847,N_20242,N_25653);
nand U34848 (N_34848,N_28714,N_29430);
nand U34849 (N_34849,N_25469,N_26129);
and U34850 (N_34850,N_27571,N_20031);
nand U34851 (N_34851,N_25471,N_22804);
xnor U34852 (N_34852,N_21952,N_22404);
and U34853 (N_34853,N_23373,N_28802);
nor U34854 (N_34854,N_21229,N_29995);
or U34855 (N_34855,N_21546,N_20037);
nor U34856 (N_34856,N_27501,N_23539);
xor U34857 (N_34857,N_24005,N_23382);
and U34858 (N_34858,N_21004,N_21489);
and U34859 (N_34859,N_22960,N_27366);
or U34860 (N_34860,N_20290,N_22310);
xnor U34861 (N_34861,N_23601,N_20424);
and U34862 (N_34862,N_27751,N_20536);
and U34863 (N_34863,N_25674,N_22051);
nor U34864 (N_34864,N_26312,N_29204);
xnor U34865 (N_34865,N_27992,N_23358);
and U34866 (N_34866,N_27231,N_29515);
nand U34867 (N_34867,N_27053,N_22352);
or U34868 (N_34868,N_27858,N_23848);
or U34869 (N_34869,N_27070,N_21466);
or U34870 (N_34870,N_20836,N_29243);
nand U34871 (N_34871,N_22695,N_21483);
nor U34872 (N_34872,N_21518,N_26391);
or U34873 (N_34873,N_25947,N_29242);
nor U34874 (N_34874,N_26706,N_21910);
nand U34875 (N_34875,N_22027,N_25193);
nor U34876 (N_34876,N_24055,N_28422);
or U34877 (N_34877,N_22569,N_27656);
or U34878 (N_34878,N_25486,N_26451);
and U34879 (N_34879,N_22945,N_24988);
xnor U34880 (N_34880,N_23854,N_20084);
nand U34881 (N_34881,N_29913,N_27342);
nand U34882 (N_34882,N_20367,N_25923);
xor U34883 (N_34883,N_23334,N_25456);
and U34884 (N_34884,N_20160,N_23435);
nor U34885 (N_34885,N_29845,N_25358);
and U34886 (N_34886,N_22264,N_25014);
and U34887 (N_34887,N_23432,N_20003);
nor U34888 (N_34888,N_21002,N_29495);
or U34889 (N_34889,N_21929,N_29883);
and U34890 (N_34890,N_25848,N_28460);
nand U34891 (N_34891,N_27424,N_26933);
and U34892 (N_34892,N_22947,N_25298);
xnor U34893 (N_34893,N_21924,N_29566);
nor U34894 (N_34894,N_23241,N_28079);
and U34895 (N_34895,N_23421,N_24498);
nand U34896 (N_34896,N_21989,N_26447);
nand U34897 (N_34897,N_21468,N_22121);
or U34898 (N_34898,N_29710,N_20791);
and U34899 (N_34899,N_22015,N_25487);
and U34900 (N_34900,N_26133,N_23023);
xnor U34901 (N_34901,N_28078,N_22908);
nor U34902 (N_34902,N_26075,N_28035);
nor U34903 (N_34903,N_23565,N_28167);
nor U34904 (N_34904,N_20619,N_25812);
and U34905 (N_34905,N_25098,N_20861);
and U34906 (N_34906,N_27735,N_20402);
nand U34907 (N_34907,N_26516,N_21316);
xnor U34908 (N_34908,N_24923,N_25092);
nand U34909 (N_34909,N_24345,N_28509);
and U34910 (N_34910,N_26827,N_27229);
and U34911 (N_34911,N_21690,N_20891);
and U34912 (N_34912,N_23901,N_23911);
nand U34913 (N_34913,N_25025,N_20006);
and U34914 (N_34914,N_22619,N_27827);
xnor U34915 (N_34915,N_28646,N_22598);
nand U34916 (N_34916,N_20550,N_21166);
xor U34917 (N_34917,N_22802,N_20487);
or U34918 (N_34918,N_21670,N_26162);
xnor U34919 (N_34919,N_29819,N_24806);
nor U34920 (N_34920,N_29461,N_29442);
xnor U34921 (N_34921,N_20970,N_24631);
xor U34922 (N_34922,N_20783,N_22558);
and U34923 (N_34923,N_20665,N_24712);
nor U34924 (N_34924,N_28002,N_26512);
nand U34925 (N_34925,N_25783,N_25168);
nor U34926 (N_34926,N_25676,N_22937);
and U34927 (N_34927,N_27586,N_20541);
xor U34928 (N_34928,N_26535,N_27532);
xnor U34929 (N_34929,N_28433,N_23758);
nand U34930 (N_34930,N_29040,N_25883);
and U34931 (N_34931,N_28097,N_27561);
or U34932 (N_34932,N_28149,N_20057);
nor U34933 (N_34933,N_25177,N_21505);
and U34934 (N_34934,N_28462,N_21196);
nand U34935 (N_34935,N_23762,N_26376);
or U34936 (N_34936,N_25833,N_29655);
or U34937 (N_34937,N_24515,N_28176);
or U34938 (N_34938,N_28976,N_20744);
nand U34939 (N_34939,N_24730,N_29607);
or U34940 (N_34940,N_27860,N_22007);
nand U34941 (N_34941,N_21250,N_20376);
nand U34942 (N_34942,N_27535,N_23184);
or U34943 (N_34943,N_21523,N_24943);
xor U34944 (N_34944,N_26772,N_29483);
nor U34945 (N_34945,N_24483,N_29177);
xor U34946 (N_34946,N_20502,N_23760);
nand U34947 (N_34947,N_29895,N_24399);
nand U34948 (N_34948,N_21387,N_28379);
and U34949 (N_34949,N_27497,N_27286);
nand U34950 (N_34950,N_24897,N_22970);
nor U34951 (N_34951,N_20811,N_22683);
nor U34952 (N_34952,N_27235,N_28318);
nand U34953 (N_34953,N_23158,N_25311);
nand U34954 (N_34954,N_28594,N_22024);
nand U34955 (N_34955,N_25433,N_25439);
nand U34956 (N_34956,N_24092,N_20491);
nor U34957 (N_34957,N_25915,N_21491);
and U34958 (N_34958,N_29514,N_20341);
or U34959 (N_34959,N_22416,N_24497);
xor U34960 (N_34960,N_29149,N_21969);
nand U34961 (N_34961,N_21191,N_28157);
xnor U34962 (N_34962,N_24670,N_26218);
nand U34963 (N_34963,N_21586,N_26149);
nand U34964 (N_34964,N_26125,N_25461);
nand U34965 (N_34965,N_28360,N_22258);
xnor U34966 (N_34966,N_22103,N_25131);
and U34967 (N_34967,N_20060,N_20176);
and U34968 (N_34968,N_28533,N_27559);
nor U34969 (N_34969,N_26596,N_26057);
and U34970 (N_34970,N_20569,N_26164);
xor U34971 (N_34971,N_21612,N_29125);
xnor U34972 (N_34972,N_20777,N_25345);
nand U34973 (N_34973,N_21751,N_28982);
nand U34974 (N_34974,N_25868,N_28541);
xnor U34975 (N_34975,N_26631,N_26183);
nand U34976 (N_34976,N_23471,N_23502);
and U34977 (N_34977,N_26928,N_28939);
nand U34978 (N_34978,N_28199,N_22865);
nand U34979 (N_34979,N_23575,N_27048);
or U34980 (N_34980,N_27639,N_27196);
nor U34981 (N_34981,N_22510,N_24341);
nand U34982 (N_34982,N_26283,N_22686);
nand U34983 (N_34983,N_25593,N_22411);
xor U34984 (N_34984,N_27859,N_21951);
nand U34985 (N_34985,N_20933,N_24725);
nor U34986 (N_34986,N_25961,N_24394);
nor U34987 (N_34987,N_25762,N_28941);
nor U34988 (N_34988,N_26540,N_26398);
nand U34989 (N_34989,N_26616,N_29844);
or U34990 (N_34990,N_22090,N_24929);
xor U34991 (N_34991,N_28932,N_28416);
or U34992 (N_34992,N_20879,N_20028);
or U34993 (N_34993,N_25792,N_22185);
nand U34994 (N_34994,N_21984,N_24905);
or U34995 (N_34995,N_21440,N_21562);
nand U34996 (N_34996,N_29746,N_26279);
and U34997 (N_34997,N_23260,N_28277);
and U34998 (N_34998,N_22561,N_25663);
or U34999 (N_34999,N_26609,N_29985);
or U35000 (N_35000,N_23948,N_26294);
and U35001 (N_35001,N_26416,N_23563);
xor U35002 (N_35002,N_26900,N_26616);
and U35003 (N_35003,N_21779,N_22031);
and U35004 (N_35004,N_22969,N_20652);
nand U35005 (N_35005,N_22894,N_28916);
or U35006 (N_35006,N_21609,N_25983);
nor U35007 (N_35007,N_29030,N_29246);
or U35008 (N_35008,N_24931,N_28008);
xnor U35009 (N_35009,N_29856,N_26419);
or U35010 (N_35010,N_27344,N_23456);
xor U35011 (N_35011,N_22243,N_27395);
xor U35012 (N_35012,N_20195,N_22458);
nor U35013 (N_35013,N_21477,N_21565);
nor U35014 (N_35014,N_21371,N_26642);
xor U35015 (N_35015,N_22066,N_24407);
xnor U35016 (N_35016,N_20273,N_26073);
nor U35017 (N_35017,N_25026,N_29089);
nor U35018 (N_35018,N_25355,N_22397);
nor U35019 (N_35019,N_26709,N_28500);
or U35020 (N_35020,N_23727,N_20993);
and U35021 (N_35021,N_23407,N_21650);
or U35022 (N_35022,N_23982,N_24158);
nand U35023 (N_35023,N_20796,N_24156);
and U35024 (N_35024,N_28167,N_22909);
and U35025 (N_35025,N_25175,N_22134);
nand U35026 (N_35026,N_26384,N_21429);
xor U35027 (N_35027,N_26111,N_21465);
nand U35028 (N_35028,N_24403,N_24534);
nor U35029 (N_35029,N_22709,N_24112);
and U35030 (N_35030,N_23408,N_28169);
xnor U35031 (N_35031,N_28500,N_20355);
nor U35032 (N_35032,N_28289,N_24604);
nand U35033 (N_35033,N_29963,N_22332);
nor U35034 (N_35034,N_25061,N_28867);
nor U35035 (N_35035,N_28740,N_26447);
nand U35036 (N_35036,N_26913,N_23665);
and U35037 (N_35037,N_25398,N_21827);
nand U35038 (N_35038,N_20530,N_27387);
and U35039 (N_35039,N_21564,N_25603);
xor U35040 (N_35040,N_21840,N_27194);
or U35041 (N_35041,N_24368,N_27515);
and U35042 (N_35042,N_25518,N_29982);
or U35043 (N_35043,N_29130,N_26075);
nand U35044 (N_35044,N_27101,N_29801);
and U35045 (N_35045,N_25738,N_25140);
nor U35046 (N_35046,N_24665,N_21198);
nand U35047 (N_35047,N_26088,N_27989);
or U35048 (N_35048,N_23469,N_27929);
nand U35049 (N_35049,N_25128,N_21991);
xor U35050 (N_35050,N_26290,N_22110);
or U35051 (N_35051,N_25164,N_21442);
xnor U35052 (N_35052,N_28372,N_20418);
xnor U35053 (N_35053,N_20425,N_22089);
xnor U35054 (N_35054,N_24819,N_21875);
and U35055 (N_35055,N_22820,N_25090);
xor U35056 (N_35056,N_27108,N_23653);
and U35057 (N_35057,N_22556,N_27590);
nand U35058 (N_35058,N_25564,N_29151);
nor U35059 (N_35059,N_28522,N_27254);
or U35060 (N_35060,N_26475,N_28539);
and U35061 (N_35061,N_22990,N_20578);
nand U35062 (N_35062,N_23315,N_29264);
nand U35063 (N_35063,N_23090,N_21452);
nand U35064 (N_35064,N_22767,N_28710);
and U35065 (N_35065,N_29140,N_25375);
xor U35066 (N_35066,N_25034,N_23664);
xor U35067 (N_35067,N_27248,N_20268);
and U35068 (N_35068,N_29703,N_23121);
nand U35069 (N_35069,N_24552,N_24670);
nand U35070 (N_35070,N_28279,N_23598);
and U35071 (N_35071,N_20608,N_29042);
nor U35072 (N_35072,N_28927,N_22700);
xor U35073 (N_35073,N_27376,N_27836);
or U35074 (N_35074,N_23268,N_28754);
or U35075 (N_35075,N_24455,N_25066);
xor U35076 (N_35076,N_24045,N_21328);
and U35077 (N_35077,N_25697,N_24998);
nand U35078 (N_35078,N_20632,N_22694);
nand U35079 (N_35079,N_22121,N_29575);
nor U35080 (N_35080,N_24524,N_21732);
xor U35081 (N_35081,N_25331,N_21988);
nand U35082 (N_35082,N_20005,N_24474);
nor U35083 (N_35083,N_29710,N_21581);
xnor U35084 (N_35084,N_28131,N_28769);
and U35085 (N_35085,N_20755,N_25284);
nor U35086 (N_35086,N_29346,N_28024);
nor U35087 (N_35087,N_24099,N_26149);
or U35088 (N_35088,N_20402,N_23800);
and U35089 (N_35089,N_23004,N_28863);
xnor U35090 (N_35090,N_29765,N_21849);
or U35091 (N_35091,N_24064,N_24319);
nor U35092 (N_35092,N_25213,N_24015);
or U35093 (N_35093,N_20295,N_24903);
nor U35094 (N_35094,N_26674,N_20632);
and U35095 (N_35095,N_20231,N_23406);
and U35096 (N_35096,N_28697,N_24472);
nor U35097 (N_35097,N_21336,N_27941);
or U35098 (N_35098,N_26717,N_28352);
nor U35099 (N_35099,N_22167,N_27371);
nor U35100 (N_35100,N_24230,N_27112);
xor U35101 (N_35101,N_21488,N_23528);
nand U35102 (N_35102,N_27615,N_27427);
xor U35103 (N_35103,N_24308,N_20637);
xor U35104 (N_35104,N_23784,N_26856);
xnor U35105 (N_35105,N_28662,N_20910);
xor U35106 (N_35106,N_20766,N_24382);
nor U35107 (N_35107,N_21048,N_29514);
and U35108 (N_35108,N_20464,N_23791);
and U35109 (N_35109,N_29525,N_22821);
nor U35110 (N_35110,N_24225,N_23850);
nand U35111 (N_35111,N_28020,N_22975);
xor U35112 (N_35112,N_23958,N_22994);
xor U35113 (N_35113,N_22298,N_22926);
or U35114 (N_35114,N_20177,N_26560);
or U35115 (N_35115,N_27123,N_23663);
xnor U35116 (N_35116,N_20080,N_21321);
or U35117 (N_35117,N_21164,N_26940);
xor U35118 (N_35118,N_21177,N_27176);
xnor U35119 (N_35119,N_22093,N_28485);
nand U35120 (N_35120,N_23254,N_23158);
and U35121 (N_35121,N_24256,N_25232);
and U35122 (N_35122,N_28510,N_26337);
or U35123 (N_35123,N_26659,N_22708);
xnor U35124 (N_35124,N_25929,N_29384);
and U35125 (N_35125,N_26769,N_21432);
nor U35126 (N_35126,N_27180,N_20594);
xor U35127 (N_35127,N_22862,N_26917);
nand U35128 (N_35128,N_23727,N_23850);
nand U35129 (N_35129,N_22246,N_29641);
nand U35130 (N_35130,N_25286,N_23225);
or U35131 (N_35131,N_22350,N_29733);
xor U35132 (N_35132,N_23517,N_22268);
nand U35133 (N_35133,N_20149,N_26291);
nand U35134 (N_35134,N_27773,N_28949);
and U35135 (N_35135,N_27364,N_20405);
nand U35136 (N_35136,N_29970,N_29283);
nand U35137 (N_35137,N_21489,N_22458);
xnor U35138 (N_35138,N_25214,N_22604);
nor U35139 (N_35139,N_29111,N_21984);
nand U35140 (N_35140,N_24103,N_28847);
or U35141 (N_35141,N_20383,N_28079);
xor U35142 (N_35142,N_23026,N_22946);
nor U35143 (N_35143,N_26327,N_24969);
xnor U35144 (N_35144,N_20646,N_23651);
and U35145 (N_35145,N_26246,N_27238);
xor U35146 (N_35146,N_29684,N_20328);
nand U35147 (N_35147,N_23102,N_20956);
nand U35148 (N_35148,N_21003,N_20355);
nand U35149 (N_35149,N_20914,N_26484);
xnor U35150 (N_35150,N_24782,N_20900);
nand U35151 (N_35151,N_27317,N_20065);
and U35152 (N_35152,N_20989,N_26416);
nor U35153 (N_35153,N_25474,N_20972);
or U35154 (N_35154,N_20700,N_21203);
nand U35155 (N_35155,N_21746,N_21814);
nand U35156 (N_35156,N_22637,N_20780);
xor U35157 (N_35157,N_24988,N_28158);
nand U35158 (N_35158,N_26244,N_28291);
nand U35159 (N_35159,N_21838,N_25934);
nor U35160 (N_35160,N_24242,N_20602);
or U35161 (N_35161,N_27142,N_28086);
or U35162 (N_35162,N_22720,N_22895);
and U35163 (N_35163,N_22973,N_25281);
xor U35164 (N_35164,N_25359,N_28522);
and U35165 (N_35165,N_21719,N_27718);
or U35166 (N_35166,N_24690,N_28920);
nand U35167 (N_35167,N_22530,N_25880);
or U35168 (N_35168,N_21940,N_29061);
or U35169 (N_35169,N_24466,N_25129);
and U35170 (N_35170,N_28269,N_24776);
nand U35171 (N_35171,N_24285,N_23255);
nand U35172 (N_35172,N_23592,N_25027);
xor U35173 (N_35173,N_29790,N_23442);
xnor U35174 (N_35174,N_23357,N_23653);
or U35175 (N_35175,N_24313,N_20556);
nor U35176 (N_35176,N_20882,N_20829);
or U35177 (N_35177,N_21599,N_24693);
or U35178 (N_35178,N_29439,N_22407);
or U35179 (N_35179,N_26265,N_29171);
and U35180 (N_35180,N_20550,N_22503);
xnor U35181 (N_35181,N_26939,N_27668);
nand U35182 (N_35182,N_21539,N_23312);
or U35183 (N_35183,N_22075,N_22742);
and U35184 (N_35184,N_27129,N_20299);
and U35185 (N_35185,N_23930,N_29946);
xor U35186 (N_35186,N_21437,N_25223);
nor U35187 (N_35187,N_26818,N_29363);
or U35188 (N_35188,N_28680,N_23338);
xnor U35189 (N_35189,N_25333,N_20094);
nor U35190 (N_35190,N_27105,N_20020);
nor U35191 (N_35191,N_25443,N_23570);
nand U35192 (N_35192,N_22565,N_29087);
xor U35193 (N_35193,N_29295,N_27041);
and U35194 (N_35194,N_29207,N_23840);
xnor U35195 (N_35195,N_22540,N_26182);
xnor U35196 (N_35196,N_28584,N_24483);
xnor U35197 (N_35197,N_25967,N_27886);
and U35198 (N_35198,N_27138,N_21331);
nor U35199 (N_35199,N_29579,N_28947);
and U35200 (N_35200,N_27335,N_28055);
nand U35201 (N_35201,N_24407,N_25002);
and U35202 (N_35202,N_21083,N_25908);
xor U35203 (N_35203,N_25877,N_28095);
nand U35204 (N_35204,N_23224,N_20741);
nor U35205 (N_35205,N_29408,N_25734);
or U35206 (N_35206,N_25047,N_22585);
xor U35207 (N_35207,N_24455,N_21919);
and U35208 (N_35208,N_26946,N_20511);
nand U35209 (N_35209,N_26740,N_27823);
nor U35210 (N_35210,N_29238,N_22437);
nor U35211 (N_35211,N_27078,N_23389);
and U35212 (N_35212,N_23291,N_23060);
or U35213 (N_35213,N_24965,N_28944);
nand U35214 (N_35214,N_24317,N_20351);
nor U35215 (N_35215,N_28523,N_27750);
nor U35216 (N_35216,N_29698,N_20340);
and U35217 (N_35217,N_22864,N_28077);
xnor U35218 (N_35218,N_29619,N_25689);
nor U35219 (N_35219,N_21205,N_20543);
nor U35220 (N_35220,N_24099,N_20035);
and U35221 (N_35221,N_20027,N_27176);
nor U35222 (N_35222,N_26174,N_27307);
nor U35223 (N_35223,N_28764,N_20277);
xor U35224 (N_35224,N_23433,N_28570);
or U35225 (N_35225,N_28100,N_25362);
xnor U35226 (N_35226,N_24142,N_23143);
nand U35227 (N_35227,N_29158,N_28427);
or U35228 (N_35228,N_27704,N_23780);
nand U35229 (N_35229,N_24008,N_21935);
xnor U35230 (N_35230,N_20625,N_28074);
nand U35231 (N_35231,N_29278,N_21553);
nor U35232 (N_35232,N_20510,N_21504);
nor U35233 (N_35233,N_24972,N_28826);
nand U35234 (N_35234,N_26618,N_22415);
or U35235 (N_35235,N_29201,N_20950);
nor U35236 (N_35236,N_20720,N_25274);
nand U35237 (N_35237,N_25589,N_23858);
nand U35238 (N_35238,N_28586,N_21437);
nor U35239 (N_35239,N_23618,N_27763);
xnor U35240 (N_35240,N_21476,N_25872);
xor U35241 (N_35241,N_28501,N_23924);
and U35242 (N_35242,N_28901,N_28645);
xor U35243 (N_35243,N_29198,N_22738);
nand U35244 (N_35244,N_26221,N_21248);
nand U35245 (N_35245,N_27454,N_25540);
and U35246 (N_35246,N_28031,N_20066);
and U35247 (N_35247,N_20960,N_20278);
nand U35248 (N_35248,N_20333,N_24044);
xnor U35249 (N_35249,N_28025,N_24532);
nor U35250 (N_35250,N_21215,N_20565);
or U35251 (N_35251,N_24211,N_28672);
xnor U35252 (N_35252,N_26510,N_24729);
nor U35253 (N_35253,N_22618,N_26377);
xnor U35254 (N_35254,N_27294,N_27931);
nand U35255 (N_35255,N_20959,N_24722);
xnor U35256 (N_35256,N_25500,N_25551);
and U35257 (N_35257,N_22976,N_24739);
and U35258 (N_35258,N_21863,N_29312);
or U35259 (N_35259,N_28424,N_21868);
xnor U35260 (N_35260,N_28510,N_23240);
nor U35261 (N_35261,N_20878,N_20830);
xnor U35262 (N_35262,N_27483,N_29511);
or U35263 (N_35263,N_25475,N_20251);
and U35264 (N_35264,N_20944,N_22611);
nand U35265 (N_35265,N_26734,N_26490);
nand U35266 (N_35266,N_24010,N_26698);
nand U35267 (N_35267,N_25428,N_27782);
xnor U35268 (N_35268,N_20111,N_20775);
nor U35269 (N_35269,N_20438,N_24091);
nor U35270 (N_35270,N_25083,N_26945);
nor U35271 (N_35271,N_22142,N_27766);
xor U35272 (N_35272,N_26726,N_29677);
and U35273 (N_35273,N_20756,N_20049);
xnor U35274 (N_35274,N_27211,N_22914);
xor U35275 (N_35275,N_25932,N_23037);
xnor U35276 (N_35276,N_27845,N_27725);
nand U35277 (N_35277,N_26521,N_20011);
nand U35278 (N_35278,N_20248,N_21352);
or U35279 (N_35279,N_26682,N_26475);
nor U35280 (N_35280,N_25127,N_29582);
or U35281 (N_35281,N_24086,N_29751);
or U35282 (N_35282,N_28064,N_20923);
nor U35283 (N_35283,N_21435,N_24615);
and U35284 (N_35284,N_22171,N_20975);
nor U35285 (N_35285,N_20578,N_22290);
nand U35286 (N_35286,N_28961,N_20285);
nor U35287 (N_35287,N_26497,N_26774);
nor U35288 (N_35288,N_20233,N_29849);
nor U35289 (N_35289,N_20748,N_25650);
and U35290 (N_35290,N_22390,N_29305);
xor U35291 (N_35291,N_27553,N_26053);
xor U35292 (N_35292,N_21247,N_21312);
nor U35293 (N_35293,N_24528,N_23830);
or U35294 (N_35294,N_29099,N_28726);
and U35295 (N_35295,N_28191,N_23005);
nand U35296 (N_35296,N_24056,N_24943);
nand U35297 (N_35297,N_26918,N_28806);
nor U35298 (N_35298,N_27763,N_25789);
nand U35299 (N_35299,N_28117,N_20119);
xnor U35300 (N_35300,N_23521,N_24694);
xnor U35301 (N_35301,N_27843,N_21957);
nand U35302 (N_35302,N_25150,N_21780);
nor U35303 (N_35303,N_27164,N_23296);
or U35304 (N_35304,N_27279,N_20611);
xnor U35305 (N_35305,N_25473,N_23194);
and U35306 (N_35306,N_21085,N_22010);
or U35307 (N_35307,N_25300,N_28555);
and U35308 (N_35308,N_26222,N_20947);
nor U35309 (N_35309,N_22080,N_22505);
nand U35310 (N_35310,N_27002,N_20097);
nor U35311 (N_35311,N_20289,N_21450);
xor U35312 (N_35312,N_29440,N_20147);
and U35313 (N_35313,N_26584,N_26107);
xnor U35314 (N_35314,N_25017,N_22981);
or U35315 (N_35315,N_23128,N_22115);
nand U35316 (N_35316,N_23738,N_25426);
nor U35317 (N_35317,N_25221,N_25479);
and U35318 (N_35318,N_29091,N_28499);
or U35319 (N_35319,N_28830,N_24749);
nand U35320 (N_35320,N_29023,N_26067);
nand U35321 (N_35321,N_23323,N_23799);
xor U35322 (N_35322,N_20855,N_25585);
nor U35323 (N_35323,N_26601,N_21783);
and U35324 (N_35324,N_23840,N_29280);
or U35325 (N_35325,N_26414,N_28382);
nand U35326 (N_35326,N_28314,N_29488);
nor U35327 (N_35327,N_26610,N_22170);
and U35328 (N_35328,N_23650,N_27987);
and U35329 (N_35329,N_29214,N_23361);
nor U35330 (N_35330,N_25597,N_21705);
and U35331 (N_35331,N_23367,N_27042);
or U35332 (N_35332,N_23785,N_21716);
nand U35333 (N_35333,N_21935,N_20643);
and U35334 (N_35334,N_29263,N_22527);
xor U35335 (N_35335,N_24858,N_24624);
nand U35336 (N_35336,N_26393,N_20248);
xnor U35337 (N_35337,N_26233,N_25416);
and U35338 (N_35338,N_28848,N_22619);
nor U35339 (N_35339,N_27052,N_24556);
nand U35340 (N_35340,N_24363,N_28204);
xnor U35341 (N_35341,N_27544,N_29293);
nor U35342 (N_35342,N_20646,N_23444);
or U35343 (N_35343,N_27864,N_27405);
nor U35344 (N_35344,N_27811,N_28199);
nand U35345 (N_35345,N_22157,N_23621);
or U35346 (N_35346,N_23730,N_28022);
nor U35347 (N_35347,N_21244,N_29448);
nor U35348 (N_35348,N_29040,N_23938);
nor U35349 (N_35349,N_25464,N_27142);
nand U35350 (N_35350,N_27819,N_25237);
xnor U35351 (N_35351,N_23248,N_29224);
and U35352 (N_35352,N_21563,N_26329);
nand U35353 (N_35353,N_26069,N_20370);
xor U35354 (N_35354,N_25168,N_28770);
nand U35355 (N_35355,N_22193,N_24801);
nor U35356 (N_35356,N_24045,N_27191);
nand U35357 (N_35357,N_22772,N_27919);
or U35358 (N_35358,N_24572,N_21655);
xnor U35359 (N_35359,N_29679,N_28247);
xor U35360 (N_35360,N_28992,N_25044);
nor U35361 (N_35361,N_23638,N_23818);
and U35362 (N_35362,N_22443,N_27229);
and U35363 (N_35363,N_25504,N_24261);
and U35364 (N_35364,N_27225,N_24373);
nand U35365 (N_35365,N_20849,N_29553);
nor U35366 (N_35366,N_26108,N_29587);
xor U35367 (N_35367,N_23428,N_20070);
nor U35368 (N_35368,N_20396,N_21180);
and U35369 (N_35369,N_25878,N_21132);
and U35370 (N_35370,N_24293,N_28475);
or U35371 (N_35371,N_20217,N_21587);
and U35372 (N_35372,N_28846,N_28733);
or U35373 (N_35373,N_20388,N_20590);
nand U35374 (N_35374,N_27473,N_25450);
xnor U35375 (N_35375,N_26483,N_24134);
nand U35376 (N_35376,N_25542,N_27617);
xor U35377 (N_35377,N_26414,N_20499);
xnor U35378 (N_35378,N_27311,N_27608);
and U35379 (N_35379,N_23164,N_21247);
nand U35380 (N_35380,N_20433,N_24633);
xor U35381 (N_35381,N_23504,N_23855);
or U35382 (N_35382,N_29953,N_28301);
nor U35383 (N_35383,N_26267,N_23477);
and U35384 (N_35384,N_23013,N_20507);
nand U35385 (N_35385,N_29244,N_26275);
nor U35386 (N_35386,N_20031,N_20049);
nand U35387 (N_35387,N_20668,N_27463);
nor U35388 (N_35388,N_20179,N_26011);
xnor U35389 (N_35389,N_26653,N_27434);
or U35390 (N_35390,N_20546,N_25714);
nor U35391 (N_35391,N_28337,N_23099);
xnor U35392 (N_35392,N_27690,N_25081);
xor U35393 (N_35393,N_26671,N_25708);
and U35394 (N_35394,N_20851,N_24674);
xnor U35395 (N_35395,N_22130,N_23486);
nor U35396 (N_35396,N_27641,N_29970);
and U35397 (N_35397,N_20684,N_29129);
or U35398 (N_35398,N_22075,N_23779);
or U35399 (N_35399,N_28671,N_27197);
xnor U35400 (N_35400,N_22239,N_22852);
and U35401 (N_35401,N_29833,N_23554);
or U35402 (N_35402,N_27526,N_23736);
nor U35403 (N_35403,N_20688,N_22060);
and U35404 (N_35404,N_24991,N_25335);
nand U35405 (N_35405,N_20396,N_24432);
nand U35406 (N_35406,N_24811,N_21346);
nor U35407 (N_35407,N_29537,N_23208);
nand U35408 (N_35408,N_29750,N_20821);
nor U35409 (N_35409,N_27309,N_27351);
xor U35410 (N_35410,N_29051,N_23744);
and U35411 (N_35411,N_28695,N_22867);
and U35412 (N_35412,N_27919,N_27250);
nor U35413 (N_35413,N_25192,N_27601);
nand U35414 (N_35414,N_27131,N_27746);
and U35415 (N_35415,N_25306,N_29329);
nand U35416 (N_35416,N_28566,N_28025);
or U35417 (N_35417,N_20045,N_26368);
xor U35418 (N_35418,N_21480,N_23931);
nand U35419 (N_35419,N_21813,N_25677);
or U35420 (N_35420,N_28012,N_26210);
or U35421 (N_35421,N_21235,N_26633);
nand U35422 (N_35422,N_22070,N_21182);
nor U35423 (N_35423,N_20259,N_20324);
and U35424 (N_35424,N_25213,N_21006);
and U35425 (N_35425,N_27430,N_27426);
and U35426 (N_35426,N_27006,N_25244);
nor U35427 (N_35427,N_22686,N_23226);
nand U35428 (N_35428,N_22050,N_29244);
nand U35429 (N_35429,N_20338,N_28159);
and U35430 (N_35430,N_27540,N_27723);
and U35431 (N_35431,N_29839,N_25562);
nor U35432 (N_35432,N_29324,N_26727);
and U35433 (N_35433,N_23263,N_20047);
xnor U35434 (N_35434,N_23753,N_23630);
and U35435 (N_35435,N_29842,N_22971);
and U35436 (N_35436,N_27441,N_23579);
and U35437 (N_35437,N_20704,N_21447);
xnor U35438 (N_35438,N_23596,N_20595);
xor U35439 (N_35439,N_25453,N_29042);
nand U35440 (N_35440,N_20897,N_28121);
nand U35441 (N_35441,N_23835,N_22201);
or U35442 (N_35442,N_28434,N_24658);
nor U35443 (N_35443,N_23837,N_21428);
or U35444 (N_35444,N_24435,N_23628);
xnor U35445 (N_35445,N_27427,N_20545);
or U35446 (N_35446,N_23934,N_25271);
nor U35447 (N_35447,N_29174,N_29940);
and U35448 (N_35448,N_22209,N_28638);
or U35449 (N_35449,N_24589,N_27060);
xor U35450 (N_35450,N_25682,N_20503);
xnor U35451 (N_35451,N_29696,N_23570);
and U35452 (N_35452,N_21231,N_23164);
nor U35453 (N_35453,N_28155,N_26950);
nand U35454 (N_35454,N_29673,N_29612);
or U35455 (N_35455,N_24300,N_28888);
nor U35456 (N_35456,N_26119,N_25569);
nor U35457 (N_35457,N_20943,N_29134);
and U35458 (N_35458,N_22201,N_22602);
or U35459 (N_35459,N_29696,N_22223);
xor U35460 (N_35460,N_27202,N_29522);
and U35461 (N_35461,N_24736,N_20174);
or U35462 (N_35462,N_26792,N_28986);
nand U35463 (N_35463,N_25062,N_23687);
xnor U35464 (N_35464,N_26053,N_24842);
and U35465 (N_35465,N_27407,N_25832);
and U35466 (N_35466,N_21329,N_27632);
and U35467 (N_35467,N_26591,N_29291);
and U35468 (N_35468,N_25885,N_24635);
or U35469 (N_35469,N_21143,N_26699);
or U35470 (N_35470,N_24368,N_26969);
nor U35471 (N_35471,N_20270,N_23821);
nand U35472 (N_35472,N_22420,N_27664);
nand U35473 (N_35473,N_23845,N_29506);
and U35474 (N_35474,N_27841,N_29589);
or U35475 (N_35475,N_20910,N_22712);
and U35476 (N_35476,N_20526,N_24754);
and U35477 (N_35477,N_22942,N_21115);
and U35478 (N_35478,N_27503,N_25379);
or U35479 (N_35479,N_20070,N_22579);
nand U35480 (N_35480,N_22198,N_23367);
and U35481 (N_35481,N_29007,N_22891);
and U35482 (N_35482,N_24531,N_27356);
nor U35483 (N_35483,N_25366,N_29942);
and U35484 (N_35484,N_24038,N_22778);
or U35485 (N_35485,N_23991,N_26652);
and U35486 (N_35486,N_26009,N_29825);
or U35487 (N_35487,N_24602,N_28282);
xor U35488 (N_35488,N_23038,N_29940);
and U35489 (N_35489,N_27689,N_22367);
nand U35490 (N_35490,N_29378,N_27116);
and U35491 (N_35491,N_21088,N_20107);
nor U35492 (N_35492,N_29527,N_21074);
or U35493 (N_35493,N_22414,N_25853);
or U35494 (N_35494,N_25711,N_29078);
nor U35495 (N_35495,N_25393,N_27978);
or U35496 (N_35496,N_23627,N_25428);
nor U35497 (N_35497,N_29934,N_20113);
nor U35498 (N_35498,N_29690,N_25176);
xor U35499 (N_35499,N_22881,N_23123);
xnor U35500 (N_35500,N_26772,N_24950);
xnor U35501 (N_35501,N_20308,N_29711);
and U35502 (N_35502,N_26764,N_21233);
and U35503 (N_35503,N_24690,N_21635);
and U35504 (N_35504,N_25228,N_20984);
xor U35505 (N_35505,N_21506,N_29522);
xor U35506 (N_35506,N_25684,N_23014);
nand U35507 (N_35507,N_24645,N_26286);
nand U35508 (N_35508,N_22887,N_26767);
or U35509 (N_35509,N_25950,N_27799);
and U35510 (N_35510,N_21814,N_25470);
or U35511 (N_35511,N_23339,N_28285);
xnor U35512 (N_35512,N_27537,N_27347);
nor U35513 (N_35513,N_22011,N_28805);
nand U35514 (N_35514,N_21128,N_22046);
or U35515 (N_35515,N_26968,N_20806);
and U35516 (N_35516,N_25328,N_21565);
xnor U35517 (N_35517,N_20408,N_20416);
or U35518 (N_35518,N_26215,N_22144);
xor U35519 (N_35519,N_23360,N_20001);
nor U35520 (N_35520,N_29030,N_29646);
nand U35521 (N_35521,N_25068,N_25248);
or U35522 (N_35522,N_26981,N_20992);
nor U35523 (N_35523,N_27701,N_20213);
or U35524 (N_35524,N_27609,N_22010);
nor U35525 (N_35525,N_20913,N_24494);
nor U35526 (N_35526,N_25851,N_22219);
nand U35527 (N_35527,N_22851,N_22019);
nor U35528 (N_35528,N_27298,N_21916);
nand U35529 (N_35529,N_20964,N_22245);
or U35530 (N_35530,N_29684,N_21606);
or U35531 (N_35531,N_29880,N_23372);
xnor U35532 (N_35532,N_28630,N_27519);
and U35533 (N_35533,N_27784,N_26711);
xnor U35534 (N_35534,N_24736,N_24861);
and U35535 (N_35535,N_21053,N_20885);
nor U35536 (N_35536,N_20125,N_28928);
nor U35537 (N_35537,N_23417,N_22918);
or U35538 (N_35538,N_22863,N_20275);
xnor U35539 (N_35539,N_28041,N_24199);
xor U35540 (N_35540,N_23412,N_22868);
nand U35541 (N_35541,N_29907,N_29623);
nor U35542 (N_35542,N_27325,N_29921);
nor U35543 (N_35543,N_26147,N_23394);
and U35544 (N_35544,N_25409,N_26595);
nor U35545 (N_35545,N_28170,N_29815);
or U35546 (N_35546,N_22039,N_22542);
and U35547 (N_35547,N_21492,N_26754);
nor U35548 (N_35548,N_25722,N_24678);
xor U35549 (N_35549,N_27019,N_26297);
or U35550 (N_35550,N_26320,N_28645);
or U35551 (N_35551,N_20519,N_20352);
nor U35552 (N_35552,N_27806,N_23597);
or U35553 (N_35553,N_27597,N_23490);
and U35554 (N_35554,N_20067,N_28348);
xnor U35555 (N_35555,N_24714,N_27090);
nor U35556 (N_35556,N_21323,N_28758);
and U35557 (N_35557,N_21577,N_21421);
nand U35558 (N_35558,N_28959,N_25514);
and U35559 (N_35559,N_26553,N_20076);
nand U35560 (N_35560,N_20364,N_28115);
xor U35561 (N_35561,N_24060,N_26997);
and U35562 (N_35562,N_20385,N_27816);
nand U35563 (N_35563,N_22770,N_21890);
and U35564 (N_35564,N_28001,N_22149);
or U35565 (N_35565,N_20084,N_21101);
xor U35566 (N_35566,N_28874,N_25743);
or U35567 (N_35567,N_22719,N_23534);
xnor U35568 (N_35568,N_25987,N_25641);
xor U35569 (N_35569,N_24404,N_21349);
or U35570 (N_35570,N_21551,N_25002);
and U35571 (N_35571,N_22397,N_27789);
nor U35572 (N_35572,N_23077,N_24043);
or U35573 (N_35573,N_23231,N_26930);
or U35574 (N_35574,N_29426,N_21812);
xnor U35575 (N_35575,N_25838,N_24550);
xnor U35576 (N_35576,N_27453,N_23937);
nor U35577 (N_35577,N_22081,N_23938);
nand U35578 (N_35578,N_24342,N_22102);
or U35579 (N_35579,N_21642,N_26708);
xor U35580 (N_35580,N_28228,N_26443);
or U35581 (N_35581,N_25277,N_27831);
xor U35582 (N_35582,N_26657,N_28705);
and U35583 (N_35583,N_25716,N_24933);
or U35584 (N_35584,N_29560,N_21082);
and U35585 (N_35585,N_25449,N_24160);
and U35586 (N_35586,N_25062,N_21362);
or U35587 (N_35587,N_22543,N_25555);
or U35588 (N_35588,N_28305,N_21134);
or U35589 (N_35589,N_20667,N_25544);
nor U35590 (N_35590,N_24283,N_26230);
nand U35591 (N_35591,N_29516,N_27242);
and U35592 (N_35592,N_25219,N_21515);
nand U35593 (N_35593,N_20222,N_24751);
xnor U35594 (N_35594,N_26212,N_24409);
or U35595 (N_35595,N_27731,N_20510);
and U35596 (N_35596,N_20378,N_24319);
nor U35597 (N_35597,N_20325,N_25396);
or U35598 (N_35598,N_29915,N_27185);
xnor U35599 (N_35599,N_21791,N_21446);
and U35600 (N_35600,N_24164,N_28510);
or U35601 (N_35601,N_21184,N_26706);
or U35602 (N_35602,N_23024,N_20930);
xnor U35603 (N_35603,N_26962,N_29982);
nand U35604 (N_35604,N_23531,N_20814);
or U35605 (N_35605,N_21566,N_24345);
or U35606 (N_35606,N_24165,N_27472);
and U35607 (N_35607,N_29680,N_20589);
and U35608 (N_35608,N_21229,N_26431);
and U35609 (N_35609,N_23437,N_23490);
and U35610 (N_35610,N_26801,N_23621);
nand U35611 (N_35611,N_29183,N_22715);
and U35612 (N_35612,N_21220,N_26821);
nand U35613 (N_35613,N_25751,N_20181);
xnor U35614 (N_35614,N_28077,N_24259);
or U35615 (N_35615,N_21057,N_22707);
xnor U35616 (N_35616,N_20441,N_23632);
nand U35617 (N_35617,N_28809,N_21459);
nand U35618 (N_35618,N_23899,N_26536);
xor U35619 (N_35619,N_28361,N_23867);
and U35620 (N_35620,N_23023,N_24627);
nand U35621 (N_35621,N_25074,N_20373);
or U35622 (N_35622,N_21384,N_20566);
nor U35623 (N_35623,N_25017,N_21070);
and U35624 (N_35624,N_24733,N_21261);
nand U35625 (N_35625,N_24145,N_22630);
nand U35626 (N_35626,N_29939,N_20438);
nand U35627 (N_35627,N_29302,N_27733);
nand U35628 (N_35628,N_22885,N_23311);
or U35629 (N_35629,N_29096,N_28810);
and U35630 (N_35630,N_27096,N_24161);
or U35631 (N_35631,N_21770,N_26941);
xnor U35632 (N_35632,N_27952,N_26983);
xor U35633 (N_35633,N_23230,N_22669);
nor U35634 (N_35634,N_27813,N_23866);
and U35635 (N_35635,N_21437,N_24857);
and U35636 (N_35636,N_24674,N_22117);
and U35637 (N_35637,N_25468,N_22784);
or U35638 (N_35638,N_27304,N_22103);
xnor U35639 (N_35639,N_24929,N_26445);
xnor U35640 (N_35640,N_28085,N_22565);
or U35641 (N_35641,N_26445,N_24601);
or U35642 (N_35642,N_24373,N_29401);
and U35643 (N_35643,N_22399,N_26760);
or U35644 (N_35644,N_20086,N_20276);
xnor U35645 (N_35645,N_21518,N_28435);
nor U35646 (N_35646,N_26792,N_20376);
or U35647 (N_35647,N_21918,N_28258);
and U35648 (N_35648,N_24973,N_22221);
xor U35649 (N_35649,N_27502,N_24265);
nand U35650 (N_35650,N_25635,N_29028);
and U35651 (N_35651,N_28279,N_20946);
or U35652 (N_35652,N_27817,N_22687);
and U35653 (N_35653,N_26929,N_29771);
xnor U35654 (N_35654,N_27951,N_22656);
xor U35655 (N_35655,N_22692,N_20902);
nor U35656 (N_35656,N_20404,N_29887);
nand U35657 (N_35657,N_24159,N_24014);
nor U35658 (N_35658,N_20496,N_20224);
xor U35659 (N_35659,N_20177,N_28238);
or U35660 (N_35660,N_27037,N_25727);
or U35661 (N_35661,N_20690,N_27531);
and U35662 (N_35662,N_21600,N_21032);
nor U35663 (N_35663,N_26644,N_25032);
nand U35664 (N_35664,N_21755,N_23925);
and U35665 (N_35665,N_20406,N_27059);
and U35666 (N_35666,N_20434,N_22704);
xor U35667 (N_35667,N_28468,N_28229);
or U35668 (N_35668,N_24809,N_24119);
and U35669 (N_35669,N_29650,N_26661);
xnor U35670 (N_35670,N_20782,N_22682);
and U35671 (N_35671,N_24591,N_26000);
nor U35672 (N_35672,N_25925,N_23351);
and U35673 (N_35673,N_22405,N_23723);
nand U35674 (N_35674,N_22804,N_22852);
and U35675 (N_35675,N_26646,N_23151);
or U35676 (N_35676,N_28906,N_24029);
or U35677 (N_35677,N_21420,N_23960);
nand U35678 (N_35678,N_29618,N_27390);
nand U35679 (N_35679,N_27682,N_22046);
or U35680 (N_35680,N_20625,N_21563);
xnor U35681 (N_35681,N_25846,N_25393);
xor U35682 (N_35682,N_26165,N_24884);
and U35683 (N_35683,N_21056,N_25246);
xor U35684 (N_35684,N_22409,N_29627);
and U35685 (N_35685,N_26235,N_27138);
nand U35686 (N_35686,N_28410,N_26072);
or U35687 (N_35687,N_23388,N_23235);
nand U35688 (N_35688,N_21597,N_28243);
and U35689 (N_35689,N_20382,N_27170);
nand U35690 (N_35690,N_29822,N_23160);
or U35691 (N_35691,N_29021,N_28676);
or U35692 (N_35692,N_23238,N_20178);
xnor U35693 (N_35693,N_21661,N_23498);
or U35694 (N_35694,N_22433,N_27210);
and U35695 (N_35695,N_28800,N_28758);
or U35696 (N_35696,N_26667,N_26058);
or U35697 (N_35697,N_22239,N_26448);
nor U35698 (N_35698,N_21911,N_22123);
xor U35699 (N_35699,N_23769,N_22050);
nor U35700 (N_35700,N_23739,N_26354);
or U35701 (N_35701,N_27990,N_23436);
nand U35702 (N_35702,N_27912,N_23668);
and U35703 (N_35703,N_27972,N_28659);
nor U35704 (N_35704,N_23603,N_27060);
nor U35705 (N_35705,N_24037,N_22517);
xor U35706 (N_35706,N_28964,N_22095);
nand U35707 (N_35707,N_26798,N_27257);
or U35708 (N_35708,N_20101,N_22357);
nor U35709 (N_35709,N_27528,N_25387);
nor U35710 (N_35710,N_20252,N_27435);
xor U35711 (N_35711,N_29744,N_29726);
xnor U35712 (N_35712,N_29245,N_22138);
nand U35713 (N_35713,N_24459,N_26795);
nor U35714 (N_35714,N_24768,N_20976);
nor U35715 (N_35715,N_29402,N_21271);
or U35716 (N_35716,N_25834,N_26875);
or U35717 (N_35717,N_27210,N_27003);
nor U35718 (N_35718,N_21825,N_21006);
nand U35719 (N_35719,N_24092,N_20355);
or U35720 (N_35720,N_23527,N_21270);
nand U35721 (N_35721,N_26017,N_20750);
or U35722 (N_35722,N_26896,N_29101);
nor U35723 (N_35723,N_28765,N_27947);
nand U35724 (N_35724,N_23467,N_22712);
or U35725 (N_35725,N_20446,N_21358);
nand U35726 (N_35726,N_23517,N_20159);
nand U35727 (N_35727,N_20072,N_23201);
or U35728 (N_35728,N_23143,N_26106);
and U35729 (N_35729,N_25372,N_21322);
nor U35730 (N_35730,N_29427,N_26055);
and U35731 (N_35731,N_26464,N_22792);
or U35732 (N_35732,N_26992,N_26677);
nor U35733 (N_35733,N_22844,N_27716);
nand U35734 (N_35734,N_28250,N_25180);
or U35735 (N_35735,N_23281,N_27773);
nand U35736 (N_35736,N_23922,N_27501);
nand U35737 (N_35737,N_20354,N_25020);
and U35738 (N_35738,N_20104,N_21081);
nor U35739 (N_35739,N_28759,N_21971);
nand U35740 (N_35740,N_24853,N_22524);
nor U35741 (N_35741,N_23987,N_20303);
and U35742 (N_35742,N_22164,N_21995);
nand U35743 (N_35743,N_28360,N_23900);
or U35744 (N_35744,N_24400,N_21358);
and U35745 (N_35745,N_21907,N_20698);
and U35746 (N_35746,N_24789,N_20395);
xnor U35747 (N_35747,N_20954,N_25084);
and U35748 (N_35748,N_28279,N_27540);
nor U35749 (N_35749,N_29175,N_28582);
nand U35750 (N_35750,N_23072,N_22217);
and U35751 (N_35751,N_23444,N_22715);
xor U35752 (N_35752,N_22678,N_26744);
nor U35753 (N_35753,N_26762,N_22510);
and U35754 (N_35754,N_25514,N_21181);
or U35755 (N_35755,N_25921,N_21921);
xor U35756 (N_35756,N_28247,N_21934);
nand U35757 (N_35757,N_23132,N_25183);
or U35758 (N_35758,N_21630,N_27159);
or U35759 (N_35759,N_24629,N_26299);
or U35760 (N_35760,N_23171,N_20064);
or U35761 (N_35761,N_26012,N_23165);
nand U35762 (N_35762,N_29508,N_20036);
nand U35763 (N_35763,N_20084,N_29797);
and U35764 (N_35764,N_27258,N_21787);
nand U35765 (N_35765,N_23811,N_21992);
nand U35766 (N_35766,N_28177,N_28772);
xor U35767 (N_35767,N_25846,N_28139);
nand U35768 (N_35768,N_22061,N_26520);
nor U35769 (N_35769,N_24025,N_21274);
xor U35770 (N_35770,N_27870,N_21347);
and U35771 (N_35771,N_22497,N_25887);
nand U35772 (N_35772,N_22369,N_28698);
nand U35773 (N_35773,N_24659,N_23687);
or U35774 (N_35774,N_25255,N_27149);
xor U35775 (N_35775,N_25083,N_29265);
nand U35776 (N_35776,N_26447,N_28669);
nand U35777 (N_35777,N_23132,N_29911);
or U35778 (N_35778,N_20339,N_21529);
nand U35779 (N_35779,N_26270,N_26582);
or U35780 (N_35780,N_28272,N_28706);
nor U35781 (N_35781,N_27758,N_24064);
nor U35782 (N_35782,N_26479,N_25609);
nor U35783 (N_35783,N_26973,N_27247);
and U35784 (N_35784,N_22174,N_29617);
nand U35785 (N_35785,N_25037,N_21823);
nor U35786 (N_35786,N_25927,N_23700);
nand U35787 (N_35787,N_24378,N_20661);
nand U35788 (N_35788,N_25114,N_27926);
nand U35789 (N_35789,N_25245,N_21075);
and U35790 (N_35790,N_20870,N_28555);
and U35791 (N_35791,N_27968,N_27241);
nor U35792 (N_35792,N_24832,N_29849);
xnor U35793 (N_35793,N_26417,N_23682);
nor U35794 (N_35794,N_27603,N_20995);
nor U35795 (N_35795,N_29717,N_22823);
nand U35796 (N_35796,N_28973,N_24029);
nand U35797 (N_35797,N_26088,N_22029);
or U35798 (N_35798,N_23640,N_24086);
nand U35799 (N_35799,N_24943,N_24577);
xnor U35800 (N_35800,N_21046,N_25863);
xnor U35801 (N_35801,N_22700,N_22805);
nand U35802 (N_35802,N_23392,N_23644);
and U35803 (N_35803,N_24258,N_29219);
nor U35804 (N_35804,N_25216,N_23957);
xor U35805 (N_35805,N_22098,N_21368);
xor U35806 (N_35806,N_26623,N_26569);
xor U35807 (N_35807,N_22040,N_22778);
nand U35808 (N_35808,N_25899,N_28294);
nand U35809 (N_35809,N_25189,N_29447);
xor U35810 (N_35810,N_27952,N_25463);
or U35811 (N_35811,N_20532,N_28236);
xnor U35812 (N_35812,N_27549,N_26824);
nand U35813 (N_35813,N_23469,N_21017);
and U35814 (N_35814,N_27627,N_29799);
nand U35815 (N_35815,N_26069,N_27247);
nand U35816 (N_35816,N_21867,N_24343);
and U35817 (N_35817,N_24164,N_23657);
nand U35818 (N_35818,N_27294,N_28264);
xor U35819 (N_35819,N_28385,N_22644);
nand U35820 (N_35820,N_20750,N_23909);
nor U35821 (N_35821,N_24766,N_27448);
nand U35822 (N_35822,N_24851,N_21651);
xnor U35823 (N_35823,N_28096,N_28831);
nor U35824 (N_35824,N_29046,N_22222);
nor U35825 (N_35825,N_26452,N_27592);
and U35826 (N_35826,N_20569,N_26035);
and U35827 (N_35827,N_28805,N_20821);
nor U35828 (N_35828,N_26936,N_22258);
and U35829 (N_35829,N_22361,N_25261);
and U35830 (N_35830,N_28511,N_25016);
or U35831 (N_35831,N_25989,N_25810);
xnor U35832 (N_35832,N_26524,N_27507);
or U35833 (N_35833,N_27169,N_22283);
or U35834 (N_35834,N_23440,N_22291);
or U35835 (N_35835,N_21933,N_24958);
or U35836 (N_35836,N_23099,N_20984);
and U35837 (N_35837,N_22040,N_25111);
xor U35838 (N_35838,N_21704,N_26195);
and U35839 (N_35839,N_23933,N_28755);
and U35840 (N_35840,N_21845,N_26907);
and U35841 (N_35841,N_25462,N_27648);
xor U35842 (N_35842,N_26149,N_24310);
or U35843 (N_35843,N_26631,N_29874);
or U35844 (N_35844,N_26817,N_27507);
xnor U35845 (N_35845,N_28287,N_22367);
nor U35846 (N_35846,N_28158,N_24510);
and U35847 (N_35847,N_28539,N_22093);
or U35848 (N_35848,N_27978,N_22178);
nand U35849 (N_35849,N_25290,N_22516);
nor U35850 (N_35850,N_28508,N_29089);
nand U35851 (N_35851,N_20667,N_29545);
xor U35852 (N_35852,N_27112,N_27216);
nor U35853 (N_35853,N_28000,N_21649);
and U35854 (N_35854,N_29750,N_27553);
xor U35855 (N_35855,N_28503,N_20172);
and U35856 (N_35856,N_29565,N_26374);
and U35857 (N_35857,N_26121,N_21841);
nor U35858 (N_35858,N_23127,N_28538);
nand U35859 (N_35859,N_22274,N_21713);
xor U35860 (N_35860,N_29244,N_26674);
nor U35861 (N_35861,N_26976,N_21539);
nand U35862 (N_35862,N_27555,N_25616);
and U35863 (N_35863,N_20724,N_26842);
nand U35864 (N_35864,N_24692,N_22719);
nand U35865 (N_35865,N_28898,N_23615);
nor U35866 (N_35866,N_28590,N_28316);
and U35867 (N_35867,N_23152,N_20685);
nor U35868 (N_35868,N_27911,N_29099);
nor U35869 (N_35869,N_23195,N_28915);
xnor U35870 (N_35870,N_26049,N_22195);
or U35871 (N_35871,N_27520,N_23560);
or U35872 (N_35872,N_23849,N_21671);
nor U35873 (N_35873,N_22175,N_28206);
xnor U35874 (N_35874,N_22574,N_28721);
nor U35875 (N_35875,N_29642,N_23203);
and U35876 (N_35876,N_27944,N_22919);
and U35877 (N_35877,N_20695,N_26143);
or U35878 (N_35878,N_28716,N_26075);
or U35879 (N_35879,N_24711,N_29022);
nor U35880 (N_35880,N_26626,N_29888);
nor U35881 (N_35881,N_21713,N_27699);
and U35882 (N_35882,N_25737,N_22737);
nor U35883 (N_35883,N_26279,N_21988);
xor U35884 (N_35884,N_22564,N_24558);
nor U35885 (N_35885,N_28518,N_25471);
or U35886 (N_35886,N_28408,N_24833);
nor U35887 (N_35887,N_27850,N_22737);
or U35888 (N_35888,N_20514,N_26739);
nor U35889 (N_35889,N_22407,N_29568);
xor U35890 (N_35890,N_28734,N_23171);
xnor U35891 (N_35891,N_21182,N_25077);
nor U35892 (N_35892,N_21821,N_29731);
or U35893 (N_35893,N_27810,N_29362);
and U35894 (N_35894,N_21211,N_27344);
or U35895 (N_35895,N_27430,N_25609);
xnor U35896 (N_35896,N_20684,N_24473);
nand U35897 (N_35897,N_29935,N_27972);
nor U35898 (N_35898,N_22700,N_26346);
and U35899 (N_35899,N_20668,N_21630);
or U35900 (N_35900,N_26830,N_28890);
or U35901 (N_35901,N_22968,N_29248);
nand U35902 (N_35902,N_26258,N_22335);
and U35903 (N_35903,N_28985,N_23862);
xnor U35904 (N_35904,N_21300,N_28079);
nor U35905 (N_35905,N_27378,N_24929);
and U35906 (N_35906,N_27202,N_26629);
and U35907 (N_35907,N_29821,N_27637);
nand U35908 (N_35908,N_25412,N_25109);
nand U35909 (N_35909,N_25730,N_23026);
and U35910 (N_35910,N_21897,N_26057);
nand U35911 (N_35911,N_24295,N_27752);
and U35912 (N_35912,N_26447,N_22682);
nor U35913 (N_35913,N_24809,N_21574);
nor U35914 (N_35914,N_24742,N_28605);
and U35915 (N_35915,N_21089,N_29844);
nand U35916 (N_35916,N_22989,N_25015);
nor U35917 (N_35917,N_29438,N_22151);
or U35918 (N_35918,N_25692,N_29286);
and U35919 (N_35919,N_23789,N_23379);
and U35920 (N_35920,N_29856,N_25431);
nand U35921 (N_35921,N_22161,N_28347);
and U35922 (N_35922,N_22724,N_25786);
and U35923 (N_35923,N_20992,N_23611);
or U35924 (N_35924,N_21313,N_21578);
nand U35925 (N_35925,N_22596,N_21678);
and U35926 (N_35926,N_26203,N_24172);
xnor U35927 (N_35927,N_21981,N_25334);
or U35928 (N_35928,N_20045,N_25243);
nor U35929 (N_35929,N_28209,N_28789);
or U35930 (N_35930,N_29368,N_28456);
or U35931 (N_35931,N_24236,N_20852);
or U35932 (N_35932,N_21079,N_25670);
nor U35933 (N_35933,N_26035,N_24750);
xor U35934 (N_35934,N_22792,N_29438);
or U35935 (N_35935,N_29600,N_29122);
or U35936 (N_35936,N_27343,N_27027);
or U35937 (N_35937,N_21700,N_24562);
nand U35938 (N_35938,N_26887,N_22925);
and U35939 (N_35939,N_23971,N_23724);
nand U35940 (N_35940,N_20769,N_25043);
nor U35941 (N_35941,N_24224,N_22022);
nor U35942 (N_35942,N_25815,N_23255);
nand U35943 (N_35943,N_29449,N_27910);
xnor U35944 (N_35944,N_22833,N_24153);
nand U35945 (N_35945,N_24607,N_27739);
nor U35946 (N_35946,N_22288,N_22029);
nand U35947 (N_35947,N_20202,N_25067);
nor U35948 (N_35948,N_24091,N_26419);
xor U35949 (N_35949,N_27322,N_22629);
nor U35950 (N_35950,N_20323,N_26334);
nand U35951 (N_35951,N_26886,N_27926);
and U35952 (N_35952,N_29936,N_23651);
or U35953 (N_35953,N_21601,N_25686);
nand U35954 (N_35954,N_21209,N_28945);
xnor U35955 (N_35955,N_28086,N_23727);
xor U35956 (N_35956,N_28456,N_23622);
or U35957 (N_35957,N_24997,N_25146);
nor U35958 (N_35958,N_29384,N_29421);
xnor U35959 (N_35959,N_23484,N_23935);
or U35960 (N_35960,N_28080,N_22499);
nor U35961 (N_35961,N_21093,N_20406);
xor U35962 (N_35962,N_29748,N_27734);
and U35963 (N_35963,N_24275,N_22214);
and U35964 (N_35964,N_21145,N_22849);
nand U35965 (N_35965,N_21093,N_28964);
nand U35966 (N_35966,N_24706,N_27445);
nand U35967 (N_35967,N_23291,N_20462);
xnor U35968 (N_35968,N_24528,N_29180);
or U35969 (N_35969,N_20018,N_25336);
xor U35970 (N_35970,N_21145,N_26672);
nor U35971 (N_35971,N_24239,N_22541);
nor U35972 (N_35972,N_23113,N_27918);
and U35973 (N_35973,N_24571,N_23302);
or U35974 (N_35974,N_25399,N_24396);
nand U35975 (N_35975,N_28301,N_21258);
nand U35976 (N_35976,N_20015,N_23713);
or U35977 (N_35977,N_20787,N_24850);
or U35978 (N_35978,N_23299,N_29245);
xnor U35979 (N_35979,N_20862,N_22052);
nand U35980 (N_35980,N_27758,N_27336);
and U35981 (N_35981,N_27315,N_27311);
nor U35982 (N_35982,N_26328,N_28730);
and U35983 (N_35983,N_22147,N_23480);
or U35984 (N_35984,N_25235,N_21561);
nor U35985 (N_35985,N_20682,N_26107);
nand U35986 (N_35986,N_24780,N_23999);
or U35987 (N_35987,N_24027,N_25745);
nor U35988 (N_35988,N_20965,N_28549);
nor U35989 (N_35989,N_29077,N_27922);
and U35990 (N_35990,N_25232,N_27846);
nand U35991 (N_35991,N_21849,N_23231);
nand U35992 (N_35992,N_21697,N_22510);
and U35993 (N_35993,N_20582,N_22068);
nor U35994 (N_35994,N_24789,N_22032);
and U35995 (N_35995,N_23401,N_25634);
nand U35996 (N_35996,N_29773,N_24770);
nand U35997 (N_35997,N_20667,N_24813);
or U35998 (N_35998,N_28852,N_20438);
xor U35999 (N_35999,N_29197,N_20897);
nor U36000 (N_36000,N_21805,N_22890);
or U36001 (N_36001,N_28602,N_22114);
or U36002 (N_36002,N_22630,N_28080);
or U36003 (N_36003,N_26284,N_24130);
or U36004 (N_36004,N_22016,N_20089);
and U36005 (N_36005,N_23711,N_24227);
nor U36006 (N_36006,N_23774,N_28055);
and U36007 (N_36007,N_26678,N_21219);
xor U36008 (N_36008,N_25760,N_25587);
nand U36009 (N_36009,N_21560,N_26696);
nand U36010 (N_36010,N_28545,N_27272);
or U36011 (N_36011,N_21598,N_24368);
or U36012 (N_36012,N_28308,N_20745);
nand U36013 (N_36013,N_29884,N_26097);
and U36014 (N_36014,N_25371,N_27351);
and U36015 (N_36015,N_27641,N_23137);
or U36016 (N_36016,N_24901,N_23161);
and U36017 (N_36017,N_24380,N_23410);
or U36018 (N_36018,N_23246,N_21777);
nor U36019 (N_36019,N_21144,N_21093);
nor U36020 (N_36020,N_20553,N_24511);
nor U36021 (N_36021,N_20827,N_23677);
or U36022 (N_36022,N_20215,N_22599);
nor U36023 (N_36023,N_27087,N_20030);
or U36024 (N_36024,N_22882,N_26371);
nor U36025 (N_36025,N_25947,N_21845);
and U36026 (N_36026,N_20270,N_23562);
or U36027 (N_36027,N_26014,N_21936);
xnor U36028 (N_36028,N_26042,N_25762);
or U36029 (N_36029,N_22366,N_22667);
or U36030 (N_36030,N_21890,N_29191);
and U36031 (N_36031,N_20134,N_24835);
nand U36032 (N_36032,N_23082,N_26044);
and U36033 (N_36033,N_29562,N_26130);
nand U36034 (N_36034,N_28080,N_25049);
nand U36035 (N_36035,N_23788,N_23526);
or U36036 (N_36036,N_23131,N_22906);
nor U36037 (N_36037,N_29506,N_22437);
xor U36038 (N_36038,N_20915,N_27199);
or U36039 (N_36039,N_29654,N_29346);
nor U36040 (N_36040,N_28175,N_29855);
nand U36041 (N_36041,N_22719,N_24082);
or U36042 (N_36042,N_20953,N_28318);
or U36043 (N_36043,N_27986,N_20131);
and U36044 (N_36044,N_22853,N_29359);
nand U36045 (N_36045,N_21568,N_28527);
and U36046 (N_36046,N_28089,N_23997);
and U36047 (N_36047,N_24178,N_22499);
nor U36048 (N_36048,N_21105,N_24425);
nor U36049 (N_36049,N_23459,N_26494);
nor U36050 (N_36050,N_26494,N_24980);
nand U36051 (N_36051,N_21651,N_25231);
or U36052 (N_36052,N_27447,N_25454);
xnor U36053 (N_36053,N_26698,N_28700);
nand U36054 (N_36054,N_20822,N_27507);
xnor U36055 (N_36055,N_20258,N_29265);
nor U36056 (N_36056,N_27765,N_24433);
nand U36057 (N_36057,N_29957,N_27371);
or U36058 (N_36058,N_21747,N_27950);
nand U36059 (N_36059,N_25985,N_25644);
nand U36060 (N_36060,N_27290,N_27259);
or U36061 (N_36061,N_27900,N_20984);
and U36062 (N_36062,N_27855,N_26751);
or U36063 (N_36063,N_26452,N_27566);
xor U36064 (N_36064,N_22203,N_23746);
nor U36065 (N_36065,N_28781,N_20545);
nor U36066 (N_36066,N_27978,N_21730);
and U36067 (N_36067,N_26339,N_27584);
nor U36068 (N_36068,N_29639,N_28047);
xor U36069 (N_36069,N_23783,N_20334);
nor U36070 (N_36070,N_25862,N_29105);
xor U36071 (N_36071,N_25199,N_23289);
and U36072 (N_36072,N_20673,N_24773);
nand U36073 (N_36073,N_25876,N_27748);
and U36074 (N_36074,N_21198,N_21176);
xor U36075 (N_36075,N_24994,N_21319);
nand U36076 (N_36076,N_21292,N_24383);
xor U36077 (N_36077,N_23144,N_28164);
xor U36078 (N_36078,N_22762,N_24248);
and U36079 (N_36079,N_24103,N_20616);
and U36080 (N_36080,N_26878,N_29088);
nor U36081 (N_36081,N_26542,N_22894);
and U36082 (N_36082,N_22985,N_21150);
nand U36083 (N_36083,N_22544,N_21148);
xnor U36084 (N_36084,N_29736,N_29828);
xor U36085 (N_36085,N_23717,N_24179);
xnor U36086 (N_36086,N_26415,N_26669);
or U36087 (N_36087,N_29116,N_27548);
nand U36088 (N_36088,N_20035,N_25389);
nand U36089 (N_36089,N_25250,N_26256);
and U36090 (N_36090,N_23443,N_27399);
and U36091 (N_36091,N_24265,N_29864);
xnor U36092 (N_36092,N_27464,N_23623);
nor U36093 (N_36093,N_27513,N_23345);
xnor U36094 (N_36094,N_24659,N_24793);
nand U36095 (N_36095,N_29679,N_21351);
nor U36096 (N_36096,N_22144,N_25253);
nand U36097 (N_36097,N_23787,N_23079);
xnor U36098 (N_36098,N_25697,N_29536);
nand U36099 (N_36099,N_27859,N_23015);
nor U36100 (N_36100,N_28830,N_22683);
xor U36101 (N_36101,N_28167,N_20006);
or U36102 (N_36102,N_28823,N_28836);
or U36103 (N_36103,N_25517,N_24257);
xnor U36104 (N_36104,N_22697,N_24412);
and U36105 (N_36105,N_21375,N_22424);
or U36106 (N_36106,N_20283,N_28078);
or U36107 (N_36107,N_28781,N_26246);
nand U36108 (N_36108,N_22175,N_27040);
or U36109 (N_36109,N_27565,N_23258);
nand U36110 (N_36110,N_23390,N_24020);
xor U36111 (N_36111,N_29263,N_21484);
or U36112 (N_36112,N_22656,N_26889);
xor U36113 (N_36113,N_28502,N_22667);
or U36114 (N_36114,N_28739,N_28439);
xnor U36115 (N_36115,N_22379,N_26316);
and U36116 (N_36116,N_21946,N_21723);
and U36117 (N_36117,N_24681,N_21769);
nand U36118 (N_36118,N_21797,N_23749);
nor U36119 (N_36119,N_23005,N_22844);
nor U36120 (N_36120,N_29188,N_26240);
nor U36121 (N_36121,N_20110,N_20222);
nand U36122 (N_36122,N_27078,N_28614);
or U36123 (N_36123,N_25277,N_21137);
xnor U36124 (N_36124,N_26835,N_22998);
nand U36125 (N_36125,N_21634,N_25309);
xor U36126 (N_36126,N_26732,N_25542);
or U36127 (N_36127,N_24878,N_26678);
nor U36128 (N_36128,N_29102,N_27662);
nand U36129 (N_36129,N_23569,N_27800);
xnor U36130 (N_36130,N_27553,N_28203);
and U36131 (N_36131,N_28987,N_22138);
nor U36132 (N_36132,N_27969,N_22840);
or U36133 (N_36133,N_26965,N_23794);
nand U36134 (N_36134,N_28999,N_20634);
or U36135 (N_36135,N_26062,N_27368);
and U36136 (N_36136,N_21986,N_28559);
and U36137 (N_36137,N_27201,N_24604);
nand U36138 (N_36138,N_27354,N_26537);
and U36139 (N_36139,N_27715,N_23879);
nor U36140 (N_36140,N_24947,N_21641);
xnor U36141 (N_36141,N_28703,N_23952);
or U36142 (N_36142,N_29620,N_28301);
xor U36143 (N_36143,N_27826,N_24889);
nor U36144 (N_36144,N_26152,N_28010);
or U36145 (N_36145,N_25961,N_25348);
nand U36146 (N_36146,N_29853,N_28117);
and U36147 (N_36147,N_26150,N_26747);
nand U36148 (N_36148,N_24775,N_21213);
or U36149 (N_36149,N_27873,N_27558);
or U36150 (N_36150,N_25042,N_22278);
xnor U36151 (N_36151,N_26781,N_27178);
nand U36152 (N_36152,N_27874,N_27096);
and U36153 (N_36153,N_24864,N_25644);
nand U36154 (N_36154,N_25599,N_25461);
xor U36155 (N_36155,N_27613,N_20270);
nand U36156 (N_36156,N_22611,N_28616);
xor U36157 (N_36157,N_23567,N_27561);
or U36158 (N_36158,N_23338,N_20683);
and U36159 (N_36159,N_27485,N_23041);
or U36160 (N_36160,N_26146,N_22646);
nand U36161 (N_36161,N_29523,N_28220);
nor U36162 (N_36162,N_24321,N_22605);
nand U36163 (N_36163,N_23517,N_29762);
nand U36164 (N_36164,N_29799,N_21542);
xor U36165 (N_36165,N_23638,N_21489);
nand U36166 (N_36166,N_24810,N_26543);
nor U36167 (N_36167,N_25636,N_26817);
nor U36168 (N_36168,N_25079,N_27698);
nand U36169 (N_36169,N_23484,N_20482);
nor U36170 (N_36170,N_20461,N_21170);
nor U36171 (N_36171,N_28178,N_21419);
or U36172 (N_36172,N_22105,N_25871);
or U36173 (N_36173,N_21666,N_21898);
nand U36174 (N_36174,N_20215,N_22261);
or U36175 (N_36175,N_22187,N_25839);
nand U36176 (N_36176,N_21829,N_21271);
nand U36177 (N_36177,N_27207,N_22345);
or U36178 (N_36178,N_23998,N_25843);
nor U36179 (N_36179,N_23315,N_20588);
or U36180 (N_36180,N_26136,N_26033);
or U36181 (N_36181,N_23797,N_23480);
nand U36182 (N_36182,N_29216,N_24021);
nor U36183 (N_36183,N_25647,N_21359);
and U36184 (N_36184,N_25696,N_20729);
or U36185 (N_36185,N_22237,N_22271);
or U36186 (N_36186,N_21746,N_21311);
xnor U36187 (N_36187,N_25262,N_21672);
or U36188 (N_36188,N_26125,N_28479);
xnor U36189 (N_36189,N_27016,N_23909);
or U36190 (N_36190,N_24854,N_26940);
nor U36191 (N_36191,N_24388,N_20181);
nand U36192 (N_36192,N_29531,N_25994);
or U36193 (N_36193,N_26918,N_21442);
nor U36194 (N_36194,N_27157,N_26271);
nor U36195 (N_36195,N_28712,N_26707);
or U36196 (N_36196,N_25534,N_22976);
or U36197 (N_36197,N_21351,N_21786);
and U36198 (N_36198,N_22988,N_23091);
nand U36199 (N_36199,N_28419,N_29568);
nor U36200 (N_36200,N_21733,N_20693);
xor U36201 (N_36201,N_28602,N_22874);
and U36202 (N_36202,N_25095,N_25269);
or U36203 (N_36203,N_23315,N_24424);
nor U36204 (N_36204,N_24058,N_22750);
and U36205 (N_36205,N_20083,N_21997);
nor U36206 (N_36206,N_22191,N_22741);
nand U36207 (N_36207,N_24716,N_28699);
and U36208 (N_36208,N_29922,N_21069);
xnor U36209 (N_36209,N_23255,N_20990);
nor U36210 (N_36210,N_21630,N_22858);
and U36211 (N_36211,N_20297,N_20370);
nand U36212 (N_36212,N_21143,N_25463);
nor U36213 (N_36213,N_25875,N_26665);
and U36214 (N_36214,N_27871,N_25605);
nand U36215 (N_36215,N_28696,N_23768);
nand U36216 (N_36216,N_25839,N_20125);
or U36217 (N_36217,N_23086,N_25859);
or U36218 (N_36218,N_24218,N_25768);
or U36219 (N_36219,N_25728,N_24251);
nand U36220 (N_36220,N_22952,N_29328);
or U36221 (N_36221,N_21535,N_24522);
or U36222 (N_36222,N_29491,N_22990);
and U36223 (N_36223,N_26072,N_29702);
xor U36224 (N_36224,N_28703,N_21765);
nor U36225 (N_36225,N_24226,N_22207);
xnor U36226 (N_36226,N_23322,N_21852);
nor U36227 (N_36227,N_27243,N_21565);
nor U36228 (N_36228,N_23589,N_24867);
and U36229 (N_36229,N_25984,N_27207);
xnor U36230 (N_36230,N_23717,N_24763);
xnor U36231 (N_36231,N_25996,N_25229);
nor U36232 (N_36232,N_24896,N_26842);
xnor U36233 (N_36233,N_29809,N_27883);
nor U36234 (N_36234,N_26049,N_22397);
and U36235 (N_36235,N_26031,N_27220);
or U36236 (N_36236,N_26479,N_26661);
nor U36237 (N_36237,N_20970,N_22560);
xnor U36238 (N_36238,N_22924,N_22842);
and U36239 (N_36239,N_23863,N_29798);
and U36240 (N_36240,N_28796,N_25701);
nand U36241 (N_36241,N_28561,N_25579);
nand U36242 (N_36242,N_28179,N_25100);
and U36243 (N_36243,N_27586,N_23483);
and U36244 (N_36244,N_24886,N_29632);
nand U36245 (N_36245,N_21252,N_26714);
or U36246 (N_36246,N_26768,N_21230);
xor U36247 (N_36247,N_26406,N_20633);
nor U36248 (N_36248,N_23758,N_29441);
or U36249 (N_36249,N_28810,N_20812);
nor U36250 (N_36250,N_21534,N_24698);
nor U36251 (N_36251,N_28023,N_28067);
and U36252 (N_36252,N_29161,N_27734);
and U36253 (N_36253,N_21649,N_24718);
nand U36254 (N_36254,N_27242,N_24497);
xor U36255 (N_36255,N_20627,N_27478);
nand U36256 (N_36256,N_21635,N_21555);
or U36257 (N_36257,N_23111,N_21038);
nand U36258 (N_36258,N_25765,N_25578);
or U36259 (N_36259,N_20998,N_26654);
nand U36260 (N_36260,N_28553,N_29995);
and U36261 (N_36261,N_25742,N_25319);
nand U36262 (N_36262,N_20022,N_27430);
or U36263 (N_36263,N_27533,N_26357);
nand U36264 (N_36264,N_20403,N_24190);
nor U36265 (N_36265,N_23872,N_26844);
nand U36266 (N_36266,N_27829,N_21932);
nor U36267 (N_36267,N_23164,N_24304);
xor U36268 (N_36268,N_29822,N_25048);
nand U36269 (N_36269,N_21374,N_22629);
xor U36270 (N_36270,N_28812,N_23981);
nand U36271 (N_36271,N_27865,N_21496);
nor U36272 (N_36272,N_21565,N_23254);
nor U36273 (N_36273,N_23169,N_20154);
and U36274 (N_36274,N_27259,N_24506);
nor U36275 (N_36275,N_29641,N_29751);
and U36276 (N_36276,N_25494,N_26871);
or U36277 (N_36277,N_20442,N_21285);
xor U36278 (N_36278,N_28766,N_22256);
or U36279 (N_36279,N_20595,N_29985);
xor U36280 (N_36280,N_26302,N_27155);
nand U36281 (N_36281,N_22562,N_27589);
xnor U36282 (N_36282,N_27273,N_20784);
nor U36283 (N_36283,N_26426,N_24087);
nor U36284 (N_36284,N_28530,N_20439);
nand U36285 (N_36285,N_22887,N_27840);
xnor U36286 (N_36286,N_23061,N_29922);
nor U36287 (N_36287,N_25336,N_26804);
nand U36288 (N_36288,N_20581,N_24815);
nand U36289 (N_36289,N_22510,N_25331);
nor U36290 (N_36290,N_28923,N_29428);
or U36291 (N_36291,N_29010,N_28493);
or U36292 (N_36292,N_21558,N_22232);
nand U36293 (N_36293,N_20847,N_23518);
nand U36294 (N_36294,N_24227,N_25661);
xnor U36295 (N_36295,N_24916,N_23970);
xnor U36296 (N_36296,N_23080,N_29608);
nor U36297 (N_36297,N_27574,N_24391);
or U36298 (N_36298,N_25081,N_28050);
nor U36299 (N_36299,N_29712,N_27884);
xnor U36300 (N_36300,N_21632,N_28253);
or U36301 (N_36301,N_25429,N_22918);
and U36302 (N_36302,N_27555,N_25480);
and U36303 (N_36303,N_28000,N_20438);
nor U36304 (N_36304,N_22179,N_22171);
or U36305 (N_36305,N_24632,N_22422);
or U36306 (N_36306,N_25373,N_25534);
xnor U36307 (N_36307,N_25886,N_28060);
nand U36308 (N_36308,N_25997,N_20460);
nor U36309 (N_36309,N_28438,N_27283);
nand U36310 (N_36310,N_24821,N_22808);
and U36311 (N_36311,N_22168,N_21994);
and U36312 (N_36312,N_20627,N_27844);
nand U36313 (N_36313,N_26819,N_22882);
and U36314 (N_36314,N_22763,N_20402);
xor U36315 (N_36315,N_21921,N_23438);
and U36316 (N_36316,N_28146,N_25630);
nor U36317 (N_36317,N_24545,N_26807);
xnor U36318 (N_36318,N_26504,N_22748);
xnor U36319 (N_36319,N_25698,N_26270);
xor U36320 (N_36320,N_21819,N_25466);
or U36321 (N_36321,N_22936,N_20764);
nor U36322 (N_36322,N_22937,N_28660);
and U36323 (N_36323,N_26143,N_26166);
or U36324 (N_36324,N_29972,N_27849);
xnor U36325 (N_36325,N_26825,N_25311);
nor U36326 (N_36326,N_20686,N_29431);
and U36327 (N_36327,N_28634,N_29573);
or U36328 (N_36328,N_27879,N_28424);
nor U36329 (N_36329,N_21335,N_23401);
nor U36330 (N_36330,N_28175,N_23623);
nor U36331 (N_36331,N_26244,N_27130);
or U36332 (N_36332,N_23625,N_24759);
or U36333 (N_36333,N_27400,N_24365);
xor U36334 (N_36334,N_29233,N_23471);
nand U36335 (N_36335,N_25220,N_24003);
or U36336 (N_36336,N_23833,N_29414);
or U36337 (N_36337,N_23744,N_20434);
xor U36338 (N_36338,N_29640,N_20278);
xnor U36339 (N_36339,N_22554,N_27651);
and U36340 (N_36340,N_23225,N_23523);
nand U36341 (N_36341,N_21362,N_21374);
nand U36342 (N_36342,N_28269,N_21106);
nand U36343 (N_36343,N_24173,N_22197);
xnor U36344 (N_36344,N_28696,N_22001);
nor U36345 (N_36345,N_23906,N_20161);
nor U36346 (N_36346,N_26542,N_23749);
nand U36347 (N_36347,N_27559,N_26668);
or U36348 (N_36348,N_25470,N_24044);
xor U36349 (N_36349,N_21861,N_27608);
or U36350 (N_36350,N_25148,N_24573);
and U36351 (N_36351,N_26501,N_29450);
or U36352 (N_36352,N_25646,N_24445);
and U36353 (N_36353,N_27601,N_24775);
or U36354 (N_36354,N_24342,N_21749);
nor U36355 (N_36355,N_24779,N_27578);
or U36356 (N_36356,N_29597,N_28751);
and U36357 (N_36357,N_24357,N_26198);
nor U36358 (N_36358,N_23447,N_20568);
and U36359 (N_36359,N_21248,N_25480);
xnor U36360 (N_36360,N_26856,N_27443);
xnor U36361 (N_36361,N_29973,N_28257);
xnor U36362 (N_36362,N_22361,N_27857);
or U36363 (N_36363,N_27278,N_27646);
and U36364 (N_36364,N_28415,N_21176);
nand U36365 (N_36365,N_23358,N_29840);
nor U36366 (N_36366,N_22848,N_22890);
xor U36367 (N_36367,N_28242,N_29747);
xor U36368 (N_36368,N_23605,N_27209);
nor U36369 (N_36369,N_20165,N_24895);
nand U36370 (N_36370,N_28702,N_24008);
or U36371 (N_36371,N_26209,N_25515);
nand U36372 (N_36372,N_29510,N_22077);
and U36373 (N_36373,N_23189,N_21052);
xnor U36374 (N_36374,N_24797,N_23338);
xor U36375 (N_36375,N_24536,N_24653);
nor U36376 (N_36376,N_26387,N_24853);
and U36377 (N_36377,N_29867,N_20046);
nor U36378 (N_36378,N_23548,N_28116);
nor U36379 (N_36379,N_23877,N_22820);
xnor U36380 (N_36380,N_25503,N_29606);
or U36381 (N_36381,N_20341,N_26374);
nand U36382 (N_36382,N_20964,N_29043);
xor U36383 (N_36383,N_29842,N_23777);
xor U36384 (N_36384,N_21908,N_25889);
nor U36385 (N_36385,N_25572,N_27656);
xor U36386 (N_36386,N_23131,N_20823);
or U36387 (N_36387,N_22288,N_21523);
or U36388 (N_36388,N_28966,N_26664);
or U36389 (N_36389,N_29594,N_21124);
xor U36390 (N_36390,N_22085,N_24077);
and U36391 (N_36391,N_24020,N_29278);
and U36392 (N_36392,N_22436,N_27533);
or U36393 (N_36393,N_20728,N_29893);
nor U36394 (N_36394,N_25637,N_26669);
nand U36395 (N_36395,N_22361,N_20490);
nand U36396 (N_36396,N_28218,N_20133);
and U36397 (N_36397,N_27770,N_20697);
and U36398 (N_36398,N_24666,N_25595);
and U36399 (N_36399,N_24528,N_24049);
nor U36400 (N_36400,N_22668,N_27275);
xor U36401 (N_36401,N_21221,N_20548);
or U36402 (N_36402,N_20946,N_21016);
nor U36403 (N_36403,N_24831,N_25172);
nor U36404 (N_36404,N_21025,N_25482);
and U36405 (N_36405,N_24855,N_24617);
and U36406 (N_36406,N_25481,N_21679);
xor U36407 (N_36407,N_24533,N_27888);
nand U36408 (N_36408,N_21756,N_24052);
nor U36409 (N_36409,N_21452,N_24343);
nor U36410 (N_36410,N_24363,N_23079);
and U36411 (N_36411,N_27106,N_27783);
or U36412 (N_36412,N_28645,N_24433);
nor U36413 (N_36413,N_23514,N_28066);
or U36414 (N_36414,N_28200,N_24279);
nand U36415 (N_36415,N_29490,N_28180);
and U36416 (N_36416,N_28485,N_24075);
xor U36417 (N_36417,N_20003,N_27214);
xnor U36418 (N_36418,N_20606,N_23244);
or U36419 (N_36419,N_21217,N_23322);
xnor U36420 (N_36420,N_26540,N_24219);
or U36421 (N_36421,N_22599,N_20366);
and U36422 (N_36422,N_29673,N_22415);
xor U36423 (N_36423,N_25292,N_27711);
or U36424 (N_36424,N_27995,N_21785);
nand U36425 (N_36425,N_28055,N_20612);
nor U36426 (N_36426,N_27299,N_22610);
and U36427 (N_36427,N_27868,N_28334);
or U36428 (N_36428,N_24153,N_24911);
or U36429 (N_36429,N_24494,N_29573);
nor U36430 (N_36430,N_23283,N_27296);
nand U36431 (N_36431,N_24219,N_23594);
or U36432 (N_36432,N_22669,N_21513);
xnor U36433 (N_36433,N_22934,N_28688);
nor U36434 (N_36434,N_20735,N_22074);
xor U36435 (N_36435,N_24292,N_22762);
xor U36436 (N_36436,N_21998,N_26180);
or U36437 (N_36437,N_29832,N_24929);
nor U36438 (N_36438,N_24619,N_20090);
and U36439 (N_36439,N_29039,N_29385);
and U36440 (N_36440,N_20288,N_25328);
and U36441 (N_36441,N_29253,N_20398);
or U36442 (N_36442,N_24954,N_26014);
or U36443 (N_36443,N_27609,N_27790);
or U36444 (N_36444,N_28736,N_27319);
and U36445 (N_36445,N_25927,N_22938);
and U36446 (N_36446,N_20574,N_25324);
nand U36447 (N_36447,N_27147,N_27449);
and U36448 (N_36448,N_21833,N_23516);
and U36449 (N_36449,N_22909,N_23448);
and U36450 (N_36450,N_22621,N_20895);
or U36451 (N_36451,N_21016,N_25962);
xor U36452 (N_36452,N_29372,N_27479);
or U36453 (N_36453,N_26443,N_20618);
and U36454 (N_36454,N_28760,N_26814);
nand U36455 (N_36455,N_29742,N_28269);
and U36456 (N_36456,N_20201,N_26325);
nand U36457 (N_36457,N_21414,N_25392);
and U36458 (N_36458,N_24382,N_23380);
or U36459 (N_36459,N_29839,N_29001);
xor U36460 (N_36460,N_28720,N_27460);
or U36461 (N_36461,N_24575,N_21772);
or U36462 (N_36462,N_20959,N_27416);
xor U36463 (N_36463,N_23896,N_24458);
and U36464 (N_36464,N_26992,N_24499);
nor U36465 (N_36465,N_24753,N_26219);
nor U36466 (N_36466,N_26189,N_29703);
and U36467 (N_36467,N_20982,N_29642);
or U36468 (N_36468,N_20262,N_28156);
or U36469 (N_36469,N_20797,N_27077);
nand U36470 (N_36470,N_27803,N_26108);
nand U36471 (N_36471,N_29134,N_24266);
xor U36472 (N_36472,N_26956,N_26942);
nor U36473 (N_36473,N_28541,N_26987);
xor U36474 (N_36474,N_28367,N_29696);
xor U36475 (N_36475,N_26296,N_26074);
or U36476 (N_36476,N_21027,N_25549);
xnor U36477 (N_36477,N_20781,N_21864);
nand U36478 (N_36478,N_29923,N_23128);
and U36479 (N_36479,N_21896,N_20248);
or U36480 (N_36480,N_23709,N_22043);
xnor U36481 (N_36481,N_23158,N_27198);
nand U36482 (N_36482,N_23720,N_22131);
nand U36483 (N_36483,N_28303,N_23398);
nor U36484 (N_36484,N_21594,N_29519);
nor U36485 (N_36485,N_27019,N_22631);
or U36486 (N_36486,N_27525,N_29272);
xnor U36487 (N_36487,N_20009,N_21652);
or U36488 (N_36488,N_27510,N_25938);
and U36489 (N_36489,N_20892,N_22049);
nand U36490 (N_36490,N_20507,N_28326);
and U36491 (N_36491,N_23036,N_23312);
and U36492 (N_36492,N_28947,N_27767);
or U36493 (N_36493,N_23012,N_29964);
and U36494 (N_36494,N_24286,N_22750);
or U36495 (N_36495,N_27034,N_27075);
nand U36496 (N_36496,N_25922,N_29840);
xnor U36497 (N_36497,N_24616,N_27544);
nand U36498 (N_36498,N_27961,N_26473);
or U36499 (N_36499,N_29161,N_29620);
and U36500 (N_36500,N_22305,N_21020);
nor U36501 (N_36501,N_24629,N_29060);
xnor U36502 (N_36502,N_27747,N_29794);
nand U36503 (N_36503,N_25306,N_27742);
nand U36504 (N_36504,N_28688,N_20061);
and U36505 (N_36505,N_23050,N_20853);
xnor U36506 (N_36506,N_24340,N_24858);
nand U36507 (N_36507,N_24867,N_29314);
nand U36508 (N_36508,N_20629,N_21277);
and U36509 (N_36509,N_20046,N_22036);
nand U36510 (N_36510,N_26250,N_22971);
nor U36511 (N_36511,N_27598,N_23775);
nand U36512 (N_36512,N_20787,N_22219);
nor U36513 (N_36513,N_25694,N_29082);
and U36514 (N_36514,N_22519,N_25450);
nor U36515 (N_36515,N_21103,N_21128);
or U36516 (N_36516,N_28522,N_25420);
xnor U36517 (N_36517,N_20139,N_28936);
nand U36518 (N_36518,N_21829,N_29212);
or U36519 (N_36519,N_26477,N_29279);
nand U36520 (N_36520,N_28308,N_20132);
nand U36521 (N_36521,N_22246,N_21433);
nand U36522 (N_36522,N_24050,N_25693);
xnor U36523 (N_36523,N_22111,N_26003);
nor U36524 (N_36524,N_26868,N_24865);
xnor U36525 (N_36525,N_29751,N_24377);
and U36526 (N_36526,N_21438,N_22201);
xnor U36527 (N_36527,N_27157,N_21951);
xor U36528 (N_36528,N_26635,N_20790);
nand U36529 (N_36529,N_24901,N_27547);
or U36530 (N_36530,N_22174,N_23073);
or U36531 (N_36531,N_29031,N_22065);
nor U36532 (N_36532,N_28086,N_21353);
xnor U36533 (N_36533,N_23507,N_20764);
and U36534 (N_36534,N_24077,N_21682);
and U36535 (N_36535,N_25961,N_24915);
nor U36536 (N_36536,N_23328,N_21549);
and U36537 (N_36537,N_21157,N_29786);
nor U36538 (N_36538,N_24401,N_25091);
nor U36539 (N_36539,N_28475,N_26431);
nand U36540 (N_36540,N_28141,N_29251);
xnor U36541 (N_36541,N_27095,N_23415);
or U36542 (N_36542,N_22660,N_24814);
or U36543 (N_36543,N_27481,N_21120);
nand U36544 (N_36544,N_24935,N_24798);
xor U36545 (N_36545,N_28401,N_27258);
nand U36546 (N_36546,N_21699,N_27419);
and U36547 (N_36547,N_28810,N_25454);
or U36548 (N_36548,N_21726,N_20902);
nand U36549 (N_36549,N_23574,N_26476);
nand U36550 (N_36550,N_22376,N_27237);
or U36551 (N_36551,N_26971,N_25698);
xor U36552 (N_36552,N_29707,N_25166);
xnor U36553 (N_36553,N_20589,N_24000);
nand U36554 (N_36554,N_20542,N_27045);
or U36555 (N_36555,N_24994,N_21850);
xnor U36556 (N_36556,N_29476,N_29467);
nand U36557 (N_36557,N_24936,N_20098);
nor U36558 (N_36558,N_29136,N_29939);
and U36559 (N_36559,N_26176,N_22476);
or U36560 (N_36560,N_22935,N_22840);
and U36561 (N_36561,N_28868,N_23846);
xor U36562 (N_36562,N_27958,N_24695);
xor U36563 (N_36563,N_27180,N_26890);
nor U36564 (N_36564,N_20541,N_20870);
or U36565 (N_36565,N_23425,N_27459);
or U36566 (N_36566,N_21278,N_23792);
and U36567 (N_36567,N_23934,N_28783);
and U36568 (N_36568,N_23862,N_23963);
xor U36569 (N_36569,N_28711,N_25447);
nand U36570 (N_36570,N_27385,N_27645);
and U36571 (N_36571,N_25128,N_27913);
nor U36572 (N_36572,N_22902,N_25431);
nand U36573 (N_36573,N_25830,N_23848);
and U36574 (N_36574,N_29205,N_29440);
and U36575 (N_36575,N_27643,N_25441);
and U36576 (N_36576,N_27133,N_20894);
xnor U36577 (N_36577,N_24272,N_21586);
or U36578 (N_36578,N_22517,N_26358);
nand U36579 (N_36579,N_20824,N_22768);
or U36580 (N_36580,N_21216,N_22948);
nand U36581 (N_36581,N_24539,N_21431);
nor U36582 (N_36582,N_23609,N_22145);
xor U36583 (N_36583,N_22971,N_26942);
xor U36584 (N_36584,N_21969,N_24274);
or U36585 (N_36585,N_22711,N_21309);
and U36586 (N_36586,N_28873,N_20991);
nor U36587 (N_36587,N_25037,N_22767);
nor U36588 (N_36588,N_28857,N_22458);
xor U36589 (N_36589,N_27195,N_28686);
nor U36590 (N_36590,N_29680,N_21570);
xor U36591 (N_36591,N_26906,N_29998);
nor U36592 (N_36592,N_24601,N_24354);
nand U36593 (N_36593,N_23202,N_21996);
or U36594 (N_36594,N_21940,N_22184);
xnor U36595 (N_36595,N_20285,N_20232);
xnor U36596 (N_36596,N_24243,N_20548);
xor U36597 (N_36597,N_22499,N_26662);
or U36598 (N_36598,N_25117,N_21728);
or U36599 (N_36599,N_26566,N_22544);
nand U36600 (N_36600,N_22622,N_28922);
xor U36601 (N_36601,N_26045,N_21714);
nand U36602 (N_36602,N_29218,N_28088);
nor U36603 (N_36603,N_29923,N_20746);
nor U36604 (N_36604,N_26064,N_26579);
or U36605 (N_36605,N_23932,N_28330);
xnor U36606 (N_36606,N_26685,N_27654);
or U36607 (N_36607,N_21258,N_29585);
nor U36608 (N_36608,N_27547,N_27665);
or U36609 (N_36609,N_27242,N_20874);
nand U36610 (N_36610,N_23378,N_20111);
nand U36611 (N_36611,N_21875,N_24511);
nor U36612 (N_36612,N_22024,N_26193);
or U36613 (N_36613,N_24306,N_22690);
nor U36614 (N_36614,N_24312,N_21571);
nand U36615 (N_36615,N_21725,N_25114);
and U36616 (N_36616,N_21704,N_27890);
or U36617 (N_36617,N_23592,N_24927);
and U36618 (N_36618,N_22931,N_23593);
nand U36619 (N_36619,N_24012,N_24984);
xor U36620 (N_36620,N_21520,N_21948);
or U36621 (N_36621,N_20042,N_20767);
and U36622 (N_36622,N_24816,N_25561);
or U36623 (N_36623,N_24680,N_23312);
xnor U36624 (N_36624,N_23980,N_21626);
nor U36625 (N_36625,N_26728,N_25417);
nand U36626 (N_36626,N_26688,N_23831);
nor U36627 (N_36627,N_27660,N_20654);
xnor U36628 (N_36628,N_24506,N_21642);
and U36629 (N_36629,N_23253,N_20097);
xor U36630 (N_36630,N_25633,N_29107);
xnor U36631 (N_36631,N_21560,N_26172);
xnor U36632 (N_36632,N_25569,N_27915);
and U36633 (N_36633,N_26404,N_27735);
nor U36634 (N_36634,N_20249,N_22355);
nand U36635 (N_36635,N_25314,N_27937);
nand U36636 (N_36636,N_27817,N_20882);
nor U36637 (N_36637,N_27647,N_25913);
and U36638 (N_36638,N_20406,N_20357);
and U36639 (N_36639,N_25877,N_24303);
or U36640 (N_36640,N_21132,N_23748);
or U36641 (N_36641,N_23581,N_25836);
xor U36642 (N_36642,N_28352,N_27042);
nand U36643 (N_36643,N_27597,N_27204);
nor U36644 (N_36644,N_24489,N_23661);
xor U36645 (N_36645,N_27002,N_28399);
nor U36646 (N_36646,N_26470,N_21749);
or U36647 (N_36647,N_21523,N_25397);
xor U36648 (N_36648,N_24248,N_28582);
nand U36649 (N_36649,N_21097,N_28366);
nor U36650 (N_36650,N_23903,N_27495);
nand U36651 (N_36651,N_27432,N_21380);
xor U36652 (N_36652,N_23793,N_26227);
nor U36653 (N_36653,N_26897,N_26906);
or U36654 (N_36654,N_26220,N_28261);
or U36655 (N_36655,N_20165,N_27853);
nor U36656 (N_36656,N_25251,N_23109);
or U36657 (N_36657,N_27862,N_23703);
xor U36658 (N_36658,N_27434,N_21188);
and U36659 (N_36659,N_20171,N_23338);
nand U36660 (N_36660,N_20170,N_23940);
or U36661 (N_36661,N_24600,N_23515);
nand U36662 (N_36662,N_28266,N_20274);
and U36663 (N_36663,N_22508,N_27444);
xnor U36664 (N_36664,N_22169,N_21640);
nor U36665 (N_36665,N_27593,N_22805);
and U36666 (N_36666,N_26245,N_22311);
xnor U36667 (N_36667,N_26494,N_21309);
xor U36668 (N_36668,N_21457,N_29874);
nor U36669 (N_36669,N_29528,N_29849);
xor U36670 (N_36670,N_20213,N_24342);
nand U36671 (N_36671,N_26894,N_24552);
or U36672 (N_36672,N_26493,N_24970);
nor U36673 (N_36673,N_27976,N_23021);
xor U36674 (N_36674,N_25220,N_20188);
and U36675 (N_36675,N_29687,N_26078);
nand U36676 (N_36676,N_28566,N_27771);
nand U36677 (N_36677,N_21608,N_23819);
and U36678 (N_36678,N_23021,N_28724);
nor U36679 (N_36679,N_24433,N_29583);
or U36680 (N_36680,N_21204,N_24135);
or U36681 (N_36681,N_21243,N_25362);
and U36682 (N_36682,N_26245,N_29981);
nor U36683 (N_36683,N_20875,N_26051);
nor U36684 (N_36684,N_25578,N_22501);
or U36685 (N_36685,N_23480,N_24015);
nor U36686 (N_36686,N_29968,N_28831);
or U36687 (N_36687,N_29308,N_20090);
and U36688 (N_36688,N_27801,N_23517);
nor U36689 (N_36689,N_23564,N_28683);
and U36690 (N_36690,N_29081,N_26747);
and U36691 (N_36691,N_22594,N_21453);
nor U36692 (N_36692,N_23885,N_27142);
xor U36693 (N_36693,N_24750,N_28225);
nand U36694 (N_36694,N_23808,N_21766);
xnor U36695 (N_36695,N_23281,N_21596);
xor U36696 (N_36696,N_23479,N_21076);
nor U36697 (N_36697,N_26462,N_27150);
and U36698 (N_36698,N_27952,N_26618);
xnor U36699 (N_36699,N_27878,N_23129);
xor U36700 (N_36700,N_22600,N_27255);
and U36701 (N_36701,N_24356,N_29702);
and U36702 (N_36702,N_21731,N_27777);
xor U36703 (N_36703,N_22273,N_29076);
or U36704 (N_36704,N_25918,N_25916);
xnor U36705 (N_36705,N_21370,N_29624);
nand U36706 (N_36706,N_23491,N_25999);
xnor U36707 (N_36707,N_21784,N_22017);
nand U36708 (N_36708,N_28601,N_22209);
nor U36709 (N_36709,N_28000,N_28665);
or U36710 (N_36710,N_26670,N_23772);
or U36711 (N_36711,N_26004,N_26677);
xor U36712 (N_36712,N_25940,N_28118);
and U36713 (N_36713,N_27951,N_21364);
nand U36714 (N_36714,N_25016,N_26590);
nand U36715 (N_36715,N_21562,N_22468);
or U36716 (N_36716,N_21716,N_29404);
nor U36717 (N_36717,N_23135,N_26508);
and U36718 (N_36718,N_20469,N_21743);
xnor U36719 (N_36719,N_21663,N_22002);
and U36720 (N_36720,N_27943,N_22745);
and U36721 (N_36721,N_20455,N_27991);
xor U36722 (N_36722,N_25047,N_26251);
nor U36723 (N_36723,N_24542,N_25672);
xnor U36724 (N_36724,N_21664,N_24929);
nor U36725 (N_36725,N_20674,N_28303);
xor U36726 (N_36726,N_29153,N_25342);
nand U36727 (N_36727,N_28822,N_29340);
and U36728 (N_36728,N_28629,N_28217);
nand U36729 (N_36729,N_22896,N_24137);
nand U36730 (N_36730,N_26285,N_21314);
nand U36731 (N_36731,N_29919,N_26900);
and U36732 (N_36732,N_21569,N_29225);
xor U36733 (N_36733,N_25551,N_21434);
nand U36734 (N_36734,N_29083,N_21192);
nand U36735 (N_36735,N_26629,N_20436);
or U36736 (N_36736,N_25143,N_22448);
xnor U36737 (N_36737,N_29610,N_22747);
nor U36738 (N_36738,N_23584,N_21466);
nand U36739 (N_36739,N_28345,N_29160);
xor U36740 (N_36740,N_26707,N_20443);
xnor U36741 (N_36741,N_23422,N_22551);
nand U36742 (N_36742,N_23056,N_20198);
nand U36743 (N_36743,N_24684,N_22127);
nand U36744 (N_36744,N_21977,N_27734);
or U36745 (N_36745,N_22698,N_27249);
xnor U36746 (N_36746,N_25320,N_21731);
nand U36747 (N_36747,N_28199,N_25493);
xnor U36748 (N_36748,N_21760,N_21634);
nand U36749 (N_36749,N_24181,N_22620);
or U36750 (N_36750,N_23900,N_24830);
and U36751 (N_36751,N_21803,N_27324);
xnor U36752 (N_36752,N_29584,N_25438);
or U36753 (N_36753,N_23309,N_21806);
nor U36754 (N_36754,N_27554,N_23048);
xnor U36755 (N_36755,N_26983,N_21070);
and U36756 (N_36756,N_23526,N_29053);
and U36757 (N_36757,N_23325,N_25229);
nand U36758 (N_36758,N_25428,N_23217);
and U36759 (N_36759,N_22591,N_26442);
and U36760 (N_36760,N_20863,N_20099);
nand U36761 (N_36761,N_20206,N_20996);
or U36762 (N_36762,N_20708,N_24508);
nor U36763 (N_36763,N_27972,N_26556);
nand U36764 (N_36764,N_28972,N_28567);
nor U36765 (N_36765,N_23488,N_29605);
xor U36766 (N_36766,N_24848,N_28547);
or U36767 (N_36767,N_20589,N_26184);
and U36768 (N_36768,N_28784,N_23292);
or U36769 (N_36769,N_21660,N_28596);
nand U36770 (N_36770,N_28229,N_25250);
and U36771 (N_36771,N_22519,N_20093);
and U36772 (N_36772,N_21930,N_29703);
or U36773 (N_36773,N_20025,N_25268);
nand U36774 (N_36774,N_24847,N_22936);
xor U36775 (N_36775,N_27340,N_26665);
nor U36776 (N_36776,N_22631,N_20959);
and U36777 (N_36777,N_26523,N_27741);
xnor U36778 (N_36778,N_21731,N_23828);
xor U36779 (N_36779,N_28111,N_26257);
nor U36780 (N_36780,N_25271,N_25162);
xnor U36781 (N_36781,N_21211,N_21528);
xor U36782 (N_36782,N_24322,N_21465);
or U36783 (N_36783,N_24743,N_22905);
xnor U36784 (N_36784,N_23730,N_25541);
nor U36785 (N_36785,N_24485,N_23881);
xor U36786 (N_36786,N_29159,N_27865);
and U36787 (N_36787,N_27205,N_26707);
nor U36788 (N_36788,N_28864,N_28196);
nand U36789 (N_36789,N_25815,N_23003);
and U36790 (N_36790,N_27576,N_28824);
and U36791 (N_36791,N_21859,N_29566);
nor U36792 (N_36792,N_22858,N_21434);
xor U36793 (N_36793,N_21678,N_27957);
or U36794 (N_36794,N_29394,N_26683);
nor U36795 (N_36795,N_26496,N_20464);
nand U36796 (N_36796,N_27677,N_28678);
nor U36797 (N_36797,N_25327,N_24789);
nand U36798 (N_36798,N_22335,N_29592);
or U36799 (N_36799,N_26956,N_27197);
nor U36800 (N_36800,N_20252,N_29618);
xor U36801 (N_36801,N_29529,N_29371);
xnor U36802 (N_36802,N_23609,N_28158);
and U36803 (N_36803,N_28477,N_21312);
xor U36804 (N_36804,N_23508,N_25549);
or U36805 (N_36805,N_25954,N_27250);
and U36806 (N_36806,N_20139,N_21753);
or U36807 (N_36807,N_23518,N_22019);
nor U36808 (N_36808,N_23643,N_20452);
or U36809 (N_36809,N_23523,N_21954);
nor U36810 (N_36810,N_25843,N_24517);
xor U36811 (N_36811,N_28097,N_21026);
xnor U36812 (N_36812,N_25891,N_21993);
nand U36813 (N_36813,N_22531,N_27344);
or U36814 (N_36814,N_28082,N_22079);
nand U36815 (N_36815,N_24803,N_26276);
or U36816 (N_36816,N_23522,N_29085);
or U36817 (N_36817,N_28272,N_28225);
and U36818 (N_36818,N_20919,N_29320);
or U36819 (N_36819,N_25572,N_26822);
and U36820 (N_36820,N_22187,N_21282);
or U36821 (N_36821,N_21298,N_26258);
and U36822 (N_36822,N_23705,N_21079);
and U36823 (N_36823,N_21660,N_29427);
xnor U36824 (N_36824,N_25608,N_23651);
or U36825 (N_36825,N_29055,N_26265);
xnor U36826 (N_36826,N_24395,N_22966);
xor U36827 (N_36827,N_28965,N_20526);
nor U36828 (N_36828,N_26486,N_21956);
or U36829 (N_36829,N_25696,N_28431);
and U36830 (N_36830,N_27988,N_26440);
xnor U36831 (N_36831,N_23045,N_28648);
nand U36832 (N_36832,N_28779,N_26046);
nand U36833 (N_36833,N_25306,N_28144);
and U36834 (N_36834,N_20885,N_28859);
xor U36835 (N_36835,N_24958,N_24985);
or U36836 (N_36836,N_20323,N_25587);
xnor U36837 (N_36837,N_26970,N_21923);
and U36838 (N_36838,N_21734,N_20352);
or U36839 (N_36839,N_29738,N_21656);
and U36840 (N_36840,N_24826,N_21742);
xnor U36841 (N_36841,N_23364,N_29691);
nand U36842 (N_36842,N_22650,N_20540);
nor U36843 (N_36843,N_22234,N_27642);
and U36844 (N_36844,N_26292,N_27389);
or U36845 (N_36845,N_26905,N_28015);
nand U36846 (N_36846,N_24080,N_21741);
xnor U36847 (N_36847,N_29895,N_27547);
or U36848 (N_36848,N_24740,N_22948);
nor U36849 (N_36849,N_25600,N_20096);
and U36850 (N_36850,N_24907,N_26299);
nor U36851 (N_36851,N_22178,N_26568);
and U36852 (N_36852,N_26955,N_24170);
and U36853 (N_36853,N_25996,N_29528);
nand U36854 (N_36854,N_28088,N_24276);
nor U36855 (N_36855,N_25440,N_23576);
xor U36856 (N_36856,N_26993,N_26476);
xnor U36857 (N_36857,N_29614,N_22694);
nor U36858 (N_36858,N_20360,N_23975);
nand U36859 (N_36859,N_22057,N_28057);
nand U36860 (N_36860,N_23739,N_23108);
nor U36861 (N_36861,N_20651,N_26490);
xor U36862 (N_36862,N_29819,N_28728);
nand U36863 (N_36863,N_24272,N_21819);
or U36864 (N_36864,N_27906,N_21652);
and U36865 (N_36865,N_28307,N_24927);
and U36866 (N_36866,N_27743,N_24851);
xnor U36867 (N_36867,N_25650,N_24033);
nand U36868 (N_36868,N_29072,N_27546);
nor U36869 (N_36869,N_24975,N_29492);
nand U36870 (N_36870,N_20488,N_28627);
xnor U36871 (N_36871,N_22881,N_24168);
nand U36872 (N_36872,N_27353,N_25758);
nand U36873 (N_36873,N_22080,N_21826);
nand U36874 (N_36874,N_27389,N_27841);
nand U36875 (N_36875,N_29188,N_21873);
nor U36876 (N_36876,N_25059,N_23083);
nor U36877 (N_36877,N_29311,N_24215);
or U36878 (N_36878,N_25105,N_29760);
xnor U36879 (N_36879,N_22462,N_26307);
nand U36880 (N_36880,N_24870,N_26053);
nand U36881 (N_36881,N_26785,N_21491);
xnor U36882 (N_36882,N_21849,N_24195);
xnor U36883 (N_36883,N_28805,N_23450);
or U36884 (N_36884,N_28539,N_23113);
and U36885 (N_36885,N_28781,N_25391);
and U36886 (N_36886,N_29157,N_29759);
or U36887 (N_36887,N_22813,N_24432);
or U36888 (N_36888,N_29411,N_26408);
nand U36889 (N_36889,N_25685,N_23129);
or U36890 (N_36890,N_29475,N_24670);
nor U36891 (N_36891,N_21499,N_22201);
and U36892 (N_36892,N_21354,N_25234);
xor U36893 (N_36893,N_24759,N_26198);
nand U36894 (N_36894,N_29297,N_23884);
or U36895 (N_36895,N_23077,N_23720);
xor U36896 (N_36896,N_29418,N_27798);
nor U36897 (N_36897,N_24578,N_23447);
nand U36898 (N_36898,N_28735,N_28212);
xor U36899 (N_36899,N_27472,N_26181);
nor U36900 (N_36900,N_28453,N_28066);
and U36901 (N_36901,N_21489,N_24862);
nand U36902 (N_36902,N_25859,N_29129);
or U36903 (N_36903,N_22264,N_21566);
nor U36904 (N_36904,N_27350,N_29876);
nor U36905 (N_36905,N_23866,N_29584);
nand U36906 (N_36906,N_23714,N_25403);
xor U36907 (N_36907,N_29587,N_20542);
nor U36908 (N_36908,N_29673,N_20345);
nor U36909 (N_36909,N_25185,N_22012);
nand U36910 (N_36910,N_21155,N_20709);
nand U36911 (N_36911,N_28666,N_26517);
nor U36912 (N_36912,N_29986,N_21467);
nand U36913 (N_36913,N_29035,N_24084);
and U36914 (N_36914,N_24922,N_29080);
nand U36915 (N_36915,N_25854,N_29627);
and U36916 (N_36916,N_29015,N_27038);
and U36917 (N_36917,N_22078,N_23826);
xnor U36918 (N_36918,N_24198,N_26646);
nand U36919 (N_36919,N_27818,N_23337);
or U36920 (N_36920,N_28589,N_24397);
nor U36921 (N_36921,N_28420,N_22295);
nand U36922 (N_36922,N_23093,N_21105);
or U36923 (N_36923,N_26099,N_22875);
or U36924 (N_36924,N_21599,N_28720);
xor U36925 (N_36925,N_28279,N_20940);
xor U36926 (N_36926,N_24205,N_20373);
xor U36927 (N_36927,N_25804,N_24246);
nand U36928 (N_36928,N_28087,N_25747);
or U36929 (N_36929,N_25208,N_29238);
xor U36930 (N_36930,N_22420,N_21306);
and U36931 (N_36931,N_27279,N_26518);
nor U36932 (N_36932,N_23076,N_27907);
nor U36933 (N_36933,N_23266,N_26549);
nor U36934 (N_36934,N_27802,N_25747);
and U36935 (N_36935,N_27286,N_23047);
and U36936 (N_36936,N_27740,N_26491);
xor U36937 (N_36937,N_23309,N_20794);
xnor U36938 (N_36938,N_25324,N_21612);
or U36939 (N_36939,N_29182,N_25135);
xnor U36940 (N_36940,N_28285,N_26494);
nand U36941 (N_36941,N_23621,N_22067);
and U36942 (N_36942,N_23395,N_24906);
and U36943 (N_36943,N_20381,N_24002);
or U36944 (N_36944,N_21551,N_28625);
nor U36945 (N_36945,N_27936,N_22664);
nor U36946 (N_36946,N_22430,N_21503);
nand U36947 (N_36947,N_28803,N_26234);
xor U36948 (N_36948,N_28829,N_29395);
xnor U36949 (N_36949,N_25098,N_24855);
nor U36950 (N_36950,N_26847,N_27783);
nand U36951 (N_36951,N_25078,N_27805);
or U36952 (N_36952,N_23934,N_20254);
or U36953 (N_36953,N_21129,N_20179);
nand U36954 (N_36954,N_21744,N_21362);
nor U36955 (N_36955,N_24991,N_28728);
or U36956 (N_36956,N_24536,N_28531);
nor U36957 (N_36957,N_22110,N_23134);
nor U36958 (N_36958,N_21294,N_22252);
and U36959 (N_36959,N_20732,N_22737);
or U36960 (N_36960,N_24640,N_22928);
and U36961 (N_36961,N_27295,N_27832);
or U36962 (N_36962,N_23407,N_22857);
xnor U36963 (N_36963,N_21219,N_27115);
nand U36964 (N_36964,N_26845,N_24331);
nor U36965 (N_36965,N_24003,N_23197);
nor U36966 (N_36966,N_28222,N_27921);
and U36967 (N_36967,N_26553,N_20881);
xor U36968 (N_36968,N_24754,N_26276);
or U36969 (N_36969,N_28684,N_21389);
or U36970 (N_36970,N_26505,N_28210);
or U36971 (N_36971,N_27781,N_29788);
xnor U36972 (N_36972,N_28584,N_29116);
nor U36973 (N_36973,N_21879,N_26291);
xor U36974 (N_36974,N_20109,N_23994);
or U36975 (N_36975,N_28658,N_22614);
nand U36976 (N_36976,N_28787,N_23721);
nand U36977 (N_36977,N_26853,N_27016);
or U36978 (N_36978,N_26620,N_20317);
or U36979 (N_36979,N_29049,N_27691);
or U36980 (N_36980,N_27950,N_25323);
xor U36981 (N_36981,N_24139,N_28451);
nor U36982 (N_36982,N_26844,N_22110);
xor U36983 (N_36983,N_21602,N_26601);
nor U36984 (N_36984,N_27117,N_22961);
or U36985 (N_36985,N_22056,N_23678);
nand U36986 (N_36986,N_21559,N_25773);
xnor U36987 (N_36987,N_24665,N_24327);
nor U36988 (N_36988,N_21264,N_25436);
nand U36989 (N_36989,N_20537,N_21591);
or U36990 (N_36990,N_24848,N_25426);
or U36991 (N_36991,N_26294,N_26124);
xor U36992 (N_36992,N_23648,N_20606);
nor U36993 (N_36993,N_20936,N_26486);
and U36994 (N_36994,N_24908,N_27593);
nand U36995 (N_36995,N_22649,N_23085);
nand U36996 (N_36996,N_26391,N_29930);
nand U36997 (N_36997,N_25577,N_26862);
xor U36998 (N_36998,N_24699,N_25034);
or U36999 (N_36999,N_28550,N_22874);
or U37000 (N_37000,N_26481,N_20877);
xnor U37001 (N_37001,N_28812,N_25580);
nand U37002 (N_37002,N_21602,N_24614);
or U37003 (N_37003,N_20103,N_20574);
and U37004 (N_37004,N_20296,N_26728);
xor U37005 (N_37005,N_23911,N_29928);
nor U37006 (N_37006,N_20131,N_26354);
nor U37007 (N_37007,N_23423,N_22422);
xor U37008 (N_37008,N_24770,N_25001);
nor U37009 (N_37009,N_28585,N_28983);
xor U37010 (N_37010,N_28952,N_20842);
nand U37011 (N_37011,N_21931,N_29856);
and U37012 (N_37012,N_25594,N_29857);
or U37013 (N_37013,N_29979,N_27100);
and U37014 (N_37014,N_25126,N_21017);
xnor U37015 (N_37015,N_22369,N_20656);
xnor U37016 (N_37016,N_24075,N_27246);
or U37017 (N_37017,N_29427,N_24957);
and U37018 (N_37018,N_20698,N_24157);
nor U37019 (N_37019,N_21217,N_29124);
or U37020 (N_37020,N_29287,N_21604);
or U37021 (N_37021,N_27403,N_25401);
and U37022 (N_37022,N_26370,N_29221);
nor U37023 (N_37023,N_28187,N_20806);
nand U37024 (N_37024,N_26652,N_27540);
xor U37025 (N_37025,N_26305,N_25318);
xor U37026 (N_37026,N_23118,N_26040);
nand U37027 (N_37027,N_28925,N_23234);
nor U37028 (N_37028,N_21846,N_27330);
and U37029 (N_37029,N_22682,N_29394);
nor U37030 (N_37030,N_20253,N_27226);
or U37031 (N_37031,N_20207,N_22903);
nor U37032 (N_37032,N_26828,N_27656);
nand U37033 (N_37033,N_29423,N_20643);
xnor U37034 (N_37034,N_29542,N_23198);
and U37035 (N_37035,N_23449,N_23421);
or U37036 (N_37036,N_20117,N_23701);
or U37037 (N_37037,N_29463,N_27117);
xor U37038 (N_37038,N_25914,N_22392);
nand U37039 (N_37039,N_22876,N_22325);
nor U37040 (N_37040,N_29845,N_27616);
xor U37041 (N_37041,N_22504,N_27450);
nand U37042 (N_37042,N_28207,N_21805);
xnor U37043 (N_37043,N_23288,N_21415);
nand U37044 (N_37044,N_27028,N_21889);
and U37045 (N_37045,N_26948,N_29541);
or U37046 (N_37046,N_27694,N_25157);
and U37047 (N_37047,N_26606,N_22079);
or U37048 (N_37048,N_24485,N_28503);
and U37049 (N_37049,N_25071,N_25152);
or U37050 (N_37050,N_29476,N_23497);
nor U37051 (N_37051,N_26195,N_25408);
nor U37052 (N_37052,N_29609,N_24086);
xnor U37053 (N_37053,N_27945,N_29312);
nand U37054 (N_37054,N_24159,N_20317);
nand U37055 (N_37055,N_26666,N_24879);
xnor U37056 (N_37056,N_23659,N_22403);
and U37057 (N_37057,N_23203,N_20567);
or U37058 (N_37058,N_28470,N_27492);
nor U37059 (N_37059,N_27812,N_20002);
and U37060 (N_37060,N_24315,N_29901);
and U37061 (N_37061,N_28262,N_25219);
nand U37062 (N_37062,N_28421,N_29795);
xnor U37063 (N_37063,N_23819,N_29375);
nand U37064 (N_37064,N_22599,N_22499);
nor U37065 (N_37065,N_25403,N_26803);
xor U37066 (N_37066,N_26402,N_25093);
and U37067 (N_37067,N_20377,N_22902);
xnor U37068 (N_37068,N_22493,N_29371);
or U37069 (N_37069,N_29010,N_23001);
xor U37070 (N_37070,N_28506,N_24454);
xnor U37071 (N_37071,N_22571,N_27774);
xnor U37072 (N_37072,N_21838,N_24813);
xnor U37073 (N_37073,N_23711,N_24797);
and U37074 (N_37074,N_25412,N_28692);
nor U37075 (N_37075,N_24116,N_24624);
xor U37076 (N_37076,N_24008,N_26228);
xor U37077 (N_37077,N_22305,N_26866);
or U37078 (N_37078,N_27892,N_22884);
nand U37079 (N_37079,N_22940,N_24348);
xnor U37080 (N_37080,N_25524,N_25866);
xnor U37081 (N_37081,N_20295,N_23118);
nor U37082 (N_37082,N_26242,N_21008);
nor U37083 (N_37083,N_21916,N_27070);
nand U37084 (N_37084,N_25092,N_24936);
nand U37085 (N_37085,N_23748,N_21057);
xor U37086 (N_37086,N_29230,N_27672);
nor U37087 (N_37087,N_25338,N_23515);
or U37088 (N_37088,N_23704,N_24193);
and U37089 (N_37089,N_25010,N_27075);
nor U37090 (N_37090,N_23809,N_28750);
and U37091 (N_37091,N_21337,N_27798);
xor U37092 (N_37092,N_28279,N_29725);
and U37093 (N_37093,N_27157,N_24223);
xnor U37094 (N_37094,N_28340,N_25080);
nand U37095 (N_37095,N_28578,N_24255);
nand U37096 (N_37096,N_24034,N_27749);
xor U37097 (N_37097,N_22291,N_28844);
or U37098 (N_37098,N_28857,N_28808);
nand U37099 (N_37099,N_27744,N_26230);
xnor U37100 (N_37100,N_20416,N_28944);
or U37101 (N_37101,N_23915,N_29688);
nand U37102 (N_37102,N_28675,N_21697);
or U37103 (N_37103,N_22258,N_21137);
or U37104 (N_37104,N_25604,N_21884);
xor U37105 (N_37105,N_24205,N_25087);
xnor U37106 (N_37106,N_20708,N_21086);
or U37107 (N_37107,N_22286,N_23093);
and U37108 (N_37108,N_24663,N_27167);
nand U37109 (N_37109,N_26897,N_25831);
and U37110 (N_37110,N_26691,N_27990);
and U37111 (N_37111,N_27923,N_23846);
nand U37112 (N_37112,N_28438,N_20733);
nor U37113 (N_37113,N_24894,N_25458);
xnor U37114 (N_37114,N_24966,N_28546);
nand U37115 (N_37115,N_28231,N_28721);
xor U37116 (N_37116,N_23872,N_28961);
xnor U37117 (N_37117,N_24980,N_21484);
xnor U37118 (N_37118,N_26340,N_21126);
and U37119 (N_37119,N_28932,N_24570);
or U37120 (N_37120,N_28612,N_27307);
nor U37121 (N_37121,N_25545,N_27512);
nand U37122 (N_37122,N_24293,N_23847);
nand U37123 (N_37123,N_27768,N_20848);
xnor U37124 (N_37124,N_20040,N_20378);
and U37125 (N_37125,N_27108,N_23366);
nor U37126 (N_37126,N_25942,N_29433);
xnor U37127 (N_37127,N_24544,N_26843);
or U37128 (N_37128,N_26165,N_28889);
or U37129 (N_37129,N_23769,N_20437);
or U37130 (N_37130,N_25206,N_24714);
nor U37131 (N_37131,N_28267,N_29387);
and U37132 (N_37132,N_26297,N_21858);
nand U37133 (N_37133,N_29132,N_20562);
xor U37134 (N_37134,N_24410,N_25758);
nor U37135 (N_37135,N_25202,N_20573);
nor U37136 (N_37136,N_21348,N_26251);
and U37137 (N_37137,N_24666,N_20066);
and U37138 (N_37138,N_25466,N_29509);
or U37139 (N_37139,N_27010,N_22703);
and U37140 (N_37140,N_24994,N_29213);
nand U37141 (N_37141,N_24610,N_24573);
nor U37142 (N_37142,N_25274,N_25180);
nor U37143 (N_37143,N_20564,N_20098);
xor U37144 (N_37144,N_23078,N_26628);
xnor U37145 (N_37145,N_22038,N_21953);
xnor U37146 (N_37146,N_24043,N_21799);
nor U37147 (N_37147,N_28095,N_26873);
nand U37148 (N_37148,N_22007,N_29784);
nor U37149 (N_37149,N_29498,N_27694);
xnor U37150 (N_37150,N_26971,N_20504);
xnor U37151 (N_37151,N_29034,N_24352);
nand U37152 (N_37152,N_28473,N_26385);
nor U37153 (N_37153,N_23923,N_26807);
nand U37154 (N_37154,N_22048,N_27274);
or U37155 (N_37155,N_27986,N_21610);
nand U37156 (N_37156,N_29299,N_23977);
nand U37157 (N_37157,N_29063,N_20091);
or U37158 (N_37158,N_27034,N_23900);
nor U37159 (N_37159,N_21678,N_26295);
nand U37160 (N_37160,N_20137,N_23322);
or U37161 (N_37161,N_27271,N_27617);
and U37162 (N_37162,N_29249,N_28434);
or U37163 (N_37163,N_27133,N_22473);
nor U37164 (N_37164,N_24169,N_21097);
nor U37165 (N_37165,N_29559,N_25634);
nand U37166 (N_37166,N_22787,N_23879);
and U37167 (N_37167,N_27136,N_26060);
and U37168 (N_37168,N_25531,N_23459);
nor U37169 (N_37169,N_28880,N_28950);
nand U37170 (N_37170,N_25161,N_22422);
nor U37171 (N_37171,N_27243,N_23130);
and U37172 (N_37172,N_22742,N_23458);
or U37173 (N_37173,N_26566,N_27281);
nor U37174 (N_37174,N_21722,N_24750);
and U37175 (N_37175,N_25035,N_25498);
nand U37176 (N_37176,N_26895,N_24464);
or U37177 (N_37177,N_25518,N_26713);
nand U37178 (N_37178,N_21445,N_25109);
or U37179 (N_37179,N_24070,N_22718);
or U37180 (N_37180,N_22115,N_25981);
and U37181 (N_37181,N_26989,N_25375);
and U37182 (N_37182,N_25671,N_24498);
nand U37183 (N_37183,N_22832,N_20166);
nor U37184 (N_37184,N_27560,N_26106);
or U37185 (N_37185,N_21021,N_20904);
nor U37186 (N_37186,N_23680,N_21954);
nand U37187 (N_37187,N_27015,N_24278);
nor U37188 (N_37188,N_25948,N_28678);
and U37189 (N_37189,N_26065,N_21011);
nand U37190 (N_37190,N_24490,N_27100);
nor U37191 (N_37191,N_20989,N_29575);
xnor U37192 (N_37192,N_27294,N_20773);
xnor U37193 (N_37193,N_24356,N_24386);
nand U37194 (N_37194,N_22653,N_27995);
nor U37195 (N_37195,N_22060,N_22156);
nor U37196 (N_37196,N_21311,N_29721);
or U37197 (N_37197,N_28186,N_28563);
nor U37198 (N_37198,N_26248,N_25749);
and U37199 (N_37199,N_28516,N_20029);
nand U37200 (N_37200,N_25134,N_25007);
nor U37201 (N_37201,N_27804,N_21647);
nor U37202 (N_37202,N_28339,N_21941);
xnor U37203 (N_37203,N_29972,N_23551);
nor U37204 (N_37204,N_29096,N_21867);
nor U37205 (N_37205,N_29930,N_20927);
nand U37206 (N_37206,N_26268,N_21739);
xnor U37207 (N_37207,N_27739,N_25248);
and U37208 (N_37208,N_27296,N_29689);
xnor U37209 (N_37209,N_20941,N_27795);
nand U37210 (N_37210,N_27667,N_28932);
or U37211 (N_37211,N_29359,N_21802);
nand U37212 (N_37212,N_20376,N_27015);
xnor U37213 (N_37213,N_25414,N_25348);
and U37214 (N_37214,N_27144,N_25146);
xnor U37215 (N_37215,N_26077,N_21928);
or U37216 (N_37216,N_29676,N_21033);
and U37217 (N_37217,N_23808,N_22981);
or U37218 (N_37218,N_22615,N_28312);
nand U37219 (N_37219,N_21539,N_26597);
or U37220 (N_37220,N_26058,N_25948);
nor U37221 (N_37221,N_25723,N_28267);
nand U37222 (N_37222,N_26709,N_20983);
or U37223 (N_37223,N_27868,N_20462);
xor U37224 (N_37224,N_27607,N_24287);
and U37225 (N_37225,N_22612,N_26423);
and U37226 (N_37226,N_26991,N_26680);
and U37227 (N_37227,N_22160,N_20124);
or U37228 (N_37228,N_28459,N_25244);
nand U37229 (N_37229,N_29319,N_24475);
nand U37230 (N_37230,N_21990,N_22907);
and U37231 (N_37231,N_27068,N_28140);
and U37232 (N_37232,N_20397,N_20070);
and U37233 (N_37233,N_25070,N_26150);
xor U37234 (N_37234,N_29691,N_28756);
nand U37235 (N_37235,N_26454,N_25713);
nand U37236 (N_37236,N_25568,N_20972);
and U37237 (N_37237,N_20159,N_22712);
nor U37238 (N_37238,N_24337,N_26218);
and U37239 (N_37239,N_27251,N_22428);
or U37240 (N_37240,N_20633,N_29057);
xnor U37241 (N_37241,N_29973,N_25066);
nor U37242 (N_37242,N_27046,N_23088);
nor U37243 (N_37243,N_25306,N_20651);
nand U37244 (N_37244,N_29593,N_26740);
xnor U37245 (N_37245,N_22735,N_25422);
nand U37246 (N_37246,N_22495,N_25825);
nand U37247 (N_37247,N_28163,N_24887);
nand U37248 (N_37248,N_28181,N_24211);
or U37249 (N_37249,N_28197,N_20836);
and U37250 (N_37250,N_27786,N_20630);
or U37251 (N_37251,N_23787,N_28853);
or U37252 (N_37252,N_26929,N_25213);
xor U37253 (N_37253,N_23760,N_28175);
or U37254 (N_37254,N_25016,N_24807);
or U37255 (N_37255,N_26205,N_24249);
or U37256 (N_37256,N_27429,N_29639);
and U37257 (N_37257,N_21992,N_29859);
xor U37258 (N_37258,N_21472,N_27562);
nand U37259 (N_37259,N_24848,N_26700);
nor U37260 (N_37260,N_24257,N_21920);
xnor U37261 (N_37261,N_21699,N_22039);
and U37262 (N_37262,N_27890,N_27012);
xor U37263 (N_37263,N_27247,N_24070);
and U37264 (N_37264,N_26921,N_24809);
and U37265 (N_37265,N_21262,N_21659);
nand U37266 (N_37266,N_26790,N_25654);
xnor U37267 (N_37267,N_23798,N_20837);
xor U37268 (N_37268,N_26411,N_25233);
or U37269 (N_37269,N_21687,N_28374);
or U37270 (N_37270,N_29606,N_22010);
nor U37271 (N_37271,N_23308,N_23805);
nand U37272 (N_37272,N_27805,N_20149);
and U37273 (N_37273,N_20909,N_23972);
and U37274 (N_37274,N_22052,N_24646);
or U37275 (N_37275,N_22951,N_23350);
xnor U37276 (N_37276,N_26153,N_29872);
xor U37277 (N_37277,N_24270,N_22038);
nand U37278 (N_37278,N_27003,N_25265);
or U37279 (N_37279,N_21240,N_20240);
or U37280 (N_37280,N_26397,N_22873);
and U37281 (N_37281,N_20197,N_23231);
nor U37282 (N_37282,N_29605,N_23741);
xnor U37283 (N_37283,N_28561,N_24129);
nand U37284 (N_37284,N_23927,N_26295);
xor U37285 (N_37285,N_23497,N_26252);
or U37286 (N_37286,N_27662,N_29043);
and U37287 (N_37287,N_27976,N_25261);
and U37288 (N_37288,N_23507,N_22345);
or U37289 (N_37289,N_27820,N_24689);
and U37290 (N_37290,N_25030,N_25536);
and U37291 (N_37291,N_29538,N_26947);
xor U37292 (N_37292,N_23291,N_22645);
nor U37293 (N_37293,N_24366,N_24923);
nor U37294 (N_37294,N_20484,N_24481);
or U37295 (N_37295,N_26749,N_27751);
nand U37296 (N_37296,N_26839,N_21596);
and U37297 (N_37297,N_23070,N_25451);
xor U37298 (N_37298,N_21585,N_24754);
nand U37299 (N_37299,N_23467,N_20242);
xnor U37300 (N_37300,N_20909,N_25616);
nand U37301 (N_37301,N_22178,N_20330);
or U37302 (N_37302,N_28959,N_22962);
nand U37303 (N_37303,N_22776,N_28398);
and U37304 (N_37304,N_24969,N_21096);
xor U37305 (N_37305,N_27053,N_27151);
xnor U37306 (N_37306,N_27666,N_29428);
or U37307 (N_37307,N_23455,N_21237);
and U37308 (N_37308,N_28058,N_26047);
nor U37309 (N_37309,N_27214,N_28267);
and U37310 (N_37310,N_25354,N_23430);
nor U37311 (N_37311,N_20251,N_21061);
and U37312 (N_37312,N_25044,N_24343);
or U37313 (N_37313,N_26663,N_29999);
or U37314 (N_37314,N_21713,N_23941);
and U37315 (N_37315,N_24685,N_21267);
xor U37316 (N_37316,N_27760,N_21571);
nand U37317 (N_37317,N_21891,N_20398);
xnor U37318 (N_37318,N_20705,N_22061);
or U37319 (N_37319,N_26047,N_23780);
nor U37320 (N_37320,N_27446,N_23661);
nor U37321 (N_37321,N_25370,N_24576);
or U37322 (N_37322,N_24347,N_21425);
and U37323 (N_37323,N_21477,N_22072);
nand U37324 (N_37324,N_25532,N_29657);
or U37325 (N_37325,N_28376,N_20543);
xor U37326 (N_37326,N_27717,N_23397);
nor U37327 (N_37327,N_28856,N_20519);
and U37328 (N_37328,N_27983,N_29175);
nand U37329 (N_37329,N_20389,N_29602);
and U37330 (N_37330,N_26720,N_28483);
nor U37331 (N_37331,N_28008,N_26639);
nor U37332 (N_37332,N_22188,N_27452);
nor U37333 (N_37333,N_22315,N_20868);
nand U37334 (N_37334,N_25535,N_25521);
xnor U37335 (N_37335,N_29065,N_25127);
and U37336 (N_37336,N_22383,N_27845);
and U37337 (N_37337,N_26155,N_20095);
and U37338 (N_37338,N_22989,N_20391);
or U37339 (N_37339,N_26859,N_24650);
xnor U37340 (N_37340,N_29464,N_26922);
nor U37341 (N_37341,N_27363,N_27066);
nor U37342 (N_37342,N_29185,N_27840);
or U37343 (N_37343,N_20318,N_26440);
nand U37344 (N_37344,N_26967,N_26844);
and U37345 (N_37345,N_27754,N_21791);
nor U37346 (N_37346,N_26115,N_29729);
and U37347 (N_37347,N_26890,N_20409);
xor U37348 (N_37348,N_27609,N_23809);
xor U37349 (N_37349,N_27772,N_24830);
nor U37350 (N_37350,N_27425,N_20873);
xor U37351 (N_37351,N_23537,N_29566);
nand U37352 (N_37352,N_24336,N_23664);
nor U37353 (N_37353,N_27145,N_20588);
nand U37354 (N_37354,N_28224,N_26481);
nand U37355 (N_37355,N_26141,N_22812);
nor U37356 (N_37356,N_21994,N_28370);
xnor U37357 (N_37357,N_21860,N_26536);
nand U37358 (N_37358,N_23975,N_25676);
nor U37359 (N_37359,N_23518,N_22712);
nand U37360 (N_37360,N_25320,N_20813);
or U37361 (N_37361,N_28069,N_28926);
nor U37362 (N_37362,N_20511,N_28270);
nor U37363 (N_37363,N_29998,N_24387);
nor U37364 (N_37364,N_26425,N_27611);
nor U37365 (N_37365,N_23811,N_22655);
xnor U37366 (N_37366,N_29466,N_22882);
and U37367 (N_37367,N_24214,N_21477);
nand U37368 (N_37368,N_24917,N_29493);
and U37369 (N_37369,N_24397,N_20473);
or U37370 (N_37370,N_21400,N_28481);
nor U37371 (N_37371,N_28476,N_25914);
nand U37372 (N_37372,N_28225,N_22153);
xnor U37373 (N_37373,N_25907,N_26086);
nand U37374 (N_37374,N_26302,N_25908);
nor U37375 (N_37375,N_29489,N_24643);
nor U37376 (N_37376,N_24902,N_27867);
or U37377 (N_37377,N_26808,N_27880);
nor U37378 (N_37378,N_20326,N_24172);
nor U37379 (N_37379,N_25551,N_22142);
xnor U37380 (N_37380,N_20900,N_29439);
nor U37381 (N_37381,N_22986,N_21800);
and U37382 (N_37382,N_21010,N_21000);
and U37383 (N_37383,N_25603,N_21128);
or U37384 (N_37384,N_26383,N_25406);
or U37385 (N_37385,N_26177,N_24687);
xnor U37386 (N_37386,N_27690,N_25957);
nand U37387 (N_37387,N_21424,N_29667);
or U37388 (N_37388,N_26223,N_20613);
or U37389 (N_37389,N_20460,N_29956);
or U37390 (N_37390,N_21528,N_21899);
nor U37391 (N_37391,N_28067,N_25645);
or U37392 (N_37392,N_20166,N_27153);
xnor U37393 (N_37393,N_29238,N_26117);
and U37394 (N_37394,N_24327,N_23368);
xnor U37395 (N_37395,N_27387,N_28767);
and U37396 (N_37396,N_24227,N_29967);
or U37397 (N_37397,N_29965,N_24230);
nor U37398 (N_37398,N_26716,N_21857);
nand U37399 (N_37399,N_26118,N_22002);
nor U37400 (N_37400,N_27014,N_20766);
nor U37401 (N_37401,N_28991,N_23295);
nand U37402 (N_37402,N_28607,N_26167);
and U37403 (N_37403,N_22624,N_26953);
and U37404 (N_37404,N_27878,N_26361);
xor U37405 (N_37405,N_20664,N_27726);
nor U37406 (N_37406,N_29171,N_27471);
xnor U37407 (N_37407,N_21107,N_22241);
and U37408 (N_37408,N_24336,N_26159);
nand U37409 (N_37409,N_24932,N_25518);
and U37410 (N_37410,N_26787,N_27736);
or U37411 (N_37411,N_23129,N_24291);
xnor U37412 (N_37412,N_29844,N_27013);
xnor U37413 (N_37413,N_25571,N_29695);
nand U37414 (N_37414,N_26304,N_22262);
or U37415 (N_37415,N_25933,N_27472);
xnor U37416 (N_37416,N_20538,N_29276);
nand U37417 (N_37417,N_25759,N_26086);
nand U37418 (N_37418,N_24770,N_23504);
or U37419 (N_37419,N_27994,N_28826);
and U37420 (N_37420,N_24784,N_22810);
or U37421 (N_37421,N_24786,N_21418);
and U37422 (N_37422,N_27546,N_29633);
or U37423 (N_37423,N_28396,N_27783);
nand U37424 (N_37424,N_26075,N_27837);
and U37425 (N_37425,N_24957,N_24161);
nand U37426 (N_37426,N_20210,N_26029);
and U37427 (N_37427,N_22094,N_29592);
or U37428 (N_37428,N_25272,N_22851);
or U37429 (N_37429,N_21585,N_25948);
nor U37430 (N_37430,N_21674,N_21946);
or U37431 (N_37431,N_22561,N_23169);
or U37432 (N_37432,N_23674,N_23939);
or U37433 (N_37433,N_27835,N_26261);
or U37434 (N_37434,N_20573,N_28601);
and U37435 (N_37435,N_27395,N_24457);
nand U37436 (N_37436,N_20898,N_25866);
nand U37437 (N_37437,N_22465,N_27238);
or U37438 (N_37438,N_29974,N_23610);
nor U37439 (N_37439,N_27898,N_25935);
nor U37440 (N_37440,N_26048,N_21900);
nand U37441 (N_37441,N_21390,N_20427);
xor U37442 (N_37442,N_24789,N_29949);
and U37443 (N_37443,N_22008,N_26848);
xor U37444 (N_37444,N_23199,N_25379);
nor U37445 (N_37445,N_22692,N_23332);
or U37446 (N_37446,N_28879,N_21017);
or U37447 (N_37447,N_26799,N_20977);
nor U37448 (N_37448,N_26632,N_25504);
nand U37449 (N_37449,N_28592,N_23792);
nor U37450 (N_37450,N_28497,N_20857);
nor U37451 (N_37451,N_22147,N_27707);
nor U37452 (N_37452,N_28151,N_26851);
xnor U37453 (N_37453,N_27162,N_21256);
xor U37454 (N_37454,N_29873,N_25272);
or U37455 (N_37455,N_29624,N_22132);
nand U37456 (N_37456,N_28668,N_24070);
xnor U37457 (N_37457,N_20620,N_27957);
nor U37458 (N_37458,N_28028,N_20084);
or U37459 (N_37459,N_28097,N_29316);
xnor U37460 (N_37460,N_28520,N_25052);
or U37461 (N_37461,N_26432,N_29946);
nand U37462 (N_37462,N_29852,N_20517);
or U37463 (N_37463,N_28272,N_26648);
nor U37464 (N_37464,N_28804,N_24751);
or U37465 (N_37465,N_26907,N_28297);
nor U37466 (N_37466,N_22497,N_28489);
nor U37467 (N_37467,N_27923,N_22320);
nand U37468 (N_37468,N_23659,N_22722);
nand U37469 (N_37469,N_27004,N_28487);
nand U37470 (N_37470,N_25233,N_25752);
nor U37471 (N_37471,N_21378,N_20270);
or U37472 (N_37472,N_27881,N_23275);
xor U37473 (N_37473,N_22620,N_22107);
and U37474 (N_37474,N_28698,N_29693);
and U37475 (N_37475,N_24446,N_25022);
or U37476 (N_37476,N_26813,N_22743);
and U37477 (N_37477,N_22580,N_27204);
xnor U37478 (N_37478,N_21058,N_21678);
and U37479 (N_37479,N_29558,N_22394);
and U37480 (N_37480,N_25823,N_29934);
xnor U37481 (N_37481,N_29177,N_21778);
and U37482 (N_37482,N_26064,N_26939);
or U37483 (N_37483,N_22861,N_20386);
nand U37484 (N_37484,N_26260,N_20462);
nand U37485 (N_37485,N_20461,N_20668);
xor U37486 (N_37486,N_20747,N_22074);
xor U37487 (N_37487,N_24655,N_23450);
and U37488 (N_37488,N_25992,N_22289);
and U37489 (N_37489,N_25671,N_21830);
xor U37490 (N_37490,N_23884,N_22342);
or U37491 (N_37491,N_26417,N_22122);
nand U37492 (N_37492,N_20710,N_24362);
xor U37493 (N_37493,N_23008,N_23893);
and U37494 (N_37494,N_29737,N_22505);
or U37495 (N_37495,N_26828,N_29606);
or U37496 (N_37496,N_25216,N_20570);
xnor U37497 (N_37497,N_26927,N_26092);
nor U37498 (N_37498,N_22331,N_25655);
nor U37499 (N_37499,N_25555,N_24172);
nor U37500 (N_37500,N_24733,N_26005);
xnor U37501 (N_37501,N_29137,N_27692);
nor U37502 (N_37502,N_21283,N_27161);
xnor U37503 (N_37503,N_21141,N_21395);
and U37504 (N_37504,N_23010,N_20351);
and U37505 (N_37505,N_26916,N_24444);
and U37506 (N_37506,N_22340,N_26011);
nor U37507 (N_37507,N_21152,N_26053);
nor U37508 (N_37508,N_23660,N_26117);
or U37509 (N_37509,N_25536,N_29469);
nand U37510 (N_37510,N_22920,N_29979);
and U37511 (N_37511,N_21656,N_22494);
xnor U37512 (N_37512,N_22978,N_29766);
or U37513 (N_37513,N_28173,N_22311);
nor U37514 (N_37514,N_27874,N_25319);
nand U37515 (N_37515,N_23642,N_24660);
xor U37516 (N_37516,N_29149,N_26648);
nor U37517 (N_37517,N_29964,N_28840);
and U37518 (N_37518,N_29182,N_21328);
xor U37519 (N_37519,N_27735,N_22469);
xor U37520 (N_37520,N_26440,N_29620);
and U37521 (N_37521,N_24930,N_23459);
and U37522 (N_37522,N_24189,N_20713);
or U37523 (N_37523,N_28843,N_29259);
nand U37524 (N_37524,N_20813,N_28009);
or U37525 (N_37525,N_23388,N_24783);
or U37526 (N_37526,N_26862,N_24386);
xnor U37527 (N_37527,N_20145,N_27684);
xnor U37528 (N_37528,N_25017,N_25390);
and U37529 (N_37529,N_25586,N_24588);
and U37530 (N_37530,N_20309,N_23611);
and U37531 (N_37531,N_28187,N_27856);
nor U37532 (N_37532,N_23670,N_24703);
nor U37533 (N_37533,N_21021,N_24245);
and U37534 (N_37534,N_21587,N_29108);
nor U37535 (N_37535,N_22211,N_22396);
nand U37536 (N_37536,N_20061,N_29112);
xor U37537 (N_37537,N_25376,N_27400);
xor U37538 (N_37538,N_22411,N_23916);
nor U37539 (N_37539,N_24448,N_20202);
or U37540 (N_37540,N_22958,N_23157);
nor U37541 (N_37541,N_20908,N_23340);
and U37542 (N_37542,N_23592,N_20746);
nand U37543 (N_37543,N_26560,N_29368);
nor U37544 (N_37544,N_24889,N_21327);
xor U37545 (N_37545,N_25006,N_27110);
nor U37546 (N_37546,N_24130,N_29611);
or U37547 (N_37547,N_26135,N_20253);
nor U37548 (N_37548,N_21000,N_28582);
nand U37549 (N_37549,N_20833,N_25162);
or U37550 (N_37550,N_21554,N_24529);
and U37551 (N_37551,N_29281,N_20979);
nor U37552 (N_37552,N_28597,N_21010);
nor U37553 (N_37553,N_25912,N_21517);
nor U37554 (N_37554,N_20487,N_20061);
nand U37555 (N_37555,N_21292,N_26498);
or U37556 (N_37556,N_29210,N_24694);
nand U37557 (N_37557,N_25512,N_20671);
nand U37558 (N_37558,N_21466,N_20064);
and U37559 (N_37559,N_28037,N_21607);
and U37560 (N_37560,N_22399,N_21681);
xnor U37561 (N_37561,N_23793,N_21626);
nand U37562 (N_37562,N_28235,N_24554);
xnor U37563 (N_37563,N_27632,N_20147);
or U37564 (N_37564,N_22776,N_25316);
xor U37565 (N_37565,N_20506,N_28739);
or U37566 (N_37566,N_29701,N_25700);
or U37567 (N_37567,N_20110,N_29139);
or U37568 (N_37568,N_26804,N_20106);
nand U37569 (N_37569,N_23175,N_29015);
nand U37570 (N_37570,N_28495,N_26570);
xnor U37571 (N_37571,N_29961,N_21805);
xnor U37572 (N_37572,N_29617,N_27434);
xnor U37573 (N_37573,N_29911,N_20834);
or U37574 (N_37574,N_26373,N_28295);
and U37575 (N_37575,N_25094,N_28759);
or U37576 (N_37576,N_23806,N_28580);
or U37577 (N_37577,N_22960,N_23507);
and U37578 (N_37578,N_25937,N_27754);
or U37579 (N_37579,N_26039,N_24195);
nor U37580 (N_37580,N_24300,N_23498);
and U37581 (N_37581,N_23270,N_29704);
nand U37582 (N_37582,N_24999,N_23491);
and U37583 (N_37583,N_22768,N_20363);
xnor U37584 (N_37584,N_25268,N_25904);
xor U37585 (N_37585,N_23093,N_27047);
xor U37586 (N_37586,N_22968,N_28076);
xor U37587 (N_37587,N_25809,N_28884);
nand U37588 (N_37588,N_22662,N_23123);
and U37589 (N_37589,N_28862,N_24772);
and U37590 (N_37590,N_27892,N_29921);
nor U37591 (N_37591,N_26764,N_23899);
xnor U37592 (N_37592,N_24591,N_24736);
and U37593 (N_37593,N_28401,N_26988);
nor U37594 (N_37594,N_29851,N_29913);
or U37595 (N_37595,N_21874,N_21176);
nand U37596 (N_37596,N_25581,N_22421);
or U37597 (N_37597,N_23291,N_26760);
nor U37598 (N_37598,N_25953,N_22606);
nand U37599 (N_37599,N_27513,N_21353);
nand U37600 (N_37600,N_25230,N_26273);
or U37601 (N_37601,N_28328,N_24322);
or U37602 (N_37602,N_28765,N_20512);
xnor U37603 (N_37603,N_21278,N_22630);
or U37604 (N_37604,N_28781,N_21705);
nor U37605 (N_37605,N_26063,N_27460);
nor U37606 (N_37606,N_23926,N_27248);
nand U37607 (N_37607,N_20255,N_28119);
nor U37608 (N_37608,N_26035,N_24691);
nand U37609 (N_37609,N_23064,N_29584);
nand U37610 (N_37610,N_25896,N_23703);
or U37611 (N_37611,N_20617,N_29899);
nor U37612 (N_37612,N_26771,N_20373);
xnor U37613 (N_37613,N_26537,N_21281);
or U37614 (N_37614,N_20783,N_29609);
nor U37615 (N_37615,N_27092,N_23423);
or U37616 (N_37616,N_26573,N_29840);
nor U37617 (N_37617,N_20710,N_24425);
and U37618 (N_37618,N_24548,N_26434);
and U37619 (N_37619,N_28718,N_29426);
or U37620 (N_37620,N_26148,N_26229);
xor U37621 (N_37621,N_27042,N_20738);
and U37622 (N_37622,N_25974,N_29286);
and U37623 (N_37623,N_25635,N_22777);
nand U37624 (N_37624,N_23372,N_24169);
nor U37625 (N_37625,N_26449,N_29625);
and U37626 (N_37626,N_22135,N_28292);
nor U37627 (N_37627,N_24119,N_29955);
nand U37628 (N_37628,N_20530,N_27818);
nor U37629 (N_37629,N_22335,N_25492);
nand U37630 (N_37630,N_22353,N_21432);
xnor U37631 (N_37631,N_26152,N_25115);
or U37632 (N_37632,N_27037,N_23415);
nand U37633 (N_37633,N_26716,N_20944);
xnor U37634 (N_37634,N_21376,N_20813);
and U37635 (N_37635,N_29479,N_22828);
xor U37636 (N_37636,N_27006,N_22018);
nor U37637 (N_37637,N_26158,N_22837);
and U37638 (N_37638,N_22814,N_24441);
and U37639 (N_37639,N_28729,N_20026);
and U37640 (N_37640,N_26537,N_21115);
or U37641 (N_37641,N_25467,N_25618);
nand U37642 (N_37642,N_29941,N_25301);
xor U37643 (N_37643,N_25084,N_24662);
and U37644 (N_37644,N_24928,N_27860);
and U37645 (N_37645,N_26511,N_28710);
xnor U37646 (N_37646,N_23274,N_25839);
nand U37647 (N_37647,N_29951,N_21539);
nand U37648 (N_37648,N_25581,N_25256);
or U37649 (N_37649,N_29075,N_24860);
and U37650 (N_37650,N_21318,N_22469);
or U37651 (N_37651,N_23702,N_20096);
nand U37652 (N_37652,N_20213,N_26672);
nor U37653 (N_37653,N_22226,N_28540);
nor U37654 (N_37654,N_26759,N_24881);
nor U37655 (N_37655,N_28540,N_25451);
and U37656 (N_37656,N_21250,N_24966);
nand U37657 (N_37657,N_29204,N_29403);
nand U37658 (N_37658,N_21436,N_26512);
or U37659 (N_37659,N_23730,N_24330);
xor U37660 (N_37660,N_25148,N_26166);
and U37661 (N_37661,N_20971,N_25449);
nor U37662 (N_37662,N_29816,N_26303);
or U37663 (N_37663,N_25310,N_27527);
nor U37664 (N_37664,N_28076,N_28487);
xnor U37665 (N_37665,N_20256,N_28277);
nor U37666 (N_37666,N_24483,N_26258);
or U37667 (N_37667,N_25888,N_27102);
or U37668 (N_37668,N_27719,N_29197);
xor U37669 (N_37669,N_21364,N_22273);
nor U37670 (N_37670,N_24814,N_23212);
or U37671 (N_37671,N_24456,N_22155);
and U37672 (N_37672,N_23554,N_25996);
nor U37673 (N_37673,N_29316,N_22439);
nand U37674 (N_37674,N_28997,N_29299);
or U37675 (N_37675,N_25491,N_22967);
nand U37676 (N_37676,N_20543,N_24554);
nand U37677 (N_37677,N_24109,N_26824);
or U37678 (N_37678,N_21915,N_28581);
nor U37679 (N_37679,N_29709,N_24825);
or U37680 (N_37680,N_23066,N_27386);
nor U37681 (N_37681,N_23414,N_23132);
nor U37682 (N_37682,N_26390,N_25903);
xor U37683 (N_37683,N_22785,N_22038);
nor U37684 (N_37684,N_26056,N_26918);
xor U37685 (N_37685,N_25476,N_20080);
nor U37686 (N_37686,N_23214,N_22354);
xnor U37687 (N_37687,N_22435,N_27762);
nor U37688 (N_37688,N_29878,N_28658);
or U37689 (N_37689,N_29398,N_27470);
nand U37690 (N_37690,N_26174,N_20406);
or U37691 (N_37691,N_26406,N_20052);
xnor U37692 (N_37692,N_21626,N_25089);
and U37693 (N_37693,N_26000,N_23960);
or U37694 (N_37694,N_21331,N_26003);
nor U37695 (N_37695,N_20957,N_29476);
nor U37696 (N_37696,N_22841,N_28789);
nand U37697 (N_37697,N_29832,N_22687);
nor U37698 (N_37698,N_20510,N_23180);
nand U37699 (N_37699,N_27217,N_27875);
and U37700 (N_37700,N_25558,N_21650);
or U37701 (N_37701,N_22327,N_25313);
nor U37702 (N_37702,N_25297,N_20330);
or U37703 (N_37703,N_27322,N_21822);
and U37704 (N_37704,N_22384,N_24187);
or U37705 (N_37705,N_23698,N_20943);
nor U37706 (N_37706,N_25751,N_20980);
and U37707 (N_37707,N_25097,N_29897);
nor U37708 (N_37708,N_29178,N_24022);
and U37709 (N_37709,N_27083,N_29827);
xnor U37710 (N_37710,N_22543,N_24072);
or U37711 (N_37711,N_24258,N_24448);
nand U37712 (N_37712,N_26792,N_23622);
or U37713 (N_37713,N_24094,N_22789);
or U37714 (N_37714,N_23333,N_22084);
or U37715 (N_37715,N_26101,N_23700);
nor U37716 (N_37716,N_28716,N_21941);
nor U37717 (N_37717,N_20754,N_28639);
nand U37718 (N_37718,N_24867,N_29469);
nor U37719 (N_37719,N_28000,N_26188);
nor U37720 (N_37720,N_26716,N_24068);
or U37721 (N_37721,N_22880,N_23213);
nand U37722 (N_37722,N_21457,N_21402);
xor U37723 (N_37723,N_25885,N_27091);
and U37724 (N_37724,N_29619,N_29803);
nor U37725 (N_37725,N_26400,N_23392);
nor U37726 (N_37726,N_22739,N_21040);
nor U37727 (N_37727,N_25479,N_24417);
nand U37728 (N_37728,N_22326,N_23494);
xor U37729 (N_37729,N_28835,N_21352);
nor U37730 (N_37730,N_24511,N_28099);
xor U37731 (N_37731,N_29216,N_27899);
xnor U37732 (N_37732,N_25463,N_28564);
and U37733 (N_37733,N_20768,N_26802);
nand U37734 (N_37734,N_28779,N_20124);
nand U37735 (N_37735,N_29394,N_27148);
nand U37736 (N_37736,N_21289,N_20421);
xnor U37737 (N_37737,N_29848,N_22246);
nor U37738 (N_37738,N_27424,N_22627);
nor U37739 (N_37739,N_26473,N_26570);
nand U37740 (N_37740,N_20797,N_20834);
and U37741 (N_37741,N_27803,N_20628);
nand U37742 (N_37742,N_23616,N_23515);
xnor U37743 (N_37743,N_25265,N_25387);
nor U37744 (N_37744,N_25459,N_23900);
nand U37745 (N_37745,N_26891,N_26509);
and U37746 (N_37746,N_20574,N_25893);
xnor U37747 (N_37747,N_28916,N_27719);
or U37748 (N_37748,N_24220,N_21493);
nand U37749 (N_37749,N_24724,N_28756);
nor U37750 (N_37750,N_29788,N_22877);
xor U37751 (N_37751,N_21012,N_20282);
xnor U37752 (N_37752,N_23951,N_21806);
and U37753 (N_37753,N_22559,N_27312);
or U37754 (N_37754,N_29995,N_23373);
or U37755 (N_37755,N_24727,N_20493);
xor U37756 (N_37756,N_21414,N_20341);
and U37757 (N_37757,N_23363,N_20531);
and U37758 (N_37758,N_29430,N_24433);
nor U37759 (N_37759,N_29503,N_23075);
nand U37760 (N_37760,N_23311,N_25878);
and U37761 (N_37761,N_20638,N_22877);
nand U37762 (N_37762,N_20899,N_20046);
and U37763 (N_37763,N_27624,N_21723);
xnor U37764 (N_37764,N_28547,N_29054);
and U37765 (N_37765,N_21491,N_26499);
and U37766 (N_37766,N_24289,N_25157);
nor U37767 (N_37767,N_29391,N_22058);
or U37768 (N_37768,N_26592,N_26208);
or U37769 (N_37769,N_25538,N_27706);
and U37770 (N_37770,N_28686,N_21057);
xor U37771 (N_37771,N_27696,N_27840);
nand U37772 (N_37772,N_29062,N_26537);
nor U37773 (N_37773,N_25648,N_28176);
nor U37774 (N_37774,N_20933,N_29116);
or U37775 (N_37775,N_27327,N_26764);
and U37776 (N_37776,N_27819,N_26787);
xor U37777 (N_37777,N_21689,N_29931);
and U37778 (N_37778,N_21617,N_25797);
nor U37779 (N_37779,N_20317,N_26286);
xnor U37780 (N_37780,N_29747,N_20162);
nor U37781 (N_37781,N_26254,N_28308);
xor U37782 (N_37782,N_23460,N_21655);
or U37783 (N_37783,N_29009,N_24348);
and U37784 (N_37784,N_28520,N_23687);
nor U37785 (N_37785,N_23162,N_25472);
xor U37786 (N_37786,N_29735,N_21493);
or U37787 (N_37787,N_29695,N_22298);
nor U37788 (N_37788,N_20268,N_21289);
nor U37789 (N_37789,N_20465,N_28383);
and U37790 (N_37790,N_23012,N_29794);
nand U37791 (N_37791,N_29269,N_24901);
nor U37792 (N_37792,N_28433,N_24955);
and U37793 (N_37793,N_28921,N_27007);
xor U37794 (N_37794,N_25829,N_26421);
and U37795 (N_37795,N_26749,N_24455);
and U37796 (N_37796,N_20704,N_29994);
xnor U37797 (N_37797,N_29683,N_29051);
nand U37798 (N_37798,N_26618,N_21242);
xor U37799 (N_37799,N_29763,N_24237);
and U37800 (N_37800,N_22191,N_20874);
or U37801 (N_37801,N_29173,N_29364);
nand U37802 (N_37802,N_29523,N_27062);
xnor U37803 (N_37803,N_26324,N_23130);
xor U37804 (N_37804,N_24071,N_24218);
or U37805 (N_37805,N_28273,N_25689);
and U37806 (N_37806,N_27564,N_27670);
nor U37807 (N_37807,N_21705,N_26789);
and U37808 (N_37808,N_22186,N_28153);
or U37809 (N_37809,N_28609,N_26785);
or U37810 (N_37810,N_22593,N_24697);
nand U37811 (N_37811,N_23850,N_29496);
nand U37812 (N_37812,N_25259,N_29614);
xor U37813 (N_37813,N_22899,N_24473);
and U37814 (N_37814,N_27390,N_21106);
nand U37815 (N_37815,N_20846,N_27542);
and U37816 (N_37816,N_27870,N_23535);
xor U37817 (N_37817,N_22913,N_22560);
and U37818 (N_37818,N_28213,N_21297);
and U37819 (N_37819,N_22422,N_22097);
and U37820 (N_37820,N_26707,N_27728);
nor U37821 (N_37821,N_22474,N_21698);
or U37822 (N_37822,N_20550,N_20842);
nand U37823 (N_37823,N_26090,N_25366);
and U37824 (N_37824,N_25004,N_20371);
nand U37825 (N_37825,N_28057,N_21774);
nand U37826 (N_37826,N_22498,N_29048);
and U37827 (N_37827,N_26522,N_26630);
nor U37828 (N_37828,N_29930,N_23816);
nor U37829 (N_37829,N_28039,N_21713);
nor U37830 (N_37830,N_27978,N_25214);
or U37831 (N_37831,N_28617,N_23569);
and U37832 (N_37832,N_29259,N_24693);
xnor U37833 (N_37833,N_26582,N_27387);
nor U37834 (N_37834,N_26355,N_20105);
and U37835 (N_37835,N_28426,N_29439);
nand U37836 (N_37836,N_25327,N_25315);
nor U37837 (N_37837,N_29438,N_21222);
nand U37838 (N_37838,N_28497,N_29961);
nand U37839 (N_37839,N_21503,N_22956);
and U37840 (N_37840,N_24196,N_22451);
nand U37841 (N_37841,N_27661,N_25341);
and U37842 (N_37842,N_23456,N_27449);
and U37843 (N_37843,N_20836,N_27966);
nand U37844 (N_37844,N_23352,N_27669);
nor U37845 (N_37845,N_24893,N_25541);
and U37846 (N_37846,N_28951,N_25214);
nor U37847 (N_37847,N_22613,N_27287);
nand U37848 (N_37848,N_22166,N_21423);
nor U37849 (N_37849,N_28501,N_22010);
nand U37850 (N_37850,N_25064,N_25847);
and U37851 (N_37851,N_24865,N_29833);
and U37852 (N_37852,N_28868,N_22204);
nand U37853 (N_37853,N_26271,N_21558);
nor U37854 (N_37854,N_23305,N_26914);
or U37855 (N_37855,N_25410,N_26842);
or U37856 (N_37856,N_24034,N_25618);
or U37857 (N_37857,N_28730,N_22972);
and U37858 (N_37858,N_29386,N_28709);
nor U37859 (N_37859,N_27356,N_24004);
and U37860 (N_37860,N_29286,N_28558);
xnor U37861 (N_37861,N_28422,N_24862);
nand U37862 (N_37862,N_20816,N_23537);
nand U37863 (N_37863,N_25278,N_28220);
nor U37864 (N_37864,N_29269,N_22930);
nand U37865 (N_37865,N_22725,N_29354);
nand U37866 (N_37866,N_29437,N_20756);
or U37867 (N_37867,N_20420,N_24064);
xnor U37868 (N_37868,N_23533,N_29372);
nor U37869 (N_37869,N_20571,N_23751);
and U37870 (N_37870,N_25388,N_24150);
nand U37871 (N_37871,N_23168,N_23120);
nand U37872 (N_37872,N_27504,N_21990);
nor U37873 (N_37873,N_22762,N_24483);
nand U37874 (N_37874,N_26112,N_24341);
and U37875 (N_37875,N_28914,N_24431);
nor U37876 (N_37876,N_27601,N_20445);
xor U37877 (N_37877,N_22878,N_26640);
xor U37878 (N_37878,N_27169,N_23945);
and U37879 (N_37879,N_21337,N_23629);
nor U37880 (N_37880,N_25083,N_28622);
xnor U37881 (N_37881,N_24974,N_28637);
nand U37882 (N_37882,N_21426,N_26745);
xor U37883 (N_37883,N_29106,N_25635);
nor U37884 (N_37884,N_24763,N_24012);
xor U37885 (N_37885,N_20599,N_29154);
or U37886 (N_37886,N_27970,N_23076);
or U37887 (N_37887,N_20995,N_21060);
nand U37888 (N_37888,N_26121,N_25507);
or U37889 (N_37889,N_29971,N_23346);
and U37890 (N_37890,N_25102,N_29836);
nand U37891 (N_37891,N_22161,N_27420);
nor U37892 (N_37892,N_21397,N_22675);
or U37893 (N_37893,N_27738,N_27932);
nand U37894 (N_37894,N_28188,N_26413);
or U37895 (N_37895,N_21258,N_28994);
xor U37896 (N_37896,N_22331,N_28499);
xor U37897 (N_37897,N_21582,N_25270);
nand U37898 (N_37898,N_29184,N_25248);
nand U37899 (N_37899,N_27433,N_24434);
xor U37900 (N_37900,N_22475,N_20581);
or U37901 (N_37901,N_29961,N_24905);
nand U37902 (N_37902,N_28963,N_22739);
nand U37903 (N_37903,N_20980,N_25136);
nor U37904 (N_37904,N_23419,N_21246);
and U37905 (N_37905,N_22617,N_26501);
or U37906 (N_37906,N_24850,N_25488);
nor U37907 (N_37907,N_20069,N_24982);
nor U37908 (N_37908,N_26627,N_20134);
xor U37909 (N_37909,N_22252,N_29163);
nor U37910 (N_37910,N_26760,N_29294);
nand U37911 (N_37911,N_24104,N_29590);
and U37912 (N_37912,N_27130,N_27656);
or U37913 (N_37913,N_23042,N_26714);
or U37914 (N_37914,N_27121,N_24283);
or U37915 (N_37915,N_29081,N_27339);
xor U37916 (N_37916,N_25939,N_23252);
and U37917 (N_37917,N_25857,N_27832);
nor U37918 (N_37918,N_20567,N_27018);
and U37919 (N_37919,N_23336,N_28552);
nor U37920 (N_37920,N_23244,N_28997);
and U37921 (N_37921,N_21353,N_22087);
xnor U37922 (N_37922,N_24913,N_24967);
xor U37923 (N_37923,N_23619,N_26689);
xnor U37924 (N_37924,N_28068,N_27816);
nor U37925 (N_37925,N_24109,N_29381);
or U37926 (N_37926,N_28929,N_20745);
xnor U37927 (N_37927,N_20011,N_20533);
or U37928 (N_37928,N_21755,N_24566);
nand U37929 (N_37929,N_29473,N_22744);
or U37930 (N_37930,N_27210,N_22144);
or U37931 (N_37931,N_20343,N_28050);
and U37932 (N_37932,N_20622,N_20540);
and U37933 (N_37933,N_28768,N_24134);
or U37934 (N_37934,N_21790,N_25481);
nor U37935 (N_37935,N_26407,N_27706);
nand U37936 (N_37936,N_23138,N_26082);
or U37937 (N_37937,N_28418,N_28730);
or U37938 (N_37938,N_22443,N_26323);
nor U37939 (N_37939,N_26814,N_27564);
or U37940 (N_37940,N_24497,N_28360);
xnor U37941 (N_37941,N_29100,N_24018);
xnor U37942 (N_37942,N_21203,N_23945);
and U37943 (N_37943,N_23297,N_27019);
nor U37944 (N_37944,N_23977,N_29421);
and U37945 (N_37945,N_21677,N_28981);
or U37946 (N_37946,N_22272,N_22255);
xnor U37947 (N_37947,N_23386,N_21874);
and U37948 (N_37948,N_24857,N_20397);
nor U37949 (N_37949,N_26224,N_20624);
or U37950 (N_37950,N_25761,N_20596);
nor U37951 (N_37951,N_27812,N_25127);
and U37952 (N_37952,N_26887,N_28993);
nand U37953 (N_37953,N_22741,N_25816);
or U37954 (N_37954,N_28388,N_25559);
nand U37955 (N_37955,N_25042,N_23402);
or U37956 (N_37956,N_21141,N_28678);
xnor U37957 (N_37957,N_29618,N_24092);
nor U37958 (N_37958,N_25586,N_28132);
xor U37959 (N_37959,N_24384,N_27018);
and U37960 (N_37960,N_26670,N_22861);
and U37961 (N_37961,N_27526,N_25360);
nand U37962 (N_37962,N_25922,N_26493);
and U37963 (N_37963,N_23241,N_29281);
xnor U37964 (N_37964,N_23113,N_24886);
nand U37965 (N_37965,N_26018,N_24732);
xor U37966 (N_37966,N_24770,N_29153);
xnor U37967 (N_37967,N_21480,N_20085);
xnor U37968 (N_37968,N_23026,N_21857);
nor U37969 (N_37969,N_26925,N_22717);
nand U37970 (N_37970,N_27819,N_25453);
nand U37971 (N_37971,N_29689,N_27662);
nor U37972 (N_37972,N_20664,N_25481);
and U37973 (N_37973,N_21963,N_27999);
and U37974 (N_37974,N_24717,N_20198);
nand U37975 (N_37975,N_27784,N_24357);
xnor U37976 (N_37976,N_29263,N_28724);
nor U37977 (N_37977,N_26581,N_25659);
xnor U37978 (N_37978,N_20526,N_25197);
and U37979 (N_37979,N_25920,N_26346);
xor U37980 (N_37980,N_21559,N_25549);
xnor U37981 (N_37981,N_24571,N_24707);
or U37982 (N_37982,N_27314,N_27366);
or U37983 (N_37983,N_27034,N_29837);
nor U37984 (N_37984,N_26066,N_28428);
nand U37985 (N_37985,N_25354,N_22160);
and U37986 (N_37986,N_20732,N_20397);
xor U37987 (N_37987,N_26682,N_28961);
nor U37988 (N_37988,N_22783,N_25429);
and U37989 (N_37989,N_28654,N_28268);
nand U37990 (N_37990,N_28677,N_22764);
nand U37991 (N_37991,N_20507,N_29615);
and U37992 (N_37992,N_21391,N_24531);
nor U37993 (N_37993,N_20306,N_27806);
nor U37994 (N_37994,N_23989,N_28277);
xnor U37995 (N_37995,N_25534,N_20075);
nand U37996 (N_37996,N_22704,N_27158);
nand U37997 (N_37997,N_21515,N_24684);
and U37998 (N_37998,N_26270,N_20100);
nand U37999 (N_37999,N_29620,N_25885);
nor U38000 (N_38000,N_21080,N_23746);
nor U38001 (N_38001,N_24813,N_27081);
or U38002 (N_38002,N_26853,N_26948);
or U38003 (N_38003,N_28423,N_23855);
xor U38004 (N_38004,N_20110,N_24618);
xnor U38005 (N_38005,N_29026,N_24327);
or U38006 (N_38006,N_24927,N_27084);
xnor U38007 (N_38007,N_24564,N_27175);
or U38008 (N_38008,N_25065,N_26441);
and U38009 (N_38009,N_24507,N_26631);
nand U38010 (N_38010,N_24655,N_26013);
nand U38011 (N_38011,N_25990,N_25498);
or U38012 (N_38012,N_28254,N_20656);
xor U38013 (N_38013,N_28538,N_24244);
nand U38014 (N_38014,N_29894,N_25940);
or U38015 (N_38015,N_27944,N_22002);
nand U38016 (N_38016,N_23511,N_23835);
or U38017 (N_38017,N_27014,N_27938);
and U38018 (N_38018,N_22965,N_28986);
xnor U38019 (N_38019,N_23385,N_25758);
nand U38020 (N_38020,N_20419,N_22669);
nor U38021 (N_38021,N_22314,N_25886);
nand U38022 (N_38022,N_28141,N_23947);
nor U38023 (N_38023,N_25209,N_25892);
xor U38024 (N_38024,N_24513,N_24572);
nor U38025 (N_38025,N_21408,N_26195);
and U38026 (N_38026,N_28664,N_23167);
nor U38027 (N_38027,N_24397,N_22943);
xor U38028 (N_38028,N_25569,N_20163);
and U38029 (N_38029,N_26410,N_27077);
and U38030 (N_38030,N_23352,N_29923);
or U38031 (N_38031,N_29520,N_27922);
nand U38032 (N_38032,N_22049,N_24769);
xor U38033 (N_38033,N_22430,N_27447);
and U38034 (N_38034,N_27870,N_22361);
and U38035 (N_38035,N_29861,N_28980);
xor U38036 (N_38036,N_22195,N_24968);
xor U38037 (N_38037,N_28657,N_21863);
xnor U38038 (N_38038,N_22086,N_21944);
xor U38039 (N_38039,N_22571,N_24886);
nand U38040 (N_38040,N_22192,N_22074);
nor U38041 (N_38041,N_23975,N_23427);
nor U38042 (N_38042,N_24934,N_23216);
nor U38043 (N_38043,N_24244,N_26034);
and U38044 (N_38044,N_23297,N_24535);
or U38045 (N_38045,N_24038,N_25899);
xor U38046 (N_38046,N_25054,N_20073);
and U38047 (N_38047,N_28525,N_28885);
nand U38048 (N_38048,N_27509,N_23652);
nand U38049 (N_38049,N_22324,N_22662);
nor U38050 (N_38050,N_24773,N_21202);
xor U38051 (N_38051,N_28629,N_25886);
or U38052 (N_38052,N_24729,N_20316);
nor U38053 (N_38053,N_29779,N_25960);
and U38054 (N_38054,N_21953,N_21150);
or U38055 (N_38055,N_20809,N_27671);
and U38056 (N_38056,N_23122,N_21022);
nand U38057 (N_38057,N_25231,N_21104);
and U38058 (N_38058,N_22315,N_23408);
nand U38059 (N_38059,N_23676,N_21340);
and U38060 (N_38060,N_20668,N_26367);
nor U38061 (N_38061,N_20038,N_29055);
xnor U38062 (N_38062,N_29699,N_23150);
or U38063 (N_38063,N_28455,N_23499);
and U38064 (N_38064,N_21702,N_28899);
and U38065 (N_38065,N_26157,N_29838);
xnor U38066 (N_38066,N_23547,N_23610);
and U38067 (N_38067,N_25624,N_26452);
nand U38068 (N_38068,N_24178,N_26783);
and U38069 (N_38069,N_23812,N_25135);
nand U38070 (N_38070,N_27948,N_29469);
or U38071 (N_38071,N_22389,N_29516);
or U38072 (N_38072,N_21112,N_26684);
nor U38073 (N_38073,N_24328,N_23664);
xor U38074 (N_38074,N_20628,N_20835);
nand U38075 (N_38075,N_28769,N_22261);
and U38076 (N_38076,N_21279,N_28616);
nand U38077 (N_38077,N_21852,N_25377);
xor U38078 (N_38078,N_20763,N_29845);
nand U38079 (N_38079,N_20207,N_29128);
nand U38080 (N_38080,N_24284,N_29454);
and U38081 (N_38081,N_21110,N_24984);
or U38082 (N_38082,N_22319,N_28098);
xnor U38083 (N_38083,N_21846,N_28078);
or U38084 (N_38084,N_21513,N_26079);
or U38085 (N_38085,N_23967,N_20345);
nand U38086 (N_38086,N_29288,N_21139);
xor U38087 (N_38087,N_27578,N_28561);
and U38088 (N_38088,N_27298,N_29326);
nand U38089 (N_38089,N_29161,N_27498);
nand U38090 (N_38090,N_21737,N_27937);
and U38091 (N_38091,N_22846,N_25198);
xor U38092 (N_38092,N_28031,N_24125);
nor U38093 (N_38093,N_28338,N_23022);
nand U38094 (N_38094,N_24772,N_27524);
or U38095 (N_38095,N_22821,N_20697);
or U38096 (N_38096,N_26944,N_25823);
nand U38097 (N_38097,N_26505,N_29006);
or U38098 (N_38098,N_29887,N_29448);
nor U38099 (N_38099,N_28908,N_25659);
and U38100 (N_38100,N_24038,N_23066);
nor U38101 (N_38101,N_22949,N_23415);
xnor U38102 (N_38102,N_23511,N_26825);
or U38103 (N_38103,N_29707,N_28731);
xnor U38104 (N_38104,N_22019,N_28926);
nand U38105 (N_38105,N_24471,N_20219);
nor U38106 (N_38106,N_26161,N_29048);
xnor U38107 (N_38107,N_23145,N_23040);
nand U38108 (N_38108,N_24418,N_29003);
xor U38109 (N_38109,N_26511,N_24915);
nand U38110 (N_38110,N_20222,N_22301);
or U38111 (N_38111,N_29874,N_23634);
nor U38112 (N_38112,N_25328,N_22044);
xnor U38113 (N_38113,N_23806,N_26858);
or U38114 (N_38114,N_27184,N_24094);
nand U38115 (N_38115,N_27357,N_24830);
or U38116 (N_38116,N_20566,N_26068);
xor U38117 (N_38117,N_24636,N_26587);
xor U38118 (N_38118,N_27089,N_23684);
nor U38119 (N_38119,N_21233,N_28331);
or U38120 (N_38120,N_25455,N_20799);
nor U38121 (N_38121,N_23540,N_24788);
and U38122 (N_38122,N_23133,N_23051);
nor U38123 (N_38123,N_28297,N_26228);
nand U38124 (N_38124,N_22058,N_29518);
nand U38125 (N_38125,N_22269,N_28634);
nand U38126 (N_38126,N_25589,N_25016);
nand U38127 (N_38127,N_27902,N_21326);
or U38128 (N_38128,N_27027,N_26612);
xor U38129 (N_38129,N_23548,N_20096);
and U38130 (N_38130,N_20774,N_21314);
and U38131 (N_38131,N_21222,N_20933);
nand U38132 (N_38132,N_29897,N_26637);
nor U38133 (N_38133,N_21282,N_21596);
nand U38134 (N_38134,N_27917,N_29682);
xnor U38135 (N_38135,N_28022,N_23864);
and U38136 (N_38136,N_22459,N_25287);
or U38137 (N_38137,N_25045,N_25455);
nor U38138 (N_38138,N_25006,N_29815);
nand U38139 (N_38139,N_21857,N_25913);
and U38140 (N_38140,N_28771,N_24868);
and U38141 (N_38141,N_24432,N_26974);
or U38142 (N_38142,N_22163,N_22132);
xnor U38143 (N_38143,N_26152,N_29194);
and U38144 (N_38144,N_22488,N_29924);
nand U38145 (N_38145,N_24667,N_27036);
xor U38146 (N_38146,N_26547,N_26250);
nor U38147 (N_38147,N_21669,N_26819);
nor U38148 (N_38148,N_21643,N_21258);
nand U38149 (N_38149,N_22638,N_20255);
nor U38150 (N_38150,N_22551,N_27599);
or U38151 (N_38151,N_20137,N_29311);
and U38152 (N_38152,N_28816,N_23618);
nand U38153 (N_38153,N_20158,N_23545);
or U38154 (N_38154,N_24512,N_28796);
nor U38155 (N_38155,N_23017,N_25884);
or U38156 (N_38156,N_22157,N_29994);
xnor U38157 (N_38157,N_23480,N_21870);
nand U38158 (N_38158,N_21400,N_20461);
and U38159 (N_38159,N_22034,N_22724);
and U38160 (N_38160,N_26178,N_23566);
or U38161 (N_38161,N_23514,N_24711);
or U38162 (N_38162,N_23696,N_25786);
or U38163 (N_38163,N_26555,N_20606);
nand U38164 (N_38164,N_21145,N_23056);
nand U38165 (N_38165,N_24527,N_22322);
and U38166 (N_38166,N_20475,N_26904);
nor U38167 (N_38167,N_23769,N_25513);
xor U38168 (N_38168,N_23694,N_27999);
nor U38169 (N_38169,N_27521,N_22771);
and U38170 (N_38170,N_21748,N_22246);
nand U38171 (N_38171,N_28340,N_21711);
nand U38172 (N_38172,N_23630,N_29410);
nor U38173 (N_38173,N_22024,N_25282);
nand U38174 (N_38174,N_20192,N_26178);
nand U38175 (N_38175,N_21706,N_28160);
and U38176 (N_38176,N_26717,N_25929);
nor U38177 (N_38177,N_26867,N_24008);
nor U38178 (N_38178,N_24382,N_25495);
nand U38179 (N_38179,N_21912,N_23693);
nor U38180 (N_38180,N_28582,N_21137);
and U38181 (N_38181,N_26506,N_24690);
or U38182 (N_38182,N_29570,N_21483);
nor U38183 (N_38183,N_21516,N_24930);
xor U38184 (N_38184,N_25243,N_23172);
xnor U38185 (N_38185,N_21747,N_24920);
xnor U38186 (N_38186,N_24231,N_27453);
nand U38187 (N_38187,N_27555,N_29530);
xnor U38188 (N_38188,N_21973,N_21237);
xor U38189 (N_38189,N_24039,N_26513);
nand U38190 (N_38190,N_21157,N_28064);
nor U38191 (N_38191,N_29041,N_27332);
xnor U38192 (N_38192,N_21424,N_21832);
or U38193 (N_38193,N_20661,N_26355);
or U38194 (N_38194,N_22392,N_29151);
nor U38195 (N_38195,N_21977,N_25138);
and U38196 (N_38196,N_26074,N_29055);
nor U38197 (N_38197,N_28811,N_21192);
xnor U38198 (N_38198,N_27965,N_25180);
or U38199 (N_38199,N_26387,N_26027);
nand U38200 (N_38200,N_27231,N_25348);
nor U38201 (N_38201,N_23421,N_23775);
and U38202 (N_38202,N_24817,N_27899);
nor U38203 (N_38203,N_26709,N_29303);
nand U38204 (N_38204,N_23577,N_23300);
nand U38205 (N_38205,N_22384,N_25370);
nand U38206 (N_38206,N_26798,N_29469);
nor U38207 (N_38207,N_25386,N_20905);
or U38208 (N_38208,N_24995,N_20563);
and U38209 (N_38209,N_27481,N_24447);
nor U38210 (N_38210,N_24766,N_27713);
nand U38211 (N_38211,N_26119,N_21732);
and U38212 (N_38212,N_23289,N_28778);
xor U38213 (N_38213,N_27693,N_29781);
nand U38214 (N_38214,N_23980,N_28366);
and U38215 (N_38215,N_26042,N_26142);
nor U38216 (N_38216,N_22695,N_26733);
and U38217 (N_38217,N_24880,N_29789);
xor U38218 (N_38218,N_28242,N_27026);
or U38219 (N_38219,N_22332,N_22834);
nand U38220 (N_38220,N_20246,N_27451);
and U38221 (N_38221,N_29042,N_21915);
and U38222 (N_38222,N_26166,N_24074);
or U38223 (N_38223,N_27393,N_22526);
nor U38224 (N_38224,N_25140,N_22291);
nand U38225 (N_38225,N_24954,N_28267);
nand U38226 (N_38226,N_26978,N_28656);
or U38227 (N_38227,N_24495,N_22254);
nand U38228 (N_38228,N_23938,N_23557);
and U38229 (N_38229,N_24913,N_27699);
xor U38230 (N_38230,N_26883,N_26080);
nor U38231 (N_38231,N_21366,N_21956);
nand U38232 (N_38232,N_22092,N_20519);
nand U38233 (N_38233,N_25911,N_27545);
nor U38234 (N_38234,N_21915,N_29879);
and U38235 (N_38235,N_25499,N_27343);
nand U38236 (N_38236,N_21724,N_23231);
nand U38237 (N_38237,N_29863,N_28961);
and U38238 (N_38238,N_26727,N_28011);
or U38239 (N_38239,N_25169,N_20459);
nand U38240 (N_38240,N_20769,N_23752);
xnor U38241 (N_38241,N_20228,N_25028);
nand U38242 (N_38242,N_24464,N_29193);
or U38243 (N_38243,N_26502,N_29529);
nor U38244 (N_38244,N_28079,N_23820);
nand U38245 (N_38245,N_24258,N_23621);
nor U38246 (N_38246,N_22975,N_25520);
xor U38247 (N_38247,N_23970,N_23463);
nand U38248 (N_38248,N_22760,N_22911);
and U38249 (N_38249,N_20196,N_21177);
and U38250 (N_38250,N_24902,N_29214);
xor U38251 (N_38251,N_24614,N_28171);
nor U38252 (N_38252,N_26366,N_28282);
xnor U38253 (N_38253,N_21085,N_27765);
nand U38254 (N_38254,N_22008,N_22562);
and U38255 (N_38255,N_24811,N_27122);
or U38256 (N_38256,N_27981,N_29647);
xnor U38257 (N_38257,N_27503,N_20542);
or U38258 (N_38258,N_27218,N_24442);
nand U38259 (N_38259,N_24283,N_25852);
xnor U38260 (N_38260,N_27308,N_22061);
or U38261 (N_38261,N_26102,N_27793);
and U38262 (N_38262,N_22861,N_29566);
or U38263 (N_38263,N_22224,N_23906);
nor U38264 (N_38264,N_24102,N_26465);
and U38265 (N_38265,N_25121,N_26603);
or U38266 (N_38266,N_22128,N_25428);
and U38267 (N_38267,N_27320,N_21658);
or U38268 (N_38268,N_25729,N_23506);
or U38269 (N_38269,N_27267,N_26434);
nand U38270 (N_38270,N_27091,N_28671);
and U38271 (N_38271,N_21891,N_23469);
and U38272 (N_38272,N_24672,N_23487);
and U38273 (N_38273,N_24977,N_27368);
xor U38274 (N_38274,N_24409,N_20815);
and U38275 (N_38275,N_24079,N_20019);
or U38276 (N_38276,N_27723,N_27000);
or U38277 (N_38277,N_23844,N_26852);
nor U38278 (N_38278,N_23358,N_24175);
xor U38279 (N_38279,N_24433,N_29618);
or U38280 (N_38280,N_25769,N_23036);
nor U38281 (N_38281,N_25026,N_20466);
and U38282 (N_38282,N_26292,N_27477);
xnor U38283 (N_38283,N_26562,N_29472);
or U38284 (N_38284,N_20368,N_22675);
or U38285 (N_38285,N_26756,N_20917);
nand U38286 (N_38286,N_29901,N_26341);
nor U38287 (N_38287,N_29764,N_20953);
and U38288 (N_38288,N_27025,N_24348);
xnor U38289 (N_38289,N_26834,N_29537);
and U38290 (N_38290,N_22997,N_24718);
xor U38291 (N_38291,N_22735,N_27312);
xnor U38292 (N_38292,N_28501,N_28155);
nor U38293 (N_38293,N_27425,N_25962);
nor U38294 (N_38294,N_20367,N_28718);
and U38295 (N_38295,N_25620,N_26767);
xor U38296 (N_38296,N_22959,N_24500);
and U38297 (N_38297,N_21070,N_23280);
or U38298 (N_38298,N_25628,N_27800);
or U38299 (N_38299,N_23407,N_23965);
or U38300 (N_38300,N_29045,N_28794);
xor U38301 (N_38301,N_28604,N_26015);
xnor U38302 (N_38302,N_22467,N_28041);
and U38303 (N_38303,N_29163,N_24999);
or U38304 (N_38304,N_20711,N_28841);
nor U38305 (N_38305,N_24570,N_28995);
nand U38306 (N_38306,N_26759,N_23706);
xor U38307 (N_38307,N_21740,N_20814);
xor U38308 (N_38308,N_25728,N_29573);
nand U38309 (N_38309,N_23778,N_28533);
and U38310 (N_38310,N_22631,N_24658);
or U38311 (N_38311,N_26391,N_20881);
and U38312 (N_38312,N_27164,N_24592);
nor U38313 (N_38313,N_23699,N_21320);
and U38314 (N_38314,N_27869,N_23687);
and U38315 (N_38315,N_25793,N_24048);
nor U38316 (N_38316,N_29303,N_24095);
nor U38317 (N_38317,N_25118,N_21501);
xnor U38318 (N_38318,N_22052,N_27751);
or U38319 (N_38319,N_24036,N_24791);
nor U38320 (N_38320,N_26893,N_28059);
xor U38321 (N_38321,N_28847,N_21970);
and U38322 (N_38322,N_26306,N_22001);
xor U38323 (N_38323,N_24136,N_28929);
nand U38324 (N_38324,N_24565,N_23934);
or U38325 (N_38325,N_26976,N_22225);
nor U38326 (N_38326,N_23182,N_27664);
nand U38327 (N_38327,N_21141,N_26392);
nand U38328 (N_38328,N_21264,N_25983);
nor U38329 (N_38329,N_27142,N_20844);
and U38330 (N_38330,N_25502,N_20655);
xor U38331 (N_38331,N_28490,N_21199);
xor U38332 (N_38332,N_25938,N_22694);
xor U38333 (N_38333,N_29027,N_25661);
xor U38334 (N_38334,N_20473,N_28934);
nor U38335 (N_38335,N_22382,N_21491);
nor U38336 (N_38336,N_24713,N_21639);
nor U38337 (N_38337,N_20241,N_20410);
and U38338 (N_38338,N_24952,N_28540);
and U38339 (N_38339,N_21869,N_22435);
or U38340 (N_38340,N_20074,N_24010);
or U38341 (N_38341,N_28894,N_23601);
or U38342 (N_38342,N_24027,N_23257);
or U38343 (N_38343,N_23142,N_24178);
and U38344 (N_38344,N_21849,N_21286);
nor U38345 (N_38345,N_29851,N_20217);
xnor U38346 (N_38346,N_29252,N_27076);
and U38347 (N_38347,N_23767,N_20051);
and U38348 (N_38348,N_25951,N_25886);
nor U38349 (N_38349,N_22855,N_21840);
and U38350 (N_38350,N_27937,N_26115);
nand U38351 (N_38351,N_28609,N_24481);
nand U38352 (N_38352,N_23158,N_24054);
nand U38353 (N_38353,N_20056,N_26712);
xnor U38354 (N_38354,N_28051,N_24479);
or U38355 (N_38355,N_24932,N_29217);
nor U38356 (N_38356,N_24501,N_29911);
and U38357 (N_38357,N_26263,N_29720);
nor U38358 (N_38358,N_22488,N_25962);
nor U38359 (N_38359,N_29321,N_26409);
nand U38360 (N_38360,N_26722,N_24573);
and U38361 (N_38361,N_22675,N_28667);
xor U38362 (N_38362,N_26861,N_24672);
nand U38363 (N_38363,N_27241,N_27891);
nand U38364 (N_38364,N_29558,N_29797);
xnor U38365 (N_38365,N_23044,N_25321);
and U38366 (N_38366,N_21479,N_21011);
or U38367 (N_38367,N_28244,N_20985);
and U38368 (N_38368,N_22126,N_29441);
and U38369 (N_38369,N_26350,N_20178);
xnor U38370 (N_38370,N_20602,N_26169);
or U38371 (N_38371,N_20010,N_26914);
nor U38372 (N_38372,N_20069,N_24446);
nand U38373 (N_38373,N_28601,N_27782);
or U38374 (N_38374,N_29335,N_26589);
nand U38375 (N_38375,N_29345,N_26130);
and U38376 (N_38376,N_22482,N_24105);
and U38377 (N_38377,N_26105,N_21770);
or U38378 (N_38378,N_27386,N_27280);
or U38379 (N_38379,N_26018,N_29275);
nand U38380 (N_38380,N_25459,N_24157);
nor U38381 (N_38381,N_23297,N_23379);
xnor U38382 (N_38382,N_23413,N_26233);
and U38383 (N_38383,N_28031,N_21999);
nand U38384 (N_38384,N_23249,N_22176);
xor U38385 (N_38385,N_26373,N_29199);
nor U38386 (N_38386,N_25744,N_21388);
and U38387 (N_38387,N_23655,N_28486);
nor U38388 (N_38388,N_25540,N_24895);
xor U38389 (N_38389,N_26355,N_23491);
or U38390 (N_38390,N_24049,N_22356);
or U38391 (N_38391,N_24591,N_29885);
nand U38392 (N_38392,N_23451,N_26184);
or U38393 (N_38393,N_25636,N_26945);
nor U38394 (N_38394,N_28917,N_27174);
nor U38395 (N_38395,N_20275,N_25226);
nand U38396 (N_38396,N_22157,N_26928);
nand U38397 (N_38397,N_23895,N_24299);
and U38398 (N_38398,N_28817,N_20316);
xnor U38399 (N_38399,N_20973,N_27074);
xor U38400 (N_38400,N_28135,N_25667);
or U38401 (N_38401,N_21122,N_20603);
nand U38402 (N_38402,N_21111,N_26954);
nor U38403 (N_38403,N_28489,N_24314);
xor U38404 (N_38404,N_21223,N_22992);
nor U38405 (N_38405,N_23581,N_23524);
xnor U38406 (N_38406,N_29414,N_21859);
and U38407 (N_38407,N_21221,N_26027);
xor U38408 (N_38408,N_21737,N_22880);
or U38409 (N_38409,N_21597,N_23179);
nor U38410 (N_38410,N_23766,N_28456);
xor U38411 (N_38411,N_26764,N_29788);
xor U38412 (N_38412,N_22476,N_28845);
nand U38413 (N_38413,N_22608,N_23407);
or U38414 (N_38414,N_24321,N_21594);
nand U38415 (N_38415,N_27205,N_28490);
nand U38416 (N_38416,N_21162,N_27634);
nor U38417 (N_38417,N_20777,N_27334);
nand U38418 (N_38418,N_20811,N_23874);
or U38419 (N_38419,N_29450,N_20383);
nor U38420 (N_38420,N_22244,N_26165);
xnor U38421 (N_38421,N_27494,N_20400);
and U38422 (N_38422,N_25961,N_22927);
or U38423 (N_38423,N_25743,N_27841);
nand U38424 (N_38424,N_23498,N_24208);
or U38425 (N_38425,N_20031,N_27762);
nand U38426 (N_38426,N_27642,N_20046);
nor U38427 (N_38427,N_20654,N_29010);
nor U38428 (N_38428,N_25484,N_26679);
and U38429 (N_38429,N_20058,N_26101);
or U38430 (N_38430,N_29377,N_25316);
or U38431 (N_38431,N_22123,N_24719);
nor U38432 (N_38432,N_25315,N_21532);
nor U38433 (N_38433,N_28450,N_27068);
and U38434 (N_38434,N_29798,N_26254);
nor U38435 (N_38435,N_23388,N_20719);
nand U38436 (N_38436,N_21305,N_23834);
and U38437 (N_38437,N_24612,N_20876);
and U38438 (N_38438,N_29707,N_26608);
xor U38439 (N_38439,N_29388,N_27313);
nand U38440 (N_38440,N_29798,N_28719);
xor U38441 (N_38441,N_24053,N_28600);
and U38442 (N_38442,N_24488,N_21477);
and U38443 (N_38443,N_29086,N_25179);
and U38444 (N_38444,N_24961,N_29859);
nor U38445 (N_38445,N_21748,N_28787);
nand U38446 (N_38446,N_29011,N_24844);
nand U38447 (N_38447,N_21821,N_29063);
nor U38448 (N_38448,N_27699,N_26294);
xor U38449 (N_38449,N_21547,N_21793);
and U38450 (N_38450,N_24780,N_28532);
nor U38451 (N_38451,N_27427,N_23508);
nor U38452 (N_38452,N_22294,N_27113);
or U38453 (N_38453,N_25852,N_23009);
or U38454 (N_38454,N_24656,N_22065);
xor U38455 (N_38455,N_26648,N_25251);
nor U38456 (N_38456,N_29529,N_22220);
or U38457 (N_38457,N_23023,N_21440);
nand U38458 (N_38458,N_29617,N_29671);
nor U38459 (N_38459,N_22195,N_26972);
and U38460 (N_38460,N_26646,N_20991);
or U38461 (N_38461,N_25881,N_23159);
nand U38462 (N_38462,N_23633,N_24695);
nor U38463 (N_38463,N_24195,N_22679);
nand U38464 (N_38464,N_29995,N_22388);
and U38465 (N_38465,N_29656,N_29614);
nand U38466 (N_38466,N_27065,N_27156);
xnor U38467 (N_38467,N_24488,N_28906);
or U38468 (N_38468,N_26593,N_29311);
xor U38469 (N_38469,N_25038,N_21876);
nor U38470 (N_38470,N_28990,N_23394);
nor U38471 (N_38471,N_22143,N_28263);
or U38472 (N_38472,N_21452,N_21193);
and U38473 (N_38473,N_23996,N_20783);
and U38474 (N_38474,N_27291,N_25545);
and U38475 (N_38475,N_27383,N_23376);
and U38476 (N_38476,N_29386,N_23684);
xor U38477 (N_38477,N_22869,N_25571);
xnor U38478 (N_38478,N_20775,N_20349);
nor U38479 (N_38479,N_20283,N_24532);
nor U38480 (N_38480,N_21094,N_22168);
xnor U38481 (N_38481,N_27053,N_22695);
nor U38482 (N_38482,N_27224,N_21897);
nor U38483 (N_38483,N_20674,N_23110);
and U38484 (N_38484,N_23906,N_26783);
or U38485 (N_38485,N_28964,N_24020);
nand U38486 (N_38486,N_20677,N_24130);
xor U38487 (N_38487,N_22399,N_28143);
and U38488 (N_38488,N_26256,N_20987);
nand U38489 (N_38489,N_29785,N_27951);
or U38490 (N_38490,N_25545,N_20434);
nand U38491 (N_38491,N_29102,N_22836);
xnor U38492 (N_38492,N_28530,N_29180);
nand U38493 (N_38493,N_26296,N_22468);
and U38494 (N_38494,N_22161,N_27315);
nor U38495 (N_38495,N_22905,N_20929);
nor U38496 (N_38496,N_28824,N_21263);
and U38497 (N_38497,N_21694,N_23092);
xor U38498 (N_38498,N_22760,N_20964);
nor U38499 (N_38499,N_29044,N_23223);
nand U38500 (N_38500,N_21304,N_20358);
and U38501 (N_38501,N_22641,N_23395);
or U38502 (N_38502,N_21174,N_25350);
xor U38503 (N_38503,N_21234,N_25224);
xnor U38504 (N_38504,N_25301,N_28179);
or U38505 (N_38505,N_26784,N_27019);
and U38506 (N_38506,N_23358,N_23598);
xor U38507 (N_38507,N_25021,N_25773);
nor U38508 (N_38508,N_20897,N_20633);
nand U38509 (N_38509,N_25316,N_28177);
and U38510 (N_38510,N_26840,N_29897);
or U38511 (N_38511,N_24882,N_29814);
or U38512 (N_38512,N_27058,N_29229);
nor U38513 (N_38513,N_25913,N_29496);
nor U38514 (N_38514,N_24976,N_23279);
nand U38515 (N_38515,N_28778,N_29469);
nor U38516 (N_38516,N_25724,N_29560);
nor U38517 (N_38517,N_27803,N_20997);
or U38518 (N_38518,N_23745,N_29797);
nand U38519 (N_38519,N_28408,N_27600);
nor U38520 (N_38520,N_29053,N_25496);
xnor U38521 (N_38521,N_29135,N_26966);
nor U38522 (N_38522,N_21398,N_26159);
nand U38523 (N_38523,N_20485,N_27982);
xor U38524 (N_38524,N_20892,N_21640);
and U38525 (N_38525,N_22818,N_26977);
and U38526 (N_38526,N_22291,N_23054);
xor U38527 (N_38527,N_22507,N_26366);
xnor U38528 (N_38528,N_23127,N_23565);
nor U38529 (N_38529,N_22409,N_22915);
and U38530 (N_38530,N_26940,N_23161);
xor U38531 (N_38531,N_25232,N_20015);
nand U38532 (N_38532,N_24771,N_29184);
or U38533 (N_38533,N_24423,N_27568);
xor U38534 (N_38534,N_20223,N_24366);
xnor U38535 (N_38535,N_23161,N_27780);
and U38536 (N_38536,N_28517,N_26235);
nand U38537 (N_38537,N_20627,N_27613);
or U38538 (N_38538,N_21549,N_28305);
xor U38539 (N_38539,N_20456,N_25071);
nand U38540 (N_38540,N_26942,N_24783);
nor U38541 (N_38541,N_24096,N_20595);
and U38542 (N_38542,N_25084,N_24449);
nor U38543 (N_38543,N_25353,N_23526);
xor U38544 (N_38544,N_25822,N_21522);
or U38545 (N_38545,N_20214,N_20479);
or U38546 (N_38546,N_27986,N_23572);
nand U38547 (N_38547,N_24334,N_24436);
nand U38548 (N_38548,N_22228,N_27513);
and U38549 (N_38549,N_26871,N_24687);
xor U38550 (N_38550,N_28647,N_27067);
and U38551 (N_38551,N_29698,N_24632);
or U38552 (N_38552,N_21850,N_24647);
nor U38553 (N_38553,N_26309,N_27426);
or U38554 (N_38554,N_28187,N_23483);
xor U38555 (N_38555,N_24650,N_22455);
xnor U38556 (N_38556,N_25181,N_27679);
nor U38557 (N_38557,N_28850,N_20145);
nor U38558 (N_38558,N_24126,N_27991);
or U38559 (N_38559,N_22276,N_22067);
and U38560 (N_38560,N_25106,N_22796);
or U38561 (N_38561,N_29543,N_27515);
or U38562 (N_38562,N_24397,N_26271);
nand U38563 (N_38563,N_20174,N_21682);
and U38564 (N_38564,N_23856,N_29067);
nand U38565 (N_38565,N_28762,N_23242);
nand U38566 (N_38566,N_23188,N_20114);
and U38567 (N_38567,N_26697,N_27569);
xnor U38568 (N_38568,N_20326,N_29804);
or U38569 (N_38569,N_23412,N_22535);
xnor U38570 (N_38570,N_20436,N_24619);
nor U38571 (N_38571,N_20127,N_25605);
xor U38572 (N_38572,N_27360,N_21298);
xnor U38573 (N_38573,N_26165,N_21461);
nor U38574 (N_38574,N_20362,N_29025);
or U38575 (N_38575,N_26479,N_26113);
and U38576 (N_38576,N_23399,N_27441);
nand U38577 (N_38577,N_23457,N_28253);
and U38578 (N_38578,N_21079,N_28772);
nor U38579 (N_38579,N_29298,N_28442);
or U38580 (N_38580,N_29182,N_25830);
and U38581 (N_38581,N_28571,N_24109);
and U38582 (N_38582,N_28194,N_27684);
nor U38583 (N_38583,N_24483,N_25794);
nor U38584 (N_38584,N_29932,N_25883);
and U38585 (N_38585,N_24338,N_26226);
and U38586 (N_38586,N_21722,N_28043);
nand U38587 (N_38587,N_27092,N_21978);
or U38588 (N_38588,N_21929,N_24787);
xor U38589 (N_38589,N_28270,N_28643);
nor U38590 (N_38590,N_22164,N_21723);
or U38591 (N_38591,N_25561,N_22978);
nand U38592 (N_38592,N_21978,N_27336);
xor U38593 (N_38593,N_22853,N_27547);
or U38594 (N_38594,N_25339,N_25535);
nor U38595 (N_38595,N_25633,N_25573);
nand U38596 (N_38596,N_25130,N_22335);
xnor U38597 (N_38597,N_20855,N_26896);
or U38598 (N_38598,N_23718,N_29983);
and U38599 (N_38599,N_27681,N_20594);
nor U38600 (N_38600,N_29359,N_23903);
nor U38601 (N_38601,N_23262,N_21316);
xnor U38602 (N_38602,N_21178,N_23351);
xor U38603 (N_38603,N_21140,N_22149);
nor U38604 (N_38604,N_28744,N_29249);
nand U38605 (N_38605,N_29347,N_25681);
nand U38606 (N_38606,N_26893,N_27833);
xor U38607 (N_38607,N_25270,N_24220);
or U38608 (N_38608,N_20598,N_26810);
and U38609 (N_38609,N_25992,N_22837);
or U38610 (N_38610,N_29625,N_28308);
or U38611 (N_38611,N_27064,N_27754);
nor U38612 (N_38612,N_20412,N_23683);
and U38613 (N_38613,N_26030,N_24404);
and U38614 (N_38614,N_27103,N_25250);
nor U38615 (N_38615,N_25406,N_24338);
xor U38616 (N_38616,N_27440,N_29721);
and U38617 (N_38617,N_28360,N_27529);
xnor U38618 (N_38618,N_20194,N_27768);
or U38619 (N_38619,N_20619,N_23028);
or U38620 (N_38620,N_24198,N_28028);
and U38621 (N_38621,N_28440,N_26455);
xor U38622 (N_38622,N_22320,N_27833);
nor U38623 (N_38623,N_21497,N_28371);
nor U38624 (N_38624,N_28595,N_22692);
and U38625 (N_38625,N_20313,N_27646);
nor U38626 (N_38626,N_27304,N_24513);
and U38627 (N_38627,N_23893,N_28885);
nor U38628 (N_38628,N_24360,N_23192);
nor U38629 (N_38629,N_22189,N_20963);
and U38630 (N_38630,N_29419,N_26290);
nor U38631 (N_38631,N_25651,N_21191);
xor U38632 (N_38632,N_28498,N_21882);
nor U38633 (N_38633,N_20991,N_23596);
and U38634 (N_38634,N_25482,N_26758);
or U38635 (N_38635,N_24145,N_21948);
and U38636 (N_38636,N_29801,N_21283);
or U38637 (N_38637,N_26779,N_26961);
or U38638 (N_38638,N_21318,N_24663);
and U38639 (N_38639,N_28306,N_27943);
or U38640 (N_38640,N_28295,N_20749);
xor U38641 (N_38641,N_23769,N_27847);
or U38642 (N_38642,N_22321,N_25260);
or U38643 (N_38643,N_23241,N_24354);
or U38644 (N_38644,N_26019,N_25223);
nor U38645 (N_38645,N_21833,N_20709);
xor U38646 (N_38646,N_27842,N_20738);
nor U38647 (N_38647,N_20613,N_28208);
nor U38648 (N_38648,N_25378,N_27918);
nand U38649 (N_38649,N_20523,N_22559);
and U38650 (N_38650,N_25972,N_21785);
nor U38651 (N_38651,N_23041,N_25130);
nor U38652 (N_38652,N_25939,N_27927);
and U38653 (N_38653,N_27687,N_25182);
and U38654 (N_38654,N_27640,N_26142);
nor U38655 (N_38655,N_26369,N_27410);
nor U38656 (N_38656,N_28417,N_20566);
nor U38657 (N_38657,N_23224,N_29122);
and U38658 (N_38658,N_28807,N_23819);
and U38659 (N_38659,N_20418,N_21647);
or U38660 (N_38660,N_26983,N_21482);
xor U38661 (N_38661,N_24558,N_22485);
nand U38662 (N_38662,N_23331,N_26180);
and U38663 (N_38663,N_20399,N_29943);
nor U38664 (N_38664,N_25137,N_20325);
xor U38665 (N_38665,N_29104,N_24991);
xor U38666 (N_38666,N_21539,N_21543);
nand U38667 (N_38667,N_21757,N_26467);
nor U38668 (N_38668,N_22151,N_26758);
nand U38669 (N_38669,N_29475,N_26900);
xor U38670 (N_38670,N_27347,N_23843);
or U38671 (N_38671,N_20155,N_29717);
or U38672 (N_38672,N_21245,N_20879);
nand U38673 (N_38673,N_28190,N_25525);
xor U38674 (N_38674,N_26954,N_28419);
nand U38675 (N_38675,N_22985,N_25160);
nand U38676 (N_38676,N_25206,N_25502);
xor U38677 (N_38677,N_21080,N_28433);
xor U38678 (N_38678,N_28052,N_20649);
and U38679 (N_38679,N_20227,N_25306);
or U38680 (N_38680,N_26541,N_21344);
nand U38681 (N_38681,N_27038,N_27583);
or U38682 (N_38682,N_29455,N_29186);
nor U38683 (N_38683,N_26429,N_25281);
or U38684 (N_38684,N_21576,N_27999);
and U38685 (N_38685,N_27827,N_25521);
nand U38686 (N_38686,N_26075,N_21400);
xor U38687 (N_38687,N_24433,N_25857);
nand U38688 (N_38688,N_25377,N_25988);
or U38689 (N_38689,N_27526,N_24232);
nor U38690 (N_38690,N_27304,N_29791);
nor U38691 (N_38691,N_29006,N_21351);
nand U38692 (N_38692,N_21636,N_22674);
nor U38693 (N_38693,N_26291,N_20600);
xnor U38694 (N_38694,N_26879,N_26277);
and U38695 (N_38695,N_21681,N_20843);
xnor U38696 (N_38696,N_20951,N_23380);
nand U38697 (N_38697,N_21256,N_24913);
nor U38698 (N_38698,N_28835,N_20233);
and U38699 (N_38699,N_28794,N_20373);
and U38700 (N_38700,N_25149,N_28815);
and U38701 (N_38701,N_23279,N_23624);
xor U38702 (N_38702,N_26956,N_26503);
nand U38703 (N_38703,N_26768,N_23440);
nor U38704 (N_38704,N_28715,N_29677);
and U38705 (N_38705,N_20697,N_27844);
nand U38706 (N_38706,N_26000,N_26237);
nand U38707 (N_38707,N_21959,N_24545);
nand U38708 (N_38708,N_23511,N_22231);
or U38709 (N_38709,N_28275,N_28702);
or U38710 (N_38710,N_23337,N_29396);
nand U38711 (N_38711,N_22564,N_21054);
and U38712 (N_38712,N_28253,N_23124);
nor U38713 (N_38713,N_24726,N_24377);
or U38714 (N_38714,N_24525,N_27878);
xnor U38715 (N_38715,N_22978,N_25697);
nand U38716 (N_38716,N_26609,N_21336);
and U38717 (N_38717,N_24933,N_26732);
nand U38718 (N_38718,N_22620,N_24309);
nor U38719 (N_38719,N_24854,N_28118);
xnor U38720 (N_38720,N_25159,N_21448);
nor U38721 (N_38721,N_20770,N_22813);
nand U38722 (N_38722,N_28221,N_27520);
and U38723 (N_38723,N_28946,N_22391);
nor U38724 (N_38724,N_21754,N_28573);
or U38725 (N_38725,N_24563,N_28010);
or U38726 (N_38726,N_20199,N_23782);
and U38727 (N_38727,N_21134,N_28620);
xor U38728 (N_38728,N_24800,N_26241);
xor U38729 (N_38729,N_28180,N_25160);
nand U38730 (N_38730,N_25556,N_23992);
or U38731 (N_38731,N_22982,N_20229);
xnor U38732 (N_38732,N_21676,N_20646);
or U38733 (N_38733,N_26889,N_29226);
nor U38734 (N_38734,N_20207,N_20001);
xor U38735 (N_38735,N_27499,N_28344);
or U38736 (N_38736,N_25469,N_25586);
or U38737 (N_38737,N_29196,N_22636);
or U38738 (N_38738,N_24438,N_23009);
xnor U38739 (N_38739,N_24431,N_20103);
xor U38740 (N_38740,N_21974,N_25328);
nand U38741 (N_38741,N_22969,N_21098);
or U38742 (N_38742,N_27421,N_25514);
xor U38743 (N_38743,N_25675,N_20094);
and U38744 (N_38744,N_23283,N_24422);
xor U38745 (N_38745,N_25176,N_27342);
nand U38746 (N_38746,N_27438,N_29257);
nand U38747 (N_38747,N_23352,N_22824);
and U38748 (N_38748,N_28604,N_25982);
xnor U38749 (N_38749,N_22160,N_27991);
nand U38750 (N_38750,N_28656,N_21854);
xor U38751 (N_38751,N_23449,N_22816);
nand U38752 (N_38752,N_29740,N_26556);
and U38753 (N_38753,N_20548,N_29430);
nand U38754 (N_38754,N_22127,N_27205);
or U38755 (N_38755,N_27021,N_24358);
xnor U38756 (N_38756,N_28639,N_21566);
and U38757 (N_38757,N_20362,N_21307);
or U38758 (N_38758,N_23381,N_29900);
xor U38759 (N_38759,N_23416,N_24015);
xnor U38760 (N_38760,N_24927,N_21569);
and U38761 (N_38761,N_27578,N_28128);
xnor U38762 (N_38762,N_28651,N_29335);
and U38763 (N_38763,N_23467,N_24830);
or U38764 (N_38764,N_26752,N_27748);
and U38765 (N_38765,N_27028,N_21053);
nor U38766 (N_38766,N_22174,N_29636);
or U38767 (N_38767,N_20696,N_25436);
nor U38768 (N_38768,N_22415,N_20555);
or U38769 (N_38769,N_21041,N_20298);
and U38770 (N_38770,N_20544,N_29903);
nor U38771 (N_38771,N_28132,N_29264);
xor U38772 (N_38772,N_20505,N_27675);
or U38773 (N_38773,N_21226,N_25372);
xor U38774 (N_38774,N_28812,N_27917);
or U38775 (N_38775,N_24979,N_29022);
and U38776 (N_38776,N_29337,N_26550);
or U38777 (N_38777,N_22201,N_29830);
or U38778 (N_38778,N_25691,N_26710);
nor U38779 (N_38779,N_21005,N_22160);
nand U38780 (N_38780,N_28614,N_26258);
nand U38781 (N_38781,N_25692,N_20280);
nand U38782 (N_38782,N_20790,N_23110);
and U38783 (N_38783,N_22115,N_26817);
nor U38784 (N_38784,N_29348,N_25089);
or U38785 (N_38785,N_22902,N_27237);
nor U38786 (N_38786,N_20020,N_28634);
nand U38787 (N_38787,N_20309,N_27293);
and U38788 (N_38788,N_22918,N_26975);
nand U38789 (N_38789,N_29431,N_21432);
nor U38790 (N_38790,N_28954,N_25135);
nand U38791 (N_38791,N_20953,N_20400);
nor U38792 (N_38792,N_21929,N_26411);
xor U38793 (N_38793,N_28902,N_26272);
xnor U38794 (N_38794,N_23804,N_26888);
and U38795 (N_38795,N_28618,N_28660);
xnor U38796 (N_38796,N_29099,N_22738);
nor U38797 (N_38797,N_28889,N_24079);
and U38798 (N_38798,N_27271,N_27299);
nand U38799 (N_38799,N_29881,N_26441);
nor U38800 (N_38800,N_27703,N_25582);
nor U38801 (N_38801,N_26149,N_26344);
nand U38802 (N_38802,N_21595,N_22560);
and U38803 (N_38803,N_21956,N_22014);
and U38804 (N_38804,N_27700,N_23626);
or U38805 (N_38805,N_26349,N_26847);
or U38806 (N_38806,N_24845,N_21063);
nand U38807 (N_38807,N_26149,N_22868);
nand U38808 (N_38808,N_22606,N_20838);
nand U38809 (N_38809,N_26811,N_24995);
nor U38810 (N_38810,N_27794,N_23759);
or U38811 (N_38811,N_24346,N_25361);
nand U38812 (N_38812,N_29598,N_25117);
or U38813 (N_38813,N_21970,N_28758);
and U38814 (N_38814,N_28911,N_26962);
nor U38815 (N_38815,N_21860,N_29350);
or U38816 (N_38816,N_26209,N_22475);
or U38817 (N_38817,N_24521,N_20437);
or U38818 (N_38818,N_22795,N_28520);
and U38819 (N_38819,N_23622,N_25398);
or U38820 (N_38820,N_28243,N_24137);
and U38821 (N_38821,N_28048,N_24414);
and U38822 (N_38822,N_26680,N_22406);
and U38823 (N_38823,N_23044,N_22535);
nand U38824 (N_38824,N_22537,N_27231);
and U38825 (N_38825,N_21165,N_26291);
nor U38826 (N_38826,N_23407,N_25193);
or U38827 (N_38827,N_25943,N_23497);
and U38828 (N_38828,N_29191,N_23513);
and U38829 (N_38829,N_29704,N_29271);
nand U38830 (N_38830,N_21675,N_25190);
or U38831 (N_38831,N_24375,N_27962);
or U38832 (N_38832,N_29317,N_27952);
xnor U38833 (N_38833,N_26810,N_27330);
nand U38834 (N_38834,N_22146,N_28793);
xor U38835 (N_38835,N_27163,N_24087);
xnor U38836 (N_38836,N_23841,N_25824);
nor U38837 (N_38837,N_21535,N_21419);
and U38838 (N_38838,N_21041,N_28435);
or U38839 (N_38839,N_24782,N_24464);
xnor U38840 (N_38840,N_25332,N_20915);
xor U38841 (N_38841,N_25459,N_28392);
nand U38842 (N_38842,N_21953,N_29170);
nand U38843 (N_38843,N_27288,N_22082);
nor U38844 (N_38844,N_26767,N_21209);
nand U38845 (N_38845,N_29365,N_25474);
xnor U38846 (N_38846,N_21023,N_25898);
nand U38847 (N_38847,N_26146,N_28735);
and U38848 (N_38848,N_27584,N_26298);
nand U38849 (N_38849,N_27175,N_20587);
or U38850 (N_38850,N_22848,N_28193);
and U38851 (N_38851,N_21205,N_22924);
xnor U38852 (N_38852,N_20126,N_26832);
or U38853 (N_38853,N_27383,N_26752);
xor U38854 (N_38854,N_28276,N_24279);
xor U38855 (N_38855,N_26079,N_28572);
and U38856 (N_38856,N_25194,N_28345);
nand U38857 (N_38857,N_25182,N_21872);
nor U38858 (N_38858,N_24526,N_28634);
nor U38859 (N_38859,N_28573,N_25181);
xor U38860 (N_38860,N_29786,N_28816);
and U38861 (N_38861,N_29586,N_23027);
and U38862 (N_38862,N_23704,N_24169);
xor U38863 (N_38863,N_27472,N_20617);
nor U38864 (N_38864,N_20829,N_27679);
or U38865 (N_38865,N_24010,N_23167);
or U38866 (N_38866,N_29504,N_28391);
and U38867 (N_38867,N_20951,N_27706);
nand U38868 (N_38868,N_20999,N_29370);
xor U38869 (N_38869,N_23729,N_21194);
and U38870 (N_38870,N_28101,N_26017);
or U38871 (N_38871,N_25843,N_22294);
nand U38872 (N_38872,N_26648,N_26777);
or U38873 (N_38873,N_23196,N_27286);
or U38874 (N_38874,N_20689,N_24873);
and U38875 (N_38875,N_27163,N_22356);
xnor U38876 (N_38876,N_23889,N_23962);
xor U38877 (N_38877,N_21574,N_24001);
or U38878 (N_38878,N_29296,N_29189);
or U38879 (N_38879,N_25030,N_25675);
or U38880 (N_38880,N_20517,N_22848);
or U38881 (N_38881,N_20421,N_23801);
nand U38882 (N_38882,N_21143,N_22513);
and U38883 (N_38883,N_24521,N_28463);
xnor U38884 (N_38884,N_23996,N_22858);
nand U38885 (N_38885,N_27952,N_23460);
nand U38886 (N_38886,N_24341,N_24906);
xnor U38887 (N_38887,N_29272,N_27112);
xor U38888 (N_38888,N_25567,N_28272);
nand U38889 (N_38889,N_29214,N_20163);
xor U38890 (N_38890,N_20394,N_27762);
or U38891 (N_38891,N_28071,N_21318);
xnor U38892 (N_38892,N_20228,N_26868);
and U38893 (N_38893,N_20790,N_29297);
or U38894 (N_38894,N_23422,N_20693);
nand U38895 (N_38895,N_21233,N_24664);
nor U38896 (N_38896,N_27007,N_26918);
xnor U38897 (N_38897,N_29535,N_26046);
nor U38898 (N_38898,N_27830,N_24095);
or U38899 (N_38899,N_26240,N_29772);
or U38900 (N_38900,N_21684,N_26757);
nor U38901 (N_38901,N_29444,N_23116);
or U38902 (N_38902,N_21869,N_29151);
or U38903 (N_38903,N_22409,N_27873);
nor U38904 (N_38904,N_24798,N_26763);
nand U38905 (N_38905,N_25270,N_23587);
xnor U38906 (N_38906,N_29504,N_20802);
xnor U38907 (N_38907,N_20184,N_28839);
nor U38908 (N_38908,N_28320,N_27389);
nand U38909 (N_38909,N_20725,N_28371);
nand U38910 (N_38910,N_21987,N_25564);
nand U38911 (N_38911,N_26171,N_25927);
xor U38912 (N_38912,N_21341,N_22348);
nand U38913 (N_38913,N_20258,N_22940);
nand U38914 (N_38914,N_28982,N_24379);
and U38915 (N_38915,N_24128,N_20161);
or U38916 (N_38916,N_24603,N_26896);
and U38917 (N_38917,N_25585,N_20936);
nand U38918 (N_38918,N_22224,N_22072);
or U38919 (N_38919,N_20908,N_28062);
nor U38920 (N_38920,N_24211,N_29214);
and U38921 (N_38921,N_23025,N_22124);
or U38922 (N_38922,N_28334,N_22179);
nand U38923 (N_38923,N_27486,N_21504);
or U38924 (N_38924,N_21816,N_24350);
or U38925 (N_38925,N_23251,N_27027);
nand U38926 (N_38926,N_24842,N_23802);
xnor U38927 (N_38927,N_27392,N_20238);
nor U38928 (N_38928,N_25447,N_29704);
nor U38929 (N_38929,N_25526,N_22249);
nand U38930 (N_38930,N_20155,N_26184);
nor U38931 (N_38931,N_24100,N_29319);
or U38932 (N_38932,N_28196,N_25119);
or U38933 (N_38933,N_21217,N_28601);
xnor U38934 (N_38934,N_29185,N_24783);
and U38935 (N_38935,N_29714,N_26258);
and U38936 (N_38936,N_21525,N_28785);
and U38937 (N_38937,N_25510,N_20409);
nand U38938 (N_38938,N_26126,N_27490);
and U38939 (N_38939,N_22711,N_28409);
xor U38940 (N_38940,N_23691,N_28204);
nand U38941 (N_38941,N_28615,N_27916);
and U38942 (N_38942,N_24566,N_21580);
nor U38943 (N_38943,N_21121,N_28334);
or U38944 (N_38944,N_24800,N_23247);
or U38945 (N_38945,N_21799,N_21769);
and U38946 (N_38946,N_27600,N_20337);
and U38947 (N_38947,N_23518,N_22405);
and U38948 (N_38948,N_26984,N_28821);
nand U38949 (N_38949,N_27676,N_26639);
nand U38950 (N_38950,N_29487,N_21373);
or U38951 (N_38951,N_22791,N_27734);
or U38952 (N_38952,N_22152,N_22617);
nor U38953 (N_38953,N_23996,N_29997);
nand U38954 (N_38954,N_20908,N_26862);
or U38955 (N_38955,N_26494,N_24418);
nor U38956 (N_38956,N_29328,N_25262);
nor U38957 (N_38957,N_21837,N_26723);
and U38958 (N_38958,N_26723,N_29554);
nand U38959 (N_38959,N_28376,N_22799);
or U38960 (N_38960,N_25436,N_23394);
xor U38961 (N_38961,N_28740,N_24004);
and U38962 (N_38962,N_23901,N_24835);
xor U38963 (N_38963,N_29927,N_23953);
nor U38964 (N_38964,N_20498,N_25171);
or U38965 (N_38965,N_29663,N_25480);
xnor U38966 (N_38966,N_28082,N_24125);
nand U38967 (N_38967,N_21642,N_21787);
and U38968 (N_38968,N_29466,N_25366);
xor U38969 (N_38969,N_23392,N_29857);
nand U38970 (N_38970,N_25357,N_27529);
nand U38971 (N_38971,N_28215,N_25257);
xnor U38972 (N_38972,N_26131,N_26332);
nor U38973 (N_38973,N_27646,N_22557);
nor U38974 (N_38974,N_26105,N_21480);
nand U38975 (N_38975,N_29062,N_28650);
or U38976 (N_38976,N_20993,N_22264);
or U38977 (N_38977,N_28369,N_29759);
xor U38978 (N_38978,N_29374,N_25519);
nand U38979 (N_38979,N_29004,N_23003);
and U38980 (N_38980,N_26260,N_26787);
and U38981 (N_38981,N_27978,N_29756);
nand U38982 (N_38982,N_24925,N_20588);
nand U38983 (N_38983,N_20121,N_25776);
nand U38984 (N_38984,N_20091,N_23426);
nor U38985 (N_38985,N_22631,N_29470);
nand U38986 (N_38986,N_22740,N_22891);
nand U38987 (N_38987,N_27203,N_26943);
nand U38988 (N_38988,N_24051,N_29970);
or U38989 (N_38989,N_24039,N_26870);
or U38990 (N_38990,N_29625,N_22325);
nor U38991 (N_38991,N_28341,N_22273);
xor U38992 (N_38992,N_20453,N_29131);
nor U38993 (N_38993,N_29705,N_22092);
nand U38994 (N_38994,N_23359,N_27130);
nand U38995 (N_38995,N_27977,N_20918);
nand U38996 (N_38996,N_20872,N_29434);
and U38997 (N_38997,N_23358,N_24541);
and U38998 (N_38998,N_28074,N_22999);
and U38999 (N_38999,N_23898,N_22256);
nor U39000 (N_39000,N_25046,N_25824);
and U39001 (N_39001,N_21702,N_23917);
or U39002 (N_39002,N_29569,N_24363);
xor U39003 (N_39003,N_28824,N_23698);
nor U39004 (N_39004,N_26898,N_22666);
nand U39005 (N_39005,N_28016,N_25797);
and U39006 (N_39006,N_27524,N_29246);
xnor U39007 (N_39007,N_27596,N_21483);
xor U39008 (N_39008,N_29857,N_22020);
xor U39009 (N_39009,N_27482,N_27876);
xnor U39010 (N_39010,N_24568,N_23940);
and U39011 (N_39011,N_25673,N_21293);
and U39012 (N_39012,N_24204,N_21935);
and U39013 (N_39013,N_28448,N_26525);
nor U39014 (N_39014,N_24841,N_24303);
or U39015 (N_39015,N_23802,N_22341);
or U39016 (N_39016,N_20754,N_24074);
nor U39017 (N_39017,N_26141,N_21794);
and U39018 (N_39018,N_27801,N_25896);
xnor U39019 (N_39019,N_21144,N_22041);
nor U39020 (N_39020,N_22098,N_26870);
xor U39021 (N_39021,N_29778,N_21969);
nand U39022 (N_39022,N_25850,N_22035);
xor U39023 (N_39023,N_20879,N_23931);
nor U39024 (N_39024,N_26796,N_23991);
nand U39025 (N_39025,N_29360,N_22449);
or U39026 (N_39026,N_24695,N_23231);
xnor U39027 (N_39027,N_26434,N_20408);
nor U39028 (N_39028,N_29503,N_20961);
xor U39029 (N_39029,N_24766,N_22350);
xor U39030 (N_39030,N_25319,N_29191);
nand U39031 (N_39031,N_24952,N_27174);
xnor U39032 (N_39032,N_23158,N_27943);
nor U39033 (N_39033,N_23034,N_24317);
nor U39034 (N_39034,N_21690,N_28463);
and U39035 (N_39035,N_27009,N_28118);
nand U39036 (N_39036,N_25133,N_24823);
and U39037 (N_39037,N_26403,N_23904);
or U39038 (N_39038,N_29552,N_25887);
or U39039 (N_39039,N_20329,N_23835);
or U39040 (N_39040,N_23746,N_22971);
nor U39041 (N_39041,N_22728,N_22224);
or U39042 (N_39042,N_23109,N_29385);
nor U39043 (N_39043,N_29125,N_27367);
nand U39044 (N_39044,N_23903,N_27272);
and U39045 (N_39045,N_23019,N_29050);
xnor U39046 (N_39046,N_27439,N_25641);
xnor U39047 (N_39047,N_21341,N_20273);
or U39048 (N_39048,N_26954,N_21966);
nand U39049 (N_39049,N_22615,N_21037);
nand U39050 (N_39050,N_28165,N_27518);
nor U39051 (N_39051,N_23631,N_23186);
xnor U39052 (N_39052,N_22436,N_21382);
nor U39053 (N_39053,N_21911,N_22730);
and U39054 (N_39054,N_28518,N_26375);
and U39055 (N_39055,N_25727,N_28366);
nand U39056 (N_39056,N_21081,N_29705);
nor U39057 (N_39057,N_26452,N_24896);
xor U39058 (N_39058,N_29971,N_28440);
nand U39059 (N_39059,N_20300,N_24956);
nor U39060 (N_39060,N_27733,N_29092);
nor U39061 (N_39061,N_20928,N_24222);
and U39062 (N_39062,N_21417,N_20365);
and U39063 (N_39063,N_21767,N_23097);
or U39064 (N_39064,N_21345,N_22021);
xor U39065 (N_39065,N_26668,N_25526);
nor U39066 (N_39066,N_25287,N_23038);
xnor U39067 (N_39067,N_29356,N_23229);
or U39068 (N_39068,N_23554,N_24592);
nor U39069 (N_39069,N_25153,N_24122);
nor U39070 (N_39070,N_25531,N_22513);
nand U39071 (N_39071,N_21112,N_26046);
xor U39072 (N_39072,N_24582,N_27566);
nor U39073 (N_39073,N_20088,N_22523);
xor U39074 (N_39074,N_26977,N_25943);
and U39075 (N_39075,N_26020,N_21400);
nor U39076 (N_39076,N_29063,N_23989);
and U39077 (N_39077,N_28430,N_24601);
and U39078 (N_39078,N_25338,N_27947);
or U39079 (N_39079,N_26405,N_21906);
and U39080 (N_39080,N_20506,N_28574);
nand U39081 (N_39081,N_21236,N_25917);
nor U39082 (N_39082,N_27395,N_22723);
nand U39083 (N_39083,N_27238,N_21972);
xnor U39084 (N_39084,N_25108,N_21340);
or U39085 (N_39085,N_29200,N_24996);
and U39086 (N_39086,N_28407,N_20561);
and U39087 (N_39087,N_24502,N_22143);
nor U39088 (N_39088,N_24956,N_20506);
or U39089 (N_39089,N_29496,N_23989);
or U39090 (N_39090,N_23157,N_20217);
xor U39091 (N_39091,N_29977,N_20463);
nand U39092 (N_39092,N_23322,N_29619);
xnor U39093 (N_39093,N_29050,N_20147);
xnor U39094 (N_39094,N_23236,N_28902);
xor U39095 (N_39095,N_27570,N_21797);
or U39096 (N_39096,N_22205,N_28803);
xor U39097 (N_39097,N_24300,N_24156);
nand U39098 (N_39098,N_21908,N_26268);
nand U39099 (N_39099,N_22298,N_25250);
nor U39100 (N_39100,N_25478,N_28055);
xor U39101 (N_39101,N_22064,N_21209);
or U39102 (N_39102,N_25264,N_20477);
and U39103 (N_39103,N_21975,N_21804);
or U39104 (N_39104,N_25468,N_28826);
and U39105 (N_39105,N_26743,N_29387);
or U39106 (N_39106,N_21383,N_26756);
and U39107 (N_39107,N_28003,N_29258);
xor U39108 (N_39108,N_22076,N_24665);
and U39109 (N_39109,N_22645,N_28282);
nand U39110 (N_39110,N_22587,N_21229);
xor U39111 (N_39111,N_21208,N_29410);
nor U39112 (N_39112,N_28212,N_29857);
nand U39113 (N_39113,N_26335,N_24322);
nand U39114 (N_39114,N_27674,N_25877);
nand U39115 (N_39115,N_24568,N_21995);
xor U39116 (N_39116,N_25748,N_29126);
xnor U39117 (N_39117,N_26944,N_29787);
xor U39118 (N_39118,N_29788,N_22284);
nand U39119 (N_39119,N_21899,N_20149);
xnor U39120 (N_39120,N_27809,N_29571);
nor U39121 (N_39121,N_29872,N_27229);
and U39122 (N_39122,N_26116,N_27215);
nor U39123 (N_39123,N_25223,N_28838);
xor U39124 (N_39124,N_25497,N_21068);
xnor U39125 (N_39125,N_21413,N_28937);
nand U39126 (N_39126,N_28811,N_26455);
and U39127 (N_39127,N_22190,N_24274);
or U39128 (N_39128,N_26203,N_24231);
nor U39129 (N_39129,N_21688,N_25330);
xor U39130 (N_39130,N_21533,N_28848);
or U39131 (N_39131,N_20757,N_23816);
and U39132 (N_39132,N_23858,N_22558);
xor U39133 (N_39133,N_24404,N_27507);
nor U39134 (N_39134,N_24005,N_28051);
xnor U39135 (N_39135,N_28174,N_23399);
or U39136 (N_39136,N_24576,N_26732);
and U39137 (N_39137,N_21487,N_24271);
nor U39138 (N_39138,N_26781,N_21990);
and U39139 (N_39139,N_29251,N_28688);
nand U39140 (N_39140,N_26528,N_29704);
nor U39141 (N_39141,N_23207,N_28527);
nand U39142 (N_39142,N_26938,N_22498);
nor U39143 (N_39143,N_20367,N_24453);
xor U39144 (N_39144,N_28979,N_21939);
and U39145 (N_39145,N_28372,N_25153);
and U39146 (N_39146,N_23339,N_21289);
xnor U39147 (N_39147,N_24100,N_22265);
nand U39148 (N_39148,N_28852,N_26174);
nand U39149 (N_39149,N_29077,N_25822);
and U39150 (N_39150,N_23804,N_20353);
and U39151 (N_39151,N_26580,N_24522);
or U39152 (N_39152,N_27733,N_24789);
nand U39153 (N_39153,N_25396,N_27550);
xor U39154 (N_39154,N_21296,N_23720);
nor U39155 (N_39155,N_24604,N_26370);
xnor U39156 (N_39156,N_26451,N_20101);
or U39157 (N_39157,N_22474,N_20293);
nor U39158 (N_39158,N_21882,N_26240);
or U39159 (N_39159,N_23583,N_21988);
or U39160 (N_39160,N_23772,N_27352);
and U39161 (N_39161,N_29370,N_29711);
nor U39162 (N_39162,N_25882,N_22373);
and U39163 (N_39163,N_20937,N_21078);
nand U39164 (N_39164,N_26359,N_26395);
xnor U39165 (N_39165,N_26436,N_22058);
or U39166 (N_39166,N_27193,N_27318);
nand U39167 (N_39167,N_25016,N_26800);
or U39168 (N_39168,N_29200,N_24457);
nor U39169 (N_39169,N_21454,N_22095);
nand U39170 (N_39170,N_20564,N_26929);
xor U39171 (N_39171,N_21620,N_29541);
nor U39172 (N_39172,N_25238,N_23136);
or U39173 (N_39173,N_29504,N_21611);
nor U39174 (N_39174,N_20782,N_23332);
nand U39175 (N_39175,N_23185,N_28095);
xor U39176 (N_39176,N_22337,N_26396);
and U39177 (N_39177,N_21927,N_20316);
or U39178 (N_39178,N_22315,N_29329);
nand U39179 (N_39179,N_27903,N_20106);
or U39180 (N_39180,N_20680,N_24107);
nand U39181 (N_39181,N_26475,N_29120);
and U39182 (N_39182,N_26679,N_28689);
xnor U39183 (N_39183,N_27966,N_29845);
nand U39184 (N_39184,N_21397,N_21377);
or U39185 (N_39185,N_25933,N_25148);
or U39186 (N_39186,N_26112,N_23270);
or U39187 (N_39187,N_24838,N_27924);
nor U39188 (N_39188,N_26716,N_21388);
nor U39189 (N_39189,N_28296,N_24443);
and U39190 (N_39190,N_27792,N_21740);
nor U39191 (N_39191,N_28481,N_20764);
or U39192 (N_39192,N_28592,N_22531);
or U39193 (N_39193,N_25155,N_21199);
nor U39194 (N_39194,N_20857,N_24290);
nor U39195 (N_39195,N_24516,N_21381);
nand U39196 (N_39196,N_20973,N_23493);
and U39197 (N_39197,N_26986,N_27557);
xor U39198 (N_39198,N_23627,N_22609);
nand U39199 (N_39199,N_25630,N_21478);
nand U39200 (N_39200,N_26132,N_20868);
nor U39201 (N_39201,N_27474,N_27817);
nor U39202 (N_39202,N_27206,N_29516);
and U39203 (N_39203,N_24914,N_21878);
xnor U39204 (N_39204,N_20935,N_20678);
xor U39205 (N_39205,N_26846,N_25176);
nor U39206 (N_39206,N_24369,N_22654);
xnor U39207 (N_39207,N_27227,N_27485);
or U39208 (N_39208,N_20204,N_25203);
xnor U39209 (N_39209,N_23285,N_24609);
or U39210 (N_39210,N_27525,N_23888);
nand U39211 (N_39211,N_23234,N_24619);
xor U39212 (N_39212,N_28994,N_22751);
xnor U39213 (N_39213,N_21780,N_22585);
or U39214 (N_39214,N_27335,N_29512);
and U39215 (N_39215,N_26083,N_21212);
xor U39216 (N_39216,N_20943,N_29491);
or U39217 (N_39217,N_21546,N_20432);
nor U39218 (N_39218,N_29850,N_23255);
and U39219 (N_39219,N_26945,N_26334);
nor U39220 (N_39220,N_27053,N_24062);
nor U39221 (N_39221,N_23989,N_23954);
nand U39222 (N_39222,N_25175,N_29313);
nand U39223 (N_39223,N_25626,N_24615);
nor U39224 (N_39224,N_20605,N_28855);
or U39225 (N_39225,N_26249,N_22178);
nand U39226 (N_39226,N_27945,N_23531);
xor U39227 (N_39227,N_29544,N_22397);
nand U39228 (N_39228,N_21083,N_25558);
and U39229 (N_39229,N_21594,N_25571);
xnor U39230 (N_39230,N_24963,N_24988);
nor U39231 (N_39231,N_25924,N_28659);
xnor U39232 (N_39232,N_21061,N_26354);
nor U39233 (N_39233,N_22603,N_22944);
nor U39234 (N_39234,N_21079,N_27630);
xor U39235 (N_39235,N_28241,N_26511);
nand U39236 (N_39236,N_27758,N_24265);
and U39237 (N_39237,N_21956,N_24235);
nor U39238 (N_39238,N_25649,N_20609);
and U39239 (N_39239,N_24182,N_28300);
nand U39240 (N_39240,N_20267,N_27770);
nor U39241 (N_39241,N_26585,N_27347);
and U39242 (N_39242,N_22377,N_24883);
nand U39243 (N_39243,N_29593,N_23021);
and U39244 (N_39244,N_20201,N_28268);
xor U39245 (N_39245,N_24855,N_20141);
or U39246 (N_39246,N_26620,N_20216);
and U39247 (N_39247,N_26433,N_25731);
or U39248 (N_39248,N_24564,N_23789);
xnor U39249 (N_39249,N_27716,N_28757);
xnor U39250 (N_39250,N_21755,N_25119);
xor U39251 (N_39251,N_21170,N_25832);
and U39252 (N_39252,N_27238,N_26649);
and U39253 (N_39253,N_29442,N_29169);
or U39254 (N_39254,N_22241,N_25774);
nand U39255 (N_39255,N_23595,N_28249);
xnor U39256 (N_39256,N_27816,N_26635);
nand U39257 (N_39257,N_29176,N_28502);
and U39258 (N_39258,N_21688,N_22675);
xnor U39259 (N_39259,N_25145,N_24033);
xor U39260 (N_39260,N_21902,N_25074);
nand U39261 (N_39261,N_28667,N_27277);
nor U39262 (N_39262,N_21564,N_29322);
nand U39263 (N_39263,N_21072,N_23521);
nor U39264 (N_39264,N_27915,N_28610);
nand U39265 (N_39265,N_20188,N_28397);
nor U39266 (N_39266,N_23192,N_25903);
nor U39267 (N_39267,N_28522,N_27210);
xor U39268 (N_39268,N_24306,N_27539);
nand U39269 (N_39269,N_20574,N_26955);
xor U39270 (N_39270,N_24128,N_25053);
nand U39271 (N_39271,N_28169,N_25862);
or U39272 (N_39272,N_29732,N_22044);
xnor U39273 (N_39273,N_28027,N_22632);
nand U39274 (N_39274,N_21119,N_21170);
xnor U39275 (N_39275,N_28871,N_27398);
or U39276 (N_39276,N_25440,N_24350);
nor U39277 (N_39277,N_29339,N_21782);
or U39278 (N_39278,N_26575,N_24927);
and U39279 (N_39279,N_25583,N_28075);
xnor U39280 (N_39280,N_28127,N_25191);
and U39281 (N_39281,N_24766,N_24656);
nand U39282 (N_39282,N_21503,N_28137);
nor U39283 (N_39283,N_25845,N_25870);
and U39284 (N_39284,N_27852,N_22356);
or U39285 (N_39285,N_28877,N_24707);
and U39286 (N_39286,N_26007,N_27773);
nand U39287 (N_39287,N_27237,N_28297);
nand U39288 (N_39288,N_25817,N_22401);
nand U39289 (N_39289,N_23483,N_22005);
nand U39290 (N_39290,N_26507,N_25288);
nand U39291 (N_39291,N_20162,N_20673);
and U39292 (N_39292,N_23522,N_21476);
or U39293 (N_39293,N_26829,N_25246);
nand U39294 (N_39294,N_23550,N_28276);
xnor U39295 (N_39295,N_25619,N_29852);
nor U39296 (N_39296,N_29784,N_24115);
and U39297 (N_39297,N_28573,N_22416);
and U39298 (N_39298,N_24644,N_29519);
nor U39299 (N_39299,N_24632,N_21375);
or U39300 (N_39300,N_20438,N_20332);
or U39301 (N_39301,N_25701,N_27538);
or U39302 (N_39302,N_29816,N_20114);
nor U39303 (N_39303,N_28682,N_29413);
and U39304 (N_39304,N_23627,N_20421);
or U39305 (N_39305,N_24643,N_21353);
and U39306 (N_39306,N_25728,N_22344);
xor U39307 (N_39307,N_23466,N_24297);
nor U39308 (N_39308,N_23549,N_29859);
nor U39309 (N_39309,N_20046,N_29943);
and U39310 (N_39310,N_29136,N_23898);
xnor U39311 (N_39311,N_20909,N_28301);
nor U39312 (N_39312,N_27381,N_29230);
or U39313 (N_39313,N_26533,N_26913);
nand U39314 (N_39314,N_23446,N_20397);
or U39315 (N_39315,N_23148,N_22217);
xnor U39316 (N_39316,N_24394,N_23939);
nand U39317 (N_39317,N_20642,N_25992);
nand U39318 (N_39318,N_20158,N_21965);
xnor U39319 (N_39319,N_22930,N_28324);
xnor U39320 (N_39320,N_20889,N_26580);
xor U39321 (N_39321,N_22028,N_20202);
xnor U39322 (N_39322,N_25190,N_24293);
or U39323 (N_39323,N_22823,N_29499);
xor U39324 (N_39324,N_23890,N_26964);
nand U39325 (N_39325,N_23177,N_26516);
xor U39326 (N_39326,N_22091,N_22941);
nor U39327 (N_39327,N_29484,N_27005);
xor U39328 (N_39328,N_27021,N_25546);
or U39329 (N_39329,N_26880,N_23726);
nand U39330 (N_39330,N_27692,N_23507);
nor U39331 (N_39331,N_27484,N_29129);
and U39332 (N_39332,N_26944,N_25876);
xor U39333 (N_39333,N_20373,N_29234);
nor U39334 (N_39334,N_21669,N_28913);
or U39335 (N_39335,N_21333,N_26261);
nor U39336 (N_39336,N_21630,N_24486);
and U39337 (N_39337,N_26036,N_29924);
xnor U39338 (N_39338,N_22207,N_21627);
or U39339 (N_39339,N_23632,N_29921);
or U39340 (N_39340,N_22123,N_23961);
xnor U39341 (N_39341,N_21897,N_27075);
nand U39342 (N_39342,N_20811,N_24797);
nand U39343 (N_39343,N_22952,N_27661);
xnor U39344 (N_39344,N_28676,N_22961);
and U39345 (N_39345,N_27675,N_23099);
xor U39346 (N_39346,N_25515,N_20301);
and U39347 (N_39347,N_25473,N_21550);
nor U39348 (N_39348,N_25566,N_24266);
and U39349 (N_39349,N_27774,N_27440);
nor U39350 (N_39350,N_28987,N_20464);
or U39351 (N_39351,N_27607,N_20336);
nand U39352 (N_39352,N_28006,N_22751);
or U39353 (N_39353,N_28576,N_25203);
nor U39354 (N_39354,N_28894,N_21351);
xor U39355 (N_39355,N_20653,N_20194);
nor U39356 (N_39356,N_20290,N_28082);
nand U39357 (N_39357,N_25490,N_20863);
xor U39358 (N_39358,N_24847,N_28455);
nand U39359 (N_39359,N_28309,N_20667);
and U39360 (N_39360,N_25072,N_25222);
nand U39361 (N_39361,N_21792,N_29727);
nor U39362 (N_39362,N_23125,N_22215);
nor U39363 (N_39363,N_23108,N_25618);
and U39364 (N_39364,N_28893,N_26749);
nor U39365 (N_39365,N_21653,N_28968);
nor U39366 (N_39366,N_23618,N_26596);
nand U39367 (N_39367,N_22431,N_26862);
nor U39368 (N_39368,N_25054,N_21200);
or U39369 (N_39369,N_27938,N_29471);
xor U39370 (N_39370,N_24409,N_22502);
and U39371 (N_39371,N_24358,N_24765);
nand U39372 (N_39372,N_20748,N_20677);
xor U39373 (N_39373,N_20952,N_20618);
nor U39374 (N_39374,N_22643,N_28500);
nor U39375 (N_39375,N_20623,N_28414);
nor U39376 (N_39376,N_24424,N_22969);
nand U39377 (N_39377,N_23012,N_28362);
nand U39378 (N_39378,N_24209,N_24257);
and U39379 (N_39379,N_26462,N_26047);
or U39380 (N_39380,N_20218,N_26482);
xor U39381 (N_39381,N_24893,N_20059);
and U39382 (N_39382,N_27784,N_24571);
xor U39383 (N_39383,N_27355,N_22482);
and U39384 (N_39384,N_28738,N_22235);
xnor U39385 (N_39385,N_29332,N_25928);
nand U39386 (N_39386,N_25032,N_25174);
and U39387 (N_39387,N_29641,N_28804);
xor U39388 (N_39388,N_24313,N_25232);
and U39389 (N_39389,N_21550,N_27989);
and U39390 (N_39390,N_26261,N_21893);
or U39391 (N_39391,N_22738,N_29915);
and U39392 (N_39392,N_21352,N_29822);
nor U39393 (N_39393,N_29975,N_23437);
nand U39394 (N_39394,N_20422,N_25771);
nand U39395 (N_39395,N_21974,N_27019);
or U39396 (N_39396,N_29973,N_28481);
and U39397 (N_39397,N_20121,N_21828);
nand U39398 (N_39398,N_24394,N_24559);
xor U39399 (N_39399,N_22917,N_28094);
nand U39400 (N_39400,N_28965,N_21436);
xor U39401 (N_39401,N_27369,N_26843);
nor U39402 (N_39402,N_26456,N_27569);
nand U39403 (N_39403,N_27152,N_20347);
or U39404 (N_39404,N_29938,N_25868);
xor U39405 (N_39405,N_21886,N_22827);
nand U39406 (N_39406,N_27616,N_21081);
nor U39407 (N_39407,N_29677,N_22918);
xor U39408 (N_39408,N_21211,N_29098);
and U39409 (N_39409,N_25977,N_28132);
and U39410 (N_39410,N_29082,N_20401);
and U39411 (N_39411,N_20015,N_29743);
nand U39412 (N_39412,N_29224,N_20369);
nor U39413 (N_39413,N_29077,N_20874);
nor U39414 (N_39414,N_23028,N_21891);
nand U39415 (N_39415,N_24134,N_22088);
xnor U39416 (N_39416,N_27787,N_23084);
xnor U39417 (N_39417,N_27158,N_24914);
and U39418 (N_39418,N_22948,N_21344);
nand U39419 (N_39419,N_21401,N_28467);
xor U39420 (N_39420,N_20961,N_27919);
or U39421 (N_39421,N_25926,N_22059);
or U39422 (N_39422,N_21089,N_28150);
nand U39423 (N_39423,N_25123,N_21953);
or U39424 (N_39424,N_21138,N_29412);
and U39425 (N_39425,N_28569,N_21214);
or U39426 (N_39426,N_25998,N_25282);
xnor U39427 (N_39427,N_29755,N_22240);
and U39428 (N_39428,N_28041,N_26600);
xor U39429 (N_39429,N_24208,N_27731);
nor U39430 (N_39430,N_25268,N_23739);
nand U39431 (N_39431,N_29936,N_22726);
xnor U39432 (N_39432,N_28739,N_28980);
and U39433 (N_39433,N_20871,N_28108);
xnor U39434 (N_39434,N_21201,N_29207);
or U39435 (N_39435,N_29122,N_25422);
or U39436 (N_39436,N_23225,N_25540);
and U39437 (N_39437,N_27362,N_26875);
and U39438 (N_39438,N_20561,N_21638);
nand U39439 (N_39439,N_25325,N_20549);
or U39440 (N_39440,N_24856,N_29506);
nor U39441 (N_39441,N_20760,N_21102);
nand U39442 (N_39442,N_24933,N_29163);
and U39443 (N_39443,N_24533,N_24198);
xor U39444 (N_39444,N_25628,N_25311);
nor U39445 (N_39445,N_26334,N_22959);
nand U39446 (N_39446,N_25114,N_28929);
and U39447 (N_39447,N_26985,N_24146);
nor U39448 (N_39448,N_22632,N_28918);
nand U39449 (N_39449,N_27578,N_23703);
and U39450 (N_39450,N_24705,N_24284);
and U39451 (N_39451,N_26320,N_26558);
nor U39452 (N_39452,N_27652,N_28617);
nor U39453 (N_39453,N_26810,N_28976);
nand U39454 (N_39454,N_24201,N_25781);
or U39455 (N_39455,N_22644,N_28376);
xnor U39456 (N_39456,N_20150,N_28234);
nor U39457 (N_39457,N_20336,N_20390);
or U39458 (N_39458,N_28600,N_22753);
nor U39459 (N_39459,N_22673,N_21487);
or U39460 (N_39460,N_27423,N_23443);
xor U39461 (N_39461,N_20239,N_28644);
nand U39462 (N_39462,N_27240,N_21443);
nand U39463 (N_39463,N_27024,N_28127);
nand U39464 (N_39464,N_22598,N_23136);
nand U39465 (N_39465,N_20745,N_23787);
and U39466 (N_39466,N_27697,N_21440);
nand U39467 (N_39467,N_27043,N_26160);
or U39468 (N_39468,N_24259,N_29489);
xor U39469 (N_39469,N_20013,N_23391);
nand U39470 (N_39470,N_25036,N_23644);
or U39471 (N_39471,N_26257,N_21630);
or U39472 (N_39472,N_21536,N_25379);
nand U39473 (N_39473,N_23208,N_21716);
or U39474 (N_39474,N_29387,N_24506);
nor U39475 (N_39475,N_20451,N_29524);
nor U39476 (N_39476,N_29249,N_29721);
xor U39477 (N_39477,N_29248,N_29482);
or U39478 (N_39478,N_25331,N_26762);
nand U39479 (N_39479,N_28975,N_26611);
xor U39480 (N_39480,N_20162,N_20401);
and U39481 (N_39481,N_27210,N_21461);
nand U39482 (N_39482,N_23201,N_20798);
xnor U39483 (N_39483,N_24335,N_21057);
and U39484 (N_39484,N_29932,N_27058);
or U39485 (N_39485,N_28107,N_22963);
and U39486 (N_39486,N_26474,N_23439);
and U39487 (N_39487,N_29754,N_26448);
and U39488 (N_39488,N_24452,N_27295);
or U39489 (N_39489,N_22279,N_29864);
nand U39490 (N_39490,N_21610,N_22137);
xnor U39491 (N_39491,N_29160,N_29539);
xnor U39492 (N_39492,N_27504,N_25050);
xnor U39493 (N_39493,N_22424,N_27987);
or U39494 (N_39494,N_21893,N_22325);
nand U39495 (N_39495,N_28649,N_24142);
or U39496 (N_39496,N_26931,N_23619);
nor U39497 (N_39497,N_22936,N_29280);
nand U39498 (N_39498,N_29339,N_26372);
xnor U39499 (N_39499,N_21672,N_23150);
and U39500 (N_39500,N_24091,N_24225);
nand U39501 (N_39501,N_24672,N_23116);
nand U39502 (N_39502,N_23916,N_27236);
xor U39503 (N_39503,N_20596,N_20812);
or U39504 (N_39504,N_26956,N_23943);
xnor U39505 (N_39505,N_23218,N_29583);
or U39506 (N_39506,N_25512,N_26144);
or U39507 (N_39507,N_28165,N_21740);
and U39508 (N_39508,N_26186,N_20764);
nor U39509 (N_39509,N_28111,N_24029);
xnor U39510 (N_39510,N_27527,N_24357);
xor U39511 (N_39511,N_20073,N_21697);
nor U39512 (N_39512,N_27537,N_26347);
nand U39513 (N_39513,N_22769,N_25262);
or U39514 (N_39514,N_25986,N_27464);
nand U39515 (N_39515,N_26269,N_28475);
xnor U39516 (N_39516,N_26475,N_25995);
xor U39517 (N_39517,N_28019,N_27536);
nor U39518 (N_39518,N_23989,N_20175);
nand U39519 (N_39519,N_29425,N_23008);
nor U39520 (N_39520,N_24944,N_24193);
nand U39521 (N_39521,N_28923,N_29180);
and U39522 (N_39522,N_28315,N_21396);
nor U39523 (N_39523,N_29797,N_21988);
nand U39524 (N_39524,N_22946,N_24494);
nand U39525 (N_39525,N_26004,N_27487);
xor U39526 (N_39526,N_29535,N_26674);
or U39527 (N_39527,N_23844,N_25925);
or U39528 (N_39528,N_25130,N_29956);
nor U39529 (N_39529,N_27679,N_21726);
or U39530 (N_39530,N_26077,N_23437);
nand U39531 (N_39531,N_25575,N_25262);
or U39532 (N_39532,N_27344,N_21039);
or U39533 (N_39533,N_29006,N_29065);
and U39534 (N_39534,N_23008,N_23924);
nor U39535 (N_39535,N_20928,N_20800);
and U39536 (N_39536,N_25342,N_22997);
xnor U39537 (N_39537,N_21344,N_26109);
nand U39538 (N_39538,N_23310,N_29001);
nand U39539 (N_39539,N_23521,N_20882);
and U39540 (N_39540,N_24303,N_21002);
xnor U39541 (N_39541,N_29919,N_24514);
and U39542 (N_39542,N_26512,N_27343);
nand U39543 (N_39543,N_26726,N_29837);
nor U39544 (N_39544,N_22170,N_27834);
xor U39545 (N_39545,N_29881,N_23108);
and U39546 (N_39546,N_20354,N_21659);
and U39547 (N_39547,N_26769,N_27925);
and U39548 (N_39548,N_28443,N_28466);
and U39549 (N_39549,N_26192,N_20567);
nor U39550 (N_39550,N_25001,N_26449);
nand U39551 (N_39551,N_23636,N_29452);
xnor U39552 (N_39552,N_25541,N_21551);
or U39553 (N_39553,N_22670,N_26952);
and U39554 (N_39554,N_25595,N_24045);
xor U39555 (N_39555,N_29059,N_29681);
nand U39556 (N_39556,N_29330,N_28904);
xnor U39557 (N_39557,N_22067,N_29469);
xor U39558 (N_39558,N_26011,N_25754);
and U39559 (N_39559,N_26679,N_21359);
xor U39560 (N_39560,N_20599,N_26690);
and U39561 (N_39561,N_23559,N_20780);
xnor U39562 (N_39562,N_21818,N_28314);
and U39563 (N_39563,N_26021,N_26434);
nand U39564 (N_39564,N_29486,N_23300);
or U39565 (N_39565,N_28207,N_25963);
or U39566 (N_39566,N_23669,N_25001);
and U39567 (N_39567,N_27574,N_28575);
and U39568 (N_39568,N_22357,N_23603);
or U39569 (N_39569,N_22945,N_24803);
nor U39570 (N_39570,N_21015,N_25113);
nand U39571 (N_39571,N_23637,N_24198);
xor U39572 (N_39572,N_22053,N_28802);
and U39573 (N_39573,N_26928,N_24044);
xor U39574 (N_39574,N_23445,N_21921);
xor U39575 (N_39575,N_20756,N_27628);
nand U39576 (N_39576,N_20629,N_25518);
and U39577 (N_39577,N_21545,N_23912);
nor U39578 (N_39578,N_29965,N_24112);
and U39579 (N_39579,N_29858,N_20952);
xor U39580 (N_39580,N_29928,N_24650);
xnor U39581 (N_39581,N_21192,N_27622);
and U39582 (N_39582,N_28208,N_20968);
nor U39583 (N_39583,N_28801,N_26477);
or U39584 (N_39584,N_20844,N_28040);
xnor U39585 (N_39585,N_27876,N_26517);
xnor U39586 (N_39586,N_27780,N_29947);
nor U39587 (N_39587,N_23558,N_24285);
nor U39588 (N_39588,N_20336,N_24375);
nand U39589 (N_39589,N_27135,N_26979);
or U39590 (N_39590,N_26377,N_20092);
or U39591 (N_39591,N_28711,N_27956);
or U39592 (N_39592,N_24148,N_20228);
nor U39593 (N_39593,N_26832,N_29918);
or U39594 (N_39594,N_29248,N_22322);
or U39595 (N_39595,N_21343,N_27388);
nor U39596 (N_39596,N_20762,N_26867);
nor U39597 (N_39597,N_26774,N_25367);
or U39598 (N_39598,N_23088,N_20029);
xnor U39599 (N_39599,N_23272,N_23393);
or U39600 (N_39600,N_21382,N_27599);
nand U39601 (N_39601,N_24275,N_20280);
xor U39602 (N_39602,N_27748,N_25845);
nand U39603 (N_39603,N_28116,N_21838);
or U39604 (N_39604,N_28450,N_20945);
or U39605 (N_39605,N_21118,N_22152);
nor U39606 (N_39606,N_26683,N_24429);
or U39607 (N_39607,N_25217,N_28720);
or U39608 (N_39608,N_20743,N_25466);
nor U39609 (N_39609,N_24119,N_26785);
or U39610 (N_39610,N_26435,N_26500);
xor U39611 (N_39611,N_24689,N_23523);
or U39612 (N_39612,N_23602,N_28413);
nor U39613 (N_39613,N_28090,N_22960);
or U39614 (N_39614,N_26961,N_20066);
nand U39615 (N_39615,N_26243,N_28523);
nor U39616 (N_39616,N_29355,N_23298);
and U39617 (N_39617,N_26578,N_22806);
xnor U39618 (N_39618,N_23440,N_26067);
nor U39619 (N_39619,N_22450,N_28269);
or U39620 (N_39620,N_26003,N_24643);
or U39621 (N_39621,N_24255,N_25183);
nor U39622 (N_39622,N_22968,N_27777);
or U39623 (N_39623,N_20773,N_27734);
nand U39624 (N_39624,N_23327,N_20439);
nand U39625 (N_39625,N_26573,N_23741);
xnor U39626 (N_39626,N_23652,N_25045);
and U39627 (N_39627,N_23287,N_22764);
and U39628 (N_39628,N_20804,N_21655);
xor U39629 (N_39629,N_28951,N_23394);
nand U39630 (N_39630,N_24155,N_28802);
or U39631 (N_39631,N_24536,N_27194);
and U39632 (N_39632,N_22395,N_22353);
and U39633 (N_39633,N_26927,N_29459);
and U39634 (N_39634,N_21852,N_22796);
nor U39635 (N_39635,N_25985,N_21488);
or U39636 (N_39636,N_29591,N_21575);
xor U39637 (N_39637,N_24702,N_20890);
nand U39638 (N_39638,N_22742,N_29351);
nand U39639 (N_39639,N_23513,N_21428);
or U39640 (N_39640,N_29587,N_24312);
nand U39641 (N_39641,N_23245,N_20632);
and U39642 (N_39642,N_27189,N_25399);
or U39643 (N_39643,N_27375,N_21641);
and U39644 (N_39644,N_29097,N_24384);
nor U39645 (N_39645,N_29348,N_23666);
nor U39646 (N_39646,N_23313,N_20243);
nand U39647 (N_39647,N_26059,N_20961);
and U39648 (N_39648,N_27834,N_28794);
nand U39649 (N_39649,N_24784,N_20641);
nor U39650 (N_39650,N_26259,N_20598);
nand U39651 (N_39651,N_20349,N_28176);
nor U39652 (N_39652,N_21908,N_25315);
and U39653 (N_39653,N_25549,N_21498);
nand U39654 (N_39654,N_26953,N_28504);
xnor U39655 (N_39655,N_24908,N_22495);
nor U39656 (N_39656,N_25792,N_21640);
nand U39657 (N_39657,N_22221,N_23201);
nand U39658 (N_39658,N_27181,N_21151);
nor U39659 (N_39659,N_23581,N_27263);
nand U39660 (N_39660,N_28251,N_26114);
xor U39661 (N_39661,N_25434,N_28719);
or U39662 (N_39662,N_20520,N_29336);
or U39663 (N_39663,N_20872,N_24335);
nor U39664 (N_39664,N_29708,N_26824);
nor U39665 (N_39665,N_27616,N_22237);
nor U39666 (N_39666,N_22209,N_23492);
and U39667 (N_39667,N_24220,N_25869);
or U39668 (N_39668,N_28366,N_28743);
nor U39669 (N_39669,N_23469,N_23201);
or U39670 (N_39670,N_28062,N_27253);
xor U39671 (N_39671,N_26476,N_28832);
and U39672 (N_39672,N_25489,N_23573);
nor U39673 (N_39673,N_21511,N_22065);
or U39674 (N_39674,N_25534,N_20104);
nand U39675 (N_39675,N_23579,N_26930);
nor U39676 (N_39676,N_27119,N_21471);
nand U39677 (N_39677,N_22240,N_25843);
xnor U39678 (N_39678,N_20278,N_21757);
xnor U39679 (N_39679,N_26518,N_24517);
nand U39680 (N_39680,N_26963,N_24719);
and U39681 (N_39681,N_22854,N_23202);
nor U39682 (N_39682,N_21328,N_22933);
or U39683 (N_39683,N_21458,N_29730);
or U39684 (N_39684,N_23365,N_20032);
nor U39685 (N_39685,N_27731,N_20164);
or U39686 (N_39686,N_27137,N_25448);
xnor U39687 (N_39687,N_21042,N_21617);
nand U39688 (N_39688,N_22155,N_26089);
xor U39689 (N_39689,N_28572,N_27284);
xor U39690 (N_39690,N_27501,N_29182);
nor U39691 (N_39691,N_28446,N_25570);
and U39692 (N_39692,N_28036,N_21492);
nand U39693 (N_39693,N_29854,N_24530);
nor U39694 (N_39694,N_21842,N_25187);
xnor U39695 (N_39695,N_24804,N_27095);
xnor U39696 (N_39696,N_28150,N_22758);
nor U39697 (N_39697,N_20949,N_24527);
nor U39698 (N_39698,N_29901,N_24566);
and U39699 (N_39699,N_23263,N_28197);
and U39700 (N_39700,N_28232,N_23531);
xor U39701 (N_39701,N_25998,N_21720);
and U39702 (N_39702,N_28988,N_21190);
nand U39703 (N_39703,N_27561,N_24815);
nor U39704 (N_39704,N_22593,N_23572);
and U39705 (N_39705,N_29257,N_28404);
xor U39706 (N_39706,N_20077,N_23322);
and U39707 (N_39707,N_26068,N_20946);
or U39708 (N_39708,N_22356,N_21044);
and U39709 (N_39709,N_26205,N_22812);
or U39710 (N_39710,N_23122,N_29462);
and U39711 (N_39711,N_25917,N_24497);
xor U39712 (N_39712,N_26773,N_26728);
or U39713 (N_39713,N_27081,N_21158);
or U39714 (N_39714,N_24988,N_21917);
xnor U39715 (N_39715,N_29497,N_26373);
or U39716 (N_39716,N_23975,N_21702);
and U39717 (N_39717,N_22238,N_27294);
nand U39718 (N_39718,N_20565,N_21244);
nand U39719 (N_39719,N_22213,N_29684);
nand U39720 (N_39720,N_27776,N_26268);
and U39721 (N_39721,N_25015,N_27163);
or U39722 (N_39722,N_23919,N_21018);
or U39723 (N_39723,N_23662,N_25872);
xnor U39724 (N_39724,N_27178,N_26550);
nand U39725 (N_39725,N_28922,N_23171);
and U39726 (N_39726,N_21182,N_28711);
nand U39727 (N_39727,N_26786,N_25844);
nor U39728 (N_39728,N_29393,N_21110);
nor U39729 (N_39729,N_27049,N_26481);
nor U39730 (N_39730,N_29667,N_26736);
nor U39731 (N_39731,N_29515,N_25635);
nand U39732 (N_39732,N_25871,N_22463);
or U39733 (N_39733,N_28170,N_24740);
and U39734 (N_39734,N_26703,N_27466);
nor U39735 (N_39735,N_25443,N_20021);
and U39736 (N_39736,N_27293,N_29906);
xnor U39737 (N_39737,N_26730,N_26505);
and U39738 (N_39738,N_26764,N_22366);
nor U39739 (N_39739,N_25959,N_26976);
nor U39740 (N_39740,N_27626,N_26006);
or U39741 (N_39741,N_26789,N_21838);
nor U39742 (N_39742,N_21376,N_24448);
nand U39743 (N_39743,N_21223,N_22068);
nand U39744 (N_39744,N_25505,N_24587);
nor U39745 (N_39745,N_20715,N_29735);
or U39746 (N_39746,N_21348,N_26794);
xnor U39747 (N_39747,N_24005,N_22742);
xor U39748 (N_39748,N_21493,N_27118);
nand U39749 (N_39749,N_28025,N_28085);
xnor U39750 (N_39750,N_23453,N_22772);
and U39751 (N_39751,N_22046,N_28518);
and U39752 (N_39752,N_26529,N_29782);
xor U39753 (N_39753,N_20093,N_29030);
nand U39754 (N_39754,N_21688,N_26330);
xnor U39755 (N_39755,N_26353,N_21356);
nor U39756 (N_39756,N_20085,N_20608);
and U39757 (N_39757,N_26459,N_20986);
xnor U39758 (N_39758,N_27403,N_21119);
xor U39759 (N_39759,N_23542,N_28782);
nor U39760 (N_39760,N_27643,N_25942);
xnor U39761 (N_39761,N_22721,N_21709);
nor U39762 (N_39762,N_26438,N_27743);
xor U39763 (N_39763,N_25896,N_22758);
or U39764 (N_39764,N_25279,N_28859);
nand U39765 (N_39765,N_24617,N_21925);
xor U39766 (N_39766,N_23114,N_29251);
and U39767 (N_39767,N_24699,N_21735);
xnor U39768 (N_39768,N_26722,N_20983);
and U39769 (N_39769,N_28361,N_27294);
or U39770 (N_39770,N_25645,N_24374);
nor U39771 (N_39771,N_20207,N_25865);
nor U39772 (N_39772,N_24227,N_23762);
xor U39773 (N_39773,N_22612,N_21499);
xnor U39774 (N_39774,N_26209,N_24069);
nor U39775 (N_39775,N_22939,N_29542);
nand U39776 (N_39776,N_29361,N_23382);
nand U39777 (N_39777,N_26966,N_23860);
and U39778 (N_39778,N_28348,N_23000);
nand U39779 (N_39779,N_27059,N_21826);
xor U39780 (N_39780,N_26600,N_20430);
nor U39781 (N_39781,N_24969,N_26824);
or U39782 (N_39782,N_24678,N_23311);
nor U39783 (N_39783,N_21959,N_24585);
or U39784 (N_39784,N_25458,N_25966);
nor U39785 (N_39785,N_23829,N_28136);
and U39786 (N_39786,N_23595,N_26183);
xnor U39787 (N_39787,N_20296,N_29413);
or U39788 (N_39788,N_27655,N_23715);
xnor U39789 (N_39789,N_21007,N_27714);
nand U39790 (N_39790,N_20628,N_29848);
and U39791 (N_39791,N_21067,N_29979);
nand U39792 (N_39792,N_26909,N_20440);
nand U39793 (N_39793,N_27650,N_25433);
xor U39794 (N_39794,N_25374,N_26638);
and U39795 (N_39795,N_25528,N_27839);
or U39796 (N_39796,N_20248,N_22645);
or U39797 (N_39797,N_27943,N_23712);
and U39798 (N_39798,N_25628,N_25503);
nor U39799 (N_39799,N_22560,N_25095);
xor U39800 (N_39800,N_21201,N_25470);
nor U39801 (N_39801,N_22612,N_22292);
xor U39802 (N_39802,N_22790,N_23245);
xnor U39803 (N_39803,N_27767,N_28532);
xnor U39804 (N_39804,N_28249,N_22596);
or U39805 (N_39805,N_24281,N_24491);
and U39806 (N_39806,N_27376,N_26666);
nand U39807 (N_39807,N_22539,N_29045);
or U39808 (N_39808,N_25156,N_24923);
xor U39809 (N_39809,N_24413,N_27104);
xnor U39810 (N_39810,N_27873,N_27301);
or U39811 (N_39811,N_29440,N_24215);
nor U39812 (N_39812,N_21327,N_24652);
xnor U39813 (N_39813,N_22088,N_24314);
nand U39814 (N_39814,N_24654,N_25124);
nor U39815 (N_39815,N_29742,N_21711);
nand U39816 (N_39816,N_24393,N_27949);
nor U39817 (N_39817,N_25969,N_28679);
nand U39818 (N_39818,N_24033,N_20535);
nor U39819 (N_39819,N_27383,N_29161);
and U39820 (N_39820,N_21354,N_26363);
xnor U39821 (N_39821,N_28328,N_24152);
and U39822 (N_39822,N_27655,N_29364);
or U39823 (N_39823,N_27820,N_24706);
nor U39824 (N_39824,N_28059,N_24816);
and U39825 (N_39825,N_28234,N_26020);
xnor U39826 (N_39826,N_20400,N_26981);
and U39827 (N_39827,N_27978,N_22384);
xor U39828 (N_39828,N_27487,N_27110);
nand U39829 (N_39829,N_25619,N_27542);
xnor U39830 (N_39830,N_25966,N_28977);
nor U39831 (N_39831,N_29020,N_23280);
and U39832 (N_39832,N_22088,N_24915);
nor U39833 (N_39833,N_24845,N_26943);
nand U39834 (N_39834,N_21251,N_24968);
and U39835 (N_39835,N_23311,N_23625);
nor U39836 (N_39836,N_23605,N_26982);
or U39837 (N_39837,N_26687,N_27497);
xnor U39838 (N_39838,N_24273,N_29530);
or U39839 (N_39839,N_25368,N_27232);
and U39840 (N_39840,N_27470,N_29823);
nand U39841 (N_39841,N_24803,N_26774);
nand U39842 (N_39842,N_20514,N_20161);
nand U39843 (N_39843,N_29533,N_29029);
and U39844 (N_39844,N_28103,N_23459);
or U39845 (N_39845,N_28556,N_20148);
xor U39846 (N_39846,N_26583,N_29916);
or U39847 (N_39847,N_25349,N_23544);
xor U39848 (N_39848,N_27428,N_26463);
or U39849 (N_39849,N_25186,N_29030);
xnor U39850 (N_39850,N_21923,N_26698);
or U39851 (N_39851,N_22114,N_23539);
nor U39852 (N_39852,N_22715,N_29575);
nand U39853 (N_39853,N_22075,N_26271);
and U39854 (N_39854,N_26794,N_22232);
nor U39855 (N_39855,N_28591,N_22602);
or U39856 (N_39856,N_28779,N_27649);
nor U39857 (N_39857,N_22674,N_21717);
nor U39858 (N_39858,N_28270,N_23935);
xnor U39859 (N_39859,N_24552,N_28869);
and U39860 (N_39860,N_23771,N_22793);
xnor U39861 (N_39861,N_22222,N_20356);
or U39862 (N_39862,N_29385,N_27511);
or U39863 (N_39863,N_20672,N_26433);
xnor U39864 (N_39864,N_23350,N_20264);
nor U39865 (N_39865,N_21386,N_20975);
nand U39866 (N_39866,N_22371,N_25519);
xnor U39867 (N_39867,N_29751,N_28436);
nand U39868 (N_39868,N_22409,N_29476);
xor U39869 (N_39869,N_26000,N_21387);
or U39870 (N_39870,N_20317,N_25665);
or U39871 (N_39871,N_22411,N_20751);
and U39872 (N_39872,N_25345,N_25038);
nand U39873 (N_39873,N_28541,N_24563);
nand U39874 (N_39874,N_25204,N_25709);
nor U39875 (N_39875,N_24561,N_27453);
and U39876 (N_39876,N_25075,N_29151);
nand U39877 (N_39877,N_26227,N_23588);
or U39878 (N_39878,N_26506,N_21647);
nor U39879 (N_39879,N_26286,N_20386);
nor U39880 (N_39880,N_29085,N_25189);
and U39881 (N_39881,N_22065,N_28064);
xor U39882 (N_39882,N_27955,N_28871);
xnor U39883 (N_39883,N_20842,N_28777);
and U39884 (N_39884,N_24442,N_26719);
nand U39885 (N_39885,N_29558,N_27613);
nand U39886 (N_39886,N_25060,N_24348);
or U39887 (N_39887,N_20835,N_20655);
xor U39888 (N_39888,N_22029,N_24422);
or U39889 (N_39889,N_21706,N_28809);
and U39890 (N_39890,N_24211,N_23863);
nand U39891 (N_39891,N_21312,N_20365);
and U39892 (N_39892,N_24951,N_20677);
xor U39893 (N_39893,N_29579,N_23281);
xnor U39894 (N_39894,N_23801,N_24303);
nor U39895 (N_39895,N_24278,N_29463);
nand U39896 (N_39896,N_23301,N_24177);
and U39897 (N_39897,N_28227,N_26330);
nand U39898 (N_39898,N_25634,N_27032);
nand U39899 (N_39899,N_29082,N_29961);
nand U39900 (N_39900,N_21519,N_22159);
nor U39901 (N_39901,N_24143,N_25941);
nand U39902 (N_39902,N_28833,N_22271);
or U39903 (N_39903,N_28252,N_25098);
and U39904 (N_39904,N_29883,N_25868);
nor U39905 (N_39905,N_26918,N_22364);
xnor U39906 (N_39906,N_27130,N_22604);
nand U39907 (N_39907,N_28825,N_21505);
and U39908 (N_39908,N_22515,N_22411);
nand U39909 (N_39909,N_25091,N_20617);
and U39910 (N_39910,N_28884,N_23494);
nand U39911 (N_39911,N_23192,N_26147);
and U39912 (N_39912,N_25125,N_29152);
and U39913 (N_39913,N_28123,N_29947);
or U39914 (N_39914,N_28254,N_28137);
or U39915 (N_39915,N_22601,N_24421);
nand U39916 (N_39916,N_26733,N_25421);
xnor U39917 (N_39917,N_25931,N_25455);
and U39918 (N_39918,N_23828,N_27510);
nand U39919 (N_39919,N_28648,N_21155);
xor U39920 (N_39920,N_26573,N_28864);
or U39921 (N_39921,N_26216,N_23623);
xor U39922 (N_39922,N_26189,N_24546);
and U39923 (N_39923,N_23328,N_21192);
and U39924 (N_39924,N_28681,N_20166);
xor U39925 (N_39925,N_22886,N_25995);
or U39926 (N_39926,N_25976,N_26424);
nand U39927 (N_39927,N_24625,N_29607);
or U39928 (N_39928,N_20566,N_26416);
nor U39929 (N_39929,N_28779,N_20100);
nor U39930 (N_39930,N_24209,N_24835);
or U39931 (N_39931,N_26717,N_25293);
and U39932 (N_39932,N_28890,N_22229);
or U39933 (N_39933,N_25405,N_23165);
or U39934 (N_39934,N_25732,N_22059);
nor U39935 (N_39935,N_25171,N_28546);
nor U39936 (N_39936,N_23129,N_25337);
xnor U39937 (N_39937,N_29611,N_23140);
xor U39938 (N_39938,N_29322,N_20624);
and U39939 (N_39939,N_28128,N_29433);
nand U39940 (N_39940,N_29401,N_26968);
or U39941 (N_39941,N_29418,N_28461);
and U39942 (N_39942,N_28754,N_20822);
nand U39943 (N_39943,N_29788,N_29687);
and U39944 (N_39944,N_22860,N_29904);
nand U39945 (N_39945,N_23286,N_23370);
or U39946 (N_39946,N_23490,N_21258);
nand U39947 (N_39947,N_24498,N_27732);
and U39948 (N_39948,N_22687,N_29432);
xnor U39949 (N_39949,N_29441,N_29957);
or U39950 (N_39950,N_29882,N_23145);
and U39951 (N_39951,N_25128,N_23761);
nand U39952 (N_39952,N_22265,N_28666);
and U39953 (N_39953,N_22428,N_26172);
nand U39954 (N_39954,N_27878,N_21134);
nor U39955 (N_39955,N_22584,N_21205);
nor U39956 (N_39956,N_21057,N_29440);
nor U39957 (N_39957,N_29470,N_26860);
or U39958 (N_39958,N_23409,N_25775);
xor U39959 (N_39959,N_28351,N_25174);
xor U39960 (N_39960,N_21100,N_23142);
nor U39961 (N_39961,N_29634,N_29512);
and U39962 (N_39962,N_23827,N_23140);
nor U39963 (N_39963,N_20346,N_22559);
nand U39964 (N_39964,N_26122,N_22831);
and U39965 (N_39965,N_26493,N_23576);
or U39966 (N_39966,N_25061,N_24466);
and U39967 (N_39967,N_22418,N_27652);
nand U39968 (N_39968,N_28199,N_25009);
xnor U39969 (N_39969,N_23766,N_22568);
xnor U39970 (N_39970,N_28752,N_28549);
or U39971 (N_39971,N_24709,N_27964);
nor U39972 (N_39972,N_23676,N_20579);
xnor U39973 (N_39973,N_21535,N_27604);
xor U39974 (N_39974,N_29889,N_23003);
or U39975 (N_39975,N_22184,N_25484);
and U39976 (N_39976,N_26152,N_22649);
nand U39977 (N_39977,N_22401,N_27011);
or U39978 (N_39978,N_26572,N_28603);
xnor U39979 (N_39979,N_28006,N_27735);
nand U39980 (N_39980,N_20602,N_28559);
nand U39981 (N_39981,N_27542,N_28638);
and U39982 (N_39982,N_24449,N_23173);
nor U39983 (N_39983,N_20095,N_25458);
nor U39984 (N_39984,N_26388,N_26827);
nand U39985 (N_39985,N_25654,N_28974);
and U39986 (N_39986,N_29338,N_20907);
and U39987 (N_39987,N_25584,N_20330);
and U39988 (N_39988,N_23029,N_29378);
nand U39989 (N_39989,N_20011,N_24040);
nand U39990 (N_39990,N_29503,N_28446);
xnor U39991 (N_39991,N_20198,N_20517);
and U39992 (N_39992,N_29625,N_27200);
nor U39993 (N_39993,N_28377,N_29962);
nand U39994 (N_39994,N_27354,N_23642);
nand U39995 (N_39995,N_26551,N_20295);
nor U39996 (N_39996,N_26532,N_21070);
nand U39997 (N_39997,N_27385,N_23321);
xnor U39998 (N_39998,N_20175,N_26056);
xor U39999 (N_39999,N_27000,N_29185);
nor U40000 (N_40000,N_31200,N_34982);
nand U40001 (N_40001,N_37369,N_30973);
or U40002 (N_40002,N_36183,N_38981);
and U40003 (N_40003,N_33008,N_35489);
nor U40004 (N_40004,N_38502,N_39145);
nand U40005 (N_40005,N_38027,N_35551);
nor U40006 (N_40006,N_34465,N_31079);
or U40007 (N_40007,N_35510,N_35618);
or U40008 (N_40008,N_31952,N_34218);
nand U40009 (N_40009,N_39226,N_35022);
and U40010 (N_40010,N_35784,N_39267);
or U40011 (N_40011,N_30408,N_32980);
and U40012 (N_40012,N_39628,N_32345);
nand U40013 (N_40013,N_34859,N_31787);
nand U40014 (N_40014,N_30981,N_34140);
nor U40015 (N_40015,N_35668,N_36964);
nor U40016 (N_40016,N_38052,N_31886);
and U40017 (N_40017,N_38221,N_32985);
and U40018 (N_40018,N_32979,N_37873);
or U40019 (N_40019,N_39564,N_34122);
nor U40020 (N_40020,N_30027,N_35805);
or U40021 (N_40021,N_36893,N_33286);
nand U40022 (N_40022,N_34346,N_30497);
nand U40023 (N_40023,N_39653,N_39565);
or U40024 (N_40024,N_38846,N_39197);
nand U40025 (N_40025,N_36093,N_32337);
xnor U40026 (N_40026,N_30582,N_38580);
and U40027 (N_40027,N_37843,N_30054);
nand U40028 (N_40028,N_33303,N_33032);
and U40029 (N_40029,N_38178,N_35928);
nor U40030 (N_40030,N_36648,N_33479);
xnor U40031 (N_40031,N_36220,N_38646);
nor U40032 (N_40032,N_35274,N_30307);
and U40033 (N_40033,N_36352,N_34498);
and U40034 (N_40034,N_35909,N_31915);
xor U40035 (N_40035,N_35925,N_38789);
nand U40036 (N_40036,N_38160,N_30227);
nand U40037 (N_40037,N_32615,N_31578);
nor U40038 (N_40038,N_39804,N_33381);
nand U40039 (N_40039,N_31209,N_34503);
and U40040 (N_40040,N_39613,N_37007);
nor U40041 (N_40041,N_37317,N_32503);
nand U40042 (N_40042,N_32565,N_36585);
nand U40043 (N_40043,N_33807,N_33680);
nor U40044 (N_40044,N_34413,N_31740);
xor U40045 (N_40045,N_39905,N_34713);
xor U40046 (N_40046,N_32784,N_35678);
nand U40047 (N_40047,N_36849,N_36588);
xor U40048 (N_40048,N_36187,N_37472);
and U40049 (N_40049,N_37959,N_38222);
xnor U40050 (N_40050,N_39797,N_36786);
xor U40051 (N_40051,N_30924,N_32425);
and U40052 (N_40052,N_33865,N_39160);
xor U40053 (N_40053,N_31705,N_38405);
nand U40054 (N_40054,N_33079,N_32636);
and U40055 (N_40055,N_37347,N_36767);
nand U40056 (N_40056,N_36025,N_33159);
xnor U40057 (N_40057,N_35082,N_33380);
nor U40058 (N_40058,N_38121,N_36682);
and U40059 (N_40059,N_32163,N_37449);
and U40060 (N_40060,N_30739,N_34221);
and U40061 (N_40061,N_30695,N_39987);
and U40062 (N_40062,N_34394,N_33369);
or U40063 (N_40063,N_31130,N_38835);
or U40064 (N_40064,N_38182,N_30690);
nand U40065 (N_40065,N_33267,N_32827);
or U40066 (N_40066,N_38584,N_39654);
or U40067 (N_40067,N_35964,N_32941);
nor U40068 (N_40068,N_37920,N_30637);
nor U40069 (N_40069,N_32710,N_35977);
and U40070 (N_40070,N_36481,N_34743);
xnor U40071 (N_40071,N_38251,N_38320);
nand U40072 (N_40072,N_37470,N_37571);
and U40073 (N_40073,N_37029,N_32222);
nand U40074 (N_40074,N_31711,N_30544);
xnor U40075 (N_40075,N_36185,N_33167);
nand U40076 (N_40076,N_33953,N_30671);
nor U40077 (N_40077,N_33900,N_33641);
nor U40078 (N_40078,N_36621,N_32690);
or U40079 (N_40079,N_31908,N_34078);
xnor U40080 (N_40080,N_30795,N_38073);
xor U40081 (N_40081,N_32706,N_36766);
nor U40082 (N_40082,N_39468,N_39580);
nor U40083 (N_40083,N_36542,N_38562);
and U40084 (N_40084,N_31172,N_30771);
nand U40085 (N_40085,N_38598,N_31272);
or U40086 (N_40086,N_39360,N_34044);
and U40087 (N_40087,N_38089,N_31728);
or U40088 (N_40088,N_30567,N_33270);
xor U40089 (N_40089,N_31628,N_32386);
or U40090 (N_40090,N_32878,N_33876);
xnor U40091 (N_40091,N_30630,N_35782);
nor U40092 (N_40092,N_30491,N_33040);
xnor U40093 (N_40093,N_34393,N_34883);
nor U40094 (N_40094,N_33868,N_36083);
or U40095 (N_40095,N_32803,N_35326);
xor U40096 (N_40096,N_38837,N_33986);
nand U40097 (N_40097,N_31790,N_30235);
xor U40098 (N_40098,N_30918,N_36781);
nand U40099 (N_40099,N_36644,N_36795);
or U40100 (N_40100,N_31599,N_38015);
and U40101 (N_40101,N_31005,N_33813);
nand U40102 (N_40102,N_38504,N_39415);
and U40103 (N_40103,N_37366,N_38613);
and U40104 (N_40104,N_35521,N_33170);
or U40105 (N_40105,N_33190,N_33098);
and U40106 (N_40106,N_38625,N_39984);
nor U40107 (N_40107,N_30500,N_31271);
or U40108 (N_40108,N_34478,N_31540);
xnor U40109 (N_40109,N_32852,N_34266);
xor U40110 (N_40110,N_39213,N_37821);
xor U40111 (N_40111,N_33587,N_37950);
and U40112 (N_40112,N_39029,N_35239);
and U40113 (N_40113,N_30167,N_36649);
and U40114 (N_40114,N_39394,N_34911);
nor U40115 (N_40115,N_38208,N_39132);
nor U40116 (N_40116,N_30681,N_35077);
or U40117 (N_40117,N_38334,N_39115);
xor U40118 (N_40118,N_33637,N_30756);
or U40119 (N_40119,N_36802,N_32914);
xnor U40120 (N_40120,N_30657,N_30745);
nand U40121 (N_40121,N_39273,N_36404);
xnor U40122 (N_40122,N_37953,N_34546);
and U40123 (N_40123,N_35089,N_31888);
xnor U40124 (N_40124,N_32007,N_33514);
and U40125 (N_40125,N_36854,N_33858);
xnor U40126 (N_40126,N_37636,N_32071);
or U40127 (N_40127,N_37324,N_33217);
nor U40128 (N_40128,N_34695,N_33921);
nand U40129 (N_40129,N_34572,N_39966);
or U40130 (N_40130,N_32483,N_31409);
xnor U40131 (N_40131,N_34702,N_35137);
or U40132 (N_40132,N_34967,N_35148);
and U40133 (N_40133,N_36527,N_35943);
nor U40134 (N_40134,N_39007,N_30705);
xnor U40135 (N_40135,N_39419,N_36623);
and U40136 (N_40136,N_31587,N_30653);
and U40137 (N_40137,N_32265,N_37424);
and U40138 (N_40138,N_30153,N_30996);
or U40139 (N_40139,N_34398,N_32667);
or U40140 (N_40140,N_34903,N_37010);
xor U40141 (N_40141,N_31820,N_32373);
and U40142 (N_40142,N_33423,N_33745);
and U40143 (N_40143,N_30203,N_31712);
nor U40144 (N_40144,N_37397,N_31563);
nor U40145 (N_40145,N_36656,N_36968);
nor U40146 (N_40146,N_34821,N_34952);
nor U40147 (N_40147,N_38751,N_35395);
xor U40148 (N_40148,N_39489,N_30737);
nand U40149 (N_40149,N_37591,N_32928);
and U40150 (N_40150,N_33545,N_31547);
or U40151 (N_40151,N_39340,N_37130);
nand U40152 (N_40152,N_31354,N_37274);
and U40153 (N_40153,N_36094,N_33864);
nand U40154 (N_40154,N_34583,N_37185);
nor U40155 (N_40155,N_31962,N_34048);
and U40156 (N_40156,N_32591,N_33259);
nor U40157 (N_40157,N_34373,N_30589);
xor U40158 (N_40158,N_30309,N_36713);
nor U40159 (N_40159,N_30724,N_30856);
nor U40160 (N_40160,N_36301,N_34388);
xor U40161 (N_40161,N_38002,N_37404);
or U40162 (N_40162,N_32095,N_37705);
or U40163 (N_40163,N_39519,N_39480);
nand U40164 (N_40164,N_38949,N_39182);
and U40165 (N_40165,N_37801,N_39546);
xor U40166 (N_40166,N_32216,N_31708);
xnor U40167 (N_40167,N_39586,N_35789);
or U40168 (N_40168,N_31045,N_38220);
or U40169 (N_40169,N_36023,N_32974);
or U40170 (N_40170,N_34097,N_30947);
nor U40171 (N_40171,N_36561,N_31286);
or U40172 (N_40172,N_39710,N_35992);
and U40173 (N_40173,N_38753,N_34231);
and U40174 (N_40174,N_30162,N_35453);
xnor U40175 (N_40175,N_33851,N_31054);
or U40176 (N_40176,N_35593,N_35216);
nand U40177 (N_40177,N_31604,N_33561);
nand U40178 (N_40178,N_34375,N_36941);
and U40179 (N_40179,N_32254,N_34772);
nand U40180 (N_40180,N_31610,N_35259);
or U40181 (N_40181,N_30905,N_31679);
and U40182 (N_40182,N_30257,N_30489);
and U40183 (N_40183,N_34654,N_31469);
nand U40184 (N_40184,N_33461,N_36919);
and U40185 (N_40185,N_31698,N_31710);
xor U40186 (N_40186,N_35336,N_39682);
xnor U40187 (N_40187,N_33172,N_39245);
or U40188 (N_40188,N_34685,N_35266);
nor U40189 (N_40189,N_35986,N_31407);
nor U40190 (N_40190,N_35529,N_37910);
xor U40191 (N_40191,N_30259,N_31458);
or U40192 (N_40192,N_38352,N_32211);
nor U40193 (N_40193,N_37878,N_38577);
and U40194 (N_40194,N_31828,N_37171);
xor U40195 (N_40195,N_37462,N_32574);
nand U40196 (N_40196,N_39951,N_34367);
nand U40197 (N_40197,N_37118,N_32282);
nand U40198 (N_40198,N_35778,N_31903);
xor U40199 (N_40199,N_30382,N_36653);
or U40200 (N_40200,N_38275,N_35276);
or U40201 (N_40201,N_37429,N_32610);
or U40202 (N_40202,N_35287,N_35217);
or U40203 (N_40203,N_38488,N_33766);
and U40204 (N_40204,N_38303,N_37524);
nand U40205 (N_40205,N_38711,N_33700);
xnor U40206 (N_40206,N_32444,N_38268);
nand U40207 (N_40207,N_32209,N_36909);
nand U40208 (N_40208,N_36006,N_31389);
nand U40209 (N_40209,N_38650,N_31012);
or U40210 (N_40210,N_35306,N_32634);
nor U40211 (N_40211,N_34604,N_38940);
nand U40212 (N_40212,N_33354,N_38219);
or U40213 (N_40213,N_37218,N_31373);
xnor U40214 (N_40214,N_30201,N_36333);
xor U40215 (N_40215,N_34189,N_34141);
or U40216 (N_40216,N_32837,N_33444);
nand U40217 (N_40217,N_39277,N_30777);
xor U40218 (N_40218,N_36855,N_30691);
or U40219 (N_40219,N_39610,N_39749);
nor U40220 (N_40220,N_35153,N_38771);
or U40221 (N_40221,N_38133,N_35588);
nor U40222 (N_40222,N_30999,N_39672);
nor U40223 (N_40223,N_37780,N_31117);
xnor U40224 (N_40224,N_33704,N_31572);
nand U40225 (N_40225,N_33201,N_37901);
xor U40226 (N_40226,N_34828,N_31185);
xnor U40227 (N_40227,N_39379,N_36271);
and U40228 (N_40228,N_33944,N_35172);
xnor U40229 (N_40229,N_38935,N_35008);
nor U40230 (N_40230,N_32724,N_39406);
xor U40231 (N_40231,N_37507,N_32056);
xor U40232 (N_40232,N_38954,N_31028);
nor U40233 (N_40233,N_37284,N_30110);
or U40234 (N_40234,N_39057,N_33243);
or U40235 (N_40235,N_33260,N_34247);
xor U40236 (N_40236,N_33186,N_33847);
nor U40237 (N_40237,N_35712,N_32664);
and U40238 (N_40238,N_32622,N_35779);
xor U40239 (N_40239,N_36759,N_33178);
nand U40240 (N_40240,N_36839,N_34721);
and U40241 (N_40241,N_32929,N_36138);
xnor U40242 (N_40242,N_35987,N_32896);
or U40243 (N_40243,N_30010,N_35398);
nand U40244 (N_40244,N_30868,N_30013);
nand U40245 (N_40245,N_32665,N_32795);
or U40246 (N_40246,N_35941,N_37802);
or U40247 (N_40247,N_30564,N_37501);
nor U40248 (N_40248,N_31143,N_37204);
nand U40249 (N_40249,N_35623,N_34165);
nand U40250 (N_40250,N_32934,N_31244);
or U40251 (N_40251,N_39673,N_35454);
and U40252 (N_40252,N_31967,N_36295);
nand U40253 (N_40253,N_34149,N_34423);
or U40254 (N_40254,N_34009,N_36632);
nor U40255 (N_40255,N_31279,N_30654);
or U40256 (N_40256,N_30772,N_30387);
and U40257 (N_40257,N_37476,N_35360);
nand U40258 (N_40258,N_38083,N_35114);
and U40259 (N_40259,N_39113,N_36077);
and U40260 (N_40260,N_36449,N_38541);
and U40261 (N_40261,N_39471,N_35702);
and U40262 (N_40262,N_35798,N_37673);
xor U40263 (N_40263,N_37653,N_35818);
xor U40264 (N_40264,N_33645,N_34178);
and U40265 (N_40265,N_31062,N_34219);
xnor U40266 (N_40266,N_37156,N_39879);
nor U40267 (N_40267,N_33878,N_32783);
nor U40268 (N_40268,N_35598,N_38399);
and U40269 (N_40269,N_38026,N_34853);
or U40270 (N_40270,N_36895,N_37083);
or U40271 (N_40271,N_30007,N_33211);
xnor U40272 (N_40272,N_36709,N_34244);
nand U40273 (N_40273,N_38462,N_36514);
or U40274 (N_40274,N_33279,N_39860);
or U40275 (N_40275,N_31731,N_31568);
nand U40276 (N_40276,N_30329,N_36190);
nand U40277 (N_40277,N_31529,N_35837);
or U40278 (N_40278,N_34961,N_33435);
or U40279 (N_40279,N_39956,N_30849);
nor U40280 (N_40280,N_37051,N_34310);
xnor U40281 (N_40281,N_35636,N_37893);
nand U40282 (N_40282,N_34723,N_30910);
or U40283 (N_40283,N_32383,N_31307);
and U40284 (N_40284,N_34698,N_35093);
nor U40285 (N_40285,N_35700,N_30244);
nor U40286 (N_40286,N_32108,N_33375);
nor U40287 (N_40287,N_39947,N_31894);
and U40288 (N_40288,N_35536,N_37818);
or U40289 (N_40289,N_30119,N_31614);
nand U40290 (N_40290,N_38469,N_32918);
or U40291 (N_40291,N_30289,N_33215);
and U40292 (N_40292,N_36060,N_34860);
xnor U40293 (N_40293,N_35099,N_31796);
nor U40294 (N_40294,N_37842,N_39412);
nand U40295 (N_40295,N_32192,N_37666);
nor U40296 (N_40296,N_32736,N_37278);
xor U40297 (N_40297,N_31589,N_30620);
nand U40298 (N_40298,N_35205,N_35751);
nand U40299 (N_40299,N_39618,N_34060);
or U40300 (N_40300,N_30149,N_31371);
or U40301 (N_40301,N_35955,N_30002);
xor U40302 (N_40302,N_36371,N_38226);
nor U40303 (N_40303,N_31672,N_33440);
nor U40304 (N_40304,N_35686,N_36834);
nor U40305 (N_40305,N_31717,N_35547);
or U40306 (N_40306,N_33465,N_35300);
nor U40307 (N_40307,N_30080,N_37048);
and U40308 (N_40308,N_37725,N_33432);
nand U40309 (N_40309,N_32335,N_33065);
nor U40310 (N_40310,N_32280,N_36901);
and U40311 (N_40311,N_33484,N_35182);
and U40312 (N_40312,N_34386,N_39961);
or U40313 (N_40313,N_36926,N_39402);
nor U40314 (N_40314,N_32332,N_36616);
or U40315 (N_40315,N_33036,N_31619);
nand U40316 (N_40316,N_34443,N_31817);
xor U40317 (N_40317,N_33742,N_36646);
or U40318 (N_40318,N_35029,N_30135);
nand U40319 (N_40319,N_32704,N_39025);
nor U40320 (N_40320,N_36873,N_37327);
or U40321 (N_40321,N_32291,N_35476);
xnor U40322 (N_40322,N_38156,N_35797);
xnor U40323 (N_40323,N_30262,N_31632);
and U40324 (N_40324,N_30369,N_30018);
or U40325 (N_40325,N_31352,N_38225);
and U40326 (N_40326,N_32489,N_37542);
nor U40327 (N_40327,N_34703,N_36576);
or U40328 (N_40328,N_30593,N_32517);
and U40329 (N_40329,N_34670,N_34552);
nor U40330 (N_40330,N_35851,N_33650);
xnor U40331 (N_40331,N_32708,N_30578);
xor U40332 (N_40332,N_32589,N_33725);
and U40333 (N_40333,N_36385,N_34493);
nor U40334 (N_40334,N_34612,N_36988);
or U40335 (N_40335,N_39851,N_34599);
xnor U40336 (N_40336,N_38941,N_39497);
nand U40337 (N_40337,N_36108,N_30912);
and U40338 (N_40338,N_32417,N_38984);
and U40339 (N_40339,N_39271,N_38523);
xor U40340 (N_40340,N_31532,N_39623);
or U40341 (N_40341,N_38030,N_36638);
or U40342 (N_40342,N_33760,N_32014);
nand U40343 (N_40343,N_31982,N_35225);
nor U40344 (N_40344,N_37151,N_37415);
xor U40345 (N_40345,N_33928,N_36176);
nand U40346 (N_40346,N_36177,N_32462);
xnor U40347 (N_40347,N_37305,N_37798);
and U40348 (N_40348,N_34979,N_32801);
or U40349 (N_40349,N_37581,N_32968);
xnor U40350 (N_40350,N_35738,N_38195);
or U40351 (N_40351,N_32476,N_39488);
nand U40352 (N_40352,N_37764,N_36038);
xnor U40353 (N_40353,N_38687,N_34035);
nor U40354 (N_40354,N_31812,N_36381);
nor U40355 (N_40355,N_37858,N_37441);
xnor U40356 (N_40356,N_35256,N_37761);
xnor U40357 (N_40357,N_37732,N_37238);
or U40358 (N_40358,N_31440,N_37769);
or U40359 (N_40359,N_36262,N_32131);
and U40360 (N_40360,N_35905,N_39469);
and U40361 (N_40361,N_30076,N_35260);
nor U40362 (N_40362,N_33671,N_38209);
nor U40363 (N_40363,N_32697,N_31378);
xnor U40364 (N_40364,N_33175,N_31350);
nand U40365 (N_40365,N_33984,N_37304);
xor U40366 (N_40366,N_33802,N_31797);
and U40367 (N_40367,N_31385,N_36003);
nand U40368 (N_40368,N_36175,N_39002);
and U40369 (N_40369,N_38433,N_37286);
or U40370 (N_40370,N_38332,N_37019);
xnor U40371 (N_40371,N_34145,N_36056);
or U40372 (N_40372,N_30379,N_34638);
nor U40373 (N_40373,N_38546,N_36881);
nor U40374 (N_40374,N_30386,N_32454);
nand U40375 (N_40375,N_36523,N_31224);
xor U40376 (N_40376,N_30875,N_35139);
and U40377 (N_40377,N_39850,N_34773);
xnor U40378 (N_40378,N_31370,N_30755);
xnor U40379 (N_40379,N_39411,N_34639);
nor U40380 (N_40380,N_35760,N_33198);
nor U40381 (N_40381,N_31659,N_39819);
or U40382 (N_40382,N_38977,N_31933);
nand U40383 (N_40383,N_37241,N_36956);
nor U40384 (N_40384,N_36594,N_32668);
xor U40385 (N_40385,N_33805,N_30870);
and U40386 (N_40386,N_38725,N_31753);
and U40387 (N_40387,N_35045,N_32945);
xnor U40388 (N_40388,N_30732,N_38250);
nand U40389 (N_40389,N_36206,N_30655);
xnor U40390 (N_40390,N_31822,N_32375);
and U40391 (N_40391,N_34069,N_33604);
nand U40392 (N_40392,N_37200,N_32174);
and U40393 (N_40393,N_30042,N_39349);
nand U40394 (N_40394,N_31754,N_32515);
or U40395 (N_40395,N_33195,N_33787);
nand U40396 (N_40396,N_31436,N_33930);
and U40397 (N_40397,N_30452,N_36857);
xor U40398 (N_40398,N_38590,N_33843);
or U40399 (N_40399,N_35606,N_37789);
and U40400 (N_40400,N_30299,N_34964);
xnor U40401 (N_40401,N_37303,N_32558);
or U40402 (N_40402,N_38989,N_38813);
nor U40403 (N_40403,N_32315,N_34487);
or U40404 (N_40404,N_32448,N_31818);
xnor U40405 (N_40405,N_35007,N_34428);
or U40406 (N_40406,N_31678,N_35413);
and U40407 (N_40407,N_39269,N_36885);
nand U40408 (N_40408,N_30885,N_32686);
nand U40409 (N_40409,N_36686,N_31420);
nand U40410 (N_40410,N_37714,N_32092);
and U40411 (N_40411,N_38588,N_32362);
and U40412 (N_40412,N_39764,N_36667);
nor U40413 (N_40413,N_34623,N_34819);
and U40414 (N_40414,N_30722,N_35040);
xnor U40415 (N_40415,N_30952,N_31463);
xor U40416 (N_40416,N_34115,N_35497);
and U40417 (N_40417,N_31432,N_38899);
or U40418 (N_40418,N_39936,N_38128);
nand U40419 (N_40419,N_34368,N_39446);
nand U40420 (N_40420,N_39972,N_31037);
xor U40421 (N_40421,N_35802,N_38384);
or U40422 (N_40422,N_31376,N_38126);
nor U40423 (N_40423,N_32182,N_37747);
and U40424 (N_40424,N_37941,N_37917);
xor U40425 (N_40425,N_38418,N_36461);
or U40426 (N_40426,N_31153,N_35060);
nand U40427 (N_40427,N_39552,N_36101);
nand U40428 (N_40428,N_38634,N_39278);
nor U40429 (N_40429,N_31823,N_33516);
or U40430 (N_40430,N_31391,N_32862);
or U40431 (N_40431,N_35534,N_32432);
nand U40432 (N_40432,N_39615,N_36118);
nand U40433 (N_40433,N_39490,N_30381);
and U40434 (N_40434,N_39733,N_33564);
nor U40435 (N_40435,N_34354,N_36146);
nor U40436 (N_40436,N_38997,N_34725);
or U40437 (N_40437,N_37315,N_36473);
nor U40438 (N_40438,N_33710,N_38183);
xnor U40439 (N_40439,N_35615,N_37318);
nor U40440 (N_40440,N_31039,N_30432);
or U40441 (N_40441,N_31422,N_35243);
xor U40442 (N_40442,N_30711,N_38563);
xor U40443 (N_40443,N_30635,N_39513);
and U40444 (N_40444,N_34616,N_39449);
xor U40445 (N_40445,N_32104,N_34361);
xor U40446 (N_40446,N_33397,N_36607);
and U40447 (N_40447,N_34876,N_33829);
xor U40448 (N_40448,N_34212,N_38144);
nand U40449 (N_40449,N_37273,N_35848);
and U40450 (N_40450,N_33255,N_35537);
or U40451 (N_40451,N_33971,N_38094);
nor U40452 (N_40452,N_30368,N_37183);
nor U40453 (N_40453,N_32946,N_37096);
or U40454 (N_40454,N_33368,N_34512);
nand U40455 (N_40455,N_34433,N_33887);
nand U40456 (N_40456,N_35825,N_36595);
xnor U40457 (N_40457,N_38186,N_30922);
and U40458 (N_40458,N_36580,N_30089);
and U40459 (N_40459,N_33532,N_36812);
or U40460 (N_40460,N_33044,N_33227);
and U40461 (N_40461,N_37452,N_32381);
and U40462 (N_40462,N_39219,N_37353);
and U40463 (N_40463,N_35111,N_32537);
and U40464 (N_40464,N_38873,N_36522);
xnor U40465 (N_40465,N_38608,N_36807);
nand U40466 (N_40466,N_34481,N_30983);
nand U40467 (N_40467,N_34249,N_38441);
xnor U40468 (N_40468,N_37937,N_36972);
and U40469 (N_40469,N_34809,N_39712);
xnor U40470 (N_40470,N_35186,N_38555);
and U40471 (N_40471,N_32618,N_35303);
nor U40472 (N_40472,N_39233,N_33747);
and U40473 (N_40473,N_32998,N_38050);
and U40474 (N_40474,N_35996,N_35516);
nor U40475 (N_40475,N_35811,N_33819);
xor U40476 (N_40476,N_38335,N_34613);
or U40477 (N_40477,N_30537,N_37936);
nor U40478 (N_40478,N_33622,N_31538);
and U40479 (N_40479,N_32146,N_30156);
and U40480 (N_40480,N_35620,N_31963);
or U40481 (N_40481,N_35822,N_39403);
xor U40482 (N_40482,N_31355,N_33798);
or U40483 (N_40483,N_35875,N_30137);
nand U40484 (N_40484,N_33827,N_32765);
or U40485 (N_40485,N_37627,N_38012);
nand U40486 (N_40486,N_36128,N_31556);
or U40487 (N_40487,N_35292,N_39999);
nand U40488 (N_40488,N_36102,N_36293);
xnor U40489 (N_40489,N_35419,N_32798);
nand U40490 (N_40490,N_38680,N_35471);
xnor U40491 (N_40491,N_30323,N_34383);
nor U40492 (N_40492,N_34091,N_35860);
nand U40493 (N_40493,N_32437,N_39205);
and U40494 (N_40494,N_35664,N_38848);
and U40495 (N_40495,N_33750,N_37425);
nor U40496 (N_40496,N_34061,N_38174);
nor U40497 (N_40497,N_39933,N_31236);
or U40498 (N_40498,N_36770,N_37513);
nand U40499 (N_40499,N_32225,N_36229);
xor U40500 (N_40500,N_38436,N_35404);
nor U40501 (N_40501,N_37423,N_33653);
and U40502 (N_40502,N_37328,N_37003);
nand U40503 (N_40503,N_34569,N_39801);
nor U40504 (N_40504,N_38594,N_34730);
nand U40505 (N_40505,N_30033,N_38459);
nand U40506 (N_40506,N_39056,N_36558);
or U40507 (N_40507,N_36470,N_37488);
and U40508 (N_40508,N_36858,N_37307);
or U40509 (N_40509,N_38678,N_36552);
or U40510 (N_40510,N_39846,N_37430);
nand U40511 (N_40511,N_35242,N_39042);
nand U40512 (N_40512,N_34691,N_32077);
and U40513 (N_40513,N_31398,N_30072);
xor U40514 (N_40514,N_39162,N_33307);
nand U40515 (N_40515,N_33646,N_35590);
xnor U40516 (N_40516,N_36911,N_38581);
nor U40517 (N_40517,N_39494,N_38467);
and U40518 (N_40518,N_39916,N_31521);
nand U40519 (N_40519,N_32231,N_37793);
or U40520 (N_40520,N_32267,N_38326);
and U40521 (N_40521,N_35118,N_37965);
nand U40522 (N_40522,N_30385,N_33180);
and U40523 (N_40523,N_35204,N_30768);
and U40524 (N_40524,N_37296,N_36029);
nand U40525 (N_40525,N_35214,N_33959);
xnor U40526 (N_40526,N_31720,N_35602);
xor U40527 (N_40527,N_37987,N_32106);
nand U40528 (N_40528,N_30793,N_30456);
nand U40529 (N_40529,N_36776,N_39980);
nand U40530 (N_40530,N_31218,N_36297);
or U40531 (N_40531,N_35241,N_35610);
and U40532 (N_40532,N_34309,N_38814);
or U40533 (N_40533,N_34484,N_33919);
nor U40534 (N_40534,N_32983,N_38454);
and U40535 (N_40535,N_30233,N_33755);
or U40536 (N_40536,N_34777,N_33816);
xnor U40537 (N_40537,N_36427,N_36285);
xor U40538 (N_40538,N_37316,N_37925);
nor U40539 (N_40539,N_33464,N_36084);
and U40540 (N_40540,N_30474,N_31663);
nor U40541 (N_40541,N_38783,N_31779);
or U40542 (N_40542,N_37514,N_37825);
nand U40543 (N_40543,N_32172,N_32497);
xnor U40544 (N_40544,N_31113,N_33705);
nor U40545 (N_40545,N_32204,N_30371);
or U40546 (N_40546,N_36946,N_32505);
and U40547 (N_40547,N_35673,N_35016);
nor U40548 (N_40548,N_37639,N_30079);
xnor U40549 (N_40549,N_34621,N_37129);
nand U40550 (N_40550,N_36135,N_32694);
xor U40551 (N_40551,N_30675,N_38716);
nand U40552 (N_40552,N_32042,N_33883);
and U40553 (N_40553,N_35876,N_38606);
nand U40554 (N_40554,N_34513,N_31023);
xor U40555 (N_40555,N_31329,N_30208);
xor U40556 (N_40556,N_30694,N_38471);
nand U40557 (N_40557,N_39135,N_33200);
nor U40558 (N_40558,N_31989,N_35849);
nand U40559 (N_40559,N_38491,N_30021);
or U40560 (N_40560,N_36195,N_35991);
and U40561 (N_40561,N_35084,N_39664);
and U40562 (N_40562,N_34053,N_33149);
nor U40563 (N_40563,N_39152,N_35919);
nor U40564 (N_40564,N_35059,N_34357);
or U40565 (N_40565,N_38752,N_31332);
nand U40566 (N_40566,N_32898,N_36609);
or U40567 (N_40567,N_34565,N_39667);
xor U40568 (N_40568,N_30660,N_30180);
nand U40569 (N_40569,N_38920,N_31294);
xor U40570 (N_40570,N_33226,N_31722);
nor U40571 (N_40571,N_36401,N_31732);
and U40572 (N_40572,N_35714,N_30372);
xor U40573 (N_40573,N_30787,N_39676);
nor U40574 (N_40574,N_37615,N_30025);
or U40575 (N_40575,N_38693,N_33158);
and U40576 (N_40576,N_36921,N_31121);
and U40577 (N_40577,N_30396,N_39910);
xnor U40578 (N_40578,N_32812,N_35250);
nand U40579 (N_40579,N_31778,N_34811);
and U40580 (N_40580,N_37489,N_35423);
nor U40581 (N_40581,N_38232,N_39888);
nand U40582 (N_40582,N_36537,N_34798);
and U40583 (N_40583,N_37892,N_37240);
nor U40584 (N_40584,N_39295,N_36441);
xor U40585 (N_40585,N_30056,N_32126);
nand U40586 (N_40586,N_33312,N_38736);
and U40587 (N_40587,N_32623,N_38850);
nor U40588 (N_40588,N_35405,N_30282);
xnor U40589 (N_40589,N_34041,N_35385);
nand U40590 (N_40590,N_35512,N_38018);
and U40591 (N_40591,N_38522,N_32240);
and U40592 (N_40592,N_31773,N_36502);
xor U40593 (N_40593,N_39230,N_37811);
and U40594 (N_40594,N_37043,N_33462);
nand U40595 (N_40595,N_39895,N_37313);
nor U40596 (N_40596,N_31048,N_38858);
nand U40597 (N_40597,N_35530,N_37877);
or U40598 (N_40598,N_30374,N_30826);
or U40599 (N_40599,N_32224,N_34297);
xnor U40600 (N_40600,N_33061,N_34332);
nor U40601 (N_40601,N_37223,N_36104);
and U40602 (N_40602,N_34619,N_39080);
xnor U40603 (N_40603,N_36991,N_38602);
and U40604 (N_40604,N_31449,N_34066);
nand U40605 (N_40605,N_30211,N_38582);
nand U40606 (N_40606,N_36129,N_30909);
and U40607 (N_40607,N_33165,N_35427);
or U40608 (N_40608,N_36891,N_37845);
nor U40609 (N_40609,N_31445,N_30170);
and U40610 (N_40610,N_39831,N_39440);
or U40611 (N_40611,N_34410,N_30831);
xnor U40612 (N_40612,N_38517,N_38793);
and U40613 (N_40613,N_39803,N_39404);
or U40614 (N_40614,N_38872,N_35683);
nor U40615 (N_40615,N_36331,N_36396);
or U40616 (N_40616,N_38379,N_39642);
xnor U40617 (N_40617,N_31999,N_38368);
xor U40618 (N_40618,N_35430,N_33762);
xor U40619 (N_40619,N_39914,N_32203);
xnor U40620 (N_40620,N_33800,N_30407);
or U40621 (N_40621,N_31363,N_34273);
xor U40622 (N_40622,N_35278,N_36947);
or U40623 (N_40623,N_38342,N_38897);
nand U40624 (N_40624,N_39796,N_34420);
and U40625 (N_40625,N_32633,N_33445);
or U40626 (N_40626,N_37493,N_31608);
or U40627 (N_40627,N_38743,N_32804);
or U40628 (N_40628,N_36861,N_36364);
or U40629 (N_40629,N_30406,N_33018);
or U40630 (N_40630,N_35904,N_36618);
xnor U40631 (N_40631,N_34714,N_36288);
and U40632 (N_40632,N_36902,N_31955);
nand U40633 (N_40633,N_31132,N_32494);
xnor U40634 (N_40634,N_35467,N_38794);
xnor U40635 (N_40635,N_31145,N_39159);
xnor U40636 (N_40636,N_35305,N_30642);
nand U40637 (N_40637,N_32097,N_38688);
nor U40638 (N_40638,N_32284,N_38139);
nor U40639 (N_40639,N_34192,N_37537);
or U40640 (N_40640,N_32175,N_36725);
xor U40641 (N_40641,N_37589,N_38686);
nor U40642 (N_40642,N_31405,N_37219);
xnor U40643 (N_40643,N_38315,N_39147);
or U40644 (N_40644,N_37836,N_34002);
and U40645 (N_40645,N_36530,N_36905);
or U40646 (N_40646,N_30286,N_36106);
nand U40647 (N_40647,N_34677,N_38003);
nand U40648 (N_40648,N_37143,N_36308);
nand U40649 (N_40649,N_32367,N_35792);
xnor U40650 (N_40650,N_34399,N_30444);
xnor U40651 (N_40651,N_38511,N_36156);
nand U40652 (N_40652,N_39014,N_32248);
and U40653 (N_40653,N_31040,N_30362);
and U40654 (N_40654,N_33081,N_33669);
nor U40655 (N_40655,N_32654,N_33916);
nor U40656 (N_40656,N_31890,N_34530);
xnor U40657 (N_40657,N_37086,N_32900);
nor U40658 (N_40658,N_32559,N_37203);
or U40659 (N_40659,N_30492,N_31262);
xor U40660 (N_40660,N_35473,N_31509);
and U40661 (N_40661,N_31671,N_31860);
and U40662 (N_40662,N_37257,N_33021);
and U40663 (N_40663,N_36290,N_36727);
nor U40664 (N_40664,N_32196,N_36645);
or U40665 (N_40665,N_35684,N_35251);
xnor U40666 (N_40666,N_38492,N_31416);
xor U40667 (N_40667,N_33523,N_33495);
nor U40668 (N_40668,N_33583,N_33230);
and U40669 (N_40669,N_36843,N_34268);
and U40670 (N_40670,N_36097,N_39968);
xor U40671 (N_40671,N_31758,N_34298);
xor U40672 (N_40672,N_39032,N_37603);
xor U40673 (N_40673,N_33360,N_38189);
xor U40674 (N_40674,N_31086,N_35807);
or U40675 (N_40675,N_37750,N_39690);
nand U40676 (N_40676,N_37822,N_31634);
xor U40677 (N_40677,N_34666,N_33912);
and U40678 (N_40678,N_36322,N_38891);
nor U40679 (N_40679,N_37464,N_32150);
nand U40680 (N_40680,N_36382,N_33911);
nand U40681 (N_40681,N_30879,N_37482);
nand U40682 (N_40682,N_36388,N_31240);
or U40683 (N_40683,N_35483,N_39929);
and U40684 (N_40684,N_33977,N_31781);
xor U40685 (N_40685,N_38708,N_30941);
xnor U40686 (N_40686,N_38715,N_35572);
xnor U40687 (N_40687,N_38329,N_34977);
xor U40688 (N_40688,N_39711,N_33426);
or U40689 (N_40689,N_34058,N_32817);
and U40690 (N_40690,N_34645,N_30632);
nor U40691 (N_40691,N_35525,N_38938);
nor U40692 (N_40692,N_34585,N_38262);
or U40693 (N_40693,N_39518,N_30084);
or U40694 (N_40694,N_30330,N_35795);
and U40695 (N_40695,N_34889,N_32889);
nand U40696 (N_40696,N_35841,N_30161);
nor U40697 (N_40697,N_39707,N_36330);
nor U40698 (N_40698,N_35183,N_34391);
xor U40699 (N_40699,N_37710,N_35762);
nor U40700 (N_40700,N_37080,N_38904);
xnor U40701 (N_40701,N_32321,N_35761);
nand U40702 (N_40702,N_30907,N_39304);
nor U40703 (N_40703,N_32268,N_37054);
nand U40704 (N_40704,N_31110,N_36779);
xnor U40705 (N_40705,N_36240,N_38704);
or U40706 (N_40706,N_37442,N_36850);
nand U40707 (N_40707,N_31533,N_39436);
and U40708 (N_40708,N_30623,N_32145);
nand U40709 (N_40709,N_38973,N_39288);
nor U40710 (N_40710,N_34028,N_38440);
xnor U40711 (N_40711,N_34021,N_38870);
nand U40712 (N_40712,N_35307,N_35485);
nand U40713 (N_40713,N_38991,N_39723);
nor U40714 (N_40714,N_38346,N_32261);
and U40715 (N_40715,N_39268,N_34700);
and U40716 (N_40716,N_34735,N_36434);
xor U40717 (N_40717,N_39859,N_32745);
and U40718 (N_40718,N_33262,N_38506);
nor U40719 (N_40719,N_38957,N_30015);
or U40720 (N_40720,N_32960,N_39670);
or U40721 (N_40721,N_33535,N_34681);
xnor U40722 (N_40722,N_31270,N_31615);
nand U40723 (N_40723,N_35188,N_34788);
xor U40724 (N_40724,N_31633,N_35028);
or U40725 (N_40725,N_32709,N_30780);
or U40726 (N_40726,N_38916,N_32075);
nor U40727 (N_40727,N_35175,N_36662);
or U40728 (N_40728,N_32156,N_34079);
nor U40729 (N_40729,N_35581,N_33914);
nor U40730 (N_40730,N_32865,N_31120);
or U40731 (N_40731,N_33676,N_39261);
xnor U40732 (N_40732,N_34366,N_32897);
xnor U40733 (N_40733,N_30339,N_33038);
and U40734 (N_40734,N_36378,N_33196);
nor U40735 (N_40735,N_34760,N_34157);
and U40736 (N_40736,N_30895,N_31058);
or U40737 (N_40737,N_36785,N_33739);
xnor U40738 (N_40738,N_37352,N_38675);
nand U40739 (N_40739,N_32627,N_36751);
nand U40740 (N_40740,N_37235,N_39010);
xnor U40741 (N_40741,N_32008,N_31383);
and U40742 (N_40742,N_30220,N_32607);
or U40743 (N_40743,N_32933,N_30442);
and U40744 (N_40744,N_33734,N_30168);
nand U40745 (N_40745,N_30569,N_31193);
and U40746 (N_40746,N_34992,N_30792);
or U40747 (N_40747,N_36248,N_36701);
nand U40748 (N_40748,N_36734,N_31049);
nor U40749 (N_40749,N_36139,N_31435);
xnor U40750 (N_40750,N_35388,N_37896);
nand U40751 (N_40751,N_39187,N_36316);
nor U40752 (N_40752,N_39775,N_33970);
nand U40753 (N_40753,N_31924,N_35578);
nand U40754 (N_40754,N_39039,N_30968);
or U40755 (N_40755,N_30140,N_36245);
or U40756 (N_40756,N_33400,N_39371);
nand U40757 (N_40757,N_39104,N_35505);
xnor U40758 (N_40758,N_34215,N_31553);
xnor U40759 (N_40759,N_35715,N_39109);
and U40760 (N_40760,N_32395,N_38896);
and U40761 (N_40761,N_34881,N_36620);
and U40762 (N_40762,N_37028,N_38391);
or U40763 (N_40763,N_37862,N_32651);
xnor U40764 (N_40764,N_36680,N_34658);
nand U40765 (N_40765,N_30803,N_34930);
xor U40766 (N_40766,N_36318,N_31176);
xnor U40767 (N_40767,N_31163,N_33643);
or U40768 (N_40768,N_30783,N_37414);
or U40769 (N_40769,N_32543,N_30752);
nor U40770 (N_40770,N_33621,N_31554);
nand U40771 (N_40771,N_33933,N_35874);
and U40772 (N_40772,N_35074,N_32158);
or U40773 (N_40773,N_33003,N_31300);
and U40774 (N_40774,N_38035,N_35226);
or U40775 (N_40775,N_35727,N_38819);
xor U40776 (N_40776,N_39852,N_32028);
or U40777 (N_40777,N_39001,N_34749);
nor U40778 (N_40778,N_33893,N_31139);
nand U40779 (N_40779,N_33804,N_30828);
nand U40780 (N_40780,N_34514,N_31815);
nand U40781 (N_40781,N_30916,N_34832);
or U40782 (N_40782,N_35020,N_31555);
nor U40783 (N_40783,N_31131,N_39834);
or U40784 (N_40784,N_33620,N_37428);
nand U40785 (N_40785,N_36916,N_33988);
xnor U40786 (N_40786,N_31791,N_38874);
nor U40787 (N_40787,N_39313,N_32685);
xor U40788 (N_40788,N_30754,N_37245);
and U40789 (N_40789,N_31020,N_37014);
nand U40790 (N_40790,N_38475,N_34653);
nand U40791 (N_40791,N_34676,N_35426);
and U40792 (N_40792,N_30672,N_33095);
nand U40793 (N_40793,N_34454,N_32420);
or U40794 (N_40794,N_32347,N_34574);
xor U40795 (N_40795,N_31939,N_30292);
nor U40796 (N_40796,N_39781,N_38966);
xor U40797 (N_40797,N_36944,N_39948);
nor U40798 (N_40798,N_30397,N_32996);
or U40799 (N_40799,N_34921,N_37232);
or U40800 (N_40800,N_38767,N_38747);
or U40801 (N_40801,N_30011,N_30345);
nor U40802 (N_40802,N_37009,N_37735);
nand U40803 (N_40803,N_39847,N_31053);
nor U40804 (N_40804,N_30682,N_34027);
nand U40805 (N_40805,N_32953,N_32757);
and U40806 (N_40806,N_31609,N_37450);
nand U40807 (N_40807,N_37549,N_35132);
nand U40808 (N_40808,N_32047,N_32061);
and U40809 (N_40809,N_37373,N_38354);
and U40810 (N_40810,N_30940,N_37295);
nor U40811 (N_40811,N_39338,N_38109);
nand U40812 (N_40812,N_32500,N_33455);
nor U40813 (N_40813,N_37724,N_39514);
xor U40814 (N_40814,N_39060,N_38672);
and U40815 (N_40815,N_33473,N_37065);
or U40816 (N_40816,N_33963,N_37258);
xnor U40817 (N_40817,N_30852,N_35138);
xor U40818 (N_40818,N_38132,N_35043);
xor U40819 (N_40819,N_31212,N_37656);
nand U40820 (N_40820,N_31896,N_37282);
nand U40821 (N_40821,N_31395,N_37053);
and U40822 (N_40822,N_38472,N_32727);
nand U40823 (N_40823,N_31508,N_37351);
or U40824 (N_40824,N_38213,N_36081);
nand U40825 (N_40825,N_34699,N_39149);
nand U40826 (N_40826,N_32663,N_38371);
nor U40827 (N_40827,N_38773,N_33503);
xor U40828 (N_40828,N_32774,N_37640);
nand U40829 (N_40829,N_35156,N_39927);
or U40830 (N_40830,N_34688,N_35364);
xnor U40831 (N_40831,N_30716,N_39325);
xnor U40832 (N_40832,N_35554,N_34731);
or U40833 (N_40833,N_35609,N_32257);
or U40834 (N_40834,N_39757,N_37005);
nor U40835 (N_40835,N_32759,N_38072);
nor U40836 (N_40836,N_35567,N_34323);
nor U40837 (N_40837,N_33501,N_32966);
xor U40838 (N_40838,N_34683,N_35327);
or U40839 (N_40839,N_34918,N_32921);
and U40840 (N_40840,N_35648,N_31769);
nand U40841 (N_40841,N_31208,N_35444);
and U40842 (N_40842,N_31308,N_31761);
and U40843 (N_40843,N_34606,N_35299);
or U40844 (N_40844,N_33403,N_38053);
nand U40845 (N_40845,N_39028,N_37114);
and U40846 (N_40846,N_34563,N_33335);
or U40847 (N_40847,N_34342,N_31617);
nor U40848 (N_40848,N_37601,N_31495);
nand U40849 (N_40849,N_37991,N_33140);
and U40850 (N_40850,N_35363,N_31341);
xnor U40851 (N_40851,N_35154,N_38843);
nand U40852 (N_40852,N_38062,N_33906);
nor U40853 (N_40853,N_36815,N_32465);
nor U40854 (N_40854,N_34136,N_37742);
xnor U40855 (N_40855,N_36133,N_38754);
and U40856 (N_40856,N_37881,N_30517);
and U40857 (N_40857,N_35515,N_36452);
nor U40858 (N_40858,N_39279,N_35642);
and U40859 (N_40859,N_38415,N_31199);
xor U40860 (N_40860,N_38283,N_39157);
xnor U40861 (N_40861,N_34134,N_38212);
nand U40862 (N_40862,N_33995,N_30989);
nor U40863 (N_40863,N_38447,N_36016);
and U40864 (N_40864,N_32939,N_34595);
or U40865 (N_40865,N_38007,N_32002);
and U40866 (N_40866,N_36835,N_35233);
xnor U40867 (N_40867,N_35109,N_37456);
or U40868 (N_40868,N_37684,N_32385);
nor U40869 (N_40869,N_34990,N_34919);
xnor U40870 (N_40870,N_33996,N_37722);
nand U40871 (N_40871,N_39068,N_38671);
nand U40872 (N_40872,N_34006,N_32809);
or U40873 (N_40873,N_39254,N_38385);
nand U40874 (N_40874,N_34709,N_36661);
nand U40875 (N_40875,N_30876,N_30440);
and U40876 (N_40876,N_36043,N_34596);
or U40877 (N_40877,N_33774,N_31311);
xor U40878 (N_40878,N_34877,N_31653);
nor U40879 (N_40879,N_30401,N_37062);
nand U40880 (N_40880,N_39487,N_39397);
and U40881 (N_40881,N_39878,N_38880);
and U40882 (N_40882,N_32021,N_34640);
nand U40883 (N_40883,N_30643,N_39637);
and U40884 (N_40884,N_38311,N_35195);
nand U40885 (N_40885,N_32141,N_31424);
nand U40886 (N_40886,N_38365,N_36897);
and U40887 (N_40887,N_39958,N_33388);
nor U40888 (N_40888,N_34167,N_32931);
or U40889 (N_40889,N_34665,N_33771);
nor U40890 (N_40890,N_35071,N_39035);
xnor U40891 (N_40891,N_37582,N_31685);
and U40892 (N_40892,N_36405,N_39408);
or U40893 (N_40893,N_31080,N_35549);
or U40894 (N_40894,N_35746,N_39201);
nor U40895 (N_40895,N_38804,N_31805);
and U40896 (N_40896,N_32626,N_30351);
nor U40897 (N_40897,N_37672,N_34897);
xnor U40898 (N_40898,N_35754,N_32228);
xor U40899 (N_40899,N_35934,N_30625);
nand U40900 (N_40900,N_32036,N_37808);
nor U40901 (N_40901,N_37746,N_33063);
nor U40902 (N_40902,N_36920,N_34225);
xor U40903 (N_40903,N_36982,N_35966);
nand U40904 (N_40904,N_37576,N_33130);
xor U40905 (N_40905,N_31210,N_30427);
xnor U40906 (N_40906,N_30773,N_34003);
xor U40907 (N_40907,N_32886,N_34950);
or U40908 (N_40908,N_34151,N_31724);
nand U40909 (N_40909,N_39036,N_34885);
nand U40910 (N_40910,N_35026,N_33456);
or U40911 (N_40911,N_39299,N_32760);
nor U40912 (N_40912,N_38300,N_38493);
or U40913 (N_40913,N_38520,N_38692);
nor U40914 (N_40914,N_36343,N_37326);
nand U40915 (N_40915,N_34063,N_38982);
or U40916 (N_40916,N_34084,N_34893);
nand U40917 (N_40917,N_31531,N_37586);
nand U40918 (N_40918,N_36910,N_34684);
or U40919 (N_40919,N_38974,N_34100);
nor U40920 (N_40920,N_32445,N_34808);
or U40921 (N_40921,N_37588,N_38122);
and U40922 (N_40922,N_30175,N_39820);
xnor U40923 (N_40923,N_31052,N_38064);
nor U40924 (N_40924,N_32122,N_38495);
xnor U40925 (N_40925,N_30581,N_30844);
nand U40926 (N_40926,N_38239,N_32649);
nor U40927 (N_40927,N_38527,N_34951);
or U40928 (N_40928,N_33134,N_35270);
or U40929 (N_40929,N_32981,N_30866);
and U40930 (N_40930,N_34195,N_32466);
nand U40931 (N_40931,N_34659,N_38599);
xor U40932 (N_40932,N_30835,N_36145);
xor U40933 (N_40933,N_33688,N_33852);
nor U40934 (N_40934,N_35386,N_36863);
nand U40935 (N_40935,N_35318,N_30059);
nand U40936 (N_40936,N_38867,N_36304);
and U40937 (N_40937,N_35261,N_37418);
or U40938 (N_40938,N_31222,N_32070);
or U40939 (N_40939,N_31953,N_37367);
xnor U40940 (N_40940,N_30719,N_38294);
nor U40941 (N_40941,N_34187,N_30585);
or U40942 (N_40942,N_33777,N_33909);
nand U40943 (N_40943,N_30158,N_33253);
nand U40944 (N_40944,N_38292,N_38269);
nor U40945 (N_40945,N_34379,N_34865);
and U40946 (N_40946,N_37596,N_33191);
xor U40947 (N_40947,N_35335,N_32582);
and U40948 (N_40948,N_36821,N_30880);
nor U40949 (N_40949,N_34830,N_39466);
and U40950 (N_40950,N_37133,N_35940);
xnor U40951 (N_40951,N_36965,N_37851);
nor U40952 (N_40952,N_32726,N_33706);
and U40953 (N_40953,N_31642,N_37108);
and U40954 (N_40954,N_38259,N_34854);
and U40955 (N_40955,N_36057,N_38951);
and U40956 (N_40956,N_36173,N_35269);
nor U40957 (N_40957,N_33917,N_34016);
xnor U40958 (N_40958,N_34937,N_31987);
and U40959 (N_40959,N_33782,N_39681);
and U40960 (N_40960,N_37349,N_32777);
and U40961 (N_40961,N_35633,N_31015);
nor U40962 (N_40962,N_34159,N_39907);
nand U40963 (N_40963,N_34193,N_30480);
or U40964 (N_40964,N_39008,N_38758);
nand U40965 (N_40965,N_37743,N_36237);
nand U40966 (N_40966,N_33707,N_34204);
or U40967 (N_40967,N_34781,N_31124);
nand U40968 (N_40968,N_39320,N_39345);
or U40969 (N_40969,N_35375,N_36814);
nor U40970 (N_40970,N_33836,N_38583);
xnor U40971 (N_40971,N_36384,N_30342);
nor U40972 (N_40972,N_39248,N_39901);
nor U40973 (N_40973,N_34741,N_30595);
nand U40974 (N_40974,N_32331,N_38587);
and U40975 (N_40975,N_31973,N_37626);
nor U40976 (N_40976,N_35331,N_32118);
xnor U40977 (N_40977,N_37188,N_30889);
or U40978 (N_40978,N_36975,N_33453);
nand U40979 (N_40979,N_34649,N_32739);
nand U40980 (N_40980,N_36247,N_32620);
nand U40981 (N_40981,N_35675,N_37061);
xnor U40982 (N_40982,N_37723,N_36718);
or U40983 (N_40983,N_39204,N_37115);
nor U40984 (N_40984,N_38382,N_34008);
and U40985 (N_40985,N_38424,N_37810);
nor U40986 (N_40986,N_30520,N_37336);
and U40987 (N_40987,N_31594,N_35196);
nand U40988 (N_40988,N_33387,N_31768);
nor U40989 (N_40989,N_32344,N_33664);
xor U40990 (N_40990,N_34096,N_32394);
nor U40991 (N_40991,N_34722,N_32130);
nand U40992 (N_40992,N_30350,N_34584);
or U40993 (N_40993,N_37616,N_33960);
or U40994 (N_40994,N_33266,N_35157);
or U40995 (N_40995,N_38654,N_34780);
nor U40996 (N_40996,N_32155,N_33123);
and U40997 (N_40997,N_34230,N_37147);
or U40998 (N_40998,N_30225,N_37827);
nand U40999 (N_40999,N_39047,N_36504);
xor U41000 (N_41000,N_37727,N_39370);
and U41001 (N_41001,N_34243,N_30893);
xnor U41002 (N_41002,N_31180,N_39456);
and U41003 (N_41003,N_35123,N_32140);
and U41004 (N_41004,N_32229,N_39744);
nand U41005 (N_41005,N_34175,N_31873);
or U41006 (N_41006,N_35144,N_33736);
nand U41007 (N_41007,N_30109,N_31995);
xnor U41008 (N_41008,N_36179,N_38243);
xor U41009 (N_41009,N_34597,N_39046);
and U41010 (N_41010,N_35094,N_32081);
xnor U41011 (N_41011,N_39356,N_35351);
or U41012 (N_41012,N_36960,N_34888);
and U41013 (N_41013,N_37809,N_37760);
xor U41014 (N_41014,N_33629,N_34954);
nand U41015 (N_41015,N_33678,N_39125);
or U41016 (N_41016,N_38701,N_39309);
and U41017 (N_41017,N_36311,N_36619);
nor U41018 (N_41018,N_36410,N_38760);
or U41019 (N_41019,N_36406,N_32419);
nand U41020 (N_41020,N_36197,N_36468);
or U41021 (N_41021,N_32453,N_38430);
and U41022 (N_41022,N_38862,N_38683);
or U41023 (N_41023,N_32421,N_39875);
and U41024 (N_41024,N_39702,N_35218);
nand U41025 (N_41025,N_30806,N_34030);
or U41026 (N_41026,N_34086,N_37078);
nor U41027 (N_41027,N_30124,N_32656);
or U41028 (N_41028,N_30953,N_39116);
and U41029 (N_41029,N_30321,N_33176);
nor U41030 (N_41030,N_32835,N_31887);
nor U41031 (N_41031,N_39387,N_38287);
and U41032 (N_41032,N_30923,N_31412);
and U41033 (N_41033,N_32348,N_34406);
nand U41034 (N_41034,N_37981,N_36862);
xnor U41035 (N_41035,N_30847,N_38503);
and U41036 (N_41036,N_35990,N_30531);
nor U41037 (N_41037,N_34010,N_35119);
or U41038 (N_41038,N_36035,N_35277);
nand U41039 (N_41039,N_39990,N_39357);
nand U41040 (N_41040,N_36001,N_36225);
xnor U41041 (N_41041,N_32217,N_37852);
nand U41042 (N_41042,N_37134,N_36672);
nor U41043 (N_41043,N_37337,N_37125);
nand U41044 (N_41044,N_33152,N_36847);
xor U41045 (N_41045,N_38871,N_31974);
or U41046 (N_41046,N_34341,N_31794);
nand U41047 (N_41047,N_36574,N_31441);
xnor U41048 (N_41048,N_35095,N_33619);
nand U41049 (N_41049,N_39168,N_38333);
or U41050 (N_41050,N_38578,N_31179);
nand U41051 (N_41051,N_35692,N_39858);
or U41052 (N_41052,N_31889,N_35150);
or U41053 (N_41053,N_38673,N_35744);
nand U41054 (N_41054,N_37035,N_38130);
xnor U41055 (N_41055,N_30721,N_31447);
nand U41056 (N_41056,N_39545,N_38075);
and U41057 (N_41057,N_35629,N_39183);
nor U41058 (N_41058,N_37122,N_32890);
nand U41059 (N_41059,N_37655,N_38965);
nand U41060 (N_41060,N_37268,N_36124);
or U41061 (N_41061,N_32397,N_32382);
xor U41062 (N_41062,N_37469,N_35532);
and U41063 (N_41063,N_34000,N_30949);
nor U41064 (N_41064,N_34704,N_37157);
or U41065 (N_41065,N_33428,N_39114);
xor U41066 (N_41066,N_30570,N_33339);
nor U41067 (N_41067,N_35930,N_30670);
or U41068 (N_41068,N_31168,N_37380);
nand U41069 (N_41069,N_39903,N_35687);
nand U41070 (N_41070,N_32920,N_32750);
and U41071 (N_41071,N_37995,N_30431);
nand U41072 (N_41072,N_31843,N_35349);
nor U41073 (N_41073,N_33687,N_36610);
xnor U41074 (N_41074,N_34632,N_39374);
nand U41075 (N_41075,N_34737,N_37057);
nor U41076 (N_41076,N_36876,N_38633);
and U41077 (N_41077,N_37164,N_36739);
nor U41078 (N_41078,N_32879,N_34932);
nand U41079 (N_41079,N_32040,N_37641);
nor U41080 (N_41080,N_39142,N_35637);
xor U41081 (N_41081,N_32187,N_32201);
nand U41082 (N_41082,N_30577,N_33316);
nor U41083 (N_41083,N_33305,N_30888);
and U41084 (N_41084,N_32424,N_30120);
nand U41085 (N_41085,N_33124,N_35176);
and U41086 (N_41086,N_38785,N_30301);
or U41087 (N_41087,N_35401,N_30993);
xor U41088 (N_41088,N_31536,N_38074);
and U41089 (N_41089,N_34040,N_34316);
and U41090 (N_41090,N_39687,N_35420);
nand U41091 (N_41091,N_36398,N_39641);
nand U41092 (N_41092,N_33298,N_36797);
nor U41093 (N_41093,N_33261,N_31497);
or U41094 (N_41094,N_32718,N_32866);
xnor U41095 (N_41095,N_31410,N_34186);
xor U41096 (N_41096,N_37523,N_38458);
or U41097 (N_41097,N_39809,N_35038);
xor U41098 (N_41098,N_36743,N_38099);
or U41099 (N_41099,N_39407,N_39881);
or U41100 (N_41100,N_31907,N_35603);
and U41101 (N_41101,N_36278,N_38496);
nor U41102 (N_41102,N_34745,N_36268);
or U41103 (N_41103,N_31517,N_30248);
and U41104 (N_41104,N_34171,N_34324);
and U41105 (N_41105,N_30547,N_30882);
nor U41106 (N_41106,N_35691,N_34125);
and U41107 (N_41107,N_31074,N_39095);
or U41108 (N_41108,N_39312,N_39957);
xnor U41109 (N_41109,N_33025,N_34024);
nor U41110 (N_41110,N_37325,N_38317);
nand U41111 (N_41111,N_32734,N_35294);
and U41112 (N_41112,N_35671,N_33931);
and U41113 (N_41113,N_32134,N_31116);
xnor U41114 (N_41114,N_35387,N_30782);
or U41115 (N_41115,N_32082,N_30946);
nand U41116 (N_41116,N_36257,N_32511);
nor U41117 (N_41117,N_35376,N_33880);
or U41118 (N_41118,N_33673,N_37280);
or U41119 (N_41119,N_30428,N_39083);
xnor U41120 (N_41120,N_39952,N_33666);
nor U41121 (N_41121,N_38185,N_30041);
nor U41122 (N_41122,N_35667,N_39735);
nor U41123 (N_41123,N_36120,N_31804);
and U41124 (N_41124,N_39194,N_31806);
xnor U41125 (N_41125,N_36886,N_38784);
nor U41126 (N_41126,N_35236,N_35826);
and U41127 (N_41127,N_31275,N_34769);
xor U41128 (N_41128,N_36544,N_39608);
or U41129 (N_41129,N_31969,N_35644);
nor U41130 (N_41130,N_35005,N_39003);
or U41131 (N_41131,N_39376,N_34094);
or U41132 (N_41132,N_35935,N_36702);
or U41133 (N_41133,N_30053,N_31423);
nor U41134 (N_41134,N_39599,N_37231);
nor U41135 (N_41135,N_30533,N_38696);
nor U41136 (N_41136,N_35238,N_39574);
or U41137 (N_41137,N_31909,N_31714);
nor U41138 (N_41138,N_33527,N_32144);
or U41139 (N_41139,N_30316,N_31838);
nand U41140 (N_41140,N_32251,N_33835);
nor U41141 (N_41141,N_31322,N_31611);
or U41142 (N_41142,N_37984,N_32363);
nor U41143 (N_41143,N_31507,N_32086);
nor U41144 (N_41144,N_32792,N_31102);
and U41145 (N_41145,N_31365,N_33487);
nor U41146 (N_41146,N_31390,N_33187);
nor U41147 (N_41147,N_32279,N_36737);
xor U41148 (N_41148,N_33806,N_30253);
nor U41149 (N_41149,N_33578,N_31160);
xnor U41150 (N_41150,N_34320,N_31786);
xnor U41151 (N_41151,N_39004,N_37199);
or U41152 (N_41152,N_30159,N_30726);
xor U41153 (N_41153,N_31936,N_33737);
nand U41154 (N_41154,N_31635,N_36426);
nand U41155 (N_41155,N_31837,N_38264);
nand U41156 (N_41156,N_33202,N_33315);
nand U41157 (N_41157,N_30047,N_37686);
or U41158 (N_41158,N_30978,N_36437);
nor U41159 (N_41159,N_30781,N_32524);
or U41160 (N_41160,N_37580,N_38412);
xor U41161 (N_41161,N_32183,N_33746);
and U41162 (N_41162,N_33317,N_37267);
or U41163 (N_41163,N_39611,N_32899);
and U41164 (N_41164,N_38227,N_33251);
nor U41165 (N_41165,N_32924,N_36899);
nor U41166 (N_41166,N_35145,N_35129);
nor U41167 (N_41167,N_38224,N_35415);
xor U41168 (N_41168,N_35605,N_39937);
nand U41169 (N_41169,N_30945,N_36940);
xnor U41170 (N_41170,N_31188,N_37229);
nand U41171 (N_41171,N_34282,N_32304);
and U41172 (N_41172,N_37176,N_39912);
nand U41173 (N_41173,N_39055,N_39347);
and U41174 (N_41174,N_37455,N_37620);
nand U41175 (N_41175,N_31127,N_30160);
and U41176 (N_41176,N_39249,N_37649);
xnor U41177 (N_41177,N_34042,N_34211);
nor U41178 (N_41178,N_36466,N_30060);
or U41179 (N_41179,N_32746,N_39420);
nand U41180 (N_41180,N_36641,N_32551);
or U41181 (N_41181,N_38341,N_37668);
or U41182 (N_41182,N_32881,N_32301);
nor U41183 (N_41183,N_30975,N_31387);
nor U41184 (N_41184,N_37988,N_37622);
nand U41185 (N_41185,N_31811,N_39662);
and U41186 (N_41186,N_38642,N_37839);
or U41187 (N_41187,N_39836,N_38187);
nor U41188 (N_41188,N_36037,N_31918);
nor U41189 (N_41189,N_30213,N_33100);
and U41190 (N_41190,N_34912,N_31287);
xor U41191 (N_41191,N_38795,N_31119);
nand U41192 (N_41192,N_35468,N_38349);
and U41193 (N_41193,N_35121,N_36669);
or U41194 (N_41194,N_34339,N_37478);
and U41195 (N_41195,N_30731,N_38319);
nor U41196 (N_41196,N_32103,N_36286);
nor U41197 (N_41197,N_30238,N_33975);
and U41198 (N_41198,N_39018,N_37017);
xor U41199 (N_41199,N_32180,N_36987);
nand U41200 (N_41200,N_30129,N_34748);
nand U41201 (N_41201,N_35063,N_38923);
xnor U41202 (N_41202,N_39303,N_32022);
or U41203 (N_41203,N_36184,N_34432);
nor U41204 (N_41204,N_32471,N_31269);
nor U41205 (N_41205,N_31979,N_36819);
nor U41206 (N_41206,N_34356,N_31418);
or U41207 (N_41207,N_34669,N_37826);
xor U41208 (N_41208,N_37401,N_35539);
nand U41209 (N_41209,N_36178,N_33069);
nor U41210 (N_41210,N_34517,N_31225);
nor U41211 (N_41211,N_35142,N_33670);
nor U41212 (N_41212,N_32190,N_36358);
or U41213 (N_41213,N_35203,N_36579);
and U41214 (N_41214,N_39005,N_36306);
nor U41215 (N_41215,N_35293,N_32836);
or U41216 (N_41216,N_36624,N_38297);
and U41217 (N_41217,N_33498,N_32460);
nand U41218 (N_41218,N_38856,N_30437);
nor U41219 (N_41219,N_35290,N_36071);
nand U41220 (N_41220,N_30827,N_34833);
or U41221 (N_41221,N_31154,N_36313);
nand U41222 (N_41222,N_33273,N_39740);
or U41223 (N_41223,N_36224,N_37270);
nand U41224 (N_41224,N_34172,N_34052);
or U41225 (N_41225,N_38735,N_30209);
xnor U41226 (N_41226,N_32354,N_39953);
nand U41227 (N_41227,N_38907,N_31402);
xor U41228 (N_41228,N_31727,N_30647);
xor U41229 (N_41229,N_37000,N_32318);
nand U41230 (N_41230,N_32659,N_36511);
xnor U41231 (N_41231,N_35252,N_37868);
and U41232 (N_41232,N_30926,N_34858);
and U41233 (N_41233,N_33731,N_31282);
xnor U41234 (N_41234,N_33655,N_33005);
xnor U41235 (N_41235,N_32833,N_36232);
xnor U41236 (N_41236,N_38994,N_37277);
nor U41237 (N_41237,N_37645,N_35948);
nor U41238 (N_41238,N_30516,N_32396);
and U41239 (N_41239,N_33882,N_33035);
or U41240 (N_41240,N_31871,N_35333);
nor U41241 (N_41241,N_32379,N_37494);
nand U41242 (N_41242,N_38609,N_33558);
nor U41243 (N_41243,N_34600,N_34543);
or U41244 (N_41244,N_36186,N_33872);
or U41245 (N_41245,N_39917,N_31216);
or U41246 (N_41246,N_34031,N_30813);
or U41247 (N_41247,N_35611,N_30098);
and U41248 (N_41248,N_30504,N_36844);
nand U41249 (N_41249,N_31149,N_35308);
nor U41250 (N_41250,N_33064,N_37160);
or U41251 (N_41251,N_35908,N_35222);
nand U41252 (N_41252,N_38398,N_32053);
nand U41253 (N_41253,N_31340,N_33757);
nand U41254 (N_41254,N_39464,N_35076);
and U41255 (N_41255,N_33054,N_32868);
nor U41256 (N_41256,N_36143,N_34696);
nand U41257 (N_41257,N_37720,N_31158);
xor U41258 (N_41258,N_39353,N_30505);
and U41259 (N_41259,N_36979,N_37184);
nor U41260 (N_41260,N_32915,N_30356);
nand U41261 (N_41261,N_30065,N_36165);
and U41262 (N_41262,N_35640,N_32193);
nor U41263 (N_41263,N_31841,N_30877);
xor U41264 (N_41264,N_37602,N_30106);
and U41265 (N_41265,N_32262,N_36205);
nor U41266 (N_41266,N_31783,N_32883);
and U41267 (N_41267,N_36103,N_30583);
nand U41268 (N_41268,N_38271,N_32372);
and U41269 (N_41269,N_37331,N_37234);
nand U41270 (N_41270,N_36772,N_36731);
nand U41271 (N_41271,N_37661,N_34005);
nor U41272 (N_41272,N_37186,N_33998);
nand U41273 (N_41273,N_36409,N_38828);
and U41274 (N_41274,N_30166,N_35034);
nor U41275 (N_41275,N_38810,N_39922);
or U41276 (N_41276,N_39048,N_34138);
xor U41277 (N_41277,N_34820,N_38131);
or U41278 (N_41278,N_39199,N_32776);
and U41279 (N_41279,N_37486,N_37105);
or U41280 (N_41280,N_31134,N_33471);
xor U41281 (N_41281,N_38805,N_33492);
xnor U41282 (N_41282,N_30933,N_38059);
or U41283 (N_41283,N_39037,N_37390);
and U41284 (N_41284,N_37828,N_33560);
xnor U41285 (N_41285,N_31613,N_33659);
nor U41286 (N_41286,N_38676,N_33433);
xnor U41287 (N_41287,N_34804,N_36199);
and U41288 (N_41288,N_30536,N_32737);
nor U41289 (N_41289,N_39923,N_38939);
nor U41290 (N_41290,N_31988,N_30255);
nor U41291 (N_41291,N_36282,N_32907);
xnor U41292 (N_41292,N_36705,N_30744);
nand U41293 (N_41293,N_38895,N_39945);
nand U41294 (N_41294,N_36207,N_37567);
nand U41295 (N_41295,N_39989,N_37956);
or U41296 (N_41296,N_31099,N_37895);
nor U41297 (N_41297,N_35669,N_30740);
nor U41298 (N_41298,N_34185,N_39943);
nor U41299 (N_41299,N_38181,N_34459);
xor U41300 (N_41300,N_35463,N_34445);
xor U41301 (N_41301,N_30503,N_30256);
or U41302 (N_41302,N_36215,N_36668);
xnor U41303 (N_41303,N_34121,N_36892);
xor U41304 (N_41304,N_35281,N_37874);
and U41305 (N_41305,N_39703,N_33551);
or U41306 (N_41306,N_38104,N_35689);
xnor U41307 (N_41307,N_32539,N_31093);
or U41308 (N_41308,N_36719,N_38145);
xor U41309 (N_41309,N_36780,N_34983);
and U41310 (N_41310,N_31094,N_35945);
nor U41311 (N_41311,N_35509,N_36048);
nor U41312 (N_41312,N_34689,N_34706);
and U41313 (N_41313,N_30384,N_36688);
nor U41314 (N_41314,N_30090,N_35450);
nand U41315 (N_41315,N_39550,N_31431);
and U41316 (N_41316,N_32903,N_34625);
xor U41317 (N_41317,N_39427,N_38597);
xnor U41318 (N_41318,N_31091,N_36818);
and U41319 (N_41319,N_36493,N_31438);
nand U41320 (N_41320,N_34318,N_31226);
nor U41321 (N_41321,N_37831,N_32679);
and U41322 (N_41322,N_36073,N_30651);
xor U41323 (N_41323,N_36629,N_32010);
or U41324 (N_41324,N_39600,N_32220);
nor U41325 (N_41325,N_32311,N_37614);
or U41326 (N_41326,N_34515,N_32857);
or U41327 (N_41327,N_30728,N_38797);
nor U41328 (N_41328,N_36099,N_39181);
nand U41329 (N_41329,N_30606,N_32423);
and U41330 (N_41330,N_35801,N_36570);
nand U41331 (N_41331,N_33042,N_30734);
xnor U41332 (N_41332,N_32109,N_37396);
nor U41333 (N_41333,N_35445,N_38930);
or U41334 (N_41334,N_31621,N_32431);
and U41335 (N_41335,N_31031,N_32018);
or U41336 (N_41336,N_37505,N_39825);
nor U41337 (N_41337,N_33855,N_36435);
xnor U41338 (N_41338,N_36582,N_34518);
and U41339 (N_41339,N_34789,N_30906);
or U41340 (N_41340,N_34262,N_39027);
and U41341 (N_41341,N_30434,N_30467);
nand U41342 (N_41342,N_33031,N_39567);
and U41343 (N_41343,N_32611,N_38877);
and U41344 (N_41344,N_38627,N_31239);
or U41345 (N_41345,N_37967,N_33857);
or U41346 (N_41346,N_33717,N_34349);
nand U41347 (N_41347,N_34286,N_36294);
xnor U41348 (N_41348,N_38800,N_31959);
xnor U41349 (N_41349,N_31900,N_32356);
nor U41350 (N_41350,N_30069,N_39067);
or U41351 (N_41351,N_36307,N_34794);
or U41352 (N_41352,N_32937,N_34419);
xor U41353 (N_41353,N_33509,N_34707);
xor U41354 (N_41354,N_37659,N_33401);
xnor U41355 (N_41355,N_36211,N_36317);
xnor U41356 (N_41356,N_34784,N_31235);
nor U41357 (N_41357,N_35296,N_35732);
nand U41358 (N_41358,N_36280,N_31638);
nand U41359 (N_41359,N_30294,N_37421);
nand U41360 (N_41360,N_31802,N_30260);
nand U41361 (N_41361,N_30839,N_37985);
xnor U41362 (N_41362,N_33580,N_35448);
xor U41363 (N_41363,N_31709,N_33087);
xor U41364 (N_41364,N_32711,N_32822);
and U41365 (N_41365,N_32705,N_37497);
and U41366 (N_41366,N_33788,N_31298);
nor U41367 (N_41367,N_37243,N_37529);
xor U41368 (N_41368,N_33232,N_33677);
nand U41369 (N_41369,N_34166,N_39626);
and U41370 (N_41370,N_33460,N_32554);
and U41371 (N_41371,N_32255,N_38845);
nor U41372 (N_41372,N_36497,N_30295);
nand U41373 (N_41373,N_37990,N_39900);
and U41374 (N_41374,N_32410,N_35550);
nand U41375 (N_41375,N_38591,N_31381);
xor U41376 (N_41376,N_35168,N_34150);
nand U41377 (N_41377,N_34474,N_38684);
nand U41378 (N_41378,N_39732,N_36433);
or U41379 (N_41379,N_39169,N_35049);
or U41380 (N_41380,N_30114,N_37948);
or U41381 (N_41381,N_34989,N_37136);
or U41382 (N_41382,N_34587,N_35612);
or U41383 (N_41383,N_31114,N_38058);
nand U41384 (N_41384,N_39701,N_30174);
xnor U41385 (N_41385,N_32599,N_39133);
or U41386 (N_41386,N_31510,N_38639);
xor U41387 (N_41387,N_34261,N_35619);
and U41388 (N_41388,N_32206,N_34796);
and U41389 (N_41389,N_30343,N_36281);
and U41390 (N_41390,N_33414,N_37149);
and U41391 (N_41391,N_31035,N_38351);
and U41392 (N_41392,N_33174,N_33332);
xor U41393 (N_41393,N_35937,N_38276);
and U41394 (N_41394,N_36046,N_38727);
nor U41395 (N_41395,N_31874,N_38223);
nor U41396 (N_41396,N_36550,N_36879);
or U41397 (N_41397,N_38586,N_37555);
nand U41398 (N_41398,N_38049,N_32060);
or U41399 (N_41399,N_35235,N_36860);
or U41400 (N_41400,N_32457,N_30157);
nand U41401 (N_41401,N_37225,N_38595);
or U41402 (N_41402,N_33926,N_34213);
xor U41403 (N_41403,N_35127,N_30426);
xnor U41404 (N_41404,N_35149,N_39192);
nor U41405 (N_41405,N_36796,N_36336);
or U41406 (N_41406,N_37757,N_33765);
and U41407 (N_41407,N_34756,N_34852);
or U41408 (N_41408,N_33358,N_38726);
or U41409 (N_41409,N_34935,N_38318);
xor U41410 (N_41410,N_37144,N_34545);
xor U41411 (N_41411,N_39659,N_33790);
or U41412 (N_41412,N_36977,N_37364);
or U41413 (N_41413,N_34389,N_33588);
or U41414 (N_41414,N_37777,N_33045);
and U41415 (N_41415,N_35163,N_32033);
and U41416 (N_41416,N_33030,N_33631);
nor U41417 (N_41417,N_35117,N_33966);
xnor U41418 (N_41418,N_30100,N_34074);
xor U41419 (N_41419,N_31809,N_35255);
nand U41420 (N_41420,N_32849,N_36353);
xor U41421 (N_41421,N_33699,N_37568);
or U41422 (N_41422,N_32290,N_34610);
or U41423 (N_41423,N_32212,N_33184);
xnor U41424 (N_41424,N_36039,N_30811);
nor U41425 (N_41425,N_36069,N_38665);
nand U41426 (N_41426,N_35938,N_33886);
nand U41427 (N_41427,N_31169,N_36208);
nand U41428 (N_41428,N_36791,N_36925);
nor U41429 (N_41429,N_38494,N_39395);
and U41430 (N_41430,N_34553,N_36429);
nor U41431 (N_41431,N_39076,N_38394);
nor U41432 (N_41432,N_35091,N_31142);
nor U41433 (N_41433,N_31751,N_37463);
xor U41434 (N_41434,N_31782,N_38051);
and U41435 (N_41435,N_36367,N_38501);
nand U41436 (N_41436,N_30769,N_36707);
nand U41437 (N_41437,N_37251,N_33119);
and U41438 (N_41438,N_35482,N_39709);
nor U41439 (N_41439,N_32604,N_36214);
or U41440 (N_41440,N_31689,N_37692);
or U41441 (N_41441,N_38031,N_36521);
nor U41442 (N_41442,N_38863,N_33037);
xor U41443 (N_41443,N_30030,N_30964);
nor U41444 (N_41444,N_35545,N_37104);
nand U41445 (N_41445,N_39166,N_33566);
and U41446 (N_41446,N_32324,N_35481);
nor U41447 (N_41447,N_35396,N_30424);
or U41448 (N_41448,N_33961,N_36721);
xnor U41449 (N_41449,N_37730,N_35209);
xnor U41450 (N_41450,N_39594,N_31388);
nor U41451 (N_41451,N_37946,N_31831);
or U41452 (N_41452,N_37420,N_35041);
or U41453 (N_41453,N_37044,N_37427);
and U41454 (N_41454,N_34827,N_37553);
and U41455 (N_41455,N_38241,N_35081);
or U41456 (N_41456,N_36908,N_33656);
nand U41457 (N_41457,N_31629,N_30858);
xnor U41458 (N_41458,N_30693,N_36223);
and U41459 (N_41459,N_32984,N_31303);
xnor U41460 (N_41460,N_39996,N_32648);
nor U41461 (N_41461,N_33552,N_30990);
xor U41462 (N_41462,N_30074,N_36708);
xor U41463 (N_41463,N_38034,N_30997);
and U41464 (N_41464,N_32317,N_33744);
nor U41465 (N_41465,N_36567,N_38060);
nor U41466 (N_41466,N_38150,N_37275);
or U41467 (N_41467,N_38006,N_32287);
nor U41468 (N_41468,N_32510,N_39582);
nand U41469 (N_41469,N_35519,N_39789);
or U41470 (N_41470,N_39084,N_31111);
or U41471 (N_41471,N_34381,N_34516);
and U41472 (N_41472,N_38404,N_32752);
nand U41473 (N_41473,N_35389,N_38924);
nand U41474 (N_41474,N_37914,N_39242);
and U41475 (N_41475,N_35210,N_39829);
and U41476 (N_41476,N_35570,N_35984);
nand U41477 (N_41477,N_36447,N_34064);
or U41478 (N_41478,N_30967,N_34770);
nand U41479 (N_41479,N_33826,N_31106);
or U41480 (N_41480,N_38434,N_37983);
and U41481 (N_41481,N_32605,N_39341);
nand U41482 (N_41482,N_38955,N_37957);
or U41483 (N_41483,N_30496,N_36758);
nand U41484 (N_41484,N_38437,N_34751);
xnor U41485 (N_41485,N_31241,N_32073);
xnor U41486 (N_41486,N_31000,N_34686);
nor U41487 (N_41487,N_31316,N_30837);
or U41488 (N_41488,N_39237,N_38906);
and U41489 (N_41489,N_32434,N_30854);
nand U41490 (N_41490,N_34559,N_30324);
and U41491 (N_41491,N_38993,N_36997);
or U41492 (N_41492,N_39643,N_32975);
nand U41493 (N_41493,N_30917,N_31687);
xor U41494 (N_41494,N_35859,N_39554);
nor U41495 (N_41495,N_35369,N_37037);
xor U41496 (N_41496,N_33322,N_36485);
nor U41497 (N_41497,N_36230,N_37215);
xor U41498 (N_41498,N_30818,N_30662);
nor U41499 (N_41499,N_30699,N_39380);
xnor U41500 (N_41500,N_39902,N_30057);
nand U41501 (N_41501,N_39521,N_31657);
nor U41502 (N_41502,N_32567,N_30484);
or U41503 (N_41503,N_37454,N_36115);
or U41504 (N_41504,N_30197,N_31257);
nor U41505 (N_41505,N_39297,N_33638);
and U41506 (N_41506,N_39492,N_38547);
nor U41507 (N_41507,N_37535,N_32035);
nor U41508 (N_41508,N_38310,N_31348);
and U41509 (N_41509,N_39782,N_36872);
nor U41510 (N_41510,N_36439,N_33326);
nand U41511 (N_41511,N_34558,N_39429);
xor U41512 (N_41512,N_39118,N_36299);
xor U41513 (N_41513,N_31243,N_31735);
or U41514 (N_41514,N_31926,N_34156);
or U41515 (N_41515,N_38201,N_35722);
xnor U41516 (N_41516,N_38231,N_33531);
nand U41517 (N_41517,N_38288,N_33962);
xnor U41518 (N_41518,N_33470,N_36853);
and U41519 (N_41519,N_31704,N_38387);
nor U41520 (N_41520,N_33173,N_33181);
and U41521 (N_41521,N_39507,N_36492);
xor U41522 (N_41522,N_35584,N_31515);
nor U41523 (N_41523,N_30900,N_33529);
and U41524 (N_41524,N_38528,N_30627);
nor U41525 (N_41525,N_34435,N_36602);
xor U41526 (N_41526,N_35518,N_38662);
and U41527 (N_41527,N_36999,N_32436);
or U41528 (N_41528,N_33562,N_30601);
and U41529 (N_41529,N_37498,N_37515);
xor U41530 (N_41530,N_36869,N_36811);
nor U41531 (N_41531,N_33336,N_35312);
nand U41532 (N_41532,N_37702,N_39172);
nand U41533 (N_41533,N_35372,N_36076);
or U41534 (N_41534,N_30760,N_30528);
nand U41535 (N_41535,N_35165,N_35263);
xor U41536 (N_41536,N_38776,N_34365);
or U41537 (N_41537,N_30749,N_39583);
xor U41538 (N_41538,N_35164,N_32590);
and U41539 (N_41539,N_37342,N_39899);
xor U41540 (N_41540,N_38129,N_34523);
and U41541 (N_41541,N_35075,N_31073);
nor U41542 (N_41542,N_30152,N_36494);
nand U41543 (N_41543,N_31644,N_37124);
xnor U41544 (N_41544,N_35211,N_30820);
nand U41545 (N_41545,N_32577,N_39678);
nor U41546 (N_41546,N_33695,N_36121);
nand U41547 (N_41547,N_39280,N_37871);
and U41548 (N_41548,N_34085,N_30944);
nor U41549 (N_41549,N_33665,N_39111);
nand U41550 (N_41550,N_35416,N_36744);
nor U41551 (N_41551,N_33794,N_35230);
nand U41552 (N_41552,N_35985,N_38151);
nand U41553 (N_41553,N_31895,N_38668);
or U41554 (N_41554,N_31789,N_36393);
and U41555 (N_41555,N_38047,N_30142);
or U41556 (N_41556,N_32514,N_34968);
nand U41557 (N_41557,N_32179,N_36746);
nor U41558 (N_41558,N_36394,N_38568);
and U41559 (N_41559,N_39414,N_35929);
nor U41560 (N_41560,N_33939,N_30358);
xnor U41561 (N_41561,N_32278,N_39274);
nor U41562 (N_41562,N_31213,N_31878);
and U41563 (N_41563,N_30048,N_35208);
nand U41564 (N_41564,N_36374,N_37127);
or U41565 (N_41565,N_31366,N_31742);
nand U41566 (N_41566,N_35495,N_31723);
nand U41567 (N_41567,N_32164,N_33136);
xor U41568 (N_41568,N_34535,N_33754);
or U41569 (N_41569,N_33614,N_39434);
nand U41570 (N_41570,N_32684,N_32389);
or U41571 (N_41571,N_39281,N_39616);
and U41572 (N_41572,N_38807,N_37861);
nor U41573 (N_41573,N_35048,N_36877);
nand U41574 (N_41574,N_32219,N_38111);
nand U41575 (N_41575,N_36875,N_39719);
nor U41576 (N_41576,N_34288,N_38397);
or U41577 (N_41577,N_30250,N_37559);
xor U41578 (N_41578,N_39134,N_39119);
nand U41579 (N_41579,N_32547,N_39470);
xnor U41580 (N_41580,N_39959,N_31317);
or U41581 (N_41581,N_31957,N_34953);
nor U41582 (N_41582,N_34763,N_34430);
nor U41583 (N_41583,N_36303,N_34894);
nor U41584 (N_41584,N_30483,N_32549);
xor U41585 (N_41585,N_31103,N_38868);
nand U41586 (N_41586,N_31931,N_38569);
and U41587 (N_41587,N_34088,N_34657);
xnor U41588 (N_41588,N_39636,N_39649);
or U41589 (N_41589,N_34527,N_37632);
or U41590 (N_41590,N_33965,N_33884);
nand U41591 (N_41591,N_30738,N_36086);
nor U41592 (N_41592,N_38647,N_33398);
or U41593 (N_41593,N_36569,N_36557);
nor U41594 (N_41594,N_39986,N_30753);
nor U41595 (N_41595,N_35910,N_37971);
nand U41596 (N_41596,N_33818,N_38008);
xnor U41597 (N_41597,N_33001,N_34650);
and U41598 (N_41598,N_33382,N_39761);
or U41599 (N_41599,N_33896,N_32305);
and U41600 (N_41600,N_32873,N_35069);
and U41601 (N_41601,N_35000,N_39071);
or U41602 (N_41602,N_30064,N_39426);
and U41603 (N_41603,N_31276,N_30308);
nand U41604 (N_41604,N_36325,N_37708);
nor U41605 (N_41605,N_33177,N_37804);
or U41606 (N_41606,N_39337,N_38557);
nand U41607 (N_41607,N_32446,N_32658);
nor U41608 (N_41608,N_36747,N_35656);
xor U41609 (N_41609,N_31417,N_39246);
nand U41610 (N_41610,N_36851,N_35528);
and U41611 (N_41611,N_31442,N_39252);
xnor U41612 (N_41612,N_32038,N_32078);
nand U41613 (N_41613,N_31428,N_37379);
xnor U41614 (N_41614,N_36203,N_37973);
and U41615 (N_41615,N_39572,N_33541);
or U41616 (N_41616,N_30388,N_39024);
nand U41617 (N_41617,N_34358,N_33443);
nor U41618 (N_41618,N_33446,N_39276);
or U41619 (N_41619,N_37403,N_33987);
xor U41620 (N_41620,N_34844,N_31283);
nand U41621 (N_41621,N_31092,N_35693);
nor U41622 (N_41622,N_35046,N_33416);
nand U41623 (N_41623,N_34442,N_39301);
xnor U41624 (N_41624,N_35989,N_31299);
or U41625 (N_41625,N_39607,N_30807);
nand U41626 (N_41626,N_39603,N_33280);
or U41627 (N_41627,N_37958,N_35756);
nand U41628 (N_41628,N_30116,N_35979);
nand U41629 (N_41629,N_39000,N_39919);
or U41630 (N_41630,N_30049,N_35594);
xnor U41631 (N_41631,N_35742,N_33768);
nor U41632 (N_41632,N_33311,N_35442);
or U41633 (N_41633,N_36421,N_37736);
nor U41634 (N_41634,N_34179,N_39644);
or U41635 (N_41635,N_33974,N_30347);
nand U41636 (N_41636,N_30534,N_30802);
or U41637 (N_41637,N_32501,N_37069);
nand U41638 (N_41638,N_31607,N_30215);
or U41639 (N_41639,N_35339,N_31135);
or U41640 (N_41640,N_32252,N_35745);
xor U41641 (N_41641,N_38140,N_31750);
or U41642 (N_41642,N_36568,N_30915);
or U41643 (N_41643,N_35490,N_31993);
or U41644 (N_41644,N_36227,N_39096);
nand U41645 (N_41645,N_30190,N_32368);
xor U41646 (N_41646,N_34814,N_37419);
and U41647 (N_41647,N_34208,N_35104);
nor U41648 (N_41648,N_37908,N_37406);
nand U41649 (N_41649,N_35643,N_38014);
nand U41650 (N_41650,N_32581,N_31845);
or U41651 (N_41651,N_32198,N_35130);
or U41652 (N_41652,N_33002,N_36415);
and U41653 (N_41653,N_31479,N_37332);
or U41654 (N_41654,N_36321,N_32281);
and U41655 (N_41655,N_35835,N_32869);
or U41656 (N_41656,N_39774,N_34114);
nor U41657 (N_41657,N_37775,N_32909);
xnor U41658 (N_41658,N_35604,N_33272);
xnor U41659 (N_41659,N_37859,N_39476);
or U41660 (N_41660,N_35126,N_34462);
nand U41661 (N_41661,N_30062,N_31675);
nand U41662 (N_41662,N_32119,N_32571);
and U41663 (N_41663,N_34664,N_34614);
or U41664 (N_41664,N_33937,N_37031);
nor U41665 (N_41665,N_37208,N_38401);
or U41666 (N_41666,N_39786,N_31063);
nand U41667 (N_41667,N_31452,N_33936);
or U41668 (N_41668,N_30554,N_33749);
and U41669 (N_41669,N_35674,N_31833);
or U41670 (N_41670,N_30034,N_33957);
xnor U41671 (N_41671,N_37085,N_39220);
xor U41672 (N_41672,N_35133,N_32025);
nand U41673 (N_41673,N_31879,N_32538);
xor U41674 (N_41674,N_31668,N_35431);
nor U41675 (N_41675,N_32491,N_32391);
and U41676 (N_41676,N_33089,N_36284);
or U41677 (N_41677,N_31658,N_33321);
xor U41678 (N_41678,N_33365,N_38943);
xor U41679 (N_41679,N_36715,N_37358);
or U41680 (N_41680,N_34327,N_31763);
nand U41681 (N_41681,N_30597,N_39713);
nor U41682 (N_41682,N_38550,N_33759);
nor U41683 (N_41683,N_31523,N_36825);
or U41684 (N_41684,N_30476,N_37527);
nor U41685 (N_41685,N_32294,N_33978);
nand U41686 (N_41686,N_31129,N_30704);
or U41687 (N_41687,N_31688,N_37694);
nand U41688 (N_41688,N_32116,N_39146);
nor U41689 (N_41689,N_36928,N_35562);
or U41690 (N_41690,N_34506,N_33425);
nor U41691 (N_41691,N_30629,N_38695);
xor U41692 (N_41692,N_33927,N_31846);
and U41693 (N_41693,N_39423,N_33633);
nor U41694 (N_41694,N_38420,N_31484);
and U41695 (N_41695,N_30584,N_30224);
and U41696 (N_41696,N_32264,N_39935);
and U41697 (N_41697,N_33589,N_31151);
nand U41698 (N_41698,N_36958,N_30155);
nor U41699 (N_41699,N_34602,N_31520);
nor U41700 (N_41700,N_36088,N_31670);
nand U41701 (N_41701,N_30982,N_30898);
and U41702 (N_41702,N_39294,N_31788);
xor U41703 (N_41703,N_34325,N_38256);
and U41704 (N_41704,N_33569,N_33841);
or U41705 (N_41705,N_32613,N_38466);
or U41706 (N_41706,N_37712,N_30638);
xor U41707 (N_41707,N_36957,N_35506);
nor U41708 (N_41708,N_37329,N_33407);
and U41709 (N_41709,N_35158,N_35220);
xnor U41710 (N_41710,N_31932,N_35999);
xor U41711 (N_41711,N_30809,N_31898);
and U41712 (N_41712,N_37883,N_30628);
or U41713 (N_41713,N_34717,N_33076);
xnor U41714 (N_41714,N_33185,N_34047);
or U41715 (N_41715,N_37292,N_35963);
or U41716 (N_41716,N_38890,N_33879);
nor U41717 (N_41717,N_30556,N_35439);
xnor U41718 (N_41718,N_33854,N_38285);
xnor U41719 (N_41719,N_39816,N_31925);
xnor U41720 (N_41720,N_34112,N_35670);
xnor U41721 (N_41721,N_34592,N_37765);
nor U41722 (N_41722,N_31403,N_38887);
or U41723 (N_41723,N_32691,N_32823);
or U41724 (N_41724,N_30896,N_30884);
nor U41725 (N_41725,N_39453,N_38624);
xor U41726 (N_41726,N_37791,N_34938);
nand U41727 (N_41727,N_34104,N_39975);
nor U41728 (N_41728,N_35737,N_31280);
or U41729 (N_41729,N_34544,N_31592);
nand U41730 (N_41730,N_35847,N_34697);
nor U41731 (N_41731,N_38381,N_34862);
or U41732 (N_41732,N_37903,N_32153);
nor U41733 (N_41733,N_33409,N_30370);
nor U41734 (N_41734,N_36831,N_34843);
or U41735 (N_41735,N_34720,N_35983);
nor U41736 (N_41736,N_36636,N_31337);
or U41737 (N_41737,N_35804,N_31462);
and U41738 (N_41738,N_38953,N_32189);
xor U41739 (N_41739,N_35098,N_38022);
and U41740 (N_41740,N_32655,N_34305);
xor U41741 (N_41741,N_34496,N_30036);
nor U41742 (N_41742,N_37032,N_33642);
nor U41743 (N_41743,N_38902,N_36465);
xor U41744 (N_41744,N_38745,N_38933);
xor U41745 (N_41745,N_32687,N_30927);
nor U41746 (N_41746,N_34539,N_37363);
or U41747 (N_41747,N_36491,N_38607);
xor U41748 (N_41748,N_30234,N_30853);
nor U41749 (N_41749,N_36191,N_35055);
or U41750 (N_41750,N_36061,N_39870);
and U41751 (N_41751,N_37994,N_34328);
nand U41752 (N_41752,N_34840,N_37041);
nor U41753 (N_41753,N_36856,N_39988);
nor U41754 (N_41754,N_36370,N_36112);
xor U41755 (N_41755,N_39663,N_34815);
nand U41756 (N_41756,N_31305,N_35544);
nor U41757 (N_41757,N_37726,N_37701);
and U41758 (N_41758,N_38124,N_38823);
and U41759 (N_41759,N_37664,N_34874);
nor U41760 (N_41760,N_32162,N_30645);
xor U41761 (N_41761,N_37001,N_32763);
and U41762 (N_41762,N_32753,N_35759);
xor U41763 (N_41763,N_31036,N_31162);
nor U41764 (N_41764,N_35933,N_35758);
xor U41765 (N_41765,N_37613,N_36937);
xor U41766 (N_41766,N_38901,N_38023);
or U41767 (N_41767,N_37511,N_37865);
xnor U41768 (N_41768,N_31327,N_35976);
nor U41769 (N_41769,N_36064,N_32606);
and U41770 (N_41770,N_34554,N_39178);
nor U41771 (N_41771,N_36501,N_32947);
xor U41772 (N_41772,N_36546,N_30099);
nor U41773 (N_41773,N_36943,N_31516);
xnor U41774 (N_41774,N_32443,N_34510);
nand U41775 (N_41775,N_34169,N_32484);
xnor U41776 (N_41776,N_36509,N_33257);
nor U41777 (N_41777,N_36584,N_35178);
and U41778 (N_41778,N_31984,N_32111);
xor U41779 (N_41779,N_36959,N_31865);
nor U41780 (N_41780,N_33093,N_33160);
and U41781 (N_41781,N_35806,N_33067);
and U41782 (N_41782,N_34301,N_36898);
or U41783 (N_41783,N_35872,N_32965);
or U41784 (N_41784,N_37335,N_39843);
xnor U41785 (N_41785,N_36267,N_35721);
xnor U41786 (N_41786,N_32525,N_37510);
or U41787 (N_41787,N_37563,N_39396);
and U41788 (N_41788,N_32695,N_36407);
and U41789 (N_41789,N_30326,N_33915);
or U41790 (N_41790,N_32556,N_37201);
nand U41791 (N_41791,N_39443,N_38033);
nand U41792 (N_41792,N_33051,N_31443);
and U41793 (N_41793,N_39725,N_38742);
nand U41794 (N_41794,N_36592,N_39066);
nand U41795 (N_41795,N_33833,N_33505);
or U41796 (N_41796,N_35855,N_36687);
nand U41797 (N_41797,N_34996,N_36418);
or U41798 (N_41798,N_38037,N_31576);
xor U41799 (N_41799,N_30498,N_31259);
and U41800 (N_41800,N_32244,N_37704);
nand U41801 (N_41801,N_37837,N_36813);
xor U41802 (N_41802,N_39648,N_38498);
xor U41803 (N_41803,N_39509,N_33599);
nand U41804 (N_41804,N_31205,N_34378);
and U41805 (N_41805,N_31491,N_33340);
or U41806 (N_41806,N_30380,N_31258);
xor U41807 (N_41807,N_30836,N_32428);
and U41808 (N_41808,N_37197,N_31595);
nand U41809 (N_41809,N_36079,N_33553);
and U41810 (N_41810,N_34184,N_36324);
nand U41811 (N_41811,N_38092,N_36172);
xnor U41812 (N_41812,N_33000,N_31839);
nor U41813 (N_41813,N_35116,N_31051);
nand U41814 (N_41814,N_30267,N_33824);
and U41815 (N_41815,N_31602,N_35054);
xor U41816 (N_41816,N_31902,N_31813);
or U41817 (N_41817,N_33969,N_35024);
nor U41818 (N_41818,N_33720,N_38674);
or U41819 (N_41819,N_34340,N_30361);
or U41820 (N_41820,N_36274,N_39754);
and U41821 (N_41821,N_37533,N_33903);
nand U41822 (N_41822,N_38432,N_30333);
and U41823 (N_41823,N_39300,N_34233);
nand U41824 (N_41824,N_32408,N_37781);
or U41825 (N_41825,N_38105,N_37495);
nand U41826 (N_41826,N_36122,N_35796);
nand U41827 (N_41827,N_33929,N_30804);
or U41828 (N_41828,N_31574,N_35212);
xor U41829 (N_41829,N_32940,N_31567);
xnor U41830 (N_41830,N_39335,N_38958);
xnor U41831 (N_41831,N_34491,N_34825);
nor U41832 (N_41832,N_32856,N_38421);
nor U41833 (N_41833,N_31152,N_30091);
or U41834 (N_41834,N_34668,N_33162);
nand U41835 (N_41835,N_34038,N_31799);
or U41836 (N_41836,N_31648,N_32562);
xnor U41837 (N_41837,N_38061,N_36253);
nor U41838 (N_41838,N_34906,N_35546);
nor U41839 (N_41839,N_39731,N_39848);
nand U41840 (N_41840,N_30663,N_35839);
or U41841 (N_41841,N_31315,N_37900);
and U41842 (N_41842,N_37362,N_32972);
nor U41843 (N_41843,N_31667,N_39382);
nor U41844 (N_41844,N_32191,N_37158);
and U41845 (N_41845,N_37771,N_31816);
xor U41846 (N_41846,N_30293,N_30730);
xnor U41847 (N_41847,N_36399,N_34451);
nand U41848 (N_41848,N_37468,N_34147);
xor U41849 (N_41849,N_33539,N_38818);
and U41850 (N_41850,N_37749,N_30003);
or U41851 (N_41851,N_39638,N_38024);
or U41852 (N_41852,N_35414,N_35087);
nand U41853 (N_41853,N_37531,N_35200);
nor U41854 (N_41854,N_36263,N_32115);
nor U41855 (N_41855,N_35244,N_35329);
xor U41856 (N_41856,N_33497,N_37131);
and U41857 (N_41857,N_33041,N_34018);
and U41858 (N_41858,N_30004,N_32339);
xnor U41859 (N_41859,N_39236,N_36967);
or U41860 (N_41860,N_39049,N_34469);
and U41861 (N_41861,N_33224,N_31514);
and U41862 (N_41862,N_32870,N_36742);
nand U41863 (N_41863,N_33654,N_34936);
or U41864 (N_41864,N_39698,N_34974);
and U41865 (N_41865,N_30263,N_32875);
nand U41866 (N_41866,N_38612,N_33010);
xnor U41867 (N_41867,N_30085,N_37678);
or U41868 (N_41868,N_32957,N_30095);
nand U41869 (N_41869,N_32729,N_31927);
xor U41870 (N_41870,N_36355,N_30762);
and U41871 (N_41871,N_37467,N_32672);
or U41872 (N_41872,N_37117,N_38085);
nor U41873 (N_41873,N_34013,N_30146);
nor U41874 (N_41874,N_34593,N_34724);
and U41875 (N_41875,N_37599,N_31450);
and U41876 (N_41876,N_35106,N_31256);
nor U41877 (N_41877,N_32221,N_32359);
nor U41878 (N_41878,N_39841,N_30133);
or U41879 (N_41879,N_32820,N_38542);
or U41880 (N_41880,N_31089,N_38299);
xor U41881 (N_41881,N_37089,N_39331);
xor U41882 (N_41882,N_36900,N_34312);
or U41883 (N_41883,N_36458,N_33099);
xnor U41884 (N_41884,N_33925,N_37190);
or U41885 (N_41885,N_34263,N_35097);
nor U41886 (N_41886,N_32063,N_31868);
nor U41887 (N_41887,N_33803,N_35790);
nand U41888 (N_41888,N_35650,N_37520);
and U41889 (N_41889,N_37795,N_30720);
or U41890 (N_41890,N_35542,N_33738);
or U41891 (N_41891,N_36440,N_30921);
nor U41892 (N_41892,N_30713,N_36840);
nor U41893 (N_41893,N_36516,N_38812);
and U41894 (N_41894,N_39444,N_34577);
xor U41895 (N_41895,N_32380,N_36455);
nand U41896 (N_41896,N_37323,N_37787);
xor U41897 (N_41897,N_34146,N_35039);
xnor U41898 (N_41898,N_39896,N_31994);
or U41899 (N_41899,N_37288,N_38682);
xnor U41900 (N_41900,N_36302,N_32277);
or U41901 (N_41901,N_36244,N_36019);
nor U41902 (N_41902,N_34200,N_36938);
or U41903 (N_41903,N_34421,N_38443);
nor U41904 (N_41904,N_38106,N_33304);
or U41905 (N_41905,N_35834,N_37823);
nor U41906 (N_41906,N_39525,N_32011);
xor U41907 (N_41907,N_34922,N_38617);
xor U41908 (N_41908,N_30788,N_34991);
nand U41909 (N_41909,N_34162,N_34127);
xnor U41910 (N_41910,N_31369,N_33171);
nand U41911 (N_41911,N_33668,N_30210);
xnor U41912 (N_41912,N_37899,N_34624);
and U41913 (N_41913,N_31157,N_30086);
nor U41914 (N_41914,N_32859,N_33517);
nor U41915 (N_41915,N_33817,N_38543);
xor U41916 (N_41916,N_37786,N_36783);
nor U41917 (N_41917,N_35334,N_31930);
nand U41918 (N_41918,N_36673,N_38361);
or U41919 (N_41919,N_31466,N_31476);
xor U41920 (N_41920,N_34995,N_31593);
or U41921 (N_41921,N_32233,N_37679);
nor U41922 (N_41922,N_39137,N_35936);
or U41923 (N_41923,N_33330,N_30328);
and U41924 (N_41924,N_35538,N_32026);
or U41925 (N_41925,N_39921,N_32341);
and U41926 (N_41926,N_35799,N_33724);
and U41927 (N_41927,N_32442,N_35914);
or U41928 (N_41928,N_33946,N_30859);
and U41929 (N_41929,N_35301,N_34397);
xor U41930 (N_41930,N_38377,N_35092);
nor U41931 (N_41931,N_30966,N_33060);
nor U41932 (N_41932,N_32548,N_32169);
and U41933 (N_41933,N_34351,N_30962);
nand U41934 (N_41934,N_31859,N_34627);
xor U41935 (N_41935,N_34447,N_35617);
and U41936 (N_41936,N_33644,N_32499);
xor U41937 (N_41937,N_39241,N_31486);
nand U41938 (N_41938,N_36745,N_36379);
nand U41939 (N_41939,N_35350,N_36008);
nand U41940 (N_41940,N_31561,N_33952);
nand U41941 (N_41941,N_34492,N_36603);
nand U41942 (N_41942,N_37738,N_32485);
xor U41943 (N_41943,N_39742,N_33116);
xnor U41944 (N_41944,N_39944,N_38188);
nor U41945 (N_41945,N_37026,N_35017);
and U41946 (N_41946,N_36148,N_38497);
or U41947 (N_41947,N_31940,N_30702);
or U41948 (N_41948,N_38847,N_37547);
or U41949 (N_41949,N_35552,N_38775);
and U41950 (N_41950,N_39780,N_32961);
and U41951 (N_41951,N_34071,N_32560);
and U41952 (N_41952,N_34224,N_31880);
nor U41953 (N_41953,N_32816,N_31097);
and U41954 (N_41954,N_30043,N_31203);
or U41955 (N_41955,N_38865,N_31739);
nand U41956 (N_41956,N_32194,N_34588);
or U41957 (N_41957,N_35553,N_32545);
nand U41958 (N_41958,N_33415,N_33533);
nor U41959 (N_41959,N_36011,N_33214);
nand U41960 (N_41960,N_31557,N_32901);
or U41961 (N_41961,N_31569,N_35819);
and U41962 (N_41962,N_37261,N_36838);
or U41963 (N_41963,N_34020,N_37436);
or U41964 (N_41964,N_38159,N_34130);
xnor U41965 (N_41965,N_32592,N_39877);
nor U41966 (N_41966,N_33419,N_38446);
nor U41967 (N_41967,N_34073,N_31627);
nand U41968 (N_41968,N_30774,N_38796);
nand U41969 (N_41969,N_39333,N_35901);
or U41970 (N_41970,N_37206,N_31856);
or U41971 (N_41971,N_37526,N_30950);
nor U41972 (N_41972,N_35032,N_39884);
nor U41973 (N_41973,N_33991,N_32799);
nand U41974 (N_41974,N_36671,N_36323);
nand U41975 (N_41975,N_35895,N_34557);
nor U41976 (N_41976,N_31897,N_30150);
nand U41977 (N_41977,N_36914,N_33576);
nor U41978 (N_41978,N_30366,N_31234);
nor U41979 (N_41979,N_33848,N_39695);
nand U41980 (N_41980,N_37579,N_31683);
xor U41981 (N_41981,N_37139,N_30392);
nor U41982 (N_41982,N_38852,N_37473);
nor U41983 (N_41983,N_39171,N_39026);
nor U41984 (N_41984,N_37979,N_38210);
or U41985 (N_41985,N_37330,N_30354);
or U41986 (N_41986,N_39085,N_37393);
xnor U41987 (N_41987,N_35357,N_35765);
nand U41988 (N_41988,N_38386,N_39339);
or U41989 (N_41989,N_34126,N_34573);
and U41990 (N_41990,N_34847,N_38664);
and U41991 (N_41991,N_38926,N_31018);
xor U41992 (N_41992,N_32027,N_39398);
nand U41993 (N_41993,N_30867,N_35881);
or U41994 (N_41994,N_32640,N_30561);
and U41995 (N_41995,N_35191,N_33856);
and U41996 (N_41996,N_30414,N_36260);
nand U41997 (N_41997,N_30277,N_39536);
and U41998 (N_41998,N_39573,N_33842);
nor U41999 (N_41999,N_31490,N_36283);
and U42000 (N_42000,N_33660,N_33066);
nor U42001 (N_42001,N_37371,N_30816);
nand U42002 (N_42002,N_30834,N_38838);
and U42003 (N_42003,N_39620,N_37338);
nor U42004 (N_42004,N_37438,N_37426);
nand U42005 (N_42005,N_35501,N_35786);
nand U42006 (N_42006,N_30840,N_30462);
nor U42007 (N_42007,N_31938,N_31851);
nand U42008 (N_42008,N_33732,N_38526);
nand U42009 (N_42009,N_35747,N_39807);
nand U42010 (N_42010,N_33314,N_32275);
xnor U42011 (N_42011,N_31339,N_37145);
or U42012 (N_42012,N_34628,N_36059);
and U42013 (N_42013,N_32670,N_39495);
xnor U42014 (N_42014,N_37926,N_35950);
xor U42015 (N_42015,N_34168,N_32161);
xnor U42016 (N_42016,N_38658,N_32643);
and U42017 (N_42017,N_38603,N_39211);
and U42018 (N_42018,N_30865,N_36704);
nand U42019 (N_42019,N_36517,N_37466);
and U42020 (N_42020,N_36717,N_32967);
or U42021 (N_42021,N_32714,N_35769);
xnor U42022 (N_42022,N_33112,N_33510);
nand U42023 (N_42023,N_36004,N_37911);
or U42024 (N_42024,N_38165,N_36228);
and U42025 (N_42025,N_36350,N_36438);
nor U42026 (N_42026,N_37168,N_32842);
xor U42027 (N_42027,N_32580,N_30472);
nand U42028 (N_42028,N_32066,N_33447);
or U42029 (N_42029,N_36445,N_37630);
nand U42030 (N_42030,N_30107,N_30542);
and U42031 (N_42031,N_35560,N_37011);
or U42032 (N_42032,N_37646,N_34232);
nand U42033 (N_42033,N_31681,N_32426);
nor U42034 (N_42034,N_36460,N_35917);
xor U42035 (N_42035,N_30486,N_31580);
or U42036 (N_42036,N_30890,N_36801);
xnor U42037 (N_42037,N_33530,N_34183);
nor U42038 (N_42038,N_32438,N_32702);
or U42039 (N_42039,N_36417,N_30559);
nor U42040 (N_42040,N_37875,N_35021);
xor U42041 (N_42041,N_30482,N_30273);
or U42042 (N_42042,N_38799,N_31293);
xnor U42043 (N_42043,N_34785,N_31004);
nor U42044 (N_42044,N_33869,N_38855);
or U42045 (N_42045,N_38802,N_39609);
or U42046 (N_42046,N_38507,N_39330);
nand U42047 (N_42047,N_33013,N_34429);
nor U42048 (N_42048,N_33649,N_35829);
xnor U42049 (N_42049,N_38830,N_34637);
or U42050 (N_42050,N_39139,N_38535);
nand U42051 (N_42051,N_33596,N_36154);
nand U42052 (N_42052,N_38566,N_35575);
and U42053 (N_42053,N_37447,N_37887);
or U42054 (N_42054,N_38738,N_32926);
and U42055 (N_42055,N_37696,N_38766);
or U42056 (N_42056,N_30367,N_34878);
or U42057 (N_42057,N_32353,N_30318);
or U42058 (N_42058,N_32302,N_32245);
xnor U42059 (N_42059,N_37597,N_38169);
nor U42060 (N_42060,N_39867,N_32971);
nor U42061 (N_42061,N_31693,N_34801);
nor U42062 (N_42062,N_34500,N_31992);
nor U42063 (N_42063,N_39188,N_37753);
xor U42064 (N_42064,N_37063,N_32841);
and U42065 (N_42065,N_35726,N_33772);
and U42066 (N_42066,N_39633,N_34181);
nor U42067 (N_42067,N_32067,N_37440);
nor U42068 (N_42068,N_36750,N_38019);
or U42069 (N_42069,N_32433,N_38362);
xor U42070 (N_42070,N_34849,N_32223);
xor U42071 (N_42071,N_36264,N_38095);
or U42072 (N_42072,N_31264,N_30709);
and U42073 (N_42073,N_35411,N_37382);
or U42074 (N_42074,N_36216,N_39697);
and U42075 (N_42075,N_35565,N_37886);
nand U42076 (N_42076,N_35682,N_33121);
or U42077 (N_42077,N_39323,N_32214);
nand U42078 (N_42078,N_32930,N_33179);
or U42079 (N_42079,N_39217,N_38833);
nand U42080 (N_42080,N_38614,N_36140);
and U42081 (N_42081,N_37123,N_36652);
xnor U42082 (N_42082,N_33519,N_35541);
or U42083 (N_42083,N_30266,N_33485);
nand U42084 (N_42084,N_33870,N_36487);
or U42085 (N_42085,N_38643,N_39210);
or U42086 (N_42086,N_32490,N_32089);
and U42087 (N_42087,N_31911,N_31112);
nor U42088 (N_42088,N_32520,N_37813);
or U42089 (N_42089,N_33613,N_39344);
nand U42090 (N_42090,N_35050,N_34267);
nand U42091 (N_42091,N_36666,N_33371);
and U42092 (N_42092,N_36500,N_35014);
nor U42093 (N_42093,N_33997,N_39551);
or U42094 (N_42094,N_30078,N_37374);
xor U42095 (N_42095,N_30684,N_39270);
xor U42096 (N_42096,N_36728,N_39793);
nand U42097 (N_42097,N_37660,N_33216);
xor U42098 (N_42098,N_31544,N_37141);
xor U42099 (N_42099,N_31749,N_35474);
nor U42100 (N_42100,N_32675,N_37070);
nand U42101 (N_42101,N_31460,N_35035);
nand U42102 (N_42102,N_36513,N_38400);
xnor U42103 (N_42103,N_32578,N_36508);
xor U42104 (N_42104,N_32568,N_38565);
and U42105 (N_42105,N_32413,N_37739);
nand U42106 (N_42106,N_32260,N_36349);
xor U42107 (N_42107,N_30139,N_37260);
nand U42108 (N_42108,N_37838,N_38344);
nor U42109 (N_42109,N_38713,N_35229);
nor U42110 (N_42110,N_32781,N_31038);
or U42111 (N_42111,N_30748,N_37230);
or U42112 (N_42112,N_37492,N_30070);
nor U42113 (N_42113,N_35622,N_39346);
xor U42114 (N_42114,N_32452,N_38254);
xnor U42115 (N_42115,N_34182,N_31958);
or U42116 (N_42116,N_36564,N_35981);
nor U42117 (N_42117,N_34037,N_32780);
nor U42118 (N_42118,N_37593,N_38261);
and U42119 (N_42119,N_32249,N_38689);
or U42120 (N_42120,N_32314,N_30470);
nand U42121 (N_42121,N_32700,N_33127);
nand U42122 (N_42122,N_31944,N_31494);
nand U42123 (N_42123,N_35374,N_30147);
or U42124 (N_42124,N_37587,N_33384);
and U42125 (N_42125,N_36116,N_30296);
and U42126 (N_42126,N_32579,N_39629);
nand U42127 (N_42127,N_33451,N_38453);
nand U42128 (N_42128,N_33325,N_38001);
and U42129 (N_42129,N_35272,N_32906);
or U42130 (N_42130,N_39343,N_37099);
or U42131 (N_42131,N_30592,N_34370);
and U42132 (N_42132,N_32519,N_38040);
nand U42133 (N_42133,N_32787,N_33153);
xor U42134 (N_42134,N_31996,N_39537);
nand U42135 (N_42135,N_31606,N_33107);
xor U42136 (N_42136,N_39275,N_37024);
or U42137 (N_42137,N_30071,N_34142);
and U42138 (N_42138,N_36314,N_38967);
xnor U42139 (N_42139,N_39995,N_36442);
or U42140 (N_42140,N_36340,N_35628);
and U42141 (N_42141,N_30279,N_38171);
or U42142 (N_42142,N_36158,N_31446);
and U42143 (N_42143,N_33518,N_36390);
xor U42144 (N_42144,N_34272,N_33651);
and U42145 (N_42145,N_36436,N_32893);
nand U42146 (N_42146,N_35882,N_35997);
or U42147 (N_42147,N_36111,N_37624);
or U42148 (N_42148,N_39177,N_37381);
nor U42149 (N_42149,N_30864,N_30513);
nand U42150 (N_42150,N_31425,N_38477);
xnor U42151 (N_42151,N_30943,N_38272);
or U42152 (N_42152,N_36696,N_36730);
nand U42153 (N_42153,N_36805,N_34934);
nor U42154 (N_42154,N_30435,N_31487);
nand U42155 (N_42155,N_33168,N_36261);
or U42156 (N_42156,N_31844,N_35962);
and U42157 (N_42157,N_39655,N_32597);
or U42158 (N_42158,N_38556,N_38772);
and U42159 (N_42159,N_35858,N_36930);
nand U42160 (N_42160,N_34279,N_33758);
and U42161 (N_42161,N_33405,N_32285);
xnor U42162 (N_42162,N_36345,N_39127);
nand U42163 (N_42163,N_30925,N_32205);
or U42164 (N_42164,N_31030,N_36369);
xor U42165 (N_42165,N_30810,N_34499);
xnor U42166 (N_42166,N_30618,N_34065);
nor U42167 (N_42167,N_39155,N_39472);
or U42168 (N_42168,N_35067,N_30808);
or U42169 (N_42169,N_30450,N_32782);
or U42170 (N_42170,N_30052,N_35461);
or U42171 (N_42171,N_36917,N_34925);
nand U42172 (N_42172,N_38077,N_34959);
and U42173 (N_42173,N_33502,N_37256);
nand U42174 (N_42174,N_36031,N_31186);
xor U42175 (N_42175,N_30121,N_38616);
nand U42176 (N_42176,N_38829,N_39072);
nand U42177 (N_42177,N_30763,N_31498);
or U42178 (N_42178,N_37068,N_33348);
or U42179 (N_42179,N_32826,N_30219);
nand U42180 (N_42180,N_36351,N_36962);
and U42181 (N_42181,N_31970,N_34417);
or U42182 (N_42182,N_30609,N_34344);
xor U42183 (N_42183,N_33342,N_34480);
xor U42184 (N_42184,N_31760,N_37986);
nor U42185 (N_42185,N_37211,N_36472);
nand U42186 (N_42186,N_33075,N_35500);
or U42187 (N_42187,N_32463,N_37052);
xnor U42188 (N_42188,N_30477,N_39122);
nand U42189 (N_42189,N_34082,N_37848);
nand U42190 (N_42190,N_38207,N_32683);
xnor U42191 (N_42191,N_32326,N_33269);
nor U42192 (N_42192,N_33288,N_35513);
nand U42193 (N_42193,N_33183,N_32512);
and U42194 (N_42194,N_36222,N_38029);
nand U42195 (N_42195,N_39112,N_34489);
nor U42196 (N_42196,N_38946,N_31819);
nor U42197 (N_42197,N_30473,N_38305);
and U42198 (N_42198,N_38553,N_38202);
and U42199 (N_42199,N_34736,N_32609);
nand U42200 (N_42200,N_33976,N_37909);
nand U42201 (N_42201,N_34025,N_34851);
xor U42202 (N_42202,N_35856,N_32197);
xnor U42203 (N_42203,N_34004,N_32065);
and U42204 (N_42204,N_37376,N_39758);
nor U42205 (N_42205,N_32045,N_36201);
xnor U42206 (N_42206,N_39766,N_32819);
and U42207 (N_42207,N_34810,N_38127);
nor U42208 (N_42208,N_38530,N_31150);
xnor U42209 (N_42209,N_33395,N_36600);
nor U42210 (N_42210,N_34456,N_35019);
xnor U42211 (N_42211,N_38622,N_31736);
nand U42212 (N_42212,N_34080,N_33810);
xor U42213 (N_42213,N_35630,N_30766);
xor U42214 (N_42214,N_30871,N_37212);
xnor U42215 (N_42215,N_37935,N_35740);
nand U42216 (N_42216,N_36412,N_34329);
or U42217 (N_42217,N_35317,N_36678);
and U42218 (N_42218,N_34940,N_39368);
xnor U42219 (N_42219,N_35112,N_33689);
xnor U42220 (N_42220,N_39908,N_37162);
and U42221 (N_42221,N_30206,N_39741);
or U42222 (N_42222,N_34965,N_38732);
or U42223 (N_42223,N_35867,N_38205);
nor U42224 (N_42224,N_39840,N_37699);
and U42225 (N_42225,N_37584,N_39045);
nor U42226 (N_42226,N_31161,N_39868);
and U42227 (N_42227,N_32388,N_30676);
nand U42228 (N_42228,N_30987,N_31645);
xor U42229 (N_42229,N_30665,N_30919);
nand U42230 (N_42230,N_31284,N_38778);
nand U42231 (N_42231,N_37500,N_30687);
xnor U42232 (N_42232,N_32584,N_39605);
nand U42233 (N_42233,N_30992,N_30764);
or U42234 (N_42234,N_34087,N_30032);
nor U42235 (N_42235,N_39302,N_31297);
nand U42236 (N_42236,N_32769,N_35265);
nand U42237 (N_42237,N_35969,N_33053);
nand U42238 (N_42238,N_34655,N_36075);
xnor U42239 (N_42239,N_39153,N_39287);
or U42240 (N_42240,N_30746,N_33376);
xnor U42241 (N_42241,N_39838,N_35451);
xor U42242 (N_42242,N_31231,N_35135);
and U42243 (N_42243,N_38359,N_36665);
nand U42244 (N_42244,N_31800,N_33364);
or U42245 (N_42245,N_33143,N_36051);
nor U42246 (N_42246,N_32062,N_39421);
nand U42247 (N_42247,N_31485,N_31743);
nand U42248 (N_42248,N_31002,N_35122);
xor U42249 (N_42249,N_35771,N_37819);
or U42250 (N_42250,N_39973,N_30144);
nor U42251 (N_42251,N_39215,N_39876);
nor U42252 (N_42252,N_33942,N_38229);
and U42253 (N_42253,N_31726,N_32493);
nor U42254 (N_42254,N_37392,N_34902);
nand U42255 (N_42255,N_32796,N_32942);
nand U42256 (N_42256,N_33616,N_34928);
nand U42257 (N_42257,N_36193,N_37322);
xor U42258 (N_42258,N_35056,N_34275);
xor U42259 (N_42259,N_34555,N_33867);
and U42260 (N_42260,N_30961,N_31155);
xnor U42261 (N_42261,N_35507,N_35703);
or U42262 (N_42262,N_36180,N_36476);
and U42263 (N_42263,N_36192,N_33828);
and U42264 (N_42264,N_39505,N_38720);
nor U42265 (N_42265,N_35780,N_38413);
nor U42266 (N_42266,N_36736,N_39791);
and U42267 (N_42267,N_36150,N_30894);
nand U42268 (N_42268,N_33237,N_31542);
or U42269 (N_42269,N_33791,N_37972);
xnor U42270 (N_42270,N_33413,N_34806);
or U42271 (N_42271,N_33235,N_38055);
and U42272 (N_42272,N_35660,N_37855);
xnor U42273 (N_42273,N_39358,N_35072);
nor U42274 (N_42274,N_32237,N_37897);
or U42275 (N_42275,N_33389,N_34755);
or U42276 (N_42276,N_32015,N_36740);
nand U42277 (N_42277,N_36483,N_33681);
and U42278 (N_42278,N_33721,N_31492);
nand U42279 (N_42279,N_30499,N_37551);
nand U42280 (N_42280,N_32614,N_39547);
nor U42281 (N_42281,N_38076,N_33712);
nor U42282 (N_42282,N_35152,N_38425);
and U42283 (N_42283,N_36477,N_31034);
nand U42284 (N_42284,N_37343,N_35555);
nand U42285 (N_42285,N_30526,N_36775);
or U42286 (N_42286,N_32096,N_34475);
or U42287 (N_42287,N_34068,N_35488);
xor U42288 (N_42288,N_38107,N_34729);
nand U42289 (N_42289,N_33015,N_39082);
or U42290 (N_42290,N_34626,N_37799);
or U42291 (N_42291,N_34822,N_30814);
nand U42292 (N_42292,N_36799,N_30016);
nand U42293 (N_42293,N_32970,N_30664);
nand U42294 (N_42294,N_32296,N_38719);
nor U42295 (N_42295,N_39668,N_35358);
nand U42296 (N_42296,N_34153,N_36723);
nand U42297 (N_42297,N_38921,N_33394);
or U42298 (N_42298,N_37982,N_35701);
xor U42299 (N_42299,N_30232,N_37642);
and U42300 (N_42300,N_30184,N_35070);
and U42301 (N_42301,N_39811,N_34284);
or U42302 (N_42302,N_35772,N_31948);
or U42303 (N_42303,N_34099,N_30378);
nand U42304 (N_42304,N_35078,N_33350);
nand U42305 (N_42305,N_33449,N_31686);
nand U42306 (N_42306,N_37259,N_38521);
nand U42307 (N_42307,N_35031,N_36276);
nand U42308 (N_42308,N_37071,N_31716);
nor U42309 (N_42309,N_35514,N_34617);
nor U42310 (N_42310,N_32447,N_31849);
nand U42311 (N_42311,N_39997,N_31107);
nand U42312 (N_42312,N_33264,N_38500);
and U42313 (N_42313,N_34753,N_31267);
nor U42314 (N_42314,N_37196,N_38763);
nand U42315 (N_42315,N_31401,N_35764);
or U42316 (N_42316,N_38826,N_31126);
and U42317 (N_42317,N_33821,N_33150);
nand U42318 (N_42318,N_39893,N_38849);
xor U42319 (N_42319,N_34334,N_34719);
nand U42320 (N_42320,N_34505,N_38102);
nor U42321 (N_42321,N_34803,N_36188);
xor U42322 (N_42322,N_34414,N_35247);
nand U42323 (N_42323,N_30192,N_37092);
nand U42324 (N_42324,N_32845,N_39175);
and U42325 (N_42325,N_35922,N_37400);
nand U42326 (N_42326,N_35370,N_31312);
nand U42327 (N_42327,N_31905,N_32916);
or U42328 (N_42328,N_31399,N_37539);
and U42329 (N_42329,N_36080,N_38806);
nand U42330 (N_42330,N_38963,N_36296);
xnor U42331 (N_42331,N_35520,N_34537);
or U42332 (N_42332,N_38948,N_35365);
xor U42333 (N_42333,N_37360,N_39061);
xnor U42334 (N_42334,N_32136,N_37252);
nand U42335 (N_42335,N_32473,N_34732);
nand U42336 (N_42336,N_39627,N_36647);
xor U42337 (N_42337,N_34904,N_30830);
nor U42338 (N_42338,N_38600,N_31980);
nor U42339 (N_42339,N_35564,N_33718);
or U42340 (N_42340,N_34139,N_36036);
nand U42341 (N_42341,N_39452,N_36490);
nand U42342 (N_42342,N_36520,N_38277);
nand U42343 (N_42343,N_39955,N_34643);
nand U42344 (N_42344,N_39170,N_37609);
xnor U42345 (N_42345,N_37389,N_34315);
or U42346 (N_42346,N_36559,N_32404);
nor U42347 (N_42347,N_32936,N_34708);
nor U42348 (N_42348,N_36087,N_35472);
xor U42349 (N_42349,N_36670,N_32647);
nand U42350 (N_42350,N_32698,N_31703);
or U42351 (N_42351,N_33077,N_39062);
nand U42352 (N_42352,N_32091,N_36589);
nor U42353 (N_42353,N_39386,N_38919);
nor U42354 (N_42354,N_37479,N_36049);
nor U42355 (N_42355,N_37824,N_30648);
or U42356 (N_42356,N_39393,N_38101);
nand U42357 (N_42357,N_38481,N_34384);
nand U42358 (N_42358,N_39286,N_31945);
xor U42359 (N_42359,N_31375,N_39777);
or U42360 (N_42360,N_38898,N_33601);
and U42361 (N_42361,N_33698,N_34534);
nand U42362 (N_42362,N_38589,N_34441);
nand U42363 (N_42363,N_32963,N_32641);
xnor U42364 (N_42364,N_36332,N_32468);
xor U42365 (N_42365,N_39110,N_36733);
and U42366 (N_42366,N_31075,N_33556);
and U42367 (N_42367,N_35649,N_35113);
and U42368 (N_42368,N_34779,N_37907);
nor U42369 (N_42369,N_36066,N_33091);
or U42370 (N_42370,N_33427,N_33072);
xnor U42371 (N_42371,N_34256,N_30761);
xor U42372 (N_42372,N_33597,N_35563);
and U42373 (N_42373,N_30000,N_35583);
or U42374 (N_42374,N_35921,N_30524);
nor U42375 (N_42375,N_30817,N_33770);
nand U42376 (N_42376,N_36894,N_37191);
xor U42377 (N_42377,N_31537,N_32309);
xnor U42378 (N_42378,N_38900,N_39348);
nor U42379 (N_42379,N_32495,N_36896);
or U42380 (N_42380,N_30420,N_31221);
and U42381 (N_42381,N_34872,N_35750);
xnor U42382 (N_42382,N_35891,N_39882);
nand U42383 (N_42383,N_39151,N_32377);
nand U42384 (N_42384,N_35582,N_38657);
or U42385 (N_42385,N_30799,N_37002);
and U42386 (N_42386,N_32744,N_32270);
and U42387 (N_42387,N_30650,N_38066);
or U42388 (N_42388,N_39208,N_36888);
or U42389 (N_42389,N_37538,N_39101);
and U42390 (N_42390,N_35809,N_37807);
or U42391 (N_42391,N_35730,N_35368);
or U42392 (N_42392,N_30419,N_31691);
and U42393 (N_42393,N_30096,N_38166);
and U42394 (N_42394,N_35004,N_37059);
and U42395 (N_42395,N_36030,N_38876);
and U42396 (N_42396,N_30596,N_32596);
xor U42397 (N_42397,N_39593,N_36651);
or U42398 (N_42398,N_33520,N_38724);
xnor U42399 (N_42399,N_39728,N_33345);
and U42400 (N_42400,N_32236,N_39355);
nor U42401 (N_42401,N_36845,N_38851);
nor U42402 (N_42402,N_34163,N_39523);
nor U42403 (N_42403,N_34412,N_30574);
and U42404 (N_42404,N_39727,N_32546);
nand U42405 (N_42405,N_35190,N_30904);
xor U42406 (N_42406,N_32832,N_39124);
nand U42407 (N_42407,N_31793,N_34629);
nand U42408 (N_42408,N_34765,N_31744);
and U42409 (N_42409,N_37706,N_39063);
xnor U42410 (N_42410,N_31910,N_36067);
nor U42411 (N_42411,N_33786,N_30959);
xor U42412 (N_42412,N_35646,N_36887);
xor U42413 (N_42413,N_34245,N_35659);
and U42414 (N_42414,N_37155,N_35707);
and U42415 (N_42415,N_36252,N_38927);
xnor U42416 (N_42416,N_38463,N_33268);
nand U42417 (N_42417,N_32526,N_35672);
and U42418 (N_42418,N_34490,N_34152);
xnor U42419 (N_42419,N_36927,N_30087);
xor U42420 (N_42420,N_33439,N_39479);
nand U42421 (N_42421,N_34229,N_31477);
nor U42422 (N_42422,N_38999,N_30507);
nand U42423 (N_42423,N_34238,N_38774);
xnor U42424 (N_42424,N_31848,N_31579);
nand U42425 (N_42425,N_33683,N_37082);
or U42426 (N_42426,N_30430,N_31292);
and U42427 (N_42427,N_38378,N_36022);
or U42428 (N_42428,N_30535,N_35655);
nand U42429 (N_42429,N_35587,N_39558);
and U42430 (N_42430,N_36243,N_34390);
xnor U42431 (N_42431,N_32246,N_36538);
nor U42432 (N_42432,N_35180,N_36387);
nor U42433 (N_42433,N_37923,N_32298);
or U42434 (N_42434,N_38690,N_36615);
xnor U42435 (N_42435,N_33299,N_30661);
or U42436 (N_42436,N_34283,N_35323);
nor U42437 (N_42437,N_30723,N_34034);
nor U42438 (N_42438,N_31978,N_38154);
or U42439 (N_42439,N_33954,N_34868);
xnor U42440 (N_42440,N_37916,N_33809);
or U42441 (N_42441,N_37340,N_39184);
nor U42442 (N_42442,N_36464,N_33491);
nand U42443 (N_42443,N_36315,N_31330);
and U42444 (N_42444,N_36044,N_38032);
nor U42445 (N_42445,N_37453,N_34019);
nand U42446 (N_42446,N_35181,N_32678);
or U42447 (N_42447,N_33310,N_36362);
nand U42448 (N_42448,N_36346,N_35189);
nor U42449 (N_42449,N_37921,N_38560);
xor U42450 (N_42450,N_38042,N_35479);
nor U42451 (N_42451,N_39883,N_35972);
or U42452 (N_42452,N_31396,N_32486);
or U42453 (N_42453,N_33667,N_31068);
and U42454 (N_42454,N_38218,N_31669);
nand U42455 (N_42455,N_35381,N_33618);
and U42456 (N_42456,N_32595,N_35624);
xor U42457 (N_42457,N_35224,N_37140);
xnor U42458 (N_42458,N_38380,N_31085);
or U42459 (N_42459,N_37888,N_32958);
or U42460 (N_42460,N_35234,N_37138);
nand U42461 (N_42461,N_38438,N_37302);
and U42462 (N_42462,N_35321,N_39530);
xnor U42463 (N_42463,N_36289,N_30506);
nand U42464 (N_42464,N_31676,N_34981);
and U42465 (N_42465,N_38252,N_35194);
nand U42466 (N_42466,N_31115,N_33793);
or U42467 (N_42467,N_33374,N_30394);
xor U42468 (N_42468,N_30550,N_30689);
nand U42469 (N_42469,N_37481,N_37662);
xor U42470 (N_42470,N_37060,N_39739);
nor U42471 (N_42471,N_33424,N_37577);
or U42472 (N_42472,N_33542,N_30541);
or U42473 (N_42473,N_39305,N_34392);
xor U42474 (N_42474,N_32049,N_36804);
nor U42475 (N_42475,N_37820,N_31087);
nand U42476 (N_42476,N_36507,N_34896);
xnor U42477 (N_42477,N_30454,N_37913);
nor U42478 (N_42478,N_38143,N_30640);
or U42479 (N_42479,N_39515,N_38114);
nor U42480 (N_42480,N_30538,N_38721);
nand U42481 (N_42481,N_35932,N_36174);
nand U42482 (N_42482,N_38043,N_35923);
nor U42483 (N_42483,N_35337,N_30199);
xnor U42484 (N_42484,N_34321,N_33934);
xor U42485 (N_42485,N_34113,N_30566);
or U42486 (N_42486,N_30741,N_33297);
nor U42487 (N_42487,N_34701,N_38240);
or U42488 (N_42488,N_39503,N_33661);
and U42489 (N_42489,N_30221,N_39795);
xnor U42490 (N_42490,N_33538,N_32619);
and U42491 (N_42491,N_37077,N_37585);
nand U42492 (N_42492,N_34742,N_33228);
nand U42493 (N_42493,N_30173,N_36078);
or U42494 (N_42494,N_34768,N_32361);
xor U42495 (N_42495,N_32733,N_30320);
or U42496 (N_42496,N_30717,N_37796);
nor U42497 (N_42497,N_36980,N_39231);
nor U42498 (N_42498,N_32884,N_31232);
or U42499 (N_42499,N_33331,N_36657);
xor U42500 (N_42500,N_38885,N_32072);
and U42501 (N_42501,N_36361,N_37794);
xor U42502 (N_42502,N_34675,N_36735);
and U42503 (N_42503,N_36971,N_30451);
nor U42504 (N_42504,N_32343,N_35103);
and U42505 (N_42505,N_37928,N_35047);
or U42506 (N_42506,N_37311,N_36774);
or U42507 (N_42507,N_31021,N_35558);
and U42508 (N_42508,N_33904,N_34251);
xnor U42509 (N_42509,N_39871,N_32995);
xor U42510 (N_42510,N_37737,N_38889);
nand U42511 (N_42511,N_34914,N_35688);
or U42512 (N_42512,N_34055,N_31666);
nor U42513 (N_42513,N_31318,N_30558);
xnor U42514 (N_42514,N_38932,N_31834);
xor U42515 (N_42515,N_37090,N_31384);
nand U42516 (N_42516,N_39073,N_35470);
nor U42517 (N_42517,N_35980,N_35264);
xnor U42518 (N_42518,N_30832,N_31803);
and U42519 (N_42519,N_31095,N_38540);
or U42520 (N_42520,N_31374,N_37192);
nand U42521 (N_42521,N_35253,N_39597);
or U42522 (N_42522,N_31055,N_37744);
or U42523 (N_42523,N_30035,N_39332);
nor U42524 (N_42524,N_30659,N_32482);
xor U42525 (N_42525,N_37119,N_33337);
nand U42526 (N_42526,N_33684,N_30902);
nor U42527 (N_42527,N_36554,N_31525);
xor U42528 (N_42528,N_38118,N_32810);
nor U42529 (N_42529,N_38339,N_33469);
nor U42530 (N_42530,N_35173,N_39314);
nand U42531 (N_42531,N_39794,N_33743);
xor U42532 (N_42532,N_31664,N_32807);
xnor U42533 (N_42533,N_37687,N_35601);
nor U42534 (N_42534,N_33139,N_32715);
and U42535 (N_42535,N_34817,N_39652);
xnor U42536 (N_42536,N_30800,N_30970);
or U42537 (N_42537,N_33101,N_33229);
or U42538 (N_42538,N_33799,N_30412);
nor U42539 (N_42539,N_33897,N_38395);
xnor U42540 (N_42540,N_30290,N_37778);
nand U42541 (N_42541,N_35739,N_35868);
nand U42542 (N_42542,N_38787,N_39863);
and U42543 (N_42543,N_32661,N_39650);
or U42544 (N_42544,N_35393,N_36820);
nand U42545 (N_42545,N_39013,N_33059);
xor U42546 (N_42546,N_38857,N_31404);
xnor U42547 (N_42547,N_31174,N_36540);
nand U42548 (N_42548,N_33047,N_37451);
nor U42549 (N_42549,N_37605,N_35863);
xor U42550 (N_42550,N_35464,N_34108);
or U42551 (N_42551,N_34622,N_31056);
and U42552 (N_42552,N_37444,N_37194);
or U42553 (N_42553,N_34471,N_31891);
or U42554 (N_42554,N_36871,N_37226);
xor U42555 (N_42555,N_36065,N_30821);
and U42556 (N_42556,N_30563,N_33715);
and U42557 (N_42557,N_34164,N_33967);
nand U42558 (N_42558,N_39806,N_31247);
xor U42559 (N_42559,N_31072,N_35184);
or U42560 (N_42560,N_33727,N_35377);
nor U42561 (N_42561,N_38473,N_37964);
nand U42562 (N_42562,N_39578,N_37633);
nand U42563 (N_42563,N_36903,N_34799);
or U42564 (N_42564,N_37882,N_34740);
xnor U42565 (N_42565,N_33521,N_30485);
or U42566 (N_42566,N_34800,N_33548);
nor U42567 (N_42567,N_34987,N_31882);
nor U42568 (N_42568,N_36119,N_33385);
or U42569 (N_42569,N_30779,N_35635);
nor U42570 (N_42570,N_35346,N_34360);
xor U42571 (N_42571,N_35787,N_32469);
or U42572 (N_42572,N_35459,N_39891);
and U42573 (N_42573,N_33463,N_33242);
nor U42574 (N_42574,N_35221,N_37805);
or U42575 (N_42575,N_30271,N_35627);
nor U42576 (N_42576,N_36771,N_30182);
and U42577 (N_42577,N_34609,N_36769);
or U42578 (N_42578,N_31400,N_36416);
xnor U42579 (N_42579,N_36234,N_36788);
and U42580 (N_42580,N_32121,N_30228);
xnor U42581 (N_42581,N_32242,N_35924);
nand U42582 (N_42582,N_32911,N_33951);
and U42583 (N_42583,N_38004,N_38295);
or U42584 (N_42584,N_34494,N_37889);
and U42585 (N_42585,N_37866,N_35108);
or U42586 (N_42586,N_34076,N_39354);
or U42587 (N_42587,N_30674,N_36953);
or U42588 (N_42588,N_31289,N_30718);
and U42589 (N_42589,N_31325,N_39706);
nor U42590 (N_42590,N_35947,N_32023);
nand U42591 (N_42591,N_39229,N_35927);
and U42592 (N_42592,N_38067,N_37417);
nor U42593 (N_42593,N_33474,N_32110);
and U42594 (N_42594,N_37341,N_30715);
and U42595 (N_42595,N_37146,N_35814);
nor U42596 (N_42596,N_39531,N_30824);
xor U42597 (N_42597,N_32208,N_36906);
and U42598 (N_42598,N_32677,N_30006);
nor U42599 (N_42599,N_30391,N_36525);
xor U42600 (N_42600,N_36716,N_31752);
nand U42601 (N_42601,N_39751,N_39542);
and U42602 (N_42602,N_35065,N_35728);
nand U42603 (N_42603,N_32168,N_38913);
and U42604 (N_42604,N_37294,N_37954);
or U42605 (N_42605,N_35353,N_35231);
and U42606 (N_42606,N_35639,N_32722);
nor U42607 (N_42607,N_33377,N_37187);
and U42608 (N_42608,N_33441,N_31414);
and U42609 (N_42609,N_37927,N_31066);
and U42610 (N_42610,N_32400,N_31565);
nand U42611 (N_42611,N_38345,N_33034);
or U42612 (N_42612,N_37233,N_31394);
nor U42613 (N_42613,N_30815,N_33639);
nand U42614 (N_42614,N_33431,N_34385);
nor U42615 (N_42615,N_32773,N_32518);
xnor U42616 (N_42616,N_32725,N_36058);
or U42617 (N_42617,N_35456,N_35663);
nand U42618 (N_42618,N_35652,N_32226);
nand U42619 (N_42619,N_39458,N_36695);
nor U42620 (N_42620,N_33352,N_38879);
nor U42621 (N_42621,N_34407,N_37519);
and U42622 (N_42622,N_38312,N_31518);
and U42623 (N_42623,N_37628,N_35591);
xor U42624 (N_42624,N_32502,N_35729);
nand U42625 (N_42625,N_37018,N_30441);
xor U42626 (N_42626,N_39324,N_38142);
xnor U42627 (N_42627,N_30154,N_38348);
nor U42628 (N_42628,N_36933,N_31349);
and U42629 (N_42629,N_38649,N_34246);
or U42630 (N_42630,N_35645,N_38980);
xnor U42631 (N_42631,N_33941,N_30373);
nor U42632 (N_42632,N_34682,N_35679);
nor U42633 (N_42633,N_30928,N_36823);
nand U42634 (N_42634,N_32703,N_31546);
nor U42635 (N_42635,N_32699,N_39684);
nor U42636 (N_42636,N_30969,N_36622);
xnor U42637 (N_42637,N_31104,N_36235);
nor U42638 (N_42638,N_30751,N_34109);
nand U42639 (N_42639,N_32253,N_37412);
nor U42640 (N_42640,N_33797,N_36784);
or U42641 (N_42641,N_33109,N_36375);
or U42642 (N_42642,N_37922,N_30994);
xnor U42643 (N_42643,N_30051,N_31195);
or U42644 (N_42644,N_30591,N_39422);
or U42645 (N_42645,N_39070,N_31682);
nand U42646 (N_42646,N_32895,N_38733);
or U42647 (N_42647,N_37355,N_31060);
or U42648 (N_42648,N_32576,N_31229);
nor U42649 (N_42649,N_33058,N_30903);
or U42650 (N_42650,N_33225,N_33947);
or U42651 (N_42651,N_32555,N_33111);
nor U42652 (N_42652,N_33083,N_36213);
and U42653 (N_42653,N_39289,N_37713);
or U42654 (N_42654,N_37039,N_38162);
or U42655 (N_42655,N_31214,N_38739);
nand U42656 (N_42656,N_39367,N_37534);
and U42657 (N_42657,N_36258,N_30395);
nand U42658 (N_42658,N_34319,N_34564);
nand U42659 (N_42659,N_34377,N_39885);
or U42660 (N_42660,N_38703,N_33024);
or U42661 (N_42661,N_34001,N_35036);
nor U42662 (N_42662,N_33417,N_38258);
or U42663 (N_42663,N_30571,N_39435);
xnor U42664 (N_42664,N_36720,N_31360);
nand U42665 (N_42665,N_39481,N_37690);
and U42666 (N_42666,N_31964,N_31853);
nor U42667 (N_42667,N_32055,N_38464);
nand U42668 (N_42668,N_32333,N_39856);
nand U42669 (N_42669,N_30191,N_31774);
and U42670 (N_42670,N_33238,N_36547);
nor U42671 (N_42671,N_39675,N_35009);
and U42672 (N_42672,N_37707,N_38931);
xor U42673 (N_42673,N_37578,N_34191);
xor U42674 (N_42674,N_37179,N_32480);
and U42675 (N_42675,N_33849,N_39691);
xor U42676 (N_42676,N_31656,N_36992);
or U42677 (N_42677,N_33105,N_31519);
and U42678 (N_42678,N_36984,N_33565);
and U42679 (N_42679,N_32987,N_39239);
or U42680 (N_42680,N_32696,N_34636);
and U42681 (N_42681,N_30448,N_34776);
or U42682 (N_42682,N_32415,N_31545);
xor U42683 (N_42683,N_34747,N_31601);
or U42684 (N_42684,N_34416,N_36430);
nand U42685 (N_42685,N_37308,N_35257);
nor U42686 (N_42686,N_37484,N_38860);
xor U42687 (N_42687,N_39798,N_39257);
nand U42688 (N_42688,N_39158,N_34867);
or U42689 (N_42689,N_34452,N_34562);
nand U42690 (N_42690,N_33088,N_36816);
xnor U42691 (N_42691,N_35237,N_32761);
nor U42692 (N_42692,N_32384,N_31261);
nor U42693 (N_42693,N_30088,N_31122);
xnor U42694 (N_42694,N_34972,N_37098);
nand U42695 (N_42695,N_31976,N_30703);
xor U42696 (N_42696,N_38120,N_32720);
nand U42697 (N_42697,N_39994,N_37772);
nand U42698 (N_42698,N_34646,N_38456);
or U42699 (N_42699,N_35131,N_33071);
and U42700 (N_42700,N_32338,N_31033);
nor U42701 (N_42701,N_31981,N_36874);
xnor U42702 (N_42702,N_30615,N_34641);
nor U42703 (N_42703,N_38439,N_34281);
nor U42704 (N_42704,N_30163,N_30196);
xnor U42705 (N_42705,N_35793,N_32334);
nor U42706 (N_42706,N_37857,N_38364);
or U42707 (N_42707,N_34845,N_32084);
and U42708 (N_42708,N_36239,N_33480);
nor U42709 (N_42709,N_35027,N_39665);
or U42710 (N_42710,N_31274,N_39106);
nor U42711 (N_42711,N_32635,N_39853);
xor U42712 (N_42712,N_30193,N_38769);
or U42713 (N_42713,N_33528,N_36007);
nand U42714 (N_42714,N_38661,N_39622);
or U42715 (N_42715,N_34278,N_38929);
nor U42716 (N_42716,N_36181,N_30621);
or U42717 (N_42717,N_33092,N_32785);
or U42718 (N_42718,N_39164,N_32716);
nand U42719 (N_42719,N_33240,N_38623);
or U42720 (N_42720,N_30453,N_31397);
and U42721 (N_42721,N_37612,N_39817);
nor U42722 (N_42722,N_30189,N_34353);
or U42723 (N_42723,N_38816,N_34975);
or U42724 (N_42724,N_33049,N_35942);
or U42725 (N_42725,N_30024,N_34726);
nand U42726 (N_42726,N_32263,N_31700);
xor U42727 (N_42727,N_38864,N_37695);
nor U42728 (N_42728,N_37540,N_36344);
nor U42729 (N_42729,N_34586,N_33188);
or U42730 (N_42730,N_36456,N_36830);
and U42731 (N_42731,N_35083,N_39043);
nor U42732 (N_42732,N_36563,N_38192);
or U42733 (N_42733,N_32451,N_36630);
and U42734 (N_42734,N_37487,N_37969);
nand U42735 (N_42735,N_37058,N_32775);
and U42736 (N_42736,N_32207,N_30963);
or U42737 (N_42737,N_31876,N_37161);
or U42738 (N_42738,N_38825,N_30117);
nor U42739 (N_42739,N_39934,N_36994);
xor U42740 (N_42740,N_34205,N_35284);
and U42741 (N_42741,N_39224,N_30127);
and U42742 (N_42742,N_31343,N_31238);
nor U42743 (N_42743,N_32234,N_30862);
or U42744 (N_42744,N_32954,N_33838);
and U42745 (N_42745,N_35912,N_31323);
and U42746 (N_42746,N_31512,N_30305);
xor U42747 (N_42747,N_37266,N_35821);
or U42748 (N_42748,N_31956,N_35348);
and U42749 (N_42749,N_36787,N_32831);
or U42750 (N_42750,N_38619,N_37110);
nand U42751 (N_42751,N_36706,N_38282);
nor U42752 (N_42752,N_32107,N_35641);
nand U42753 (N_42753,N_34467,N_30417);
and U42754 (N_42754,N_34733,N_34287);
or U42755 (N_42755,N_39108,N_37491);
xnor U42756 (N_42756,N_32102,N_30797);
or U42757 (N_42757,N_38925,N_31899);
or U42758 (N_42758,N_33822,N_38552);
nand U42759 (N_42759,N_31990,N_34866);
nor U42760 (N_42760,N_38750,N_34910);
or U42761 (N_42761,N_35884,N_32387);
or U42762 (N_42762,N_30325,N_32533);
and U42763 (N_42763,N_30611,N_34532);
and U42764 (N_42764,N_30178,N_30466);
nand U42765 (N_42765,N_33362,N_31309);
and U42766 (N_42766,N_33102,N_31022);
nor U42767 (N_42767,N_32910,N_35232);
or U42768 (N_42768,N_35088,N_38956);
nor U42769 (N_42769,N_39647,N_38936);
nand U42770 (N_42770,N_34836,N_31597);
and U42771 (N_42771,N_30522,N_37004);
nand U42772 (N_42772,N_38036,N_34824);
nor U42773 (N_42773,N_36040,N_35390);
and U42774 (N_42774,N_35322,N_39924);
nor U42775 (N_42775,N_38892,N_31643);
nor U42776 (N_42776,N_34107,N_33275);
nor U42777 (N_42777,N_39264,N_31043);
xor U42778 (N_42778,N_37617,N_33735);
nor U42779 (N_42779,N_39486,N_33493);
xnor U42780 (N_42780,N_32090,N_35906);
nand U42781 (N_42781,N_31219,N_39978);
nor U42782 (N_42782,N_34678,N_32401);
xor U42783 (N_42783,N_34615,N_34007);
nand U42784 (N_42784,N_34956,N_39461);
or U42785 (N_42785,N_36132,N_32306);
and U42786 (N_42786,N_39087,N_39431);
and U42787 (N_42787,N_39467,N_35494);
or U42788 (N_42788,N_30285,N_34457);
or U42789 (N_42789,N_35107,N_39322);
or U42790 (N_42790,N_39854,N_30532);
and U42791 (N_42791,N_37833,N_38179);
or U42792 (N_42792,N_38204,N_34495);
xnor U42793 (N_42793,N_30767,N_37919);
xor U42794 (N_42794,N_39658,N_34578);
xnor U42795 (N_42795,N_30254,N_38968);
nor U42796 (N_42796,N_30336,N_36605);
xor U42797 (N_42797,N_34274,N_36085);
and U42798 (N_42798,N_33244,N_34188);
nand U42799 (N_42799,N_30599,N_35658);
and U42800 (N_42800,N_34202,N_35267);
and U42801 (N_42801,N_38431,N_39463);
nand U42802 (N_42802,N_39033,N_33861);
nand U42803 (N_42803,N_32250,N_38660);
or U42804 (N_42804,N_37446,N_33477);
xnor U42805 (N_42805,N_31003,N_35724);
xor U42806 (N_42806,N_37306,N_34908);
and U42807 (N_42807,N_32600,N_30819);
and U42808 (N_42808,N_31419,N_33135);
nand U42809 (N_42809,N_33730,N_32312);
nor U42810 (N_42810,N_32402,N_32764);
and U42811 (N_42811,N_38513,N_36929);
xnor U42812 (N_42812,N_37773,N_33920);
nor U42813 (N_42813,N_30708,N_37359);
nand U42814 (N_42814,N_35815,N_37113);
xnor U42815 (N_42815,N_37460,N_30548);
or U42816 (N_42816,N_39460,N_34873);
nor U42817 (N_42817,N_33593,N_35228);
xnor U42818 (N_42818,N_33396,N_35085);
or U42819 (N_42819,N_37797,N_36403);
xor U42820 (N_42820,N_35566,N_37175);
nor U42821 (N_42821,N_37357,N_36015);
xor U42822 (N_42822,N_39253,N_31810);
or U42823 (N_42823,N_31046,N_34472);
and U42824 (N_42824,N_32083,N_36697);
xor U42825 (N_42825,N_35890,N_37598);
and U42826 (N_42826,N_36948,N_37876);
nand U42827 (N_42827,N_31997,N_37265);
nand U42828 (N_42828,N_35681,N_30598);
xnor U42829 (N_42829,N_32719,N_38427);
nor U42830 (N_42830,N_39930,N_37731);
xor U42831 (N_42831,N_39504,N_35697);
nand U42832 (N_42832,N_30490,N_38516);
nand U42833 (N_42833,N_34359,N_37508);
nand U42834 (N_42834,N_30920,N_35634);
and U42835 (N_42835,N_34767,N_33370);
nand U42836 (N_42836,N_35429,N_39454);
nand U42837 (N_42837,N_39075,N_30020);
and U42838 (N_42838,N_32561,N_31623);
or U42839 (N_42839,N_32662,N_32994);
or U42840 (N_42840,N_33740,N_36643);
nand U42841 (N_42841,N_39750,N_33582);
xor U42842 (N_42842,N_32989,N_36241);
and U42843 (N_42843,N_30495,N_30265);
nor U42844 (N_42844,N_39327,N_35713);
and U42845 (N_42845,N_36236,N_31227);
nor U42846 (N_42846,N_33442,N_33506);
xnor U42847 (N_42847,N_33554,N_31260);
and U42848 (N_42848,N_35053,N_37768);
nor U42849 (N_42849,N_33247,N_36270);
and U42850 (N_42850,N_30322,N_34081);
nor U42851 (N_42851,N_39428,N_34032);
or U42852 (N_42852,N_30341,N_35447);
and U42853 (N_42853,N_35589,N_39447);
or U42854 (N_42854,N_33274,N_32034);
or U42855 (N_42855,N_32789,N_38296);
nand U42856 (N_42856,N_39310,N_36889);
or U42857 (N_42857,N_38248,N_35304);
or U42858 (N_42858,N_33890,N_35147);
or U42859 (N_42859,N_33390,N_37216);
nor U42860 (N_42860,N_35695,N_39180);
nor U42861 (N_42861,N_37512,N_35356);
xor U42862 (N_42862,N_38298,N_32666);
nand U42863 (N_42863,N_37552,N_35595);
and U42864 (N_42864,N_33363,N_39880);
xor U42865 (N_42865,N_32323,N_30300);
nand U42866 (N_42866,N_36402,N_33144);
xor U42867 (N_42867,N_35400,N_37242);
and U42868 (N_42868,N_34110,N_30082);
nor U42869 (N_42869,N_31883,N_33296);
or U42870 (N_42870,N_38710,N_33048);
nand U42871 (N_42871,N_34051,N_30360);
nor U42872 (N_42872,N_33526,N_37654);
xnor U42873 (N_42873,N_30576,N_33634);
or U42874 (N_42874,N_34986,N_39553);
and U42875 (N_42875,N_39251,N_37321);
nor U42876 (N_42876,N_35899,N_36045);
nand U42877 (N_42877,N_31041,N_32532);
nand U42878 (N_42878,N_38422,N_32741);
and U42879 (N_42879,N_39019,N_30252);
nand U42880 (N_42880,N_36699,N_31624);
xnor U42881 (N_42881,N_32673,N_34958);
or U42882 (N_42882,N_37651,N_34405);
xnor U42883 (N_42883,N_36273,N_36803);
or U42884 (N_42884,N_39839,N_36882);
or U42885 (N_42885,N_38373,N_38490);
xor U42886 (N_42886,N_39015,N_36684);
nand U42887 (N_42887,N_39539,N_33956);
nor U42888 (N_42888,N_30786,N_34880);
and U42889 (N_42889,N_37142,N_30881);
nand U42890 (N_42890,N_32477,N_36954);
and U42891 (N_42891,N_30812,N_36627);
xor U42892 (N_42892,N_35030,N_31543);
or U42893 (N_42893,N_35638,N_30553);
and U42894 (N_42894,N_39260,N_38698);
or U42895 (N_42895,N_37416,N_31146);
nand U42896 (N_42896,N_32210,N_30187);
nand U42897 (N_42897,N_38723,N_37766);
xor U42898 (N_42898,N_35665,N_37854);
nor U42899 (N_42899,N_31457,N_39747);
and U42900 (N_42900,N_30200,N_39954);
and U42901 (N_42901,N_33993,N_39259);
nand U42902 (N_42902,N_38666,N_34293);
nand U42903 (N_42903,N_37715,N_36292);
and U42904 (N_42904,N_31737,N_31503);
nand U42905 (N_42905,N_34960,N_33682);
or U42906 (N_42906,N_33832,N_31123);
or U42907 (N_42907,N_35974,N_30848);
nand U42908 (N_42908,N_35803,N_35044);
nand U42909 (N_42909,N_36471,N_39418);
and U42910 (N_42910,N_33459,N_38551);
xor U42911 (N_42911,N_30633,N_31771);
nor U42912 (N_42912,N_36878,N_36613);
or U42913 (N_42913,N_38998,N_38820);
nor U42914 (N_42914,N_36642,N_39985);
and U42915 (N_42915,N_34792,N_39656);
nand U42916 (N_42916,N_37522,N_32052);
nand U42917 (N_42917,N_39410,N_35951);
nand U42918 (N_42918,N_30005,N_30376);
or U42919 (N_42919,N_31721,N_37097);
and U42920 (N_42920,N_35061,N_33356);
xnor U42921 (N_42921,N_39967,N_34962);
xnor U42922 (N_42922,N_33057,N_32913);
nand U42923 (N_42923,N_33329,N_39272);
nand U42924 (N_42924,N_35438,N_36432);
xnor U42925 (N_42925,N_39156,N_38632);
and U42926 (N_42926,N_35161,N_30222);
and U42927 (N_42927,N_37841,N_33823);
xor U42928 (N_42928,N_34119,N_39778);
and U42929 (N_42929,N_35215,N_32522);
nor U42930 (N_42930,N_36130,N_32440);
xor U42931 (N_42931,N_39940,N_37244);
nor U42932 (N_42932,N_31170,N_36238);
xnor U42933 (N_42933,N_34236,N_37152);
nor U42934 (N_42934,N_38172,N_34254);
nor U42935 (N_42935,N_38086,N_31133);
and U42936 (N_42936,N_35654,N_31662);
and U42937 (N_42937,N_30202,N_38572);
nand U42938 (N_42938,N_38255,N_39677);
xor U42939 (N_42939,N_39439,N_38667);
and U42940 (N_42940,N_39508,N_36639);
xor U42941 (N_42941,N_33282,N_39292);
nand U42942 (N_42942,N_32157,N_33043);
nand U42943 (N_42943,N_36693,N_33910);
or U42944 (N_42944,N_31801,N_38749);
or U42945 (N_42945,N_35971,N_33948);
or U42946 (N_42946,N_30075,N_36182);
nor U42947 (N_42947,N_39962,N_32171);
xor U42948 (N_42948,N_32017,N_33276);
or U42949 (N_42949,N_35458,N_33980);
xor U42950 (N_42950,N_33271,N_35931);
or U42951 (N_42951,N_30546,N_31108);
nand U42952 (N_42952,N_32922,N_38134);
xnor U42953 (N_42953,N_38618,N_36391);
and U42954 (N_42954,N_37518,N_31321);
or U42955 (N_42955,N_35953,N_35223);
or U42956 (N_42956,N_32128,N_31808);
nand U42957 (N_42957,N_37050,N_32853);
xor U42958 (N_42958,N_38021,N_39316);
or U42959 (N_42959,N_38460,N_30112);
xor U42960 (N_42960,N_38722,N_39050);
xnor U42961 (N_42961,N_38834,N_38198);
and U42962 (N_42962,N_33579,N_30044);
or U42963 (N_42963,N_39657,N_37276);
and U42964 (N_42964,N_36310,N_34993);
or U42965 (N_42965,N_34738,N_30138);
nand U42966 (N_42966,N_37671,N_35731);
xor U42967 (N_42967,N_30736,N_33723);
or U42968 (N_42968,N_32624,N_34348);
xor U42969 (N_42969,N_37249,N_38167);
nor U42970 (N_42970,N_33901,N_39640);
nor U42971 (N_42971,N_30518,N_33281);
xor U42972 (N_42972,N_33029,N_38260);
nand U42973 (N_42973,N_34620,N_35412);
xor U42974 (N_42974,N_39756,N_31064);
xnor U42975 (N_42975,N_36565,N_37457);
nor U42976 (N_42976,N_39890,N_38952);
nor U42977 (N_42977,N_37670,N_39619);
and U42978 (N_42978,N_38233,N_30393);
or U42979 (N_42979,N_31968,N_32986);
and U42980 (N_42980,N_33213,N_37128);
xnor U42981 (N_42981,N_37748,N_34582);
and U42982 (N_42982,N_37562,N_31032);
nor U42983 (N_42983,N_30487,N_34511);
nor U42984 (N_42984,N_34382,N_34271);
or U42985 (N_42985,N_33785,N_35770);
or U42986 (N_42986,N_37869,N_30481);
and U42987 (N_42987,N_35328,N_36153);
and U42988 (N_42988,N_36660,N_30310);
nor U42989 (N_42989,N_36113,N_31175);
and U42990 (N_42990,N_35719,N_35613);
xnor U42991 (N_42991,N_31356,N_32988);
and U42992 (N_42992,N_33007,N_35967);
and U42993 (N_42993,N_33204,N_31719);
nor U42994 (N_42994,N_38570,N_30179);
or U42995 (N_42995,N_30607,N_31725);
nand U42996 (N_42996,N_30588,N_38069);
and U42997 (N_42997,N_39822,N_37410);
and U42998 (N_42998,N_35569,N_35124);
or U42999 (N_42999,N_33550,N_36778);
nor U43000 (N_43000,N_37924,N_38164);
nand U43001 (N_43001,N_38313,N_37088);
nor U43002 (N_43002,N_33246,N_39913);
and U43003 (N_43003,N_34631,N_35523);
nand U43004 (N_43004,N_36924,N_36664);
and U43005 (N_43005,N_36915,N_36806);
and U43006 (N_43006,N_34884,N_31067);
nor U43007 (N_43007,N_31575,N_31921);
nor U43008 (N_43008,N_37849,N_32689);
xnor U43009 (N_43009,N_34540,N_32872);
nand U43010 (N_43010,N_33945,N_32892);
or U43011 (N_43011,N_33437,N_38986);
nor U43012 (N_43012,N_35853,N_36828);
or U43013 (N_43013,N_30937,N_32572);
xor U43014 (N_43014,N_32479,N_37045);
nor U43015 (N_43015,N_35240,N_38367);
and U43016 (N_43016,N_36865,N_31333);
nor U43017 (N_43017,N_34855,N_34196);
nor U43018 (N_43018,N_31421,N_33575);
xor U43019 (N_43019,N_39592,N_33709);
nor U43020 (N_43020,N_32997,N_33486);
nand U43021 (N_43021,N_32300,N_35279);
nor U43022 (N_43022,N_38626,N_37997);
nor U43023 (N_43023,N_34036,N_39755);
nor U43024 (N_43024,N_30683,N_31626);
xor U43025 (N_43025,N_32138,N_38918);
nand U43026 (N_43026,N_37502,N_31858);
or U43027 (N_43027,N_38697,N_37222);
and U43028 (N_43028,N_30641,N_30775);
xnor U43029 (N_43029,N_37283,N_30055);
xnor U43030 (N_43030,N_35342,N_34712);
xor U43031 (N_43031,N_31125,N_35141);
nor U43032 (N_43032,N_36545,N_34343);
xnor U43033 (N_43033,N_37170,N_30707);
or U43034 (N_43034,N_39117,N_30540);
nor U43035 (N_43035,N_33584,N_36354);
or U43036 (N_43036,N_34190,N_32238);
nand U43037 (N_43037,N_30829,N_35062);
and U43038 (N_43038,N_38532,N_35757);
and U43039 (N_43039,N_30415,N_37546);
nor U43040 (N_43040,N_36541,N_31566);
nor U43041 (N_43041,N_33308,N_32218);
xor U43042 (N_43042,N_33438,N_35616);
and U43043 (N_43043,N_37741,N_30679);
and U43044 (N_43044,N_30148,N_36110);
and U43045 (N_43045,N_30438,N_39372);
nor U43046 (N_43046,N_38369,N_30046);
nor U43047 (N_43047,N_33346,N_37955);
and U43048 (N_43048,N_31765,N_34556);
nor U43049 (N_43049,N_34927,N_35820);
nand U43050 (N_43050,N_39465,N_36233);
nor U43051 (N_43051,N_31029,N_37172);
xnor U43052 (N_43052,N_34520,N_30805);
xnor U43053 (N_43053,N_31406,N_31862);
or U43054 (N_43054,N_36868,N_31869);
xnor U43055 (N_43055,N_31451,N_36912);
or U43056 (N_43056,N_39785,N_39193);
nand U43057 (N_43057,N_30790,N_34829);
nor U43058 (N_43058,N_33722,N_39736);
nor U43059 (N_43059,N_33128,N_33922);
and U43060 (N_43060,N_32778,N_31919);
xnor U43061 (N_43061,N_32041,N_35170);
nor U43062 (N_43062,N_31526,N_34269);
xnor U43063 (N_43063,N_32813,N_36020);
nand U43064 (N_43064,N_30863,N_35994);
xor U43065 (N_43065,N_32992,N_35493);
xor U43066 (N_43066,N_34839,N_39185);
nand U43067 (N_43067,N_33454,N_31335);
and U43068 (N_43068,N_30188,N_39779);
or U43069 (N_43069,N_36221,N_37461);
or U43070 (N_43070,N_33507,N_33313);
nand U43071 (N_43071,N_38444,N_33623);
xnor U43072 (N_43072,N_30976,N_30247);
nand U43073 (N_43073,N_36423,N_38343);
nor U43074 (N_43074,N_30105,N_39225);
nand U43075 (N_43075,N_39163,N_37975);
and U43076 (N_43076,N_36444,N_32637);
and U43077 (N_43077,N_36305,N_32132);
and U43078 (N_43078,N_30258,N_35192);
or U43079 (N_43079,N_33686,N_37076);
and U43080 (N_43080,N_36529,N_32013);
xor U43081 (N_43081,N_37395,N_39983);
and U43082 (N_43082,N_38230,N_37569);
and U43083 (N_43083,N_36359,N_31807);
nor U43084 (N_43084,N_34497,N_33691);
or U43085 (N_43085,N_36633,N_35854);
xor U43086 (N_43086,N_38281,N_30404);
or U43087 (N_43087,N_30245,N_31767);
xor U43088 (N_43088,N_38670,N_37181);
xor U43089 (N_43089,N_31747,N_30995);
nor U43090 (N_43090,N_33898,N_35862);
and U43091 (N_43091,N_35651,N_36951);
and U43092 (N_43092,N_32509,N_33708);
xor U43093 (N_43093,N_38190,N_38629);
xor U43094 (N_43094,N_32603,N_33287);
xnor U43095 (N_43095,N_38478,N_37618);
and U43096 (N_43096,N_35894,N_30375);
nor U43097 (N_43097,N_30017,N_35954);
nor U43098 (N_43098,N_35219,N_36724);
or U43099 (N_43099,N_30626,N_34661);
nor U43100 (N_43100,N_31306,N_39748);
nor U43101 (N_43101,N_30701,N_36562);
or U43102 (N_43102,N_38959,N_32616);
xor U43103 (N_43103,N_32742,N_37506);
xor U43104 (N_43104,N_31877,N_34376);
xnor U43105 (N_43105,N_30104,N_31367);
nor U43106 (N_43106,N_34177,N_34404);
xnor U43107 (N_43107,N_31430,N_39053);
and U43108 (N_43108,N_36170,N_33602);
or U43109 (N_43109,N_38228,N_39813);
or U43110 (N_43110,N_35579,N_33338);
or U43111 (N_43111,N_36338,N_39207);
and U43112 (N_43112,N_30742,N_33249);
or U43113 (N_43113,N_36637,N_31266);
nor U43114 (N_43114,N_35543,N_38428);
nor U43115 (N_43115,N_36512,N_31511);
xor U43116 (N_43116,N_33741,N_38419);
xnor U43117 (N_43117,N_35824,N_30735);
or U43118 (N_43118,N_32507,N_30479);
nand U43119 (N_43119,N_30061,N_30610);
nor U43120 (N_43120,N_38942,N_39538);
or U43121 (N_43121,N_32213,N_31904);
xnor U43122 (N_43122,N_32492,N_39283);
xor U43123 (N_43123,N_30402,N_38193);
and U43124 (N_43124,N_30710,N_34455);
or U43125 (N_43125,N_36368,N_34905);
nand U43126 (N_43126,N_36373,N_34372);
nand U43127 (N_43127,N_32376,N_35418);
nand U43128 (N_43128,N_31674,N_34939);
nand U43129 (N_43129,N_39198,N_38136);
xor U43130 (N_43130,N_30446,N_34591);
nor U43131 (N_43131,N_32867,N_35073);
and U43132 (N_43132,N_30557,N_34705);
and U43133 (N_43133,N_36551,N_36462);
nor U43134 (N_43134,N_32818,N_32105);
and U43135 (N_43135,N_34093,N_36474);
xnor U43136 (N_43136,N_31461,N_39150);
xnor U43137 (N_43137,N_39950,N_34891);
xor U43138 (N_43138,N_31042,N_38079);
nor U43139 (N_43139,N_37894,N_30039);
and U43140 (N_43140,N_38505,N_34915);
xnor U43141 (N_43141,N_37968,N_36164);
xnor U43142 (N_43142,N_32058,N_39679);
nand U43143 (N_43143,N_37783,N_35491);
nand U43144 (N_43144,N_38445,N_39250);
and U43145 (N_43145,N_34608,N_36002);
nand U43146 (N_43146,N_34257,N_37174);
nor U43147 (N_43147,N_36127,N_31488);
or U43148 (N_43148,N_35262,N_30352);
and U43149 (N_43149,N_39052,N_38170);
and U43150 (N_43150,N_31854,N_37604);
nor U43151 (N_43151,N_38564,N_39938);
or U43152 (N_43152,N_38808,N_32564);
nor U43153 (N_43153,N_36042,N_38709);
or U43154 (N_43154,N_33753,N_33118);
nand U43155 (N_43155,N_39462,N_32874);
nor U43156 (N_43156,N_34973,N_36161);
xnor U43157 (N_43157,N_33781,N_39981);
and U43158 (N_43158,N_32674,N_31612);
nor U43159 (N_43159,N_35873,N_30493);
xnor U43160 (N_43160,N_37594,N_35012);
nand U43161 (N_43161,N_37237,N_34240);
nand U43162 (N_43162,N_32730,N_38576);
xor U43163 (N_43163,N_33234,N_32405);
nand U43164 (N_43164,N_35557,N_36836);
xor U43165 (N_43165,N_36674,N_30280);
xnor U43166 (N_43166,N_34059,N_39568);
xnor U43167 (N_43167,N_35066,N_32048);
xor U43168 (N_43168,N_32170,N_37247);
nand U43169 (N_43169,N_36209,N_36137);
or U43170 (N_43170,N_36163,N_38148);
nand U43171 (N_43171,N_31605,N_30971);
nor U43172 (N_43172,N_35823,N_30688);
nor U43173 (N_43173,N_38266,N_36117);
nor U43174 (N_43174,N_33694,N_33540);
nand U43175 (N_43175,N_36327,N_32475);
nand U43176 (N_43176,N_35441,N_37365);
nand U43177 (N_43177,N_37471,N_31729);
nor U43178 (N_43178,N_39475,N_36420);
xor U43179 (N_43179,N_39493,N_31237);
or U43180 (N_43180,N_37483,N_38822);
nand U43181 (N_43181,N_39520,N_35886);
xnor U43182 (N_43182,N_36425,N_39624);
or U43183 (N_43183,N_37271,N_35833);
nand U43184 (N_43184,N_38824,N_37015);
or U43185 (N_43185,N_31651,N_30413);
xnor U43186 (N_43186,N_35838,N_35155);
nor U43187 (N_43187,N_37354,N_39845);
nand U43188 (N_43188,N_35916,N_30126);
xor U43189 (N_43189,N_33716,N_35090);
nand U43190 (N_43190,N_39430,N_35965);
nand U43191 (N_43191,N_39543,N_34863);
and U43192 (N_43192,N_31346,N_39100);
xor U43193 (N_43193,N_32076,N_31998);
nand U43194 (N_43194,N_35831,N_34744);
xnor U43195 (N_43195,N_33126,N_39373);
nor U43196 (N_43196,N_37864,N_33475);
nand U43197 (N_43197,N_38917,N_30355);
nor U43198 (N_43198,N_31776,N_32342);
and U43199 (N_43199,N_37066,N_38841);
xor U43200 (N_43200,N_34786,N_33349);
or U43201 (N_43201,N_33719,N_30029);
xor U43202 (N_43202,N_37544,N_36985);
nor U43203 (N_43203,N_38605,N_31302);
nand U43204 (N_43204,N_38579,N_31582);
nand U43205 (N_43205,N_34448,N_34525);
nor U43206 (N_43206,N_36166,N_34561);
nor U43207 (N_43207,N_31759,N_33378);
and U43208 (N_43208,N_31929,N_31591);
nand U43209 (N_43209,N_37650,N_36342);
nand U43210 (N_43210,N_35310,N_32701);
xnor U43211 (N_43211,N_35626,N_35496);
nor U43212 (N_43212,N_37368,N_33411);
and U43213 (N_43213,N_39478,N_31140);
nor U43214 (N_43214,N_38455,N_38350);
or U43215 (N_43215,N_39595,N_38544);
nor U43216 (N_43216,N_36337,N_36764);
and U43217 (N_43217,N_36918,N_36973);
xnor U43218 (N_43218,N_31530,N_36219);
nand U43219 (N_43219,N_35096,N_31427);
or U43220 (N_43220,N_35711,N_31581);
and U43221 (N_43221,N_31631,N_31171);
nand U43222 (N_43222,N_31875,N_32805);
and U43223 (N_43223,N_37279,N_37025);
or U43224 (N_43224,N_38465,N_39284);
xor U43225 (N_43225,N_30261,N_36756);
xnor U43226 (N_43226,N_35535,N_36591);
xnor U43227 (N_43227,N_38017,N_30957);
nand U43228 (N_43228,N_35315,N_36217);
and U43229 (N_43229,N_33662,N_35830);
or U43230 (N_43230,N_32149,N_35449);
or U43231 (N_43231,N_31971,N_33300);
xnor U43232 (N_43232,N_38468,N_30685);
and U43233 (N_43233,N_31230,N_34504);
nand U43234 (N_43234,N_36196,N_34120);
and U43235 (N_43235,N_30860,N_32184);
and U43236 (N_43236,N_34969,N_38304);
xnor U43237 (N_43237,N_38791,N_34533);
nor U43238 (N_43238,N_35462,N_35866);
xor U43239 (N_43239,N_36495,N_33019);
nor U43240 (N_43240,N_30236,N_33245);
and U43241 (N_43241,N_34529,N_39319);
or U43242 (N_43242,N_36089,N_32644);
and U43243 (N_43243,N_32059,N_31892);
nand U43244 (N_43244,N_33319,N_37485);
nand U43245 (N_43245,N_36026,N_32529);
nand U43246 (N_43246,N_36922,N_37717);
nand U43247 (N_43247,N_32098,N_34971);
xnor U43248 (N_43248,N_30605,N_38123);
nand U43249 (N_43249,N_37073,N_30288);
and U43250 (N_43250,N_34671,N_39409);
nor U43251 (N_43251,N_30838,N_30899);
nor U43252 (N_43252,N_36141,N_34400);
xnor U43253 (N_43253,N_33142,N_33534);
and U43254 (N_43254,N_36478,N_38416);
nor U43255 (N_43255,N_37572,N_31991);
or U43256 (N_43256,N_37756,N_36298);
or U43257 (N_43257,N_38279,N_39631);
xnor U43258 (N_43258,N_36549,N_32474);
and U43259 (N_43259,N_35160,N_34758);
nand U43260 (N_43260,N_36628,N_37458);
or U43261 (N_43261,N_33366,N_32148);
nor U43262 (N_43262,N_39051,N_30398);
xnor U43263 (N_43263,N_32137,N_32908);
and U43264 (N_43264,N_35295,N_32638);
and U43265 (N_43265,N_30552,N_34946);
and U43266 (N_43266,N_35596,N_35748);
nand U43267 (N_43267,N_36328,N_30617);
nand U43268 (N_43268,N_33052,N_34509);
or U43269 (N_43269,N_37202,N_35961);
nor U43270 (N_43270,N_36970,N_36790);
or U43271 (N_43271,N_30383,N_39510);
xnor U43272 (N_43272,N_38922,N_35373);
nor U43273 (N_43273,N_33860,N_33074);
nand U43274 (N_43274,N_30508,N_32743);
xnor U43275 (N_43275,N_37022,N_34929);
nor U43276 (N_43276,N_30298,N_39038);
or U43277 (N_43277,N_34790,N_36599);
xor U43278 (N_43278,N_32441,N_33056);
nor U43279 (N_43279,N_33333,N_39293);
nor U43280 (N_43280,N_30857,N_37703);
xor U43281 (N_43281,N_38908,N_31090);
xnor U43282 (N_43282,N_37751,N_34280);
and U43283 (N_43283,N_35177,N_30778);
xor U43284 (N_43284,N_32293,N_30433);
nand U43285 (N_43285,N_32166,N_30269);
and U43286 (N_43286,N_35949,N_33863);
and U43287 (N_43287,N_32977,N_38893);
xor U43288 (N_43288,N_39549,N_38324);
xnor U43289 (N_43289,N_31551,N_34135);
and U43290 (N_43290,N_31692,N_31147);
xor U43291 (N_43291,N_38567,N_38515);
nor U43292 (N_43292,N_32829,N_34223);
xnor U43293 (N_43293,N_30658,N_37870);
xnor U43294 (N_43294,N_39991,N_35268);
nor U43295 (N_43295,N_38355,N_36800);
nand U43296 (N_43296,N_36998,N_36047);
nor U43297 (N_43297,N_37711,N_33568);
nor U43298 (N_43298,N_31148,N_33068);
and U43299 (N_43299,N_30680,N_33212);
xnor U43300 (N_43300,N_33598,N_32755);
and U43301 (N_43301,N_30614,N_35354);
nand U43302 (N_43302,N_32243,N_39291);
nand U43303 (N_43303,N_38450,N_36063);
nand U43304 (N_43304,N_36950,N_38604);
xnor U43305 (N_43305,N_33586,N_36741);
nor U43306 (N_43306,N_39165,N_31570);
and U43307 (N_43307,N_31393,N_38717);
nor U43308 (N_43308,N_31502,N_38011);
nand U43309 (N_43309,N_30094,N_35568);
or U43310 (N_43310,N_39760,N_39364);
xnor U43311 (N_43311,N_38996,N_37677);
xnor U43312 (N_43312,N_33853,N_32735);
or U43313 (N_43313,N_33982,N_36694);
nor U43314 (N_43314,N_35499,N_37830);
or U43315 (N_43315,N_36242,N_39581);
nand U43316 (N_43316,N_34043,N_39692);
and U43317 (N_43317,N_31741,N_31934);
nand U43318 (N_43318,N_38699,N_35052);
nor U43319 (N_43319,N_34444,N_34761);
or U43320 (N_43320,N_38910,N_30706);
nor U43321 (N_43321,N_30111,N_34598);
and U43322 (N_43322,N_34762,N_37644);
nand U43323 (N_43323,N_31549,N_33222);
nand U43324 (N_43324,N_33488,N_36531);
or U43325 (N_43325,N_35371,N_30461);
nor U43326 (N_43326,N_30733,N_34739);
and U43327 (N_43327,N_37667,N_37978);
nand U43328 (N_43328,N_33223,N_38414);
nor U43329 (N_43329,N_37792,N_32575);
nand U43330 (N_43330,N_36383,N_32863);
nand U43331 (N_43331,N_30230,N_31603);
xor U43332 (N_43332,N_34757,N_35832);
and U43333 (N_43333,N_37800,N_34449);
or U43334 (N_43334,N_34270,N_37217);
and U43335 (N_43335,N_38314,N_32371);
and U43336 (N_43336,N_31641,N_39753);
xnor U43337 (N_43337,N_30616,N_35366);
and U43338 (N_43338,N_37779,N_36450);
and U43339 (N_43339,N_34092,N_31766);
or U43340 (N_43340,N_34823,N_33658);
nand U43341 (N_43341,N_32688,N_39459);
or U43342 (N_43342,N_30667,N_32508);
or U43343 (N_43343,N_34479,N_37996);
or U43344 (N_43344,N_39318,N_36626);
and U43345 (N_43345,N_37385,N_34966);
nor U43346 (N_43346,N_38065,N_32276);
nor U43347 (N_43347,N_35527,N_38601);
nor U43348 (N_43348,N_37759,N_37269);
nor U43349 (N_43349,N_31730,N_30510);
and U43350 (N_43350,N_34057,N_36677);
nor U43351 (N_43351,N_30335,N_37963);
and U43352 (N_43352,N_36018,N_33940);
nor U43353 (N_43353,N_37846,N_34947);
nor U43354 (N_43354,N_35666,N_35718);
xnor U43355 (N_43355,N_33989,N_32521);
nor U43356 (N_43356,N_33907,N_39646);
xnor U43357 (N_43357,N_35382,N_35676);
and U43358 (N_43358,N_39960,N_33888);
nor U43359 (N_43359,N_32418,N_31359);
nor U43360 (N_43360,N_37904,N_30551);
and U43361 (N_43361,N_32241,N_37951);
and U43362 (N_43362,N_36334,N_38482);
nor U43363 (N_43363,N_38746,N_39898);
or U43364 (N_43364,N_39442,N_35486);
or U43365 (N_43365,N_37949,N_35435);
nand U43366 (N_43366,N_39588,N_39689);
and U43367 (N_43367,N_35245,N_32427);
or U43368 (N_43368,N_35892,N_34345);
and U43369 (N_43369,N_38146,N_39857);
xnor U43370 (N_43370,N_34352,N_33630);
nand U43371 (N_43371,N_37504,N_36526);
or U43372 (N_43372,N_32316,N_31541);
xnor U43373 (N_43373,N_33923,N_37652);
nor U43374 (N_43374,N_34882,N_38119);
nand U43375 (N_43375,N_31453,N_33291);
and U43376 (N_43376,N_37465,N_31128);
or U43377 (N_43377,N_37663,N_38110);
xor U43378 (N_43378,N_33844,N_36319);
xor U43379 (N_43379,N_31249,N_35561);
and U43380 (N_43380,N_39200,N_31001);
nor U43381 (N_43381,N_39571,N_36169);
xnor U43382 (N_43382,N_38108,N_37016);
or U43383 (N_43383,N_37375,N_32012);
xor U43384 (N_43384,N_34694,N_38180);
xor U43385 (N_43385,N_35647,N_38039);
nand U43386 (N_43386,N_37698,N_39328);
nor U43387 (N_43387,N_34795,N_36005);
and U43388 (N_43388,N_34314,N_31764);
or U43389 (N_43389,N_31884,N_37093);
xnor U43390 (N_43390,N_31983,N_36935);
nand U43391 (N_43391,N_37844,N_38325);
xor U43392 (N_43392,N_39074,N_38406);
nor U43393 (N_43393,N_31942,N_31937);
xor U43394 (N_43394,N_38573,N_33155);
nand U43395 (N_43395,N_34260,N_39635);
xnor U43396 (N_43396,N_32912,N_32858);
nor U43397 (N_43397,N_30656,N_38376);
or U43398 (N_43398,N_32009,N_30519);
xnor U43399 (N_43399,N_30019,N_37683);
and U43400 (N_43400,N_33679,N_32286);
xor U43401 (N_43401,N_30842,N_37752);
nand U43402 (N_43402,N_34778,N_33895);
or U43403 (N_43403,N_31913,N_32165);
or U43404 (N_43404,N_32093,N_36147);
xnor U43405 (N_43405,N_35051,N_37665);
nand U43406 (N_43406,N_31245,N_39266);
xnor U43407 (N_43407,N_37021,N_33935);
nand U43408 (N_43408,N_35720,N_33557);
and U43409 (N_43409,N_35125,N_31137);
or U43410 (N_43410,N_30747,N_34861);
and U43411 (N_43411,N_31190,N_30093);
xor U43412 (N_43412,N_32176,N_32758);
nor U43413 (N_43413,N_38798,N_34941);
xnor U43414 (N_43414,N_39770,N_30887);
and U43415 (N_43415,N_30604,N_36098);
or U43416 (N_43416,N_31654,N_32959);
nand U43417 (N_43417,N_39625,N_31006);
xor U43418 (N_43418,N_30083,N_32406);
xnor U43419 (N_43419,N_35791,N_36974);
nand U43420 (N_43420,N_30560,N_33062);
xnor U43421 (N_43421,N_30231,N_37182);
nor U43422 (N_43422,N_32200,N_35422);
nor U43423 (N_43423,N_34470,N_33131);
nand U43424 (N_43424,N_36109,N_37729);
xnor U43425 (N_43425,N_33355,N_36789);
nor U43426 (N_43426,N_39438,N_36376);
and U43427 (N_43427,N_31746,N_33881);
xor U43428 (N_43428,N_38652,N_38235);
and U43429 (N_43429,N_31646,N_34576);
xnor U43430 (N_43430,N_39256,N_30037);
nor U43431 (N_43431,N_37934,N_32788);
xnor U43432 (N_43432,N_30955,N_39186);
and U43433 (N_43433,N_33138,N_31217);
or U43434 (N_43434,N_32188,N_38402);
xor U43435 (N_43435,N_30014,N_39810);
nand U43436 (N_43436,N_31772,N_37600);
or U43437 (N_43437,N_32598,N_38184);
nand U43438 (N_43438,N_35716,N_33761);
or U43439 (N_43439,N_31083,N_32905);
or U43440 (N_43440,N_39485,N_32006);
xnor U43441 (N_43441,N_33972,N_32851);
nand U43442 (N_43442,N_32531,N_35781);
xor U43443 (N_43443,N_30066,N_31253);
or U43444 (N_43444,N_31278,N_39445);
nand U43445 (N_43445,N_39081,N_39088);
xor U43446 (N_43446,N_30204,N_30972);
nand U43447 (N_43447,N_39258,N_33318);
xnor U43448 (N_43448,N_33386,N_37287);
or U43449 (N_43449,N_39362,N_34594);
nor U43450 (N_43450,N_37674,N_36829);
nand U43451 (N_43451,N_38451,N_35817);
nand U43452 (N_43452,N_30226,N_35526);
and U43453 (N_43453,N_31057,N_38663);
or U43454 (N_43454,N_34901,N_34362);
xor U43455 (N_43455,N_33751,N_31361);
xor U43456 (N_43456,N_32357,N_35959);
nor U43457 (N_43457,N_30337,N_37545);
or U43458 (N_43458,N_30521,N_32650);
nor U43459 (N_43459,N_32467,N_31426);
xor U43460 (N_43460,N_36617,N_32422);
and U43461 (N_43461,N_34607,N_39688);
and U43462 (N_43462,N_30284,N_30214);
nand U43463 (N_43463,N_38641,N_33697);
nor U43464 (N_43464,N_34237,N_39721);
and U43465 (N_43465,N_33086,N_31144);
and U43466 (N_43466,N_37992,N_30539);
xnor U43467 (N_43467,N_39556,N_30270);
and U43468 (N_43468,N_30846,N_30725);
or U43469 (N_43469,N_37583,N_37433);
xnor U43470 (N_43470,N_39012,N_35475);
nand U43471 (N_43471,N_30872,N_30696);
and U43472 (N_43472,N_31472,N_39144);
and U43473 (N_43473,N_31564,N_30457);
nand U43474 (N_43474,N_34326,N_35502);
and U43475 (N_43475,N_39926,N_37067);
nand U43476 (N_43476,N_38979,N_37528);
or U43477 (N_43477,N_35440,N_37774);
or U43478 (N_43478,N_34426,N_31706);
nand U43479 (N_43479,N_39738,N_32258);
and U43480 (N_43480,N_31977,N_39006);
or U43481 (N_43481,N_38374,N_35169);
nand U43482 (N_43482,N_33137,N_32247);
and U43483 (N_43483,N_35309,N_36072);
and U43484 (N_43484,N_32585,N_33248);
nand U43485 (N_43485,N_35166,N_34526);
or U43486 (N_43486,N_39265,N_36710);
nand U43487 (N_43487,N_38410,N_36027);
nor U43488 (N_43488,N_33205,N_30509);
nor U43489 (N_43489,N_38842,N_36422);
xor U43490 (N_43490,N_36300,N_32496);
and U43491 (N_43491,N_30851,N_36413);
nor U43492 (N_43492,N_35903,N_32340);
nand U43493 (N_43493,N_32645,N_38702);
nand U43494 (N_43494,N_31314,N_38449);
and U43495 (N_43495,N_35379,N_34255);
nor U43496 (N_43496,N_39993,N_38426);
nor U43497 (N_43497,N_35741,N_31975);
or U43498 (N_43498,N_34630,N_31182);
nand U43499 (N_43499,N_30411,N_32019);
nor U43500 (N_43500,N_34252,N_35625);
nor U43501 (N_43501,N_35775,N_38016);
xnor U43502 (N_43502,N_39823,N_39474);
and U43503 (N_43503,N_37762,N_37890);
nor U43504 (N_43504,N_39815,N_36489);
or U43505 (N_43505,N_34567,N_39746);
nand U43506 (N_43506,N_39214,N_35079);
and U43507 (N_43507,N_35828,N_36533);
or U43508 (N_43508,N_33795,N_38215);
nor U43509 (N_43509,N_34090,N_35755);
nand U43510 (N_43510,N_37880,N_38238);
and U43511 (N_43511,N_32030,N_33748);
and U43512 (N_43512,N_33393,N_39579);
and U43513 (N_43513,N_38046,N_33399);
xor U43514 (N_43514,N_32621,N_39704);
and U43515 (N_43515,N_31324,N_30833);
nor U43516 (N_43516,N_33924,N_32583);
or U43517 (N_43517,N_35752,N_34787);
nor U43518 (N_43518,N_39602,N_33990);
xor U43519 (N_43519,N_37565,N_34302);
nand U43520 (N_43520,N_34106,N_32978);
nor U43521 (N_43521,N_35006,N_30525);
xor U43522 (N_43522,N_31290,N_33197);
and U43523 (N_43523,N_32786,N_30334);
xor U43524 (N_43524,N_38125,N_34285);
and U43525 (N_43525,N_33892,N_31748);
or U43526 (N_43526,N_32127,N_34330);
nand U43527 (N_43527,N_37906,N_38163);
nor U43528 (N_43528,N_34336,N_39560);
xnor U43529 (N_43529,N_30423,N_38452);
xnor U43530 (N_43530,N_39866,N_31017);
and U43531 (N_43531,N_36249,N_38088);
or U43532 (N_43532,N_39079,N_34045);
nor U43533 (N_43533,N_38964,N_32037);
and U43534 (N_43534,N_39441,N_32112);
nand U43535 (N_43535,N_38483,N_36832);
nor U43536 (N_43536,N_34988,N_38071);
and U43537 (N_43537,N_31136,N_34473);
nand U43538 (N_43538,N_31600,N_37432);
nor U43539 (N_43539,N_37952,N_34248);
and U43540 (N_43540,N_34217,N_37570);
nand U43541 (N_43541,N_37816,N_37300);
or U43542 (N_43542,N_38790,N_36760);
xor U43543 (N_43543,N_37709,N_34687);
nor U43544 (N_43544,N_33294,N_31985);
nor U43545 (N_43545,N_32129,N_36277);
or U43546 (N_43546,N_37619,N_35767);
nand U43547 (N_43547,N_33846,N_36256);
and U43548 (N_43548,N_36096,N_39862);
and U43549 (N_43549,N_38764,N_37788);
or U43550 (N_43550,N_31596,N_38571);
or U43551 (N_43551,N_39457,N_32167);
nand U43552 (N_43552,N_32779,N_32181);
xor U43553 (N_43553,N_38289,N_35436);
nor U43554 (N_43554,N_32449,N_31949);
and U43555 (N_43555,N_35248,N_30349);
nor U43556 (N_43556,N_31499,N_39783);
nand U43557 (N_43557,N_36028,N_37932);
xor U43558 (N_43558,N_34290,N_38866);
or U43559 (N_43559,N_39524,N_35708);
nor U43560 (N_43560,N_35407,N_34313);
or U43561 (N_43561,N_32133,N_35733);
xor U43562 (N_43562,N_36536,N_39548);
or U43563 (N_43563,N_39391,N_30934);
nand U43564 (N_43564,N_34077,N_34501);
or U43565 (N_43565,N_35275,N_38978);
and U43566 (N_43566,N_39683,N_30960);
or U43567 (N_43567,N_30181,N_31650);
nand U43568 (N_43568,N_31864,N_33525);
nor U43569 (N_43569,N_38005,N_30891);
or U43570 (N_43570,N_33039,N_39190);
xor U43571 (N_43571,N_32586,N_33703);
and U43572 (N_43572,N_37521,N_35592);
nand U43573 (N_43573,N_32411,N_36612);
xnor U43574 (N_43574,N_34201,N_31336);
and U43575 (N_43575,N_38206,N_35944);
nor U43576 (N_43576,N_39768,N_34369);
or U43577 (N_43577,N_35580,N_30249);
xnor U43578 (N_43578,N_37087,N_38961);
or U43579 (N_43579,N_35199,N_32693);
and U43580 (N_43580,N_32504,N_34440);
and U43581 (N_43581,N_35734,N_34870);
nand U43582 (N_43582,N_39021,N_35201);
and U43583 (N_43583,N_35338,N_30958);
nand U43584 (N_43584,N_32800,N_37081);
or U43585 (N_43585,N_32350,N_34446);
nand U43586 (N_43586,N_37079,N_39381);
and U43587 (N_43587,N_34158,N_30377);
and U43588 (N_43588,N_37993,N_30092);
nor U43589 (N_43589,N_30714,N_30113);
or U43590 (N_43590,N_30951,N_34111);
or U43591 (N_43591,N_30956,N_34746);
nor U43592 (N_43592,N_37135,N_32173);
and U43593 (N_43593,N_38519,N_34771);
nand U43594 (N_43594,N_30038,N_33078);
and U43595 (N_43595,N_34292,N_32631);
nand U43596 (N_43596,N_32046,N_39499);
or U43597 (N_43597,N_34837,N_35443);
or U43598 (N_43598,N_39925,N_31694);
and U43599 (N_43599,N_36168,N_33193);
nor U43600 (N_43600,N_33626,N_36218);
and U43601 (N_43601,N_37574,N_31201);
or U43602 (N_43602,N_39734,N_38280);
nor U43603 (N_43603,N_38915,N_36532);
and U43604 (N_43604,N_36539,N_39932);
and U43605 (N_43605,N_30103,N_32101);
nor U43606 (N_43606,N_39243,N_31273);
and U43607 (N_43607,N_32806,N_31785);
xor U43608 (N_43608,N_36467,N_32815);
nand U43609 (N_43609,N_37530,N_35367);
nor U43610 (N_43610,N_34933,N_31696);
nor U43611 (N_43611,N_34029,N_37111);
or U43612 (N_43612,N_37590,N_31920);
nor U43613 (N_43613,N_34581,N_30878);
or U43614 (N_43614,N_35556,N_38990);
nor U43615 (N_43615,N_31295,N_35347);
nor U43616 (N_43616,N_36773,N_30475);
or U43617 (N_43617,N_30636,N_37847);
nand U43618 (N_43618,N_37153,N_33905);
xor U43619 (N_43619,N_36755,N_35861);
nor U43620 (N_43620,N_37320,N_36596);
nand U43621 (N_43621,N_35410,N_34460);
and U43622 (N_43622,N_33546,N_33885);
or U43623 (N_43623,N_38270,N_34835);
nand U43624 (N_43624,N_33467,N_35893);
or U43625 (N_43625,N_35207,N_32738);
and U43626 (N_43626,N_33825,N_30590);
nor U43627 (N_43627,N_37960,N_32016);
or U43628 (N_43628,N_32962,N_32932);
or U43629 (N_43629,N_33943,N_33522);
and U43630 (N_43630,N_35743,N_31456);
nand U43631 (N_43631,N_30164,N_34203);
nand U43632 (N_43632,N_34458,N_38486);
nor U43633 (N_43633,N_39685,N_39092);
and U43634 (N_43634,N_31640,N_36431);
xor U43635 (N_43635,N_32943,N_37239);
nor U43636 (N_43636,N_38214,N_33023);
nor U43637 (N_43637,N_35850,N_30023);
xnor U43638 (N_43638,N_32094,N_39715);
xnor U43639 (N_43639,N_33458,N_37929);
and U43640 (N_43640,N_30908,N_35254);
and U43641 (N_43641,N_33104,N_34957);
or U43642 (N_43642,N_37236,N_35001);
or U43643 (N_43643,N_30586,N_39964);
nor U43644 (N_43644,N_35361,N_34380);
and U43645 (N_43645,N_33320,N_34816);
nor U43646 (N_43646,N_30327,N_33866);
nor U43647 (N_43647,N_35902,N_36822);
xnor U43648 (N_43648,N_36032,N_33302);
or U43649 (N_43649,N_31065,N_32358);
nor U43650 (N_43650,N_36105,N_36722);
xnor U43651 (N_43651,N_33429,N_32044);
or U43652 (N_43652,N_38882,N_38366);
and U43653 (N_43653,N_33343,N_36251);
and U43654 (N_43654,N_35973,N_35283);
nand U43655 (N_43655,N_31347,N_35982);
and U43656 (N_43656,N_37532,N_36488);
nand U43657 (N_43657,N_35198,N_33603);
nor U43658 (N_43658,N_32630,N_39971);
xor U43659 (N_43659,N_36142,N_30634);
xnor U43660 (N_43660,N_31548,N_34887);
nand U43661 (N_43661,N_33577,N_31755);
nand U43662 (N_43662,N_39792,N_36762);
nor U43663 (N_43663,N_39931,N_31762);
nor U43664 (N_43664,N_34466,N_32731);
and U43665 (N_43665,N_39671,N_35785);
or U43666 (N_43666,N_31215,N_36479);
xnor U43667 (N_43667,N_33729,N_37384);
and U43668 (N_43668,N_31223,N_36255);
nor U43669 (N_43669,N_36597,N_31019);
and U43670 (N_43670,N_36454,N_35524);
xnor U43671 (N_43671,N_35015,N_36510);
nor U43672 (N_43672,N_32470,N_30108);
xnor U43673 (N_43673,N_38970,N_35889);
and U43674 (N_43674,N_30785,N_34834);
and U43675 (N_43675,N_37543,N_34477);
and U43676 (N_43676,N_35013,N_30913);
xnor U43677 (N_43677,N_38928,N_32074);
nor U43678 (N_43678,N_33122,N_36726);
nor U43679 (N_43679,N_39378,N_35657);
xnor U43680 (N_43680,N_37101,N_30874);
nor U43681 (N_43681,N_30171,N_37102);
xor U43682 (N_43682,N_30331,N_30449);
nand U43683 (N_43683,N_33421,N_34782);
nand U43684 (N_43684,N_36162,N_38741);
and U43685 (N_43685,N_34437,N_32982);
xor U43686 (N_43686,N_30613,N_33615);
nor U43687 (N_43687,N_36160,N_32487);
nand U43688 (N_43688,N_32756,N_33769);
or U43689 (N_43689,N_35736,N_34601);
nor U43690 (N_43690,N_38536,N_33544);
or U43691 (N_43691,N_31836,N_34590);
and U43692 (N_43692,N_32528,N_34680);
and U43693 (N_43693,N_39308,N_35725);
nor U43694 (N_43694,N_32652,N_34879);
and U43695 (N_43695,N_36356,N_35508);
nor U43696 (N_43696,N_31413,N_32186);
or U43697 (N_43697,N_34253,N_32707);
and U43698 (N_43698,N_32877,N_33713);
nor U43699 (N_43699,N_31821,N_37812);
or U43700 (N_43700,N_39722,N_37556);
or U43701 (N_43701,N_37610,N_31504);
nor U43702 (N_43702,N_38336,N_37856);
nand U43703 (N_43703,N_34062,N_37042);
and U43704 (N_43704,N_39946,N_35845);
or U43705 (N_43705,N_31250,N_31756);
and U43706 (N_43706,N_33585,N_31684);
and U43707 (N_43707,N_39861,N_35206);
or U43708 (N_43708,N_36377,N_32821);
or U43709 (N_43709,N_34679,N_35378);
or U43710 (N_43710,N_31281,N_34672);
or U43711 (N_43711,N_38508,N_34072);
and U43712 (N_43712,N_39450,N_31181);
nor U43713 (N_43713,N_32202,N_33373);
nor U43714 (N_43714,N_38091,N_32527);
xor U43715 (N_43715,N_36052,N_37770);
nor U43716 (N_43716,N_36945,N_39528);
nor U43717 (N_43717,N_36226,N_33696);
or U43718 (N_43718,N_38284,N_33648);
nand U43719 (N_43719,N_34980,N_32329);
xnor U43720 (N_43720,N_34235,N_32794);
nand U43721 (N_43721,N_36703,N_38585);
or U43722 (N_43722,N_34337,N_39498);
or U43723 (N_43723,N_38610,N_33324);
and U43724 (N_43724,N_34180,N_30869);
xnor U43725 (N_43725,N_32612,N_36246);
or U43726 (N_43726,N_39455,N_32751);
or U43727 (N_43727,N_30131,N_30977);
nor U43728 (N_43728,N_39992,N_38487);
and U43729 (N_43729,N_34674,N_35717);
xnor U43730 (N_43730,N_39666,N_33504);
or U43731 (N_43731,N_36366,N_37503);
xor U43732 (N_43732,N_36125,N_32274);
xnor U43733 (N_43733,N_35600,N_38728);
nor U43734 (N_43734,N_34715,N_30008);
nand U43735 (N_43735,N_33106,N_31207);
or U43736 (N_43736,N_32952,N_33252);
or U43737 (N_43737,N_38135,N_30251);
and U43738 (N_43738,N_34802,N_30936);
or U43739 (N_43739,N_31830,N_38700);
nand U43740 (N_43740,N_39375,N_34418);
nand U43741 (N_43741,N_34605,N_35193);
or U43742 (N_43742,N_34895,N_32409);
nand U43743 (N_43743,N_37163,N_38937);
nor U43744 (N_43744,N_31928,N_38740);
and U43745 (N_43745,N_36152,N_39827);
or U43746 (N_43746,N_38859,N_31008);
xnor U43747 (N_43747,N_36167,N_37558);
and U43748 (N_43748,N_36942,N_33120);
or U43749 (N_43749,N_30488,N_31320);
xnor U43750 (N_43750,N_38911,N_35571);
nor U43751 (N_43751,N_38786,N_33379);
nor U43752 (N_43752,N_31480,N_36469);
or U43753 (N_43753,N_30668,N_34207);
or U43754 (N_43754,N_32976,N_31522);
and U43755 (N_43755,N_38302,N_39203);
or U43756 (N_43756,N_33476,N_32272);
or U43757 (N_43757,N_36194,N_38388);
or U43758 (N_43758,N_37372,N_36486);
xnor U43759 (N_43759,N_30911,N_37814);
xor U43760 (N_43760,N_35662,N_39604);
nand U43761 (N_43761,N_32310,N_34663);
xnor U43762 (N_43762,N_35003,N_39196);
and U43763 (N_43763,N_38236,N_35316);
xor U43764 (N_43764,N_33609,N_32713);
and U43765 (N_43765,N_37719,N_31960);
xnor U43766 (N_43766,N_37370,N_30523);
or U43767 (N_43767,N_38323,N_32159);
or U43768 (N_43768,N_32050,N_37606);
nor U43769 (N_43769,N_32364,N_36159);
xnor U43770 (N_43770,N_37137,N_33992);
nor U43771 (N_43771,N_31202,N_32235);
and U43772 (N_43772,N_33148,N_36134);
xnor U43773 (N_43773,N_31795,N_37055);
and U43774 (N_43774,N_36348,N_31101);
nand U43775 (N_43775,N_34101,N_39405);
and U43776 (N_43776,N_32793,N_35425);
or U43777 (N_43777,N_31798,N_34039);
or U43778 (N_43778,N_32864,N_39562);
and U43779 (N_43779,N_34519,N_38574);
or U43780 (N_43780,N_34395,N_36691);
and U43781 (N_43781,N_35314,N_35698);
xnor U43782 (N_43782,N_33209,N_38792);
xnor U43783 (N_43783,N_32114,N_39123);
or U43784 (N_43784,N_34476,N_37685);
or U43785 (N_43785,N_32100,N_37754);
and U43786 (N_43786,N_33006,N_39491);
and U43787 (N_43787,N_38631,N_35788);
nand U43788 (N_43788,N_30081,N_34117);
or U43789 (N_43789,N_35774,N_33594);
xor U43790 (N_43790,N_30418,N_36571);
nor U43791 (N_43791,N_34197,N_34015);
or U43792 (N_43792,N_30825,N_34899);
nand U43793 (N_43793,N_39417,N_33500);
xor U43794 (N_43794,N_38087,N_30729);
xnor U43795 (N_43795,N_30141,N_36269);
or U43796 (N_43796,N_39844,N_31061);
or U43797 (N_43797,N_34486,N_38706);
or U43798 (N_43798,N_33617,N_31699);
or U43799 (N_43799,N_30306,N_31326);
nor U43800 (N_43800,N_32646,N_38141);
and U43801 (N_43801,N_32374,N_33254);
nand U43802 (N_43802,N_30077,N_39563);
nand U43803 (N_43803,N_39020,N_31304);
nor U43804 (N_43804,N_34734,N_35042);
nand U43805 (N_43805,N_30776,N_37745);
nand U43806 (N_43806,N_30151,N_31014);
xor U43807 (N_43807,N_35213,N_32552);
or U43808 (N_43808,N_37013,N_38196);
or U43809 (N_43809,N_33241,N_33657);
nor U43810 (N_43810,N_30469,N_33549);
nand U43811 (N_43811,N_34924,N_34635);
xor U43812 (N_43812,N_32790,N_35898);
nand U43813 (N_43813,N_37250,N_38780);
xnor U43814 (N_43814,N_38596,N_34998);
xor U43815 (N_43815,N_35574,N_34485);
xnor U43816 (N_43816,N_38869,N_36347);
nor U43817 (N_43817,N_33141,N_32435);
xnor U43818 (N_43818,N_38878,N_36535);
or U43819 (N_43819,N_31941,N_33207);
nand U43820 (N_43820,N_37782,N_35511);
nand U43821 (N_43821,N_37193,N_37721);
or U43822 (N_43822,N_36496,N_36939);
and U43823 (N_43823,N_38041,N_39570);
xnor U43824 (N_43824,N_37350,N_30439);
nor U43825 (N_43825,N_32902,N_37228);
nor U43826 (N_43826,N_38056,N_33607);
nor U43827 (N_43827,N_37734,N_38013);
xnor U43828 (N_43828,N_32349,N_33938);
nor U43829 (N_43829,N_39976,N_36395);
nor U43830 (N_43830,N_31639,N_36100);
and U43831 (N_43831,N_38286,N_34173);
nor U43832 (N_43832,N_33301,N_32319);
nand U43833 (N_43833,N_36989,N_34403);
or U43834 (N_43834,N_31242,N_33090);
nor U43835 (N_43835,N_30185,N_30274);
or U43836 (N_43836,N_34056,N_30068);
or U43837 (N_43837,N_38817,N_39103);
and U43838 (N_43838,N_39501,N_33096);
or U43839 (N_43839,N_37998,N_31109);
xnor U43840 (N_43840,N_39897,N_33968);
and U43841 (N_43841,N_38694,N_38779);
nand U43842 (N_43842,N_35392,N_32430);
and U43843 (N_43843,N_33515,N_36608);
and U43844 (N_43844,N_36936,N_39247);
xor U43845 (N_43845,N_37064,N_30841);
xor U43846 (N_43846,N_31251,N_31464);
xor U43847 (N_43847,N_32087,N_39017);
and U43848 (N_43848,N_32232,N_39928);
or U43849 (N_43849,N_39094,N_32039);
xnor U43850 (N_43850,N_31024,N_36050);
and U43851 (N_43851,N_33899,N_39730);
xor U43852 (N_43852,N_37344,N_33406);
and U43853 (N_43853,N_35631,N_38554);
and U43854 (N_43854,N_34220,N_37405);
nor U43855 (N_43855,N_36463,N_39855);
xnor U43856 (N_43856,N_34521,N_31636);
xor U43857 (N_43857,N_39660,N_37398);
and U43858 (N_43858,N_31501,N_37940);
nand U43859 (N_43859,N_31840,N_37607);
or U43860 (N_43860,N_39724,N_37548);
and U43861 (N_43861,N_38423,N_33489);
or U43862 (N_43862,N_38158,N_32772);
xnor U43863 (N_43863,N_37207,N_38840);
and U43864 (N_43864,N_33250,N_37850);
nor U43865 (N_43865,N_38000,N_33094);
xor U43866 (N_43866,N_30348,N_33543);
nand U43867 (N_43867,N_38098,N_30399);
xor U43868 (N_43868,N_38685,N_30843);
nand U43869 (N_43869,N_37264,N_37860);
or U43870 (N_43870,N_34131,N_35171);
xor U43871 (N_43871,N_36548,N_33859);
xnor U43872 (N_43872,N_35185,N_37312);
xnor U43873 (N_43873,N_33323,N_31047);
nand U43874 (N_43874,N_35810,N_33410);
xnor U43875 (N_43875,N_39699,N_33157);
nor U43876 (N_43876,N_34350,N_34547);
and U43877 (N_43877,N_38237,N_38992);
nor U43878 (N_43878,N_33231,N_34900);
nand U43879 (N_43879,N_31473,N_39078);
xnor U43880 (N_43880,N_31866,N_30468);
and U43881 (N_43881,N_37033,N_32085);
nand U43882 (N_43882,N_31192,N_32951);
or U43883 (N_43883,N_30464,N_34548);
nor U43884 (N_43884,N_37755,N_37595);
nand U43885 (N_43885,N_36663,N_38103);
xnor U43886 (N_43886,N_32553,N_36000);
nand U43887 (N_43887,N_32414,N_36515);
nand U43888 (N_43888,N_35406,N_34774);
nor U43889 (N_43889,N_35417,N_31372);
nand U43890 (N_43890,N_39366,N_39336);
nand U43891 (N_43891,N_36700,N_34999);
nand U43892 (N_43892,N_30965,N_33027);
nor U43893 (N_43893,N_31059,N_36408);
nor U43894 (N_43894,N_38803,N_32770);
nor U43895 (N_43895,N_33328,N_33114);
xor U43896 (N_43896,N_35037,N_32393);
xnor U43897 (N_43897,N_39176,N_35960);
xor U43898 (N_43898,N_37214,N_35773);
and U43899 (N_43899,N_35710,N_32669);
nor U43900 (N_43900,N_37408,N_39743);
xor U43901 (N_43901,N_39970,N_35167);
nand U43902 (N_43902,N_34300,N_38525);
xnor U43903 (N_43903,N_34692,N_31351);
xnor U43904 (N_43904,N_33434,N_37178);
nand U43905 (N_43905,N_30622,N_39102);
and U43906 (N_43906,N_38611,N_30389);
nor U43907 (N_43907,N_31177,N_32949);
nor U43908 (N_43908,N_39577,N_33567);
xor U43909 (N_43909,N_39621,N_30458);
xor U43910 (N_43910,N_38831,N_32723);
nand U43911 (N_43911,N_33236,N_34618);
and U43912 (N_43912,N_32043,N_33796);
xnor U43913 (N_43913,N_30143,N_39179);
or U43914 (N_43914,N_33125,N_37980);
or U43915 (N_43915,N_31870,N_35970);
and U43916 (N_43916,N_31707,N_36114);
xor U43917 (N_43917,N_39167,N_34531);
or U43918 (N_43918,N_39138,N_30991);
xnor U43919 (N_43919,N_32378,N_31775);
or U43920 (N_43920,N_30303,N_32370);
and U43921 (N_43921,N_31433,N_38651);
nand U43922 (N_43922,N_34143,N_38659);
nand U43923 (N_43923,N_39696,N_39661);
nand U43924 (N_43924,N_38759,N_37608);
or U43925 (N_43925,N_33452,N_32871);
and U43926 (N_43926,N_36753,N_30264);
and U43927 (N_43927,N_32068,N_30128);
nand U43928 (N_43928,N_39589,N_30136);
or U43929 (N_43929,N_30914,N_37688);
xnor U43930 (N_43930,N_36932,N_39824);
and U43931 (N_43931,N_38645,N_32771);
nand U43932 (N_43932,N_31459,N_34507);
or U43933 (N_43933,N_39031,N_38615);
nor U43934 (N_43934,N_38309,N_33422);
nor U43935 (N_43935,N_30031,N_32054);
and U43936 (N_43936,N_36136,N_38194);
xnor U43937 (N_43937,N_37445,N_33070);
xor U43938 (N_43938,N_34656,N_37944);
and U43939 (N_43939,N_37676,N_31288);
and U43940 (N_43940,N_37422,N_35585);
or U43941 (N_43941,N_34296,N_35946);
or U43942 (N_43942,N_39040,N_38975);
nand U43943 (N_43943,N_32925,N_37517);
or U43944 (N_43944,N_33840,N_35939);
and U43945 (N_43945,N_36761,N_30101);
or U43946 (N_43946,N_39227,N_38063);
and U43947 (N_43947,N_38777,N_33145);
nor U43948 (N_43948,N_31088,N_36090);
nand U43949 (N_43949,N_37976,N_33693);
xnor U43950 (N_43950,N_32215,N_38253);
xor U43951 (N_43951,N_34886,N_38549);
or U43952 (N_43952,N_30359,N_36519);
nand U43953 (N_43953,N_36446,N_37879);
and U43954 (N_43954,N_35437,N_36952);
nand U43955 (N_43955,N_30123,N_39086);
xnor U43956 (N_43956,N_39522,N_36451);
xnor U43957 (N_43957,N_37853,N_34424);
and U43958 (N_43958,N_39614,N_37561);
nand U43959 (N_43959,N_30063,N_31362);
nand U43960 (N_43960,N_37835,N_34818);
xor U43961 (N_43961,N_32123,N_32416);
and U43962 (N_43962,N_34250,N_34955);
nand U43963 (N_43963,N_31078,N_34907);
nor U43964 (N_43964,N_30897,N_39235);
nand U43965 (N_43965,N_33359,N_38474);
nand U43966 (N_43966,N_31893,N_32919);
nor U43967 (N_43967,N_39054,N_37448);
and U43968 (N_43968,N_30572,N_36683);
nand U43969 (N_43969,N_39161,N_38081);
or U43970 (N_43970,N_31392,N_35394);
and U43971 (N_43971,N_30855,N_39189);
xor U43972 (N_43972,N_36250,N_33219);
nor U43973 (N_43973,N_35776,N_39232);
or U43974 (N_43974,N_30217,N_32292);
or U43975 (N_43975,N_33690,N_39920);
nand U43976 (N_43976,N_39598,N_33277);
or U43977 (N_43977,N_39771,N_35911);
and U43978 (N_43978,N_34850,N_36499);
xnor U43979 (N_43979,N_35978,N_38592);
nand U43980 (N_43980,N_34331,N_32488);
nor U43981 (N_43981,N_33783,N_30727);
xor U43982 (N_43982,N_33468,N_30998);
and U43983 (N_43983,N_31745,N_36650);
nand U43984 (N_43984,N_34580,N_37434);
nand U43985 (N_43985,N_36640,N_39818);
nor U43986 (N_43986,N_31358,N_36411);
or U43987 (N_43987,N_33932,N_39557);
nor U43988 (N_43988,N_32472,N_34098);
nand U43989 (N_43989,N_35685,N_33097);
nand U43990 (N_43990,N_32259,N_32740);
and U43991 (N_43991,N_37166,N_32269);
xnor U43992 (N_43992,N_34871,N_30436);
xnor U43993 (N_43993,N_34807,N_32802);
and U43994 (N_43994,N_36995,N_33163);
nand U43995 (N_43995,N_33874,N_32369);
and U43996 (N_43996,N_31081,N_31071);
or U43997 (N_43997,N_36503,N_33605);
nand U43998 (N_43998,N_31535,N_34347);
nor U43999 (N_43999,N_34210,N_38821);
xnor U44000 (N_44000,N_39206,N_37740);
nand U44001 (N_44001,N_30529,N_34728);
nand U44002 (N_44002,N_30243,N_30501);
nand U44003 (N_44003,N_31733,N_32185);
and U44004 (N_44004,N_31923,N_34311);
and U44005 (N_44005,N_35466,N_37189);
nor U44006 (N_44006,N_35249,N_32692);
or U44007 (N_44007,N_35469,N_33591);
nor U44008 (N_44008,N_39720,N_38057);
nor U44009 (N_44009,N_39982,N_34438);
xor U44010 (N_44010,N_30205,N_37220);
nand U44011 (N_44011,N_39473,N_37074);
nand U44012 (N_44012,N_39864,N_38757);
nor U44013 (N_44013,N_33026,N_38718);
or U44014 (N_44014,N_33391,N_32513);
nand U44015 (N_44015,N_34011,N_36824);
and U44016 (N_44016,N_37121,N_31588);
xor U44017 (N_44017,N_34690,N_32885);
nor U44018 (N_44018,N_32728,N_31814);
nor U44019 (N_44019,N_39433,N_33194);
nor U44020 (N_44020,N_30511,N_32563);
nor U44021 (N_44021,N_35661,N_33132);
and U44022 (N_44022,N_36913,N_33595);
xor U44023 (N_44023,N_38524,N_39645);
nor U44024 (N_44024,N_36014,N_39575);
and U44025 (N_44025,N_37030,N_35975);
and U44026 (N_44026,N_38263,N_35311);
nor U44027 (N_44027,N_38811,N_39030);
nor U44028 (N_44028,N_37109,N_31196);
xor U44029 (N_44029,N_33113,N_36400);
or U44030 (N_44030,N_34409,N_39788);
xor U44031 (N_44031,N_32064,N_32566);
nand U44032 (N_44032,N_37697,N_35517);
and U44033 (N_44033,N_33490,N_34374);
nand U44034 (N_44034,N_36890,N_39359);
or U44035 (N_44035,N_32882,N_35285);
nor U44036 (N_44036,N_36692,N_39714);
nor U44037 (N_44037,N_38357,N_39516);
and U44038 (N_44038,N_37132,N_33220);
xor U44039 (N_44039,N_35522,N_34103);
or U44040 (N_44040,N_37767,N_38306);
and U44041 (N_44041,N_36969,N_31382);
xnor U44042 (N_44042,N_39401,N_33482);
or U44043 (N_44043,N_39977,N_34322);
xnor U44044 (N_44044,N_38983,N_30886);
nor U44045 (N_44045,N_36625,N_37103);
nor U44046 (N_44046,N_35432,N_31301);
nor U44047 (N_44047,N_33263,N_37056);
nor U44048 (N_44048,N_30974,N_36859);
nor U44049 (N_44049,N_36598,N_30686);
and U44050 (N_44050,N_38048,N_34303);
xor U44051 (N_44051,N_34502,N_30026);
nor U44052 (N_44052,N_31861,N_36189);
nor U44053 (N_44053,N_31558,N_30759);
and U44054 (N_44054,N_36794,N_37319);
nand U44055 (N_44055,N_33831,N_31649);
nor U44056 (N_44056,N_37107,N_35576);
xnor U44057 (N_44057,N_33559,N_34299);
xor U44058 (N_44058,N_32336,N_34550);
nand U44059 (N_44059,N_32366,N_32227);
xor U44060 (N_44060,N_37345,N_35159);
xnor U44061 (N_44061,N_33210,N_30796);
and U44062 (N_44062,N_36070,N_31296);
and U44063 (N_44063,N_32766,N_32923);
and U44064 (N_44064,N_39321,N_34017);
nor U44065 (N_44065,N_31571,N_37634);
xor U44066 (N_44066,N_39416,N_34206);
nand U44067 (N_44067,N_35766,N_32721);
xor U44068 (N_44068,N_35068,N_38096);
or U44069 (N_44069,N_37154,N_38080);
nand U44070 (N_44070,N_38338,N_33949);
and U44071 (N_44071,N_36428,N_38987);
xnor U44072 (N_44072,N_31665,N_33902);
xor U44073 (N_44073,N_39195,N_35677);
nand U44074 (N_44074,N_38322,N_39874);
xnor U44075 (N_44075,N_35258,N_32177);
xor U44076 (N_44076,N_34898,N_34892);
or U44077 (N_44077,N_33792,N_39669);
nor U44078 (N_44078,N_33206,N_38894);
xor U44079 (N_44079,N_39290,N_35621);
nor U44080 (N_44080,N_38489,N_35136);
xor U44081 (N_44081,N_31411,N_33877);
and U44082 (N_44082,N_38370,N_37629);
xnor U44083 (N_44083,N_32848,N_32461);
nand U44084 (N_44084,N_39535,N_32273);
nand U44085 (N_44085,N_35064,N_30338);
nand U44086 (N_44086,N_35836,N_30097);
nand U44087 (N_44087,N_35487,N_39837);
or U44088 (N_44088,N_35607,N_33367);
nor U44089 (N_44089,N_33973,N_32569);
xor U44090 (N_44090,N_30312,N_33151);
nor U44091 (N_44091,N_39154,N_33117);
and U44092 (N_44092,N_37625,N_39700);
or U44093 (N_44093,N_30207,N_36748);
nor U44094 (N_44094,N_34258,N_35355);
and U44095 (N_44095,N_36837,N_30549);
nor U44096 (N_44096,N_36793,N_34176);
and U44097 (N_44097,N_32544,N_33306);
nand U44098 (N_44098,N_37648,N_34049);
nand U44099 (N_44099,N_34335,N_34137);
nand U44100 (N_44100,N_35151,N_37411);
and U44101 (N_44101,N_35900,N_34228);
xor U44102 (N_44102,N_31847,N_33082);
nand U44103 (N_44103,N_35573,N_33764);
or U44104 (N_44104,N_36923,N_33985);
and U44105 (N_44105,N_35887,N_39533);
and U44106 (N_44106,N_32327,N_33499);
and U44107 (N_44107,N_38363,N_37474);
and U44108 (N_44108,N_31647,N_34431);
nor U44109 (N_44109,N_35877,N_32464);
nor U44110 (N_44110,N_34831,N_31482);
and U44111 (N_44111,N_32051,N_31489);
or U44112 (N_44112,N_37038,N_32398);
nor U44113 (N_44113,N_36556,N_32001);
and U44114 (N_44114,N_31483,N_39090);
xnor U44115 (N_44115,N_38176,N_36202);
xnor U44116 (N_44116,N_37023,N_30409);
or U44117 (N_44117,N_35352,N_37943);
or U44118 (N_44118,N_37657,N_30692);
and U44119 (N_44119,N_37566,N_31357);
xor U44120 (N_44120,N_36448,N_31655);
or U44121 (N_44121,N_38301,N_32587);
nor U44122 (N_44122,N_34422,N_39448);
nor U44123 (N_44123,N_34542,N_30195);
or U44124 (N_44124,N_35885,N_30186);
nor U44125 (N_44125,N_36357,N_33012);
or U44126 (N_44126,N_35324,N_31916);
xnor U44127 (N_44127,N_34289,N_31673);
nand U44128 (N_44128,N_34242,N_39752);
xnor U44129 (N_44129,N_34716,N_32506);
xor U44130 (N_44130,N_38972,N_31220);
nand U44131 (N_44131,N_37947,N_30353);
nand U44132 (N_44132,N_36698,N_35869);
xnor U44133 (N_44133,N_38175,N_37637);
nor U44134 (N_44134,N_31159,N_31986);
nand U44135 (N_44135,N_36654,N_35871);
and U44136 (N_44136,N_37246,N_31291);
xnor U44137 (N_44137,N_33524,N_38744);
or U44138 (N_44138,N_39540,N_33436);
or U44139 (N_44139,N_32308,N_37106);
or U44140 (N_44140,N_30619,N_33555);
or U44141 (N_44141,N_37148,N_35018);
nand U44142 (N_44142,N_31319,N_31524);
xnor U44143 (N_44143,N_35280,N_35800);
nand U44144 (N_44144,N_38781,N_39140);
nor U44145 (N_44145,N_35227,N_30861);
and U44146 (N_44146,N_34075,N_36010);
and U44147 (N_44147,N_32601,N_37210);
nand U44148 (N_44148,N_34667,N_32322);
nand U44149 (N_44149,N_35362,N_37040);
and U44150 (N_44150,N_36659,N_37399);
and U44151 (N_44151,N_37413,N_39016);
nor U44152 (N_44152,N_37682,N_31922);
or U44153 (N_44153,N_36587,N_31228);
nor U44154 (N_44154,N_30988,N_31500);
or U44155 (N_44155,N_36231,N_35883);
or U44156 (N_44156,N_36792,N_30463);
xor U44157 (N_44157,N_37034,N_30624);
and U44158 (N_44158,N_34144,N_31077);
and U44159 (N_44159,N_35704,N_32099);
xnor U44160 (N_44160,N_37020,N_39532);
or U44161 (N_44161,N_30883,N_33767);
nor U44162 (N_44162,N_31252,N_32303);
and U44163 (N_44163,N_36981,N_33612);
xnor U44164 (N_44164,N_37221,N_33733);
nand U44165 (N_44165,N_38761,N_33611);
or U44166 (N_44166,N_39566,N_37669);
nand U44167 (N_44167,N_36107,N_38653);
and U44168 (N_44168,N_35952,N_38947);
and U44169 (N_44169,N_35403,N_34364);
nor U44170 (N_44170,N_35827,N_36131);
xnor U44171 (N_44171,N_39762,N_32154);
nand U44172 (N_44172,N_39821,N_39483);
nand U44173 (N_44173,N_38137,N_35958);
or U44174 (N_44174,N_38962,N_30579);
nand U44175 (N_44175,N_34401,N_39098);
nor U44176 (N_44176,N_33014,N_34402);
xnor U44177 (N_44177,N_39216,N_33466);
nor U44178 (N_44178,N_38257,N_39282);
xnor U44179 (N_44179,N_39963,N_35434);
xor U44180 (N_44180,N_30587,N_39383);
nand U44181 (N_44181,N_35477,N_31943);
and U44182 (N_44182,N_34434,N_33189);
and U44183 (N_44183,N_37227,N_39223);
nor U44184 (N_44184,N_36808,N_39228);
or U44185 (N_44185,N_38340,N_33845);
nor U44186 (N_44186,N_39601,N_30757);
nor U44187 (N_44187,N_33182,N_36763);
and U44188 (N_44188,N_39800,N_38914);
nor U44189 (N_44189,N_32834,N_38113);
nor U44190 (N_44190,N_33775,N_30422);
nand U44191 (N_44191,N_32355,N_30134);
and U44192 (N_44192,N_38197,N_31141);
nor U44193 (N_44193,N_39058,N_32639);
nand U44194 (N_44194,N_32838,N_31164);
nand U44195 (N_44195,N_37209,N_37872);
nor U44196 (N_44196,N_34154,N_35540);
nand U44197 (N_44197,N_36586,N_30272);
or U44198 (N_44198,N_36151,N_33478);
and U44199 (N_44199,N_39942,N_37285);
xnor U44200 (N_44200,N_35998,N_32498);
nand U44201 (N_44201,N_32732,N_36414);
xnor U44202 (N_44202,N_34216,N_33295);
xnor U44203 (N_44203,N_33022,N_37126);
nor U44204 (N_44204,N_32993,N_30850);
or U44205 (N_44205,N_39632,N_30403);
or U44206 (N_44206,N_38383,N_30697);
nand U44207 (N_44207,N_32230,N_30001);
nand U44208 (N_44208,N_38656,N_30471);
nand U44209 (N_44209,N_30067,N_38909);
nor U44210 (N_44210,N_33199,N_31661);
xor U44211 (N_44211,N_36265,N_39511);
xor U44212 (N_44212,N_31702,N_31191);
and U44213 (N_44213,N_31770,N_37989);
and U44214 (N_44214,N_32676,N_31697);
or U44215 (N_44215,N_37356,N_35465);
nor U44216 (N_44216,N_36480,N_33811);
and U44217 (N_44217,N_38861,N_31434);
xnor U44218 (N_44218,N_36810,N_35291);
nor U44219 (N_44219,N_38768,N_33289);
nor U44220 (N_44220,N_38117,N_36738);
or U44221 (N_44221,N_35480,N_33752);
nor U44222 (N_44222,N_37334,N_32588);
nor U44223 (N_44223,N_35533,N_38200);
nor U44224 (N_44224,N_38832,N_39011);
or U44225 (N_44225,N_36782,N_37333);
xor U44226 (N_44226,N_31577,N_37536);
and U44227 (N_44227,N_33955,N_38950);
or U44228 (N_44228,N_39512,N_36949);
nand U44229 (N_44229,N_30986,N_30012);
and U44230 (N_44230,N_31951,N_31027);
nand U44231 (N_44231,N_36993,N_39716);
and U44232 (N_44232,N_33164,N_37939);
nand U44233 (N_44233,N_33701,N_35913);
or U44234 (N_44234,N_36809,N_30317);
nand U44235 (N_44235,N_31044,N_34644);
nand U44236 (N_44236,N_35341,N_33285);
xor U44237 (N_44237,N_38782,N_34923);
nand U44238 (N_44238,N_35286,N_34944);
nand U44239 (N_44239,N_37377,N_35813);
xor U44240 (N_44240,N_33408,N_35484);
nand U44241 (N_44241,N_37198,N_34920);
nor U44242 (N_44242,N_34522,N_33820);
nor U44243 (N_44243,N_37205,N_32938);
nor U44244 (N_44244,N_33981,N_32117);
xor U44245 (N_44245,N_30291,N_34913);
and U44246 (N_44246,N_30281,N_39212);
xor U44247 (N_44247,N_39892,N_39826);
and U44248 (N_44248,N_30246,N_36757);
and U44249 (N_44249,N_39832,N_39099);
or U44250 (N_44250,N_30644,N_39384);
or U44251 (N_44251,N_30058,N_38969);
xor U44252 (N_44252,N_35870,N_38912);
and U44253 (N_44253,N_39808,N_33256);
and U44254 (N_44254,N_33161,N_35320);
xnor U44255 (N_44255,N_33784,N_38476);
nor U44256 (N_44256,N_33652,N_36983);
and U44257 (N_44257,N_36870,N_31076);
nor U44258 (N_44258,N_32570,N_35086);
or U44259 (N_44259,N_31285,N_39904);
nand U44260 (N_44260,N_36604,N_38620);
or U44261 (N_44261,N_30938,N_39240);
xnor U44262 (N_44262,N_30344,N_31246);
and U44263 (N_44263,N_31792,N_37884);
and U44264 (N_44264,N_36934,N_39432);
and U44265 (N_44265,N_30194,N_37966);
nand U44266 (N_44266,N_34387,N_31827);
xor U44267 (N_44267,N_37905,N_31586);
nand U44268 (N_44268,N_34759,N_35653);
nand U44269 (N_44269,N_31590,N_31585);
or U44270 (N_44270,N_38539,N_38442);
nor U44271 (N_44271,N_39585,N_37180);
or U44272 (N_44272,N_31206,N_37095);
or U44273 (N_44273,N_35597,N_31559);
nand U44274 (N_44274,N_37437,N_37611);
and U44275 (N_44275,N_39044,N_36679);
or U44276 (N_44276,N_33692,N_31825);
or U44277 (N_44277,N_35146,N_34942);
nor U44278 (N_44278,N_39872,N_31534);
and U44279 (N_44279,N_33834,N_30278);
nand U44280 (N_44280,N_33146,N_38881);
or U44281 (N_44281,N_39787,N_35865);
nor U44282 (N_44282,N_36017,N_34842);
and U44283 (N_44283,N_39191,N_34308);
xor U44284 (N_44284,N_35577,N_37012);
xnor U44285 (N_44285,N_32955,N_32195);
and U44286 (N_44286,N_39326,N_33033);
xnor U44287 (N_44287,N_39849,N_35632);
or U44288 (N_44288,N_39915,N_33085);
xor U44289 (N_44289,N_31268,N_36055);
nand U44290 (N_44290,N_38655,N_36712);
nor U44291 (N_44291,N_37945,N_36335);
nand U44292 (N_44292,N_33776,N_36157);
or U44293 (N_44293,N_35080,N_33728);
nand U44294 (N_44294,N_31616,N_34463);
xnor U44295 (N_44295,N_35383,N_31690);
xor U44296 (N_44296,N_30677,N_33481);
nand U44297 (N_44297,N_30340,N_37475);
nand U44298 (N_44298,N_37309,N_38903);
nor U44299 (N_44299,N_38756,N_39352);
or U44300 (N_44300,N_33110,N_32439);
or U44301 (N_44301,N_36590,N_35840);
nor U44302 (N_44302,N_38097,N_36864);
xnor U44303 (N_44303,N_39399,N_35812);
xor U44304 (N_44304,N_36392,N_32542);
nor U44305 (N_44305,N_37213,N_33233);
and U44306 (N_44306,N_35559,N_32143);
xor U44307 (N_44307,N_38854,N_38217);
xor U44308 (N_44308,N_38636,N_32455);
xnor U44309 (N_44309,N_31184,N_39842);
and U44310 (N_44310,N_33073,N_34662);
xor U44311 (N_44311,N_30608,N_37301);
nand U44312 (N_44312,N_34538,N_32020);
and U44313 (N_44313,N_36573,N_31016);
xor U44314 (N_44314,N_39238,N_32891);
and U44315 (N_44315,N_33563,N_31496);
or U44316 (N_44316,N_34306,N_30365);
and U44317 (N_44317,N_34909,N_38886);
nand U44318 (N_44318,N_31552,N_31050);
or U44319 (N_44319,N_30669,N_34264);
or U44320 (N_44320,N_37806,N_37643);
nand U44321 (N_44321,N_34116,N_33862);
nor U44322 (N_44322,N_39802,N_39361);
or U44323 (N_44323,N_35918,N_32481);
xnor U44324 (N_44324,N_38448,N_33592);
nand U44325 (N_44325,N_37550,N_36752);
or U44326 (N_44326,N_30425,N_32031);
and U44327 (N_44327,N_34067,N_31165);
xnor U44328 (N_44328,N_37293,N_36009);
nand U44329 (N_44329,N_34461,N_39390);
or U44330 (N_44330,N_39388,N_37733);
and U44331 (N_44331,N_33606,N_32991);
and U44332 (N_44332,N_36996,N_30646);
or U44333 (N_44333,N_31211,N_33028);
nor U44334 (N_44334,N_30512,N_38707);
xnor U44335 (N_44335,N_33169,N_37974);
and U44336 (N_44336,N_35920,N_32814);
or U44337 (N_44337,N_30242,N_32330);
nand U44338 (N_44338,N_33430,N_36054);
or U44339 (N_44339,N_37592,N_36689);
nand U44340 (N_44340,N_37942,N_30118);
xor U44341 (N_44341,N_39772,N_36341);
nor U44342 (N_44342,N_32860,N_32844);
nand U44343 (N_44343,N_34014,N_31677);
nand U44344 (N_44344,N_33494,N_36534);
or U44345 (N_44345,N_31852,N_37573);
nand U44346 (N_44346,N_32360,N_35896);
xor U44347 (N_44347,N_38875,N_39482);
nand U44348 (N_44348,N_34022,N_37647);
and U44349 (N_44349,N_30948,N_37165);
and U44350 (N_44350,N_32671,N_36749);
nand U44351 (N_44351,N_36149,N_36614);
or U44352 (N_44352,N_30169,N_33309);
or U44353 (N_44353,N_35011,N_34589);
or U44354 (N_44354,N_34174,N_34277);
xor U44355 (N_44355,N_37962,N_31026);
nor U44356 (N_44356,N_32840,N_38009);
xnor U44357 (N_44357,N_37150,N_36842);
nand U44358 (N_44358,N_31620,N_37298);
xor U44359 (N_44359,N_32289,N_33581);
xor U44360 (N_44360,N_34647,N_32124);
xnor U44361 (N_44361,N_33711,N_31780);
and U44362 (N_44362,N_31474,N_31331);
or U44363 (N_44363,N_35749,N_34693);
nor U44364 (N_44364,N_36754,N_31255);
or U44365 (N_44365,N_37758,N_32768);
nor U44366 (N_44366,N_32450,N_33873);
nor U44367 (N_44367,N_39369,N_30873);
nor U44368 (N_44368,N_30315,N_39544);
or U44369 (N_44369,N_31637,N_39965);
or U44370 (N_44370,N_32125,N_34864);
nand U44371 (N_44371,N_31368,N_34411);
and U44372 (N_44372,N_34571,N_30939);
nand U44373 (N_44373,N_35399,N_32762);
and U44374 (N_44374,N_34611,N_38093);
and U44375 (N_44375,N_34070,N_30931);
or U44376 (N_44376,N_36631,N_37718);
xnor U44377 (N_44377,N_36254,N_31009);
xnor U44378 (N_44378,N_32412,N_30319);
nand U44379 (N_44379,N_39639,N_36033);
and U44380 (N_44380,N_38538,N_32653);
and U44381 (N_44381,N_39255,N_39998);
nand U44382 (N_44382,N_37049,N_39941);
nor U44383 (N_44383,N_35101,N_33258);
xnor U44384 (N_44384,N_32888,N_36634);
nor U44385 (N_44385,N_31738,N_37891);
xor U44386 (N_44386,N_37378,N_33166);
nor U44387 (N_44387,N_31966,N_37402);
nor U44388 (N_44388,N_33016,N_37693);
xor U44389 (N_44389,N_38307,N_34970);
nor U44390 (N_44390,N_30631,N_38809);
nor U44391 (N_44391,N_38028,N_32256);
or U44392 (N_44392,N_30527,N_35110);
nor U44393 (N_44393,N_34259,N_31842);
or U44394 (N_44394,N_39263,N_39221);
nor U44395 (N_44395,N_38960,N_34727);
nand U44396 (N_44396,N_38988,N_39244);
nor U44397 (N_44397,N_38246,N_39377);
nor U44398 (N_44398,N_36867,N_36013);
or U44399 (N_44399,N_36961,N_39097);
nand U44400 (N_44400,N_33218,N_35446);
or U44401 (N_44401,N_36498,N_35025);
and U44402 (N_44402,N_34227,N_36990);
and U44403 (N_44403,N_30892,N_37785);
xnor U44404 (N_44404,N_39596,N_37931);
or U44405 (N_44405,N_32142,N_31069);
and U44406 (N_44406,N_30460,N_33147);
xnor U44407 (N_44407,N_32747,N_31455);
or U44408 (N_44408,N_31377,N_33726);
xor U44409 (N_44409,N_38534,N_37439);
xnor U44410 (N_44410,N_34718,N_37977);
nor U44411 (N_44411,N_35332,N_30743);
nand U44412 (N_44412,N_34209,N_32029);
and U44413 (N_44413,N_35879,N_35460);
nor U44414 (N_44414,N_34917,N_33420);
xnor U44415 (N_44415,N_38330,N_31105);
nor U44416 (N_44416,N_35455,N_36505);
nand U44417 (N_44417,N_33780,N_36528);
or U44418 (N_44418,N_31826,N_38316);
nor U44419 (N_44419,N_37728,N_33964);
nor U44420 (N_44420,N_37435,N_39534);
nand U44421 (N_44421,N_30304,N_32594);
xnor U44422 (N_44422,N_30332,N_33402);
xnor U44423 (N_44423,N_34436,N_34129);
nand U44424 (N_44424,N_34128,N_32824);
or U44425 (N_44425,N_32113,N_34033);
nor U44426 (N_44426,N_38249,N_30241);
or U44427 (N_44427,N_37763,N_32320);
and U44428 (N_44428,N_31204,N_33292);
nor U44429 (N_44429,N_39969,N_30502);
or U44430 (N_44430,N_38020,N_35397);
nor U44431 (N_44431,N_32876,N_30115);
or U44432 (N_44432,N_34427,N_37289);
or U44433 (N_44433,N_37248,N_37388);
and U44434 (N_44434,N_39561,N_34012);
and U44435 (N_44435,N_33994,N_31454);
or U44436 (N_44436,N_38191,N_38010);
xor U44437 (N_44437,N_38531,N_32850);
xor U44438 (N_44438,N_31070,N_39526);
nor U44439 (N_44439,N_38358,N_39784);
or U44440 (N_44440,N_39737,N_33293);
or U44441 (N_44441,N_35343,N_37255);
or U44442 (N_44442,N_38372,N_39717);
xnor U44443 (N_44443,N_39296,N_34764);
and U44444 (N_44444,N_36593,N_34161);
xor U44445 (N_44445,N_34579,N_30603);
nor U44446 (N_44446,N_39979,N_31471);
xnor U44447 (N_44447,N_33908,N_39680);
xnor U44448 (N_44448,N_39974,N_32748);
or U44449 (N_44449,N_37623,N_33011);
or U44450 (N_44450,N_32660,N_35162);
xor U44451 (N_44451,N_38945,N_33789);
xnor U44452 (N_44452,N_37635,N_38630);
nor U44453 (N_44453,N_31444,N_31901);
nand U44454 (N_44454,N_31084,N_33457);
and U44455 (N_44455,N_31429,N_38677);
and U44456 (N_44456,N_38836,N_34123);
nand U44457 (N_44457,N_32629,N_30750);
and U44458 (N_44458,N_39413,N_31100);
xnor U44459 (N_44459,N_39306,N_37554);
and U44460 (N_44460,N_31506,N_34916);
or U44461 (N_44461,N_39569,N_34838);
nor U44462 (N_44462,N_33103,N_38470);
nor U44463 (N_44463,N_39496,N_31718);
xnor U44464 (N_44464,N_32846,N_31386);
xor U44465 (N_44465,N_31961,N_35680);
xor U44466 (N_44466,N_30416,N_36976);
or U44467 (N_44467,N_30447,N_30176);
nand U44468 (N_44468,N_32295,N_37116);
nand U44469 (N_44469,N_33221,N_30600);
nor U44470 (N_44470,N_31189,N_32808);
xnor U44471 (N_44471,N_39693,N_33627);
xnor U44472 (N_44472,N_39365,N_33496);
nor U44473 (N_44473,N_36312,N_36457);
nor U44474 (N_44474,N_37224,N_39763);
nand U44475 (N_44475,N_30177,N_39023);
nor U44476 (N_44476,N_32458,N_34095);
or U44477 (N_44477,N_34754,N_37480);
and U44478 (N_44478,N_35282,N_33334);
xor U44479 (N_44479,N_35599,N_36360);
or U44480 (N_44480,N_37863,N_39869);
and U44481 (N_44481,N_35926,N_37346);
or U44482 (N_44482,N_33129,N_33778);
and U44483 (N_44483,N_36212,N_35915);
xnor U44484 (N_44484,N_37169,N_31379);
and U44485 (N_44485,N_33815,N_39218);
nand U44486 (N_44486,N_32523,N_35384);
nor U44487 (N_44487,N_36732,N_31439);
and U44488 (N_44488,N_30565,N_36852);
nor U44489 (N_44489,N_34483,N_33635);
nor U44490 (N_44490,N_31935,N_38729);
xor U44491 (N_44491,N_33830,N_31784);
or U44492 (N_44492,N_39708,N_30555);
and U44493 (N_44493,N_36259,N_39617);
nand U44494 (N_44494,N_34673,N_36978);
nand U44495 (N_44495,N_36482,N_37262);
or U44496 (N_44496,N_32887,N_39148);
or U44497 (N_44497,N_35864,N_30794);
or U44498 (N_44498,N_39342,N_35492);
or U44499 (N_44499,N_35100,N_37621);
and U44500 (N_44500,N_31881,N_33511);
or U44501 (N_44501,N_31867,N_31328);
nor U44502 (N_44502,N_39765,N_39121);
nand U44503 (N_44503,N_32266,N_36883);
nor U44504 (N_44504,N_32541,N_33050);
or U44505 (N_44505,N_36884,N_38762);
nor U44506 (N_44506,N_33814,N_35115);
and U44507 (N_44507,N_30240,N_36817);
xnor U44508 (N_44508,N_34869,N_37689);
and U44509 (N_44509,N_30040,N_31513);
nor U44510 (N_44510,N_30594,N_39591);
or U44511 (N_44511,N_31481,N_37815);
and U44512 (N_44512,N_36841,N_33450);
nor U44513 (N_44513,N_36866,N_33351);
or U44514 (N_44514,N_32855,N_31863);
nand U44515 (N_44515,N_33572,N_36729);
or U44516 (N_44516,N_35271,N_36611);
nor U44517 (N_44517,N_34752,N_35002);
and U44518 (N_44518,N_37499,N_37915);
and U44519 (N_44519,N_32239,N_37681);
nand U44520 (N_44520,N_32530,N_34826);
nor U44521 (N_44521,N_34841,N_31954);
nand U44522 (N_44522,N_32392,N_30357);
and U44523 (N_44523,N_33600,N_31734);
nand U44524 (N_44524,N_38328,N_31598);
xor U44525 (N_44525,N_39351,N_36363);
nor U44526 (N_44526,N_32990,N_36062);
or U44527 (N_44527,N_31408,N_38801);
and U44528 (N_44528,N_38274,N_35768);
xnor U44529 (N_44529,N_31082,N_34488);
nor U44530 (N_44530,N_30314,N_32079);
and U44531 (N_44531,N_38537,N_31630);
and U44532 (N_44532,N_39729,N_30223);
xnor U44533 (N_44533,N_33763,N_38321);
nand U44534 (N_44534,N_38038,N_31187);
nand U44535 (N_44535,N_36453,N_35134);
nand U44536 (N_44536,N_39584,N_35143);
nand U44537 (N_44537,N_37999,N_30573);
or U44538 (N_44538,N_39130,N_31342);
or U44539 (N_44539,N_36204,N_37348);
or U44540 (N_44540,N_31777,N_33837);
and U44541 (N_44541,N_37716,N_35174);
or U44542 (N_44542,N_39812,N_37173);
or U44543 (N_44543,N_30410,N_32828);
nor U44544 (N_44544,N_35878,N_31652);
nor U44545 (N_44545,N_38389,N_30429);
or U44546 (N_44546,N_35202,N_34943);
nand U44547 (N_44547,N_30798,N_32843);
xor U44548 (N_44548,N_36443,N_32657);
xnor U44549 (N_44549,N_37961,N_38815);
or U44550 (N_44550,N_33004,N_38561);
xor U44551 (N_44551,N_35503,N_30478);
and U44552 (N_44552,N_32825,N_36365);
or U44553 (N_44553,N_36074,N_38203);
nand U44554 (N_44554,N_39502,N_34783);
nor U44555 (N_44555,N_39694,N_32307);
xnor U44556 (N_44556,N_32557,N_33418);
xnor U44557 (N_44557,N_33773,N_33372);
or U44558 (N_44558,N_33536,N_39143);
nor U44559 (N_44559,N_30346,N_35057);
or U44560 (N_44560,N_39814,N_39911);
nor U44561 (N_44561,N_31265,N_33284);
xnor U44562 (N_44562,N_30122,N_32927);
xor U44563 (N_44563,N_30009,N_30145);
xor U44564 (N_44564,N_38514,N_31972);
nand U44565 (N_44565,N_36655,N_33108);
nor U44566 (N_44566,N_38173,N_32680);
nand U44567 (N_44567,N_33574,N_38155);
and U44568 (N_44568,N_37084,N_32005);
nor U44569 (N_44569,N_31096,N_37477);
xnor U44570 (N_44570,N_33412,N_32352);
xnor U44571 (N_44571,N_37263,N_31965);
and U44572 (N_44572,N_36095,N_38638);
or U44573 (N_44573,N_38293,N_35705);
and U44574 (N_44574,N_37299,N_35957);
nor U44575 (N_44575,N_33361,N_35696);
and U44576 (N_44576,N_35128,N_37784);
and U44577 (N_44577,N_37700,N_35428);
xnor U44578 (N_44578,N_37100,N_33913);
nor U44579 (N_44579,N_30125,N_34194);
xnor U44580 (N_44580,N_31528,N_38149);
or U44581 (N_44581,N_38529,N_33875);
nor U44582 (N_44582,N_34660,N_30275);
nand U44583 (N_44583,N_30465,N_38712);
and U44584 (N_44584,N_32346,N_33894);
xor U44585 (N_44585,N_36144,N_33674);
and U44586 (N_44586,N_32839,N_34711);
xor U44587 (N_44587,N_30218,N_39805);
or U44588 (N_44588,N_31194,N_38356);
nand U44589 (N_44589,N_35844,N_38484);
nor U44590 (N_44590,N_36389,N_35694);
nor U44591 (N_44591,N_38308,N_36459);
xor U44592 (N_44592,N_32313,N_31625);
xnor U44593 (N_44593,N_35857,N_37387);
or U44594 (N_44594,N_36082,N_36091);
or U44595 (N_44595,N_33357,N_31010);
nand U44596 (N_44596,N_31950,N_36171);
or U44597 (N_44597,N_31467,N_32944);
or U44598 (N_44598,N_35288,N_31478);
nor U44599 (N_44599,N_38360,N_37509);
or U44600 (N_44600,N_39136,N_31832);
nor U44601 (N_44601,N_39329,N_32178);
nand U44602 (N_44602,N_31334,N_31025);
xnor U44603 (N_44603,N_38090,N_34118);
xnor U44604 (N_44604,N_38375,N_37516);
nor U44605 (N_44605,N_33265,N_32328);
nor U44606 (N_44606,N_31947,N_36053);
and U44607 (N_44607,N_30045,N_36484);
or U44608 (N_44608,N_33640,N_33046);
xnor U44609 (N_44609,N_39126,N_33203);
xor U44610 (N_44610,N_30459,N_38731);
and U44611 (N_44611,N_32935,N_34214);
nand U44612 (N_44612,N_37541,N_39173);
or U44613 (N_44613,N_34102,N_38705);
or U44614 (N_44614,N_30297,N_34226);
xor U44615 (N_44615,N_37803,N_30172);
or U44616 (N_44616,N_32593,N_32271);
and U44617 (N_44617,N_35699,N_33513);
xnor U44618 (N_44618,N_34570,N_34775);
or U44619 (N_44619,N_36041,N_39555);
nor U44620 (N_44620,N_32459,N_38291);
xnor U44621 (N_44621,N_35794,N_38273);
nor U44622 (N_44622,N_30985,N_35457);
nor U44623 (N_44623,N_31197,N_30979);
and U44624 (N_44624,N_37680,N_38084);
and U44625 (N_44625,N_38888,N_32536);
and U44626 (N_44626,N_32152,N_30421);
and U44627 (N_44627,N_38499,N_30514);
nand U44628 (N_44628,N_35548,N_38161);
nor U44629 (N_44629,N_35880,N_32139);
and U44630 (N_44630,N_37832,N_32811);
nor U44631 (N_44631,N_32478,N_30239);
or U44632 (N_44632,N_32854,N_38593);
xor U44633 (N_44633,N_34363,N_33756);
and U44634 (N_44634,N_35380,N_39759);
nor U44635 (N_44635,N_39651,N_36833);
nor U44636 (N_44636,N_35421,N_37918);
xnor U44637 (N_44637,N_33392,N_38347);
nand U44638 (N_44638,N_37902,N_32004);
or U44639 (N_44639,N_32573,N_36955);
xor U44640 (N_44640,N_39886,N_32754);
or U44641 (N_44641,N_39541,N_36543);
or U44642 (N_44642,N_38417,N_35197);
or U44643 (N_44643,N_30700,N_30363);
nand U44644 (N_44644,N_33472,N_32681);
xor U44645 (N_44645,N_36777,N_31465);
or U44646 (N_44646,N_31660,N_39209);
or U44647 (N_44647,N_39587,N_37177);
nand U44648 (N_44648,N_33685,N_36827);
xnor U44649 (N_44649,N_38883,N_34528);
and U44650 (N_44650,N_39105,N_36581);
nand U44651 (N_44651,N_34132,N_32550);
and U44652 (N_44652,N_37557,N_31198);
nor U44653 (N_44653,N_35297,N_37525);
xnor U44654 (N_44654,N_39576,N_39091);
or U44655 (N_44655,N_31173,N_35424);
xor U44656 (N_44656,N_30932,N_36560);
nand U44657 (N_44657,N_32456,N_30652);
nand U44658 (N_44658,N_38327,N_34985);
nand U44659 (N_44659,N_34482,N_31695);
xnor U44660 (N_44660,N_31622,N_32904);
nor U44661 (N_44661,N_39726,N_39385);
xor U44662 (N_44662,N_32080,N_32399);
nand U44663 (N_44663,N_30649,N_38265);
and U44664 (N_44664,N_36419,N_33208);
nor U44665 (N_44665,N_37631,N_33508);
xor U44666 (N_44666,N_33950,N_33891);
xor U44667 (N_44667,N_31013,N_38245);
xor U44668 (N_44668,N_36380,N_31618);
xnor U44669 (N_44669,N_30364,N_34408);
and U44670 (N_44670,N_32917,N_32325);
or U44671 (N_44671,N_37047,N_38177);
nor U44672 (N_44672,N_39009,N_36768);
nor U44673 (N_44673,N_35010,N_32534);
nand U44674 (N_44674,N_30639,N_38147);
and U44675 (N_44675,N_39262,N_34984);
and U44676 (N_44676,N_34170,N_33779);
nor U44677 (N_44677,N_39317,N_34926);
xnor U44678 (N_44678,N_37930,N_39949);
and U44679 (N_44679,N_38714,N_31885);
nor U44680 (N_44680,N_38971,N_35888);
and U44681 (N_44681,N_34994,N_31166);
xnor U44682 (N_44682,N_34642,N_33647);
xnor U44683 (N_44683,N_33624,N_38755);
nand U44684 (N_44684,N_34317,N_31583);
nor U44685 (N_44685,N_34549,N_30515);
and U44686 (N_44686,N_33084,N_37898);
nand U44687 (N_44687,N_39141,N_30455);
and U44688 (N_44688,N_31468,N_36555);
and U44689 (N_44689,N_39686,N_36287);
nand U44690 (N_44690,N_34338,N_37091);
or U44691 (N_44691,N_34276,N_37046);
or U44692 (N_44692,N_30530,N_33628);
nand U44693 (N_44693,N_39776,N_36904);
xnor U44694 (N_44694,N_38068,N_31310);
or U44695 (N_44695,N_32880,N_36475);
xnor U44696 (N_44696,N_35995,N_37361);
nand U44697 (N_44697,N_30954,N_33239);
or U44698 (N_44698,N_30602,N_30984);
nand U44699 (N_44699,N_36092,N_38199);
nand U44700 (N_44700,N_39889,N_38512);
nand U44701 (N_44701,N_37658,N_33839);
nand U44702 (N_44702,N_38509,N_38435);
or U44703 (N_44703,N_32135,N_38331);
xnor U44704 (N_44704,N_39828,N_38045);
nand U44705 (N_44705,N_37291,N_33812);
and U44706 (N_44706,N_38409,N_37394);
nor U44707 (N_44707,N_33608,N_31527);
xor U44708 (N_44708,N_35120,N_35325);
nand U44709 (N_44709,N_32069,N_37094);
nor U44710 (N_44710,N_38353,N_34566);
nor U44711 (N_44711,N_32297,N_30822);
or U44712 (N_44712,N_38247,N_30612);
and U44713 (N_44713,N_35723,N_31562);
xnor U44714 (N_44714,N_37912,N_33512);
and U44715 (N_44715,N_39529,N_36880);
and U44716 (N_44716,N_32288,N_35706);
or U44717 (N_44717,N_38429,N_31573);
xnor U44718 (N_44718,N_34026,N_31824);
and U44719 (N_44719,N_36966,N_37885);
xnor U44720 (N_44720,N_39559,N_38461);
nand U44721 (N_44721,N_30901,N_31701);
or U44722 (N_44722,N_36798,N_39517);
nand U44723 (N_44723,N_32024,N_38216);
and U44724 (N_44724,N_39334,N_36583);
xor U44725 (N_44725,N_39906,N_35808);
xor U44726 (N_44726,N_30930,N_34046);
xor U44727 (N_44727,N_30132,N_34797);
and U44728 (N_44728,N_35402,N_39041);
nand U44729 (N_44729,N_37027,N_38116);
xor U44730 (N_44730,N_33115,N_36126);
and U44731 (N_44731,N_30935,N_37006);
or U44732 (N_44732,N_32956,N_33714);
xor U44733 (N_44733,N_34766,N_32894);
nand U44734 (N_44734,N_38485,N_34239);
and U44735 (N_44735,N_37314,N_36068);
nor U44736 (N_44736,N_36518,N_38403);
nand U44737 (N_44737,N_34295,N_37970);
xor U44738 (N_44738,N_37036,N_34198);
nand U44739 (N_44739,N_36577,N_32608);
nor U44740 (N_44740,N_33590,N_33017);
or U44741 (N_44741,N_38770,N_32830);
nor U44742 (N_44742,N_36155,N_34652);
nor U44743 (N_44743,N_34812,N_39392);
or U44744 (N_44744,N_35246,N_33290);
xnor U44745 (N_44745,N_38392,N_31254);
nor U44746 (N_44746,N_38044,N_35614);
nor U44747 (N_44747,N_37938,N_39311);
nor U44748 (N_44748,N_31560,N_38518);
nand U44749 (N_44749,N_39222,N_35140);
or U44750 (N_44750,N_38976,N_36123);
xor U44751 (N_44751,N_36711,N_30678);
and U44752 (N_44752,N_33404,N_39484);
nand U44753 (N_44753,N_32535,N_35993);
nand U44754 (N_44754,N_31098,N_34524);
nand U44755 (N_44755,N_39174,N_30130);
nor U44756 (N_44756,N_38267,N_31493);
or U44757 (N_44757,N_39069,N_39389);
nor U44758 (N_44758,N_37564,N_38628);
or U44759 (N_44759,N_35478,N_38244);
and U44760 (N_44760,N_32964,N_39527);
or U44761 (N_44761,N_35586,N_36765);
nand U44762 (N_44762,N_32712,N_39705);
nand U44763 (N_44763,N_31277,N_39129);
nor U44764 (N_44764,N_30237,N_32160);
nand U44765 (N_44765,N_34978,N_38635);
nor U44766 (N_44766,N_39909,N_32199);
xnor U44767 (N_44767,N_30845,N_38934);
and U44768 (N_44768,N_39093,N_39745);
xor U44769 (N_44769,N_34848,N_32057);
or U44770 (N_44770,N_34976,N_31156);
and U44771 (N_44771,N_30276,N_34160);
nand U44772 (N_44772,N_39307,N_33133);
nand U44773 (N_44773,N_39425,N_37691);
xor U44774 (N_44774,N_33983,N_37386);
or U44775 (N_44775,N_30311,N_38734);
or U44776 (N_44776,N_30443,N_36986);
nor U44777 (N_44777,N_38025,N_32602);
or U44778 (N_44778,N_34997,N_30313);
xor U44779 (N_44779,N_39612,N_39918);
nand U44780 (N_44780,N_34890,N_31835);
and U44781 (N_44781,N_34089,N_30028);
nor U44782 (N_44782,N_30216,N_33192);
nand U44783 (N_44783,N_35102,N_32969);
nand U44784 (N_44784,N_35344,N_35433);
nor U44785 (N_44785,N_39590,N_38242);
xor U44786 (N_44786,N_34468,N_30562);
or U44787 (N_44787,N_33571,N_31680);
xor U44788 (N_44788,N_33327,N_39773);
or U44789 (N_44789,N_37407,N_36566);
xor U44790 (N_44790,N_35783,N_30666);
nor U44791 (N_44791,N_39790,N_39350);
nand U44792 (N_44792,N_32540,N_32973);
nor U44793 (N_44793,N_34805,N_38115);
and U44794 (N_44794,N_39120,N_31715);
or U44795 (N_44795,N_38853,N_39128);
nand U44796 (N_44796,N_35504,N_38082);
or U44797 (N_44797,N_31505,N_36606);
or U44798 (N_44798,N_35690,N_32151);
nand U44799 (N_44799,N_35452,N_32429);
nand U44800 (N_44800,N_30287,N_39894);
xor U44801 (N_44801,N_31248,N_39234);
nand U44802 (N_44802,N_38533,N_37391);
or U44803 (N_44803,N_38545,N_30980);
and U44804 (N_44804,N_39131,N_33610);
nand U44805 (N_44805,N_39835,N_34023);
nor U44806 (N_44806,N_31344,N_39606);
and U44807 (N_44807,N_38168,N_31539);
and U44808 (N_44808,N_36931,N_39298);
nand U44809 (N_44809,N_34945,N_39833);
or U44810 (N_44810,N_39630,N_34948);
nand U44811 (N_44811,N_30283,N_38070);
and U44812 (N_44812,N_35842,N_33632);
and U44813 (N_44813,N_38479,N_38457);
xnor U44814 (N_44814,N_37496,N_30543);
nor U44815 (N_44815,N_31855,N_39477);
and U44816 (N_44816,N_38138,N_33448);
or U44817 (N_44817,N_34371,N_31550);
or U44818 (N_44818,N_34453,N_39437);
nor U44819 (N_44819,N_32003,N_32797);
and U44820 (N_44820,N_38691,N_35735);
and U44821 (N_44821,N_37281,N_30765);
xor U44822 (N_44822,N_34294,N_36021);
nand U44823 (N_44823,N_31757,N_36339);
or U44824 (N_44824,N_36963,N_37008);
nor U44825 (N_44825,N_39315,N_35907);
nor U44826 (N_44826,N_30712,N_33537);
xnor U44827 (N_44827,N_37829,N_31313);
and U44828 (N_44828,N_36506,N_37272);
and U44829 (N_44829,N_32767,N_31118);
and U44830 (N_44830,N_33353,N_36553);
xor U44831 (N_44831,N_31917,N_36681);
or U44832 (N_44832,N_35843,N_35187);
or U44833 (N_44833,N_34050,N_38788);
nand U44834 (N_44834,N_30405,N_38648);
nand U44835 (N_44835,N_33999,N_34793);
or U44836 (N_44836,N_38290,N_32749);
nand U44837 (N_44837,N_34291,N_32088);
nor U44838 (N_44838,N_39065,N_39363);
and U44839 (N_44839,N_39285,N_33283);
and U44840 (N_44840,N_35179,N_30942);
nor U44841 (N_44841,N_39830,N_31906);
or U44842 (N_44842,N_35289,N_33156);
and U44843 (N_44843,N_36024,N_39107);
xor U44844 (N_44844,N_37195,N_35763);
and U44845 (N_44845,N_35023,N_37459);
nor U44846 (N_44846,N_34857,N_34541);
nand U44847 (N_44847,N_38078,N_33918);
xor U44848 (N_44848,N_38637,N_32390);
xnor U44849 (N_44849,N_37560,N_33871);
or U44850 (N_44850,N_33663,N_32791);
xnor U44851 (N_44851,N_35345,N_30198);
xor U44852 (N_44852,N_33483,N_38337);
or U44853 (N_44853,N_30229,N_34791);
xnor U44854 (N_44854,N_39064,N_34083);
and U44855 (N_44855,N_31007,N_30801);
xor U44856 (N_44856,N_33020,N_33009);
and U44857 (N_44857,N_37112,N_34333);
xor U44858 (N_44858,N_37834,N_35330);
xor U44859 (N_44859,N_39424,N_34265);
nand U44860 (N_44860,N_38644,N_39022);
nor U44861 (N_44861,N_34425,N_34450);
and U44862 (N_44862,N_32283,N_34963);
nor U44863 (N_44863,N_30758,N_30073);
nor U44864 (N_44864,N_39865,N_32516);
nor U44865 (N_44865,N_37167,N_36848);
or U44866 (N_44866,N_33979,N_37254);
xor U44867 (N_44867,N_38112,N_33080);
and U44868 (N_44868,N_38393,N_34931);
and U44869 (N_44869,N_35897,N_34355);
or U44870 (N_44870,N_38278,N_38396);
nand U44871 (N_44871,N_32632,N_34750);
nor U44872 (N_44872,N_33341,N_35313);
and U44873 (N_44873,N_35105,N_31380);
and U44874 (N_44874,N_35852,N_38407);
nor U44875 (N_44875,N_38748,N_38944);
nor U44876 (N_44876,N_35531,N_35409);
and U44877 (N_44877,N_34551,N_32642);
and U44878 (N_44878,N_39077,N_30400);
or U44879 (N_44879,N_30268,N_32999);
nor U44880 (N_44880,N_34464,N_34633);
nand U44881 (N_44881,N_34155,N_30545);
and U44882 (N_44882,N_34648,N_32365);
xnor U44883 (N_44883,N_35816,N_35988);
and U44884 (N_44884,N_35846,N_33801);
and U44885 (N_44885,N_31338,N_37575);
nand U44886 (N_44886,N_31713,N_39769);
nor U44887 (N_44887,N_37120,N_38211);
or U44888 (N_44888,N_34396,N_34813);
xor U44889 (N_44889,N_31448,N_31415);
xnor U44890 (N_44890,N_36690,N_31183);
nand U44891 (N_44891,N_36524,N_37075);
xnor U44892 (N_44892,N_30791,N_38411);
and U44893 (N_44893,N_33702,N_35956);
or U44894 (N_44894,N_33636,N_33344);
or U44895 (N_44895,N_30494,N_31850);
and U44896 (N_44896,N_30929,N_32847);
xnor U44897 (N_44897,N_35709,N_39059);
or U44898 (N_44898,N_34415,N_37339);
nor U44899 (N_44899,N_35408,N_36329);
xnor U44900 (N_44900,N_32407,N_37253);
nor U44901 (N_44901,N_39202,N_33383);
xor U44902 (N_44902,N_33958,N_31475);
nand U44903 (N_44903,N_36572,N_38558);
xor U44904 (N_44904,N_36279,N_38234);
nand U44905 (N_44905,N_36601,N_37790);
nand U44906 (N_44906,N_34222,N_37290);
or U44907 (N_44907,N_31584,N_36386);
nor U44908 (N_44908,N_38730,N_38737);
and U44909 (N_44909,N_39500,N_30022);
or U44910 (N_44910,N_31829,N_34856);
and U44911 (N_44911,N_30050,N_39089);
and U44912 (N_44912,N_37840,N_38390);
nor U44913 (N_44913,N_30580,N_36034);
nor U44914 (N_44914,N_38157,N_35033);
xnor U44915 (N_44915,N_36424,N_39767);
and U44916 (N_44916,N_37675,N_36575);
and U44917 (N_44917,N_34508,N_34651);
and U44918 (N_44918,N_37443,N_35968);
nand U44919 (N_44919,N_36309,N_34875);
or U44920 (N_44920,N_32861,N_32032);
xor U44921 (N_44921,N_34199,N_36846);
and U44922 (N_44922,N_35319,N_36200);
or U44923 (N_44923,N_34307,N_34575);
or U44924 (N_44924,N_33850,N_33573);
and U44925 (N_44925,N_33154,N_36326);
nand U44926 (N_44926,N_37310,N_38548);
xnor U44927 (N_44927,N_32682,N_30575);
nand U44928 (N_44928,N_32717,N_30789);
or U44929 (N_44929,N_36275,N_33675);
xnor U44930 (N_44930,N_31011,N_34634);
or U44931 (N_44931,N_30102,N_33055);
or U44932 (N_44932,N_39400,N_34568);
xnor U44933 (N_44933,N_38905,N_38884);
nor U44934 (N_44934,N_34949,N_39451);
or U44935 (N_44935,N_33278,N_30698);
xnor U44936 (N_44936,N_32950,N_33889);
nor U44937 (N_44937,N_32628,N_32625);
xnor U44938 (N_44938,N_33808,N_31872);
or U44939 (N_44939,N_34304,N_35298);
xor U44940 (N_44940,N_34133,N_34124);
xor U44941 (N_44941,N_31912,N_37933);
or U44942 (N_44942,N_32617,N_32299);
xor U44943 (N_44943,N_34054,N_39506);
xnor U44944 (N_44944,N_31138,N_38827);
xor U44945 (N_44945,N_37867,N_38844);
nand U44946 (N_44946,N_39887,N_39718);
xor U44947 (N_44947,N_31167,N_36198);
nor U44948 (N_44948,N_30302,N_36320);
nor U44949 (N_44949,N_31364,N_34560);
and U44950 (N_44950,N_38679,N_36826);
nand U44951 (N_44951,N_38575,N_39873);
nand U44952 (N_44952,N_34603,N_38480);
and U44953 (N_44953,N_37817,N_37490);
or U44954 (N_44954,N_37776,N_37383);
nor U44955 (N_44955,N_35340,N_36675);
xor U44956 (N_44956,N_38559,N_33347);
nand U44957 (N_44957,N_32351,N_30770);
nand U44958 (N_44958,N_36685,N_30212);
and U44959 (N_44959,N_33625,N_32403);
and U44960 (N_44960,N_31857,N_38100);
or U44961 (N_44961,N_39674,N_39939);
xor U44962 (N_44962,N_33570,N_31178);
and U44963 (N_44963,N_38621,N_31233);
and U44964 (N_44964,N_34536,N_31470);
or U44965 (N_44965,N_31437,N_31353);
or U44966 (N_44966,N_39034,N_30165);
nand U44967 (N_44967,N_35302,N_34105);
xnor U44968 (N_44968,N_32948,N_35608);
and U44969 (N_44969,N_39799,N_37072);
xnor U44970 (N_44970,N_30390,N_38839);
and U44971 (N_44971,N_35777,N_37297);
xor U44972 (N_44972,N_31345,N_35058);
nand U44973 (N_44973,N_36397,N_36676);
nand U44974 (N_44974,N_36714,N_30784);
nor U44975 (N_44975,N_36012,N_30445);
xor U44976 (N_44976,N_30673,N_36266);
xor U44977 (N_44977,N_36372,N_36578);
and U44978 (N_44978,N_35753,N_34846);
nand U44979 (N_44979,N_38995,N_33672);
nor U44980 (N_44980,N_36272,N_38510);
nor U44981 (N_44981,N_37638,N_34241);
nand U44982 (N_44982,N_36907,N_33547);
nor U44983 (N_44983,N_35273,N_36291);
or U44984 (N_44984,N_36210,N_38153);
and U44985 (N_44985,N_34234,N_38152);
or U44986 (N_44986,N_37409,N_38681);
nand U44987 (N_44987,N_39634,N_32147);
nand U44988 (N_44988,N_30823,N_38985);
xnor U44989 (N_44989,N_31914,N_32120);
and U44990 (N_44990,N_36658,N_34148);
nand U44991 (N_44991,N_30568,N_32000);
and U44992 (N_44992,N_34439,N_31263);
nor U44993 (N_44993,N_38765,N_38054);
xnor U44994 (N_44994,N_37159,N_31946);
xor U44995 (N_44995,N_38408,N_35359);
or U44996 (N_44996,N_38669,N_34710);
xor U44997 (N_44997,N_35498,N_38640);
xor U44998 (N_44998,N_37431,N_35391);
or U44999 (N_44999,N_30183,N_36635);
nor U45000 (N_45000,N_35264,N_37509);
nor U45001 (N_45001,N_33488,N_30671);
or U45002 (N_45002,N_33524,N_30736);
and U45003 (N_45003,N_39378,N_31528);
nor U45004 (N_45004,N_36659,N_31650);
nor U45005 (N_45005,N_31427,N_37288);
or U45006 (N_45006,N_36698,N_33939);
or U45007 (N_45007,N_35678,N_31013);
nand U45008 (N_45008,N_38617,N_38153);
nand U45009 (N_45009,N_37550,N_35815);
nor U45010 (N_45010,N_39067,N_35031);
or U45011 (N_45011,N_37261,N_36252);
nor U45012 (N_45012,N_30221,N_37447);
and U45013 (N_45013,N_33856,N_35634);
nor U45014 (N_45014,N_38570,N_33608);
xor U45015 (N_45015,N_32654,N_32894);
nand U45016 (N_45016,N_31436,N_37138);
or U45017 (N_45017,N_37300,N_37590);
nor U45018 (N_45018,N_30897,N_31980);
xor U45019 (N_45019,N_32455,N_30634);
nor U45020 (N_45020,N_30807,N_36016);
nor U45021 (N_45021,N_30544,N_33634);
and U45022 (N_45022,N_32223,N_39540);
xnor U45023 (N_45023,N_39592,N_38373);
and U45024 (N_45024,N_31339,N_33261);
nor U45025 (N_45025,N_37852,N_33561);
nand U45026 (N_45026,N_38645,N_30568);
and U45027 (N_45027,N_38750,N_33433);
nand U45028 (N_45028,N_39943,N_34908);
nor U45029 (N_45029,N_31065,N_35912);
nand U45030 (N_45030,N_38684,N_38902);
nor U45031 (N_45031,N_30237,N_30337);
nand U45032 (N_45032,N_31616,N_36433);
and U45033 (N_45033,N_36446,N_36165);
or U45034 (N_45034,N_30032,N_30140);
and U45035 (N_45035,N_30759,N_36569);
nand U45036 (N_45036,N_32731,N_38349);
and U45037 (N_45037,N_39137,N_33281);
and U45038 (N_45038,N_30703,N_34284);
xor U45039 (N_45039,N_33625,N_33376);
nor U45040 (N_45040,N_35705,N_32232);
or U45041 (N_45041,N_36322,N_31056);
and U45042 (N_45042,N_36020,N_35323);
nor U45043 (N_45043,N_30944,N_30835);
xnor U45044 (N_45044,N_30044,N_38622);
and U45045 (N_45045,N_33876,N_32437);
and U45046 (N_45046,N_38147,N_33692);
nand U45047 (N_45047,N_38067,N_34525);
nand U45048 (N_45048,N_38229,N_38677);
nand U45049 (N_45049,N_36590,N_38791);
and U45050 (N_45050,N_37368,N_33052);
and U45051 (N_45051,N_32518,N_33549);
nor U45052 (N_45052,N_33216,N_39151);
nand U45053 (N_45053,N_33651,N_38483);
or U45054 (N_45054,N_37291,N_33543);
xor U45055 (N_45055,N_37948,N_30566);
and U45056 (N_45056,N_36304,N_30941);
xor U45057 (N_45057,N_30284,N_30659);
or U45058 (N_45058,N_36121,N_35524);
xor U45059 (N_45059,N_34807,N_39452);
nand U45060 (N_45060,N_36982,N_33794);
nor U45061 (N_45061,N_36097,N_39233);
xnor U45062 (N_45062,N_31313,N_38130);
nor U45063 (N_45063,N_39074,N_38350);
nand U45064 (N_45064,N_32622,N_31678);
xnor U45065 (N_45065,N_38186,N_37575);
or U45066 (N_45066,N_34921,N_30713);
and U45067 (N_45067,N_34989,N_37694);
or U45068 (N_45068,N_30157,N_39601);
nor U45069 (N_45069,N_34924,N_32948);
xnor U45070 (N_45070,N_36203,N_39727);
or U45071 (N_45071,N_37663,N_34575);
or U45072 (N_45072,N_30978,N_35350);
or U45073 (N_45073,N_33207,N_30042);
nor U45074 (N_45074,N_32145,N_39896);
xnor U45075 (N_45075,N_33940,N_33406);
nand U45076 (N_45076,N_37359,N_31441);
nor U45077 (N_45077,N_31598,N_38257);
xor U45078 (N_45078,N_34037,N_33176);
nand U45079 (N_45079,N_32914,N_36932);
and U45080 (N_45080,N_30806,N_33513);
or U45081 (N_45081,N_35430,N_31517);
and U45082 (N_45082,N_35637,N_33530);
xnor U45083 (N_45083,N_30475,N_36728);
nand U45084 (N_45084,N_36369,N_31292);
and U45085 (N_45085,N_35327,N_31537);
nor U45086 (N_45086,N_35277,N_39543);
or U45087 (N_45087,N_35767,N_31576);
nand U45088 (N_45088,N_39298,N_31006);
xnor U45089 (N_45089,N_33925,N_31007);
nand U45090 (N_45090,N_39262,N_35064);
or U45091 (N_45091,N_34955,N_39051);
nand U45092 (N_45092,N_36892,N_39692);
and U45093 (N_45093,N_33501,N_30278);
xnor U45094 (N_45094,N_30803,N_37701);
and U45095 (N_45095,N_37522,N_37396);
or U45096 (N_45096,N_37964,N_35597);
nand U45097 (N_45097,N_32330,N_31689);
xor U45098 (N_45098,N_32037,N_38710);
nor U45099 (N_45099,N_35019,N_34056);
and U45100 (N_45100,N_31526,N_31995);
or U45101 (N_45101,N_30334,N_34643);
nor U45102 (N_45102,N_33890,N_35183);
and U45103 (N_45103,N_34358,N_39420);
and U45104 (N_45104,N_38116,N_39918);
xnor U45105 (N_45105,N_34691,N_32692);
nand U45106 (N_45106,N_33774,N_32799);
xnor U45107 (N_45107,N_36211,N_35703);
or U45108 (N_45108,N_35834,N_35900);
nor U45109 (N_45109,N_37618,N_30366);
or U45110 (N_45110,N_33509,N_37959);
nand U45111 (N_45111,N_39183,N_37981);
and U45112 (N_45112,N_38817,N_30490);
nor U45113 (N_45113,N_38875,N_36602);
nand U45114 (N_45114,N_39992,N_34685);
nand U45115 (N_45115,N_35311,N_35160);
nor U45116 (N_45116,N_38478,N_34217);
xor U45117 (N_45117,N_39561,N_36375);
nand U45118 (N_45118,N_32496,N_31652);
or U45119 (N_45119,N_36149,N_35610);
xor U45120 (N_45120,N_37660,N_31598);
and U45121 (N_45121,N_32880,N_32434);
nand U45122 (N_45122,N_37731,N_38483);
nor U45123 (N_45123,N_34534,N_34623);
nand U45124 (N_45124,N_37561,N_38304);
xnor U45125 (N_45125,N_37641,N_34598);
or U45126 (N_45126,N_35898,N_34158);
or U45127 (N_45127,N_32761,N_38272);
or U45128 (N_45128,N_38433,N_30198);
nand U45129 (N_45129,N_36133,N_39643);
nor U45130 (N_45130,N_32986,N_33388);
nand U45131 (N_45131,N_35937,N_32476);
xor U45132 (N_45132,N_31538,N_39710);
xor U45133 (N_45133,N_39928,N_34605);
and U45134 (N_45134,N_38495,N_32854);
xor U45135 (N_45135,N_32512,N_32828);
and U45136 (N_45136,N_38662,N_33581);
nor U45137 (N_45137,N_37271,N_37322);
nor U45138 (N_45138,N_37392,N_36293);
xnor U45139 (N_45139,N_37619,N_35633);
nand U45140 (N_45140,N_33449,N_36841);
xnor U45141 (N_45141,N_30631,N_30469);
nor U45142 (N_45142,N_31339,N_39981);
nand U45143 (N_45143,N_38966,N_38190);
or U45144 (N_45144,N_39310,N_32802);
and U45145 (N_45145,N_36627,N_35465);
and U45146 (N_45146,N_33680,N_34429);
and U45147 (N_45147,N_32279,N_31927);
nand U45148 (N_45148,N_33201,N_30164);
nor U45149 (N_45149,N_39462,N_38008);
and U45150 (N_45150,N_39699,N_32963);
or U45151 (N_45151,N_30125,N_33373);
nor U45152 (N_45152,N_34394,N_36752);
or U45153 (N_45153,N_30707,N_33275);
nand U45154 (N_45154,N_37737,N_35052);
or U45155 (N_45155,N_32696,N_39949);
and U45156 (N_45156,N_32931,N_35551);
nand U45157 (N_45157,N_32934,N_35251);
nor U45158 (N_45158,N_38420,N_33499);
nor U45159 (N_45159,N_35855,N_36329);
and U45160 (N_45160,N_35600,N_31351);
and U45161 (N_45161,N_34926,N_35867);
nor U45162 (N_45162,N_39099,N_32931);
or U45163 (N_45163,N_36627,N_38584);
xor U45164 (N_45164,N_30364,N_34786);
nor U45165 (N_45165,N_31162,N_36786);
xor U45166 (N_45166,N_32352,N_37331);
nor U45167 (N_45167,N_30468,N_33297);
nor U45168 (N_45168,N_37684,N_35077);
nand U45169 (N_45169,N_34365,N_37408);
xnor U45170 (N_45170,N_37785,N_32869);
nand U45171 (N_45171,N_33954,N_31768);
nand U45172 (N_45172,N_35136,N_35642);
and U45173 (N_45173,N_35161,N_30009);
and U45174 (N_45174,N_38810,N_30352);
xnor U45175 (N_45175,N_30926,N_32326);
and U45176 (N_45176,N_30607,N_31841);
and U45177 (N_45177,N_37709,N_32744);
nand U45178 (N_45178,N_31366,N_35741);
nand U45179 (N_45179,N_31322,N_33883);
nand U45180 (N_45180,N_38524,N_38512);
xnor U45181 (N_45181,N_38422,N_30747);
or U45182 (N_45182,N_37838,N_34194);
nand U45183 (N_45183,N_37588,N_33378);
or U45184 (N_45184,N_32721,N_33775);
nor U45185 (N_45185,N_36373,N_37040);
xnor U45186 (N_45186,N_37013,N_36403);
nand U45187 (N_45187,N_39177,N_39374);
xor U45188 (N_45188,N_39939,N_30414);
nor U45189 (N_45189,N_32566,N_39711);
nor U45190 (N_45190,N_38652,N_38724);
and U45191 (N_45191,N_34201,N_31047);
nor U45192 (N_45192,N_30726,N_30097);
and U45193 (N_45193,N_30206,N_36007);
nor U45194 (N_45194,N_33758,N_32272);
or U45195 (N_45195,N_34578,N_31951);
and U45196 (N_45196,N_34448,N_35146);
nor U45197 (N_45197,N_32712,N_37614);
and U45198 (N_45198,N_36244,N_35972);
and U45199 (N_45199,N_36129,N_37934);
nor U45200 (N_45200,N_38562,N_39337);
nor U45201 (N_45201,N_39863,N_34196);
nor U45202 (N_45202,N_33411,N_38563);
nand U45203 (N_45203,N_35957,N_31671);
or U45204 (N_45204,N_36896,N_33800);
and U45205 (N_45205,N_35452,N_33623);
nand U45206 (N_45206,N_30328,N_30013);
nor U45207 (N_45207,N_36434,N_37163);
and U45208 (N_45208,N_33741,N_32847);
and U45209 (N_45209,N_34263,N_31875);
xor U45210 (N_45210,N_34531,N_35193);
or U45211 (N_45211,N_33098,N_30875);
nor U45212 (N_45212,N_30758,N_31686);
xnor U45213 (N_45213,N_37717,N_31007);
or U45214 (N_45214,N_36257,N_33109);
nor U45215 (N_45215,N_33552,N_30709);
or U45216 (N_45216,N_32559,N_37732);
xor U45217 (N_45217,N_31824,N_38456);
nand U45218 (N_45218,N_35151,N_38131);
nor U45219 (N_45219,N_33518,N_32340);
nand U45220 (N_45220,N_35510,N_38419);
nand U45221 (N_45221,N_34075,N_32454);
nand U45222 (N_45222,N_37178,N_39919);
or U45223 (N_45223,N_31389,N_36523);
nor U45224 (N_45224,N_35219,N_35775);
xor U45225 (N_45225,N_31453,N_30224);
xor U45226 (N_45226,N_30023,N_37859);
xor U45227 (N_45227,N_30212,N_34462);
nand U45228 (N_45228,N_31495,N_39022);
nor U45229 (N_45229,N_32712,N_37931);
nor U45230 (N_45230,N_31493,N_33431);
and U45231 (N_45231,N_38073,N_34829);
and U45232 (N_45232,N_39549,N_31962);
or U45233 (N_45233,N_37789,N_38173);
and U45234 (N_45234,N_31117,N_33218);
nor U45235 (N_45235,N_30682,N_35705);
xor U45236 (N_45236,N_31738,N_30356);
nor U45237 (N_45237,N_37727,N_39725);
nor U45238 (N_45238,N_30970,N_37647);
nand U45239 (N_45239,N_36872,N_32274);
and U45240 (N_45240,N_35648,N_36567);
or U45241 (N_45241,N_30341,N_36789);
nor U45242 (N_45242,N_30282,N_34528);
or U45243 (N_45243,N_31015,N_39374);
or U45244 (N_45244,N_32003,N_32575);
nand U45245 (N_45245,N_35690,N_32424);
and U45246 (N_45246,N_34983,N_33895);
or U45247 (N_45247,N_31948,N_37914);
xnor U45248 (N_45248,N_32603,N_30217);
nor U45249 (N_45249,N_36024,N_30415);
and U45250 (N_45250,N_35033,N_30339);
and U45251 (N_45251,N_37388,N_35262);
or U45252 (N_45252,N_30052,N_30974);
and U45253 (N_45253,N_39066,N_30241);
xor U45254 (N_45254,N_35857,N_34780);
nand U45255 (N_45255,N_33250,N_34945);
nor U45256 (N_45256,N_32978,N_30120);
and U45257 (N_45257,N_39398,N_36186);
and U45258 (N_45258,N_33639,N_30799);
nand U45259 (N_45259,N_31796,N_37056);
nor U45260 (N_45260,N_35099,N_36005);
nor U45261 (N_45261,N_34917,N_34643);
nor U45262 (N_45262,N_30203,N_32403);
or U45263 (N_45263,N_39440,N_39332);
or U45264 (N_45264,N_33511,N_32526);
xor U45265 (N_45265,N_35445,N_36681);
nand U45266 (N_45266,N_34491,N_30483);
xnor U45267 (N_45267,N_37114,N_36275);
and U45268 (N_45268,N_31335,N_35222);
and U45269 (N_45269,N_31617,N_33346);
and U45270 (N_45270,N_33273,N_30914);
nand U45271 (N_45271,N_32577,N_31758);
xor U45272 (N_45272,N_37894,N_31574);
nand U45273 (N_45273,N_30590,N_39532);
nand U45274 (N_45274,N_38208,N_36796);
nand U45275 (N_45275,N_32620,N_36647);
and U45276 (N_45276,N_32836,N_35446);
and U45277 (N_45277,N_33867,N_33562);
xnor U45278 (N_45278,N_30240,N_37911);
xnor U45279 (N_45279,N_32128,N_30490);
nor U45280 (N_45280,N_32132,N_34648);
and U45281 (N_45281,N_32146,N_37111);
or U45282 (N_45282,N_37644,N_33852);
or U45283 (N_45283,N_37744,N_34416);
xor U45284 (N_45284,N_35369,N_37154);
nand U45285 (N_45285,N_38179,N_36361);
xnor U45286 (N_45286,N_39792,N_34912);
nor U45287 (N_45287,N_38812,N_33438);
nor U45288 (N_45288,N_36052,N_33308);
and U45289 (N_45289,N_31004,N_33508);
or U45290 (N_45290,N_36708,N_35468);
or U45291 (N_45291,N_39073,N_31546);
nand U45292 (N_45292,N_32648,N_39223);
or U45293 (N_45293,N_31510,N_30221);
and U45294 (N_45294,N_30475,N_36932);
and U45295 (N_45295,N_39366,N_37186);
xor U45296 (N_45296,N_35603,N_33772);
or U45297 (N_45297,N_36183,N_38586);
and U45298 (N_45298,N_39764,N_36372);
or U45299 (N_45299,N_31441,N_35021);
nor U45300 (N_45300,N_30381,N_37759);
and U45301 (N_45301,N_39364,N_39297);
xnor U45302 (N_45302,N_31216,N_33970);
nand U45303 (N_45303,N_35497,N_32115);
and U45304 (N_45304,N_33616,N_39458);
and U45305 (N_45305,N_38720,N_33884);
or U45306 (N_45306,N_36695,N_30365);
xor U45307 (N_45307,N_32952,N_35038);
and U45308 (N_45308,N_32364,N_33479);
xnor U45309 (N_45309,N_35234,N_36092);
nor U45310 (N_45310,N_39320,N_32076);
nor U45311 (N_45311,N_37014,N_39797);
xnor U45312 (N_45312,N_38575,N_30023);
or U45313 (N_45313,N_33014,N_31495);
nor U45314 (N_45314,N_30184,N_32109);
and U45315 (N_45315,N_36204,N_39213);
or U45316 (N_45316,N_36055,N_32545);
nor U45317 (N_45317,N_34650,N_38309);
nand U45318 (N_45318,N_35286,N_39753);
nor U45319 (N_45319,N_33502,N_33649);
or U45320 (N_45320,N_38741,N_39243);
nand U45321 (N_45321,N_32755,N_35399);
nand U45322 (N_45322,N_33840,N_32158);
and U45323 (N_45323,N_35973,N_33800);
xor U45324 (N_45324,N_36018,N_39626);
nor U45325 (N_45325,N_36988,N_36533);
nand U45326 (N_45326,N_37737,N_35279);
xnor U45327 (N_45327,N_36217,N_38936);
nor U45328 (N_45328,N_38860,N_36160);
nand U45329 (N_45329,N_38693,N_36121);
or U45330 (N_45330,N_34421,N_35657);
nor U45331 (N_45331,N_34916,N_39353);
or U45332 (N_45332,N_34817,N_36571);
nand U45333 (N_45333,N_37417,N_31758);
nand U45334 (N_45334,N_38613,N_32532);
xnor U45335 (N_45335,N_39828,N_36694);
nor U45336 (N_45336,N_36041,N_30799);
xor U45337 (N_45337,N_38230,N_34207);
or U45338 (N_45338,N_39388,N_37382);
nand U45339 (N_45339,N_39570,N_34725);
and U45340 (N_45340,N_30198,N_32956);
nand U45341 (N_45341,N_36855,N_39536);
nand U45342 (N_45342,N_38104,N_39608);
nand U45343 (N_45343,N_32329,N_31435);
and U45344 (N_45344,N_34304,N_35195);
xor U45345 (N_45345,N_31828,N_39355);
nor U45346 (N_45346,N_37961,N_34414);
nor U45347 (N_45347,N_39880,N_31915);
nor U45348 (N_45348,N_34290,N_36678);
and U45349 (N_45349,N_30173,N_36465);
and U45350 (N_45350,N_31650,N_35692);
nand U45351 (N_45351,N_37402,N_35099);
nor U45352 (N_45352,N_36655,N_31333);
nand U45353 (N_45353,N_32789,N_30007);
or U45354 (N_45354,N_35848,N_30657);
nand U45355 (N_45355,N_39841,N_33580);
xor U45356 (N_45356,N_30109,N_30257);
nor U45357 (N_45357,N_38955,N_35035);
and U45358 (N_45358,N_30661,N_34537);
nand U45359 (N_45359,N_36035,N_37958);
or U45360 (N_45360,N_38410,N_35751);
xor U45361 (N_45361,N_32655,N_33856);
xor U45362 (N_45362,N_35284,N_35462);
nand U45363 (N_45363,N_31011,N_36636);
or U45364 (N_45364,N_35491,N_36158);
or U45365 (N_45365,N_33403,N_39944);
nor U45366 (N_45366,N_38669,N_31533);
and U45367 (N_45367,N_38990,N_30645);
nand U45368 (N_45368,N_39458,N_35643);
and U45369 (N_45369,N_30339,N_34222);
or U45370 (N_45370,N_37070,N_39921);
or U45371 (N_45371,N_37313,N_37997);
xnor U45372 (N_45372,N_38842,N_33469);
or U45373 (N_45373,N_32315,N_30871);
nor U45374 (N_45374,N_37067,N_37646);
nor U45375 (N_45375,N_34142,N_37009);
nor U45376 (N_45376,N_31213,N_34448);
nor U45377 (N_45377,N_31091,N_36442);
nand U45378 (N_45378,N_39585,N_33364);
and U45379 (N_45379,N_36061,N_31303);
or U45380 (N_45380,N_39812,N_39416);
nor U45381 (N_45381,N_39813,N_32609);
nand U45382 (N_45382,N_35584,N_32679);
or U45383 (N_45383,N_31114,N_36887);
nor U45384 (N_45384,N_38868,N_34933);
and U45385 (N_45385,N_38735,N_31409);
or U45386 (N_45386,N_39980,N_37717);
and U45387 (N_45387,N_38814,N_30524);
nor U45388 (N_45388,N_39604,N_30255);
or U45389 (N_45389,N_37661,N_33998);
xor U45390 (N_45390,N_35353,N_35450);
or U45391 (N_45391,N_34724,N_37690);
nor U45392 (N_45392,N_30130,N_35160);
nand U45393 (N_45393,N_35186,N_31962);
nor U45394 (N_45394,N_35782,N_39858);
nor U45395 (N_45395,N_34143,N_32599);
nor U45396 (N_45396,N_33389,N_37424);
xor U45397 (N_45397,N_33689,N_31412);
xnor U45398 (N_45398,N_37457,N_39435);
and U45399 (N_45399,N_36548,N_31492);
and U45400 (N_45400,N_32423,N_35719);
nor U45401 (N_45401,N_35341,N_34457);
and U45402 (N_45402,N_39863,N_35037);
and U45403 (N_45403,N_32020,N_36552);
xor U45404 (N_45404,N_34168,N_32287);
or U45405 (N_45405,N_38881,N_34326);
or U45406 (N_45406,N_37071,N_33769);
or U45407 (N_45407,N_38881,N_33261);
nor U45408 (N_45408,N_36042,N_32740);
xnor U45409 (N_45409,N_37735,N_34569);
and U45410 (N_45410,N_31094,N_32743);
or U45411 (N_45411,N_38698,N_37810);
xor U45412 (N_45412,N_35071,N_37671);
xnor U45413 (N_45413,N_37024,N_38264);
xor U45414 (N_45414,N_38500,N_36532);
xnor U45415 (N_45415,N_30880,N_37285);
and U45416 (N_45416,N_30968,N_33143);
or U45417 (N_45417,N_38066,N_32074);
and U45418 (N_45418,N_30146,N_33210);
xnor U45419 (N_45419,N_33967,N_36953);
and U45420 (N_45420,N_35568,N_37138);
nor U45421 (N_45421,N_35775,N_39782);
xnor U45422 (N_45422,N_37563,N_30980);
nor U45423 (N_45423,N_37651,N_38831);
xnor U45424 (N_45424,N_30354,N_38513);
nand U45425 (N_45425,N_35465,N_37715);
and U45426 (N_45426,N_39159,N_30378);
xnor U45427 (N_45427,N_37928,N_34672);
nand U45428 (N_45428,N_36127,N_30101);
xnor U45429 (N_45429,N_39672,N_34110);
nand U45430 (N_45430,N_39370,N_30245);
and U45431 (N_45431,N_37267,N_32068);
nand U45432 (N_45432,N_33347,N_31730);
and U45433 (N_45433,N_33370,N_35607);
xnor U45434 (N_45434,N_35906,N_32926);
and U45435 (N_45435,N_32810,N_39181);
nand U45436 (N_45436,N_37480,N_30425);
nor U45437 (N_45437,N_32045,N_33528);
nand U45438 (N_45438,N_32018,N_31416);
xor U45439 (N_45439,N_37749,N_39563);
nor U45440 (N_45440,N_39038,N_37020);
or U45441 (N_45441,N_39893,N_32877);
or U45442 (N_45442,N_31155,N_33838);
or U45443 (N_45443,N_31370,N_33565);
nor U45444 (N_45444,N_39038,N_33581);
or U45445 (N_45445,N_34868,N_32696);
xor U45446 (N_45446,N_37569,N_34283);
nand U45447 (N_45447,N_34097,N_33294);
or U45448 (N_45448,N_32228,N_39558);
and U45449 (N_45449,N_34691,N_32981);
xor U45450 (N_45450,N_37623,N_32512);
nor U45451 (N_45451,N_31830,N_37247);
xor U45452 (N_45452,N_36931,N_37265);
or U45453 (N_45453,N_37574,N_30340);
or U45454 (N_45454,N_31416,N_37470);
xor U45455 (N_45455,N_38962,N_32388);
or U45456 (N_45456,N_35228,N_30851);
nand U45457 (N_45457,N_34489,N_36260);
nor U45458 (N_45458,N_33798,N_36163);
and U45459 (N_45459,N_33198,N_31381);
nor U45460 (N_45460,N_34445,N_30888);
and U45461 (N_45461,N_34896,N_35319);
and U45462 (N_45462,N_37961,N_38566);
or U45463 (N_45463,N_32958,N_36939);
and U45464 (N_45464,N_30059,N_36953);
nand U45465 (N_45465,N_36243,N_38899);
nor U45466 (N_45466,N_32460,N_37046);
or U45467 (N_45467,N_38428,N_31159);
nor U45468 (N_45468,N_35111,N_31768);
xnor U45469 (N_45469,N_32776,N_34192);
nor U45470 (N_45470,N_39117,N_35397);
and U45471 (N_45471,N_34628,N_32539);
nor U45472 (N_45472,N_32553,N_39590);
and U45473 (N_45473,N_36440,N_39464);
xnor U45474 (N_45474,N_32176,N_36639);
xnor U45475 (N_45475,N_37280,N_34626);
and U45476 (N_45476,N_39155,N_30706);
nor U45477 (N_45477,N_30830,N_38531);
nor U45478 (N_45478,N_33581,N_37365);
xnor U45479 (N_45479,N_38059,N_37657);
nor U45480 (N_45480,N_34753,N_39680);
nand U45481 (N_45481,N_33129,N_37612);
or U45482 (N_45482,N_32689,N_30596);
nor U45483 (N_45483,N_33845,N_30886);
nor U45484 (N_45484,N_34435,N_39827);
and U45485 (N_45485,N_38447,N_37827);
xnor U45486 (N_45486,N_31135,N_33274);
nor U45487 (N_45487,N_33636,N_32130);
nand U45488 (N_45488,N_31812,N_33283);
or U45489 (N_45489,N_30800,N_30598);
and U45490 (N_45490,N_31043,N_32145);
nor U45491 (N_45491,N_34157,N_35274);
xor U45492 (N_45492,N_34537,N_39587);
and U45493 (N_45493,N_38608,N_34339);
and U45494 (N_45494,N_35422,N_31716);
and U45495 (N_45495,N_35260,N_37245);
nor U45496 (N_45496,N_33548,N_30797);
and U45497 (N_45497,N_33236,N_31386);
xnor U45498 (N_45498,N_36116,N_34143);
nand U45499 (N_45499,N_32215,N_31606);
or U45500 (N_45500,N_33488,N_37617);
nor U45501 (N_45501,N_37569,N_34947);
nor U45502 (N_45502,N_31554,N_35863);
xnor U45503 (N_45503,N_32723,N_36897);
or U45504 (N_45504,N_31966,N_36757);
or U45505 (N_45505,N_34609,N_34924);
nor U45506 (N_45506,N_38471,N_30199);
and U45507 (N_45507,N_33794,N_38466);
or U45508 (N_45508,N_35144,N_31771);
or U45509 (N_45509,N_34537,N_34338);
and U45510 (N_45510,N_33965,N_36229);
or U45511 (N_45511,N_35710,N_37542);
nor U45512 (N_45512,N_32680,N_30765);
xor U45513 (N_45513,N_36623,N_32915);
nor U45514 (N_45514,N_39690,N_30553);
nor U45515 (N_45515,N_35080,N_36210);
nand U45516 (N_45516,N_33946,N_34472);
xor U45517 (N_45517,N_34121,N_30226);
and U45518 (N_45518,N_39742,N_39478);
nor U45519 (N_45519,N_36179,N_36620);
and U45520 (N_45520,N_30443,N_37224);
xor U45521 (N_45521,N_37909,N_37628);
nor U45522 (N_45522,N_30860,N_35094);
nor U45523 (N_45523,N_34050,N_39721);
and U45524 (N_45524,N_38815,N_37268);
or U45525 (N_45525,N_31177,N_31256);
and U45526 (N_45526,N_30708,N_32113);
xnor U45527 (N_45527,N_36891,N_33917);
xnor U45528 (N_45528,N_35490,N_32181);
or U45529 (N_45529,N_32050,N_39472);
nor U45530 (N_45530,N_31391,N_34206);
or U45531 (N_45531,N_32240,N_34116);
or U45532 (N_45532,N_38258,N_34450);
nand U45533 (N_45533,N_32070,N_34829);
or U45534 (N_45534,N_36085,N_39164);
or U45535 (N_45535,N_30385,N_35349);
nand U45536 (N_45536,N_37406,N_30683);
nand U45537 (N_45537,N_34223,N_37593);
xor U45538 (N_45538,N_39906,N_32383);
nor U45539 (N_45539,N_37221,N_37212);
and U45540 (N_45540,N_37870,N_35048);
and U45541 (N_45541,N_37107,N_39460);
and U45542 (N_45542,N_35927,N_33783);
xnor U45543 (N_45543,N_31684,N_35284);
and U45544 (N_45544,N_39675,N_36612);
nand U45545 (N_45545,N_33386,N_31386);
nor U45546 (N_45546,N_38852,N_38080);
nand U45547 (N_45547,N_32606,N_32835);
xor U45548 (N_45548,N_38512,N_34083);
xnor U45549 (N_45549,N_32799,N_38504);
nor U45550 (N_45550,N_37829,N_37803);
or U45551 (N_45551,N_39233,N_35384);
nand U45552 (N_45552,N_37863,N_33307);
nand U45553 (N_45553,N_39458,N_34114);
xnor U45554 (N_45554,N_32594,N_32645);
or U45555 (N_45555,N_35515,N_32175);
nor U45556 (N_45556,N_39659,N_38027);
and U45557 (N_45557,N_34110,N_36332);
nand U45558 (N_45558,N_39842,N_33834);
nor U45559 (N_45559,N_38742,N_39910);
and U45560 (N_45560,N_39388,N_30071);
or U45561 (N_45561,N_38147,N_34180);
nand U45562 (N_45562,N_34087,N_36828);
and U45563 (N_45563,N_36867,N_33056);
or U45564 (N_45564,N_34676,N_31538);
nand U45565 (N_45565,N_30198,N_35459);
xor U45566 (N_45566,N_37029,N_31804);
or U45567 (N_45567,N_31464,N_31107);
nand U45568 (N_45568,N_37381,N_33886);
nor U45569 (N_45569,N_37998,N_39501);
xnor U45570 (N_45570,N_36343,N_32275);
or U45571 (N_45571,N_32083,N_35244);
nor U45572 (N_45572,N_39563,N_37813);
nand U45573 (N_45573,N_31722,N_39528);
and U45574 (N_45574,N_34009,N_31389);
and U45575 (N_45575,N_30807,N_33867);
nor U45576 (N_45576,N_32609,N_35176);
or U45577 (N_45577,N_31288,N_37640);
xnor U45578 (N_45578,N_38735,N_37074);
and U45579 (N_45579,N_30546,N_30469);
nand U45580 (N_45580,N_36411,N_33521);
nor U45581 (N_45581,N_39161,N_38047);
nor U45582 (N_45582,N_30563,N_36281);
nor U45583 (N_45583,N_33284,N_35121);
nor U45584 (N_45584,N_30200,N_33614);
nand U45585 (N_45585,N_34593,N_37768);
nor U45586 (N_45586,N_36656,N_37661);
nand U45587 (N_45587,N_30809,N_33078);
nand U45588 (N_45588,N_32972,N_34895);
nor U45589 (N_45589,N_33384,N_38373);
and U45590 (N_45590,N_38923,N_32107);
and U45591 (N_45591,N_31957,N_32324);
or U45592 (N_45592,N_33606,N_37397);
nor U45593 (N_45593,N_31779,N_36349);
nor U45594 (N_45594,N_38523,N_30814);
xnor U45595 (N_45595,N_32341,N_31474);
and U45596 (N_45596,N_36599,N_34150);
nand U45597 (N_45597,N_38126,N_37931);
nand U45598 (N_45598,N_38148,N_39623);
and U45599 (N_45599,N_31628,N_38175);
or U45600 (N_45600,N_36568,N_34892);
or U45601 (N_45601,N_31811,N_39439);
xor U45602 (N_45602,N_35735,N_33911);
nand U45603 (N_45603,N_34479,N_33887);
and U45604 (N_45604,N_38783,N_30747);
xor U45605 (N_45605,N_38700,N_37288);
xor U45606 (N_45606,N_34833,N_36955);
and U45607 (N_45607,N_30882,N_33057);
nand U45608 (N_45608,N_30248,N_37154);
nor U45609 (N_45609,N_37992,N_36943);
xnor U45610 (N_45610,N_36497,N_37008);
nor U45611 (N_45611,N_33840,N_30039);
and U45612 (N_45612,N_32760,N_36803);
xnor U45613 (N_45613,N_36837,N_31012);
or U45614 (N_45614,N_31837,N_38460);
nand U45615 (N_45615,N_33738,N_36638);
nand U45616 (N_45616,N_35129,N_31709);
nor U45617 (N_45617,N_36403,N_30788);
nand U45618 (N_45618,N_32359,N_37815);
xnor U45619 (N_45619,N_37371,N_36965);
xnor U45620 (N_45620,N_31056,N_31959);
nor U45621 (N_45621,N_34810,N_33370);
xnor U45622 (N_45622,N_33984,N_39981);
nand U45623 (N_45623,N_34728,N_38213);
nand U45624 (N_45624,N_37294,N_39973);
nor U45625 (N_45625,N_37219,N_38472);
xnor U45626 (N_45626,N_30432,N_33074);
nand U45627 (N_45627,N_35762,N_37656);
nand U45628 (N_45628,N_34766,N_37852);
nor U45629 (N_45629,N_31225,N_32175);
nor U45630 (N_45630,N_31058,N_30891);
nand U45631 (N_45631,N_36126,N_33973);
nand U45632 (N_45632,N_35992,N_30942);
nand U45633 (N_45633,N_32870,N_30149);
xor U45634 (N_45634,N_39367,N_32289);
and U45635 (N_45635,N_33496,N_38862);
xor U45636 (N_45636,N_36506,N_35811);
xnor U45637 (N_45637,N_34462,N_38981);
xor U45638 (N_45638,N_31750,N_31447);
or U45639 (N_45639,N_34457,N_36094);
or U45640 (N_45640,N_30720,N_30959);
nand U45641 (N_45641,N_31450,N_38213);
nand U45642 (N_45642,N_32823,N_38499);
nor U45643 (N_45643,N_38588,N_37292);
or U45644 (N_45644,N_39370,N_34219);
or U45645 (N_45645,N_37572,N_38021);
nor U45646 (N_45646,N_36974,N_32553);
xnor U45647 (N_45647,N_37284,N_30047);
or U45648 (N_45648,N_31363,N_39174);
xor U45649 (N_45649,N_33221,N_37020);
xnor U45650 (N_45650,N_32604,N_35058);
nor U45651 (N_45651,N_33168,N_31756);
xnor U45652 (N_45652,N_35552,N_35520);
nand U45653 (N_45653,N_31844,N_30506);
or U45654 (N_45654,N_36512,N_36564);
nand U45655 (N_45655,N_35625,N_34974);
xnor U45656 (N_45656,N_38793,N_36567);
and U45657 (N_45657,N_30475,N_39455);
and U45658 (N_45658,N_33893,N_38465);
and U45659 (N_45659,N_36581,N_31242);
or U45660 (N_45660,N_31231,N_35499);
nor U45661 (N_45661,N_35688,N_37174);
nor U45662 (N_45662,N_36952,N_35456);
xnor U45663 (N_45663,N_31082,N_38356);
and U45664 (N_45664,N_35533,N_37185);
or U45665 (N_45665,N_32148,N_38969);
and U45666 (N_45666,N_34140,N_33693);
or U45667 (N_45667,N_34300,N_36925);
nor U45668 (N_45668,N_33117,N_39613);
or U45669 (N_45669,N_33058,N_37229);
nor U45670 (N_45670,N_34823,N_35742);
nand U45671 (N_45671,N_39612,N_30275);
or U45672 (N_45672,N_39541,N_32623);
and U45673 (N_45673,N_35882,N_36946);
nand U45674 (N_45674,N_33825,N_36763);
and U45675 (N_45675,N_32133,N_31060);
nor U45676 (N_45676,N_33915,N_36107);
nor U45677 (N_45677,N_34150,N_30161);
and U45678 (N_45678,N_34532,N_38237);
xnor U45679 (N_45679,N_31690,N_31520);
xnor U45680 (N_45680,N_35613,N_37801);
nor U45681 (N_45681,N_39461,N_36598);
nor U45682 (N_45682,N_33947,N_31189);
nand U45683 (N_45683,N_38787,N_35769);
nor U45684 (N_45684,N_39216,N_33330);
nand U45685 (N_45685,N_34534,N_38794);
nand U45686 (N_45686,N_37394,N_30991);
or U45687 (N_45687,N_30422,N_33408);
xor U45688 (N_45688,N_33592,N_34464);
or U45689 (N_45689,N_38421,N_34582);
xnor U45690 (N_45690,N_30566,N_33147);
or U45691 (N_45691,N_34066,N_34923);
xor U45692 (N_45692,N_34620,N_33452);
and U45693 (N_45693,N_32842,N_33830);
xnor U45694 (N_45694,N_39389,N_33051);
nand U45695 (N_45695,N_32506,N_36108);
nand U45696 (N_45696,N_38558,N_38590);
xor U45697 (N_45697,N_35826,N_34061);
and U45698 (N_45698,N_31745,N_30452);
nor U45699 (N_45699,N_38772,N_33774);
and U45700 (N_45700,N_38228,N_31198);
nand U45701 (N_45701,N_32612,N_34552);
nor U45702 (N_45702,N_31785,N_31843);
or U45703 (N_45703,N_39171,N_37543);
and U45704 (N_45704,N_34366,N_38846);
nor U45705 (N_45705,N_36735,N_35080);
nor U45706 (N_45706,N_34439,N_30341);
nand U45707 (N_45707,N_37270,N_38146);
nor U45708 (N_45708,N_39919,N_38318);
nor U45709 (N_45709,N_37705,N_32010);
nor U45710 (N_45710,N_31393,N_32246);
or U45711 (N_45711,N_31098,N_30046);
xnor U45712 (N_45712,N_35931,N_36352);
nand U45713 (N_45713,N_38623,N_32357);
and U45714 (N_45714,N_33989,N_36246);
and U45715 (N_45715,N_32875,N_34586);
or U45716 (N_45716,N_31099,N_36660);
and U45717 (N_45717,N_39219,N_37248);
nor U45718 (N_45718,N_37897,N_31197);
nor U45719 (N_45719,N_36553,N_37879);
or U45720 (N_45720,N_38695,N_33545);
or U45721 (N_45721,N_32273,N_32983);
xnor U45722 (N_45722,N_38331,N_38830);
nand U45723 (N_45723,N_37858,N_33051);
nor U45724 (N_45724,N_36738,N_34915);
nor U45725 (N_45725,N_30827,N_34187);
nor U45726 (N_45726,N_34019,N_31965);
xor U45727 (N_45727,N_33297,N_38295);
and U45728 (N_45728,N_34794,N_34822);
and U45729 (N_45729,N_34223,N_37409);
xor U45730 (N_45730,N_36051,N_30829);
nor U45731 (N_45731,N_30588,N_33377);
or U45732 (N_45732,N_31192,N_32328);
xor U45733 (N_45733,N_30496,N_35568);
and U45734 (N_45734,N_39140,N_39985);
xnor U45735 (N_45735,N_32563,N_30134);
nor U45736 (N_45736,N_33221,N_35582);
and U45737 (N_45737,N_35308,N_31075);
nor U45738 (N_45738,N_34228,N_33403);
nand U45739 (N_45739,N_34581,N_31384);
nor U45740 (N_45740,N_33897,N_38190);
or U45741 (N_45741,N_35407,N_32958);
xor U45742 (N_45742,N_36208,N_37104);
nor U45743 (N_45743,N_31041,N_33400);
and U45744 (N_45744,N_33471,N_34783);
xor U45745 (N_45745,N_39087,N_36541);
and U45746 (N_45746,N_36068,N_39509);
nand U45747 (N_45747,N_35971,N_31184);
nand U45748 (N_45748,N_39804,N_31860);
xor U45749 (N_45749,N_31528,N_36767);
xor U45750 (N_45750,N_39860,N_35280);
and U45751 (N_45751,N_39607,N_31035);
nor U45752 (N_45752,N_37225,N_38055);
and U45753 (N_45753,N_33678,N_31616);
nor U45754 (N_45754,N_36341,N_38333);
and U45755 (N_45755,N_35808,N_36697);
or U45756 (N_45756,N_37653,N_33097);
xnor U45757 (N_45757,N_33646,N_36221);
nor U45758 (N_45758,N_33449,N_30424);
nor U45759 (N_45759,N_38873,N_37482);
or U45760 (N_45760,N_37831,N_37316);
or U45761 (N_45761,N_38796,N_39945);
or U45762 (N_45762,N_37780,N_35574);
or U45763 (N_45763,N_34376,N_31807);
or U45764 (N_45764,N_39853,N_36283);
xnor U45765 (N_45765,N_33084,N_39183);
and U45766 (N_45766,N_33496,N_36616);
xnor U45767 (N_45767,N_30198,N_36674);
nor U45768 (N_45768,N_32952,N_33638);
xor U45769 (N_45769,N_39956,N_37298);
nor U45770 (N_45770,N_32231,N_35952);
nor U45771 (N_45771,N_34773,N_36846);
and U45772 (N_45772,N_33632,N_39510);
nand U45773 (N_45773,N_37997,N_31257);
or U45774 (N_45774,N_30338,N_32645);
or U45775 (N_45775,N_39384,N_39888);
and U45776 (N_45776,N_36392,N_35093);
and U45777 (N_45777,N_34553,N_32687);
xnor U45778 (N_45778,N_31229,N_36513);
nor U45779 (N_45779,N_34365,N_34374);
and U45780 (N_45780,N_36548,N_32632);
xnor U45781 (N_45781,N_32242,N_38257);
nand U45782 (N_45782,N_33240,N_34334);
and U45783 (N_45783,N_34526,N_33085);
nand U45784 (N_45784,N_32000,N_37304);
and U45785 (N_45785,N_33047,N_36498);
and U45786 (N_45786,N_38133,N_35841);
or U45787 (N_45787,N_37154,N_37696);
and U45788 (N_45788,N_37241,N_32617);
and U45789 (N_45789,N_37213,N_35902);
nor U45790 (N_45790,N_30761,N_37606);
or U45791 (N_45791,N_38038,N_37251);
xnor U45792 (N_45792,N_36478,N_33043);
nand U45793 (N_45793,N_37401,N_34443);
nor U45794 (N_45794,N_37232,N_38074);
or U45795 (N_45795,N_33192,N_32365);
xor U45796 (N_45796,N_30470,N_39943);
nand U45797 (N_45797,N_30300,N_36236);
nand U45798 (N_45798,N_34043,N_33663);
xor U45799 (N_45799,N_38914,N_30970);
nand U45800 (N_45800,N_39587,N_35848);
nor U45801 (N_45801,N_31662,N_31649);
nand U45802 (N_45802,N_33032,N_34846);
or U45803 (N_45803,N_38080,N_38659);
nor U45804 (N_45804,N_39807,N_35249);
and U45805 (N_45805,N_39832,N_39650);
nand U45806 (N_45806,N_30956,N_36143);
or U45807 (N_45807,N_35837,N_30499);
nand U45808 (N_45808,N_36603,N_31213);
and U45809 (N_45809,N_35028,N_34130);
or U45810 (N_45810,N_33194,N_31212);
nand U45811 (N_45811,N_39663,N_37867);
xor U45812 (N_45812,N_32294,N_31513);
nand U45813 (N_45813,N_37783,N_37713);
and U45814 (N_45814,N_38925,N_34887);
and U45815 (N_45815,N_34342,N_34121);
xnor U45816 (N_45816,N_38355,N_37231);
nand U45817 (N_45817,N_36620,N_34417);
nor U45818 (N_45818,N_33467,N_34834);
xnor U45819 (N_45819,N_30398,N_30738);
xor U45820 (N_45820,N_37543,N_35391);
or U45821 (N_45821,N_35362,N_34597);
or U45822 (N_45822,N_32407,N_37550);
and U45823 (N_45823,N_38411,N_31275);
and U45824 (N_45824,N_30518,N_34146);
nor U45825 (N_45825,N_30758,N_33945);
xor U45826 (N_45826,N_37617,N_33195);
and U45827 (N_45827,N_36315,N_31099);
nand U45828 (N_45828,N_39324,N_35723);
or U45829 (N_45829,N_32653,N_31408);
or U45830 (N_45830,N_38065,N_38222);
nand U45831 (N_45831,N_32491,N_33373);
nand U45832 (N_45832,N_32416,N_37516);
or U45833 (N_45833,N_36785,N_36554);
xor U45834 (N_45834,N_31132,N_38492);
nand U45835 (N_45835,N_34275,N_31183);
xnor U45836 (N_45836,N_34704,N_38855);
and U45837 (N_45837,N_36186,N_33409);
and U45838 (N_45838,N_35285,N_39336);
and U45839 (N_45839,N_34423,N_31324);
and U45840 (N_45840,N_33267,N_31342);
or U45841 (N_45841,N_32356,N_39278);
and U45842 (N_45842,N_37906,N_31481);
xor U45843 (N_45843,N_37513,N_31177);
xor U45844 (N_45844,N_35792,N_34119);
or U45845 (N_45845,N_30782,N_38925);
nor U45846 (N_45846,N_33173,N_30177);
nor U45847 (N_45847,N_31569,N_32886);
xnor U45848 (N_45848,N_32848,N_31623);
nor U45849 (N_45849,N_30736,N_36260);
xor U45850 (N_45850,N_39325,N_38574);
xor U45851 (N_45851,N_35182,N_34576);
nand U45852 (N_45852,N_32501,N_37659);
nand U45853 (N_45853,N_32829,N_31009);
nor U45854 (N_45854,N_34222,N_30870);
xnor U45855 (N_45855,N_33223,N_30665);
or U45856 (N_45856,N_35752,N_32761);
or U45857 (N_45857,N_33570,N_32181);
nor U45858 (N_45858,N_33141,N_37635);
nand U45859 (N_45859,N_39370,N_33960);
nand U45860 (N_45860,N_32911,N_39664);
and U45861 (N_45861,N_39861,N_31499);
xnor U45862 (N_45862,N_34916,N_38763);
or U45863 (N_45863,N_32206,N_37189);
nand U45864 (N_45864,N_30045,N_33361);
or U45865 (N_45865,N_32981,N_37893);
or U45866 (N_45866,N_38384,N_32170);
or U45867 (N_45867,N_30123,N_37279);
nor U45868 (N_45868,N_39426,N_38588);
and U45869 (N_45869,N_39298,N_39682);
nor U45870 (N_45870,N_38399,N_32348);
xor U45871 (N_45871,N_33203,N_30912);
nor U45872 (N_45872,N_30689,N_33015);
nand U45873 (N_45873,N_31945,N_38925);
and U45874 (N_45874,N_30249,N_34566);
and U45875 (N_45875,N_39290,N_30488);
xnor U45876 (N_45876,N_32502,N_36251);
nor U45877 (N_45877,N_34820,N_30492);
and U45878 (N_45878,N_31504,N_33244);
xor U45879 (N_45879,N_39149,N_36280);
and U45880 (N_45880,N_35207,N_35139);
nand U45881 (N_45881,N_30153,N_31472);
xor U45882 (N_45882,N_32696,N_32768);
xnor U45883 (N_45883,N_36299,N_31055);
nor U45884 (N_45884,N_35213,N_32251);
nor U45885 (N_45885,N_39059,N_33275);
nor U45886 (N_45886,N_36706,N_31766);
and U45887 (N_45887,N_30344,N_32204);
or U45888 (N_45888,N_34987,N_31261);
nor U45889 (N_45889,N_39383,N_35443);
or U45890 (N_45890,N_37896,N_32658);
nor U45891 (N_45891,N_35206,N_37685);
nor U45892 (N_45892,N_39473,N_32764);
and U45893 (N_45893,N_37531,N_35162);
or U45894 (N_45894,N_34387,N_31532);
xnor U45895 (N_45895,N_38902,N_34106);
and U45896 (N_45896,N_31500,N_39501);
xor U45897 (N_45897,N_33495,N_31325);
and U45898 (N_45898,N_38844,N_39141);
nor U45899 (N_45899,N_30233,N_37098);
xnor U45900 (N_45900,N_33591,N_30060);
and U45901 (N_45901,N_30536,N_35941);
xor U45902 (N_45902,N_34244,N_35733);
or U45903 (N_45903,N_30156,N_35668);
nor U45904 (N_45904,N_37992,N_32235);
xor U45905 (N_45905,N_31944,N_34796);
and U45906 (N_45906,N_32911,N_31350);
nor U45907 (N_45907,N_33885,N_38985);
nor U45908 (N_45908,N_30921,N_30935);
or U45909 (N_45909,N_34565,N_36719);
or U45910 (N_45910,N_32308,N_34374);
nor U45911 (N_45911,N_30282,N_36941);
nor U45912 (N_45912,N_34984,N_33980);
nand U45913 (N_45913,N_37842,N_39452);
nor U45914 (N_45914,N_39067,N_32325);
and U45915 (N_45915,N_37227,N_31470);
or U45916 (N_45916,N_35762,N_33183);
nand U45917 (N_45917,N_30869,N_36970);
nor U45918 (N_45918,N_38448,N_36770);
and U45919 (N_45919,N_37584,N_35329);
nor U45920 (N_45920,N_31591,N_37213);
or U45921 (N_45921,N_30502,N_39000);
xor U45922 (N_45922,N_33584,N_35400);
xor U45923 (N_45923,N_30006,N_35674);
and U45924 (N_45924,N_35339,N_33576);
and U45925 (N_45925,N_31662,N_30126);
xnor U45926 (N_45926,N_30451,N_36011);
nor U45927 (N_45927,N_38441,N_34378);
xnor U45928 (N_45928,N_37072,N_37903);
nor U45929 (N_45929,N_32601,N_30915);
nor U45930 (N_45930,N_32114,N_32152);
and U45931 (N_45931,N_32638,N_36384);
and U45932 (N_45932,N_39955,N_31311);
nand U45933 (N_45933,N_36609,N_31251);
xnor U45934 (N_45934,N_30153,N_33970);
and U45935 (N_45935,N_30937,N_32982);
and U45936 (N_45936,N_32418,N_32652);
and U45937 (N_45937,N_31432,N_35959);
xor U45938 (N_45938,N_34432,N_33291);
nand U45939 (N_45939,N_31799,N_36285);
nand U45940 (N_45940,N_36272,N_35334);
xor U45941 (N_45941,N_39124,N_32343);
xor U45942 (N_45942,N_32759,N_37111);
or U45943 (N_45943,N_32165,N_33175);
nand U45944 (N_45944,N_34853,N_35774);
and U45945 (N_45945,N_38667,N_36818);
nand U45946 (N_45946,N_39844,N_35168);
nand U45947 (N_45947,N_37792,N_31199);
and U45948 (N_45948,N_36730,N_34412);
nor U45949 (N_45949,N_38601,N_31467);
nor U45950 (N_45950,N_30645,N_36856);
nand U45951 (N_45951,N_35792,N_31952);
xor U45952 (N_45952,N_37141,N_36565);
and U45953 (N_45953,N_34546,N_34797);
and U45954 (N_45954,N_35638,N_38646);
nor U45955 (N_45955,N_31891,N_39557);
or U45956 (N_45956,N_35706,N_34859);
nor U45957 (N_45957,N_31448,N_38487);
nand U45958 (N_45958,N_34368,N_30012);
nor U45959 (N_45959,N_36560,N_33419);
and U45960 (N_45960,N_33978,N_32856);
nand U45961 (N_45961,N_31566,N_36453);
xnor U45962 (N_45962,N_35048,N_36167);
nand U45963 (N_45963,N_36064,N_33591);
or U45964 (N_45964,N_36032,N_37939);
xor U45965 (N_45965,N_34353,N_39584);
xnor U45966 (N_45966,N_39005,N_37762);
or U45967 (N_45967,N_38644,N_39981);
nor U45968 (N_45968,N_38137,N_35462);
xor U45969 (N_45969,N_39307,N_34500);
and U45970 (N_45970,N_35790,N_39582);
xnor U45971 (N_45971,N_37526,N_34594);
or U45972 (N_45972,N_31582,N_32335);
nor U45973 (N_45973,N_34656,N_32036);
nand U45974 (N_45974,N_32845,N_34493);
xnor U45975 (N_45975,N_36610,N_30927);
nand U45976 (N_45976,N_30919,N_34274);
or U45977 (N_45977,N_39271,N_37785);
nor U45978 (N_45978,N_33273,N_34272);
nor U45979 (N_45979,N_31400,N_31959);
nor U45980 (N_45980,N_34995,N_33218);
nand U45981 (N_45981,N_35223,N_37210);
nand U45982 (N_45982,N_31065,N_30881);
or U45983 (N_45983,N_32422,N_36835);
xnor U45984 (N_45984,N_39280,N_30626);
or U45985 (N_45985,N_35914,N_33343);
nor U45986 (N_45986,N_33047,N_38550);
nand U45987 (N_45987,N_35109,N_38954);
nor U45988 (N_45988,N_37201,N_30208);
or U45989 (N_45989,N_31739,N_36309);
nand U45990 (N_45990,N_39325,N_30123);
xnor U45991 (N_45991,N_36675,N_33282);
xor U45992 (N_45992,N_36821,N_31583);
or U45993 (N_45993,N_33762,N_33764);
and U45994 (N_45994,N_30096,N_34928);
nor U45995 (N_45995,N_33202,N_39967);
nor U45996 (N_45996,N_33573,N_30057);
or U45997 (N_45997,N_36960,N_30080);
and U45998 (N_45998,N_34230,N_33351);
nand U45999 (N_45999,N_38658,N_39101);
xnor U46000 (N_46000,N_39190,N_35830);
nand U46001 (N_46001,N_35270,N_38305);
nor U46002 (N_46002,N_33337,N_34177);
or U46003 (N_46003,N_33506,N_36919);
or U46004 (N_46004,N_39331,N_34725);
nand U46005 (N_46005,N_33543,N_38945);
nor U46006 (N_46006,N_35156,N_36417);
xor U46007 (N_46007,N_33369,N_37810);
or U46008 (N_46008,N_36430,N_39882);
nor U46009 (N_46009,N_38795,N_38614);
or U46010 (N_46010,N_38313,N_34997);
nor U46011 (N_46011,N_34830,N_30589);
nand U46012 (N_46012,N_34240,N_38701);
or U46013 (N_46013,N_37893,N_35806);
and U46014 (N_46014,N_30121,N_35367);
nor U46015 (N_46015,N_31303,N_30254);
or U46016 (N_46016,N_37379,N_39496);
xnor U46017 (N_46017,N_32233,N_32487);
or U46018 (N_46018,N_30139,N_36217);
or U46019 (N_46019,N_35396,N_34429);
xor U46020 (N_46020,N_37369,N_35922);
nor U46021 (N_46021,N_34795,N_34562);
and U46022 (N_46022,N_34363,N_38049);
xnor U46023 (N_46023,N_38003,N_38883);
and U46024 (N_46024,N_32813,N_37099);
nor U46025 (N_46025,N_37690,N_30912);
or U46026 (N_46026,N_30260,N_32955);
nor U46027 (N_46027,N_34575,N_36982);
nor U46028 (N_46028,N_30137,N_34856);
and U46029 (N_46029,N_36027,N_35142);
or U46030 (N_46030,N_32908,N_33953);
xnor U46031 (N_46031,N_36311,N_35102);
and U46032 (N_46032,N_34522,N_36350);
or U46033 (N_46033,N_33389,N_37401);
xor U46034 (N_46034,N_32928,N_38041);
nor U46035 (N_46035,N_39779,N_33670);
or U46036 (N_46036,N_33246,N_36432);
and U46037 (N_46037,N_39239,N_36187);
nand U46038 (N_46038,N_34700,N_31054);
nor U46039 (N_46039,N_38152,N_32279);
and U46040 (N_46040,N_39551,N_30795);
nor U46041 (N_46041,N_34009,N_33225);
or U46042 (N_46042,N_31262,N_31277);
or U46043 (N_46043,N_39583,N_33625);
or U46044 (N_46044,N_31864,N_39493);
or U46045 (N_46045,N_32868,N_34627);
and U46046 (N_46046,N_34144,N_37314);
xor U46047 (N_46047,N_37439,N_33980);
nand U46048 (N_46048,N_38607,N_34529);
nand U46049 (N_46049,N_30847,N_32569);
and U46050 (N_46050,N_39240,N_31497);
or U46051 (N_46051,N_36334,N_38203);
nand U46052 (N_46052,N_37784,N_37129);
xor U46053 (N_46053,N_31466,N_31724);
xnor U46054 (N_46054,N_34889,N_31571);
nor U46055 (N_46055,N_30757,N_38844);
or U46056 (N_46056,N_36231,N_30506);
or U46057 (N_46057,N_34383,N_33593);
and U46058 (N_46058,N_31019,N_31941);
nor U46059 (N_46059,N_39933,N_35127);
xnor U46060 (N_46060,N_35932,N_38480);
and U46061 (N_46061,N_38865,N_34409);
nor U46062 (N_46062,N_34667,N_31070);
and U46063 (N_46063,N_33500,N_36569);
xor U46064 (N_46064,N_36139,N_35680);
nand U46065 (N_46065,N_34562,N_38075);
xnor U46066 (N_46066,N_39875,N_33002);
nand U46067 (N_46067,N_36813,N_35247);
nor U46068 (N_46068,N_37860,N_34300);
nand U46069 (N_46069,N_35089,N_36055);
nand U46070 (N_46070,N_37261,N_34054);
nand U46071 (N_46071,N_30946,N_37357);
or U46072 (N_46072,N_33213,N_35811);
nand U46073 (N_46073,N_39618,N_31326);
nor U46074 (N_46074,N_36793,N_35824);
or U46075 (N_46075,N_38848,N_33900);
nand U46076 (N_46076,N_32259,N_35602);
nor U46077 (N_46077,N_34569,N_31273);
nor U46078 (N_46078,N_32809,N_31824);
or U46079 (N_46079,N_37603,N_35894);
nand U46080 (N_46080,N_36212,N_32038);
or U46081 (N_46081,N_37051,N_39769);
nor U46082 (N_46082,N_35447,N_38108);
nor U46083 (N_46083,N_34963,N_31563);
or U46084 (N_46084,N_33498,N_34037);
and U46085 (N_46085,N_36410,N_30652);
xor U46086 (N_46086,N_35302,N_32910);
and U46087 (N_46087,N_33328,N_33537);
xnor U46088 (N_46088,N_32839,N_35395);
or U46089 (N_46089,N_32658,N_31558);
or U46090 (N_46090,N_36566,N_31517);
or U46091 (N_46091,N_35049,N_30543);
nand U46092 (N_46092,N_32363,N_35256);
nand U46093 (N_46093,N_36565,N_37774);
nor U46094 (N_46094,N_39467,N_30035);
or U46095 (N_46095,N_33567,N_39797);
and U46096 (N_46096,N_34007,N_37306);
nor U46097 (N_46097,N_39114,N_36567);
and U46098 (N_46098,N_38534,N_38713);
nand U46099 (N_46099,N_35306,N_33756);
or U46100 (N_46100,N_31007,N_37952);
xnor U46101 (N_46101,N_35982,N_31475);
nor U46102 (N_46102,N_36503,N_36415);
xnor U46103 (N_46103,N_38313,N_33964);
nand U46104 (N_46104,N_37977,N_35466);
and U46105 (N_46105,N_39371,N_38568);
or U46106 (N_46106,N_33168,N_33896);
xor U46107 (N_46107,N_36565,N_34432);
nand U46108 (N_46108,N_39133,N_36138);
and U46109 (N_46109,N_31621,N_33299);
and U46110 (N_46110,N_31493,N_37547);
nor U46111 (N_46111,N_37229,N_31505);
xor U46112 (N_46112,N_35919,N_38331);
nor U46113 (N_46113,N_31312,N_31927);
nand U46114 (N_46114,N_37606,N_30463);
and U46115 (N_46115,N_31207,N_39127);
nor U46116 (N_46116,N_34980,N_30984);
and U46117 (N_46117,N_31208,N_38071);
nor U46118 (N_46118,N_37425,N_32114);
nand U46119 (N_46119,N_39351,N_36706);
nand U46120 (N_46120,N_30404,N_33064);
or U46121 (N_46121,N_33445,N_34347);
nand U46122 (N_46122,N_35802,N_32326);
nand U46123 (N_46123,N_36667,N_38380);
nand U46124 (N_46124,N_31442,N_30271);
and U46125 (N_46125,N_33775,N_30869);
nor U46126 (N_46126,N_38853,N_31991);
or U46127 (N_46127,N_34879,N_39598);
or U46128 (N_46128,N_35345,N_39288);
and U46129 (N_46129,N_36955,N_32591);
nand U46130 (N_46130,N_39740,N_37375);
and U46131 (N_46131,N_37709,N_30861);
xor U46132 (N_46132,N_30775,N_30214);
nor U46133 (N_46133,N_31172,N_38398);
or U46134 (N_46134,N_31292,N_34767);
or U46135 (N_46135,N_39392,N_33611);
or U46136 (N_46136,N_35123,N_30175);
nor U46137 (N_46137,N_32641,N_39063);
and U46138 (N_46138,N_37843,N_30647);
nor U46139 (N_46139,N_38235,N_30188);
and U46140 (N_46140,N_37587,N_38877);
nand U46141 (N_46141,N_34225,N_34091);
or U46142 (N_46142,N_39015,N_33754);
or U46143 (N_46143,N_33365,N_36521);
nor U46144 (N_46144,N_35474,N_39673);
and U46145 (N_46145,N_32667,N_30458);
or U46146 (N_46146,N_33206,N_30634);
and U46147 (N_46147,N_35506,N_30706);
or U46148 (N_46148,N_33487,N_30664);
xor U46149 (N_46149,N_34562,N_30023);
nor U46150 (N_46150,N_32271,N_30861);
and U46151 (N_46151,N_35950,N_30191);
nor U46152 (N_46152,N_35438,N_39183);
and U46153 (N_46153,N_35537,N_35890);
nand U46154 (N_46154,N_30157,N_37783);
and U46155 (N_46155,N_31148,N_35836);
nand U46156 (N_46156,N_36600,N_30607);
nand U46157 (N_46157,N_33386,N_36614);
nand U46158 (N_46158,N_32721,N_32672);
or U46159 (N_46159,N_32684,N_36440);
or U46160 (N_46160,N_39712,N_33720);
nand U46161 (N_46161,N_34393,N_31042);
xor U46162 (N_46162,N_31861,N_37454);
or U46163 (N_46163,N_30983,N_35970);
nand U46164 (N_46164,N_37659,N_37530);
xor U46165 (N_46165,N_39325,N_32438);
nand U46166 (N_46166,N_39978,N_30202);
nand U46167 (N_46167,N_36350,N_36672);
nor U46168 (N_46168,N_39405,N_34885);
nor U46169 (N_46169,N_33963,N_30751);
and U46170 (N_46170,N_31126,N_37903);
and U46171 (N_46171,N_31964,N_39822);
and U46172 (N_46172,N_36740,N_38572);
xor U46173 (N_46173,N_34509,N_37653);
or U46174 (N_46174,N_39646,N_35979);
and U46175 (N_46175,N_36361,N_35115);
or U46176 (N_46176,N_35459,N_33935);
nor U46177 (N_46177,N_32147,N_36971);
and U46178 (N_46178,N_34196,N_33056);
nor U46179 (N_46179,N_30848,N_30258);
nand U46180 (N_46180,N_38326,N_33790);
and U46181 (N_46181,N_39626,N_34152);
or U46182 (N_46182,N_31031,N_30526);
or U46183 (N_46183,N_35377,N_31986);
and U46184 (N_46184,N_36121,N_31118);
xor U46185 (N_46185,N_34160,N_32617);
or U46186 (N_46186,N_34933,N_30303);
and U46187 (N_46187,N_34514,N_36059);
and U46188 (N_46188,N_30330,N_31818);
or U46189 (N_46189,N_39805,N_38510);
xor U46190 (N_46190,N_31011,N_30448);
nand U46191 (N_46191,N_32600,N_38344);
and U46192 (N_46192,N_30389,N_33970);
nand U46193 (N_46193,N_39970,N_33274);
nand U46194 (N_46194,N_32835,N_31705);
xnor U46195 (N_46195,N_39866,N_39858);
or U46196 (N_46196,N_35037,N_39786);
nand U46197 (N_46197,N_37576,N_30894);
or U46198 (N_46198,N_37677,N_37209);
and U46199 (N_46199,N_35107,N_38514);
or U46200 (N_46200,N_30976,N_38331);
nand U46201 (N_46201,N_36031,N_31150);
nor U46202 (N_46202,N_31655,N_39251);
xor U46203 (N_46203,N_34963,N_35938);
nor U46204 (N_46204,N_37290,N_30114);
xnor U46205 (N_46205,N_35586,N_33380);
nand U46206 (N_46206,N_38008,N_30819);
and U46207 (N_46207,N_35591,N_38204);
or U46208 (N_46208,N_31696,N_31863);
and U46209 (N_46209,N_38147,N_36338);
and U46210 (N_46210,N_34710,N_31874);
nand U46211 (N_46211,N_38250,N_36210);
nand U46212 (N_46212,N_31085,N_30944);
or U46213 (N_46213,N_34426,N_36875);
xor U46214 (N_46214,N_32739,N_35134);
or U46215 (N_46215,N_39828,N_35199);
or U46216 (N_46216,N_37121,N_39740);
xnor U46217 (N_46217,N_35681,N_37793);
or U46218 (N_46218,N_39665,N_38931);
or U46219 (N_46219,N_30425,N_36536);
nor U46220 (N_46220,N_30455,N_37502);
xor U46221 (N_46221,N_32880,N_37006);
and U46222 (N_46222,N_31358,N_37936);
or U46223 (N_46223,N_34998,N_37731);
xnor U46224 (N_46224,N_31486,N_35694);
and U46225 (N_46225,N_39549,N_37950);
nor U46226 (N_46226,N_31832,N_38636);
and U46227 (N_46227,N_34604,N_35823);
and U46228 (N_46228,N_33724,N_36468);
nor U46229 (N_46229,N_30112,N_39601);
xnor U46230 (N_46230,N_38644,N_34042);
xnor U46231 (N_46231,N_31347,N_30707);
xor U46232 (N_46232,N_30931,N_31689);
nand U46233 (N_46233,N_36422,N_33293);
nor U46234 (N_46234,N_31853,N_36494);
xor U46235 (N_46235,N_32040,N_35979);
and U46236 (N_46236,N_33516,N_31106);
and U46237 (N_46237,N_36950,N_34091);
nand U46238 (N_46238,N_31079,N_39111);
nor U46239 (N_46239,N_38953,N_30592);
nand U46240 (N_46240,N_32538,N_36211);
nor U46241 (N_46241,N_35741,N_34579);
or U46242 (N_46242,N_32284,N_31237);
nor U46243 (N_46243,N_32510,N_37087);
and U46244 (N_46244,N_36590,N_31830);
and U46245 (N_46245,N_32311,N_34447);
nor U46246 (N_46246,N_32506,N_38110);
or U46247 (N_46247,N_30729,N_33170);
or U46248 (N_46248,N_35096,N_38479);
nor U46249 (N_46249,N_38276,N_35992);
or U46250 (N_46250,N_37811,N_35822);
or U46251 (N_46251,N_30080,N_39730);
nand U46252 (N_46252,N_33318,N_36650);
or U46253 (N_46253,N_35811,N_35406);
nand U46254 (N_46254,N_31783,N_38786);
nor U46255 (N_46255,N_33195,N_36041);
or U46256 (N_46256,N_33228,N_36884);
nand U46257 (N_46257,N_32159,N_30428);
nor U46258 (N_46258,N_39547,N_38765);
or U46259 (N_46259,N_34740,N_31304);
nand U46260 (N_46260,N_30163,N_32130);
or U46261 (N_46261,N_30419,N_33590);
nor U46262 (N_46262,N_39873,N_32731);
nor U46263 (N_46263,N_38650,N_37240);
or U46264 (N_46264,N_36371,N_30149);
or U46265 (N_46265,N_39648,N_30186);
nor U46266 (N_46266,N_32509,N_35231);
nand U46267 (N_46267,N_32339,N_39217);
nor U46268 (N_46268,N_31946,N_35817);
nand U46269 (N_46269,N_34614,N_32994);
nor U46270 (N_46270,N_38328,N_39774);
and U46271 (N_46271,N_36864,N_37315);
or U46272 (N_46272,N_34310,N_35325);
nor U46273 (N_46273,N_30209,N_35687);
nand U46274 (N_46274,N_37565,N_32757);
or U46275 (N_46275,N_34117,N_34693);
and U46276 (N_46276,N_36039,N_34241);
and U46277 (N_46277,N_31236,N_35747);
or U46278 (N_46278,N_33514,N_36924);
nand U46279 (N_46279,N_31751,N_37174);
xor U46280 (N_46280,N_31446,N_35763);
nand U46281 (N_46281,N_37554,N_38781);
nand U46282 (N_46282,N_37742,N_37881);
xnor U46283 (N_46283,N_33780,N_38037);
or U46284 (N_46284,N_33576,N_30382);
and U46285 (N_46285,N_33870,N_31645);
nand U46286 (N_46286,N_30352,N_37159);
and U46287 (N_46287,N_32914,N_30456);
xnor U46288 (N_46288,N_35687,N_35211);
and U46289 (N_46289,N_39816,N_34470);
or U46290 (N_46290,N_34751,N_38539);
and U46291 (N_46291,N_31795,N_31048);
or U46292 (N_46292,N_38562,N_34675);
nor U46293 (N_46293,N_38316,N_35093);
nand U46294 (N_46294,N_31171,N_33940);
nor U46295 (N_46295,N_35253,N_35099);
and U46296 (N_46296,N_34217,N_37558);
and U46297 (N_46297,N_37189,N_35417);
and U46298 (N_46298,N_34632,N_36342);
nand U46299 (N_46299,N_33457,N_32397);
or U46300 (N_46300,N_34546,N_31973);
or U46301 (N_46301,N_32264,N_35927);
nor U46302 (N_46302,N_31667,N_32131);
or U46303 (N_46303,N_39858,N_34450);
and U46304 (N_46304,N_38938,N_36302);
nand U46305 (N_46305,N_32023,N_34871);
nor U46306 (N_46306,N_32931,N_38759);
or U46307 (N_46307,N_35713,N_33494);
or U46308 (N_46308,N_36908,N_34061);
or U46309 (N_46309,N_35986,N_32937);
or U46310 (N_46310,N_32813,N_32762);
and U46311 (N_46311,N_36999,N_34933);
nor U46312 (N_46312,N_39204,N_36103);
and U46313 (N_46313,N_39925,N_30194);
nand U46314 (N_46314,N_35096,N_35451);
xor U46315 (N_46315,N_37502,N_39148);
nand U46316 (N_46316,N_36493,N_37299);
xor U46317 (N_46317,N_30229,N_36950);
xnor U46318 (N_46318,N_30111,N_37241);
and U46319 (N_46319,N_32981,N_39428);
and U46320 (N_46320,N_32934,N_30486);
nor U46321 (N_46321,N_32357,N_37374);
nand U46322 (N_46322,N_38535,N_32178);
xnor U46323 (N_46323,N_35807,N_32198);
nor U46324 (N_46324,N_33669,N_31749);
nor U46325 (N_46325,N_39634,N_32752);
nand U46326 (N_46326,N_39631,N_33959);
xnor U46327 (N_46327,N_36979,N_31857);
and U46328 (N_46328,N_33927,N_32636);
and U46329 (N_46329,N_33441,N_35433);
nand U46330 (N_46330,N_39256,N_30546);
nand U46331 (N_46331,N_32025,N_37854);
xor U46332 (N_46332,N_30078,N_38297);
xor U46333 (N_46333,N_37864,N_35956);
and U46334 (N_46334,N_36921,N_36281);
nor U46335 (N_46335,N_37092,N_38485);
nor U46336 (N_46336,N_37106,N_34754);
nor U46337 (N_46337,N_34439,N_31643);
xnor U46338 (N_46338,N_36135,N_36555);
nand U46339 (N_46339,N_34876,N_38261);
xor U46340 (N_46340,N_34352,N_37588);
and U46341 (N_46341,N_30562,N_38345);
nand U46342 (N_46342,N_38523,N_32374);
and U46343 (N_46343,N_30303,N_38307);
nor U46344 (N_46344,N_37033,N_35892);
or U46345 (N_46345,N_37454,N_33206);
nor U46346 (N_46346,N_38933,N_34433);
nand U46347 (N_46347,N_36575,N_32670);
nor U46348 (N_46348,N_37964,N_38883);
xnor U46349 (N_46349,N_39358,N_30434);
nand U46350 (N_46350,N_35265,N_39020);
or U46351 (N_46351,N_33623,N_39507);
or U46352 (N_46352,N_37191,N_34374);
or U46353 (N_46353,N_36143,N_32057);
nor U46354 (N_46354,N_30177,N_31992);
or U46355 (N_46355,N_37272,N_34888);
nand U46356 (N_46356,N_31344,N_33388);
xnor U46357 (N_46357,N_37764,N_36264);
nand U46358 (N_46358,N_32083,N_35918);
and U46359 (N_46359,N_36088,N_33725);
xor U46360 (N_46360,N_33030,N_37260);
xnor U46361 (N_46361,N_38010,N_33325);
or U46362 (N_46362,N_35087,N_38168);
or U46363 (N_46363,N_38143,N_34962);
nor U46364 (N_46364,N_38000,N_39476);
nor U46365 (N_46365,N_31017,N_36097);
or U46366 (N_46366,N_34638,N_33578);
nand U46367 (N_46367,N_36520,N_37446);
and U46368 (N_46368,N_37135,N_39060);
nand U46369 (N_46369,N_35639,N_38007);
nand U46370 (N_46370,N_39383,N_32552);
nor U46371 (N_46371,N_34315,N_38346);
or U46372 (N_46372,N_34709,N_39795);
xor U46373 (N_46373,N_34308,N_36647);
nor U46374 (N_46374,N_39414,N_32760);
nand U46375 (N_46375,N_38572,N_31518);
nor U46376 (N_46376,N_38857,N_39869);
or U46377 (N_46377,N_38210,N_37501);
nand U46378 (N_46378,N_30323,N_37501);
xor U46379 (N_46379,N_39464,N_32002);
and U46380 (N_46380,N_37767,N_31502);
or U46381 (N_46381,N_34414,N_35744);
xor U46382 (N_46382,N_35932,N_34089);
xnor U46383 (N_46383,N_38701,N_33236);
xor U46384 (N_46384,N_31179,N_39816);
or U46385 (N_46385,N_35660,N_30100);
nand U46386 (N_46386,N_34344,N_30812);
nor U46387 (N_46387,N_37265,N_39742);
nor U46388 (N_46388,N_35053,N_35584);
or U46389 (N_46389,N_37215,N_37076);
xor U46390 (N_46390,N_39662,N_37812);
and U46391 (N_46391,N_38208,N_32794);
nand U46392 (N_46392,N_34991,N_38067);
nand U46393 (N_46393,N_31050,N_33026);
and U46394 (N_46394,N_38380,N_32832);
and U46395 (N_46395,N_34092,N_34205);
or U46396 (N_46396,N_36033,N_34676);
and U46397 (N_46397,N_32146,N_32907);
xnor U46398 (N_46398,N_31287,N_39181);
nor U46399 (N_46399,N_31992,N_36665);
nand U46400 (N_46400,N_33680,N_36455);
nand U46401 (N_46401,N_35070,N_35196);
nor U46402 (N_46402,N_38973,N_30911);
nor U46403 (N_46403,N_32800,N_34415);
xor U46404 (N_46404,N_38050,N_37527);
xor U46405 (N_46405,N_38975,N_37132);
nor U46406 (N_46406,N_36764,N_32285);
nand U46407 (N_46407,N_34511,N_38197);
nor U46408 (N_46408,N_38719,N_38005);
and U46409 (N_46409,N_30141,N_34881);
or U46410 (N_46410,N_35105,N_37621);
xnor U46411 (N_46411,N_34912,N_39966);
and U46412 (N_46412,N_36508,N_32926);
and U46413 (N_46413,N_34477,N_32727);
xnor U46414 (N_46414,N_37136,N_30899);
nor U46415 (N_46415,N_33956,N_31753);
xnor U46416 (N_46416,N_34262,N_33456);
or U46417 (N_46417,N_34179,N_37414);
nor U46418 (N_46418,N_34109,N_37018);
or U46419 (N_46419,N_30997,N_34719);
and U46420 (N_46420,N_32417,N_31240);
and U46421 (N_46421,N_31741,N_39691);
and U46422 (N_46422,N_31119,N_30859);
and U46423 (N_46423,N_36153,N_32379);
and U46424 (N_46424,N_31340,N_33380);
nand U46425 (N_46425,N_34020,N_34535);
nand U46426 (N_46426,N_33346,N_39159);
nor U46427 (N_46427,N_31571,N_33883);
and U46428 (N_46428,N_39651,N_30276);
nor U46429 (N_46429,N_30656,N_35705);
or U46430 (N_46430,N_31488,N_33934);
nand U46431 (N_46431,N_31396,N_34346);
xnor U46432 (N_46432,N_38230,N_33723);
nor U46433 (N_46433,N_38029,N_33218);
or U46434 (N_46434,N_36783,N_35666);
or U46435 (N_46435,N_30911,N_35835);
or U46436 (N_46436,N_37850,N_32300);
xor U46437 (N_46437,N_31826,N_34903);
xor U46438 (N_46438,N_31669,N_31240);
nor U46439 (N_46439,N_37854,N_37585);
nand U46440 (N_46440,N_32784,N_36080);
nor U46441 (N_46441,N_35008,N_31512);
nor U46442 (N_46442,N_36451,N_31530);
nor U46443 (N_46443,N_34071,N_37589);
or U46444 (N_46444,N_32231,N_34323);
nand U46445 (N_46445,N_32205,N_31932);
xnor U46446 (N_46446,N_35721,N_31168);
or U46447 (N_46447,N_36111,N_36346);
and U46448 (N_46448,N_35390,N_30053);
xnor U46449 (N_46449,N_30819,N_30375);
or U46450 (N_46450,N_33916,N_34488);
nand U46451 (N_46451,N_34250,N_30299);
or U46452 (N_46452,N_39057,N_36738);
nand U46453 (N_46453,N_36348,N_39290);
nand U46454 (N_46454,N_39961,N_38377);
nand U46455 (N_46455,N_39834,N_34700);
nand U46456 (N_46456,N_31043,N_34887);
xor U46457 (N_46457,N_34659,N_39034);
and U46458 (N_46458,N_37079,N_34019);
and U46459 (N_46459,N_36700,N_37068);
xnor U46460 (N_46460,N_32548,N_32542);
or U46461 (N_46461,N_35854,N_36747);
and U46462 (N_46462,N_37702,N_32086);
or U46463 (N_46463,N_36834,N_38370);
nor U46464 (N_46464,N_30155,N_36533);
or U46465 (N_46465,N_35137,N_36009);
xor U46466 (N_46466,N_38459,N_37180);
nand U46467 (N_46467,N_38366,N_34535);
nand U46468 (N_46468,N_38906,N_33918);
and U46469 (N_46469,N_30399,N_37092);
nand U46470 (N_46470,N_30300,N_36989);
nor U46471 (N_46471,N_38986,N_36249);
or U46472 (N_46472,N_37179,N_30917);
or U46473 (N_46473,N_31801,N_36041);
nand U46474 (N_46474,N_38071,N_32293);
or U46475 (N_46475,N_38361,N_35312);
and U46476 (N_46476,N_31153,N_32125);
or U46477 (N_46477,N_35289,N_34494);
or U46478 (N_46478,N_33613,N_35015);
or U46479 (N_46479,N_36655,N_31238);
or U46480 (N_46480,N_30310,N_33211);
and U46481 (N_46481,N_38343,N_37506);
xnor U46482 (N_46482,N_30188,N_37075);
xnor U46483 (N_46483,N_35097,N_37333);
and U46484 (N_46484,N_34884,N_35804);
nand U46485 (N_46485,N_30331,N_30591);
and U46486 (N_46486,N_34254,N_39507);
and U46487 (N_46487,N_39568,N_32516);
or U46488 (N_46488,N_34795,N_38235);
xor U46489 (N_46489,N_36634,N_30239);
nor U46490 (N_46490,N_32447,N_38508);
xor U46491 (N_46491,N_36062,N_36031);
or U46492 (N_46492,N_39652,N_34186);
nor U46493 (N_46493,N_39127,N_33478);
nor U46494 (N_46494,N_34878,N_31132);
nor U46495 (N_46495,N_31060,N_33425);
or U46496 (N_46496,N_36559,N_37443);
and U46497 (N_46497,N_31669,N_31700);
nand U46498 (N_46498,N_34101,N_39948);
nand U46499 (N_46499,N_32045,N_38625);
or U46500 (N_46500,N_35322,N_35839);
and U46501 (N_46501,N_30469,N_36768);
nor U46502 (N_46502,N_37410,N_39743);
or U46503 (N_46503,N_33178,N_35784);
or U46504 (N_46504,N_39818,N_35765);
nor U46505 (N_46505,N_39808,N_39486);
xor U46506 (N_46506,N_35011,N_33744);
xor U46507 (N_46507,N_34407,N_37808);
and U46508 (N_46508,N_36289,N_35421);
xnor U46509 (N_46509,N_36861,N_38403);
nand U46510 (N_46510,N_33104,N_34017);
xnor U46511 (N_46511,N_38759,N_38644);
or U46512 (N_46512,N_30277,N_37080);
nand U46513 (N_46513,N_34990,N_34243);
and U46514 (N_46514,N_32433,N_32291);
or U46515 (N_46515,N_31235,N_37460);
and U46516 (N_46516,N_37970,N_37651);
nand U46517 (N_46517,N_35757,N_34140);
and U46518 (N_46518,N_32472,N_33233);
and U46519 (N_46519,N_34550,N_30550);
nor U46520 (N_46520,N_30342,N_37301);
xnor U46521 (N_46521,N_33011,N_36972);
xnor U46522 (N_46522,N_33540,N_36961);
xnor U46523 (N_46523,N_31703,N_35737);
xor U46524 (N_46524,N_32491,N_37061);
or U46525 (N_46525,N_36059,N_35454);
nand U46526 (N_46526,N_30440,N_33330);
nand U46527 (N_46527,N_35882,N_34241);
xnor U46528 (N_46528,N_35140,N_32435);
xnor U46529 (N_46529,N_30962,N_36036);
nand U46530 (N_46530,N_32024,N_39988);
xnor U46531 (N_46531,N_35618,N_39047);
or U46532 (N_46532,N_36630,N_31574);
nor U46533 (N_46533,N_37792,N_39395);
nand U46534 (N_46534,N_39641,N_33731);
nor U46535 (N_46535,N_32913,N_38780);
nor U46536 (N_46536,N_32107,N_37603);
and U46537 (N_46537,N_30922,N_39788);
nor U46538 (N_46538,N_39319,N_39845);
or U46539 (N_46539,N_34003,N_34115);
nor U46540 (N_46540,N_31962,N_37773);
nand U46541 (N_46541,N_33726,N_36981);
nand U46542 (N_46542,N_37799,N_35027);
nand U46543 (N_46543,N_32961,N_33768);
or U46544 (N_46544,N_31525,N_36159);
and U46545 (N_46545,N_37944,N_36806);
nor U46546 (N_46546,N_37557,N_39620);
nand U46547 (N_46547,N_30250,N_36889);
or U46548 (N_46548,N_39568,N_36834);
or U46549 (N_46549,N_38762,N_37825);
and U46550 (N_46550,N_32302,N_39256);
or U46551 (N_46551,N_36098,N_30676);
and U46552 (N_46552,N_36220,N_34542);
nor U46553 (N_46553,N_31413,N_33349);
xnor U46554 (N_46554,N_31582,N_30160);
nor U46555 (N_46555,N_31422,N_30238);
and U46556 (N_46556,N_38417,N_39243);
xor U46557 (N_46557,N_31865,N_37825);
and U46558 (N_46558,N_38280,N_34842);
and U46559 (N_46559,N_39433,N_35003);
nor U46560 (N_46560,N_39046,N_38986);
and U46561 (N_46561,N_38183,N_37627);
xor U46562 (N_46562,N_30737,N_33241);
or U46563 (N_46563,N_36982,N_34330);
xor U46564 (N_46564,N_37441,N_38446);
or U46565 (N_46565,N_37341,N_32066);
or U46566 (N_46566,N_31605,N_38489);
nor U46567 (N_46567,N_35107,N_37181);
or U46568 (N_46568,N_30183,N_31181);
xnor U46569 (N_46569,N_37160,N_36753);
and U46570 (N_46570,N_38997,N_30629);
or U46571 (N_46571,N_38348,N_38535);
nor U46572 (N_46572,N_37093,N_30499);
or U46573 (N_46573,N_30549,N_32008);
and U46574 (N_46574,N_38363,N_38104);
nor U46575 (N_46575,N_31794,N_32487);
nor U46576 (N_46576,N_33450,N_37156);
xor U46577 (N_46577,N_32894,N_35261);
and U46578 (N_46578,N_37379,N_31597);
or U46579 (N_46579,N_38777,N_36903);
xor U46580 (N_46580,N_37297,N_32064);
xnor U46581 (N_46581,N_31778,N_34552);
and U46582 (N_46582,N_36460,N_31001);
or U46583 (N_46583,N_37763,N_32737);
nand U46584 (N_46584,N_32885,N_38559);
nand U46585 (N_46585,N_32865,N_31005);
nand U46586 (N_46586,N_37319,N_39365);
nand U46587 (N_46587,N_36717,N_31709);
nor U46588 (N_46588,N_35499,N_33500);
nand U46589 (N_46589,N_34243,N_35247);
nor U46590 (N_46590,N_31823,N_32806);
nand U46591 (N_46591,N_34641,N_34071);
nand U46592 (N_46592,N_36615,N_39702);
nor U46593 (N_46593,N_34903,N_35854);
nand U46594 (N_46594,N_34092,N_33316);
and U46595 (N_46595,N_37590,N_34943);
nand U46596 (N_46596,N_36280,N_34212);
nand U46597 (N_46597,N_31986,N_35760);
xnor U46598 (N_46598,N_37690,N_31711);
nor U46599 (N_46599,N_39682,N_35538);
or U46600 (N_46600,N_33544,N_35108);
nand U46601 (N_46601,N_32951,N_33174);
or U46602 (N_46602,N_31817,N_34589);
and U46603 (N_46603,N_36429,N_39860);
nor U46604 (N_46604,N_39186,N_31865);
or U46605 (N_46605,N_36147,N_30262);
and U46606 (N_46606,N_30777,N_37334);
nor U46607 (N_46607,N_32407,N_33186);
xnor U46608 (N_46608,N_36515,N_31519);
and U46609 (N_46609,N_31518,N_33405);
nand U46610 (N_46610,N_37023,N_37270);
nor U46611 (N_46611,N_39881,N_39684);
xor U46612 (N_46612,N_33742,N_30798);
or U46613 (N_46613,N_39329,N_30561);
nand U46614 (N_46614,N_39231,N_32894);
and U46615 (N_46615,N_31571,N_30710);
or U46616 (N_46616,N_31231,N_34643);
and U46617 (N_46617,N_33901,N_39711);
xor U46618 (N_46618,N_34974,N_32540);
or U46619 (N_46619,N_39302,N_33032);
nand U46620 (N_46620,N_39093,N_35459);
nor U46621 (N_46621,N_39946,N_37205);
nor U46622 (N_46622,N_37974,N_39085);
and U46623 (N_46623,N_35780,N_34723);
nor U46624 (N_46624,N_31060,N_35351);
nand U46625 (N_46625,N_32354,N_30759);
or U46626 (N_46626,N_36973,N_31357);
and U46627 (N_46627,N_33960,N_32250);
xor U46628 (N_46628,N_30811,N_35522);
and U46629 (N_46629,N_31283,N_34990);
or U46630 (N_46630,N_36924,N_33321);
or U46631 (N_46631,N_34452,N_39471);
nand U46632 (N_46632,N_33390,N_32183);
nand U46633 (N_46633,N_32014,N_31253);
and U46634 (N_46634,N_31072,N_39119);
nor U46635 (N_46635,N_33651,N_39697);
xnor U46636 (N_46636,N_37622,N_39868);
nand U46637 (N_46637,N_34698,N_30351);
xnor U46638 (N_46638,N_35117,N_33988);
nor U46639 (N_46639,N_31643,N_39368);
nor U46640 (N_46640,N_31663,N_37414);
and U46641 (N_46641,N_39936,N_34658);
or U46642 (N_46642,N_37387,N_39711);
and U46643 (N_46643,N_34165,N_30663);
xnor U46644 (N_46644,N_36436,N_30158);
nand U46645 (N_46645,N_37037,N_34628);
nor U46646 (N_46646,N_30511,N_36939);
xnor U46647 (N_46647,N_33336,N_39291);
or U46648 (N_46648,N_33124,N_34156);
or U46649 (N_46649,N_34462,N_37359);
nand U46650 (N_46650,N_37248,N_30669);
and U46651 (N_46651,N_35073,N_32678);
xnor U46652 (N_46652,N_38168,N_34824);
xor U46653 (N_46653,N_33118,N_31696);
nor U46654 (N_46654,N_32852,N_32833);
xor U46655 (N_46655,N_30341,N_31371);
and U46656 (N_46656,N_30426,N_39185);
xnor U46657 (N_46657,N_33347,N_32064);
xnor U46658 (N_46658,N_38936,N_39479);
nor U46659 (N_46659,N_36275,N_39456);
or U46660 (N_46660,N_36547,N_38057);
or U46661 (N_46661,N_33545,N_34160);
nor U46662 (N_46662,N_34751,N_36090);
or U46663 (N_46663,N_37142,N_37232);
xor U46664 (N_46664,N_39815,N_35577);
xor U46665 (N_46665,N_38909,N_38987);
or U46666 (N_46666,N_35987,N_31318);
and U46667 (N_46667,N_39650,N_30904);
or U46668 (N_46668,N_38482,N_36242);
nor U46669 (N_46669,N_39178,N_34895);
and U46670 (N_46670,N_38276,N_36506);
nor U46671 (N_46671,N_33627,N_39209);
and U46672 (N_46672,N_34089,N_34456);
nor U46673 (N_46673,N_38260,N_36871);
or U46674 (N_46674,N_39449,N_30047);
and U46675 (N_46675,N_30971,N_32225);
or U46676 (N_46676,N_33252,N_38972);
xor U46677 (N_46677,N_38751,N_32220);
nor U46678 (N_46678,N_38229,N_35174);
xnor U46679 (N_46679,N_39693,N_39628);
nor U46680 (N_46680,N_38235,N_38616);
nand U46681 (N_46681,N_31001,N_37370);
nand U46682 (N_46682,N_30035,N_37078);
and U46683 (N_46683,N_33342,N_35449);
and U46684 (N_46684,N_32893,N_30393);
xor U46685 (N_46685,N_32205,N_30564);
and U46686 (N_46686,N_31860,N_31288);
xor U46687 (N_46687,N_31026,N_35309);
nor U46688 (N_46688,N_37805,N_39201);
nor U46689 (N_46689,N_35682,N_38704);
or U46690 (N_46690,N_36355,N_39338);
nand U46691 (N_46691,N_33670,N_36317);
and U46692 (N_46692,N_35811,N_34228);
or U46693 (N_46693,N_34549,N_30852);
or U46694 (N_46694,N_32292,N_35145);
and U46695 (N_46695,N_32342,N_36437);
nor U46696 (N_46696,N_32037,N_36137);
nand U46697 (N_46697,N_38522,N_34811);
and U46698 (N_46698,N_35884,N_39041);
or U46699 (N_46699,N_36336,N_38367);
xor U46700 (N_46700,N_32902,N_33358);
or U46701 (N_46701,N_37932,N_34755);
or U46702 (N_46702,N_34725,N_30154);
xnor U46703 (N_46703,N_31822,N_36196);
and U46704 (N_46704,N_39248,N_39569);
nand U46705 (N_46705,N_31180,N_31442);
xnor U46706 (N_46706,N_33235,N_35044);
nor U46707 (N_46707,N_34774,N_38811);
xnor U46708 (N_46708,N_32040,N_34897);
nor U46709 (N_46709,N_33841,N_37776);
xor U46710 (N_46710,N_32805,N_38981);
xnor U46711 (N_46711,N_31079,N_30309);
or U46712 (N_46712,N_33507,N_32202);
xor U46713 (N_46713,N_30534,N_32121);
nor U46714 (N_46714,N_35269,N_31272);
and U46715 (N_46715,N_36458,N_37460);
xor U46716 (N_46716,N_34879,N_37440);
and U46717 (N_46717,N_36141,N_36780);
nor U46718 (N_46718,N_36066,N_35709);
and U46719 (N_46719,N_36822,N_39925);
nor U46720 (N_46720,N_30998,N_39980);
and U46721 (N_46721,N_35509,N_31973);
nor U46722 (N_46722,N_30825,N_33160);
and U46723 (N_46723,N_36367,N_32001);
xor U46724 (N_46724,N_32629,N_38547);
xor U46725 (N_46725,N_30283,N_35460);
nand U46726 (N_46726,N_37392,N_38121);
xnor U46727 (N_46727,N_39509,N_31980);
xnor U46728 (N_46728,N_33476,N_35957);
nor U46729 (N_46729,N_39721,N_34503);
nor U46730 (N_46730,N_34719,N_34828);
nor U46731 (N_46731,N_38774,N_39235);
and U46732 (N_46732,N_35297,N_37861);
xnor U46733 (N_46733,N_35787,N_33972);
and U46734 (N_46734,N_38546,N_34678);
and U46735 (N_46735,N_35523,N_30975);
and U46736 (N_46736,N_36476,N_30146);
nor U46737 (N_46737,N_33446,N_32980);
or U46738 (N_46738,N_30373,N_30598);
nor U46739 (N_46739,N_30004,N_37522);
xnor U46740 (N_46740,N_32402,N_39773);
or U46741 (N_46741,N_39474,N_39709);
and U46742 (N_46742,N_31231,N_31877);
or U46743 (N_46743,N_39221,N_34502);
xnor U46744 (N_46744,N_34910,N_31695);
nand U46745 (N_46745,N_31583,N_38488);
and U46746 (N_46746,N_37272,N_38791);
xnor U46747 (N_46747,N_34752,N_32211);
xor U46748 (N_46748,N_31352,N_37353);
and U46749 (N_46749,N_36905,N_36502);
or U46750 (N_46750,N_37621,N_35651);
and U46751 (N_46751,N_36757,N_30872);
or U46752 (N_46752,N_39102,N_32469);
xnor U46753 (N_46753,N_37282,N_30043);
xnor U46754 (N_46754,N_33951,N_34082);
and U46755 (N_46755,N_39905,N_39297);
and U46756 (N_46756,N_38162,N_37839);
or U46757 (N_46757,N_32971,N_37455);
or U46758 (N_46758,N_35320,N_32647);
nor U46759 (N_46759,N_32773,N_38099);
nor U46760 (N_46760,N_33306,N_39487);
or U46761 (N_46761,N_32464,N_36502);
or U46762 (N_46762,N_35517,N_39158);
xnor U46763 (N_46763,N_35130,N_39090);
nor U46764 (N_46764,N_38259,N_37654);
or U46765 (N_46765,N_32150,N_31570);
xnor U46766 (N_46766,N_39045,N_32393);
nor U46767 (N_46767,N_34070,N_37866);
nand U46768 (N_46768,N_32129,N_34242);
nand U46769 (N_46769,N_34561,N_30845);
or U46770 (N_46770,N_37346,N_37531);
and U46771 (N_46771,N_35979,N_34340);
and U46772 (N_46772,N_31767,N_37331);
nand U46773 (N_46773,N_36575,N_39879);
or U46774 (N_46774,N_38976,N_30379);
xnor U46775 (N_46775,N_33377,N_35382);
nand U46776 (N_46776,N_38131,N_30819);
and U46777 (N_46777,N_36801,N_38644);
or U46778 (N_46778,N_33080,N_33861);
xnor U46779 (N_46779,N_31285,N_36019);
nand U46780 (N_46780,N_31800,N_32589);
xor U46781 (N_46781,N_37737,N_30454);
nor U46782 (N_46782,N_33564,N_31972);
xnor U46783 (N_46783,N_31469,N_34921);
nor U46784 (N_46784,N_39145,N_32176);
nor U46785 (N_46785,N_35721,N_37935);
nor U46786 (N_46786,N_34014,N_34103);
nand U46787 (N_46787,N_39617,N_39145);
or U46788 (N_46788,N_34330,N_34553);
and U46789 (N_46789,N_36144,N_34167);
nor U46790 (N_46790,N_35819,N_35512);
nand U46791 (N_46791,N_37531,N_36620);
and U46792 (N_46792,N_30878,N_36690);
xnor U46793 (N_46793,N_33013,N_36642);
nand U46794 (N_46794,N_34113,N_39308);
nor U46795 (N_46795,N_31323,N_36812);
xnor U46796 (N_46796,N_39849,N_38138);
nand U46797 (N_46797,N_39178,N_39092);
or U46798 (N_46798,N_31704,N_30888);
or U46799 (N_46799,N_35049,N_37706);
or U46800 (N_46800,N_36086,N_39276);
xor U46801 (N_46801,N_32007,N_32293);
or U46802 (N_46802,N_32915,N_36947);
xor U46803 (N_46803,N_37740,N_38169);
nand U46804 (N_46804,N_34665,N_31381);
or U46805 (N_46805,N_38462,N_35159);
or U46806 (N_46806,N_33351,N_37514);
nor U46807 (N_46807,N_32034,N_30117);
nor U46808 (N_46808,N_36377,N_33615);
xor U46809 (N_46809,N_36356,N_30406);
nand U46810 (N_46810,N_34983,N_32357);
and U46811 (N_46811,N_35982,N_38434);
and U46812 (N_46812,N_39026,N_31696);
and U46813 (N_46813,N_30011,N_33514);
or U46814 (N_46814,N_33655,N_39780);
or U46815 (N_46815,N_32105,N_34549);
xnor U46816 (N_46816,N_30549,N_32214);
or U46817 (N_46817,N_31095,N_34220);
and U46818 (N_46818,N_39816,N_32170);
or U46819 (N_46819,N_37450,N_37973);
and U46820 (N_46820,N_39386,N_34228);
nand U46821 (N_46821,N_36016,N_36671);
or U46822 (N_46822,N_38857,N_30046);
nor U46823 (N_46823,N_39461,N_35503);
nand U46824 (N_46824,N_39011,N_39355);
nor U46825 (N_46825,N_36792,N_39936);
or U46826 (N_46826,N_31264,N_37906);
nor U46827 (N_46827,N_35651,N_35802);
and U46828 (N_46828,N_30553,N_32043);
xnor U46829 (N_46829,N_38830,N_31082);
nand U46830 (N_46830,N_37012,N_36894);
nor U46831 (N_46831,N_35260,N_39810);
nand U46832 (N_46832,N_37915,N_32886);
xor U46833 (N_46833,N_31365,N_31124);
and U46834 (N_46834,N_37928,N_30050);
or U46835 (N_46835,N_32844,N_32403);
nand U46836 (N_46836,N_37577,N_32297);
nor U46837 (N_46837,N_31526,N_30657);
xnor U46838 (N_46838,N_32315,N_32255);
nand U46839 (N_46839,N_39391,N_32983);
nand U46840 (N_46840,N_39015,N_31522);
and U46841 (N_46841,N_30746,N_30701);
xnor U46842 (N_46842,N_34929,N_37721);
or U46843 (N_46843,N_36045,N_35420);
nand U46844 (N_46844,N_38443,N_35252);
nor U46845 (N_46845,N_31850,N_32045);
xnor U46846 (N_46846,N_37478,N_33781);
nand U46847 (N_46847,N_32947,N_32501);
and U46848 (N_46848,N_37485,N_32645);
or U46849 (N_46849,N_30027,N_34850);
xnor U46850 (N_46850,N_32503,N_34146);
and U46851 (N_46851,N_32022,N_37080);
or U46852 (N_46852,N_37859,N_37588);
nand U46853 (N_46853,N_36299,N_32503);
nand U46854 (N_46854,N_32245,N_37721);
nand U46855 (N_46855,N_34799,N_32511);
and U46856 (N_46856,N_33650,N_34148);
or U46857 (N_46857,N_38938,N_32254);
and U46858 (N_46858,N_39372,N_30992);
nor U46859 (N_46859,N_35395,N_36665);
xnor U46860 (N_46860,N_35365,N_31023);
nand U46861 (N_46861,N_38708,N_37575);
nand U46862 (N_46862,N_33553,N_38790);
and U46863 (N_46863,N_34821,N_31172);
or U46864 (N_46864,N_31584,N_35805);
xor U46865 (N_46865,N_31196,N_30589);
xor U46866 (N_46866,N_35777,N_34793);
nand U46867 (N_46867,N_30038,N_37249);
nand U46868 (N_46868,N_37952,N_34012);
nor U46869 (N_46869,N_38885,N_34436);
or U46870 (N_46870,N_31455,N_32021);
nand U46871 (N_46871,N_35771,N_32495);
nand U46872 (N_46872,N_32457,N_31259);
xor U46873 (N_46873,N_32463,N_35477);
xor U46874 (N_46874,N_39425,N_38929);
or U46875 (N_46875,N_37215,N_38793);
nand U46876 (N_46876,N_32841,N_39080);
or U46877 (N_46877,N_34717,N_30763);
nor U46878 (N_46878,N_30930,N_33883);
nand U46879 (N_46879,N_38086,N_33638);
xor U46880 (N_46880,N_33333,N_30672);
and U46881 (N_46881,N_39654,N_30397);
nor U46882 (N_46882,N_38117,N_38044);
or U46883 (N_46883,N_38123,N_33758);
nor U46884 (N_46884,N_38698,N_30457);
nor U46885 (N_46885,N_32561,N_33485);
nand U46886 (N_46886,N_37028,N_35953);
nor U46887 (N_46887,N_30966,N_39019);
nor U46888 (N_46888,N_31745,N_33491);
or U46889 (N_46889,N_31365,N_31356);
and U46890 (N_46890,N_32209,N_35007);
and U46891 (N_46891,N_38591,N_34146);
xor U46892 (N_46892,N_35594,N_32577);
nor U46893 (N_46893,N_37487,N_39171);
or U46894 (N_46894,N_39498,N_32954);
nand U46895 (N_46895,N_39717,N_31497);
nor U46896 (N_46896,N_30041,N_36285);
xnor U46897 (N_46897,N_31416,N_34537);
or U46898 (N_46898,N_35747,N_31594);
xor U46899 (N_46899,N_34443,N_30764);
nand U46900 (N_46900,N_36672,N_37545);
xnor U46901 (N_46901,N_34987,N_38280);
nand U46902 (N_46902,N_32385,N_30841);
nor U46903 (N_46903,N_37646,N_30588);
nand U46904 (N_46904,N_30168,N_37703);
or U46905 (N_46905,N_31653,N_38823);
and U46906 (N_46906,N_30238,N_33457);
nor U46907 (N_46907,N_32444,N_35297);
nand U46908 (N_46908,N_38981,N_39176);
nor U46909 (N_46909,N_35667,N_37960);
and U46910 (N_46910,N_33374,N_31380);
and U46911 (N_46911,N_38332,N_31857);
xor U46912 (N_46912,N_39519,N_39930);
or U46913 (N_46913,N_37200,N_32139);
nor U46914 (N_46914,N_35632,N_36318);
xor U46915 (N_46915,N_38388,N_34542);
xor U46916 (N_46916,N_31475,N_39310);
and U46917 (N_46917,N_33393,N_39561);
or U46918 (N_46918,N_37279,N_36721);
and U46919 (N_46919,N_30327,N_31259);
nor U46920 (N_46920,N_33756,N_30942);
nor U46921 (N_46921,N_39037,N_36386);
and U46922 (N_46922,N_32677,N_31523);
and U46923 (N_46923,N_30127,N_39070);
nand U46924 (N_46924,N_33524,N_34044);
nand U46925 (N_46925,N_34381,N_35729);
or U46926 (N_46926,N_30421,N_35227);
nand U46927 (N_46927,N_32739,N_33194);
nor U46928 (N_46928,N_32919,N_38633);
and U46929 (N_46929,N_35395,N_33118);
nand U46930 (N_46930,N_38350,N_37938);
xnor U46931 (N_46931,N_35218,N_33484);
xor U46932 (N_46932,N_35621,N_32005);
nor U46933 (N_46933,N_39235,N_35375);
nor U46934 (N_46934,N_32609,N_37325);
xnor U46935 (N_46935,N_34669,N_36872);
and U46936 (N_46936,N_34395,N_31659);
xor U46937 (N_46937,N_35907,N_35453);
nand U46938 (N_46938,N_34085,N_31928);
or U46939 (N_46939,N_31085,N_39076);
and U46940 (N_46940,N_37670,N_37631);
nand U46941 (N_46941,N_37373,N_32449);
or U46942 (N_46942,N_39406,N_32508);
nand U46943 (N_46943,N_37587,N_30266);
or U46944 (N_46944,N_35713,N_31646);
and U46945 (N_46945,N_32592,N_39791);
nand U46946 (N_46946,N_30874,N_30765);
xnor U46947 (N_46947,N_30583,N_33562);
or U46948 (N_46948,N_38730,N_36487);
or U46949 (N_46949,N_33259,N_31381);
xnor U46950 (N_46950,N_31142,N_35574);
or U46951 (N_46951,N_38238,N_35083);
or U46952 (N_46952,N_39723,N_36035);
nor U46953 (N_46953,N_30505,N_39383);
xnor U46954 (N_46954,N_37225,N_37840);
or U46955 (N_46955,N_33721,N_39196);
and U46956 (N_46956,N_33771,N_36471);
nand U46957 (N_46957,N_34538,N_37709);
nor U46958 (N_46958,N_35604,N_37544);
nor U46959 (N_46959,N_36264,N_31223);
nor U46960 (N_46960,N_33580,N_35353);
or U46961 (N_46961,N_35795,N_36497);
nand U46962 (N_46962,N_35385,N_34785);
xnor U46963 (N_46963,N_34637,N_34899);
and U46964 (N_46964,N_32087,N_35133);
and U46965 (N_46965,N_32954,N_36619);
and U46966 (N_46966,N_32274,N_32362);
nor U46967 (N_46967,N_36930,N_36274);
or U46968 (N_46968,N_39747,N_34630);
xnor U46969 (N_46969,N_32792,N_35587);
nor U46970 (N_46970,N_36006,N_35619);
nand U46971 (N_46971,N_35901,N_37335);
and U46972 (N_46972,N_34942,N_32840);
nor U46973 (N_46973,N_33262,N_35067);
nand U46974 (N_46974,N_35812,N_33182);
nand U46975 (N_46975,N_34864,N_39582);
xnor U46976 (N_46976,N_38432,N_32736);
or U46977 (N_46977,N_37229,N_39222);
and U46978 (N_46978,N_32529,N_38179);
nand U46979 (N_46979,N_33951,N_31529);
nor U46980 (N_46980,N_31969,N_35640);
nor U46981 (N_46981,N_30257,N_35904);
or U46982 (N_46982,N_35995,N_36941);
and U46983 (N_46983,N_32255,N_34794);
nor U46984 (N_46984,N_38145,N_35481);
nand U46985 (N_46985,N_31210,N_31880);
and U46986 (N_46986,N_37501,N_36378);
and U46987 (N_46987,N_35634,N_39813);
nand U46988 (N_46988,N_30650,N_30022);
and U46989 (N_46989,N_30487,N_35118);
nor U46990 (N_46990,N_38418,N_34159);
and U46991 (N_46991,N_37523,N_35523);
or U46992 (N_46992,N_32434,N_32217);
nand U46993 (N_46993,N_33425,N_31312);
nand U46994 (N_46994,N_31591,N_35070);
nor U46995 (N_46995,N_36236,N_33257);
nor U46996 (N_46996,N_39465,N_39367);
nand U46997 (N_46997,N_30449,N_31745);
or U46998 (N_46998,N_39210,N_31724);
and U46999 (N_46999,N_32502,N_37338);
xor U47000 (N_47000,N_37924,N_34609);
nand U47001 (N_47001,N_36299,N_37080);
and U47002 (N_47002,N_37401,N_33600);
nor U47003 (N_47003,N_30699,N_30085);
nor U47004 (N_47004,N_37983,N_35824);
and U47005 (N_47005,N_32920,N_33692);
nor U47006 (N_47006,N_30208,N_34004);
xnor U47007 (N_47007,N_33815,N_35146);
nand U47008 (N_47008,N_35440,N_32635);
or U47009 (N_47009,N_33059,N_31883);
nand U47010 (N_47010,N_39127,N_36474);
nor U47011 (N_47011,N_35163,N_30688);
nor U47012 (N_47012,N_38662,N_38689);
nand U47013 (N_47013,N_32688,N_34517);
nand U47014 (N_47014,N_39065,N_39422);
or U47015 (N_47015,N_35170,N_33104);
and U47016 (N_47016,N_37452,N_35686);
and U47017 (N_47017,N_30247,N_36397);
or U47018 (N_47018,N_35056,N_35756);
or U47019 (N_47019,N_33890,N_37725);
nor U47020 (N_47020,N_36248,N_36464);
or U47021 (N_47021,N_39261,N_31909);
xor U47022 (N_47022,N_38534,N_37431);
or U47023 (N_47023,N_30494,N_37584);
and U47024 (N_47024,N_34773,N_33231);
nor U47025 (N_47025,N_31126,N_33295);
nor U47026 (N_47026,N_32069,N_30498);
or U47027 (N_47027,N_32858,N_34130);
nand U47028 (N_47028,N_34925,N_33649);
nand U47029 (N_47029,N_34824,N_36876);
and U47030 (N_47030,N_30946,N_37117);
xor U47031 (N_47031,N_37267,N_35078);
or U47032 (N_47032,N_31750,N_33212);
xnor U47033 (N_47033,N_30477,N_35330);
or U47034 (N_47034,N_39987,N_38548);
nor U47035 (N_47035,N_30088,N_35521);
or U47036 (N_47036,N_37421,N_38620);
nor U47037 (N_47037,N_34163,N_37664);
xor U47038 (N_47038,N_34664,N_36086);
nor U47039 (N_47039,N_36811,N_39328);
xnor U47040 (N_47040,N_34379,N_38102);
or U47041 (N_47041,N_30838,N_38957);
and U47042 (N_47042,N_30000,N_36955);
or U47043 (N_47043,N_35622,N_30531);
xnor U47044 (N_47044,N_39863,N_36593);
xnor U47045 (N_47045,N_38225,N_33949);
and U47046 (N_47046,N_37105,N_32934);
or U47047 (N_47047,N_31859,N_31395);
xor U47048 (N_47048,N_30977,N_37963);
or U47049 (N_47049,N_33883,N_32479);
or U47050 (N_47050,N_33554,N_39243);
nand U47051 (N_47051,N_36794,N_38062);
or U47052 (N_47052,N_36472,N_36610);
nand U47053 (N_47053,N_30903,N_33682);
and U47054 (N_47054,N_32981,N_35074);
or U47055 (N_47055,N_33102,N_34335);
nand U47056 (N_47056,N_36475,N_33024);
and U47057 (N_47057,N_33141,N_30471);
nand U47058 (N_47058,N_36229,N_30930);
or U47059 (N_47059,N_30138,N_31298);
nand U47060 (N_47060,N_31004,N_30863);
nor U47061 (N_47061,N_31593,N_30416);
or U47062 (N_47062,N_30366,N_30458);
nand U47063 (N_47063,N_38276,N_32520);
xor U47064 (N_47064,N_37606,N_37463);
or U47065 (N_47065,N_37129,N_39624);
nand U47066 (N_47066,N_33714,N_31082);
nor U47067 (N_47067,N_32770,N_35344);
and U47068 (N_47068,N_38035,N_33928);
xor U47069 (N_47069,N_33887,N_38103);
nand U47070 (N_47070,N_38178,N_37499);
nor U47071 (N_47071,N_32078,N_33380);
nor U47072 (N_47072,N_30746,N_37023);
or U47073 (N_47073,N_39748,N_36462);
nand U47074 (N_47074,N_38267,N_39761);
nor U47075 (N_47075,N_31122,N_34356);
nor U47076 (N_47076,N_38152,N_37430);
nand U47077 (N_47077,N_32095,N_39893);
and U47078 (N_47078,N_39975,N_38539);
nand U47079 (N_47079,N_39416,N_30018);
and U47080 (N_47080,N_30352,N_34632);
xnor U47081 (N_47081,N_30861,N_38837);
nor U47082 (N_47082,N_34488,N_36317);
xnor U47083 (N_47083,N_38770,N_37449);
nand U47084 (N_47084,N_33717,N_35468);
xnor U47085 (N_47085,N_30221,N_31534);
or U47086 (N_47086,N_34241,N_39719);
and U47087 (N_47087,N_31685,N_39926);
xnor U47088 (N_47088,N_37508,N_35689);
xor U47089 (N_47089,N_30352,N_34129);
nand U47090 (N_47090,N_31444,N_37678);
nor U47091 (N_47091,N_36220,N_36793);
and U47092 (N_47092,N_33630,N_39207);
and U47093 (N_47093,N_35656,N_35060);
nor U47094 (N_47094,N_38669,N_36914);
nor U47095 (N_47095,N_36596,N_30643);
or U47096 (N_47096,N_31328,N_33795);
xnor U47097 (N_47097,N_30084,N_34078);
nor U47098 (N_47098,N_31216,N_31537);
or U47099 (N_47099,N_38595,N_33609);
or U47100 (N_47100,N_39643,N_34462);
xnor U47101 (N_47101,N_38449,N_37332);
nor U47102 (N_47102,N_37615,N_30826);
or U47103 (N_47103,N_33152,N_32617);
nand U47104 (N_47104,N_35647,N_39408);
and U47105 (N_47105,N_39497,N_34056);
or U47106 (N_47106,N_32022,N_34677);
nand U47107 (N_47107,N_34675,N_31665);
or U47108 (N_47108,N_37574,N_38951);
nand U47109 (N_47109,N_31522,N_35818);
xnor U47110 (N_47110,N_33086,N_37475);
nand U47111 (N_47111,N_30324,N_33039);
xor U47112 (N_47112,N_30350,N_35638);
xnor U47113 (N_47113,N_38269,N_38705);
nor U47114 (N_47114,N_30348,N_30584);
and U47115 (N_47115,N_31413,N_39904);
nand U47116 (N_47116,N_30614,N_31989);
nand U47117 (N_47117,N_36210,N_30012);
nand U47118 (N_47118,N_30214,N_37526);
xor U47119 (N_47119,N_32300,N_31992);
nor U47120 (N_47120,N_30651,N_30615);
nand U47121 (N_47121,N_33466,N_38194);
xor U47122 (N_47122,N_36620,N_35172);
or U47123 (N_47123,N_34903,N_38481);
or U47124 (N_47124,N_33258,N_37657);
nor U47125 (N_47125,N_34512,N_39970);
or U47126 (N_47126,N_30653,N_31195);
nand U47127 (N_47127,N_33688,N_35704);
or U47128 (N_47128,N_33578,N_30799);
nand U47129 (N_47129,N_33005,N_37255);
or U47130 (N_47130,N_33174,N_31359);
xnor U47131 (N_47131,N_31023,N_38583);
and U47132 (N_47132,N_39420,N_34608);
nor U47133 (N_47133,N_37189,N_38464);
nor U47134 (N_47134,N_33910,N_32162);
nor U47135 (N_47135,N_39901,N_31472);
and U47136 (N_47136,N_36910,N_34610);
nor U47137 (N_47137,N_34289,N_31893);
nor U47138 (N_47138,N_37156,N_35812);
xnor U47139 (N_47139,N_35081,N_31050);
xnor U47140 (N_47140,N_39059,N_31737);
or U47141 (N_47141,N_37174,N_39388);
xor U47142 (N_47142,N_30733,N_33207);
and U47143 (N_47143,N_36103,N_33491);
nand U47144 (N_47144,N_38444,N_39125);
or U47145 (N_47145,N_36126,N_30578);
nand U47146 (N_47146,N_39284,N_37449);
nor U47147 (N_47147,N_36936,N_36489);
xor U47148 (N_47148,N_39060,N_35266);
xnor U47149 (N_47149,N_37675,N_39140);
or U47150 (N_47150,N_36462,N_33328);
nand U47151 (N_47151,N_37912,N_36822);
and U47152 (N_47152,N_35429,N_38559);
xnor U47153 (N_47153,N_39553,N_30404);
and U47154 (N_47154,N_39240,N_39189);
nor U47155 (N_47155,N_33760,N_33990);
and U47156 (N_47156,N_30341,N_36975);
or U47157 (N_47157,N_30022,N_36306);
and U47158 (N_47158,N_39855,N_33551);
xor U47159 (N_47159,N_35014,N_39893);
xor U47160 (N_47160,N_30062,N_33185);
or U47161 (N_47161,N_39183,N_37581);
or U47162 (N_47162,N_37665,N_30891);
nor U47163 (N_47163,N_36389,N_35905);
and U47164 (N_47164,N_38032,N_39360);
or U47165 (N_47165,N_35023,N_30924);
or U47166 (N_47166,N_38559,N_33214);
and U47167 (N_47167,N_34210,N_35900);
xnor U47168 (N_47168,N_39045,N_36271);
nor U47169 (N_47169,N_31440,N_31898);
and U47170 (N_47170,N_37656,N_32816);
xnor U47171 (N_47171,N_38620,N_34619);
or U47172 (N_47172,N_37497,N_36983);
nor U47173 (N_47173,N_34370,N_34625);
nor U47174 (N_47174,N_31232,N_37755);
xnor U47175 (N_47175,N_34331,N_32873);
nand U47176 (N_47176,N_39109,N_35229);
xnor U47177 (N_47177,N_32948,N_38575);
and U47178 (N_47178,N_30525,N_38414);
nand U47179 (N_47179,N_30957,N_37865);
nor U47180 (N_47180,N_38227,N_31822);
xnor U47181 (N_47181,N_33347,N_39494);
xor U47182 (N_47182,N_38012,N_35040);
and U47183 (N_47183,N_37978,N_37896);
and U47184 (N_47184,N_30721,N_34164);
and U47185 (N_47185,N_36057,N_31625);
or U47186 (N_47186,N_39188,N_32731);
nor U47187 (N_47187,N_30783,N_35699);
and U47188 (N_47188,N_32651,N_38782);
nand U47189 (N_47189,N_33768,N_33013);
and U47190 (N_47190,N_32251,N_34716);
nand U47191 (N_47191,N_33407,N_34883);
nand U47192 (N_47192,N_35603,N_30595);
nor U47193 (N_47193,N_37694,N_36861);
nand U47194 (N_47194,N_38082,N_33418);
nand U47195 (N_47195,N_30455,N_39660);
nand U47196 (N_47196,N_30552,N_35787);
or U47197 (N_47197,N_32661,N_33874);
and U47198 (N_47198,N_32826,N_39024);
or U47199 (N_47199,N_37486,N_36498);
nand U47200 (N_47200,N_34226,N_34212);
nor U47201 (N_47201,N_31721,N_37677);
xnor U47202 (N_47202,N_31958,N_35464);
nand U47203 (N_47203,N_37006,N_33077);
or U47204 (N_47204,N_38642,N_37156);
nor U47205 (N_47205,N_39669,N_37665);
nand U47206 (N_47206,N_32531,N_31143);
xnor U47207 (N_47207,N_39520,N_35478);
xor U47208 (N_47208,N_39948,N_39425);
or U47209 (N_47209,N_34502,N_38238);
or U47210 (N_47210,N_31430,N_31176);
and U47211 (N_47211,N_38487,N_39294);
and U47212 (N_47212,N_39167,N_32051);
nand U47213 (N_47213,N_37147,N_34429);
or U47214 (N_47214,N_31743,N_37728);
nor U47215 (N_47215,N_39960,N_35582);
xor U47216 (N_47216,N_32037,N_34920);
nand U47217 (N_47217,N_30576,N_32654);
xor U47218 (N_47218,N_33774,N_33249);
or U47219 (N_47219,N_32776,N_33741);
or U47220 (N_47220,N_34265,N_38228);
nor U47221 (N_47221,N_36086,N_39999);
nor U47222 (N_47222,N_31851,N_39607);
and U47223 (N_47223,N_36810,N_30040);
nand U47224 (N_47224,N_34993,N_39711);
nand U47225 (N_47225,N_32410,N_36003);
nor U47226 (N_47226,N_36291,N_37861);
xnor U47227 (N_47227,N_30479,N_30646);
and U47228 (N_47228,N_30627,N_35378);
nand U47229 (N_47229,N_39969,N_36642);
nor U47230 (N_47230,N_34001,N_39168);
nand U47231 (N_47231,N_33184,N_36421);
and U47232 (N_47232,N_32081,N_35187);
nand U47233 (N_47233,N_36865,N_37933);
xnor U47234 (N_47234,N_37057,N_34102);
and U47235 (N_47235,N_34377,N_35210);
xnor U47236 (N_47236,N_39746,N_33554);
nand U47237 (N_47237,N_38519,N_36014);
or U47238 (N_47238,N_34475,N_38445);
or U47239 (N_47239,N_36544,N_32029);
or U47240 (N_47240,N_35909,N_31735);
or U47241 (N_47241,N_35103,N_35070);
or U47242 (N_47242,N_39843,N_31317);
and U47243 (N_47243,N_36654,N_37988);
and U47244 (N_47244,N_36898,N_38215);
nor U47245 (N_47245,N_30461,N_35215);
xor U47246 (N_47246,N_34455,N_32309);
nand U47247 (N_47247,N_37889,N_39895);
nand U47248 (N_47248,N_36859,N_39591);
nor U47249 (N_47249,N_34956,N_31618);
nor U47250 (N_47250,N_30761,N_32829);
nand U47251 (N_47251,N_30065,N_30953);
or U47252 (N_47252,N_38598,N_39634);
nor U47253 (N_47253,N_32153,N_33692);
xnor U47254 (N_47254,N_30964,N_30487);
or U47255 (N_47255,N_31739,N_30946);
nand U47256 (N_47256,N_31339,N_36221);
xor U47257 (N_47257,N_35372,N_32236);
or U47258 (N_47258,N_35575,N_36896);
nor U47259 (N_47259,N_31423,N_32960);
xnor U47260 (N_47260,N_33998,N_35602);
and U47261 (N_47261,N_30832,N_34584);
nand U47262 (N_47262,N_32310,N_37309);
and U47263 (N_47263,N_38430,N_35408);
nand U47264 (N_47264,N_37897,N_32542);
nor U47265 (N_47265,N_39561,N_32495);
nand U47266 (N_47266,N_31759,N_31641);
nor U47267 (N_47267,N_39921,N_30442);
or U47268 (N_47268,N_33424,N_33940);
nor U47269 (N_47269,N_30793,N_30992);
xor U47270 (N_47270,N_31756,N_33126);
nand U47271 (N_47271,N_31536,N_39675);
nand U47272 (N_47272,N_35391,N_35306);
or U47273 (N_47273,N_39778,N_37852);
and U47274 (N_47274,N_37965,N_31685);
and U47275 (N_47275,N_39970,N_31342);
or U47276 (N_47276,N_37839,N_37926);
xnor U47277 (N_47277,N_33930,N_35407);
xnor U47278 (N_47278,N_31161,N_34909);
xnor U47279 (N_47279,N_36932,N_34209);
xor U47280 (N_47280,N_31380,N_39176);
and U47281 (N_47281,N_30427,N_34836);
nor U47282 (N_47282,N_37254,N_39582);
xor U47283 (N_47283,N_32907,N_35047);
nand U47284 (N_47284,N_37724,N_35127);
xor U47285 (N_47285,N_31072,N_36951);
or U47286 (N_47286,N_35471,N_32628);
and U47287 (N_47287,N_34540,N_32643);
xnor U47288 (N_47288,N_35364,N_34182);
nor U47289 (N_47289,N_33294,N_37139);
nand U47290 (N_47290,N_30367,N_30505);
or U47291 (N_47291,N_33819,N_32781);
xor U47292 (N_47292,N_34043,N_30342);
nand U47293 (N_47293,N_33465,N_30076);
xnor U47294 (N_47294,N_31374,N_38272);
and U47295 (N_47295,N_34345,N_34511);
nor U47296 (N_47296,N_35635,N_33008);
and U47297 (N_47297,N_30665,N_35813);
nand U47298 (N_47298,N_32016,N_30631);
nor U47299 (N_47299,N_33812,N_33972);
or U47300 (N_47300,N_36334,N_37924);
or U47301 (N_47301,N_32130,N_34304);
xnor U47302 (N_47302,N_35369,N_31409);
or U47303 (N_47303,N_31985,N_36445);
and U47304 (N_47304,N_37615,N_34142);
nor U47305 (N_47305,N_31174,N_38512);
or U47306 (N_47306,N_31792,N_32441);
xnor U47307 (N_47307,N_32074,N_34095);
or U47308 (N_47308,N_39878,N_36541);
or U47309 (N_47309,N_30697,N_34502);
or U47310 (N_47310,N_31011,N_37231);
or U47311 (N_47311,N_36606,N_33621);
nand U47312 (N_47312,N_39172,N_33922);
nor U47313 (N_47313,N_31669,N_30101);
and U47314 (N_47314,N_33942,N_36699);
xnor U47315 (N_47315,N_36988,N_36339);
nor U47316 (N_47316,N_35397,N_33453);
or U47317 (N_47317,N_32591,N_32262);
nor U47318 (N_47318,N_32235,N_35257);
nor U47319 (N_47319,N_31542,N_31093);
xnor U47320 (N_47320,N_34642,N_35091);
nor U47321 (N_47321,N_30317,N_32957);
and U47322 (N_47322,N_35707,N_32583);
xnor U47323 (N_47323,N_35646,N_33203);
xnor U47324 (N_47324,N_30977,N_37969);
xor U47325 (N_47325,N_36391,N_35437);
or U47326 (N_47326,N_35862,N_34782);
nand U47327 (N_47327,N_35320,N_34373);
nand U47328 (N_47328,N_37630,N_32885);
nor U47329 (N_47329,N_35039,N_30167);
nand U47330 (N_47330,N_31543,N_39597);
nor U47331 (N_47331,N_33747,N_35488);
or U47332 (N_47332,N_39018,N_35890);
xor U47333 (N_47333,N_39910,N_39363);
and U47334 (N_47334,N_34717,N_31172);
nor U47335 (N_47335,N_39587,N_33823);
nor U47336 (N_47336,N_35194,N_34690);
xnor U47337 (N_47337,N_36983,N_33239);
xor U47338 (N_47338,N_30388,N_38296);
or U47339 (N_47339,N_39733,N_33012);
nor U47340 (N_47340,N_38517,N_38108);
xnor U47341 (N_47341,N_31507,N_31646);
nor U47342 (N_47342,N_35794,N_30676);
nand U47343 (N_47343,N_30246,N_37298);
nand U47344 (N_47344,N_36663,N_38350);
nor U47345 (N_47345,N_32246,N_37813);
or U47346 (N_47346,N_35269,N_33628);
xor U47347 (N_47347,N_32365,N_32208);
nand U47348 (N_47348,N_30499,N_32803);
and U47349 (N_47349,N_32800,N_36890);
nand U47350 (N_47350,N_35447,N_31267);
xor U47351 (N_47351,N_35663,N_38023);
or U47352 (N_47352,N_30589,N_30363);
nand U47353 (N_47353,N_37550,N_36363);
xor U47354 (N_47354,N_30211,N_38434);
nor U47355 (N_47355,N_39339,N_33814);
nand U47356 (N_47356,N_35019,N_39242);
xnor U47357 (N_47357,N_34671,N_38755);
nand U47358 (N_47358,N_33603,N_39746);
xor U47359 (N_47359,N_33436,N_34866);
nor U47360 (N_47360,N_39044,N_32640);
nor U47361 (N_47361,N_39686,N_33455);
xnor U47362 (N_47362,N_30368,N_39221);
xnor U47363 (N_47363,N_37355,N_38327);
nor U47364 (N_47364,N_31238,N_35505);
or U47365 (N_47365,N_31159,N_39792);
and U47366 (N_47366,N_32784,N_30752);
xnor U47367 (N_47367,N_37056,N_32791);
xnor U47368 (N_47368,N_34645,N_38313);
xnor U47369 (N_47369,N_39804,N_33553);
and U47370 (N_47370,N_30368,N_32097);
or U47371 (N_47371,N_39704,N_36717);
xor U47372 (N_47372,N_34262,N_34875);
or U47373 (N_47373,N_39500,N_32538);
xnor U47374 (N_47374,N_36836,N_35116);
nor U47375 (N_47375,N_37988,N_32336);
xnor U47376 (N_47376,N_34432,N_31693);
and U47377 (N_47377,N_35209,N_39064);
xor U47378 (N_47378,N_32514,N_35114);
nand U47379 (N_47379,N_36277,N_39098);
nand U47380 (N_47380,N_31514,N_33161);
or U47381 (N_47381,N_34154,N_32096);
nor U47382 (N_47382,N_31210,N_32148);
nand U47383 (N_47383,N_37044,N_37932);
xor U47384 (N_47384,N_35227,N_31895);
nor U47385 (N_47385,N_34272,N_31842);
or U47386 (N_47386,N_39497,N_39318);
or U47387 (N_47387,N_32405,N_34743);
nand U47388 (N_47388,N_36097,N_37621);
nor U47389 (N_47389,N_38467,N_31309);
nand U47390 (N_47390,N_39233,N_38125);
or U47391 (N_47391,N_35491,N_37205);
xnor U47392 (N_47392,N_32979,N_36961);
nand U47393 (N_47393,N_35678,N_34709);
or U47394 (N_47394,N_38965,N_37152);
xor U47395 (N_47395,N_33835,N_34813);
nand U47396 (N_47396,N_37275,N_33813);
nor U47397 (N_47397,N_39192,N_36686);
or U47398 (N_47398,N_36337,N_36153);
xnor U47399 (N_47399,N_37672,N_35976);
xnor U47400 (N_47400,N_39649,N_33930);
nand U47401 (N_47401,N_39831,N_39012);
xnor U47402 (N_47402,N_39905,N_33023);
nor U47403 (N_47403,N_34383,N_38289);
and U47404 (N_47404,N_39095,N_30443);
xnor U47405 (N_47405,N_39002,N_30308);
nor U47406 (N_47406,N_36756,N_30978);
and U47407 (N_47407,N_37689,N_33540);
nor U47408 (N_47408,N_39565,N_35960);
nor U47409 (N_47409,N_35351,N_35644);
nor U47410 (N_47410,N_35890,N_37725);
and U47411 (N_47411,N_36628,N_34124);
and U47412 (N_47412,N_36350,N_33425);
and U47413 (N_47413,N_39042,N_36876);
xor U47414 (N_47414,N_35776,N_33031);
or U47415 (N_47415,N_35467,N_39286);
xor U47416 (N_47416,N_39764,N_30979);
or U47417 (N_47417,N_31560,N_39174);
nand U47418 (N_47418,N_38719,N_31085);
nand U47419 (N_47419,N_39984,N_39060);
nor U47420 (N_47420,N_31150,N_33366);
nand U47421 (N_47421,N_31791,N_39897);
nand U47422 (N_47422,N_33242,N_39718);
nand U47423 (N_47423,N_33854,N_37680);
and U47424 (N_47424,N_30389,N_30256);
or U47425 (N_47425,N_37211,N_36803);
and U47426 (N_47426,N_30270,N_31691);
nor U47427 (N_47427,N_32323,N_37874);
or U47428 (N_47428,N_34114,N_39503);
and U47429 (N_47429,N_32106,N_34795);
nand U47430 (N_47430,N_37625,N_36049);
xor U47431 (N_47431,N_34754,N_32313);
xnor U47432 (N_47432,N_36318,N_38091);
nor U47433 (N_47433,N_39000,N_36615);
or U47434 (N_47434,N_36635,N_35396);
and U47435 (N_47435,N_37976,N_37132);
or U47436 (N_47436,N_37298,N_39297);
nor U47437 (N_47437,N_34526,N_31996);
xnor U47438 (N_47438,N_39496,N_35815);
and U47439 (N_47439,N_31271,N_33915);
xnor U47440 (N_47440,N_33305,N_32924);
or U47441 (N_47441,N_37786,N_32481);
nand U47442 (N_47442,N_30681,N_36940);
or U47443 (N_47443,N_37076,N_38984);
and U47444 (N_47444,N_35169,N_31964);
and U47445 (N_47445,N_32451,N_31399);
and U47446 (N_47446,N_30288,N_38182);
or U47447 (N_47447,N_30877,N_33490);
and U47448 (N_47448,N_32269,N_31898);
and U47449 (N_47449,N_31094,N_31855);
nand U47450 (N_47450,N_38504,N_33050);
or U47451 (N_47451,N_31443,N_31729);
xnor U47452 (N_47452,N_36231,N_38100);
nand U47453 (N_47453,N_39094,N_37233);
xnor U47454 (N_47454,N_30265,N_30007);
and U47455 (N_47455,N_35218,N_33033);
xor U47456 (N_47456,N_33625,N_38187);
or U47457 (N_47457,N_35659,N_33861);
xor U47458 (N_47458,N_37256,N_37693);
and U47459 (N_47459,N_31199,N_37694);
and U47460 (N_47460,N_37829,N_37076);
nor U47461 (N_47461,N_36529,N_30929);
or U47462 (N_47462,N_34130,N_37790);
nand U47463 (N_47463,N_39126,N_31722);
or U47464 (N_47464,N_35779,N_32448);
xnor U47465 (N_47465,N_37113,N_30165);
or U47466 (N_47466,N_32187,N_35367);
nor U47467 (N_47467,N_34907,N_39111);
nor U47468 (N_47468,N_31982,N_37302);
and U47469 (N_47469,N_37832,N_31202);
nor U47470 (N_47470,N_36514,N_31105);
nor U47471 (N_47471,N_34855,N_38585);
nand U47472 (N_47472,N_39352,N_33505);
and U47473 (N_47473,N_32322,N_34405);
nor U47474 (N_47474,N_34677,N_38378);
or U47475 (N_47475,N_31606,N_33792);
nand U47476 (N_47476,N_33086,N_39707);
nand U47477 (N_47477,N_35684,N_31417);
and U47478 (N_47478,N_35147,N_30196);
xnor U47479 (N_47479,N_39749,N_32432);
or U47480 (N_47480,N_30644,N_35887);
nor U47481 (N_47481,N_38864,N_37298);
or U47482 (N_47482,N_38758,N_32947);
and U47483 (N_47483,N_32182,N_35773);
nand U47484 (N_47484,N_38190,N_34533);
nand U47485 (N_47485,N_31026,N_30933);
nor U47486 (N_47486,N_35999,N_33975);
xnor U47487 (N_47487,N_35611,N_38022);
or U47488 (N_47488,N_32466,N_39626);
or U47489 (N_47489,N_33295,N_31193);
nor U47490 (N_47490,N_30134,N_37030);
or U47491 (N_47491,N_33158,N_37232);
and U47492 (N_47492,N_35422,N_30199);
and U47493 (N_47493,N_38125,N_39910);
nand U47494 (N_47494,N_33346,N_33835);
and U47495 (N_47495,N_31077,N_30492);
nand U47496 (N_47496,N_30468,N_31413);
nand U47497 (N_47497,N_38837,N_38286);
nor U47498 (N_47498,N_37759,N_30523);
xor U47499 (N_47499,N_39245,N_39964);
nand U47500 (N_47500,N_30932,N_31030);
nor U47501 (N_47501,N_32212,N_38879);
nor U47502 (N_47502,N_32434,N_35043);
nor U47503 (N_47503,N_36665,N_37232);
xnor U47504 (N_47504,N_36699,N_33656);
nand U47505 (N_47505,N_35882,N_35013);
nor U47506 (N_47506,N_38206,N_30886);
xor U47507 (N_47507,N_36375,N_30714);
nand U47508 (N_47508,N_32790,N_37106);
nor U47509 (N_47509,N_35295,N_32616);
xor U47510 (N_47510,N_37601,N_39980);
nand U47511 (N_47511,N_31005,N_31736);
and U47512 (N_47512,N_33770,N_37811);
or U47513 (N_47513,N_30609,N_38430);
and U47514 (N_47514,N_34718,N_34833);
xnor U47515 (N_47515,N_33726,N_30941);
nand U47516 (N_47516,N_30714,N_35336);
and U47517 (N_47517,N_39133,N_33031);
and U47518 (N_47518,N_37332,N_32322);
nor U47519 (N_47519,N_32898,N_39801);
and U47520 (N_47520,N_31255,N_35172);
nand U47521 (N_47521,N_32422,N_30641);
and U47522 (N_47522,N_34071,N_33915);
and U47523 (N_47523,N_37363,N_32940);
and U47524 (N_47524,N_32238,N_33356);
nand U47525 (N_47525,N_36342,N_36156);
and U47526 (N_47526,N_39737,N_32731);
and U47527 (N_47527,N_37957,N_39408);
nand U47528 (N_47528,N_31331,N_33020);
and U47529 (N_47529,N_30128,N_38793);
xor U47530 (N_47530,N_35678,N_39687);
xnor U47531 (N_47531,N_36737,N_34531);
and U47532 (N_47532,N_32001,N_30393);
and U47533 (N_47533,N_30631,N_37113);
and U47534 (N_47534,N_35376,N_37655);
and U47535 (N_47535,N_35372,N_37063);
xnor U47536 (N_47536,N_31630,N_33363);
and U47537 (N_47537,N_38812,N_38778);
xnor U47538 (N_47538,N_31813,N_34906);
nor U47539 (N_47539,N_37552,N_39645);
nor U47540 (N_47540,N_30948,N_35180);
xnor U47541 (N_47541,N_32979,N_30217);
xnor U47542 (N_47542,N_32060,N_34177);
nor U47543 (N_47543,N_32529,N_32051);
nor U47544 (N_47544,N_31068,N_35144);
nand U47545 (N_47545,N_31929,N_33996);
xor U47546 (N_47546,N_37821,N_39238);
or U47547 (N_47547,N_38674,N_38655);
nor U47548 (N_47548,N_34525,N_34257);
nand U47549 (N_47549,N_31701,N_32644);
or U47550 (N_47550,N_36331,N_33173);
xnor U47551 (N_47551,N_39774,N_32896);
nor U47552 (N_47552,N_32521,N_30151);
xor U47553 (N_47553,N_38246,N_32725);
and U47554 (N_47554,N_33259,N_31383);
nand U47555 (N_47555,N_32280,N_39983);
or U47556 (N_47556,N_38921,N_32516);
or U47557 (N_47557,N_38830,N_34482);
nor U47558 (N_47558,N_35091,N_31723);
nand U47559 (N_47559,N_35045,N_35832);
and U47560 (N_47560,N_37962,N_34115);
xnor U47561 (N_47561,N_38173,N_30995);
nor U47562 (N_47562,N_36192,N_32581);
and U47563 (N_47563,N_32539,N_30613);
nand U47564 (N_47564,N_31076,N_34124);
nor U47565 (N_47565,N_32922,N_38915);
nor U47566 (N_47566,N_34445,N_33368);
and U47567 (N_47567,N_37781,N_31923);
and U47568 (N_47568,N_37050,N_36163);
nand U47569 (N_47569,N_30407,N_33317);
or U47570 (N_47570,N_39634,N_34894);
nand U47571 (N_47571,N_34092,N_39193);
or U47572 (N_47572,N_33056,N_38806);
nand U47573 (N_47573,N_36915,N_31635);
and U47574 (N_47574,N_38827,N_30294);
or U47575 (N_47575,N_39994,N_36525);
nor U47576 (N_47576,N_30279,N_34690);
and U47577 (N_47577,N_33723,N_39739);
xor U47578 (N_47578,N_33358,N_38141);
or U47579 (N_47579,N_33412,N_37994);
nand U47580 (N_47580,N_38971,N_32305);
nor U47581 (N_47581,N_37204,N_31280);
and U47582 (N_47582,N_38749,N_32667);
or U47583 (N_47583,N_34626,N_38685);
xor U47584 (N_47584,N_32199,N_38548);
nand U47585 (N_47585,N_33547,N_37221);
and U47586 (N_47586,N_30204,N_39662);
xor U47587 (N_47587,N_34292,N_31652);
nor U47588 (N_47588,N_32473,N_34874);
and U47589 (N_47589,N_36917,N_37300);
and U47590 (N_47590,N_33666,N_39322);
nand U47591 (N_47591,N_37133,N_36342);
and U47592 (N_47592,N_34800,N_37973);
and U47593 (N_47593,N_32529,N_39920);
or U47594 (N_47594,N_38843,N_31554);
xor U47595 (N_47595,N_34128,N_34166);
and U47596 (N_47596,N_34048,N_32867);
and U47597 (N_47597,N_35524,N_35970);
xnor U47598 (N_47598,N_37246,N_38922);
nor U47599 (N_47599,N_38582,N_38404);
xnor U47600 (N_47600,N_32282,N_37848);
or U47601 (N_47601,N_36725,N_32827);
xor U47602 (N_47602,N_34027,N_38699);
or U47603 (N_47603,N_36123,N_31158);
or U47604 (N_47604,N_32295,N_39057);
nor U47605 (N_47605,N_37301,N_39450);
xor U47606 (N_47606,N_35469,N_39524);
and U47607 (N_47607,N_38547,N_34167);
xnor U47608 (N_47608,N_37735,N_33302);
nand U47609 (N_47609,N_32754,N_32025);
nand U47610 (N_47610,N_36003,N_35309);
nand U47611 (N_47611,N_34175,N_31733);
nor U47612 (N_47612,N_39991,N_35260);
nor U47613 (N_47613,N_39219,N_39593);
xor U47614 (N_47614,N_35065,N_31535);
xnor U47615 (N_47615,N_36746,N_38691);
or U47616 (N_47616,N_39856,N_37547);
or U47617 (N_47617,N_32014,N_35922);
and U47618 (N_47618,N_33545,N_36274);
and U47619 (N_47619,N_38738,N_32497);
or U47620 (N_47620,N_39132,N_31439);
nor U47621 (N_47621,N_31662,N_35311);
or U47622 (N_47622,N_34767,N_32201);
or U47623 (N_47623,N_36065,N_32740);
xor U47624 (N_47624,N_35122,N_36098);
or U47625 (N_47625,N_34465,N_38372);
xnor U47626 (N_47626,N_37450,N_33171);
nand U47627 (N_47627,N_33405,N_31356);
xor U47628 (N_47628,N_38950,N_39215);
xor U47629 (N_47629,N_39996,N_32796);
xor U47630 (N_47630,N_30763,N_37790);
nor U47631 (N_47631,N_37081,N_31308);
nand U47632 (N_47632,N_35860,N_30680);
nor U47633 (N_47633,N_34229,N_30284);
and U47634 (N_47634,N_30304,N_32607);
or U47635 (N_47635,N_30083,N_36115);
and U47636 (N_47636,N_36055,N_32047);
and U47637 (N_47637,N_36847,N_35873);
and U47638 (N_47638,N_38678,N_34171);
nand U47639 (N_47639,N_31995,N_34777);
nand U47640 (N_47640,N_39925,N_36978);
and U47641 (N_47641,N_30972,N_37638);
or U47642 (N_47642,N_31158,N_31247);
nand U47643 (N_47643,N_34772,N_38134);
xnor U47644 (N_47644,N_39859,N_38236);
nand U47645 (N_47645,N_36343,N_37012);
and U47646 (N_47646,N_39404,N_31100);
nor U47647 (N_47647,N_37574,N_31818);
xnor U47648 (N_47648,N_33743,N_35225);
or U47649 (N_47649,N_35716,N_39984);
or U47650 (N_47650,N_30702,N_34277);
nor U47651 (N_47651,N_36965,N_30013);
and U47652 (N_47652,N_34643,N_32700);
nor U47653 (N_47653,N_32781,N_31089);
nor U47654 (N_47654,N_39671,N_32601);
nand U47655 (N_47655,N_34719,N_30015);
xnor U47656 (N_47656,N_33872,N_39681);
or U47657 (N_47657,N_34144,N_32194);
nor U47658 (N_47658,N_34713,N_39948);
or U47659 (N_47659,N_31268,N_39499);
nor U47660 (N_47660,N_36501,N_34299);
nor U47661 (N_47661,N_37016,N_30277);
nor U47662 (N_47662,N_32659,N_30431);
xnor U47663 (N_47663,N_32968,N_31272);
nand U47664 (N_47664,N_37790,N_36289);
nand U47665 (N_47665,N_30545,N_37978);
nor U47666 (N_47666,N_37007,N_34684);
or U47667 (N_47667,N_35353,N_30346);
nor U47668 (N_47668,N_39098,N_37541);
or U47669 (N_47669,N_38536,N_39619);
nand U47670 (N_47670,N_35853,N_39712);
nand U47671 (N_47671,N_34772,N_33528);
xor U47672 (N_47672,N_30715,N_32517);
and U47673 (N_47673,N_39926,N_35632);
xor U47674 (N_47674,N_34592,N_38210);
nand U47675 (N_47675,N_30269,N_38501);
or U47676 (N_47676,N_34834,N_37869);
and U47677 (N_47677,N_35819,N_36297);
and U47678 (N_47678,N_34799,N_35015);
and U47679 (N_47679,N_32993,N_37926);
or U47680 (N_47680,N_30072,N_35788);
nand U47681 (N_47681,N_35759,N_35967);
or U47682 (N_47682,N_38026,N_30542);
xnor U47683 (N_47683,N_36177,N_32905);
or U47684 (N_47684,N_37057,N_37279);
nand U47685 (N_47685,N_38695,N_35114);
xor U47686 (N_47686,N_31233,N_38710);
xor U47687 (N_47687,N_32118,N_37613);
xor U47688 (N_47688,N_36154,N_38867);
nor U47689 (N_47689,N_31418,N_34754);
xor U47690 (N_47690,N_32797,N_33017);
or U47691 (N_47691,N_35765,N_37993);
nand U47692 (N_47692,N_34891,N_31717);
or U47693 (N_47693,N_34905,N_39749);
nor U47694 (N_47694,N_30210,N_39598);
xor U47695 (N_47695,N_36261,N_33080);
nor U47696 (N_47696,N_32393,N_36980);
or U47697 (N_47697,N_37226,N_31692);
and U47698 (N_47698,N_34408,N_36023);
and U47699 (N_47699,N_31499,N_36246);
and U47700 (N_47700,N_35082,N_30081);
nor U47701 (N_47701,N_33017,N_31245);
nand U47702 (N_47702,N_37242,N_34308);
or U47703 (N_47703,N_34610,N_39892);
nor U47704 (N_47704,N_39695,N_33177);
or U47705 (N_47705,N_30158,N_36544);
or U47706 (N_47706,N_30751,N_30610);
and U47707 (N_47707,N_33998,N_39388);
nand U47708 (N_47708,N_36438,N_30519);
or U47709 (N_47709,N_35641,N_36621);
and U47710 (N_47710,N_33073,N_36336);
xnor U47711 (N_47711,N_34149,N_32307);
or U47712 (N_47712,N_38205,N_32895);
nand U47713 (N_47713,N_32063,N_31136);
or U47714 (N_47714,N_39176,N_36378);
and U47715 (N_47715,N_38181,N_30632);
and U47716 (N_47716,N_30569,N_31585);
and U47717 (N_47717,N_36303,N_35201);
nand U47718 (N_47718,N_35351,N_38063);
xor U47719 (N_47719,N_33931,N_38719);
and U47720 (N_47720,N_37777,N_38444);
nor U47721 (N_47721,N_37342,N_36858);
nand U47722 (N_47722,N_35398,N_35931);
or U47723 (N_47723,N_34469,N_38514);
xor U47724 (N_47724,N_39599,N_31538);
xnor U47725 (N_47725,N_36811,N_34131);
xor U47726 (N_47726,N_37934,N_38933);
or U47727 (N_47727,N_36427,N_37099);
or U47728 (N_47728,N_30797,N_32522);
or U47729 (N_47729,N_30827,N_31334);
nor U47730 (N_47730,N_39520,N_37682);
nand U47731 (N_47731,N_34550,N_33865);
xor U47732 (N_47732,N_33709,N_31188);
and U47733 (N_47733,N_34061,N_39933);
nor U47734 (N_47734,N_31126,N_33701);
or U47735 (N_47735,N_30696,N_32321);
nor U47736 (N_47736,N_38169,N_31835);
xor U47737 (N_47737,N_31578,N_32506);
nand U47738 (N_47738,N_31059,N_31076);
and U47739 (N_47739,N_35911,N_39073);
nor U47740 (N_47740,N_39420,N_36779);
nand U47741 (N_47741,N_39969,N_33364);
or U47742 (N_47742,N_31812,N_31954);
xor U47743 (N_47743,N_36152,N_35592);
and U47744 (N_47744,N_31447,N_33368);
or U47745 (N_47745,N_32235,N_38662);
nand U47746 (N_47746,N_33414,N_34433);
and U47747 (N_47747,N_33148,N_31278);
or U47748 (N_47748,N_38326,N_33952);
xnor U47749 (N_47749,N_30828,N_38445);
or U47750 (N_47750,N_34208,N_32455);
or U47751 (N_47751,N_37511,N_30615);
nand U47752 (N_47752,N_38137,N_37392);
and U47753 (N_47753,N_33088,N_32783);
or U47754 (N_47754,N_30912,N_34233);
nand U47755 (N_47755,N_30888,N_31937);
or U47756 (N_47756,N_35387,N_36653);
xor U47757 (N_47757,N_33543,N_37198);
nand U47758 (N_47758,N_33435,N_36650);
nor U47759 (N_47759,N_32036,N_30435);
or U47760 (N_47760,N_35461,N_35734);
nand U47761 (N_47761,N_38060,N_32031);
nand U47762 (N_47762,N_36459,N_34989);
nor U47763 (N_47763,N_34287,N_33153);
or U47764 (N_47764,N_33749,N_33390);
and U47765 (N_47765,N_33922,N_39939);
nand U47766 (N_47766,N_33646,N_38817);
nand U47767 (N_47767,N_31187,N_38271);
or U47768 (N_47768,N_37437,N_33976);
nand U47769 (N_47769,N_39676,N_35208);
xor U47770 (N_47770,N_36371,N_30024);
and U47771 (N_47771,N_39319,N_39351);
and U47772 (N_47772,N_31869,N_39989);
xor U47773 (N_47773,N_38020,N_33364);
xor U47774 (N_47774,N_31313,N_31693);
nand U47775 (N_47775,N_38336,N_37727);
xor U47776 (N_47776,N_38400,N_31737);
or U47777 (N_47777,N_33087,N_32770);
nand U47778 (N_47778,N_33064,N_33730);
or U47779 (N_47779,N_37262,N_30572);
and U47780 (N_47780,N_33133,N_35954);
xnor U47781 (N_47781,N_36552,N_38056);
nand U47782 (N_47782,N_35827,N_34167);
and U47783 (N_47783,N_37612,N_35865);
and U47784 (N_47784,N_32222,N_39172);
nor U47785 (N_47785,N_32659,N_38528);
nand U47786 (N_47786,N_35853,N_33156);
xnor U47787 (N_47787,N_37040,N_33871);
nand U47788 (N_47788,N_30823,N_37219);
xor U47789 (N_47789,N_30264,N_33604);
nor U47790 (N_47790,N_30472,N_33237);
nor U47791 (N_47791,N_38839,N_35656);
or U47792 (N_47792,N_34038,N_31974);
xor U47793 (N_47793,N_39421,N_36919);
and U47794 (N_47794,N_39950,N_37778);
nand U47795 (N_47795,N_31838,N_34760);
or U47796 (N_47796,N_35636,N_33615);
nand U47797 (N_47797,N_38207,N_38500);
or U47798 (N_47798,N_37281,N_32726);
and U47799 (N_47799,N_33311,N_32617);
or U47800 (N_47800,N_31445,N_39051);
or U47801 (N_47801,N_30580,N_36222);
nand U47802 (N_47802,N_38227,N_33806);
and U47803 (N_47803,N_33102,N_32976);
xnor U47804 (N_47804,N_34217,N_32757);
nand U47805 (N_47805,N_31056,N_33597);
and U47806 (N_47806,N_37132,N_32465);
or U47807 (N_47807,N_38141,N_31081);
xor U47808 (N_47808,N_37313,N_31277);
or U47809 (N_47809,N_34066,N_31148);
or U47810 (N_47810,N_34165,N_38266);
nand U47811 (N_47811,N_35119,N_36867);
nor U47812 (N_47812,N_32706,N_39801);
xnor U47813 (N_47813,N_34674,N_36530);
xor U47814 (N_47814,N_34863,N_31893);
nor U47815 (N_47815,N_33525,N_34668);
nand U47816 (N_47816,N_35829,N_36584);
nand U47817 (N_47817,N_37587,N_33461);
xnor U47818 (N_47818,N_37713,N_38759);
xnor U47819 (N_47819,N_35176,N_33235);
xor U47820 (N_47820,N_30655,N_32792);
nor U47821 (N_47821,N_38628,N_35203);
nand U47822 (N_47822,N_36873,N_38892);
xnor U47823 (N_47823,N_37830,N_30375);
xnor U47824 (N_47824,N_37379,N_35831);
or U47825 (N_47825,N_34760,N_38286);
nand U47826 (N_47826,N_30618,N_39442);
nand U47827 (N_47827,N_35226,N_30383);
and U47828 (N_47828,N_30349,N_37116);
nor U47829 (N_47829,N_39503,N_33067);
nand U47830 (N_47830,N_32534,N_34864);
nand U47831 (N_47831,N_34641,N_35289);
nand U47832 (N_47832,N_30454,N_33812);
and U47833 (N_47833,N_30351,N_30865);
and U47834 (N_47834,N_38174,N_33377);
and U47835 (N_47835,N_34279,N_35529);
nand U47836 (N_47836,N_32350,N_34422);
and U47837 (N_47837,N_37494,N_35014);
nand U47838 (N_47838,N_37754,N_34144);
and U47839 (N_47839,N_38114,N_37517);
nor U47840 (N_47840,N_39003,N_36373);
and U47841 (N_47841,N_39373,N_30576);
and U47842 (N_47842,N_39999,N_30841);
and U47843 (N_47843,N_34351,N_32790);
nand U47844 (N_47844,N_34310,N_34369);
nor U47845 (N_47845,N_36456,N_31189);
nand U47846 (N_47846,N_38648,N_36216);
or U47847 (N_47847,N_35060,N_38328);
xor U47848 (N_47848,N_36181,N_38666);
xor U47849 (N_47849,N_33499,N_36119);
nand U47850 (N_47850,N_37562,N_38437);
or U47851 (N_47851,N_34079,N_38548);
and U47852 (N_47852,N_30470,N_33807);
nor U47853 (N_47853,N_35602,N_39313);
or U47854 (N_47854,N_31796,N_38174);
nor U47855 (N_47855,N_35455,N_37355);
nand U47856 (N_47856,N_30148,N_39617);
xnor U47857 (N_47857,N_38282,N_32789);
or U47858 (N_47858,N_33315,N_32114);
or U47859 (N_47859,N_37316,N_38798);
nand U47860 (N_47860,N_33562,N_39255);
or U47861 (N_47861,N_30770,N_31917);
and U47862 (N_47862,N_34131,N_36614);
nor U47863 (N_47863,N_31256,N_39817);
nor U47864 (N_47864,N_38578,N_34715);
and U47865 (N_47865,N_31381,N_32777);
xnor U47866 (N_47866,N_30304,N_34260);
nand U47867 (N_47867,N_31842,N_37609);
and U47868 (N_47868,N_31899,N_30738);
and U47869 (N_47869,N_32788,N_37777);
nor U47870 (N_47870,N_35697,N_37282);
xnor U47871 (N_47871,N_34666,N_34519);
nand U47872 (N_47872,N_39883,N_39158);
or U47873 (N_47873,N_35883,N_35035);
nand U47874 (N_47874,N_31999,N_34301);
nand U47875 (N_47875,N_37506,N_31648);
nor U47876 (N_47876,N_38615,N_30358);
or U47877 (N_47877,N_35215,N_37659);
xnor U47878 (N_47878,N_30187,N_35817);
nor U47879 (N_47879,N_33520,N_35657);
nor U47880 (N_47880,N_35859,N_36075);
and U47881 (N_47881,N_33716,N_36914);
xnor U47882 (N_47882,N_39254,N_39320);
nor U47883 (N_47883,N_36249,N_39693);
and U47884 (N_47884,N_31947,N_38468);
nor U47885 (N_47885,N_35496,N_36357);
or U47886 (N_47886,N_33543,N_31927);
or U47887 (N_47887,N_37188,N_38140);
xnor U47888 (N_47888,N_39174,N_36950);
nand U47889 (N_47889,N_38769,N_31880);
nand U47890 (N_47890,N_37331,N_34064);
or U47891 (N_47891,N_39508,N_34723);
nor U47892 (N_47892,N_35713,N_36619);
nor U47893 (N_47893,N_39304,N_34238);
nand U47894 (N_47894,N_36965,N_30477);
or U47895 (N_47895,N_37564,N_33181);
and U47896 (N_47896,N_35801,N_37825);
xor U47897 (N_47897,N_33023,N_35863);
and U47898 (N_47898,N_32762,N_32105);
xor U47899 (N_47899,N_38362,N_33544);
and U47900 (N_47900,N_30191,N_38405);
xnor U47901 (N_47901,N_39014,N_30567);
and U47902 (N_47902,N_37373,N_35333);
nor U47903 (N_47903,N_38115,N_30529);
and U47904 (N_47904,N_30492,N_37479);
and U47905 (N_47905,N_30643,N_31578);
nor U47906 (N_47906,N_32127,N_33009);
nand U47907 (N_47907,N_37727,N_30100);
nor U47908 (N_47908,N_35444,N_38605);
or U47909 (N_47909,N_39115,N_39317);
or U47910 (N_47910,N_35659,N_38792);
nor U47911 (N_47911,N_30763,N_35758);
or U47912 (N_47912,N_32235,N_38137);
and U47913 (N_47913,N_35707,N_32568);
nand U47914 (N_47914,N_36253,N_35951);
xnor U47915 (N_47915,N_30877,N_35255);
or U47916 (N_47916,N_31644,N_39369);
xnor U47917 (N_47917,N_37791,N_30627);
xnor U47918 (N_47918,N_37183,N_38245);
or U47919 (N_47919,N_31266,N_35389);
nor U47920 (N_47920,N_34452,N_39803);
nand U47921 (N_47921,N_34733,N_30407);
and U47922 (N_47922,N_31431,N_32341);
nand U47923 (N_47923,N_35646,N_37657);
nand U47924 (N_47924,N_35650,N_39488);
nor U47925 (N_47925,N_37121,N_39486);
xnor U47926 (N_47926,N_35222,N_33340);
xnor U47927 (N_47927,N_36931,N_35319);
or U47928 (N_47928,N_35575,N_38018);
nand U47929 (N_47929,N_38138,N_35060);
or U47930 (N_47930,N_37877,N_31874);
xnor U47931 (N_47931,N_32360,N_38240);
and U47932 (N_47932,N_38269,N_34564);
and U47933 (N_47933,N_34319,N_37503);
nor U47934 (N_47934,N_32852,N_36274);
nand U47935 (N_47935,N_36634,N_39899);
xnor U47936 (N_47936,N_35472,N_35574);
xor U47937 (N_47937,N_38558,N_32885);
nand U47938 (N_47938,N_36657,N_38393);
xnor U47939 (N_47939,N_37244,N_35563);
nand U47940 (N_47940,N_38261,N_39091);
and U47941 (N_47941,N_32341,N_30237);
nor U47942 (N_47942,N_32793,N_35672);
nand U47943 (N_47943,N_38443,N_39236);
nor U47944 (N_47944,N_39818,N_37517);
or U47945 (N_47945,N_38662,N_35049);
or U47946 (N_47946,N_31959,N_39633);
and U47947 (N_47947,N_37195,N_30776);
and U47948 (N_47948,N_32823,N_33638);
nand U47949 (N_47949,N_30772,N_33644);
nor U47950 (N_47950,N_38109,N_32680);
nand U47951 (N_47951,N_38348,N_32525);
nor U47952 (N_47952,N_30963,N_33613);
or U47953 (N_47953,N_30215,N_39597);
nand U47954 (N_47954,N_32809,N_39017);
nand U47955 (N_47955,N_33450,N_38311);
nand U47956 (N_47956,N_35377,N_37592);
xor U47957 (N_47957,N_33935,N_37289);
and U47958 (N_47958,N_32297,N_32377);
and U47959 (N_47959,N_33735,N_31839);
and U47960 (N_47960,N_38853,N_35747);
xor U47961 (N_47961,N_33988,N_33623);
and U47962 (N_47962,N_34022,N_33176);
xnor U47963 (N_47963,N_33613,N_35927);
nand U47964 (N_47964,N_32164,N_37231);
or U47965 (N_47965,N_30788,N_33306);
nand U47966 (N_47966,N_39452,N_37504);
xnor U47967 (N_47967,N_34146,N_30331);
xnor U47968 (N_47968,N_31943,N_32743);
or U47969 (N_47969,N_34915,N_31236);
nor U47970 (N_47970,N_30178,N_30019);
nor U47971 (N_47971,N_30144,N_38175);
or U47972 (N_47972,N_35126,N_31713);
xor U47973 (N_47973,N_32507,N_38929);
nand U47974 (N_47974,N_33108,N_37751);
or U47975 (N_47975,N_36226,N_38969);
xor U47976 (N_47976,N_33582,N_31055);
nand U47977 (N_47977,N_32182,N_39622);
nor U47978 (N_47978,N_34206,N_31792);
xnor U47979 (N_47979,N_36401,N_37717);
nand U47980 (N_47980,N_33768,N_38646);
or U47981 (N_47981,N_32641,N_33449);
xnor U47982 (N_47982,N_37102,N_38260);
nand U47983 (N_47983,N_30623,N_30783);
xnor U47984 (N_47984,N_39461,N_33118);
and U47985 (N_47985,N_33518,N_39903);
xnor U47986 (N_47986,N_38581,N_39161);
and U47987 (N_47987,N_37440,N_30427);
nand U47988 (N_47988,N_32748,N_34439);
xnor U47989 (N_47989,N_30412,N_35320);
nor U47990 (N_47990,N_37447,N_36043);
xor U47991 (N_47991,N_30250,N_39800);
nand U47992 (N_47992,N_33885,N_30576);
nand U47993 (N_47993,N_35342,N_39127);
nand U47994 (N_47994,N_30418,N_35157);
nor U47995 (N_47995,N_30877,N_37204);
xor U47996 (N_47996,N_39869,N_33550);
and U47997 (N_47997,N_36621,N_30633);
and U47998 (N_47998,N_36221,N_38524);
or U47999 (N_47999,N_31910,N_36121);
nor U48000 (N_48000,N_33623,N_39848);
and U48001 (N_48001,N_38951,N_39611);
and U48002 (N_48002,N_34679,N_38841);
nand U48003 (N_48003,N_32055,N_30577);
and U48004 (N_48004,N_38273,N_38791);
xor U48005 (N_48005,N_34063,N_30135);
or U48006 (N_48006,N_33427,N_30231);
or U48007 (N_48007,N_33644,N_30917);
and U48008 (N_48008,N_32264,N_35377);
and U48009 (N_48009,N_37695,N_39400);
or U48010 (N_48010,N_30877,N_36002);
nor U48011 (N_48011,N_39720,N_33222);
or U48012 (N_48012,N_38415,N_39341);
nand U48013 (N_48013,N_32806,N_36991);
xnor U48014 (N_48014,N_34725,N_35630);
nor U48015 (N_48015,N_32207,N_30375);
nor U48016 (N_48016,N_32773,N_39281);
or U48017 (N_48017,N_38918,N_36701);
or U48018 (N_48018,N_37668,N_32225);
or U48019 (N_48019,N_35146,N_37546);
nor U48020 (N_48020,N_36000,N_35006);
or U48021 (N_48021,N_38685,N_39494);
xnor U48022 (N_48022,N_32288,N_36184);
and U48023 (N_48023,N_37384,N_31884);
and U48024 (N_48024,N_33820,N_36526);
and U48025 (N_48025,N_34610,N_32128);
nand U48026 (N_48026,N_37865,N_38998);
and U48027 (N_48027,N_38861,N_30832);
and U48028 (N_48028,N_32804,N_37981);
nand U48029 (N_48029,N_33714,N_39665);
nor U48030 (N_48030,N_34793,N_39914);
nor U48031 (N_48031,N_37247,N_31964);
xor U48032 (N_48032,N_38935,N_37570);
and U48033 (N_48033,N_35251,N_34049);
nor U48034 (N_48034,N_37700,N_36610);
and U48035 (N_48035,N_33510,N_33958);
nand U48036 (N_48036,N_36193,N_37868);
nor U48037 (N_48037,N_37118,N_39490);
or U48038 (N_48038,N_38767,N_30694);
nand U48039 (N_48039,N_32202,N_32143);
xor U48040 (N_48040,N_38314,N_35453);
and U48041 (N_48041,N_32975,N_33639);
nand U48042 (N_48042,N_30914,N_39671);
or U48043 (N_48043,N_32976,N_30782);
xnor U48044 (N_48044,N_37232,N_36633);
and U48045 (N_48045,N_30110,N_33623);
or U48046 (N_48046,N_31781,N_32677);
or U48047 (N_48047,N_30284,N_34842);
nor U48048 (N_48048,N_35846,N_38970);
xnor U48049 (N_48049,N_35311,N_37598);
xor U48050 (N_48050,N_30854,N_36172);
and U48051 (N_48051,N_30986,N_32420);
nand U48052 (N_48052,N_39477,N_37006);
or U48053 (N_48053,N_38356,N_31578);
nor U48054 (N_48054,N_30015,N_31482);
and U48055 (N_48055,N_32000,N_37482);
and U48056 (N_48056,N_30882,N_37441);
xor U48057 (N_48057,N_39835,N_36130);
and U48058 (N_48058,N_39358,N_31527);
nor U48059 (N_48059,N_38614,N_33893);
and U48060 (N_48060,N_37338,N_35789);
or U48061 (N_48061,N_37264,N_39308);
nand U48062 (N_48062,N_34021,N_31920);
and U48063 (N_48063,N_34701,N_37957);
xnor U48064 (N_48064,N_38994,N_35692);
nand U48065 (N_48065,N_37697,N_35967);
xnor U48066 (N_48066,N_31179,N_30473);
and U48067 (N_48067,N_34740,N_32775);
xor U48068 (N_48068,N_39246,N_36815);
or U48069 (N_48069,N_34288,N_34440);
or U48070 (N_48070,N_37558,N_36633);
nand U48071 (N_48071,N_38883,N_34078);
xnor U48072 (N_48072,N_32504,N_32864);
nand U48073 (N_48073,N_39642,N_33949);
or U48074 (N_48074,N_39548,N_35232);
or U48075 (N_48075,N_35485,N_39802);
nand U48076 (N_48076,N_37776,N_32639);
xnor U48077 (N_48077,N_38986,N_34704);
and U48078 (N_48078,N_36974,N_35104);
nor U48079 (N_48079,N_32591,N_35004);
xor U48080 (N_48080,N_36758,N_36934);
nor U48081 (N_48081,N_31339,N_30917);
nand U48082 (N_48082,N_36557,N_33613);
nor U48083 (N_48083,N_37126,N_30322);
nor U48084 (N_48084,N_39859,N_39168);
xor U48085 (N_48085,N_34127,N_37847);
and U48086 (N_48086,N_34049,N_35492);
nand U48087 (N_48087,N_38000,N_35860);
nor U48088 (N_48088,N_37311,N_37427);
xor U48089 (N_48089,N_38484,N_30793);
nand U48090 (N_48090,N_38132,N_34986);
and U48091 (N_48091,N_36128,N_39779);
nor U48092 (N_48092,N_34007,N_37170);
nor U48093 (N_48093,N_33611,N_31986);
nand U48094 (N_48094,N_33160,N_32299);
nor U48095 (N_48095,N_30094,N_35839);
xnor U48096 (N_48096,N_31898,N_37798);
xor U48097 (N_48097,N_37493,N_35811);
xnor U48098 (N_48098,N_37649,N_38450);
and U48099 (N_48099,N_37239,N_36450);
nand U48100 (N_48100,N_32887,N_37575);
nor U48101 (N_48101,N_34400,N_33119);
and U48102 (N_48102,N_35419,N_37293);
nor U48103 (N_48103,N_30746,N_38552);
or U48104 (N_48104,N_31763,N_35760);
or U48105 (N_48105,N_31400,N_37431);
and U48106 (N_48106,N_33440,N_36725);
or U48107 (N_48107,N_30207,N_35568);
nand U48108 (N_48108,N_36629,N_32060);
nand U48109 (N_48109,N_38966,N_39688);
nand U48110 (N_48110,N_35591,N_36727);
xor U48111 (N_48111,N_37057,N_37989);
nand U48112 (N_48112,N_37888,N_37613);
or U48113 (N_48113,N_34021,N_38232);
or U48114 (N_48114,N_30735,N_39103);
and U48115 (N_48115,N_38065,N_35458);
nor U48116 (N_48116,N_37000,N_30204);
xnor U48117 (N_48117,N_35955,N_33218);
xor U48118 (N_48118,N_39852,N_34969);
nand U48119 (N_48119,N_33795,N_30754);
and U48120 (N_48120,N_39365,N_34527);
xnor U48121 (N_48121,N_35943,N_32411);
nand U48122 (N_48122,N_31702,N_32055);
or U48123 (N_48123,N_38369,N_39164);
and U48124 (N_48124,N_38259,N_37198);
xnor U48125 (N_48125,N_33714,N_36174);
nor U48126 (N_48126,N_30259,N_33005);
nor U48127 (N_48127,N_34135,N_36723);
nor U48128 (N_48128,N_34493,N_31060);
nand U48129 (N_48129,N_30790,N_37396);
or U48130 (N_48130,N_35202,N_36271);
and U48131 (N_48131,N_37663,N_35210);
xor U48132 (N_48132,N_32788,N_31461);
xnor U48133 (N_48133,N_32483,N_35390);
nand U48134 (N_48134,N_32434,N_37422);
xnor U48135 (N_48135,N_35711,N_33182);
nor U48136 (N_48136,N_32367,N_39116);
or U48137 (N_48137,N_31968,N_36078);
nand U48138 (N_48138,N_37944,N_33971);
nor U48139 (N_48139,N_32952,N_38275);
nand U48140 (N_48140,N_33576,N_31074);
nor U48141 (N_48141,N_36114,N_32099);
nand U48142 (N_48142,N_33383,N_38312);
xor U48143 (N_48143,N_35739,N_33238);
nand U48144 (N_48144,N_33813,N_31962);
xor U48145 (N_48145,N_37038,N_30944);
nand U48146 (N_48146,N_35815,N_39869);
or U48147 (N_48147,N_39569,N_31464);
nor U48148 (N_48148,N_31934,N_39749);
or U48149 (N_48149,N_39390,N_32339);
nor U48150 (N_48150,N_30446,N_31766);
or U48151 (N_48151,N_31199,N_36402);
and U48152 (N_48152,N_35574,N_35404);
and U48153 (N_48153,N_32720,N_33144);
nor U48154 (N_48154,N_31319,N_33523);
and U48155 (N_48155,N_38559,N_33158);
nor U48156 (N_48156,N_39534,N_39768);
or U48157 (N_48157,N_38480,N_33073);
and U48158 (N_48158,N_30919,N_34982);
nand U48159 (N_48159,N_34509,N_31457);
or U48160 (N_48160,N_39464,N_37396);
and U48161 (N_48161,N_33611,N_33707);
and U48162 (N_48162,N_35316,N_30993);
and U48163 (N_48163,N_35668,N_34201);
xor U48164 (N_48164,N_30117,N_35627);
xnor U48165 (N_48165,N_31475,N_32103);
nand U48166 (N_48166,N_39620,N_38891);
nand U48167 (N_48167,N_33131,N_32140);
nand U48168 (N_48168,N_34397,N_37296);
nand U48169 (N_48169,N_34211,N_38922);
and U48170 (N_48170,N_31708,N_30552);
or U48171 (N_48171,N_32960,N_38141);
xnor U48172 (N_48172,N_36741,N_38342);
or U48173 (N_48173,N_33511,N_30285);
and U48174 (N_48174,N_32072,N_34999);
xnor U48175 (N_48175,N_37307,N_37962);
nand U48176 (N_48176,N_31964,N_38359);
nor U48177 (N_48177,N_38753,N_30995);
nor U48178 (N_48178,N_33787,N_35175);
xnor U48179 (N_48179,N_30003,N_39193);
nor U48180 (N_48180,N_38161,N_35069);
nor U48181 (N_48181,N_35387,N_33313);
nor U48182 (N_48182,N_36187,N_38224);
xor U48183 (N_48183,N_37561,N_34587);
or U48184 (N_48184,N_32210,N_30362);
xnor U48185 (N_48185,N_31296,N_31092);
nor U48186 (N_48186,N_38308,N_33178);
nand U48187 (N_48187,N_39432,N_32363);
or U48188 (N_48188,N_39480,N_39491);
or U48189 (N_48189,N_32758,N_33058);
nor U48190 (N_48190,N_33959,N_32804);
or U48191 (N_48191,N_38985,N_35259);
nor U48192 (N_48192,N_34078,N_31274);
xor U48193 (N_48193,N_35672,N_32896);
nor U48194 (N_48194,N_33318,N_39780);
and U48195 (N_48195,N_39962,N_31271);
nand U48196 (N_48196,N_37197,N_34819);
or U48197 (N_48197,N_30639,N_37849);
nor U48198 (N_48198,N_34443,N_39114);
and U48199 (N_48199,N_39949,N_38100);
xor U48200 (N_48200,N_39245,N_35800);
or U48201 (N_48201,N_30378,N_33375);
and U48202 (N_48202,N_38926,N_36605);
and U48203 (N_48203,N_34373,N_34338);
xor U48204 (N_48204,N_36712,N_37880);
and U48205 (N_48205,N_35041,N_36686);
or U48206 (N_48206,N_39519,N_35236);
and U48207 (N_48207,N_31312,N_37642);
or U48208 (N_48208,N_33892,N_36372);
xor U48209 (N_48209,N_30994,N_31473);
xnor U48210 (N_48210,N_31795,N_35443);
or U48211 (N_48211,N_34129,N_38479);
and U48212 (N_48212,N_31973,N_35305);
and U48213 (N_48213,N_34272,N_30837);
nor U48214 (N_48214,N_33829,N_34759);
nor U48215 (N_48215,N_37252,N_30521);
nor U48216 (N_48216,N_36428,N_37864);
and U48217 (N_48217,N_38181,N_32853);
nand U48218 (N_48218,N_34719,N_30568);
nor U48219 (N_48219,N_37109,N_35962);
or U48220 (N_48220,N_32590,N_32133);
nand U48221 (N_48221,N_35430,N_33670);
xnor U48222 (N_48222,N_31889,N_38575);
and U48223 (N_48223,N_30314,N_37118);
xor U48224 (N_48224,N_33413,N_32741);
nand U48225 (N_48225,N_34166,N_38597);
or U48226 (N_48226,N_39197,N_36579);
nand U48227 (N_48227,N_37880,N_30276);
nor U48228 (N_48228,N_35907,N_39103);
nand U48229 (N_48229,N_31209,N_37152);
xor U48230 (N_48230,N_39741,N_37771);
and U48231 (N_48231,N_34542,N_39441);
xnor U48232 (N_48232,N_34370,N_34666);
xnor U48233 (N_48233,N_36077,N_36594);
or U48234 (N_48234,N_33783,N_32155);
xnor U48235 (N_48235,N_30251,N_34193);
xor U48236 (N_48236,N_37615,N_35651);
nand U48237 (N_48237,N_38086,N_33234);
nor U48238 (N_48238,N_32602,N_30434);
and U48239 (N_48239,N_33345,N_36796);
xor U48240 (N_48240,N_31080,N_38315);
nand U48241 (N_48241,N_33296,N_39882);
xor U48242 (N_48242,N_33118,N_38927);
and U48243 (N_48243,N_37521,N_37493);
and U48244 (N_48244,N_38987,N_36971);
nor U48245 (N_48245,N_32860,N_31416);
nand U48246 (N_48246,N_37350,N_36888);
or U48247 (N_48247,N_36003,N_37283);
or U48248 (N_48248,N_39427,N_32187);
nor U48249 (N_48249,N_33348,N_31317);
nor U48250 (N_48250,N_39496,N_34141);
nor U48251 (N_48251,N_32770,N_30568);
nor U48252 (N_48252,N_33167,N_31356);
or U48253 (N_48253,N_34786,N_34117);
nor U48254 (N_48254,N_34248,N_36342);
or U48255 (N_48255,N_36335,N_36784);
and U48256 (N_48256,N_35865,N_34372);
nor U48257 (N_48257,N_38194,N_37180);
xnor U48258 (N_48258,N_39328,N_33381);
nor U48259 (N_48259,N_33978,N_39684);
or U48260 (N_48260,N_30648,N_36444);
and U48261 (N_48261,N_38571,N_39734);
xor U48262 (N_48262,N_37119,N_30325);
xor U48263 (N_48263,N_34170,N_37362);
nor U48264 (N_48264,N_38755,N_32535);
nand U48265 (N_48265,N_32892,N_36509);
or U48266 (N_48266,N_34972,N_36731);
and U48267 (N_48267,N_30452,N_30418);
or U48268 (N_48268,N_32273,N_35937);
nor U48269 (N_48269,N_33249,N_36166);
nand U48270 (N_48270,N_31512,N_31098);
nor U48271 (N_48271,N_38718,N_33232);
or U48272 (N_48272,N_33860,N_39251);
or U48273 (N_48273,N_35993,N_38200);
nor U48274 (N_48274,N_39134,N_33578);
xnor U48275 (N_48275,N_30632,N_34397);
nor U48276 (N_48276,N_33374,N_31975);
xnor U48277 (N_48277,N_37355,N_33192);
xnor U48278 (N_48278,N_37067,N_36674);
nand U48279 (N_48279,N_31153,N_33669);
and U48280 (N_48280,N_36506,N_38512);
or U48281 (N_48281,N_38375,N_30018);
xnor U48282 (N_48282,N_30271,N_34711);
and U48283 (N_48283,N_33690,N_39939);
and U48284 (N_48284,N_38690,N_32558);
nor U48285 (N_48285,N_35567,N_32016);
nor U48286 (N_48286,N_39453,N_31085);
or U48287 (N_48287,N_35156,N_37628);
and U48288 (N_48288,N_39914,N_31367);
and U48289 (N_48289,N_31738,N_38850);
nand U48290 (N_48290,N_37985,N_36650);
nand U48291 (N_48291,N_36906,N_31732);
and U48292 (N_48292,N_33321,N_30977);
or U48293 (N_48293,N_32546,N_35943);
nor U48294 (N_48294,N_38376,N_34689);
xor U48295 (N_48295,N_30318,N_34066);
xnor U48296 (N_48296,N_37095,N_30009);
or U48297 (N_48297,N_33602,N_31640);
or U48298 (N_48298,N_30827,N_38835);
nor U48299 (N_48299,N_32003,N_37543);
xor U48300 (N_48300,N_38389,N_32319);
and U48301 (N_48301,N_31043,N_36600);
or U48302 (N_48302,N_32518,N_38156);
or U48303 (N_48303,N_31028,N_35801);
nand U48304 (N_48304,N_30383,N_38175);
or U48305 (N_48305,N_32712,N_34865);
nand U48306 (N_48306,N_36354,N_35652);
and U48307 (N_48307,N_32540,N_35522);
nand U48308 (N_48308,N_31330,N_32545);
xor U48309 (N_48309,N_37361,N_30846);
or U48310 (N_48310,N_34783,N_32902);
xor U48311 (N_48311,N_35298,N_38849);
nor U48312 (N_48312,N_34210,N_30556);
nor U48313 (N_48313,N_36359,N_37933);
nor U48314 (N_48314,N_37800,N_37260);
and U48315 (N_48315,N_39438,N_38645);
nand U48316 (N_48316,N_34694,N_30087);
and U48317 (N_48317,N_32091,N_30599);
or U48318 (N_48318,N_32214,N_31863);
xnor U48319 (N_48319,N_30334,N_34311);
and U48320 (N_48320,N_35960,N_37161);
nor U48321 (N_48321,N_31861,N_34001);
nor U48322 (N_48322,N_35084,N_33353);
or U48323 (N_48323,N_31626,N_31529);
or U48324 (N_48324,N_38329,N_30565);
xor U48325 (N_48325,N_33133,N_32379);
xnor U48326 (N_48326,N_37502,N_39607);
and U48327 (N_48327,N_31360,N_32997);
nand U48328 (N_48328,N_33293,N_39404);
or U48329 (N_48329,N_33019,N_34072);
or U48330 (N_48330,N_33092,N_33593);
nand U48331 (N_48331,N_30547,N_38329);
nor U48332 (N_48332,N_35262,N_31849);
or U48333 (N_48333,N_32425,N_38256);
and U48334 (N_48334,N_31118,N_32976);
or U48335 (N_48335,N_31057,N_38915);
xor U48336 (N_48336,N_39034,N_34135);
and U48337 (N_48337,N_36107,N_38859);
or U48338 (N_48338,N_31198,N_36525);
xnor U48339 (N_48339,N_35955,N_39940);
or U48340 (N_48340,N_36940,N_30497);
xnor U48341 (N_48341,N_34674,N_37646);
nor U48342 (N_48342,N_31905,N_38187);
and U48343 (N_48343,N_39043,N_38543);
nand U48344 (N_48344,N_34937,N_30772);
or U48345 (N_48345,N_33325,N_33581);
and U48346 (N_48346,N_31098,N_32283);
or U48347 (N_48347,N_35718,N_31220);
or U48348 (N_48348,N_33580,N_30385);
nor U48349 (N_48349,N_36193,N_32687);
or U48350 (N_48350,N_33135,N_36894);
xnor U48351 (N_48351,N_31207,N_32300);
nand U48352 (N_48352,N_38192,N_35148);
xnor U48353 (N_48353,N_33451,N_34622);
and U48354 (N_48354,N_31622,N_30060);
and U48355 (N_48355,N_36387,N_38486);
xor U48356 (N_48356,N_36546,N_31299);
nand U48357 (N_48357,N_32449,N_31279);
and U48358 (N_48358,N_32146,N_34153);
or U48359 (N_48359,N_39209,N_37892);
xnor U48360 (N_48360,N_38760,N_35436);
and U48361 (N_48361,N_31009,N_39946);
nand U48362 (N_48362,N_30494,N_38363);
xor U48363 (N_48363,N_33064,N_31301);
xnor U48364 (N_48364,N_34847,N_38574);
nand U48365 (N_48365,N_36189,N_38555);
xor U48366 (N_48366,N_30719,N_36300);
nor U48367 (N_48367,N_38760,N_36109);
nor U48368 (N_48368,N_36295,N_38187);
nor U48369 (N_48369,N_35159,N_35214);
nor U48370 (N_48370,N_31445,N_30768);
or U48371 (N_48371,N_32274,N_37419);
or U48372 (N_48372,N_36303,N_35153);
xnor U48373 (N_48373,N_34409,N_36281);
xor U48374 (N_48374,N_35419,N_33980);
and U48375 (N_48375,N_31087,N_31226);
nand U48376 (N_48376,N_34390,N_31740);
or U48377 (N_48377,N_34871,N_35951);
nor U48378 (N_48378,N_38833,N_32565);
xnor U48379 (N_48379,N_34040,N_30827);
and U48380 (N_48380,N_30672,N_34388);
nand U48381 (N_48381,N_36542,N_30502);
nor U48382 (N_48382,N_35360,N_39366);
nand U48383 (N_48383,N_38702,N_37503);
or U48384 (N_48384,N_33593,N_35998);
xnor U48385 (N_48385,N_33150,N_35704);
xnor U48386 (N_48386,N_35216,N_35191);
and U48387 (N_48387,N_34816,N_32158);
nand U48388 (N_48388,N_35934,N_39956);
and U48389 (N_48389,N_34066,N_36951);
nand U48390 (N_48390,N_38894,N_30307);
nor U48391 (N_48391,N_35427,N_31953);
or U48392 (N_48392,N_39348,N_32846);
or U48393 (N_48393,N_38763,N_32311);
or U48394 (N_48394,N_38137,N_38000);
nand U48395 (N_48395,N_35983,N_39401);
or U48396 (N_48396,N_35032,N_34583);
nand U48397 (N_48397,N_39474,N_33527);
or U48398 (N_48398,N_39413,N_32811);
or U48399 (N_48399,N_31142,N_30227);
nand U48400 (N_48400,N_32922,N_39557);
xnor U48401 (N_48401,N_36120,N_34983);
xor U48402 (N_48402,N_36639,N_39506);
nand U48403 (N_48403,N_30235,N_39523);
nor U48404 (N_48404,N_37941,N_35384);
nor U48405 (N_48405,N_34060,N_35920);
nor U48406 (N_48406,N_31658,N_33651);
or U48407 (N_48407,N_34721,N_32446);
nand U48408 (N_48408,N_33281,N_35041);
nand U48409 (N_48409,N_32963,N_31214);
nand U48410 (N_48410,N_33852,N_37974);
or U48411 (N_48411,N_37692,N_31450);
nor U48412 (N_48412,N_30306,N_31851);
nand U48413 (N_48413,N_35657,N_33974);
nor U48414 (N_48414,N_34108,N_37744);
xnor U48415 (N_48415,N_32038,N_37451);
xnor U48416 (N_48416,N_38500,N_30153);
and U48417 (N_48417,N_32595,N_37016);
or U48418 (N_48418,N_35380,N_31379);
xor U48419 (N_48419,N_38304,N_33105);
xor U48420 (N_48420,N_34424,N_37847);
or U48421 (N_48421,N_35361,N_32731);
xor U48422 (N_48422,N_34156,N_39702);
nand U48423 (N_48423,N_37908,N_39562);
or U48424 (N_48424,N_30745,N_39210);
xnor U48425 (N_48425,N_31566,N_35139);
and U48426 (N_48426,N_35461,N_34592);
nand U48427 (N_48427,N_31387,N_32901);
nand U48428 (N_48428,N_39306,N_39711);
or U48429 (N_48429,N_34663,N_36786);
xor U48430 (N_48430,N_37924,N_37980);
nand U48431 (N_48431,N_35866,N_32910);
and U48432 (N_48432,N_39365,N_32758);
nand U48433 (N_48433,N_31365,N_33154);
nor U48434 (N_48434,N_36074,N_31177);
xor U48435 (N_48435,N_32581,N_35556);
or U48436 (N_48436,N_38386,N_39943);
nor U48437 (N_48437,N_35398,N_33822);
and U48438 (N_48438,N_30083,N_34295);
nor U48439 (N_48439,N_33795,N_33384);
and U48440 (N_48440,N_37222,N_30164);
and U48441 (N_48441,N_37384,N_34985);
nand U48442 (N_48442,N_39191,N_35620);
and U48443 (N_48443,N_35154,N_35086);
xor U48444 (N_48444,N_39107,N_34788);
and U48445 (N_48445,N_37073,N_35665);
nand U48446 (N_48446,N_32211,N_32150);
and U48447 (N_48447,N_38939,N_36589);
nand U48448 (N_48448,N_34481,N_36034);
or U48449 (N_48449,N_33328,N_34285);
xnor U48450 (N_48450,N_35314,N_32455);
and U48451 (N_48451,N_31289,N_39682);
nand U48452 (N_48452,N_33557,N_38012);
and U48453 (N_48453,N_39723,N_36033);
or U48454 (N_48454,N_32376,N_35613);
or U48455 (N_48455,N_31829,N_33884);
xor U48456 (N_48456,N_35395,N_38576);
or U48457 (N_48457,N_34837,N_36267);
and U48458 (N_48458,N_30460,N_33171);
xnor U48459 (N_48459,N_37997,N_37383);
nand U48460 (N_48460,N_32572,N_32810);
or U48461 (N_48461,N_37820,N_37320);
or U48462 (N_48462,N_38051,N_38984);
nand U48463 (N_48463,N_36142,N_34886);
xnor U48464 (N_48464,N_35231,N_35917);
xnor U48465 (N_48465,N_38977,N_34624);
xor U48466 (N_48466,N_30757,N_34812);
nor U48467 (N_48467,N_37193,N_33118);
nand U48468 (N_48468,N_34608,N_30104);
nand U48469 (N_48469,N_38754,N_39141);
nand U48470 (N_48470,N_36355,N_39986);
and U48471 (N_48471,N_36061,N_30017);
nand U48472 (N_48472,N_38821,N_37272);
or U48473 (N_48473,N_36104,N_37918);
nor U48474 (N_48474,N_34665,N_35399);
or U48475 (N_48475,N_32282,N_30348);
or U48476 (N_48476,N_38172,N_35183);
nand U48477 (N_48477,N_36217,N_31947);
or U48478 (N_48478,N_30053,N_32338);
or U48479 (N_48479,N_36974,N_39165);
or U48480 (N_48480,N_39962,N_37181);
nor U48481 (N_48481,N_34369,N_33659);
nor U48482 (N_48482,N_39451,N_39411);
and U48483 (N_48483,N_36055,N_35412);
or U48484 (N_48484,N_37593,N_37033);
and U48485 (N_48485,N_37532,N_38636);
or U48486 (N_48486,N_31665,N_38951);
nor U48487 (N_48487,N_34459,N_34611);
or U48488 (N_48488,N_36289,N_39141);
or U48489 (N_48489,N_38082,N_38648);
nor U48490 (N_48490,N_37011,N_39429);
or U48491 (N_48491,N_34666,N_32153);
and U48492 (N_48492,N_38825,N_30182);
and U48493 (N_48493,N_33839,N_35146);
xor U48494 (N_48494,N_39515,N_36511);
nand U48495 (N_48495,N_37663,N_32326);
and U48496 (N_48496,N_30228,N_32521);
and U48497 (N_48497,N_30804,N_39163);
xor U48498 (N_48498,N_36740,N_34829);
nor U48499 (N_48499,N_37629,N_34592);
and U48500 (N_48500,N_37851,N_37067);
nand U48501 (N_48501,N_34978,N_38082);
and U48502 (N_48502,N_30525,N_33603);
and U48503 (N_48503,N_35847,N_36480);
or U48504 (N_48504,N_33135,N_30425);
nor U48505 (N_48505,N_32004,N_34309);
and U48506 (N_48506,N_38652,N_39124);
or U48507 (N_48507,N_38190,N_35898);
nor U48508 (N_48508,N_36358,N_34279);
and U48509 (N_48509,N_36992,N_34187);
xnor U48510 (N_48510,N_33593,N_39865);
xnor U48511 (N_48511,N_33861,N_34493);
and U48512 (N_48512,N_35883,N_35555);
and U48513 (N_48513,N_30573,N_30534);
or U48514 (N_48514,N_33993,N_38836);
nor U48515 (N_48515,N_36211,N_39849);
nor U48516 (N_48516,N_38595,N_31436);
nor U48517 (N_48517,N_32778,N_38142);
and U48518 (N_48518,N_30177,N_32126);
xor U48519 (N_48519,N_32648,N_36618);
and U48520 (N_48520,N_34874,N_34253);
nor U48521 (N_48521,N_32229,N_33447);
or U48522 (N_48522,N_30908,N_35106);
and U48523 (N_48523,N_37080,N_30122);
and U48524 (N_48524,N_34162,N_37681);
or U48525 (N_48525,N_36210,N_30403);
xor U48526 (N_48526,N_35685,N_37868);
and U48527 (N_48527,N_35205,N_32834);
or U48528 (N_48528,N_36314,N_31265);
nand U48529 (N_48529,N_34473,N_32931);
nand U48530 (N_48530,N_37369,N_35934);
and U48531 (N_48531,N_36839,N_30882);
or U48532 (N_48532,N_36993,N_30588);
nor U48533 (N_48533,N_32188,N_36449);
or U48534 (N_48534,N_31798,N_33467);
and U48535 (N_48535,N_36801,N_31128);
nor U48536 (N_48536,N_36811,N_39897);
xnor U48537 (N_48537,N_39902,N_37800);
nor U48538 (N_48538,N_37652,N_37288);
nor U48539 (N_48539,N_39545,N_30054);
or U48540 (N_48540,N_31197,N_38123);
nand U48541 (N_48541,N_31864,N_36316);
xor U48542 (N_48542,N_33223,N_30322);
and U48543 (N_48543,N_33516,N_33443);
nor U48544 (N_48544,N_34508,N_38743);
xor U48545 (N_48545,N_37153,N_34369);
or U48546 (N_48546,N_31115,N_39726);
and U48547 (N_48547,N_37017,N_31295);
or U48548 (N_48548,N_39617,N_31036);
nor U48549 (N_48549,N_38833,N_37259);
xor U48550 (N_48550,N_34854,N_31315);
and U48551 (N_48551,N_34813,N_36171);
or U48552 (N_48552,N_34851,N_34339);
and U48553 (N_48553,N_38255,N_30397);
nor U48554 (N_48554,N_39106,N_30710);
and U48555 (N_48555,N_37783,N_36904);
or U48556 (N_48556,N_35704,N_35943);
or U48557 (N_48557,N_33666,N_36629);
xor U48558 (N_48558,N_36259,N_34288);
or U48559 (N_48559,N_31749,N_35019);
nor U48560 (N_48560,N_36321,N_35822);
or U48561 (N_48561,N_39956,N_39428);
xnor U48562 (N_48562,N_30839,N_31360);
or U48563 (N_48563,N_30959,N_36361);
or U48564 (N_48564,N_35314,N_39274);
or U48565 (N_48565,N_31782,N_39118);
or U48566 (N_48566,N_39490,N_35913);
nor U48567 (N_48567,N_32863,N_38952);
xor U48568 (N_48568,N_33942,N_31441);
and U48569 (N_48569,N_37419,N_35843);
nor U48570 (N_48570,N_36277,N_32902);
or U48571 (N_48571,N_32890,N_32606);
nand U48572 (N_48572,N_32061,N_35304);
and U48573 (N_48573,N_37816,N_34296);
and U48574 (N_48574,N_37055,N_33276);
nand U48575 (N_48575,N_30900,N_38953);
and U48576 (N_48576,N_39089,N_35062);
nand U48577 (N_48577,N_38491,N_36626);
nand U48578 (N_48578,N_31102,N_34943);
and U48579 (N_48579,N_36019,N_31115);
nand U48580 (N_48580,N_39128,N_30351);
and U48581 (N_48581,N_35384,N_37367);
nand U48582 (N_48582,N_34429,N_30189);
nand U48583 (N_48583,N_30189,N_37963);
nand U48584 (N_48584,N_38650,N_39321);
or U48585 (N_48585,N_32731,N_33195);
and U48586 (N_48586,N_37094,N_30971);
nand U48587 (N_48587,N_37553,N_39972);
or U48588 (N_48588,N_36341,N_39007);
xnor U48589 (N_48589,N_34219,N_36624);
or U48590 (N_48590,N_39759,N_36981);
xor U48591 (N_48591,N_39485,N_31974);
or U48592 (N_48592,N_39130,N_36054);
and U48593 (N_48593,N_32471,N_31094);
and U48594 (N_48594,N_35739,N_34145);
nand U48595 (N_48595,N_31386,N_33732);
and U48596 (N_48596,N_31154,N_34540);
xor U48597 (N_48597,N_36968,N_39569);
or U48598 (N_48598,N_37967,N_32398);
xor U48599 (N_48599,N_37195,N_30886);
nor U48600 (N_48600,N_33401,N_32776);
nor U48601 (N_48601,N_36548,N_33359);
nand U48602 (N_48602,N_33539,N_37190);
or U48603 (N_48603,N_35530,N_30858);
and U48604 (N_48604,N_39975,N_31400);
nor U48605 (N_48605,N_32406,N_33296);
and U48606 (N_48606,N_34574,N_33423);
and U48607 (N_48607,N_39429,N_32574);
or U48608 (N_48608,N_33550,N_39953);
or U48609 (N_48609,N_36243,N_35323);
and U48610 (N_48610,N_34244,N_36243);
and U48611 (N_48611,N_30806,N_30886);
nand U48612 (N_48612,N_32814,N_31453);
nand U48613 (N_48613,N_38409,N_38880);
or U48614 (N_48614,N_32371,N_33970);
or U48615 (N_48615,N_38368,N_38593);
nand U48616 (N_48616,N_32698,N_35986);
nand U48617 (N_48617,N_34362,N_30323);
nand U48618 (N_48618,N_32811,N_39036);
nand U48619 (N_48619,N_30837,N_36525);
nor U48620 (N_48620,N_31899,N_31235);
and U48621 (N_48621,N_33941,N_31931);
or U48622 (N_48622,N_31700,N_37179);
or U48623 (N_48623,N_33052,N_37585);
xnor U48624 (N_48624,N_36700,N_36175);
nand U48625 (N_48625,N_37138,N_30396);
nand U48626 (N_48626,N_31542,N_36784);
or U48627 (N_48627,N_37563,N_32391);
xnor U48628 (N_48628,N_32490,N_33219);
and U48629 (N_48629,N_39840,N_37681);
nor U48630 (N_48630,N_36109,N_35077);
and U48631 (N_48631,N_36740,N_36205);
nand U48632 (N_48632,N_36070,N_38259);
or U48633 (N_48633,N_39173,N_34084);
and U48634 (N_48634,N_32823,N_30435);
nand U48635 (N_48635,N_35705,N_33286);
xnor U48636 (N_48636,N_36317,N_34392);
nor U48637 (N_48637,N_35755,N_33426);
nor U48638 (N_48638,N_37367,N_37022);
and U48639 (N_48639,N_34089,N_30520);
nor U48640 (N_48640,N_37023,N_32436);
nor U48641 (N_48641,N_31359,N_32795);
and U48642 (N_48642,N_35513,N_30199);
and U48643 (N_48643,N_34519,N_37458);
and U48644 (N_48644,N_38668,N_37191);
nand U48645 (N_48645,N_33764,N_35363);
xor U48646 (N_48646,N_34945,N_37996);
xnor U48647 (N_48647,N_36367,N_38645);
nand U48648 (N_48648,N_36949,N_30943);
nand U48649 (N_48649,N_38945,N_31845);
nor U48650 (N_48650,N_33604,N_39694);
nand U48651 (N_48651,N_31083,N_38700);
or U48652 (N_48652,N_35817,N_30207);
and U48653 (N_48653,N_37446,N_38283);
nor U48654 (N_48654,N_30435,N_37873);
nor U48655 (N_48655,N_35324,N_32291);
and U48656 (N_48656,N_32517,N_34274);
nand U48657 (N_48657,N_31493,N_32205);
or U48658 (N_48658,N_39924,N_30270);
xor U48659 (N_48659,N_36729,N_31826);
nand U48660 (N_48660,N_32449,N_34494);
nor U48661 (N_48661,N_39071,N_34736);
nor U48662 (N_48662,N_34372,N_36287);
nand U48663 (N_48663,N_34792,N_35069);
xor U48664 (N_48664,N_36892,N_34238);
and U48665 (N_48665,N_38316,N_33713);
xnor U48666 (N_48666,N_31951,N_35643);
nand U48667 (N_48667,N_34843,N_37496);
and U48668 (N_48668,N_37824,N_33866);
nor U48669 (N_48669,N_32844,N_30287);
and U48670 (N_48670,N_39406,N_35670);
xor U48671 (N_48671,N_34728,N_36759);
xnor U48672 (N_48672,N_33667,N_32810);
nor U48673 (N_48673,N_37837,N_39064);
xnor U48674 (N_48674,N_32393,N_32545);
xor U48675 (N_48675,N_32413,N_39709);
and U48676 (N_48676,N_36263,N_35839);
nand U48677 (N_48677,N_39001,N_35793);
nor U48678 (N_48678,N_39013,N_39038);
or U48679 (N_48679,N_33011,N_38329);
and U48680 (N_48680,N_33616,N_30497);
and U48681 (N_48681,N_35831,N_33687);
nor U48682 (N_48682,N_35727,N_30856);
nand U48683 (N_48683,N_31036,N_33270);
xnor U48684 (N_48684,N_38181,N_35956);
or U48685 (N_48685,N_30070,N_34764);
or U48686 (N_48686,N_33379,N_34715);
xor U48687 (N_48687,N_31008,N_37461);
nand U48688 (N_48688,N_36755,N_33596);
nand U48689 (N_48689,N_34721,N_35645);
and U48690 (N_48690,N_39023,N_35781);
or U48691 (N_48691,N_34266,N_36002);
and U48692 (N_48692,N_38959,N_30304);
nor U48693 (N_48693,N_38598,N_34128);
or U48694 (N_48694,N_36776,N_37226);
nand U48695 (N_48695,N_36453,N_36851);
xor U48696 (N_48696,N_30825,N_37555);
nor U48697 (N_48697,N_39219,N_37276);
or U48698 (N_48698,N_34530,N_31537);
nor U48699 (N_48699,N_33970,N_35759);
nand U48700 (N_48700,N_34014,N_36176);
xnor U48701 (N_48701,N_30711,N_37577);
and U48702 (N_48702,N_32213,N_36912);
nor U48703 (N_48703,N_30474,N_32484);
nand U48704 (N_48704,N_39811,N_34764);
and U48705 (N_48705,N_33562,N_32384);
or U48706 (N_48706,N_33160,N_39105);
or U48707 (N_48707,N_32828,N_31816);
nor U48708 (N_48708,N_39442,N_31944);
and U48709 (N_48709,N_39565,N_38927);
nand U48710 (N_48710,N_30591,N_32475);
and U48711 (N_48711,N_32756,N_30941);
or U48712 (N_48712,N_34923,N_37002);
xor U48713 (N_48713,N_32686,N_33539);
nand U48714 (N_48714,N_33067,N_33655);
xnor U48715 (N_48715,N_35654,N_39277);
and U48716 (N_48716,N_39194,N_36032);
nand U48717 (N_48717,N_32786,N_36607);
nand U48718 (N_48718,N_36957,N_32310);
and U48719 (N_48719,N_35579,N_39034);
nand U48720 (N_48720,N_30650,N_37963);
xor U48721 (N_48721,N_38639,N_31330);
nor U48722 (N_48722,N_33627,N_38498);
xor U48723 (N_48723,N_36631,N_38877);
nand U48724 (N_48724,N_30334,N_30156);
xor U48725 (N_48725,N_31508,N_36020);
nor U48726 (N_48726,N_38461,N_33149);
and U48727 (N_48727,N_35346,N_38061);
or U48728 (N_48728,N_31675,N_38163);
nor U48729 (N_48729,N_33455,N_33746);
nand U48730 (N_48730,N_34874,N_37789);
xnor U48731 (N_48731,N_35972,N_38094);
or U48732 (N_48732,N_38893,N_37902);
or U48733 (N_48733,N_30010,N_37410);
nand U48734 (N_48734,N_38281,N_39642);
nor U48735 (N_48735,N_36980,N_31589);
or U48736 (N_48736,N_31734,N_30317);
and U48737 (N_48737,N_30600,N_35224);
nand U48738 (N_48738,N_37014,N_32968);
xnor U48739 (N_48739,N_36902,N_33845);
nor U48740 (N_48740,N_33718,N_31340);
and U48741 (N_48741,N_33483,N_35139);
nand U48742 (N_48742,N_30093,N_36618);
or U48743 (N_48743,N_35534,N_35285);
and U48744 (N_48744,N_33786,N_33618);
and U48745 (N_48745,N_34627,N_34755);
and U48746 (N_48746,N_32582,N_36325);
xor U48747 (N_48747,N_36806,N_39529);
nor U48748 (N_48748,N_32321,N_37496);
and U48749 (N_48749,N_36454,N_36348);
and U48750 (N_48750,N_36335,N_32070);
or U48751 (N_48751,N_32926,N_37310);
nor U48752 (N_48752,N_30454,N_35226);
xor U48753 (N_48753,N_32101,N_32724);
and U48754 (N_48754,N_36989,N_36133);
or U48755 (N_48755,N_33618,N_31047);
or U48756 (N_48756,N_34926,N_35093);
nand U48757 (N_48757,N_37026,N_33253);
nor U48758 (N_48758,N_34656,N_34038);
or U48759 (N_48759,N_31903,N_33371);
xor U48760 (N_48760,N_35037,N_37574);
and U48761 (N_48761,N_33052,N_32146);
and U48762 (N_48762,N_32656,N_38975);
xor U48763 (N_48763,N_35754,N_36809);
xor U48764 (N_48764,N_38000,N_35286);
and U48765 (N_48765,N_36358,N_38835);
and U48766 (N_48766,N_30067,N_38375);
and U48767 (N_48767,N_32193,N_36146);
or U48768 (N_48768,N_36281,N_32451);
nor U48769 (N_48769,N_36975,N_30912);
or U48770 (N_48770,N_32998,N_33870);
or U48771 (N_48771,N_39081,N_34655);
xnor U48772 (N_48772,N_34042,N_31105);
nand U48773 (N_48773,N_38864,N_39359);
or U48774 (N_48774,N_31069,N_38738);
xnor U48775 (N_48775,N_30409,N_33012);
xor U48776 (N_48776,N_37784,N_39443);
or U48777 (N_48777,N_31745,N_37125);
or U48778 (N_48778,N_32597,N_32777);
nor U48779 (N_48779,N_31452,N_39690);
nor U48780 (N_48780,N_30773,N_32660);
or U48781 (N_48781,N_36786,N_34233);
xnor U48782 (N_48782,N_38638,N_33196);
and U48783 (N_48783,N_37902,N_37289);
or U48784 (N_48784,N_32773,N_34033);
nor U48785 (N_48785,N_34199,N_34390);
or U48786 (N_48786,N_39627,N_33458);
nand U48787 (N_48787,N_31555,N_33663);
nor U48788 (N_48788,N_30347,N_35592);
nand U48789 (N_48789,N_32910,N_38597);
xor U48790 (N_48790,N_39673,N_31464);
xnor U48791 (N_48791,N_37536,N_31533);
nand U48792 (N_48792,N_30571,N_34718);
nand U48793 (N_48793,N_33733,N_35950);
xnor U48794 (N_48794,N_36286,N_30995);
nor U48795 (N_48795,N_32500,N_31576);
nor U48796 (N_48796,N_34983,N_37251);
nand U48797 (N_48797,N_38745,N_32816);
xnor U48798 (N_48798,N_33225,N_37923);
nand U48799 (N_48799,N_31421,N_30082);
or U48800 (N_48800,N_38060,N_38591);
and U48801 (N_48801,N_34855,N_30880);
nor U48802 (N_48802,N_37440,N_33113);
nor U48803 (N_48803,N_33064,N_32272);
or U48804 (N_48804,N_33631,N_30224);
nor U48805 (N_48805,N_33120,N_33751);
xnor U48806 (N_48806,N_36815,N_35239);
nor U48807 (N_48807,N_30473,N_34030);
nor U48808 (N_48808,N_33756,N_39377);
or U48809 (N_48809,N_37068,N_39027);
nor U48810 (N_48810,N_34619,N_33066);
or U48811 (N_48811,N_39844,N_33907);
nand U48812 (N_48812,N_36274,N_34944);
xor U48813 (N_48813,N_32712,N_37824);
or U48814 (N_48814,N_39230,N_35961);
xor U48815 (N_48815,N_35500,N_38106);
nand U48816 (N_48816,N_38791,N_35378);
nand U48817 (N_48817,N_30161,N_32300);
or U48818 (N_48818,N_33937,N_37374);
nand U48819 (N_48819,N_37456,N_32277);
nor U48820 (N_48820,N_33036,N_30330);
nor U48821 (N_48821,N_37364,N_33727);
or U48822 (N_48822,N_38498,N_37041);
or U48823 (N_48823,N_30079,N_34524);
nor U48824 (N_48824,N_32301,N_39357);
or U48825 (N_48825,N_31662,N_37939);
xor U48826 (N_48826,N_39408,N_37887);
nor U48827 (N_48827,N_34975,N_35074);
and U48828 (N_48828,N_34517,N_35484);
xnor U48829 (N_48829,N_36235,N_37875);
and U48830 (N_48830,N_34866,N_35655);
nor U48831 (N_48831,N_32463,N_36875);
nand U48832 (N_48832,N_35477,N_31991);
xnor U48833 (N_48833,N_35331,N_34930);
and U48834 (N_48834,N_31117,N_31422);
or U48835 (N_48835,N_38915,N_30734);
xnor U48836 (N_48836,N_39566,N_33956);
and U48837 (N_48837,N_30607,N_30161);
xnor U48838 (N_48838,N_38239,N_30755);
nand U48839 (N_48839,N_31567,N_34737);
xor U48840 (N_48840,N_38283,N_30289);
xor U48841 (N_48841,N_31173,N_31264);
xor U48842 (N_48842,N_33437,N_35641);
and U48843 (N_48843,N_31370,N_30308);
or U48844 (N_48844,N_33345,N_31546);
nand U48845 (N_48845,N_37166,N_30312);
or U48846 (N_48846,N_39170,N_31745);
nand U48847 (N_48847,N_32458,N_33410);
or U48848 (N_48848,N_35815,N_34326);
or U48849 (N_48849,N_30397,N_37296);
nand U48850 (N_48850,N_35529,N_35811);
or U48851 (N_48851,N_36813,N_36316);
and U48852 (N_48852,N_30374,N_34442);
or U48853 (N_48853,N_32021,N_31879);
nand U48854 (N_48854,N_37979,N_34904);
nand U48855 (N_48855,N_36489,N_30673);
xnor U48856 (N_48856,N_32010,N_31434);
and U48857 (N_48857,N_39265,N_37145);
xnor U48858 (N_48858,N_37695,N_31004);
xor U48859 (N_48859,N_37130,N_30987);
nand U48860 (N_48860,N_32395,N_34053);
xnor U48861 (N_48861,N_38195,N_31309);
or U48862 (N_48862,N_36464,N_32728);
nor U48863 (N_48863,N_31314,N_31427);
nand U48864 (N_48864,N_36090,N_30459);
nand U48865 (N_48865,N_33230,N_33273);
or U48866 (N_48866,N_36959,N_35839);
xor U48867 (N_48867,N_35370,N_38780);
nand U48868 (N_48868,N_34602,N_36372);
or U48869 (N_48869,N_37809,N_39172);
or U48870 (N_48870,N_39075,N_31154);
or U48871 (N_48871,N_37892,N_39766);
and U48872 (N_48872,N_38512,N_31987);
and U48873 (N_48873,N_32369,N_30105);
nor U48874 (N_48874,N_35270,N_35740);
xor U48875 (N_48875,N_34238,N_34539);
nor U48876 (N_48876,N_39755,N_35116);
or U48877 (N_48877,N_30373,N_37067);
and U48878 (N_48878,N_33994,N_37885);
and U48879 (N_48879,N_39522,N_35613);
or U48880 (N_48880,N_39675,N_30900);
xnor U48881 (N_48881,N_34210,N_31929);
or U48882 (N_48882,N_33707,N_31865);
and U48883 (N_48883,N_35458,N_34157);
nor U48884 (N_48884,N_35574,N_30813);
xnor U48885 (N_48885,N_34502,N_34237);
and U48886 (N_48886,N_36407,N_32164);
xor U48887 (N_48887,N_37659,N_38912);
or U48888 (N_48888,N_37345,N_35453);
nor U48889 (N_48889,N_35211,N_35041);
nor U48890 (N_48890,N_39013,N_39194);
and U48891 (N_48891,N_39945,N_33989);
nand U48892 (N_48892,N_39580,N_36708);
xor U48893 (N_48893,N_36753,N_38608);
nand U48894 (N_48894,N_33557,N_35730);
and U48895 (N_48895,N_30867,N_34254);
nor U48896 (N_48896,N_33080,N_35206);
and U48897 (N_48897,N_30253,N_36520);
xnor U48898 (N_48898,N_30411,N_32124);
or U48899 (N_48899,N_34058,N_32535);
or U48900 (N_48900,N_34323,N_39846);
or U48901 (N_48901,N_38733,N_34758);
xnor U48902 (N_48902,N_34206,N_37732);
nor U48903 (N_48903,N_37733,N_33545);
nand U48904 (N_48904,N_31345,N_31860);
or U48905 (N_48905,N_31704,N_39856);
xor U48906 (N_48906,N_36167,N_38997);
and U48907 (N_48907,N_31690,N_37560);
xnor U48908 (N_48908,N_38925,N_34981);
nor U48909 (N_48909,N_38180,N_36886);
xor U48910 (N_48910,N_38245,N_37903);
xnor U48911 (N_48911,N_32830,N_36754);
nor U48912 (N_48912,N_39156,N_33100);
xnor U48913 (N_48913,N_34618,N_36144);
nand U48914 (N_48914,N_36100,N_38316);
xor U48915 (N_48915,N_37927,N_38876);
nand U48916 (N_48916,N_31209,N_39432);
nand U48917 (N_48917,N_32331,N_35201);
or U48918 (N_48918,N_31262,N_33727);
xor U48919 (N_48919,N_30946,N_36561);
or U48920 (N_48920,N_31796,N_37305);
and U48921 (N_48921,N_32947,N_30893);
nor U48922 (N_48922,N_31961,N_34824);
nor U48923 (N_48923,N_38863,N_39426);
nor U48924 (N_48924,N_30368,N_36212);
xor U48925 (N_48925,N_33136,N_30595);
and U48926 (N_48926,N_36771,N_38945);
or U48927 (N_48927,N_30957,N_33003);
nand U48928 (N_48928,N_38493,N_36029);
nand U48929 (N_48929,N_34241,N_32214);
xnor U48930 (N_48930,N_30329,N_35567);
xnor U48931 (N_48931,N_34329,N_35818);
xnor U48932 (N_48932,N_34488,N_33855);
nand U48933 (N_48933,N_35312,N_38962);
or U48934 (N_48934,N_32269,N_36015);
and U48935 (N_48935,N_35647,N_30577);
nand U48936 (N_48936,N_36373,N_39188);
and U48937 (N_48937,N_31275,N_32381);
nand U48938 (N_48938,N_35774,N_38882);
xnor U48939 (N_48939,N_37469,N_32828);
and U48940 (N_48940,N_37842,N_36454);
xnor U48941 (N_48941,N_30497,N_30604);
nand U48942 (N_48942,N_31588,N_38869);
nor U48943 (N_48943,N_38096,N_37633);
or U48944 (N_48944,N_32245,N_36921);
and U48945 (N_48945,N_35170,N_36848);
nor U48946 (N_48946,N_35425,N_38158);
xor U48947 (N_48947,N_30558,N_36347);
xnor U48948 (N_48948,N_37816,N_37341);
or U48949 (N_48949,N_35006,N_30144);
nand U48950 (N_48950,N_36140,N_38041);
xor U48951 (N_48951,N_36297,N_34332);
xnor U48952 (N_48952,N_35347,N_37245);
nor U48953 (N_48953,N_33754,N_31499);
xnor U48954 (N_48954,N_35097,N_32552);
nor U48955 (N_48955,N_35590,N_38858);
or U48956 (N_48956,N_31570,N_37769);
xnor U48957 (N_48957,N_36484,N_30387);
nor U48958 (N_48958,N_37257,N_37622);
and U48959 (N_48959,N_36027,N_38017);
xor U48960 (N_48960,N_36455,N_37508);
xor U48961 (N_48961,N_31225,N_39661);
and U48962 (N_48962,N_34174,N_37237);
nor U48963 (N_48963,N_39991,N_34260);
nand U48964 (N_48964,N_31234,N_32152);
and U48965 (N_48965,N_34361,N_31849);
and U48966 (N_48966,N_32465,N_38742);
or U48967 (N_48967,N_39877,N_32888);
nand U48968 (N_48968,N_31359,N_33069);
nor U48969 (N_48969,N_38629,N_31604);
nor U48970 (N_48970,N_34596,N_38386);
or U48971 (N_48971,N_30537,N_30013);
or U48972 (N_48972,N_35431,N_33013);
xor U48973 (N_48973,N_36767,N_31637);
or U48974 (N_48974,N_38534,N_37489);
nand U48975 (N_48975,N_38792,N_39680);
and U48976 (N_48976,N_39491,N_33027);
nor U48977 (N_48977,N_30665,N_36387);
xnor U48978 (N_48978,N_38218,N_30333);
nand U48979 (N_48979,N_34313,N_35709);
xnor U48980 (N_48980,N_34920,N_33958);
and U48981 (N_48981,N_32627,N_34134);
nand U48982 (N_48982,N_33630,N_39905);
xor U48983 (N_48983,N_33663,N_32633);
xor U48984 (N_48984,N_35410,N_33858);
nor U48985 (N_48985,N_36198,N_35001);
and U48986 (N_48986,N_35437,N_39533);
or U48987 (N_48987,N_33003,N_35977);
and U48988 (N_48988,N_36685,N_32250);
nor U48989 (N_48989,N_32544,N_33942);
nand U48990 (N_48990,N_32881,N_31600);
nor U48991 (N_48991,N_34637,N_33296);
nand U48992 (N_48992,N_39851,N_38612);
nor U48993 (N_48993,N_31387,N_34546);
and U48994 (N_48994,N_38830,N_35337);
nor U48995 (N_48995,N_31397,N_30459);
nand U48996 (N_48996,N_33080,N_36864);
nor U48997 (N_48997,N_38869,N_32056);
and U48998 (N_48998,N_37769,N_36951);
nor U48999 (N_48999,N_37435,N_39167);
nor U49000 (N_49000,N_36305,N_34910);
xor U49001 (N_49001,N_38287,N_39359);
and U49002 (N_49002,N_38999,N_39137);
xor U49003 (N_49003,N_38760,N_36252);
or U49004 (N_49004,N_37254,N_37956);
and U49005 (N_49005,N_34625,N_31564);
and U49006 (N_49006,N_32514,N_35987);
nand U49007 (N_49007,N_31663,N_33212);
nor U49008 (N_49008,N_39963,N_36805);
or U49009 (N_49009,N_39172,N_33411);
xnor U49010 (N_49010,N_37863,N_32539);
or U49011 (N_49011,N_31804,N_39249);
nor U49012 (N_49012,N_36639,N_37497);
nand U49013 (N_49013,N_37422,N_37992);
nand U49014 (N_49014,N_32437,N_36951);
and U49015 (N_49015,N_30387,N_30964);
xnor U49016 (N_49016,N_38685,N_32108);
nor U49017 (N_49017,N_33764,N_34417);
nand U49018 (N_49018,N_30925,N_35093);
and U49019 (N_49019,N_38422,N_38349);
xor U49020 (N_49020,N_34135,N_36292);
or U49021 (N_49021,N_38542,N_39016);
nand U49022 (N_49022,N_30263,N_33741);
and U49023 (N_49023,N_34839,N_36532);
and U49024 (N_49024,N_32825,N_34252);
xnor U49025 (N_49025,N_32829,N_30639);
or U49026 (N_49026,N_37639,N_39090);
and U49027 (N_49027,N_31303,N_32403);
xnor U49028 (N_49028,N_32939,N_33172);
or U49029 (N_49029,N_34779,N_33326);
and U49030 (N_49030,N_33109,N_32102);
xor U49031 (N_49031,N_31703,N_33533);
nor U49032 (N_49032,N_39599,N_37038);
xor U49033 (N_49033,N_39937,N_36675);
nor U49034 (N_49034,N_32322,N_32184);
and U49035 (N_49035,N_34760,N_34799);
and U49036 (N_49036,N_37481,N_36310);
or U49037 (N_49037,N_33270,N_30337);
xnor U49038 (N_49038,N_33095,N_30662);
nor U49039 (N_49039,N_31470,N_34682);
nand U49040 (N_49040,N_38170,N_35531);
or U49041 (N_49041,N_30082,N_39545);
and U49042 (N_49042,N_39550,N_38717);
nand U49043 (N_49043,N_32243,N_34279);
nand U49044 (N_49044,N_32500,N_30708);
and U49045 (N_49045,N_38434,N_39824);
or U49046 (N_49046,N_30478,N_38612);
or U49047 (N_49047,N_36263,N_30660);
xor U49048 (N_49048,N_33312,N_37721);
nand U49049 (N_49049,N_31602,N_37197);
nand U49050 (N_49050,N_32039,N_39552);
xnor U49051 (N_49051,N_35607,N_34563);
nand U49052 (N_49052,N_34690,N_31256);
or U49053 (N_49053,N_37903,N_35319);
xor U49054 (N_49054,N_33667,N_39506);
and U49055 (N_49055,N_30182,N_39414);
nor U49056 (N_49056,N_31401,N_32349);
and U49057 (N_49057,N_38544,N_30837);
nor U49058 (N_49058,N_31996,N_31012);
nand U49059 (N_49059,N_34078,N_39129);
or U49060 (N_49060,N_36319,N_31291);
or U49061 (N_49061,N_32542,N_30585);
nand U49062 (N_49062,N_37422,N_38384);
nand U49063 (N_49063,N_32965,N_38468);
nand U49064 (N_49064,N_35192,N_37003);
xnor U49065 (N_49065,N_39301,N_32472);
nand U49066 (N_49066,N_39994,N_31140);
nor U49067 (N_49067,N_32780,N_33010);
xor U49068 (N_49068,N_36198,N_37723);
xor U49069 (N_49069,N_32640,N_38245);
or U49070 (N_49070,N_35409,N_37126);
or U49071 (N_49071,N_39288,N_38628);
and U49072 (N_49072,N_39371,N_31115);
nor U49073 (N_49073,N_39407,N_35990);
and U49074 (N_49074,N_37779,N_30940);
nor U49075 (N_49075,N_31001,N_37399);
or U49076 (N_49076,N_37361,N_30647);
xnor U49077 (N_49077,N_30792,N_37118);
or U49078 (N_49078,N_39298,N_35893);
or U49079 (N_49079,N_36147,N_31740);
nand U49080 (N_49080,N_31017,N_37154);
xor U49081 (N_49081,N_34156,N_32399);
nand U49082 (N_49082,N_37768,N_34049);
and U49083 (N_49083,N_37425,N_33683);
or U49084 (N_49084,N_37520,N_36818);
nand U49085 (N_49085,N_31316,N_39465);
xor U49086 (N_49086,N_39298,N_34596);
or U49087 (N_49087,N_31440,N_35033);
and U49088 (N_49088,N_32733,N_32393);
and U49089 (N_49089,N_35897,N_39604);
nand U49090 (N_49090,N_36190,N_38921);
or U49091 (N_49091,N_36683,N_33206);
nor U49092 (N_49092,N_31509,N_34589);
and U49093 (N_49093,N_39522,N_32158);
nand U49094 (N_49094,N_32309,N_39086);
or U49095 (N_49095,N_34830,N_38858);
nand U49096 (N_49096,N_32251,N_32184);
or U49097 (N_49097,N_32268,N_33455);
nand U49098 (N_49098,N_35835,N_33063);
nor U49099 (N_49099,N_33108,N_39680);
nand U49100 (N_49100,N_30630,N_31639);
nor U49101 (N_49101,N_34184,N_31201);
or U49102 (N_49102,N_30524,N_38218);
and U49103 (N_49103,N_35243,N_33508);
and U49104 (N_49104,N_32875,N_35502);
nor U49105 (N_49105,N_34122,N_31093);
nand U49106 (N_49106,N_36916,N_37788);
and U49107 (N_49107,N_36283,N_30538);
nand U49108 (N_49108,N_30532,N_39934);
or U49109 (N_49109,N_31206,N_37692);
or U49110 (N_49110,N_31570,N_39770);
xor U49111 (N_49111,N_32061,N_33640);
or U49112 (N_49112,N_30813,N_39407);
xnor U49113 (N_49113,N_31923,N_31551);
or U49114 (N_49114,N_30363,N_34759);
or U49115 (N_49115,N_38096,N_32342);
xor U49116 (N_49116,N_36289,N_34726);
xor U49117 (N_49117,N_35824,N_36866);
xor U49118 (N_49118,N_38128,N_34648);
and U49119 (N_49119,N_34729,N_31894);
nor U49120 (N_49120,N_36644,N_33111);
xor U49121 (N_49121,N_37927,N_34146);
xnor U49122 (N_49122,N_35015,N_37756);
or U49123 (N_49123,N_35075,N_34490);
nor U49124 (N_49124,N_35062,N_36329);
nor U49125 (N_49125,N_30711,N_30252);
or U49126 (N_49126,N_36002,N_31768);
or U49127 (N_49127,N_39716,N_31078);
or U49128 (N_49128,N_35887,N_31154);
nand U49129 (N_49129,N_30809,N_30596);
and U49130 (N_49130,N_39359,N_30343);
xnor U49131 (N_49131,N_36466,N_30710);
or U49132 (N_49132,N_33743,N_34876);
or U49133 (N_49133,N_34018,N_38985);
nand U49134 (N_49134,N_31983,N_35358);
nor U49135 (N_49135,N_39163,N_31251);
or U49136 (N_49136,N_39900,N_34400);
or U49137 (N_49137,N_33574,N_39031);
nand U49138 (N_49138,N_38247,N_30511);
nor U49139 (N_49139,N_33731,N_36765);
or U49140 (N_49140,N_33887,N_32309);
or U49141 (N_49141,N_39622,N_38156);
nor U49142 (N_49142,N_36428,N_33571);
xor U49143 (N_49143,N_38472,N_30733);
nand U49144 (N_49144,N_35344,N_35409);
and U49145 (N_49145,N_36404,N_35526);
nand U49146 (N_49146,N_37374,N_38666);
nor U49147 (N_49147,N_38914,N_32102);
xor U49148 (N_49148,N_39061,N_32387);
or U49149 (N_49149,N_38122,N_35199);
xor U49150 (N_49150,N_35278,N_35473);
or U49151 (N_49151,N_33273,N_35120);
nand U49152 (N_49152,N_33856,N_32794);
or U49153 (N_49153,N_35405,N_38863);
nor U49154 (N_49154,N_35928,N_37241);
nand U49155 (N_49155,N_38211,N_39706);
nand U49156 (N_49156,N_36049,N_38078);
or U49157 (N_49157,N_35558,N_39185);
and U49158 (N_49158,N_30395,N_31488);
xor U49159 (N_49159,N_32025,N_38941);
or U49160 (N_49160,N_34651,N_33086);
xor U49161 (N_49161,N_37408,N_33114);
nand U49162 (N_49162,N_35403,N_34251);
nor U49163 (N_49163,N_36461,N_30902);
xor U49164 (N_49164,N_37369,N_36249);
nor U49165 (N_49165,N_31323,N_32175);
and U49166 (N_49166,N_39370,N_39525);
or U49167 (N_49167,N_35189,N_38210);
and U49168 (N_49168,N_39936,N_37797);
nand U49169 (N_49169,N_34431,N_34740);
nand U49170 (N_49170,N_34972,N_37719);
nor U49171 (N_49171,N_38605,N_30010);
nor U49172 (N_49172,N_36682,N_34553);
xor U49173 (N_49173,N_34225,N_37295);
nor U49174 (N_49174,N_33098,N_30709);
nand U49175 (N_49175,N_35637,N_37471);
nor U49176 (N_49176,N_31184,N_34111);
or U49177 (N_49177,N_31739,N_32757);
and U49178 (N_49178,N_39458,N_31990);
nand U49179 (N_49179,N_34808,N_36463);
nor U49180 (N_49180,N_33747,N_33078);
nand U49181 (N_49181,N_37891,N_31215);
or U49182 (N_49182,N_36132,N_31105);
or U49183 (N_49183,N_39077,N_39832);
and U49184 (N_49184,N_30922,N_38179);
xnor U49185 (N_49185,N_35648,N_38283);
xor U49186 (N_49186,N_36748,N_39079);
xor U49187 (N_49187,N_34461,N_31823);
nor U49188 (N_49188,N_38166,N_37508);
nand U49189 (N_49189,N_30546,N_36246);
xor U49190 (N_49190,N_39627,N_38476);
nor U49191 (N_49191,N_31124,N_31855);
or U49192 (N_49192,N_31795,N_33209);
nand U49193 (N_49193,N_31591,N_30963);
nand U49194 (N_49194,N_34347,N_39820);
or U49195 (N_49195,N_30851,N_38162);
nor U49196 (N_49196,N_32450,N_39495);
or U49197 (N_49197,N_32008,N_32883);
nor U49198 (N_49198,N_32362,N_39573);
xor U49199 (N_49199,N_34429,N_31495);
nand U49200 (N_49200,N_37215,N_33228);
nand U49201 (N_49201,N_35295,N_33070);
or U49202 (N_49202,N_39009,N_39109);
nor U49203 (N_49203,N_35120,N_35106);
xor U49204 (N_49204,N_35809,N_37581);
nand U49205 (N_49205,N_34201,N_31402);
xnor U49206 (N_49206,N_32131,N_36974);
and U49207 (N_49207,N_32382,N_32309);
and U49208 (N_49208,N_35899,N_37325);
xnor U49209 (N_49209,N_32490,N_37751);
and U49210 (N_49210,N_34244,N_39937);
or U49211 (N_49211,N_37470,N_38624);
or U49212 (N_49212,N_38784,N_33456);
nand U49213 (N_49213,N_37466,N_35091);
nor U49214 (N_49214,N_37205,N_36476);
and U49215 (N_49215,N_34482,N_35294);
nor U49216 (N_49216,N_30686,N_38263);
and U49217 (N_49217,N_34455,N_37342);
nand U49218 (N_49218,N_34394,N_33297);
xnor U49219 (N_49219,N_38353,N_32823);
nor U49220 (N_49220,N_32916,N_33915);
xnor U49221 (N_49221,N_32205,N_31706);
xor U49222 (N_49222,N_39348,N_35661);
or U49223 (N_49223,N_35818,N_37490);
or U49224 (N_49224,N_38501,N_33132);
xnor U49225 (N_49225,N_35980,N_33076);
nor U49226 (N_49226,N_33128,N_38210);
nor U49227 (N_49227,N_32075,N_38534);
nand U49228 (N_49228,N_30532,N_30618);
xor U49229 (N_49229,N_32346,N_36875);
nor U49230 (N_49230,N_36925,N_34878);
nand U49231 (N_49231,N_31102,N_37075);
xor U49232 (N_49232,N_35611,N_39372);
nor U49233 (N_49233,N_34124,N_30193);
nand U49234 (N_49234,N_38509,N_39327);
or U49235 (N_49235,N_35806,N_31868);
or U49236 (N_49236,N_30774,N_33505);
xnor U49237 (N_49237,N_33964,N_33867);
nand U49238 (N_49238,N_31080,N_31763);
nand U49239 (N_49239,N_31379,N_34913);
nor U49240 (N_49240,N_37006,N_38836);
nand U49241 (N_49241,N_32438,N_38754);
and U49242 (N_49242,N_36007,N_34270);
xnor U49243 (N_49243,N_39728,N_37753);
nand U49244 (N_49244,N_31558,N_38709);
nand U49245 (N_49245,N_38644,N_30047);
nand U49246 (N_49246,N_37362,N_36491);
nand U49247 (N_49247,N_39414,N_39078);
nand U49248 (N_49248,N_34081,N_37732);
and U49249 (N_49249,N_37566,N_37259);
xnor U49250 (N_49250,N_32867,N_37264);
xor U49251 (N_49251,N_34656,N_37764);
nor U49252 (N_49252,N_32277,N_33614);
or U49253 (N_49253,N_38330,N_34403);
and U49254 (N_49254,N_38858,N_35371);
nand U49255 (N_49255,N_36008,N_33598);
and U49256 (N_49256,N_33588,N_36066);
or U49257 (N_49257,N_33313,N_36276);
nand U49258 (N_49258,N_33321,N_38391);
nor U49259 (N_49259,N_31941,N_32399);
nand U49260 (N_49260,N_39013,N_39714);
or U49261 (N_49261,N_32471,N_34602);
and U49262 (N_49262,N_38733,N_33309);
xor U49263 (N_49263,N_31815,N_38751);
and U49264 (N_49264,N_33826,N_36222);
xor U49265 (N_49265,N_33277,N_30548);
and U49266 (N_49266,N_33136,N_38033);
nor U49267 (N_49267,N_36690,N_33000);
nand U49268 (N_49268,N_37599,N_35899);
xor U49269 (N_49269,N_30559,N_35731);
xnor U49270 (N_49270,N_30508,N_32596);
and U49271 (N_49271,N_32571,N_37565);
and U49272 (N_49272,N_32748,N_32658);
xor U49273 (N_49273,N_33958,N_36494);
and U49274 (N_49274,N_32541,N_33317);
and U49275 (N_49275,N_36927,N_35128);
nand U49276 (N_49276,N_38647,N_30036);
or U49277 (N_49277,N_35714,N_38569);
and U49278 (N_49278,N_30671,N_30886);
and U49279 (N_49279,N_31465,N_37060);
nand U49280 (N_49280,N_33654,N_30732);
nand U49281 (N_49281,N_34302,N_31307);
or U49282 (N_49282,N_34742,N_37262);
nand U49283 (N_49283,N_31891,N_38590);
nand U49284 (N_49284,N_37754,N_31766);
nor U49285 (N_49285,N_38324,N_30172);
nor U49286 (N_49286,N_35389,N_35212);
xnor U49287 (N_49287,N_31382,N_34598);
or U49288 (N_49288,N_35729,N_32113);
and U49289 (N_49289,N_37835,N_35941);
xnor U49290 (N_49290,N_38856,N_39159);
nor U49291 (N_49291,N_32414,N_38086);
or U49292 (N_49292,N_37641,N_34868);
xnor U49293 (N_49293,N_39978,N_37895);
nand U49294 (N_49294,N_31030,N_32960);
nand U49295 (N_49295,N_35507,N_35272);
or U49296 (N_49296,N_32952,N_32183);
and U49297 (N_49297,N_39469,N_30277);
nor U49298 (N_49298,N_30178,N_32877);
and U49299 (N_49299,N_36027,N_34700);
and U49300 (N_49300,N_38879,N_32881);
and U49301 (N_49301,N_37494,N_30024);
xnor U49302 (N_49302,N_30636,N_31574);
or U49303 (N_49303,N_31288,N_32135);
or U49304 (N_49304,N_36061,N_33356);
nand U49305 (N_49305,N_36357,N_31740);
or U49306 (N_49306,N_32991,N_35455);
or U49307 (N_49307,N_38551,N_31578);
and U49308 (N_49308,N_31752,N_39928);
nor U49309 (N_49309,N_35063,N_39053);
and U49310 (N_49310,N_36310,N_37364);
xnor U49311 (N_49311,N_31348,N_32866);
nand U49312 (N_49312,N_36496,N_30492);
nand U49313 (N_49313,N_37015,N_33121);
and U49314 (N_49314,N_32188,N_31524);
xor U49315 (N_49315,N_37955,N_35198);
nor U49316 (N_49316,N_33259,N_32830);
or U49317 (N_49317,N_37440,N_33871);
xnor U49318 (N_49318,N_39713,N_32942);
nor U49319 (N_49319,N_31570,N_36677);
or U49320 (N_49320,N_36247,N_30011);
and U49321 (N_49321,N_35614,N_35920);
xnor U49322 (N_49322,N_39379,N_35759);
nor U49323 (N_49323,N_33878,N_36300);
and U49324 (N_49324,N_38341,N_36273);
and U49325 (N_49325,N_37960,N_39062);
xnor U49326 (N_49326,N_37833,N_38792);
or U49327 (N_49327,N_34879,N_36456);
xnor U49328 (N_49328,N_37074,N_38679);
nand U49329 (N_49329,N_31352,N_31428);
xnor U49330 (N_49330,N_37183,N_31471);
nand U49331 (N_49331,N_32840,N_35874);
or U49332 (N_49332,N_31440,N_30465);
or U49333 (N_49333,N_36717,N_34780);
or U49334 (N_49334,N_30907,N_30067);
xor U49335 (N_49335,N_38696,N_33835);
and U49336 (N_49336,N_33021,N_33526);
or U49337 (N_49337,N_37496,N_31699);
nand U49338 (N_49338,N_34075,N_30478);
nor U49339 (N_49339,N_39753,N_38909);
nor U49340 (N_49340,N_31623,N_35195);
nand U49341 (N_49341,N_37992,N_33327);
or U49342 (N_49342,N_36163,N_30833);
xor U49343 (N_49343,N_39153,N_35139);
and U49344 (N_49344,N_37555,N_38764);
or U49345 (N_49345,N_31882,N_35614);
nand U49346 (N_49346,N_37689,N_37246);
nor U49347 (N_49347,N_33676,N_31060);
and U49348 (N_49348,N_35122,N_34822);
nor U49349 (N_49349,N_37259,N_35759);
nand U49350 (N_49350,N_38921,N_35989);
nand U49351 (N_49351,N_33648,N_31995);
xor U49352 (N_49352,N_39732,N_35490);
nand U49353 (N_49353,N_36102,N_38316);
or U49354 (N_49354,N_35642,N_36667);
and U49355 (N_49355,N_33135,N_34356);
and U49356 (N_49356,N_38046,N_32688);
and U49357 (N_49357,N_31028,N_34619);
nand U49358 (N_49358,N_30588,N_31864);
or U49359 (N_49359,N_38313,N_35874);
nand U49360 (N_49360,N_31658,N_36569);
nor U49361 (N_49361,N_38371,N_33096);
and U49362 (N_49362,N_37139,N_39962);
nor U49363 (N_49363,N_32649,N_34290);
nor U49364 (N_49364,N_32709,N_34128);
nand U49365 (N_49365,N_36993,N_35282);
and U49366 (N_49366,N_37681,N_30122);
nor U49367 (N_49367,N_35142,N_35775);
nor U49368 (N_49368,N_35610,N_35389);
xor U49369 (N_49369,N_32179,N_33531);
or U49370 (N_49370,N_39313,N_35035);
and U49371 (N_49371,N_38363,N_38737);
or U49372 (N_49372,N_33359,N_37050);
and U49373 (N_49373,N_32503,N_35399);
nand U49374 (N_49374,N_37729,N_35937);
nand U49375 (N_49375,N_34338,N_33149);
nor U49376 (N_49376,N_32376,N_39661);
nor U49377 (N_49377,N_38320,N_34848);
xnor U49378 (N_49378,N_38088,N_36304);
xor U49379 (N_49379,N_32781,N_37303);
xnor U49380 (N_49380,N_38361,N_33100);
nor U49381 (N_49381,N_34079,N_38234);
xnor U49382 (N_49382,N_36193,N_38825);
or U49383 (N_49383,N_30567,N_32865);
and U49384 (N_49384,N_39021,N_34129);
or U49385 (N_49385,N_39902,N_34367);
xnor U49386 (N_49386,N_36458,N_30829);
or U49387 (N_49387,N_30953,N_33536);
xnor U49388 (N_49388,N_33989,N_33793);
and U49389 (N_49389,N_30997,N_31053);
xnor U49390 (N_49390,N_38425,N_36411);
and U49391 (N_49391,N_39462,N_30200);
nor U49392 (N_49392,N_35525,N_33503);
xor U49393 (N_49393,N_39642,N_36148);
nor U49394 (N_49394,N_31015,N_33170);
nand U49395 (N_49395,N_31123,N_37882);
or U49396 (N_49396,N_32239,N_38599);
xor U49397 (N_49397,N_35753,N_30111);
and U49398 (N_49398,N_33101,N_35544);
nor U49399 (N_49399,N_35118,N_30187);
and U49400 (N_49400,N_34642,N_35511);
or U49401 (N_49401,N_35298,N_31103);
nor U49402 (N_49402,N_37435,N_37180);
nor U49403 (N_49403,N_30603,N_35856);
nand U49404 (N_49404,N_30241,N_35114);
xnor U49405 (N_49405,N_38413,N_31183);
nand U49406 (N_49406,N_32960,N_35690);
nand U49407 (N_49407,N_33485,N_38750);
nor U49408 (N_49408,N_38032,N_31598);
nand U49409 (N_49409,N_35164,N_30888);
xor U49410 (N_49410,N_35015,N_31843);
nand U49411 (N_49411,N_32519,N_35032);
nor U49412 (N_49412,N_32997,N_39429);
and U49413 (N_49413,N_36781,N_35972);
and U49414 (N_49414,N_37389,N_34837);
nand U49415 (N_49415,N_34581,N_33298);
nor U49416 (N_49416,N_34356,N_39716);
nand U49417 (N_49417,N_35478,N_36229);
xor U49418 (N_49418,N_36707,N_39714);
nand U49419 (N_49419,N_30421,N_32928);
xor U49420 (N_49420,N_32701,N_38009);
nand U49421 (N_49421,N_35475,N_31991);
nor U49422 (N_49422,N_31205,N_33280);
and U49423 (N_49423,N_36943,N_30307);
xnor U49424 (N_49424,N_35434,N_39092);
xnor U49425 (N_49425,N_35747,N_33513);
xnor U49426 (N_49426,N_39543,N_32768);
or U49427 (N_49427,N_33718,N_35334);
and U49428 (N_49428,N_30034,N_32228);
nor U49429 (N_49429,N_38669,N_38470);
nor U49430 (N_49430,N_39887,N_31445);
and U49431 (N_49431,N_34518,N_37754);
nand U49432 (N_49432,N_35316,N_34439);
or U49433 (N_49433,N_39540,N_33802);
and U49434 (N_49434,N_30594,N_33146);
nor U49435 (N_49435,N_34820,N_38217);
xnor U49436 (N_49436,N_31542,N_38093);
xor U49437 (N_49437,N_33126,N_35360);
xor U49438 (N_49438,N_31751,N_38169);
xor U49439 (N_49439,N_36861,N_33900);
nor U49440 (N_49440,N_31512,N_35116);
xnor U49441 (N_49441,N_30659,N_31576);
or U49442 (N_49442,N_32148,N_31191);
nor U49443 (N_49443,N_35051,N_34353);
xor U49444 (N_49444,N_39637,N_30111);
nor U49445 (N_49445,N_31125,N_36334);
or U49446 (N_49446,N_34097,N_39766);
or U49447 (N_49447,N_36989,N_36993);
or U49448 (N_49448,N_39876,N_33692);
nand U49449 (N_49449,N_34355,N_31315);
nand U49450 (N_49450,N_30692,N_38712);
xor U49451 (N_49451,N_34414,N_37694);
nor U49452 (N_49452,N_37070,N_30129);
and U49453 (N_49453,N_32107,N_35933);
and U49454 (N_49454,N_34879,N_39533);
nand U49455 (N_49455,N_37674,N_31439);
and U49456 (N_49456,N_31970,N_39026);
or U49457 (N_49457,N_30843,N_34722);
and U49458 (N_49458,N_32326,N_39369);
nand U49459 (N_49459,N_30312,N_32410);
and U49460 (N_49460,N_39669,N_37455);
nor U49461 (N_49461,N_35578,N_31150);
nor U49462 (N_49462,N_38366,N_39670);
nand U49463 (N_49463,N_37921,N_33193);
nand U49464 (N_49464,N_39290,N_34007);
xor U49465 (N_49465,N_31711,N_35351);
nor U49466 (N_49466,N_38262,N_36466);
or U49467 (N_49467,N_30141,N_32988);
nand U49468 (N_49468,N_34886,N_31834);
xnor U49469 (N_49469,N_37894,N_30060);
xnor U49470 (N_49470,N_34871,N_38482);
or U49471 (N_49471,N_35018,N_38920);
nor U49472 (N_49472,N_34155,N_36874);
xnor U49473 (N_49473,N_36397,N_34315);
nand U49474 (N_49474,N_38995,N_35194);
xor U49475 (N_49475,N_31572,N_34603);
xnor U49476 (N_49476,N_34902,N_31019);
and U49477 (N_49477,N_38492,N_33465);
xnor U49478 (N_49478,N_38588,N_34719);
or U49479 (N_49479,N_35862,N_36362);
nand U49480 (N_49480,N_39188,N_39996);
nand U49481 (N_49481,N_38852,N_38906);
nand U49482 (N_49482,N_30885,N_34311);
and U49483 (N_49483,N_36870,N_33762);
nand U49484 (N_49484,N_36236,N_30048);
nor U49485 (N_49485,N_31242,N_30865);
xnor U49486 (N_49486,N_36832,N_30238);
nor U49487 (N_49487,N_35611,N_34661);
or U49488 (N_49488,N_31309,N_30390);
or U49489 (N_49489,N_30379,N_34336);
and U49490 (N_49490,N_32052,N_37347);
nand U49491 (N_49491,N_32747,N_32275);
nor U49492 (N_49492,N_36162,N_30318);
nor U49493 (N_49493,N_34792,N_35581);
nand U49494 (N_49494,N_37813,N_30685);
and U49495 (N_49495,N_39092,N_36701);
nand U49496 (N_49496,N_32625,N_31109);
nand U49497 (N_49497,N_39100,N_32421);
nor U49498 (N_49498,N_31563,N_38076);
nand U49499 (N_49499,N_39173,N_36245);
or U49500 (N_49500,N_38347,N_32722);
nor U49501 (N_49501,N_30110,N_31084);
or U49502 (N_49502,N_31012,N_35095);
or U49503 (N_49503,N_35276,N_39968);
and U49504 (N_49504,N_31668,N_39193);
xnor U49505 (N_49505,N_36806,N_33958);
nor U49506 (N_49506,N_36323,N_30706);
nor U49507 (N_49507,N_30529,N_37462);
and U49508 (N_49508,N_30942,N_33820);
or U49509 (N_49509,N_30165,N_39092);
nand U49510 (N_49510,N_38695,N_38039);
nor U49511 (N_49511,N_32953,N_38273);
or U49512 (N_49512,N_34299,N_31544);
xnor U49513 (N_49513,N_39396,N_32624);
nand U49514 (N_49514,N_35942,N_35604);
nor U49515 (N_49515,N_37293,N_30158);
or U49516 (N_49516,N_37374,N_36037);
xnor U49517 (N_49517,N_30842,N_33537);
and U49518 (N_49518,N_31279,N_31032);
nor U49519 (N_49519,N_37622,N_38531);
and U49520 (N_49520,N_34553,N_32108);
xnor U49521 (N_49521,N_37695,N_30209);
xor U49522 (N_49522,N_36382,N_38798);
nor U49523 (N_49523,N_35089,N_39264);
or U49524 (N_49524,N_36234,N_37806);
nor U49525 (N_49525,N_34921,N_35944);
or U49526 (N_49526,N_36946,N_35963);
or U49527 (N_49527,N_34780,N_39963);
and U49528 (N_49528,N_38025,N_31148);
or U49529 (N_49529,N_38073,N_30044);
xor U49530 (N_49530,N_37918,N_31770);
and U49531 (N_49531,N_32721,N_36575);
xnor U49532 (N_49532,N_32945,N_36950);
xnor U49533 (N_49533,N_34423,N_39747);
nand U49534 (N_49534,N_33167,N_33885);
and U49535 (N_49535,N_31751,N_34311);
nand U49536 (N_49536,N_34245,N_33044);
nor U49537 (N_49537,N_37114,N_37938);
nor U49538 (N_49538,N_36241,N_34490);
xor U49539 (N_49539,N_39682,N_33488);
and U49540 (N_49540,N_30450,N_37161);
nand U49541 (N_49541,N_36493,N_39405);
or U49542 (N_49542,N_33563,N_38094);
and U49543 (N_49543,N_35920,N_39627);
and U49544 (N_49544,N_36101,N_33281);
or U49545 (N_49545,N_39187,N_38200);
and U49546 (N_49546,N_34985,N_36787);
or U49547 (N_49547,N_39562,N_37544);
and U49548 (N_49548,N_31058,N_33770);
and U49549 (N_49549,N_32318,N_38730);
nand U49550 (N_49550,N_30105,N_35936);
nor U49551 (N_49551,N_38453,N_33899);
and U49552 (N_49552,N_33163,N_35079);
xor U49553 (N_49553,N_37996,N_31547);
xnor U49554 (N_49554,N_38020,N_38832);
xnor U49555 (N_49555,N_38283,N_39234);
or U49556 (N_49556,N_37766,N_35972);
nand U49557 (N_49557,N_33576,N_39596);
xor U49558 (N_49558,N_33135,N_32259);
nor U49559 (N_49559,N_31277,N_31524);
and U49560 (N_49560,N_38274,N_33824);
xnor U49561 (N_49561,N_33589,N_35540);
and U49562 (N_49562,N_39202,N_34709);
nor U49563 (N_49563,N_31590,N_37794);
nor U49564 (N_49564,N_30343,N_39739);
nand U49565 (N_49565,N_35646,N_30539);
nand U49566 (N_49566,N_37688,N_33835);
nand U49567 (N_49567,N_30874,N_32791);
or U49568 (N_49568,N_32454,N_30572);
nand U49569 (N_49569,N_38985,N_38681);
nand U49570 (N_49570,N_37553,N_31136);
xor U49571 (N_49571,N_34624,N_37086);
and U49572 (N_49572,N_39670,N_30675);
nand U49573 (N_49573,N_31341,N_30812);
or U49574 (N_49574,N_33970,N_38199);
nand U49575 (N_49575,N_39263,N_30779);
nor U49576 (N_49576,N_37593,N_35421);
and U49577 (N_49577,N_37857,N_36362);
or U49578 (N_49578,N_37297,N_34128);
nand U49579 (N_49579,N_37802,N_30874);
nand U49580 (N_49580,N_33020,N_38188);
or U49581 (N_49581,N_36259,N_31338);
or U49582 (N_49582,N_35363,N_38385);
xnor U49583 (N_49583,N_36648,N_37410);
and U49584 (N_49584,N_36143,N_33745);
nand U49585 (N_49585,N_33671,N_35293);
nor U49586 (N_49586,N_39028,N_38452);
xor U49587 (N_49587,N_38839,N_36059);
nor U49588 (N_49588,N_34790,N_37409);
or U49589 (N_49589,N_32197,N_30023);
nand U49590 (N_49590,N_34562,N_37046);
and U49591 (N_49591,N_33731,N_30089);
or U49592 (N_49592,N_36525,N_32612);
xnor U49593 (N_49593,N_32139,N_34977);
nand U49594 (N_49594,N_33184,N_34681);
nand U49595 (N_49595,N_30653,N_38771);
nor U49596 (N_49596,N_32512,N_39091);
xor U49597 (N_49597,N_30845,N_38246);
nand U49598 (N_49598,N_34836,N_36467);
or U49599 (N_49599,N_30135,N_33196);
and U49600 (N_49600,N_34822,N_38091);
nor U49601 (N_49601,N_32370,N_39056);
and U49602 (N_49602,N_30837,N_33225);
and U49603 (N_49603,N_32166,N_30883);
nand U49604 (N_49604,N_34921,N_34939);
nor U49605 (N_49605,N_37467,N_35624);
xor U49606 (N_49606,N_38865,N_34915);
or U49607 (N_49607,N_34733,N_33487);
or U49608 (N_49608,N_39869,N_38243);
nand U49609 (N_49609,N_39785,N_30591);
or U49610 (N_49610,N_34062,N_32505);
nand U49611 (N_49611,N_35480,N_30541);
and U49612 (N_49612,N_35056,N_35920);
xnor U49613 (N_49613,N_39156,N_35878);
nand U49614 (N_49614,N_30757,N_33858);
nor U49615 (N_49615,N_37016,N_32217);
and U49616 (N_49616,N_36749,N_36515);
nor U49617 (N_49617,N_31767,N_34920);
nor U49618 (N_49618,N_33205,N_39823);
xnor U49619 (N_49619,N_37687,N_37786);
or U49620 (N_49620,N_31747,N_32082);
and U49621 (N_49621,N_31281,N_34375);
nand U49622 (N_49622,N_39617,N_39695);
nand U49623 (N_49623,N_37228,N_33959);
and U49624 (N_49624,N_34608,N_39573);
or U49625 (N_49625,N_39320,N_34346);
and U49626 (N_49626,N_30800,N_39280);
xor U49627 (N_49627,N_36520,N_33654);
or U49628 (N_49628,N_30025,N_33866);
nand U49629 (N_49629,N_30716,N_38837);
or U49630 (N_49630,N_31086,N_37258);
xor U49631 (N_49631,N_30295,N_35091);
nand U49632 (N_49632,N_35514,N_38508);
nand U49633 (N_49633,N_34825,N_33284);
and U49634 (N_49634,N_32314,N_34742);
xnor U49635 (N_49635,N_32085,N_37904);
nand U49636 (N_49636,N_34269,N_32425);
nor U49637 (N_49637,N_31890,N_31174);
nor U49638 (N_49638,N_33243,N_36457);
xor U49639 (N_49639,N_38032,N_35517);
nor U49640 (N_49640,N_31473,N_39270);
and U49641 (N_49641,N_34355,N_33590);
nor U49642 (N_49642,N_30515,N_33825);
nor U49643 (N_49643,N_31098,N_32965);
xor U49644 (N_49644,N_35650,N_36556);
nor U49645 (N_49645,N_30390,N_31822);
nand U49646 (N_49646,N_35409,N_32198);
xnor U49647 (N_49647,N_39697,N_33368);
nor U49648 (N_49648,N_35627,N_35538);
nand U49649 (N_49649,N_34820,N_37357);
nor U49650 (N_49650,N_32196,N_36627);
xnor U49651 (N_49651,N_32650,N_36308);
nor U49652 (N_49652,N_30939,N_38015);
nor U49653 (N_49653,N_38982,N_31462);
nand U49654 (N_49654,N_38957,N_39700);
xor U49655 (N_49655,N_38544,N_37263);
or U49656 (N_49656,N_36178,N_32273);
and U49657 (N_49657,N_38217,N_38498);
and U49658 (N_49658,N_36979,N_37951);
nand U49659 (N_49659,N_36771,N_35228);
nor U49660 (N_49660,N_38264,N_34190);
and U49661 (N_49661,N_32056,N_37630);
and U49662 (N_49662,N_39270,N_36151);
and U49663 (N_49663,N_31657,N_30186);
nor U49664 (N_49664,N_36860,N_38787);
and U49665 (N_49665,N_38754,N_36835);
xnor U49666 (N_49666,N_38029,N_38766);
xnor U49667 (N_49667,N_38140,N_39571);
and U49668 (N_49668,N_39958,N_35502);
xor U49669 (N_49669,N_37661,N_39921);
or U49670 (N_49670,N_38075,N_30821);
nand U49671 (N_49671,N_32468,N_37722);
nand U49672 (N_49672,N_38879,N_38153);
xor U49673 (N_49673,N_38607,N_38389);
or U49674 (N_49674,N_39297,N_34263);
and U49675 (N_49675,N_32300,N_35240);
nand U49676 (N_49676,N_38157,N_32432);
nand U49677 (N_49677,N_37358,N_36032);
nand U49678 (N_49678,N_30374,N_36736);
or U49679 (N_49679,N_34917,N_36163);
nor U49680 (N_49680,N_39371,N_38426);
and U49681 (N_49681,N_32921,N_39228);
nor U49682 (N_49682,N_35396,N_31727);
or U49683 (N_49683,N_35332,N_33706);
or U49684 (N_49684,N_33672,N_38185);
and U49685 (N_49685,N_36048,N_38502);
xnor U49686 (N_49686,N_30002,N_36635);
nand U49687 (N_49687,N_32494,N_38387);
or U49688 (N_49688,N_36390,N_33737);
nor U49689 (N_49689,N_31859,N_34833);
nand U49690 (N_49690,N_32617,N_36403);
nand U49691 (N_49691,N_36660,N_31105);
nor U49692 (N_49692,N_35737,N_37987);
nand U49693 (N_49693,N_32898,N_31122);
nor U49694 (N_49694,N_31924,N_32171);
xnor U49695 (N_49695,N_36230,N_30136);
or U49696 (N_49696,N_32350,N_37209);
and U49697 (N_49697,N_30002,N_34444);
xor U49698 (N_49698,N_38331,N_37803);
and U49699 (N_49699,N_38523,N_35421);
or U49700 (N_49700,N_36229,N_30918);
or U49701 (N_49701,N_31054,N_37083);
nand U49702 (N_49702,N_37298,N_33547);
and U49703 (N_49703,N_35479,N_38156);
nor U49704 (N_49704,N_39227,N_34474);
nor U49705 (N_49705,N_35915,N_35056);
nand U49706 (N_49706,N_35293,N_33071);
nand U49707 (N_49707,N_32325,N_39003);
xnor U49708 (N_49708,N_38564,N_35392);
or U49709 (N_49709,N_33034,N_39224);
and U49710 (N_49710,N_37211,N_33820);
or U49711 (N_49711,N_36394,N_37660);
and U49712 (N_49712,N_31154,N_33034);
and U49713 (N_49713,N_38342,N_39215);
or U49714 (N_49714,N_34743,N_32694);
xnor U49715 (N_49715,N_35818,N_36123);
xnor U49716 (N_49716,N_39186,N_35391);
and U49717 (N_49717,N_37957,N_35046);
nor U49718 (N_49718,N_39138,N_39972);
nor U49719 (N_49719,N_33584,N_35663);
or U49720 (N_49720,N_30881,N_33210);
nand U49721 (N_49721,N_39166,N_36484);
nand U49722 (N_49722,N_32626,N_30431);
xnor U49723 (N_49723,N_37846,N_34801);
xor U49724 (N_49724,N_31967,N_36005);
or U49725 (N_49725,N_33947,N_35851);
or U49726 (N_49726,N_33330,N_37111);
nor U49727 (N_49727,N_31237,N_33773);
nor U49728 (N_49728,N_37722,N_36933);
nor U49729 (N_49729,N_32030,N_37798);
and U49730 (N_49730,N_32517,N_36996);
nand U49731 (N_49731,N_38394,N_31233);
or U49732 (N_49732,N_32234,N_31029);
and U49733 (N_49733,N_35569,N_30778);
nand U49734 (N_49734,N_30047,N_36568);
or U49735 (N_49735,N_39096,N_35361);
nor U49736 (N_49736,N_36444,N_37664);
nor U49737 (N_49737,N_39806,N_37221);
nor U49738 (N_49738,N_36730,N_34759);
xnor U49739 (N_49739,N_36705,N_37989);
xnor U49740 (N_49740,N_33057,N_30309);
nand U49741 (N_49741,N_38571,N_35939);
and U49742 (N_49742,N_30104,N_36004);
nand U49743 (N_49743,N_36520,N_31506);
nor U49744 (N_49744,N_35931,N_38709);
nand U49745 (N_49745,N_32177,N_33177);
and U49746 (N_49746,N_38543,N_30456);
nand U49747 (N_49747,N_39568,N_33150);
and U49748 (N_49748,N_32223,N_36654);
nand U49749 (N_49749,N_30748,N_30309);
nor U49750 (N_49750,N_31838,N_38826);
xor U49751 (N_49751,N_32116,N_39030);
nor U49752 (N_49752,N_31494,N_31496);
nor U49753 (N_49753,N_37698,N_33030);
and U49754 (N_49754,N_38263,N_34286);
xor U49755 (N_49755,N_35728,N_38417);
xor U49756 (N_49756,N_37417,N_37948);
nor U49757 (N_49757,N_37395,N_39426);
and U49758 (N_49758,N_33424,N_34988);
or U49759 (N_49759,N_32238,N_38054);
xnor U49760 (N_49760,N_33541,N_35778);
nor U49761 (N_49761,N_34601,N_39074);
and U49762 (N_49762,N_31479,N_33564);
xor U49763 (N_49763,N_39856,N_36985);
xor U49764 (N_49764,N_38832,N_33389);
and U49765 (N_49765,N_38391,N_33578);
and U49766 (N_49766,N_32654,N_35047);
or U49767 (N_49767,N_34125,N_31004);
and U49768 (N_49768,N_31193,N_30506);
xor U49769 (N_49769,N_34416,N_36696);
and U49770 (N_49770,N_36173,N_39918);
nor U49771 (N_49771,N_31389,N_33792);
nand U49772 (N_49772,N_34666,N_30128);
nand U49773 (N_49773,N_35977,N_32159);
xor U49774 (N_49774,N_39945,N_34033);
nor U49775 (N_49775,N_38954,N_38158);
and U49776 (N_49776,N_39255,N_31772);
or U49777 (N_49777,N_37274,N_39475);
nand U49778 (N_49778,N_34885,N_34865);
nor U49779 (N_49779,N_35239,N_34379);
or U49780 (N_49780,N_36277,N_36814);
xor U49781 (N_49781,N_31323,N_32061);
nor U49782 (N_49782,N_37647,N_37372);
xnor U49783 (N_49783,N_35033,N_36487);
xnor U49784 (N_49784,N_39417,N_35474);
and U49785 (N_49785,N_34517,N_30758);
or U49786 (N_49786,N_39623,N_39965);
or U49787 (N_49787,N_36027,N_37709);
and U49788 (N_49788,N_30765,N_39646);
xnor U49789 (N_49789,N_39494,N_35173);
nand U49790 (N_49790,N_36189,N_38287);
nand U49791 (N_49791,N_32416,N_36602);
nor U49792 (N_49792,N_38149,N_38843);
xor U49793 (N_49793,N_31086,N_38438);
or U49794 (N_49794,N_31413,N_36873);
or U49795 (N_49795,N_33258,N_37414);
nor U49796 (N_49796,N_35693,N_34688);
nand U49797 (N_49797,N_31933,N_39390);
nand U49798 (N_49798,N_32259,N_30447);
and U49799 (N_49799,N_33494,N_34196);
nor U49800 (N_49800,N_33699,N_33445);
nand U49801 (N_49801,N_39590,N_34071);
nor U49802 (N_49802,N_39158,N_31191);
or U49803 (N_49803,N_35784,N_35888);
nand U49804 (N_49804,N_34403,N_39042);
and U49805 (N_49805,N_34933,N_36777);
nor U49806 (N_49806,N_32274,N_38777);
or U49807 (N_49807,N_35616,N_30598);
nor U49808 (N_49808,N_35808,N_33280);
or U49809 (N_49809,N_36441,N_38193);
nand U49810 (N_49810,N_39466,N_32904);
xor U49811 (N_49811,N_34029,N_33751);
nand U49812 (N_49812,N_36363,N_32575);
nand U49813 (N_49813,N_30829,N_37096);
and U49814 (N_49814,N_35875,N_37406);
nand U49815 (N_49815,N_36485,N_34558);
nand U49816 (N_49816,N_35896,N_36688);
or U49817 (N_49817,N_35124,N_37688);
nand U49818 (N_49818,N_39660,N_38479);
nand U49819 (N_49819,N_38280,N_34837);
xnor U49820 (N_49820,N_35149,N_36012);
and U49821 (N_49821,N_37885,N_30494);
or U49822 (N_49822,N_31793,N_31343);
nor U49823 (N_49823,N_37467,N_39546);
nor U49824 (N_49824,N_33393,N_37551);
or U49825 (N_49825,N_30367,N_39982);
or U49826 (N_49826,N_34511,N_36829);
nand U49827 (N_49827,N_35378,N_37713);
and U49828 (N_49828,N_33703,N_38896);
nand U49829 (N_49829,N_38556,N_31150);
xnor U49830 (N_49830,N_31763,N_31860);
nand U49831 (N_49831,N_34938,N_31484);
and U49832 (N_49832,N_39601,N_33221);
nand U49833 (N_49833,N_37834,N_39487);
xnor U49834 (N_49834,N_37279,N_35296);
or U49835 (N_49835,N_38901,N_32166);
or U49836 (N_49836,N_37727,N_37700);
xnor U49837 (N_49837,N_36822,N_37504);
xor U49838 (N_49838,N_39024,N_31714);
nor U49839 (N_49839,N_39583,N_30326);
nor U49840 (N_49840,N_35468,N_34210);
or U49841 (N_49841,N_35581,N_38162);
xor U49842 (N_49842,N_38354,N_30334);
nand U49843 (N_49843,N_30332,N_36278);
nor U49844 (N_49844,N_38656,N_38096);
nand U49845 (N_49845,N_34397,N_37351);
xnor U49846 (N_49846,N_30302,N_37107);
nand U49847 (N_49847,N_39771,N_33179);
nand U49848 (N_49848,N_37920,N_36094);
or U49849 (N_49849,N_37635,N_35720);
and U49850 (N_49850,N_31122,N_33184);
and U49851 (N_49851,N_36833,N_34356);
xnor U49852 (N_49852,N_34137,N_35739);
nand U49853 (N_49853,N_34163,N_35372);
or U49854 (N_49854,N_37749,N_38149);
nand U49855 (N_49855,N_33169,N_37372);
xor U49856 (N_49856,N_39980,N_31100);
nand U49857 (N_49857,N_33963,N_30399);
xor U49858 (N_49858,N_34937,N_35223);
nand U49859 (N_49859,N_30770,N_31896);
or U49860 (N_49860,N_36415,N_30360);
nand U49861 (N_49861,N_38704,N_33672);
nand U49862 (N_49862,N_30011,N_31238);
xnor U49863 (N_49863,N_38745,N_35289);
and U49864 (N_49864,N_34748,N_38923);
nand U49865 (N_49865,N_34508,N_34276);
nand U49866 (N_49866,N_30213,N_39558);
xor U49867 (N_49867,N_34262,N_30060);
or U49868 (N_49868,N_31147,N_33312);
or U49869 (N_49869,N_37309,N_33576);
nand U49870 (N_49870,N_35633,N_36086);
and U49871 (N_49871,N_34364,N_33293);
nand U49872 (N_49872,N_33813,N_31772);
and U49873 (N_49873,N_31769,N_31669);
nand U49874 (N_49874,N_39900,N_38412);
xor U49875 (N_49875,N_34816,N_35948);
nand U49876 (N_49876,N_31763,N_31834);
xnor U49877 (N_49877,N_34656,N_39051);
xor U49878 (N_49878,N_34666,N_30934);
and U49879 (N_49879,N_39473,N_32444);
or U49880 (N_49880,N_31193,N_31838);
nand U49881 (N_49881,N_38046,N_30417);
or U49882 (N_49882,N_35200,N_33039);
xnor U49883 (N_49883,N_36948,N_36401);
xor U49884 (N_49884,N_34555,N_30689);
and U49885 (N_49885,N_36370,N_38809);
or U49886 (N_49886,N_33195,N_38655);
or U49887 (N_49887,N_30053,N_35832);
and U49888 (N_49888,N_36254,N_33840);
nand U49889 (N_49889,N_30269,N_30894);
xor U49890 (N_49890,N_30433,N_34045);
or U49891 (N_49891,N_31282,N_37948);
or U49892 (N_49892,N_33206,N_39629);
or U49893 (N_49893,N_31684,N_32916);
or U49894 (N_49894,N_37761,N_35323);
and U49895 (N_49895,N_35353,N_34905);
nor U49896 (N_49896,N_31067,N_33982);
nand U49897 (N_49897,N_31778,N_32184);
nand U49898 (N_49898,N_34771,N_36017);
or U49899 (N_49899,N_38878,N_37183);
xor U49900 (N_49900,N_31093,N_34001);
nor U49901 (N_49901,N_36142,N_34076);
nor U49902 (N_49902,N_34043,N_36575);
xnor U49903 (N_49903,N_39338,N_38449);
xnor U49904 (N_49904,N_38694,N_37428);
nor U49905 (N_49905,N_31630,N_30391);
or U49906 (N_49906,N_32213,N_30744);
or U49907 (N_49907,N_30865,N_31780);
xor U49908 (N_49908,N_36065,N_35516);
nor U49909 (N_49909,N_39403,N_31060);
and U49910 (N_49910,N_31345,N_38000);
nand U49911 (N_49911,N_31442,N_37162);
nor U49912 (N_49912,N_37292,N_35973);
nand U49913 (N_49913,N_37056,N_30605);
and U49914 (N_49914,N_30718,N_34244);
nor U49915 (N_49915,N_31304,N_38595);
nand U49916 (N_49916,N_34885,N_32052);
or U49917 (N_49917,N_31048,N_35781);
nand U49918 (N_49918,N_30572,N_37569);
nand U49919 (N_49919,N_37537,N_33590);
xnor U49920 (N_49920,N_31981,N_39168);
or U49921 (N_49921,N_32731,N_36639);
nand U49922 (N_49922,N_37920,N_32739);
xor U49923 (N_49923,N_38130,N_38493);
xnor U49924 (N_49924,N_37637,N_37644);
xor U49925 (N_49925,N_30389,N_30820);
xor U49926 (N_49926,N_30004,N_30898);
nor U49927 (N_49927,N_32146,N_35765);
or U49928 (N_49928,N_31021,N_32758);
or U49929 (N_49929,N_30040,N_35533);
nand U49930 (N_49930,N_31365,N_31449);
nand U49931 (N_49931,N_30121,N_36846);
or U49932 (N_49932,N_37202,N_31988);
nor U49933 (N_49933,N_35925,N_38853);
and U49934 (N_49934,N_30054,N_38777);
and U49935 (N_49935,N_35298,N_30409);
nand U49936 (N_49936,N_39264,N_34281);
xor U49937 (N_49937,N_38015,N_34671);
nand U49938 (N_49938,N_34031,N_37061);
nor U49939 (N_49939,N_31631,N_37989);
or U49940 (N_49940,N_32275,N_34865);
or U49941 (N_49941,N_34177,N_33018);
xnor U49942 (N_49942,N_38243,N_36627);
and U49943 (N_49943,N_38410,N_35012);
nor U49944 (N_49944,N_32551,N_31746);
or U49945 (N_49945,N_30668,N_38334);
xor U49946 (N_49946,N_34415,N_35975);
nand U49947 (N_49947,N_37971,N_36641);
nand U49948 (N_49948,N_35821,N_35735);
nand U49949 (N_49949,N_38560,N_35809);
nor U49950 (N_49950,N_31837,N_33940);
or U49951 (N_49951,N_39314,N_31110);
nor U49952 (N_49952,N_30273,N_38017);
and U49953 (N_49953,N_37976,N_37720);
or U49954 (N_49954,N_39841,N_30628);
and U49955 (N_49955,N_37123,N_33906);
nand U49956 (N_49956,N_39624,N_33701);
and U49957 (N_49957,N_38896,N_39729);
nor U49958 (N_49958,N_34925,N_35378);
xnor U49959 (N_49959,N_30496,N_37088);
nor U49960 (N_49960,N_35242,N_34330);
nand U49961 (N_49961,N_31221,N_30152);
xor U49962 (N_49962,N_34221,N_32074);
nor U49963 (N_49963,N_39803,N_39019);
and U49964 (N_49964,N_39683,N_35381);
and U49965 (N_49965,N_33276,N_38937);
and U49966 (N_49966,N_38476,N_33119);
or U49967 (N_49967,N_32443,N_39890);
nand U49968 (N_49968,N_35380,N_31402);
nand U49969 (N_49969,N_30156,N_30582);
or U49970 (N_49970,N_38142,N_32067);
or U49971 (N_49971,N_39390,N_32127);
or U49972 (N_49972,N_31776,N_35156);
xnor U49973 (N_49973,N_34434,N_36083);
and U49974 (N_49974,N_39769,N_39681);
and U49975 (N_49975,N_35038,N_37912);
nor U49976 (N_49976,N_36871,N_38921);
nor U49977 (N_49977,N_36197,N_37926);
nor U49978 (N_49978,N_38563,N_35895);
xor U49979 (N_49979,N_33943,N_31127);
xor U49980 (N_49980,N_35755,N_36719);
and U49981 (N_49981,N_31104,N_38118);
xor U49982 (N_49982,N_34416,N_31016);
nand U49983 (N_49983,N_33033,N_37033);
nor U49984 (N_49984,N_30395,N_31983);
or U49985 (N_49985,N_30985,N_37982);
nand U49986 (N_49986,N_30366,N_31722);
nor U49987 (N_49987,N_36654,N_35895);
nor U49988 (N_49988,N_38232,N_38273);
or U49989 (N_49989,N_34051,N_34952);
or U49990 (N_49990,N_31711,N_30102);
xor U49991 (N_49991,N_31662,N_37215);
xor U49992 (N_49992,N_37470,N_33103);
nor U49993 (N_49993,N_38954,N_31928);
and U49994 (N_49994,N_36209,N_33582);
or U49995 (N_49995,N_37503,N_38233);
xor U49996 (N_49996,N_30574,N_35297);
and U49997 (N_49997,N_34345,N_36341);
nand U49998 (N_49998,N_33057,N_37973);
and U49999 (N_49999,N_37321,N_35440);
nand UO_0 (O_0,N_48799,N_48742);
nor UO_1 (O_1,N_48804,N_46075);
nor UO_2 (O_2,N_43400,N_40637);
or UO_3 (O_3,N_43945,N_40725);
nand UO_4 (O_4,N_49245,N_48508);
nand UO_5 (O_5,N_48450,N_47790);
xor UO_6 (O_6,N_47965,N_41202);
and UO_7 (O_7,N_47676,N_40345);
or UO_8 (O_8,N_43819,N_48261);
nor UO_9 (O_9,N_45771,N_48764);
or UO_10 (O_10,N_46022,N_44791);
and UO_11 (O_11,N_49711,N_44030);
or UO_12 (O_12,N_42437,N_44837);
or UO_13 (O_13,N_43078,N_45670);
and UO_14 (O_14,N_47878,N_40610);
and UO_15 (O_15,N_45225,N_49781);
and UO_16 (O_16,N_41027,N_45743);
and UO_17 (O_17,N_41833,N_41770);
and UO_18 (O_18,N_40801,N_47182);
xor UO_19 (O_19,N_46130,N_49316);
xnor UO_20 (O_20,N_41745,N_46366);
or UO_21 (O_21,N_41434,N_40533);
nor UO_22 (O_22,N_41251,N_42548);
nand UO_23 (O_23,N_47720,N_40228);
or UO_24 (O_24,N_49833,N_46499);
nor UO_25 (O_25,N_46098,N_44854);
and UO_26 (O_26,N_40082,N_45312);
xor UO_27 (O_27,N_43603,N_44072);
nor UO_28 (O_28,N_49162,N_40844);
xor UO_29 (O_29,N_40113,N_43794);
nor UO_30 (O_30,N_49199,N_49407);
xor UO_31 (O_31,N_41402,N_41535);
nand UO_32 (O_32,N_40507,N_49487);
nand UO_33 (O_33,N_40606,N_40485);
or UO_34 (O_34,N_49665,N_46551);
or UO_35 (O_35,N_41411,N_44116);
xor UO_36 (O_36,N_46239,N_41480);
and UO_37 (O_37,N_47364,N_49518);
and UO_38 (O_38,N_46603,N_44268);
or UO_39 (O_39,N_44331,N_42027);
xor UO_40 (O_40,N_49606,N_45440);
nor UO_41 (O_41,N_41812,N_42250);
xnor UO_42 (O_42,N_42935,N_46955);
nand UO_43 (O_43,N_46771,N_47012);
nand UO_44 (O_44,N_49271,N_43408);
or UO_45 (O_45,N_45847,N_47213);
nand UO_46 (O_46,N_48451,N_42738);
xnor UO_47 (O_47,N_42219,N_44488);
and UO_48 (O_48,N_42279,N_47898);
and UO_49 (O_49,N_44957,N_42628);
or UO_50 (O_50,N_48664,N_43834);
nor UO_51 (O_51,N_41664,N_42104);
xor UO_52 (O_52,N_48863,N_42699);
nand UO_53 (O_53,N_47804,N_42569);
nor UO_54 (O_54,N_42579,N_44240);
nor UO_55 (O_55,N_43123,N_43830);
or UO_56 (O_56,N_41070,N_45173);
nor UO_57 (O_57,N_42174,N_41879);
or UO_58 (O_58,N_49340,N_45020);
nor UO_59 (O_59,N_41954,N_47848);
xnor UO_60 (O_60,N_43740,N_41238);
or UO_61 (O_61,N_41672,N_43532);
xor UO_62 (O_62,N_46480,N_40183);
nor UO_63 (O_63,N_44598,N_48579);
xnor UO_64 (O_64,N_47264,N_42102);
xnor UO_65 (O_65,N_42070,N_47097);
and UO_66 (O_66,N_41688,N_43315);
or UO_67 (O_67,N_45716,N_44784);
and UO_68 (O_68,N_48629,N_43484);
xor UO_69 (O_69,N_46731,N_44689);
and UO_70 (O_70,N_45080,N_49584);
or UO_71 (O_71,N_41586,N_49838);
and UO_72 (O_72,N_41784,N_44735);
and UO_73 (O_73,N_44098,N_47124);
nand UO_74 (O_74,N_46328,N_42732);
xnor UO_75 (O_75,N_48921,N_49338);
xnor UO_76 (O_76,N_49075,N_45539);
or UO_77 (O_77,N_44343,N_45029);
nand UO_78 (O_78,N_47415,N_42064);
nand UO_79 (O_79,N_48589,N_46755);
xor UO_80 (O_80,N_41676,N_49698);
and UO_81 (O_81,N_40056,N_44363);
or UO_82 (O_82,N_48235,N_40708);
and UO_83 (O_83,N_42260,N_45710);
or UO_84 (O_84,N_48416,N_41838);
xor UO_85 (O_85,N_42186,N_40402);
nor UO_86 (O_86,N_46833,N_46193);
nand UO_87 (O_87,N_49658,N_46386);
nor UO_88 (O_88,N_44017,N_46292);
and UO_89 (O_89,N_49125,N_43501);
nor UO_90 (O_90,N_47277,N_45501);
xor UO_91 (O_91,N_48280,N_40969);
and UO_92 (O_92,N_44053,N_47300);
and UO_93 (O_93,N_43827,N_42623);
or UO_94 (O_94,N_45134,N_45698);
nand UO_95 (O_95,N_44541,N_48350);
nand UO_96 (O_96,N_45298,N_42333);
nand UO_97 (O_97,N_49809,N_48727);
nor UO_98 (O_98,N_41796,N_48705);
and UO_99 (O_99,N_49031,N_46946);
nand UO_100 (O_100,N_40780,N_46760);
and UO_101 (O_101,N_47006,N_46536);
nand UO_102 (O_102,N_48728,N_45317);
xor UO_103 (O_103,N_48975,N_44140);
nand UO_104 (O_104,N_49250,N_49685);
or UO_105 (O_105,N_46943,N_43682);
nand UO_106 (O_106,N_45723,N_41347);
nand UO_107 (O_107,N_48906,N_45232);
and UO_108 (O_108,N_47682,N_49336);
or UO_109 (O_109,N_46883,N_42149);
nor UO_110 (O_110,N_41963,N_46406);
xor UO_111 (O_111,N_42977,N_48077);
nor UO_112 (O_112,N_43674,N_48121);
and UO_113 (O_113,N_47286,N_44913);
nor UO_114 (O_114,N_46264,N_44882);
and UO_115 (O_115,N_41523,N_43703);
and UO_116 (O_116,N_42883,N_46250);
or UO_117 (O_117,N_45850,N_47601);
nor UO_118 (O_118,N_40456,N_42600);
nand UO_119 (O_119,N_46886,N_45429);
or UO_120 (O_120,N_43082,N_41349);
or UO_121 (O_121,N_45988,N_42286);
and UO_122 (O_122,N_49703,N_48560);
and UO_123 (O_123,N_46361,N_40008);
and UO_124 (O_124,N_42014,N_49376);
nand UO_125 (O_125,N_41787,N_49810);
nand UO_126 (O_126,N_41379,N_43370);
xor UO_127 (O_127,N_44225,N_49986);
nor UO_128 (O_128,N_47108,N_44937);
nand UO_129 (O_129,N_47853,N_41038);
nand UO_130 (O_130,N_42870,N_40842);
or UO_131 (O_131,N_40006,N_48187);
nand UO_132 (O_132,N_45068,N_41339);
or UO_133 (O_133,N_49130,N_47054);
and UO_134 (O_134,N_48362,N_40119);
or UO_135 (O_135,N_49650,N_46985);
nor UO_136 (O_136,N_47971,N_46173);
nand UO_137 (O_137,N_44632,N_45144);
or UO_138 (O_138,N_49668,N_40281);
nand UO_139 (O_139,N_48564,N_41799);
nand UO_140 (O_140,N_40715,N_45923);
nor UO_141 (O_141,N_40546,N_43722);
xor UO_142 (O_142,N_41021,N_44771);
nand UO_143 (O_143,N_41320,N_40325);
or UO_144 (O_144,N_43909,N_44495);
nor UO_145 (O_145,N_49531,N_42380);
nor UO_146 (O_146,N_46839,N_46278);
nor UO_147 (O_147,N_48284,N_44533);
nor UO_148 (O_148,N_49677,N_42399);
nor UO_149 (O_149,N_44016,N_42488);
and UO_150 (O_150,N_41362,N_43994);
or UO_151 (O_151,N_44704,N_41847);
xnor UO_152 (O_152,N_49867,N_44415);
and UO_153 (O_153,N_46314,N_42118);
nor UO_154 (O_154,N_48485,N_45950);
nand UO_155 (O_155,N_43684,N_42123);
or UO_156 (O_156,N_40732,N_43153);
nor UO_157 (O_157,N_44588,N_46524);
xnor UO_158 (O_158,N_49999,N_40103);
or UO_159 (O_159,N_45782,N_40282);
nand UO_160 (O_160,N_40256,N_48269);
and UO_161 (O_161,N_41735,N_41880);
nor UO_162 (O_162,N_43912,N_46769);
xnor UO_163 (O_163,N_46368,N_43330);
and UO_164 (O_164,N_46681,N_43061);
nor UO_165 (O_165,N_45388,N_48022);
nand UO_166 (O_166,N_43218,N_42841);
nor UO_167 (O_167,N_42898,N_48957);
nor UO_168 (O_168,N_41699,N_49533);
xor UO_169 (O_169,N_44557,N_45564);
nor UO_170 (O_170,N_41080,N_42817);
nor UO_171 (O_171,N_42606,N_49847);
or UO_172 (O_172,N_49219,N_45062);
or UO_173 (O_173,N_49875,N_43428);
xnor UO_174 (O_174,N_41520,N_46349);
xor UO_175 (O_175,N_43731,N_41452);
or UO_176 (O_176,N_49649,N_40618);
and UO_177 (O_177,N_43190,N_42253);
xnor UO_178 (O_178,N_43103,N_43891);
or UO_179 (O_179,N_47693,N_42926);
nand UO_180 (O_180,N_48395,N_49737);
nand UO_181 (O_181,N_47942,N_40661);
xnor UO_182 (O_182,N_46186,N_49221);
and UO_183 (O_183,N_45686,N_48905);
nand UO_184 (O_184,N_46261,N_49390);
or UO_185 (O_185,N_47732,N_48075);
nor UO_186 (O_186,N_40540,N_41892);
and UO_187 (O_187,N_45944,N_41874);
xor UO_188 (O_188,N_46904,N_42204);
nor UO_189 (O_189,N_48273,N_49172);
nor UO_190 (O_190,N_49959,N_43583);
nor UO_191 (O_191,N_40852,N_49415);
nand UO_192 (O_192,N_48923,N_43777);
nand UO_193 (O_193,N_49149,N_41924);
xnor UO_194 (O_194,N_47196,N_45628);
nor UO_195 (O_195,N_44402,N_47259);
xnor UO_196 (O_196,N_47708,N_40355);
and UO_197 (O_197,N_46449,N_48049);
or UO_198 (O_198,N_43768,N_41162);
or UO_199 (O_199,N_40014,N_40846);
xor UO_200 (O_200,N_40531,N_42509);
nor UO_201 (O_201,N_41921,N_45302);
or UO_202 (O_202,N_44004,N_47214);
xor UO_203 (O_203,N_41648,N_43820);
and UO_204 (O_204,N_47153,N_49187);
and UO_205 (O_205,N_42630,N_43277);
xor UO_206 (O_206,N_48058,N_45049);
and UO_207 (O_207,N_47842,N_41894);
nor UO_208 (O_208,N_40127,N_41455);
and UO_209 (O_209,N_49601,N_48697);
and UO_210 (O_210,N_48237,N_42799);
nor UO_211 (O_211,N_48625,N_46573);
and UO_212 (O_212,N_44187,N_44730);
xnor UO_213 (O_213,N_43981,N_44182);
xnor UO_214 (O_214,N_47761,N_47792);
or UO_215 (O_215,N_42938,N_48402);
and UO_216 (O_216,N_48675,N_40687);
xnor UO_217 (O_217,N_47184,N_40776);
or UO_218 (O_218,N_45600,N_43558);
or UO_219 (O_219,N_45667,N_49284);
xnor UO_220 (O_220,N_49943,N_42324);
nand UO_221 (O_221,N_41476,N_42726);
nor UO_222 (O_222,N_42495,N_45665);
xor UO_223 (O_223,N_40720,N_44911);
and UO_224 (O_224,N_45088,N_40356);
or UO_225 (O_225,N_45450,N_49727);
xor UO_226 (O_226,N_40554,N_40459);
and UO_227 (O_227,N_42491,N_49528);
or UO_228 (O_228,N_40105,N_42262);
nand UO_229 (O_229,N_43470,N_49150);
xnor UO_230 (O_230,N_46209,N_47207);
xor UO_231 (O_231,N_42494,N_48860);
xnor UO_232 (O_232,N_42599,N_47465);
nand UO_233 (O_233,N_40855,N_44982);
nand UO_234 (O_234,N_44659,N_49767);
or UO_235 (O_235,N_47913,N_42216);
and UO_236 (O_236,N_40437,N_48744);
nand UO_237 (O_237,N_40481,N_40128);
nor UO_238 (O_238,N_47065,N_47657);
and UO_239 (O_239,N_40227,N_42603);
nand UO_240 (O_240,N_43813,N_45504);
xor UO_241 (O_241,N_48912,N_45683);
nor UO_242 (O_242,N_44869,N_43709);
nand UO_243 (O_243,N_41227,N_44508);
and UO_244 (O_244,N_40676,N_43495);
or UO_245 (O_245,N_46992,N_42200);
or UO_246 (O_246,N_47789,N_47231);
xnor UO_247 (O_247,N_48616,N_44699);
nand UO_248 (O_248,N_46175,N_43095);
xor UO_249 (O_249,N_42087,N_41544);
nor UO_250 (O_250,N_46854,N_46893);
nand UO_251 (O_251,N_47326,N_42355);
or UO_252 (O_252,N_45689,N_46581);
and UO_253 (O_253,N_42775,N_46652);
nor UO_254 (O_254,N_40999,N_49255);
and UO_255 (O_255,N_43167,N_45579);
or UO_256 (O_256,N_43866,N_47610);
or UO_257 (O_257,N_49917,N_46122);
nand UO_258 (O_258,N_46230,N_43225);
and UO_259 (O_259,N_44968,N_41242);
nor UO_260 (O_260,N_49530,N_47268);
nand UO_261 (O_261,N_48334,N_44696);
and UO_262 (O_262,N_49371,N_47426);
xor UO_263 (O_263,N_41607,N_42414);
or UO_264 (O_264,N_41494,N_47953);
or UO_265 (O_265,N_47532,N_44486);
and UO_266 (O_266,N_44757,N_46443);
nand UO_267 (O_267,N_44191,N_47880);
nand UO_268 (O_268,N_42939,N_48915);
nor UO_269 (O_269,N_44700,N_43630);
nand UO_270 (O_270,N_48035,N_45191);
nand UO_271 (O_271,N_42947,N_40972);
and UO_272 (O_272,N_46749,N_43179);
nor UO_273 (O_273,N_49246,N_49373);
or UO_274 (O_274,N_42221,N_43798);
and UO_275 (O_275,N_43003,N_40622);
xor UO_276 (O_276,N_45468,N_40754);
xnor UO_277 (O_277,N_45706,N_47018);
and UO_278 (O_278,N_48472,N_45864);
or UO_279 (O_279,N_48198,N_40392);
nor UO_280 (O_280,N_42681,N_45510);
nand UO_281 (O_281,N_47979,N_40552);
nor UO_282 (O_282,N_41772,N_47452);
nand UO_283 (O_283,N_43067,N_49783);
nand UO_284 (O_284,N_42465,N_41908);
nor UO_285 (O_285,N_44944,N_48342);
and UO_286 (O_286,N_46068,N_40050);
nand UO_287 (O_287,N_46432,N_45596);
xnor UO_288 (O_288,N_43520,N_46059);
or UO_289 (O_289,N_49570,N_43241);
nor UO_290 (O_290,N_41629,N_42311);
xor UO_291 (O_291,N_41791,N_43069);
xnor UO_292 (O_292,N_44774,N_43134);
nand UO_293 (O_293,N_42911,N_42398);
or UO_294 (O_294,N_46612,N_43138);
nand UO_295 (O_295,N_42301,N_46707);
xor UO_296 (O_296,N_46715,N_49561);
and UO_297 (O_297,N_42546,N_43465);
or UO_298 (O_298,N_46852,N_42659);
or UO_299 (O_299,N_45435,N_47649);
and UO_300 (O_300,N_40727,N_48977);
nor UO_301 (O_301,N_49134,N_42830);
nor UO_302 (O_302,N_40809,N_48471);
nor UO_303 (O_303,N_47162,N_45848);
nand UO_304 (O_304,N_40216,N_48248);
xnor UO_305 (O_305,N_42631,N_46564);
nand UO_306 (O_306,N_49424,N_45893);
nand UO_307 (O_307,N_44956,N_49059);
and UO_308 (O_308,N_41804,N_46004);
and UO_309 (O_309,N_49967,N_40018);
nor UO_310 (O_310,N_45476,N_43775);
and UO_311 (O_311,N_46305,N_44190);
xor UO_312 (O_312,N_48862,N_44725);
or UO_313 (O_313,N_44767,N_43662);
or UO_314 (O_314,N_41660,N_43568);
xor UO_315 (O_315,N_40423,N_45207);
or UO_316 (O_316,N_49135,N_43743);
xnor UO_317 (O_317,N_45226,N_47360);
nand UO_318 (O_318,N_49922,N_41415);
or UO_319 (O_319,N_42321,N_46620);
xnor UO_320 (O_320,N_46977,N_46017);
and UO_321 (O_321,N_46351,N_48833);
or UO_322 (O_322,N_43036,N_46509);
xor UO_323 (O_323,N_42427,N_49716);
xor UO_324 (O_324,N_47195,N_42065);
xnor UO_325 (O_325,N_48539,N_46647);
xnor UO_326 (O_326,N_45913,N_42627);
nand UO_327 (O_327,N_42275,N_47046);
xor UO_328 (O_328,N_45774,N_42902);
or UO_329 (O_329,N_45406,N_49060);
nand UO_330 (O_330,N_43156,N_49542);
nand UO_331 (O_331,N_40781,N_44890);
xnor UO_332 (O_332,N_44916,N_41895);
or UO_333 (O_333,N_47907,N_45582);
and UO_334 (O_334,N_43097,N_44277);
and UO_335 (O_335,N_42101,N_46088);
nand UO_336 (O_336,N_47467,N_49718);
or UO_337 (O_337,N_41128,N_43679);
and UO_338 (O_338,N_40884,N_40269);
nand UO_339 (O_339,N_48766,N_47189);
xor UO_340 (O_340,N_47916,N_42624);
nor UO_341 (O_341,N_42930,N_46685);
or UO_342 (O_342,N_49025,N_46665);
nand UO_343 (O_343,N_48965,N_47631);
or UO_344 (O_344,N_47509,N_46429);
or UO_345 (O_345,N_46631,N_46296);
xor UO_346 (O_346,N_48515,N_48099);
nand UO_347 (O_347,N_48120,N_46338);
nor UO_348 (O_348,N_48946,N_42928);
nand UO_349 (O_349,N_49043,N_49078);
nand UO_350 (O_350,N_40005,N_49916);
and UO_351 (O_351,N_45684,N_43851);
xnor UO_352 (O_352,N_44137,N_48790);
xnor UO_353 (O_353,N_49051,N_49450);
and UO_354 (O_354,N_41596,N_41194);
or UO_355 (O_355,N_47626,N_44170);
nand UO_356 (O_356,N_49853,N_46479);
nand UO_357 (O_357,N_45046,N_43210);
and UO_358 (O_358,N_45557,N_40155);
nor UO_359 (O_359,N_45480,N_42776);
nand UO_360 (O_360,N_40283,N_43713);
nand UO_361 (O_361,N_40527,N_45221);
or UO_362 (O_362,N_43347,N_43290);
and UO_363 (O_363,N_42580,N_45410);
nand UO_364 (O_364,N_49395,N_44946);
nand UO_365 (O_365,N_45428,N_46339);
and UO_366 (O_366,N_42474,N_42078);
or UO_367 (O_367,N_41143,N_44193);
xnor UO_368 (O_368,N_45238,N_46998);
xor UO_369 (O_369,N_46930,N_42288);
nand UO_370 (O_370,N_46326,N_44840);
and UO_371 (O_371,N_41670,N_49539);
xor UO_372 (O_372,N_46225,N_45294);
nor UO_373 (O_373,N_43320,N_43286);
and UO_374 (O_374,N_40763,N_48392);
and UO_375 (O_375,N_41108,N_47021);
nor UO_376 (O_376,N_45933,N_47681);
or UO_377 (O_377,N_48148,N_47968);
or UO_378 (O_378,N_48428,N_48888);
nor UO_379 (O_379,N_45282,N_45015);
nand UO_380 (O_380,N_43302,N_44858);
nand UO_381 (O_381,N_42910,N_46739);
nor UO_382 (O_382,N_47332,N_42593);
or UO_383 (O_383,N_41440,N_42813);
nand UO_384 (O_384,N_40002,N_47926);
nand UO_385 (O_385,N_48740,N_41208);
nor UO_386 (O_386,N_40381,N_45650);
and UO_387 (O_387,N_44104,N_44902);
xor UO_388 (O_388,N_48666,N_49864);
nand UO_389 (O_389,N_43058,N_43281);
nor UO_390 (O_390,N_48669,N_40820);
nor UO_391 (O_391,N_43178,N_43448);
nor UO_392 (O_392,N_41722,N_42236);
or UO_393 (O_393,N_47106,N_45956);
xor UO_394 (O_394,N_46084,N_48481);
nand UO_395 (O_395,N_48702,N_40466);
or UO_396 (O_396,N_43161,N_43808);
or UO_397 (O_397,N_44487,N_41114);
nor UO_398 (O_398,N_48151,N_40460);
nand UO_399 (O_399,N_46313,N_41717);
nand UO_400 (O_400,N_44069,N_46144);
xor UO_401 (O_401,N_47001,N_42337);
nor UO_402 (O_402,N_43262,N_41465);
xor UO_403 (O_403,N_45714,N_47791);
nor UO_404 (O_404,N_48465,N_40901);
and UO_405 (O_405,N_44607,N_44811);
or UO_406 (O_406,N_42093,N_43610);
and UO_407 (O_407,N_46301,N_42467);
xor UO_408 (O_408,N_46293,N_44223);
nor UO_409 (O_409,N_44953,N_47574);
and UO_410 (O_410,N_49826,N_45516);
and UO_411 (O_411,N_46216,N_46450);
nor UO_412 (O_412,N_48903,N_43666);
and UO_413 (O_413,N_40340,N_43803);
nor UO_414 (O_414,N_43734,N_41429);
nand UO_415 (O_415,N_41539,N_47174);
and UO_416 (O_416,N_45535,N_47923);
and UO_417 (O_417,N_42721,N_41158);
xor UO_418 (O_418,N_45651,N_49223);
or UO_419 (O_419,N_45407,N_47542);
nand UO_420 (O_420,N_47747,N_42743);
and UO_421 (O_421,N_49572,N_45619);
nor UO_422 (O_422,N_48880,N_47592);
and UO_423 (O_423,N_46751,N_44479);
nor UO_424 (O_424,N_49046,N_46012);
nor UO_425 (O_425,N_45140,N_49910);
nor UO_426 (O_426,N_40701,N_45443);
nand UO_427 (O_427,N_44947,N_44773);
nand UO_428 (O_428,N_48813,N_43432);
xor UO_429 (O_429,N_47352,N_41635);
and UO_430 (O_430,N_49926,N_46912);
xor UO_431 (O_431,N_40665,N_42966);
and UO_432 (O_432,N_47550,N_42673);
nor UO_433 (O_433,N_48511,N_48249);
xnor UO_434 (O_434,N_42945,N_43599);
or UO_435 (O_435,N_41538,N_46006);
and UO_436 (O_436,N_41444,N_48142);
nor UO_437 (O_437,N_41447,N_40112);
xnor UO_438 (O_438,N_41154,N_47102);
nand UO_439 (O_439,N_48476,N_47707);
xor UO_440 (O_440,N_43200,N_43533);
or UO_441 (O_441,N_42317,N_44192);
nand UO_442 (O_442,N_42396,N_47808);
nor UO_443 (O_443,N_48192,N_41926);
nand UO_444 (O_444,N_41568,N_45506);
and UO_445 (O_445,N_49388,N_44905);
nand UO_446 (O_446,N_47024,N_45425);
or UO_447 (O_447,N_44915,N_43009);
and UO_448 (O_448,N_47247,N_42995);
xor UO_449 (O_449,N_42979,N_45102);
or UO_450 (O_450,N_41861,N_41706);
nor UO_451 (O_451,N_41746,N_46360);
or UO_452 (O_452,N_45803,N_40523);
and UO_453 (O_453,N_43450,N_46824);
and UO_454 (O_454,N_41253,N_43992);
and UO_455 (O_455,N_49988,N_43787);
and UO_456 (O_456,N_46658,N_41189);
and UO_457 (O_457,N_48756,N_44395);
nor UO_458 (O_458,N_44686,N_46735);
nor UO_459 (O_459,N_42676,N_45441);
nand UO_460 (O_460,N_47407,N_44741);
xnor UO_461 (O_461,N_43964,N_40304);
and UO_462 (O_462,N_42805,N_43672);
nand UO_463 (O_463,N_42475,N_45041);
nor UO_464 (O_464,N_41293,N_42794);
nor UO_465 (O_465,N_49800,N_47941);
nor UO_466 (O_466,N_48063,N_48712);
or UO_467 (O_467,N_43223,N_49742);
nand UO_468 (O_468,N_46420,N_49356);
xnor UO_469 (O_469,N_44792,N_48635);
or UO_470 (O_470,N_45917,N_49965);
nand UO_471 (O_471,N_48798,N_42780);
xnor UO_472 (O_472,N_40859,N_49869);
and UO_473 (O_473,N_49378,N_49646);
nor UO_474 (O_474,N_44406,N_41017);
and UO_475 (O_475,N_41416,N_42556);
xor UO_476 (O_476,N_48067,N_49554);
xor UO_477 (O_477,N_48165,N_43751);
nor UO_478 (O_478,N_49144,N_40066);
nor UO_479 (O_479,N_47016,N_46947);
xnor UO_480 (O_480,N_44025,N_40782);
nor UO_481 (O_481,N_45345,N_47358);
nor UO_482 (O_482,N_44247,N_49501);
xor UO_483 (O_483,N_46910,N_48716);
nor UO_484 (O_484,N_44684,N_40992);
and UO_485 (O_485,N_44646,N_40913);
and UO_486 (O_486,N_44856,N_42130);
and UO_487 (O_487,N_46738,N_49746);
or UO_488 (O_488,N_40952,N_46692);
nor UO_489 (O_489,N_45035,N_49233);
nor UO_490 (O_490,N_49923,N_47490);
nor UO_491 (O_491,N_49169,N_47958);
or UO_492 (O_492,N_42657,N_42406);
nand UO_493 (O_493,N_44474,N_40010);
nand UO_494 (O_494,N_43585,N_41666);
nor UO_495 (O_495,N_45508,N_45204);
nor UO_496 (O_496,N_43415,N_47608);
nor UO_497 (O_497,N_49722,N_41404);
and UO_498 (O_498,N_43749,N_44466);
nand UO_499 (O_499,N_48137,N_44822);
xor UO_500 (O_500,N_45150,N_45892);
xor UO_501 (O_501,N_44350,N_48636);
nand UO_502 (O_502,N_43860,N_42063);
and UO_503 (O_503,N_43643,N_47173);
and UO_504 (O_504,N_48112,N_49799);
or UO_505 (O_505,N_47545,N_44300);
and UO_506 (O_506,N_48991,N_49322);
nor UO_507 (O_507,N_43268,N_46284);
nand UO_508 (O_508,N_45056,N_46106);
or UO_509 (O_509,N_40519,N_49311);
nand UO_510 (O_510,N_45768,N_40030);
and UO_511 (O_511,N_44385,N_40099);
nand UO_512 (O_512,N_49556,N_40871);
nand UO_513 (O_513,N_47158,N_45636);
and UO_514 (O_514,N_44745,N_40141);
nor UO_515 (O_515,N_40612,N_48300);
xnor UO_516 (O_516,N_46829,N_41530);
xnor UO_517 (O_517,N_48676,N_45172);
nor UO_518 (O_518,N_49489,N_46819);
or UO_519 (O_519,N_48305,N_40551);
and UO_520 (O_520,N_42410,N_49166);
nand UO_521 (O_521,N_47678,N_47688);
xor UO_522 (O_522,N_46444,N_45348);
and UO_523 (O_523,N_49843,N_43882);
nor UO_524 (O_524,N_41782,N_49108);
nor UO_525 (O_525,N_46931,N_49204);
nor UO_526 (O_526,N_44619,N_48167);
or UO_527 (O_527,N_41378,N_42887);
and UO_528 (O_528,N_47684,N_46909);
nor UO_529 (O_529,N_40961,N_45084);
and UO_530 (O_530,N_49890,N_47513);
or UO_531 (O_531,N_43874,N_41822);
nand UO_532 (O_532,N_43079,N_45614);
and UO_533 (O_533,N_46269,N_44942);
xnor UO_534 (O_534,N_42862,N_42851);
nor UO_535 (O_535,N_45044,N_42493);
nand UO_536 (O_536,N_42549,N_47921);
nand UO_537 (O_537,N_47483,N_41443);
or UO_538 (O_538,N_42239,N_45167);
xor UO_539 (O_539,N_41226,N_40603);
nand UO_540 (O_540,N_46661,N_45949);
nor UO_541 (O_541,N_44088,N_42590);
xor UO_542 (O_542,N_48414,N_41508);
and UO_543 (O_543,N_48045,N_48528);
nand UO_544 (O_544,N_44755,N_46873);
nand UO_545 (O_545,N_45760,N_42099);
nor UO_546 (O_546,N_46978,N_46989);
xor UO_547 (O_547,N_49588,N_46740);
and UO_548 (O_548,N_49182,N_40627);
xnor UO_549 (O_549,N_45820,N_47497);
xnor UO_550 (O_550,N_47711,N_40748);
xor UO_551 (O_551,N_49788,N_45141);
nor UO_552 (O_552,N_49260,N_42080);
and UO_553 (O_553,N_40303,N_45234);
or UO_554 (O_554,N_43870,N_49990);
and UO_555 (O_555,N_42484,N_44621);
and UO_556 (O_556,N_43243,N_40445);
and UO_557 (O_557,N_45484,N_42140);
or UO_558 (O_558,N_49014,N_45824);
xor UO_559 (O_559,N_49759,N_48190);
and UO_560 (O_560,N_49891,N_42829);
nor UO_561 (O_561,N_44967,N_42019);
nand UO_562 (O_562,N_48869,N_44812);
and UO_563 (O_563,N_47655,N_48943);
or UO_564 (O_564,N_44976,N_43116);
or UO_565 (O_565,N_41521,N_48118);
or UO_566 (O_566,N_48382,N_43496);
nand UO_567 (O_567,N_42214,N_41781);
nand UO_568 (O_568,N_43349,N_49614);
and UO_569 (O_569,N_47623,N_44929);
nand UO_570 (O_570,N_44515,N_42418);
nand UO_571 (O_571,N_45007,N_44794);
xor UO_572 (O_572,N_49414,N_49040);
or UO_573 (O_573,N_40184,N_41888);
nand UO_574 (O_574,N_40317,N_46862);
nand UO_575 (O_575,N_48150,N_41517);
xor UO_576 (O_576,N_42532,N_48442);
or UO_577 (O_577,N_41636,N_47130);
and UO_578 (O_578,N_47015,N_40953);
xnor UO_579 (O_579,N_47367,N_46503);
and UO_580 (O_580,N_41184,N_49256);
nand UO_581 (O_581,N_47679,N_42617);
or UO_582 (O_582,N_43442,N_40198);
nor UO_583 (O_583,N_48649,N_45648);
xor UO_584 (O_584,N_41369,N_41277);
xnor UO_585 (O_585,N_43598,N_40511);
nand UO_586 (O_586,N_43596,N_49710);
and UO_587 (O_587,N_45748,N_43013);
or UO_588 (O_588,N_45606,N_45158);
nand UO_589 (O_589,N_44647,N_44601);
nand UO_590 (O_590,N_47924,N_44377);
xor UO_591 (O_591,N_43064,N_46856);
nand UO_592 (O_592,N_41506,N_48461);
xor UO_593 (O_593,N_49622,N_47390);
or UO_594 (O_594,N_41509,N_41621);
nor UO_595 (O_595,N_42293,N_47448);
xor UO_596 (O_596,N_46549,N_49023);
nand UO_597 (O_597,N_46241,N_45324);
nor UO_598 (O_598,N_47354,N_43386);
and UO_599 (O_599,N_43831,N_41471);
xnor UO_600 (O_600,N_49540,N_48762);
or UO_601 (O_601,N_49196,N_40768);
and UO_602 (O_602,N_48535,N_45066);
xor UO_603 (O_603,N_41827,N_45520);
or UO_604 (O_604,N_42021,N_46513);
and UO_605 (O_605,N_44407,N_44398);
nand UO_606 (O_606,N_49849,N_48939);
and UO_607 (O_607,N_45479,N_42480);
or UO_608 (O_608,N_49748,N_42141);
nand UO_609 (O_609,N_47172,N_43507);
xor UO_610 (O_610,N_40742,N_44555);
nor UO_611 (O_611,N_49217,N_48299);
nor UO_612 (O_612,N_42458,N_43015);
xor UO_613 (O_613,N_44878,N_45011);
xnor UO_614 (O_614,N_41734,N_43293);
xor UO_615 (O_615,N_42125,N_40709);
or UO_616 (O_616,N_49386,N_46795);
xnor UO_617 (O_617,N_49112,N_44113);
or UO_618 (O_618,N_47793,N_46590);
nand UO_619 (O_619,N_44203,N_48226);
nand UO_620 (O_620,N_42561,N_43300);
or UO_621 (O_621,N_45155,N_48030);
and UO_622 (O_622,N_49253,N_41858);
and UO_623 (O_623,N_48797,N_48674);
nand UO_624 (O_624,N_44955,N_42455);
xor UO_625 (O_625,N_48751,N_47872);
or UO_626 (O_626,N_42340,N_44396);
nor UO_627 (O_627,N_43051,N_42810);
nand UO_628 (O_628,N_41317,N_40408);
nand UO_629 (O_629,N_44476,N_46858);
or UO_630 (O_630,N_44954,N_45869);
and UO_631 (O_631,N_41644,N_46981);
and UO_632 (O_632,N_43758,N_49480);
nor UO_633 (O_633,N_45076,N_40417);
nor UO_634 (O_634,N_44275,N_40578);
or UO_635 (O_635,N_45807,N_40470);
or UO_636 (O_636,N_48052,N_41802);
or UO_637 (O_637,N_49824,N_47972);
nand UO_638 (O_638,N_48757,N_43207);
xor UO_639 (O_639,N_48598,N_49403);
xor UO_640 (O_640,N_42941,N_49165);
nor UO_641 (O_641,N_47283,N_44814);
nor UO_642 (O_642,N_47593,N_41069);
or UO_643 (O_643,N_40090,N_47307);
xnor UO_644 (O_644,N_46962,N_45971);
xor UO_645 (O_645,N_46892,N_48670);
xnor UO_646 (O_646,N_43502,N_42412);
or UO_647 (O_647,N_48854,N_40563);
xnor UO_648 (O_648,N_49947,N_41939);
or UO_649 (O_649,N_49538,N_42710);
nor UO_650 (O_650,N_46580,N_46853);
xnor UO_651 (O_651,N_45727,N_43747);
nand UO_652 (O_652,N_43350,N_40258);
nand UO_653 (O_653,N_47298,N_49009);
xor UO_654 (O_654,N_47904,N_41742);
xor UO_655 (O_655,N_40851,N_44156);
nor UO_656 (O_656,N_46214,N_45091);
or UO_657 (O_657,N_45839,N_47868);
nor UO_658 (O_658,N_42518,N_43043);
nand UO_659 (O_659,N_48955,N_42405);
or UO_660 (O_660,N_40452,N_44232);
xnor UO_661 (O_661,N_43383,N_43625);
nor UO_662 (O_662,N_44471,N_48453);
nand UO_663 (O_663,N_40352,N_44020);
or UO_664 (O_664,N_44400,N_48021);
or UO_665 (O_665,N_44889,N_40226);
nand UO_666 (O_666,N_42004,N_42271);
or UO_667 (O_667,N_44510,N_46772);
and UO_668 (O_668,N_40587,N_41260);
and UO_669 (O_669,N_47546,N_42062);
or UO_670 (O_670,N_47948,N_49167);
nor UO_671 (O_671,N_40262,N_40499);
xnor UO_672 (O_672,N_44567,N_40872);
or UO_673 (O_673,N_41139,N_49892);
xor UO_674 (O_674,N_45146,N_45875);
nor UO_675 (O_675,N_43405,N_44742);
or UO_676 (O_676,N_49585,N_46598);
xnor UO_677 (O_677,N_40261,N_49859);
or UO_678 (O_678,N_46409,N_48484);
xor UO_679 (O_679,N_44802,N_41074);
nand UO_680 (O_680,N_48236,N_49281);
nor UO_681 (O_681,N_47599,N_42595);
xnor UO_682 (O_682,N_42136,N_43185);
xnor UO_683 (O_683,N_40919,N_49024);
nand UO_684 (O_684,N_42124,N_47457);
xnor UO_685 (O_685,N_45630,N_49422);
nand UO_686 (O_686,N_42225,N_47537);
nor UO_687 (O_687,N_44039,N_48095);
nand UO_688 (O_688,N_47909,N_41830);
and UO_689 (O_689,N_48298,N_49369);
or UO_690 (O_690,N_45528,N_43401);
nand UO_691 (O_691,N_44279,N_46340);
nand UO_692 (O_692,N_42198,N_47361);
nor UO_693 (O_693,N_48029,N_40971);
nand UO_694 (O_694,N_47180,N_44928);
xnor UO_695 (O_695,N_44451,N_40967);
nor UO_696 (O_696,N_45199,N_40833);
xor UO_697 (O_697,N_40858,N_48631);
or UO_698 (O_698,N_40372,N_40922);
nor UO_699 (O_699,N_40195,N_47806);
xnor UO_700 (O_700,N_40493,N_46894);
xnor UO_701 (O_701,N_45178,N_47271);
or UO_702 (O_702,N_44836,N_45680);
and UO_703 (O_703,N_44171,N_43491);
xnor UO_704 (O_704,N_42356,N_43712);
or UO_705 (O_705,N_43962,N_42079);
nand UO_706 (O_706,N_41533,N_40327);
nor UO_707 (O_707,N_44697,N_47612);
nand UO_708 (O_708,N_46454,N_46754);
nand UO_709 (O_709,N_47700,N_42615);
and UO_710 (O_710,N_43956,N_41510);
and UO_711 (O_711,N_48686,N_41424);
nand UO_712 (O_712,N_49007,N_41156);
nor UO_713 (O_713,N_44241,N_48245);
nand UO_714 (O_714,N_47920,N_46111);
and UO_715 (O_715,N_49637,N_44166);
nand UO_716 (O_716,N_45393,N_45712);
xor UO_717 (O_717,N_45057,N_47787);
nand UO_718 (O_718,N_45898,N_41460);
or UO_719 (O_719,N_44332,N_41913);
nand UO_720 (O_720,N_49069,N_49975);
nor UO_721 (O_721,N_44583,N_40984);
nand UO_722 (O_722,N_40779,N_47111);
nor UO_723 (O_723,N_46457,N_49638);
and UO_724 (O_724,N_43889,N_41200);
nor UO_725 (O_725,N_42090,N_41902);
xor UO_726 (O_726,N_43551,N_46126);
nor UO_727 (O_727,N_42755,N_48262);
xor UO_728 (O_728,N_45401,N_48657);
xnor UO_729 (O_729,N_41147,N_41964);
or UO_730 (O_730,N_40509,N_42049);
xnor UO_731 (O_731,N_42648,N_44125);
nand UO_732 (O_732,N_44142,N_43779);
or UO_733 (O_733,N_42089,N_45395);
nand UO_734 (O_734,N_45494,N_45036);
nor UO_735 (O_735,N_46714,N_48223);
nand UO_736 (O_736,N_49913,N_47396);
nand UO_737 (O_737,N_42166,N_44724);
or UO_738 (O_738,N_43812,N_41035);
nand UO_739 (O_739,N_44537,N_44260);
and UO_740 (O_740,N_49370,N_44108);
nand UO_741 (O_741,N_43675,N_47166);
and UO_742 (O_742,N_44212,N_44570);
or UO_743 (O_743,N_48518,N_40584);
xnor UO_744 (O_744,N_46747,N_48694);
nor UO_745 (O_745,N_48865,N_49073);
or UO_746 (O_746,N_47406,N_44366);
xor UO_747 (O_747,N_46042,N_47691);
nor UO_748 (O_748,N_43938,N_41840);
and UO_749 (O_749,N_47461,N_46071);
nor UO_750 (O_750,N_48530,N_41403);
or UO_751 (O_751,N_49502,N_48827);
nand UO_752 (O_752,N_45692,N_44046);
nand UO_753 (O_753,N_43670,N_45591);
nand UO_754 (O_754,N_41451,N_46506);
nand UO_755 (O_755,N_49022,N_41511);
or UO_756 (O_756,N_49699,N_48710);
nor UO_757 (O_757,N_40853,N_40968);
or UO_758 (O_758,N_42197,N_47846);
or UO_759 (O_759,N_44750,N_48733);
or UO_760 (O_760,N_48275,N_44527);
nor UO_761 (O_761,N_42604,N_47101);
nor UO_762 (O_762,N_48615,N_41944);
or UO_763 (O_763,N_47261,N_49263);
nand UO_764 (O_764,N_42771,N_46265);
or UO_765 (O_765,N_48805,N_49179);
and UO_766 (O_766,N_46836,N_49375);
xnor UO_767 (O_767,N_42900,N_44257);
nor UO_768 (O_768,N_43664,N_46234);
and UO_769 (O_769,N_43824,N_41814);
or UO_770 (O_770,N_47331,N_43114);
xnor UO_771 (O_771,N_45022,N_43530);
and UO_772 (O_772,N_43467,N_41367);
nand UO_773 (O_773,N_43724,N_43466);
nand UO_774 (O_774,N_42211,N_49270);
nor UO_775 (O_775,N_40905,N_43542);
and UO_776 (O_776,N_47372,N_43288);
or UO_777 (O_777,N_41006,N_49330);
nor UO_778 (O_778,N_48617,N_48188);
and UO_779 (O_779,N_49295,N_41282);
or UO_780 (O_780,N_48010,N_49662);
or UO_781 (O_781,N_44847,N_44126);
and UO_782 (O_782,N_41121,N_45103);
xor UO_783 (O_783,N_46686,N_43298);
or UO_784 (O_784,N_42688,N_44560);
and UO_785 (O_785,N_46746,N_43957);
and UO_786 (O_786,N_44208,N_43478);
xnor UO_787 (O_787,N_45886,N_45754);
and UO_788 (O_788,N_43042,N_42003);
or UO_789 (O_789,N_47085,N_49958);
or UO_790 (O_790,N_43660,N_44962);
xor UO_791 (O_791,N_45446,N_42728);
nor UO_792 (O_792,N_42672,N_49701);
and UO_793 (O_793,N_43100,N_47636);
and UO_794 (O_794,N_40435,N_47996);
nand UO_795 (O_795,N_46437,N_46027);
nor UO_796 (O_796,N_43772,N_46709);
or UO_797 (O_797,N_48034,N_44326);
xnor UO_798 (O_798,N_44671,N_40409);
nor UO_799 (O_799,N_43700,N_43590);
nor UO_800 (O_800,N_49980,N_47433);
or UO_801 (O_801,N_42058,N_44608);
nand UO_802 (O_802,N_48109,N_45087);
nor UO_803 (O_803,N_48089,N_49067);
nand UO_804 (O_804,N_43594,N_49019);
nand UO_805 (O_805,N_44105,N_45524);
nand UO_806 (O_806,N_47723,N_48102);
xnor UO_807 (O_807,N_41066,N_43547);
and UO_808 (O_808,N_44120,N_45125);
or UO_809 (O_809,N_46005,N_42381);
and UO_810 (O_810,N_47225,N_46418);
xor UO_811 (O_811,N_43554,N_41461);
xor UO_812 (O_812,N_44863,N_42240);
xor UO_813 (O_813,N_42416,N_42545);
xor UO_814 (O_814,N_42451,N_47391);
xnor UO_815 (O_815,N_42077,N_48871);
xor UO_816 (O_816,N_48930,N_48421);
xnor UO_817 (O_817,N_40659,N_48517);
xnor UO_818 (O_818,N_43521,N_42818);
or UO_819 (O_819,N_49731,N_43852);
xor UO_820 (O_820,N_44141,N_49095);
nand UO_821 (O_821,N_43497,N_44416);
xnor UO_822 (O_822,N_47522,N_49306);
and UO_823 (O_823,N_40154,N_41526);
and UO_824 (O_824,N_44357,N_45200);
or UO_825 (O_825,N_49930,N_41956);
or UO_826 (O_826,N_48189,N_41504);
nand UO_827 (O_827,N_47739,N_46753);
or UO_828 (O_828,N_41111,N_48580);
or UO_829 (O_829,N_48566,N_47469);
or UO_830 (O_830,N_40638,N_45709);
or UO_831 (O_831,N_47193,N_48901);
nand UO_832 (O_832,N_45632,N_43814);
and UO_833 (O_833,N_46384,N_44793);
and UO_834 (O_834,N_49618,N_40510);
xnor UO_835 (O_835,N_46407,N_47053);
nor UO_836 (O_836,N_44842,N_46375);
nand UO_837 (O_837,N_44846,N_44484);
xor UO_838 (O_838,N_44539,N_48008);
or UO_839 (O_839,N_45926,N_46558);
nor UO_840 (O_840,N_46183,N_43759);
nand UO_841 (O_841,N_48822,N_49308);
and UO_842 (O_842,N_40123,N_42431);
nor UO_843 (O_843,N_43359,N_49816);
nor UO_844 (O_844,N_41079,N_40896);
or UO_845 (O_845,N_45530,N_48231);
nand UO_846 (O_846,N_46668,N_47233);
xnor UO_847 (O_847,N_41373,N_49208);
nor UO_848 (O_848,N_40428,N_40239);
and UO_849 (O_849,N_42119,N_40678);
xnor UO_850 (O_850,N_49425,N_41546);
xnor UO_851 (O_851,N_42760,N_43869);
nor UO_852 (O_852,N_47248,N_44633);
and UO_853 (O_853,N_46831,N_43750);
or UO_854 (O_854,N_40289,N_40244);
nand UO_855 (O_855,N_48233,N_46999);
nand UO_856 (O_856,N_41315,N_49438);
xnor UO_857 (O_857,N_49586,N_47518);
and UO_858 (O_858,N_40399,N_44093);
nor UO_859 (O_859,N_47922,N_42359);
nand UO_860 (O_860,N_44804,N_40166);
xor UO_861 (O_861,N_41107,N_47379);
nand UO_862 (O_862,N_42147,N_46902);
nor UO_863 (O_863,N_43508,N_41914);
nand UO_864 (O_864,N_48129,N_41340);
nor UO_865 (O_865,N_47712,N_41947);
xnor UO_866 (O_866,N_40118,N_44391);
and UO_867 (O_867,N_43715,N_40674);
xnor UO_868 (O_868,N_40778,N_45895);
and UO_869 (O_869,N_48073,N_46434);
xnor UO_870 (O_870,N_48293,N_45903);
nand UO_871 (O_871,N_41210,N_40193);
nor UO_872 (O_872,N_47673,N_40926);
nand UO_873 (O_873,N_47910,N_41422);
and UO_874 (O_874,N_46424,N_43601);
xnor UO_875 (O_875,N_44421,N_46354);
and UO_876 (O_876,N_48962,N_46337);
or UO_877 (O_877,N_45367,N_40681);
and UO_878 (O_878,N_49074,N_44315);
nor UO_879 (O_879,N_46115,N_41639);
and UO_880 (O_880,N_49688,N_47495);
or UO_881 (O_881,N_46485,N_40569);
nor UO_882 (O_882,N_44364,N_47785);
nand UO_883 (O_883,N_49897,N_43413);
nand UO_884 (O_884,N_46788,N_46629);
or UO_885 (O_885,N_45465,N_45961);
nand UO_886 (O_886,N_45711,N_49357);
xnor UO_887 (O_887,N_43704,N_44531);
and UO_888 (O_888,N_41420,N_48981);
nor UO_889 (O_889,N_46712,N_41690);
or UO_890 (O_890,N_46089,N_43344);
xor UO_891 (O_891,N_46116,N_43693);
xor UO_892 (O_892,N_49475,N_49334);
nor UO_893 (O_893,N_45247,N_49950);
and UO_894 (O_894,N_43878,N_48181);
and UO_895 (O_895,N_43963,N_46572);
and UO_896 (O_896,N_45132,N_41571);
and UO_897 (O_897,N_43904,N_46995);
nor UO_898 (O_898,N_49969,N_46994);
xnor UO_899 (O_899,N_47480,N_42478);
or UO_900 (O_900,N_46744,N_47387);
and UO_901 (O_901,N_47564,N_40670);
nor UO_902 (O_902,N_48815,N_43736);
nor UO_903 (O_903,N_49157,N_44146);
and UO_904 (O_904,N_42944,N_42247);
and UO_905 (O_905,N_40658,N_49968);
or UO_906 (O_906,N_43658,N_46376);
and UO_907 (O_907,N_48087,N_48523);
nor UO_908 (O_908,N_46363,N_41834);
and UO_909 (O_909,N_43151,N_41793);
nor UO_910 (O_910,N_46294,N_44369);
and UO_911 (O_911,N_43430,N_43323);
and UO_912 (O_912,N_43334,N_45985);
nor UO_913 (O_913,N_40660,N_42670);
xnor UO_914 (O_914,N_48037,N_47198);
nor UO_915 (O_915,N_49011,N_43244);
xor UO_916 (O_916,N_48056,N_47930);
or UO_917 (O_917,N_46455,N_40292);
or UO_918 (O_918,N_45532,N_49151);
and UO_919 (O_919,N_44885,N_41090);
or UO_920 (O_920,N_49345,N_46167);
nand UO_921 (O_921,N_49734,N_41572);
nand UO_922 (O_922,N_49654,N_42820);
nor UO_923 (O_923,N_40232,N_42046);
and UO_924 (O_924,N_41408,N_46876);
nand UO_925 (O_925,N_45254,N_48497);
and UO_926 (O_926,N_45156,N_41694);
nand UO_927 (O_927,N_40611,N_41875);
or UO_928 (O_928,N_43388,N_49170);
and UO_929 (O_929,N_49486,N_48447);
or UO_930 (O_930,N_45649,N_49954);
xor UO_931 (O_931,N_48768,N_46942);
nand UO_932 (O_932,N_44744,N_40348);
nand UO_933 (O_933,N_41337,N_44641);
nor UO_934 (O_934,N_43695,N_43548);
xor UO_935 (O_935,N_44884,N_44222);
nor UO_936 (O_936,N_46817,N_45438);
or UO_937 (O_937,N_46276,N_43770);
nor UO_938 (O_938,N_48500,N_45851);
xor UO_939 (O_939,N_47508,N_42703);
nor UO_940 (O_940,N_47294,N_41417);
and UO_941 (O_941,N_42880,N_48394);
and UO_942 (O_942,N_40075,N_46628);
xor UO_943 (O_943,N_46049,N_40643);
nor UO_944 (O_944,N_41281,N_44721);
nand UO_945 (O_945,N_42323,N_49657);
nor UO_946 (O_946,N_41659,N_46945);
nor UO_947 (O_947,N_49055,N_48206);
and UO_948 (O_948,N_43074,N_41475);
nor UO_949 (O_949,N_45422,N_46052);
nand UO_950 (O_950,N_41064,N_43849);
nor UO_951 (O_951,N_48232,N_46201);
and UO_952 (O_952,N_46445,N_46379);
nand UO_953 (O_953,N_44040,N_42653);
nor UO_954 (O_954,N_46190,N_47009);
and UO_955 (O_955,N_49562,N_44809);
nor UO_956 (O_956,N_48672,N_45854);
nor UO_957 (O_957,N_40215,N_41807);
nor UO_958 (O_958,N_40065,N_48933);
nand UO_959 (O_959,N_47800,N_43821);
xor UO_960 (O_960,N_41945,N_49283);
nor UO_961 (O_961,N_43062,N_42685);
or UO_962 (O_962,N_47897,N_44117);
xnor UO_963 (O_963,N_40762,N_48055);
nand UO_964 (O_964,N_41262,N_40642);
xor UO_965 (O_965,N_45964,N_44835);
nor UO_966 (O_966,N_44653,N_43398);
xnor UO_967 (O_967,N_49831,N_44271);
xnor UO_968 (O_968,N_45117,N_42309);
nand UO_969 (O_969,N_44716,N_42056);
nor UO_970 (O_970,N_46887,N_44559);
nor UO_971 (O_971,N_43150,N_44614);
and UO_972 (O_972,N_48577,N_47076);
and UO_973 (O_973,N_41757,N_45693);
and UO_974 (O_974,N_46905,N_46390);
nand UO_975 (O_975,N_45384,N_49733);
and UO_976 (O_976,N_42808,N_44933);
or UO_977 (O_977,N_49963,N_43005);
nor UO_978 (O_978,N_49600,N_48741);
nor UO_979 (O_979,N_49437,N_44887);
nand UO_980 (O_980,N_42626,N_49920);
and UO_981 (O_981,N_48133,N_43489);
nor UO_982 (O_982,N_43742,N_42991);
or UO_983 (O_983,N_47828,N_47488);
nor UO_984 (O_984,N_41099,N_41274);
nand UO_985 (O_985,N_47905,N_41656);
nand UO_986 (O_986,N_45904,N_44830);
nand UO_987 (O_987,N_45588,N_42207);
nor UO_988 (O_988,N_49527,N_46495);
xnor UO_989 (O_989,N_48996,N_49081);
or UO_990 (O_990,N_44490,N_48460);
nand UO_991 (O_991,N_41132,N_47951);
nor UO_992 (O_992,N_44695,N_41542);
nor UO_993 (O_993,N_42432,N_40446);
xnor UO_994 (O_994,N_41181,N_42341);
nand UO_995 (O_995,N_47928,N_49979);
or UO_996 (O_996,N_43363,N_43031);
xnor UO_997 (O_997,N_41191,N_40873);
xor UO_998 (O_998,N_49902,N_43494);
xor UO_999 (O_999,N_41967,N_41794);
nand UO_1000 (O_1000,N_43435,N_46185);
nand UO_1001 (O_1001,N_40240,N_45452);
xor UO_1002 (O_1002,N_46378,N_41002);
and UO_1003 (O_1003,N_48032,N_46764);
nor UO_1004 (O_1004,N_40863,N_43372);
or UO_1005 (O_1005,N_45244,N_41555);
xnor UO_1006 (O_1006,N_48219,N_44806);
nor UO_1007 (O_1007,N_44964,N_41606);
xnor UO_1008 (O_1008,N_42669,N_48883);
nand UO_1009 (O_1009,N_47160,N_46848);
and UO_1010 (O_1010,N_44917,N_44150);
nand UO_1011 (O_1011,N_42441,N_47462);
or UO_1012 (O_1012,N_47871,N_43202);
xnor UO_1013 (O_1013,N_47157,N_40983);
xnor UO_1014 (O_1014,N_45107,N_41866);
nor UO_1015 (O_1015,N_40343,N_43971);
and UO_1016 (O_1016,N_48628,N_41046);
and UO_1017 (O_1017,N_42713,N_41593);
xor UO_1018 (O_1018,N_48665,N_40718);
nand UO_1019 (O_1019,N_47232,N_40266);
xnor UO_1020 (O_1020,N_41909,N_48174);
and UO_1021 (O_1021,N_44303,N_41869);
xor UO_1022 (O_1022,N_42564,N_44800);
and UO_1023 (O_1023,N_49229,N_40157);
nor UO_1024 (O_1024,N_42368,N_41992);
or UO_1025 (O_1025,N_40475,N_48760);
nor UO_1026 (O_1026,N_46317,N_48325);
xor UO_1027 (O_1027,N_40830,N_45195);
xnor UO_1028 (O_1028,N_44680,N_49429);
and UO_1029 (O_1029,N_44081,N_45750);
or UO_1030 (O_1030,N_43761,N_40697);
nand UO_1031 (O_1031,N_46031,N_46552);
and UO_1032 (O_1032,N_40451,N_48504);
or UO_1033 (O_1033,N_43688,N_42811);
nand UO_1034 (O_1034,N_45521,N_48627);
nor UO_1035 (O_1035,N_42496,N_48926);
and UO_1036 (O_1036,N_48310,N_49399);
nor UO_1037 (O_1037,N_47156,N_49402);
xnor UO_1038 (O_1038,N_40652,N_46498);
or UO_1039 (O_1039,N_48524,N_45175);
and UO_1040 (O_1040,N_47060,N_46515);
or UO_1041 (O_1041,N_48048,N_41987);
nor UO_1042 (O_1042,N_40407,N_46719);
nor UO_1043 (O_1043,N_43606,N_45762);
xnor UO_1044 (O_1044,N_44067,N_43248);
nor UO_1045 (O_1045,N_47619,N_48940);
or UO_1046 (O_1046,N_40589,N_44714);
and UO_1047 (O_1047,N_45400,N_46417);
or UO_1048 (O_1048,N_41774,N_46114);
xnor UO_1049 (O_1049,N_45663,N_41578);
or UO_1050 (O_1050,N_42954,N_42854);
and UO_1051 (O_1051,N_46451,N_47895);
xnor UO_1052 (O_1052,N_48878,N_49793);
and UO_1053 (O_1053,N_45219,N_42489);
nor UO_1054 (O_1054,N_44095,N_46514);
nand UO_1055 (O_1055,N_42609,N_44160);
and UO_1056 (O_1056,N_47609,N_47487);
and UO_1057 (O_1057,N_42577,N_44690);
and UO_1058 (O_1058,N_40007,N_47375);
xnor UO_1059 (O_1059,N_48746,N_41225);
nor UO_1060 (O_1060,N_40380,N_49262);
nand UO_1061 (O_1061,N_42719,N_48506);
nor UO_1062 (O_1062,N_42034,N_47290);
or UO_1063 (O_1063,N_48105,N_41900);
xnor UO_1064 (O_1064,N_45201,N_45366);
nor UO_1065 (O_1065,N_44542,N_40704);
nor UO_1066 (O_1066,N_46778,N_42514);
xor UO_1067 (O_1067,N_49641,N_40488);
nor UO_1068 (O_1068,N_45575,N_40561);
and UO_1069 (O_1069,N_47291,N_45414);
and UO_1070 (O_1070,N_44055,N_45602);
nor UO_1071 (O_1071,N_41005,N_44592);
and UO_1072 (O_1072,N_44226,N_45823);
xnor UO_1073 (O_1073,N_46274,N_46484);
xnor UO_1074 (O_1074,N_44123,N_47416);
xnor UO_1075 (O_1075,N_42435,N_40387);
and UO_1076 (O_1076,N_43785,N_49971);
nand UO_1077 (O_1077,N_42868,N_43894);
and UO_1078 (O_1078,N_40335,N_49707);
or UO_1079 (O_1079,N_48493,N_41412);
nand UO_1080 (O_1080,N_44023,N_46132);
and UO_1081 (O_1081,N_42861,N_48870);
and UO_1082 (O_1082,N_44934,N_48107);
nor UO_1083 (O_1083,N_43906,N_46864);
nor UO_1084 (O_1084,N_44460,N_49355);
and UO_1085 (O_1085,N_42007,N_49238);
nor UO_1086 (O_1086,N_47244,N_43165);
nand UO_1087 (O_1087,N_49602,N_41561);
nor UO_1088 (O_1088,N_46614,N_44547);
or UO_1089 (O_1089,N_49324,N_46743);
and UO_1090 (O_1090,N_44335,N_49195);
and UO_1091 (O_1091,N_40129,N_40806);
and UO_1092 (O_1092,N_47466,N_49678);
xor UO_1093 (O_1093,N_41195,N_41297);
and UO_1094 (O_1094,N_40425,N_42522);
or UO_1095 (O_1095,N_46544,N_41272);
nor UO_1096 (O_1096,N_46765,N_44269);
xor UO_1097 (O_1097,N_41284,N_45417);
nor UO_1098 (O_1098,N_41934,N_47849);
xor UO_1099 (O_1099,N_46918,N_48532);
nor UO_1100 (O_1100,N_43474,N_49610);
or UO_1101 (O_1101,N_47535,N_45730);
xnor UO_1102 (O_1102,N_42486,N_41650);
and UO_1103 (O_1103,N_45953,N_40174);
xor UO_1104 (O_1104,N_41457,N_42826);
and UO_1105 (O_1105,N_41395,N_49145);
and UO_1106 (O_1106,N_40882,N_44589);
nand UO_1107 (O_1107,N_46585,N_46896);
or UO_1108 (O_1108,N_43850,N_44501);
nor UO_1109 (O_1109,N_48005,N_40067);
and UO_1110 (O_1110,N_46604,N_40645);
or UO_1111 (O_1111,N_44365,N_47413);
or UO_1112 (O_1112,N_49696,N_42285);
xor UO_1113 (O_1113,N_43387,N_48637);
nand UO_1114 (O_1114,N_42047,N_48205);
nand UO_1115 (O_1115,N_44580,N_49131);
nand UO_1116 (O_1116,N_44347,N_44892);
nand UO_1117 (O_1117,N_45457,N_49478);
and UO_1118 (O_1118,N_49427,N_48572);
nand UO_1119 (O_1119,N_40803,N_48038);
xnor UO_1120 (O_1120,N_41288,N_48337);
nand UO_1121 (O_1121,N_46875,N_49634);
or UO_1122 (O_1122,N_48722,N_40941);
xnor UO_1123 (O_1123,N_45576,N_45413);
or UO_1124 (O_1124,N_49191,N_49363);
and UO_1125 (O_1125,N_40613,N_43118);
xor UO_1126 (O_1126,N_40060,N_48648);
xor UO_1127 (O_1127,N_43806,N_47990);
nor UO_1128 (O_1128,N_45431,N_41617);
xor UO_1129 (O_1129,N_47585,N_43106);
and UO_1130 (O_1130,N_41813,N_43246);
or UO_1131 (O_1131,N_43579,N_45309);
xnor UO_1132 (O_1132,N_44883,N_44660);
nand UO_1133 (O_1133,N_46651,N_49153);
nor UO_1134 (O_1134,N_44951,N_46399);
nand UO_1135 (O_1135,N_43504,N_48074);
nand UO_1136 (O_1136,N_44620,N_49057);
xnor UO_1137 (O_1137,N_41065,N_44949);
or UO_1138 (O_1138,N_49362,N_44164);
and UO_1139 (O_1139,N_41463,N_40827);
and UO_1140 (O_1140,N_40117,N_46745);
xnor UO_1141 (O_1141,N_46607,N_49335);
nor UO_1142 (O_1142,N_49526,N_47000);
xnor UO_1143 (O_1143,N_43708,N_44703);
nand UO_1144 (O_1144,N_46768,N_46584);
xor UO_1145 (O_1145,N_42725,N_49866);
xnor UO_1146 (O_1146,N_46837,N_40394);
or UO_1147 (O_1147,N_45746,N_46619);
nor UO_1148 (O_1148,N_49434,N_43718);
nor UO_1149 (O_1149,N_49448,N_48646);
and UO_1150 (O_1150,N_44900,N_42002);
xor UO_1151 (O_1151,N_41119,N_42469);
nor UO_1152 (O_1152,N_41037,N_44089);
xor UO_1153 (O_1153,N_48131,N_40836);
or UO_1154 (O_1154,N_47190,N_41001);
and UO_1155 (O_1155,N_47970,N_43706);
nand UO_1156 (O_1156,N_45593,N_41019);
xor UO_1157 (O_1157,N_46187,N_41470);
xor UO_1158 (O_1158,N_43121,N_46625);
nor UO_1159 (O_1159,N_43146,N_41220);
nor UO_1160 (O_1160,N_42801,N_41397);
xnor UO_1161 (O_1161,N_43360,N_48857);
nor UO_1162 (O_1162,N_41686,N_41235);
or UO_1163 (O_1163,N_45741,N_49418);
and UO_1164 (O_1164,N_40306,N_42891);
and UO_1165 (O_1165,N_41486,N_44676);
and UO_1166 (O_1166,N_49547,N_48541);
and UO_1167 (O_1167,N_47877,N_45445);
and UO_1168 (O_1168,N_49198,N_42016);
nand UO_1169 (O_1169,N_41109,N_40149);
xor UO_1170 (O_1170,N_43557,N_47603);
nor UO_1171 (O_1171,N_46809,N_40175);
nand UO_1172 (O_1172,N_46538,N_48723);
xnor UO_1173 (O_1173,N_42184,N_49745);
xor UO_1174 (O_1174,N_40991,N_41088);
nor UO_1175 (O_1175,N_45491,N_43661);
xor UO_1176 (O_1176,N_48252,N_41445);
or UO_1177 (O_1177,N_49384,N_45261);
and UO_1178 (O_1178,N_43251,N_44128);
and UO_1179 (O_1179,N_48949,N_43519);
nor UO_1180 (O_1180,N_40242,N_45797);
and UO_1181 (O_1181,N_42296,N_48684);
and UO_1182 (O_1182,N_44602,N_47345);
nand UO_1183 (O_1183,N_49141,N_41543);
and UO_1184 (O_1184,N_45586,N_42245);
xnor UO_1185 (O_1185,N_45756,N_46237);
and UO_1186 (O_1186,N_44229,N_44248);
nand UO_1187 (O_1187,N_43636,N_42454);
or UO_1188 (O_1188,N_42425,N_45830);
or UO_1189 (O_1189,N_49365,N_41854);
nand UO_1190 (O_1190,N_41033,N_44008);
xor UO_1191 (O_1191,N_47090,N_45859);
or UO_1192 (O_1192,N_49935,N_44638);
or UO_1193 (O_1193,N_44174,N_40041);
or UO_1194 (O_1194,N_41112,N_45236);
xnor UO_1195 (O_1195,N_47216,N_43488);
or UO_1196 (O_1196,N_41724,N_44899);
xor UO_1197 (O_1197,N_44825,N_42562);
nor UO_1198 (O_1198,N_48141,N_47982);
nand UO_1199 (O_1199,N_45749,N_45657);
nor UO_1200 (O_1200,N_44037,N_47389);
nand UO_1201 (O_1201,N_42039,N_42423);
and UO_1202 (O_1202,N_40686,N_46592);
nand UO_1203 (O_1203,N_42539,N_48365);
or UO_1204 (O_1204,N_47320,N_42836);
nand UO_1205 (O_1205,N_40241,N_44118);
nor UO_1206 (O_1206,N_49085,N_41665);
nor UO_1207 (O_1207,N_48576,N_44057);
and UO_1208 (O_1208,N_48084,N_48763);
xnor UO_1209 (O_1209,N_47403,N_45871);
nand UO_1210 (O_1210,N_43159,N_49498);
and UO_1211 (O_1211,N_44413,N_43702);
and UO_1212 (O_1212,N_43716,N_46330);
nor UO_1213 (O_1213,N_47822,N_44470);
and UO_1214 (O_1214,N_48216,N_47154);
nand UO_1215 (O_1215,N_44731,N_46015);
nand UO_1216 (O_1216,N_41820,N_44873);
xor UO_1217 (O_1217,N_48818,N_40954);
and UO_1218 (O_1218,N_46970,N_42193);
or UO_1219 (O_1219,N_46146,N_48103);
nor UO_1220 (O_1220,N_41115,N_42169);
nand UO_1221 (O_1221,N_43958,N_48586);
and UO_1222 (O_1222,N_45502,N_41353);
and UO_1223 (O_1223,N_46520,N_45621);
and UO_1224 (O_1224,N_41244,N_45300);
nand UO_1225 (O_1225,N_46404,N_43607);
nor UO_1226 (O_1226,N_47999,N_43045);
nor UO_1227 (O_1227,N_45004,N_45169);
nor UO_1228 (O_1228,N_44340,N_41990);
and UO_1229 (O_1229,N_40838,N_44906);
nor UO_1230 (O_1230,N_48448,N_41094);
nand UO_1231 (O_1231,N_41169,N_46787);
xor UO_1232 (O_1232,N_44290,N_45644);
nand UO_1233 (O_1233,N_44133,N_44214);
nand UO_1234 (O_1234,N_40595,N_44264);
nand UO_1235 (O_1235,N_44718,N_48071);
nand UO_1236 (O_1236,N_46486,N_45921);
or UO_1237 (O_1237,N_45262,N_44789);
or UO_1238 (O_1238,N_45890,N_44759);
xor UO_1239 (O_1239,N_45216,N_49408);
nor UO_1240 (O_1240,N_40464,N_49543);
xnor UO_1241 (O_1241,N_47066,N_42544);
and UO_1242 (O_1242,N_47031,N_45580);
xnor UO_1243 (O_1243,N_42084,N_41441);
and UO_1244 (O_1244,N_48377,N_42223);
xnor UO_1245 (O_1245,N_42985,N_45791);
and UO_1246 (O_1246,N_46195,N_42297);
or UO_1247 (O_1247,N_42351,N_40236);
xnor UO_1248 (O_1248,N_44923,N_41928);
and UO_1249 (O_1249,N_45708,N_42840);
nand UO_1250 (O_1250,N_43087,N_44544);
or UO_1251 (O_1251,N_47362,N_46706);
and UO_1252 (O_1252,N_48958,N_43104);
nor UO_1253 (O_1253,N_44420,N_47384);
and UO_1254 (O_1254,N_43192,N_41785);
xor UO_1255 (O_1255,N_48386,N_49937);
or UO_1256 (O_1256,N_40690,N_46748);
or UO_1257 (O_1257,N_46104,N_48178);
or UO_1258 (O_1258,N_46781,N_46248);
xor UO_1259 (O_1259,N_44148,N_47903);
and UO_1260 (O_1260,N_47786,N_47620);
nand UO_1261 (O_1261,N_40299,N_44634);
nand UO_1262 (O_1262,N_43748,N_46064);
nand UO_1263 (O_1263,N_43148,N_48707);
nor UO_1264 (O_1264,N_46355,N_41371);
nor UO_1265 (O_1265,N_46145,N_40794);
or UO_1266 (O_1266,N_46079,N_41695);
nand UO_1267 (O_1267,N_48110,N_40083);
or UO_1268 (O_1268,N_42585,N_44162);
nor UO_1269 (O_1269,N_42230,N_48033);
and UO_1270 (O_1270,N_48370,N_43810);
xor UO_1271 (O_1271,N_41713,N_40829);
nand UO_1272 (O_1272,N_48101,N_41754);
xnor UO_1273 (O_1273,N_49579,N_46914);
nand UO_1274 (O_1274,N_47388,N_49578);
and UO_1275 (O_1275,N_48329,N_43993);
nand UO_1276 (O_1276,N_46825,N_46783);
and UO_1277 (O_1277,N_47801,N_46285);
and UO_1278 (O_1278,N_42578,N_45183);
nand UO_1279 (O_1279,N_49995,N_43578);
xnor UO_1280 (O_1280,N_49396,N_46860);
nor UO_1281 (O_1281,N_46440,N_48956);
xor UO_1282 (O_1282,N_45289,N_47167);
xor UO_1283 (O_1283,N_41716,N_46525);
xnor UO_1284 (O_1284,N_49440,N_46227);
nand UO_1285 (O_1285,N_45010,N_45769);
nor UO_1286 (O_1286,N_45675,N_43346);
or UO_1287 (O_1287,N_43720,N_46840);
and UO_1288 (O_1288,N_45767,N_42320);
xor UO_1289 (O_1289,N_49274,N_45019);
nor UO_1290 (O_1290,N_48452,N_43905);
and UO_1291 (O_1291,N_42646,N_44296);
nor UO_1292 (O_1292,N_48040,N_43191);
nand UO_1293 (O_1293,N_47744,N_49140);
xnor UO_1294 (O_1294,N_44234,N_49687);
and UO_1295 (O_1295,N_48355,N_42879);
and UO_1296 (O_1296,N_45569,N_46123);
and UO_1297 (O_1297,N_47670,N_40532);
nand UO_1298 (O_1298,N_44217,N_48081);
and UO_1299 (O_1299,N_47686,N_44477);
and UO_1300 (O_1300,N_45064,N_42608);
nand UO_1301 (O_1301,N_44262,N_44280);
nor UO_1302 (O_1302,N_47103,N_41036);
nor UO_1303 (O_1303,N_49123,N_44574);
xor UO_1304 (O_1304,N_40766,N_47797);
nor UO_1305 (O_1305,N_48659,N_47317);
or UO_1306 (O_1306,N_46810,N_48538);
nand UO_1307 (O_1307,N_40671,N_43766);
or UO_1308 (O_1308,N_40503,N_47328);
or UO_1309 (O_1309,N_43325,N_44805);
nand UO_1310 (O_1310,N_43291,N_49557);
xor UO_1311 (O_1311,N_42557,N_41862);
and UO_1312 (O_1312,N_41172,N_42470);
nor UO_1313 (O_1313,N_47113,N_49645);
nand UO_1314 (O_1314,N_47419,N_46206);
and UO_1315 (O_1315,N_47667,N_46416);
or UO_1316 (O_1316,N_48455,N_49101);
xor UO_1317 (O_1317,N_46018,N_40864);
and UO_1318 (O_1318,N_49966,N_49317);
or UO_1319 (O_1319,N_49441,N_42092);
or UO_1320 (O_1320,N_42071,N_47222);
and UO_1321 (O_1321,N_45592,N_46823);
xnor UO_1322 (O_1322,N_47411,N_40440);
or UO_1323 (O_1323,N_44874,N_46926);
nor UO_1324 (O_1324,N_48135,N_41943);
xnor UO_1325 (O_1325,N_43412,N_42534);
nor UO_1326 (O_1326,N_46724,N_44534);
nor UO_1327 (O_1327,N_44864,N_40861);
and UO_1328 (O_1328,N_46939,N_48661);
nand UO_1329 (O_1329,N_42334,N_46782);
or UO_1330 (O_1330,N_42866,N_42942);
xnor UO_1331 (O_1331,N_44861,N_41351);
xnor UO_1332 (O_1332,N_45775,N_43310);
xnor UO_1333 (O_1333,N_45130,N_42307);
and UO_1334 (O_1334,N_47297,N_43535);
or UO_1335 (O_1335,N_44895,N_49205);
or UO_1336 (O_1336,N_44798,N_48059);
xnor UO_1337 (O_1337,N_46689,N_48801);
xnor UO_1338 (O_1338,N_49444,N_43865);
nor UO_1339 (O_1339,N_49998,N_40151);
nor UO_1340 (O_1340,N_45222,N_41860);
nand UO_1341 (O_1341,N_46900,N_41101);
nor UO_1342 (O_1342,N_49679,N_44860);
nor UO_1343 (O_1343,N_46345,N_45522);
xor UO_1344 (O_1344,N_46477,N_48168);
nand UO_1345 (O_1345,N_43854,N_48952);
xor UO_1346 (O_1346,N_46381,N_46611);
nand UO_1347 (O_1347,N_47363,N_43211);
xnor UO_1348 (O_1348,N_40739,N_40964);
nor UO_1349 (O_1349,N_44596,N_48378);
or UO_1350 (O_1350,N_44070,N_41537);
nand UO_1351 (O_1351,N_47126,N_45469);
or UO_1352 (O_1352,N_42845,N_40025);
or UO_1353 (O_1353,N_40565,N_46691);
nand UO_1354 (O_1354,N_49594,N_48132);
or UO_1355 (O_1355,N_43925,N_48507);
and UO_1356 (O_1356,N_42291,N_45124);
xor UO_1357 (O_1357,N_47175,N_41205);
xor UO_1358 (O_1358,N_42000,N_47035);
and UO_1359 (O_1359,N_42774,N_47855);
xnor UO_1360 (O_1360,N_43825,N_48464);
nor UO_1361 (O_1361,N_41502,N_49508);
nand UO_1362 (O_1362,N_43275,N_43366);
xnor UO_1363 (O_1363,N_41851,N_49267);
or UO_1364 (O_1364,N_46149,N_43928);
nor UO_1365 (O_1365,N_49563,N_40998);
nand UO_1366 (O_1366,N_46083,N_47378);
or UO_1367 (O_1367,N_42839,N_40026);
xor UO_1368 (O_1368,N_43563,N_43321);
and UO_1369 (O_1369,N_42376,N_47886);
or UO_1370 (O_1370,N_46197,N_45231);
xor UO_1371 (O_1371,N_41485,N_44064);
xnor UO_1372 (O_1372,N_46003,N_48914);
nor UO_1373 (O_1373,N_43102,N_41658);
or UO_1374 (O_1374,N_48593,N_48457);
nand UO_1375 (O_1375,N_43424,N_48338);
or UO_1376 (O_1376,N_46032,N_40689);
or UO_1377 (O_1377,N_48754,N_41582);
or UO_1378 (O_1378,N_43115,N_48850);
xnor UO_1379 (O_1379,N_45635,N_48371);
nand UO_1380 (O_1380,N_40319,N_45722);
and UO_1381 (O_1381,N_46372,N_48191);
xnor UO_1382 (O_1382,N_49524,N_40685);
and UO_1383 (O_1383,N_44872,N_47463);
nand UO_1384 (O_1384,N_41549,N_41303);
nand UO_1385 (O_1385,N_46699,N_42300);
xor UO_1386 (O_1386,N_43999,N_47197);
nand UO_1387 (O_1387,N_42152,N_42217);
or UO_1388 (O_1388,N_47178,N_46491);
nand UO_1389 (O_1389,N_49635,N_44787);
nand UO_1390 (O_1390,N_42846,N_48066);
xnor UO_1391 (O_1391,N_43616,N_49821);
nand UO_1392 (O_1392,N_49631,N_44733);
and UO_1393 (O_1393,N_46352,N_42502);
or UO_1394 (O_1394,N_43247,N_42362);
xnor UO_1395 (O_1395,N_42175,N_42889);
nand UO_1396 (O_1396,N_46562,N_45344);
nand UO_1397 (O_1397,N_47049,N_48467);
xnor UO_1398 (O_1398,N_40080,N_42159);
xnor UO_1399 (O_1399,N_45112,N_44409);
or UO_1400 (O_1400,N_45612,N_42762);
nor UO_1401 (O_1401,N_41556,N_48951);
and UO_1402 (O_1402,N_40411,N_47438);
and UO_1403 (O_1403,N_41024,N_47549);
or UO_1404 (O_1404,N_42998,N_48255);
and UO_1405 (O_1405,N_45707,N_40664);
nand UO_1406 (O_1406,N_44330,N_42692);
and UO_1407 (O_1407,N_41263,N_45059);
nand UO_1408 (O_1408,N_43980,N_40793);
nor UO_1409 (O_1409,N_48347,N_48462);
or UO_1410 (O_1410,N_40598,N_43515);
and UO_1411 (O_1411,N_48241,N_48828);
xnor UO_1412 (O_1412,N_46347,N_48227);
nor UO_1413 (O_1413,N_43959,N_45609);
xnor UO_1414 (O_1414,N_43886,N_48626);
or UO_1415 (O_1415,N_49989,N_49368);
nor UO_1416 (O_1416,N_47376,N_46016);
nand UO_1417 (O_1417,N_48512,N_48363);
or UO_1418 (O_1418,N_43564,N_45391);
and UO_1419 (O_1419,N_44513,N_48042);
and UO_1420 (O_1420,N_47408,N_43409);
nand UO_1421 (O_1421,N_45865,N_45717);
or UO_1422 (O_1422,N_43967,N_49907);
and UO_1423 (O_1423,N_40956,N_49597);
nor UO_1424 (O_1424,N_44005,N_44603);
or UO_1425 (O_1425,N_40208,N_47237);
xnor UO_1426 (O_1426,N_44995,N_48449);
and UO_1427 (O_1427,N_40350,N_45101);
xnor UO_1428 (O_1428,N_40238,N_49079);
and UO_1429 (O_1429,N_42506,N_40978);
or UO_1430 (O_1430,N_40680,N_47004);
nand UO_1431 (O_1431,N_45550,N_40102);
and UO_1432 (O_1432,N_41585,N_47005);
nor UO_1433 (O_1433,N_43101,N_46550);
or UO_1434 (O_1434,N_41949,N_44710);
nand UO_1435 (O_1435,N_40580,N_46150);
xor UO_1436 (O_1436,N_40416,N_48856);
xnor UO_1437 (O_1437,N_41647,N_44524);
xnor UO_1438 (O_1438,N_41000,N_45326);
or UO_1439 (O_1439,N_49320,N_43422);
nand UO_1440 (O_1440,N_43157,N_40211);
nor UO_1441 (O_1441,N_42401,N_49595);
or UO_1442 (O_1442,N_44651,N_42753);
nand UO_1443 (O_1443,N_49038,N_46655);
nor UO_1444 (O_1444,N_43204,N_46928);
xor UO_1445 (O_1445,N_48840,N_46442);
nand UO_1446 (O_1446,N_49109,N_48913);
and UO_1447 (O_1447,N_46957,N_45013);
or UO_1448 (O_1448,N_46147,N_40467);
nor UO_1449 (O_1449,N_43680,N_44897);
xor UO_1450 (O_1450,N_43868,N_40101);
or UO_1451 (O_1451,N_42727,N_41873);
or UO_1452 (O_1452,N_41110,N_44625);
or UO_1453 (O_1453,N_46041,N_48739);
or UO_1454 (O_1454,N_43537,N_43342);
nand UO_1455 (O_1455,N_48201,N_46038);
and UO_1456 (O_1456,N_40388,N_43974);
nand UO_1457 (O_1457,N_42052,N_47561);
or UO_1458 (O_1458,N_45920,N_41942);
xor UO_1459 (O_1459,N_44516,N_44281);
and UO_1460 (O_1460,N_40516,N_41049);
nor UO_1461 (O_1461,N_41013,N_42828);
and UO_1462 (O_1462,N_43986,N_46154);
xor UO_1463 (O_1463,N_48695,N_43828);
xor UO_1464 (O_1464,N_47431,N_42155);
or UO_1465 (O_1465,N_44870,N_46761);
xor UO_1466 (O_1466,N_49119,N_47565);
xnor UO_1467 (O_1467,N_41584,N_47325);
nand UO_1468 (O_1468,N_41850,N_48555);
xnor UO_1469 (O_1469,N_46128,N_48439);
xnor UO_1470 (O_1470,N_42633,N_43746);
and UO_1471 (O_1471,N_42266,N_40673);
and UO_1472 (O_1472,N_44904,N_48984);
and UO_1473 (O_1473,N_44086,N_45946);
and UO_1474 (O_1474,N_45470,N_40455);
or UO_1475 (O_1475,N_48335,N_43838);
nor UO_1476 (O_1476,N_41245,N_41611);
or UO_1477 (O_1477,N_41137,N_42575);
nor UO_1478 (O_1478,N_44251,N_41669);
or UO_1479 (O_1479,N_43781,N_42306);
and UO_1480 (O_1480,N_49628,N_43149);
and UO_1481 (O_1481,N_49784,N_47633);
or UO_1482 (O_1482,N_49433,N_40607);
or UO_1483 (O_1483,N_47938,N_43900);
and UO_1484 (O_1484,N_44419,N_42501);
xor UO_1485 (O_1485,N_46359,N_43738);
xor UO_1486 (O_1486,N_46540,N_48781);
or UO_1487 (O_1487,N_45180,N_41183);
nor UO_1488 (O_1488,N_46600,N_45529);
nand UO_1489 (O_1489,N_48306,N_41821);
nor UO_1490 (O_1490,N_47030,N_43186);
nand UO_1491 (O_1491,N_47136,N_45773);
nand UO_1492 (O_1492,N_43771,N_42391);
xor UO_1493 (O_1493,N_45541,N_48699);
and UO_1494 (O_1494,N_48352,N_48318);
and UO_1495 (O_1495,N_41569,N_44202);
or UO_1496 (O_1496,N_43284,N_48552);
or UO_1497 (O_1497,N_48407,N_45451);
xnor UO_1498 (O_1498,N_49765,N_42373);
nand UO_1499 (O_1499,N_48108,N_40798);
nor UO_1500 (O_1500,N_41256,N_46177);
nor UO_1501 (O_1501,N_42114,N_42888);
or UO_1502 (O_1502,N_49879,N_46319);
and UO_1503 (O_1503,N_44920,N_44154);
and UO_1504 (O_1504,N_44048,N_49955);
and UO_1505 (O_1505,N_40253,N_44188);
or UO_1506 (O_1506,N_48001,N_48277);
or UO_1507 (O_1507,N_45293,N_40695);
xnor UO_1508 (O_1508,N_46034,N_42059);
xnor UO_1509 (O_1509,N_44349,N_42796);
nand UO_1510 (O_1510,N_49580,N_44024);
nor UO_1511 (O_1511,N_41775,N_47780);
nand UO_1512 (O_1512,N_42091,N_47572);
nand UO_1513 (O_1513,N_49652,N_44237);
xnor UO_1514 (O_1514,N_49901,N_44564);
xnor UO_1515 (O_1515,N_40169,N_44468);
nand UO_1516 (O_1516,N_49842,N_47702);
and UO_1517 (O_1517,N_44036,N_42126);
or UO_1518 (O_1518,N_45323,N_42201);
or UO_1519 (O_1519,N_46423,N_46270);
xnor UO_1520 (O_1520,N_44071,N_40832);
and UO_1521 (O_1521,N_40902,N_43918);
and UO_1522 (O_1522,N_44525,N_42107);
nand UO_1523 (O_1523,N_41356,N_43203);
or UO_1524 (O_1524,N_46414,N_48775);
nand UO_1525 (O_1525,N_44001,N_40134);
nand UO_1526 (O_1526,N_41364,N_42281);
and UO_1527 (O_1527,N_48002,N_45647);
xor UO_1528 (O_1528,N_45855,N_49921);
or UO_1529 (O_1529,N_46982,N_47656);
nor UO_1530 (O_1530,N_41209,N_46533);
nor UO_1531 (O_1531,N_48968,N_44027);
nand UO_1532 (O_1532,N_43368,N_45223);
or UO_1533 (O_1533,N_45061,N_43753);
and UO_1534 (O_1534,N_42189,N_48812);
xnor UO_1535 (O_1535,N_42662,N_41084);
or UO_1536 (O_1536,N_45998,N_41276);
or UO_1537 (O_1537,N_43034,N_48677);
or UO_1538 (O_1538,N_44013,N_46395);
and UO_1539 (O_1539,N_43471,N_44765);
and UO_1540 (O_1540,N_43308,N_49214);
or UO_1541 (O_1541,N_43152,N_47131);
and UO_1542 (O_1542,N_49209,N_44151);
and UO_1543 (O_1543,N_47409,N_47575);
or UO_1544 (O_1544,N_49113,N_46630);
xor UO_1545 (O_1545,N_40617,N_48638);
or UO_1546 (O_1546,N_44677,N_41479);
and UO_1547 (O_1547,N_47351,N_45607);
and UO_1548 (O_1548,N_49490,N_41983);
or UO_1549 (O_1549,N_43694,N_43307);
nor UO_1550 (O_1550,N_46869,N_41011);
nand UO_1551 (O_1551,N_48239,N_44941);
and UO_1552 (O_1552,N_49367,N_42925);
nor UO_1553 (O_1553,N_42859,N_40837);
xnor UO_1554 (O_1554,N_48691,N_43457);
or UO_1555 (O_1555,N_40804,N_44056);
xnor UO_1556 (O_1556,N_49050,N_44772);
and UO_1557 (O_1557,N_47646,N_41577);
xnor UO_1558 (O_1558,N_45075,N_45857);
nor UO_1559 (O_1559,N_41428,N_47491);
xor UO_1560 (O_1560,N_47260,N_44627);
and UO_1561 (O_1561,N_44103,N_43676);
and UO_1562 (O_1562,N_49970,N_41298);
nand UO_1563 (O_1563,N_45459,N_45357);
and UO_1564 (O_1564,N_48786,N_41237);
nor UO_1565 (O_1565,N_48309,N_44097);
or UO_1566 (O_1566,N_40233,N_43112);
and UO_1567 (O_1567,N_41780,N_42440);
and UO_1568 (O_1568,N_45669,N_40834);
nand UO_1569 (O_1569,N_45674,N_49064);
nand UO_1570 (O_1570,N_48215,N_42984);
xor UO_1571 (O_1571,N_47424,N_46859);
nand UO_1572 (O_1572,N_42932,N_47653);
nor UO_1573 (O_1573,N_45137,N_49757);
nand UO_1574 (O_1574,N_41164,N_41196);
nand UO_1575 (O_1575,N_48459,N_40602);
nand UO_1576 (O_1576,N_49404,N_44238);
nand UO_1577 (O_1577,N_40087,N_45099);
or UO_1578 (O_1578,N_48154,N_48004);
nand UO_1579 (O_1579,N_46271,N_44719);
or UO_1580 (O_1580,N_46684,N_45795);
or UO_1581 (O_1581,N_48156,N_44152);
and UO_1582 (O_1582,N_46245,N_40084);
or UO_1583 (O_1583,N_42139,N_41406);
nand UO_1584 (O_1584,N_48267,N_41146);
or UO_1585 (O_1585,N_41155,N_42636);
nor UO_1586 (O_1586,N_42835,N_46923);
nand UO_1587 (O_1587,N_40072,N_44351);
nand UO_1588 (O_1588,N_42012,N_41081);
and UO_1589 (O_1589,N_41977,N_41175);
or UO_1590 (O_1590,N_45404,N_49193);
nand UO_1591 (O_1591,N_45098,N_47506);
nor UO_1592 (O_1592,N_43921,N_48204);
and UO_1593 (O_1593,N_45437,N_47504);
nand UO_1594 (O_1594,N_40347,N_44373);
xor UO_1595 (O_1595,N_45340,N_48916);
nor UO_1596 (O_1596,N_41472,N_40894);
nor UO_1597 (O_1597,N_45547,N_48890);
or UO_1598 (O_1598,N_44517,N_44344);
or UO_1599 (O_1599,N_48839,N_46433);
nor UO_1600 (O_1600,N_49016,N_46500);
nand UO_1601 (O_1601,N_42289,N_42923);
and UO_1602 (O_1602,N_49777,N_41015);
nand UO_1603 (O_1603,N_47757,N_45927);
or UO_1604 (O_1604,N_47728,N_45822);
nand UO_1605 (O_1605,N_44359,N_44169);
and UO_1606 (O_1606,N_41266,N_48993);
and UO_1607 (O_1607,N_46335,N_42237);
or UO_1608 (O_1608,N_48031,N_46014);
xnor UO_1609 (O_1609,N_47588,N_45745);
nand UO_1610 (O_1610,N_44079,N_41204);
nand UO_1611 (O_1611,N_49603,N_44163);
nor UO_1612 (O_1612,N_45821,N_45496);
nand UO_1613 (O_1613,N_47347,N_45783);
nand UO_1614 (O_1614,N_49643,N_48258);
xnor UO_1615 (O_1615,N_45023,N_48807);
xnor UO_1616 (O_1616,N_48516,N_47765);
xor UO_1617 (O_1617,N_41597,N_49548);
and UO_1618 (O_1618,N_41725,N_47079);
xnor UO_1619 (O_1619,N_49565,N_41490);
nand UO_1620 (O_1620,N_45661,N_40650);
or UO_1621 (O_1621,N_43242,N_49599);
and UO_1622 (O_1622,N_41045,N_45947);
xnor UO_1623 (O_1623,N_40900,N_47753);
and UO_1624 (O_1624,N_41491,N_42326);
xnor UO_1625 (O_1625,N_43402,N_42074);
or UO_1626 (O_1626,N_49961,N_42408);
nand UO_1627 (O_1627,N_47117,N_49183);
and UO_1628 (O_1628,N_49670,N_46365);
and UO_1629 (O_1629,N_44410,N_42181);
nand UO_1630 (O_1630,N_40706,N_49721);
or UO_1631 (O_1631,N_47096,N_44910);
and UO_1632 (O_1632,N_49782,N_45273);
xnor UO_1633 (O_1633,N_44324,N_49494);
nor UO_1634 (O_1634,N_41043,N_44084);
and UO_1635 (O_1635,N_41697,N_43128);
nand UO_1636 (O_1636,N_41980,N_44834);
nor UO_1637 (O_1637,N_49608,N_41435);
and UO_1638 (O_1638,N_45881,N_40486);
nand UO_1639 (O_1639,N_40897,N_47484);
and UO_1640 (O_1640,N_40711,N_40076);
nand UO_1641 (O_1641,N_49104,N_41759);
and UO_1642 (O_1642,N_48692,N_47962);
and UO_1643 (O_1643,N_47870,N_44526);
or UO_1644 (O_1644,N_46835,N_49331);
and UO_1645 (O_1645,N_40544,N_46965);
or UO_1646 (O_1646,N_48333,N_42387);
and UO_1647 (O_1647,N_40899,N_47429);
nand UO_1648 (O_1648,N_41098,N_49405);
and UO_1649 (O_1649,N_47042,N_43943);
and UO_1650 (O_1650,N_47253,N_41442);
nor UO_1651 (O_1651,N_47212,N_42364);
nand UO_1652 (O_1652,N_44297,N_42842);
xnor UO_1653 (O_1653,N_47527,N_47121);
or UO_1654 (O_1654,N_41357,N_40667);
and UO_1655 (O_1655,N_46527,N_40548);
or UO_1656 (O_1656,N_44636,N_43113);
nand UO_1657 (O_1657,N_42269,N_48612);
or UO_1658 (O_1658,N_42177,N_48967);
or UO_1659 (O_1659,N_48210,N_44207);
nor UO_1660 (O_1660,N_41072,N_42043);
or UO_1661 (O_1661,N_46474,N_49323);
nor UO_1662 (O_1662,N_47033,N_40298);
nor UO_1663 (O_1663,N_41528,N_40924);
nand UO_1664 (O_1664,N_46113,N_45735);
or UO_1665 (O_1665,N_41608,N_47851);
and UO_1666 (O_1666,N_42849,N_46780);
nand UO_1667 (O_1667,N_45161,N_42283);
nand UO_1668 (O_1668,N_40243,N_44706);
and UO_1669 (O_1669,N_40321,N_49211);
and UO_1670 (O_1670,N_44994,N_44015);
nand UO_1671 (O_1671,N_42573,N_45240);
and UO_1672 (O_1672,N_46961,N_42111);
nand UO_1673 (O_1673,N_46478,N_44109);
and UO_1674 (O_1674,N_46204,N_45763);
xnor UO_1675 (O_1675,N_46730,N_43998);
nand UO_1676 (O_1676,N_46272,N_48409);
or UO_1677 (O_1677,N_44713,N_41048);
nand UO_1678 (O_1678,N_44263,N_45213);
and UO_1679 (O_1679,N_42723,N_44418);
nand UO_1680 (O_1680,N_47873,N_44258);
xnor UO_1681 (O_1681,N_44972,N_40431);
xnor UO_1682 (O_1682,N_41917,N_46164);
and UO_1683 (O_1683,N_43864,N_43498);
or UO_1684 (O_1684,N_41999,N_41261);
or UO_1685 (O_1685,N_44753,N_43229);
nand UO_1686 (O_1686,N_41904,N_45737);
and UO_1687 (O_1687,N_48793,N_41707);
nand UO_1688 (O_1688,N_45979,N_42272);
nor UO_1689 (O_1689,N_40085,N_45043);
xor UO_1690 (O_1690,N_41948,N_44600);
nor UO_1691 (O_1691,N_47499,N_40368);
or UO_1692 (O_1692,N_42607,N_43739);
and UO_1693 (O_1693,N_40599,N_41249);
nor UO_1694 (O_1694,N_47602,N_43855);
xor UO_1695 (O_1695,N_42751,N_43534);
nand UO_1696 (O_1696,N_43587,N_47020);
nor UO_1697 (O_1697,N_49534,N_40108);
and UO_1698 (O_1698,N_44294,N_42195);
nor UO_1699 (O_1699,N_47075,N_43094);
xnor UO_1700 (O_1700,N_40231,N_49551);
nand UO_1701 (O_1701,N_43592,N_41051);
xnor UO_1702 (O_1702,N_44556,N_46066);
or UO_1703 (O_1703,N_43691,N_42020);
nand UO_1704 (O_1704,N_44504,N_48185);
nand UO_1705 (O_1705,N_42834,N_48881);
and UO_1706 (O_1706,N_47734,N_44940);
nand UO_1707 (O_1707,N_43187,N_41801);
and UO_1708 (O_1708,N_41329,N_48655);
xor UO_1709 (O_1709,N_48423,N_45817);
or UO_1710 (O_1710,N_45932,N_40196);
nand UO_1711 (O_1711,N_47310,N_45016);
or UO_1712 (O_1712,N_44445,N_40822);
xnor UO_1713 (O_1713,N_47010,N_43071);
and UO_1714 (O_1714,N_48795,N_43143);
xor UO_1715 (O_1715,N_45720,N_41343);
nor UO_1716 (O_1716,N_49178,N_44177);
xor UO_1717 (O_1717,N_42968,N_43948);
and UO_1718 (O_1718,N_46471,N_44243);
xor UO_1719 (O_1719,N_47118,N_47254);
nor UO_1720 (O_1720,N_48358,N_40936);
nor UO_1721 (O_1721,N_40615,N_49242);
or UO_1722 (O_1722,N_45968,N_47221);
or UO_1723 (O_1723,N_46667,N_48848);
nor UO_1724 (O_1724,N_48619,N_45838);
or UO_1725 (O_1725,N_40719,N_46377);
nand UO_1726 (O_1726,N_47258,N_42611);
xor UO_1727 (O_1727,N_42803,N_44624);
xnor UO_1728 (O_1728,N_43142,N_43572);
nor UO_1729 (O_1729,N_41809,N_47607);
and UO_1730 (O_1730,N_45499,N_46991);
and UO_1731 (O_1731,N_44386,N_44683);
nor UO_1732 (O_1732,N_48868,N_49732);
nand UO_1733 (O_1733,N_45965,N_41966);
xnor UO_1734 (O_1734,N_47242,N_41501);
and UO_1735 (O_1735,N_45653,N_41093);
nor UO_1736 (O_1736,N_44655,N_46676);
nand UO_1737 (O_1737,N_41075,N_48406);
and UO_1738 (O_1738,N_41230,N_46257);
or UO_1739 (O_1739,N_42560,N_48534);
xor UO_1740 (O_1740,N_48623,N_40592);
xnor UO_1741 (O_1741,N_45507,N_47002);
xnor UO_1742 (O_1742,N_46907,N_40472);
and UO_1743 (O_1743,N_43656,N_43569);
nor UO_1744 (O_1744,N_49719,N_40949);
nand UO_1745 (O_1745,N_48054,N_48014);
or UO_1746 (O_1746,N_40657,N_42893);
xnor UO_1747 (O_1747,N_47827,N_49953);
and UO_1748 (O_1748,N_46664,N_42187);
nand UO_1749 (O_1749,N_49181,N_40788);
nand UO_1750 (O_1750,N_45638,N_40297);
nor UO_1751 (O_1751,N_49818,N_46696);
and UO_1752 (O_1752,N_42453,N_46526);
and UO_1753 (O_1753,N_42809,N_42554);
xor UO_1754 (O_1754,N_45513,N_43406);
nand UO_1755 (O_1755,N_47969,N_48007);
nor UO_1756 (O_1756,N_43885,N_47027);
xor UO_1757 (O_1757,N_40092,N_49613);
nand UO_1758 (O_1758,N_48884,N_43164);
nor UO_1759 (O_1759,N_45351,N_49908);
xnor UO_1760 (O_1760,N_47273,N_48932);
xnor UO_1761 (O_1761,N_42656,N_46850);
and UO_1762 (O_1762,N_48043,N_43486);
and UO_1763 (O_1763,N_47270,N_46494);
nor UO_1764 (O_1764,N_40646,N_49305);
xor UO_1765 (O_1765,N_44656,N_44901);
nand UO_1766 (O_1766,N_46348,N_46026);
xor UO_1767 (O_1767,N_49900,N_41478);
nor UO_1768 (O_1768,N_48563,N_46388);
nor UO_1769 (O_1769,N_44623,N_46392);
nor UO_1770 (O_1770,N_49240,N_40504);
and UO_1771 (O_1771,N_42227,N_48679);
xor UO_1772 (O_1772,N_48036,N_45070);
or UO_1773 (O_1773,N_47312,N_48270);
nor UO_1774 (O_1774,N_41563,N_44678);
nand UO_1775 (O_1775,N_42955,N_40137);
nor UO_1776 (O_1776,N_42777,N_47318);
nand UO_1777 (O_1777,N_45891,N_40629);
nor UO_1778 (O_1778,N_41327,N_42264);
nor UO_1779 (O_1779,N_47120,N_42570);
or UO_1780 (O_1780,N_44764,N_42894);
xnor UO_1781 (O_1781,N_47486,N_41886);
or UO_1782 (O_1782,N_45500,N_40453);
xor UO_1783 (O_1783,N_46949,N_42674);
or UO_1784 (O_1784,N_43621,N_47366);
xor UO_1785 (O_1785,N_47964,N_41474);
nand UO_1786 (O_1786,N_40588,N_49299);
or UO_1787 (O_1787,N_41385,N_41198);
nand UO_1788 (O_1788,N_45574,N_49715);
nand UO_1789 (O_1789,N_49962,N_45165);
nand UO_1790 (O_1790,N_48696,N_47327);
xor UO_1791 (O_1791,N_47441,N_40482);
nor UO_1792 (O_1792,N_45488,N_44213);
or UO_1793 (O_1793,N_49738,N_44475);
and UO_1794 (O_1794,N_43931,N_47733);
nand UO_1795 (O_1795,N_44302,N_43059);
xor UO_1796 (O_1796,N_48399,N_40850);
xor UO_1797 (O_1797,N_49885,N_40390);
nor UO_1798 (O_1798,N_40997,N_48537);
nor UO_1799 (O_1799,N_45811,N_46727);
xor UO_1800 (O_1800,N_41077,N_43818);
and UO_1801 (O_1801,N_46693,N_44153);
and UO_1802 (O_1802,N_45641,N_49912);
and UO_1803 (O_1803,N_49560,N_45603);
nor UO_1804 (O_1804,N_46427,N_42069);
or UO_1805 (O_1805,N_47144,N_48861);
or UO_1806 (O_1806,N_46634,N_42347);
xor UO_1807 (O_1807,N_49391,N_47423);
nor UO_1808 (O_1808,N_40651,N_48971);
xor UO_1809 (O_1809,N_42524,N_45320);
nor UO_1810 (O_1810,N_46247,N_46897);
or UO_1811 (O_1811,N_48487,N_47917);
nor UO_1812 (O_1812,N_42772,N_42789);
or UO_1813 (O_1813,N_48164,N_43131);
or UO_1814 (O_1814,N_49477,N_47857);
and UO_1815 (O_1815,N_43174,N_40712);
xnor UO_1816 (O_1816,N_48899,N_45227);
nor UO_1817 (O_1817,N_44051,N_43217);
or UO_1818 (O_1818,N_47798,N_41803);
xnor UO_1819 (O_1819,N_42565,N_49387);
nor UO_1820 (O_1820,N_46734,N_48011);
nor UO_1821 (O_1821,N_44354,N_40791);
nor UO_1822 (O_1822,N_41425,N_48596);
xnor UO_1823 (O_1823,N_43482,N_46108);
nand UO_1824 (O_1824,N_42853,N_49559);
or UO_1825 (O_1825,N_41016,N_49581);
nor UO_1826 (O_1826,N_44639,N_45796);
nor UO_1827 (O_1827,N_47658,N_48259);
nand UO_1828 (O_1828,N_47044,N_46880);
nand UO_1829 (O_1829,N_49736,N_40841);
nand UO_1830 (O_1830,N_45691,N_42158);
and UO_1831 (O_1831,N_44980,N_43124);
nor UO_1832 (O_1832,N_48253,N_46832);
xor UO_1833 (O_1833,N_48327,N_45073);
nor UO_1834 (O_1834,N_43732,N_44543);
nor UO_1835 (O_1835,N_42709,N_49203);
and UO_1836 (O_1836,N_47803,N_46762);
nand UO_1837 (O_1837,N_45045,N_46040);
and UO_1838 (O_1838,N_42707,N_47760);
or UO_1839 (O_1839,N_47127,N_42731);
nor UO_1840 (O_1840,N_40420,N_43376);
nor UO_1841 (O_1841,N_40364,N_45939);
nor UO_1842 (O_1842,N_49706,N_41150);
or UO_1843 (O_1843,N_43111,N_48482);
nand UO_1844 (O_1844,N_46650,N_44519);
nor UO_1845 (O_1845,N_45633,N_43907);
nor UO_1846 (O_1846,N_43068,N_45937);
nor UO_1847 (O_1847,N_46344,N_45751);
nor UO_1848 (O_1848,N_45403,N_43924);
nand UO_1849 (O_1849,N_47485,N_41835);
nand UO_1850 (O_1850,N_45386,N_48908);
or UO_1851 (O_1851,N_48321,N_42505);
and UO_1852 (O_1852,N_41213,N_48964);
nor UO_1853 (O_1853,N_43180,N_49667);
or UO_1854 (O_1854,N_48281,N_43027);
or UO_1855 (O_1855,N_46448,N_45370);
nor UO_1856 (O_1856,N_47643,N_44866);
or UO_1857 (O_1857,N_48304,N_48565);
xor UO_1858 (O_1858,N_44986,N_47380);
nor UO_1859 (O_1859,N_42758,N_49949);
and UO_1860 (O_1860,N_48578,N_41531);
nand UO_1861 (O_1861,N_49576,N_41468);
nand UO_1862 (O_1862,N_47847,N_45910);
nor UO_1863 (O_1863,N_46021,N_44922);
nor UO_1864 (O_1864,N_49442,N_42438);
and UO_1865 (O_1865,N_47104,N_46863);
or UO_1866 (O_1866,N_40604,N_49002);
xnor UO_1867 (O_1867,N_47263,N_49529);
nor UO_1868 (O_1868,N_43705,N_40974);
nand UO_1869 (O_1869,N_47176,N_49624);
nor UO_1870 (O_1870,N_46541,N_45467);
and UO_1871 (O_1871,N_40943,N_46553);
nor UO_1872 (O_1872,N_40522,N_47336);
nand UO_1873 (O_1873,N_45911,N_49499);
nand UO_1874 (O_1874,N_46935,N_45572);
xor UO_1875 (O_1875,N_45836,N_40051);
xnor UO_1876 (O_1876,N_48525,N_45466);
nand UO_1877 (O_1877,N_48838,N_40931);
or UO_1878 (O_1878,N_47611,N_42208);
or UO_1879 (O_1879,N_40465,N_45885);
and UO_1880 (O_1880,N_44100,N_43845);
or UO_1881 (O_1881,N_43637,N_41825);
nor UO_1882 (O_1882,N_42625,N_44826);
nor UO_1883 (O_1883,N_40881,N_40001);
nor UO_1884 (O_1884,N_44401,N_48401);
and UO_1885 (O_1885,N_48961,N_44018);
or UO_1886 (O_1886,N_41950,N_46205);
xnor UO_1887 (O_1887,N_46415,N_47555);
and UO_1888 (O_1888,N_46639,N_47346);
or UO_1889 (O_1889,N_41763,N_47899);
or UO_1890 (O_1890,N_47554,N_45237);
or UO_1891 (O_1891,N_43429,N_45118);
nand UO_1892 (O_1892,N_43479,N_49148);
xor UO_1893 (O_1893,N_48928,N_46802);
nand UO_1894 (O_1894,N_43902,N_41810);
xor UO_1895 (O_1895,N_42343,N_47737);
nor UO_1896 (O_1896,N_45381,N_41113);
or UO_1897 (O_1897,N_43760,N_40753);
or UO_1898 (O_1898,N_46281,N_40413);
nor UO_1899 (O_1899,N_40889,N_48283);
xor UO_1900 (O_1900,N_42956,N_45715);
nor UO_1901 (O_1901,N_44155,N_44593);
nand UO_1902 (O_1902,N_45719,N_43194);
nor UO_1903 (O_1903,N_49801,N_42958);
or UO_1904 (O_1904,N_45477,N_40223);
nand UO_1905 (O_1905,N_40979,N_48931);
or UO_1906 (O_1906,N_45153,N_46793);
xnor UO_1907 (O_1907,N_49936,N_40079);
and UO_1908 (O_1908,N_42314,N_47783);
and UO_1909 (O_1909,N_47927,N_48755);
xnor UO_1910 (O_1910,N_42395,N_47961);
or UO_1911 (O_1911,N_44259,N_41398);
and UO_1912 (O_1912,N_42017,N_42443);
nor UO_1913 (O_1913,N_42209,N_49755);
and UO_1914 (O_1914,N_42389,N_47908);
nor UO_1915 (O_1915,N_48725,N_41055);
xnor UO_1916 (O_1916,N_49911,N_49133);
or UO_1917 (O_1917,N_41674,N_41391);
xor UO_1918 (O_1918,N_48356,N_47600);
xnor UO_1919 (O_1919,N_44376,N_47796);
or UO_1920 (O_1920,N_40710,N_49841);
and UO_1921 (O_1921,N_45951,N_47888);
or UO_1922 (O_1922,N_42735,N_43107);
nor UO_1923 (O_1923,N_49201,N_43181);
or UO_1924 (O_1924,N_44871,N_44521);
xor UO_1925 (O_1925,N_40109,N_42583);
xor UO_1926 (O_1926,N_40139,N_44127);
or UO_1927 (O_1927,N_46280,N_40662);
nand UO_1928 (O_1928,N_46481,N_43629);
xor UO_1929 (O_1929,N_45182,N_45894);
or UO_1930 (O_1930,N_48351,N_48990);
nor UO_1931 (O_1931,N_45552,N_48743);
nor UO_1932 (O_1932,N_48574,N_46815);
or UO_1933 (O_1933,N_40526,N_49772);
and UO_1934 (O_1934,N_47512,N_43437);
and UO_1935 (O_1935,N_49924,N_40738);
nor UO_1936 (O_1936,N_45805,N_47373);
xnor UO_1937 (O_1937,N_40925,N_47630);
nor UO_1938 (O_1938,N_49512,N_49054);
nor UO_1939 (O_1939,N_49756,N_42248);
xnor UO_1940 (O_1940,N_49832,N_46332);
nand UO_1941 (O_1941,N_41279,N_46641);
nor UO_1942 (O_1942,N_41645,N_49091);
nand UO_1943 (O_1943,N_41989,N_48424);
xor UO_1944 (O_1944,N_40019,N_43788);
nand UO_1945 (O_1945,N_45587,N_44423);
and UO_1946 (O_1946,N_40305,N_49037);
or UO_1947 (O_1947,N_48554,N_40758);
or UO_1948 (O_1948,N_46556,N_45024);
xor UO_1949 (O_1949,N_48313,N_49632);
and UO_1950 (O_1950,N_43836,N_43389);
or UO_1951 (O_1951,N_45512,N_42278);
and UO_1952 (O_1952,N_43936,N_47041);
and UO_1953 (O_1953,N_42770,N_47088);
nor UO_1954 (O_1954,N_49609,N_40783);
nand UO_1955 (O_1955,N_45339,N_43126);
or UO_1956 (O_1956,N_49805,N_46674);
and UO_1957 (O_1957,N_40400,N_47401);
xor UO_1958 (O_1958,N_49142,N_46063);
and UO_1959 (O_1959,N_41161,N_46371);
nor UO_1960 (O_1960,N_49671,N_41769);
nor UO_1961 (O_1961,N_49272,N_40559);
nand UO_1962 (O_1962,N_45341,N_48806);
xnor UO_1963 (O_1963,N_46095,N_45014);
nor UO_1964 (O_1964,N_46971,N_44877);
nand UO_1965 (O_1965,N_42655,N_45829);
or UO_1966 (O_1966,N_42665,N_44931);
xor UO_1967 (O_1967,N_49026,N_46690);
and UO_1968 (O_1968,N_49451,N_44138);
nand UO_1969 (O_1969,N_49708,N_43379);
or UO_1970 (O_1970,N_43857,N_42378);
nand UO_1971 (O_1971,N_41800,N_40608);
nor UO_1972 (O_1972,N_41370,N_40206);
or UO_1973 (O_1973,N_41624,N_42385);
xor UO_1974 (O_1974,N_49523,N_46889);
or UO_1975 (O_1975,N_42596,N_42276);
nor UO_1976 (O_1976,N_44681,N_41721);
xor UO_1977 (O_1977,N_49552,N_44535);
xor UO_1978 (O_1978,N_44685,N_41592);
and UO_1979 (O_1979,N_49659,N_44394);
xnor UO_1980 (O_1980,N_43671,N_46983);
or UO_1981 (O_1981,N_45634,N_40590);
or UO_1982 (O_1982,N_42095,N_41856);
and UO_1983 (O_1983,N_49174,N_44819);
and UO_1984 (O_1984,N_49813,N_41473);
xnor UO_1985 (O_1985,N_49555,N_45136);
nand UO_1986 (O_1986,N_41831,N_40818);
and UO_1987 (O_1987,N_44119,N_49471);
xor UO_1988 (O_1988,N_45974,N_45083);
and UO_1989 (O_1989,N_49510,N_46951);
nor UO_1990 (O_1990,N_45284,N_48100);
nor UO_1991 (O_1991,N_41603,N_46487);
nor UO_1992 (O_1992,N_48536,N_49904);
nor UO_1993 (O_1993,N_43169,N_44709);
and UO_1994 (O_1994,N_46522,N_48410);
nand UO_1995 (O_1995,N_48115,N_49730);
nand UO_1996 (O_1996,N_46229,N_49536);
xnor UO_1997 (O_1997,N_48437,N_44617);
nand UO_1998 (O_1998,N_49769,N_44498);
and UO_1999 (O_1999,N_41731,N_43077);
or UO_2000 (O_2000,N_44511,N_49942);
nor UO_2001 (O_2001,N_44629,N_47960);
nor UO_2002 (O_2002,N_41136,N_46085);
nor UO_2003 (O_2003,N_42081,N_47368);
xor UO_2004 (O_2004,N_47095,N_44782);
and UO_2005 (O_2005,N_44985,N_40734);
nor UO_2006 (O_2006,N_45212,N_49683);
nor UO_2007 (O_2007,N_42188,N_48250);
xnor UO_2008 (O_2008,N_41407,N_47476);
nand UO_2009 (O_2009,N_44626,N_47432);
nor UO_2010 (O_2010,N_43888,N_43561);
nand UO_2011 (O_2011,N_40904,N_40077);
and UO_2012 (O_2012,N_45853,N_47084);
or UO_2013 (O_2013,N_41673,N_43935);
xor UO_2014 (O_2014,N_40528,N_45554);
nand UO_2015 (O_2015,N_44562,N_40623);
or UO_2016 (O_2016,N_40767,N_46868);
and UO_2017 (O_2017,N_40903,N_43757);
or UO_2018 (O_2018,N_48260,N_41165);
and UO_2019 (O_2019,N_46547,N_43066);
or UO_2020 (O_2020,N_41580,N_44219);
and UO_2021 (O_2021,N_40950,N_44179);
nand UO_2022 (O_2022,N_47459,N_46152);
nor UO_2023 (O_2023,N_43137,N_49735);
xor UO_2024 (O_2024,N_42025,N_41970);
nand UO_2025 (O_2025,N_40365,N_41957);
xor UO_2026 (O_2026,N_40907,N_49269);
nand UO_2027 (O_2027,N_41922,N_40663);
nor UO_2028 (O_2028,N_49304,N_44211);
xor UO_2029 (O_2029,N_41726,N_49185);
xnor UO_2030 (O_2030,N_48296,N_49136);
and UO_2031 (O_2031,N_49612,N_41910);
and UO_2032 (O_2032,N_45217,N_40946);
nand UO_2033 (O_2033,N_47492,N_47735);
nor UO_2034 (O_2034,N_49228,N_44795);
nor UO_2035 (O_2035,N_48604,N_43949);
nor UO_2036 (O_2036,N_40656,N_48688);
and UO_2037 (O_2037,N_49780,N_42555);
xnor UO_2038 (O_2038,N_47138,N_41477);
and UO_2039 (O_2039,N_42348,N_47579);
xnor UO_2040 (O_2040,N_46316,N_44189);
nor UO_2041 (O_2041,N_49436,N_46794);
nand UO_2042 (O_2042,N_42215,N_43269);
nand UO_2043 (O_2043,N_47036,N_43403);
and UO_2044 (O_2044,N_45726,N_46037);
nand UO_2045 (O_2045,N_47357,N_40948);
and UO_2046 (O_2046,N_47397,N_48128);
and UO_2047 (O_2047,N_46885,N_40929);
and UO_2048 (O_2048,N_48438,N_44306);
xor UO_2049 (O_2049,N_49760,N_44514);
nor UO_2050 (O_2050,N_49068,N_40560);
and UO_2051 (O_2051,N_47293,N_48782);
nand UO_2052 (O_2052,N_42610,N_46143);
nand UO_2053 (O_2053,N_40585,N_47209);
or UO_2054 (O_2054,N_41844,N_49237);
xnor UO_2055 (O_2055,N_42006,N_45896);
or UO_2056 (O_2056,N_42336,N_43012);
and UO_2057 (O_2057,N_42113,N_48959);
and UO_2058 (O_2058,N_46569,N_44599);
nor UO_2059 (O_2059,N_48086,N_40412);
or UO_2060 (O_2060,N_42172,N_40880);
and UO_2061 (O_2061,N_44875,N_49629);
nor UO_2062 (O_2062,N_43763,N_48172);
nand UO_2063 (O_2063,N_46890,N_47587);
xor UO_2064 (O_2064,N_43133,N_46482);
and UO_2065 (O_2065,N_40396,N_43285);
xor UO_2066 (O_2066,N_43641,N_41595);
nor UO_2067 (O_2067,N_49114,N_48709);
xor UO_2068 (O_2068,N_42457,N_41359);
and UO_2069 (O_2069,N_45485,N_47845);
nor UO_2070 (O_2070,N_45205,N_41499);
nand UO_2071 (O_2071,N_49213,N_41973);
nor UO_2072 (O_2072,N_41760,N_43026);
xor UO_2073 (O_2073,N_41594,N_46733);
or UO_2074 (O_2074,N_45376,N_44610);
or UO_2075 (O_2075,N_42361,N_41125);
or UO_2076 (O_2076,N_40620,N_43007);
nor UO_2077 (O_2077,N_45844,N_42621);
nand UO_2078 (O_2078,N_43292,N_46822);
and UO_2079 (O_2079,N_47752,N_48062);
nor UO_2080 (O_2080,N_47883,N_41857);
nor UO_2081 (O_2081,N_46091,N_42477);
or UO_2082 (O_2082,N_45907,N_49705);
nor UO_2083 (O_2083,N_41167,N_42194);
or UO_2084 (O_2084,N_43823,N_49177);
nand UO_2085 (O_2085,N_42097,N_45209);
xor UO_2086 (O_2086,N_41765,N_43454);
and UO_2087 (O_2087,N_40391,N_40474);
nor UO_2088 (O_2088,N_46057,N_45094);
xnor UO_2089 (O_2089,N_44220,N_48477);
and UO_2090 (O_2090,N_49550,N_48643);
xor UO_2091 (O_2091,N_41719,N_45203);
xor UO_2092 (O_2092,N_43182,N_45573);
xor UO_2093 (O_2093,N_44674,N_44378);
nand UO_2094 (O_2094,N_42411,N_42164);
and UO_2095 (O_2095,N_47515,N_43896);
or UO_2096 (O_2096,N_49360,N_40172);
nor UO_2097 (O_2097,N_45258,N_45186);
or UO_2098 (O_2098,N_40641,N_46567);
or UO_2099 (O_2099,N_42075,N_47863);
or UO_2100 (O_2100,N_49741,N_43377);
xnor UO_2101 (O_2101,N_45416,N_40799);
and UO_2102 (O_2102,N_42018,N_46246);
xor UO_2103 (O_2103,N_45082,N_41848);
nand UO_2104 (O_2104,N_43531,N_41955);
or UO_2105 (O_2105,N_44311,N_42011);
nor UO_2106 (O_2106,N_44428,N_41133);
nand UO_2107 (O_2107,N_45846,N_45786);
or UO_2108 (O_2108,N_46171,N_43075);
or UO_2109 (O_2109,N_47399,N_40730);
and UO_2110 (O_2110,N_47531,N_40980);
or UO_2111 (O_2111,N_44063,N_45872);
and UO_2112 (O_2112,N_44110,N_46329);
nand UO_2113 (O_2113,N_46927,N_41168);
or UO_2114 (O_2114,N_47943,N_45133);
nand UO_2115 (O_2115,N_41832,N_47833);
xnor UO_2116 (O_2116,N_42315,N_47875);
nor UO_2117 (O_2117,N_49484,N_47302);
nand UO_2118 (O_2118,N_47474,N_46609);
and UO_2119 (O_2119,N_49032,N_48470);
nor UO_2120 (O_2120,N_48986,N_45793);
and UO_2121 (O_2121,N_40444,N_42479);
nand UO_2122 (O_2122,N_43081,N_49889);
xor UO_2123 (O_2123,N_49987,N_44810);
or UO_2124 (O_2124,N_44078,N_40694);
nor UO_2125 (O_2125,N_48549,N_44853);
nand UO_2126 (O_2126,N_46575,N_40338);
and UO_2127 (O_2127,N_44252,N_44195);
xnor UO_2128 (O_2128,N_46666,N_42734);
or UO_2129 (O_2129,N_44914,N_40181);
xnor UO_2130 (O_2130,N_41778,N_45828);
and UO_2131 (O_2131,N_45110,N_47256);
nor UO_2132 (O_2132,N_40100,N_45862);
or UO_2133 (O_2133,N_44388,N_42085);
and UO_2134 (O_2134,N_45589,N_45190);
nand UO_2135 (O_2135,N_41940,N_41959);
xnor UO_2136 (O_2136,N_43903,N_43469);
and UO_2137 (O_2137,N_45027,N_44630);
xor UO_2138 (O_2138,N_43407,N_42640);
nor UO_2139 (O_2139,N_47945,N_47544);
xor UO_2140 (O_2140,N_48844,N_43063);
and UO_2141 (O_2141,N_48473,N_49887);
nand UO_2142 (O_2142,N_40593,N_49326);
nand UO_2143 (O_2143,N_43549,N_48680);
nand UO_2144 (O_2144,N_47616,N_40021);
or UO_2145 (O_2145,N_47743,N_41628);
or UO_2146 (O_2146,N_40807,N_45527);
nand UO_2147 (O_2147,N_44012,N_47662);
xor UO_2148 (O_2148,N_42243,N_47359);
xnor UO_2149 (O_2149,N_47937,N_44338);
and UO_2150 (O_2150,N_48488,N_48641);
nor UO_2151 (O_2151,N_48104,N_48904);
nand UO_2152 (O_2152,N_47179,N_40200);
or UO_2153 (O_2153,N_47514,N_42088);
nand UO_2154 (O_2154,N_43793,N_49309);
nand UO_2155 (O_2155,N_41456,N_47503);
xor UO_2156 (O_2156,N_42686,N_44807);
nand UO_2157 (O_2157,N_41287,N_41430);
or UO_2158 (O_2158,N_48824,N_45583);
and UO_2159 (O_2159,N_42637,N_44032);
xor UO_2160 (O_2160,N_46161,N_40197);
nor UO_2161 (O_2161,N_48357,N_46473);
nor UO_2162 (O_2162,N_47963,N_49945);
xnor UO_2163 (O_2163,N_47738,N_46903);
or UO_2164 (O_2164,N_48533,N_45640);
nand UO_2165 (O_2165,N_43030,N_42048);
xor UO_2166 (O_2166,N_43473,N_49946);
and UO_2167 (O_2167,N_42235,N_41730);
and UO_2168 (O_2168,N_48924,N_45206);
nand UO_2169 (O_2169,N_42913,N_49660);
nor UO_2170 (O_2170,N_40213,N_49161);
or UO_2171 (O_2171,N_45447,N_46959);
and UO_2172 (O_2172,N_46561,N_46633);
nor UO_2173 (O_2173,N_42804,N_45676);
or UO_2174 (O_2174,N_45625,N_47334);
or UO_2175 (O_2175,N_44111,N_45387);
and UO_2176 (O_2176,N_44215,N_44939);
xor UO_2177 (O_2177,N_47381,N_40300);
nand UO_2178 (O_2178,N_42160,N_41789);
nand UO_2179 (O_2179,N_46446,N_46906);
and UO_2180 (O_2180,N_49226,N_43374);
or UO_2181 (O_2181,N_49093,N_44966);
nand UO_2182 (O_2182,N_45802,N_43117);
or UO_2183 (O_2183,N_49092,N_49417);
nand UO_2184 (O_2184,N_49312,N_40163);
and UO_2185 (O_2185,N_41738,N_48316);
nor UO_2186 (O_2186,N_45736,N_47155);
xnor UO_2187 (O_2187,N_41102,N_41991);
and UO_2188 (O_2188,N_41637,N_47591);
nand UO_2189 (O_2189,N_40449,N_40874);
nand UO_2190 (O_2190,N_41342,N_41153);
or UO_2191 (O_2191,N_48003,N_46807);
or UO_2192 (O_2192,N_44253,N_49207);
nor UO_2193 (O_2193,N_49076,N_41916);
xor UO_2194 (O_2194,N_46096,N_47634);
or UO_2195 (O_2195,N_42162,N_41776);
xor UO_2196 (O_2196,N_46129,N_46582);
and UO_2197 (O_2197,N_41661,N_45316);
and UO_2198 (O_2198,N_44612,N_43475);
nand UO_2199 (O_2199,N_47810,N_46908);
nor UO_2200 (O_2200,N_48922,N_44318);
or UO_2201 (O_2201,N_47918,N_42210);
and UO_2202 (O_2202,N_40562,N_45766);
and UO_2203 (O_2203,N_45759,N_49823);
or UO_2204 (O_2204,N_46534,N_41915);
and UO_2205 (O_2205,N_49364,N_40679);
xnor UO_2206 (O_2206,N_41192,N_45253);
xor UO_2207 (O_2207,N_40091,N_41705);
nand UO_2208 (O_2208,N_44298,N_48246);
xor UO_2209 (O_2209,N_49567,N_48486);
or UO_2210 (O_2210,N_46984,N_49275);
nand UO_2211 (O_2211,N_48175,N_45721);
or UO_2212 (O_2212,N_44035,N_47820);
and UO_2213 (O_2213,N_47321,N_43983);
nor UO_2214 (O_2214,N_47675,N_46954);
nor UO_2215 (O_2215,N_43459,N_43381);
nor UO_2216 (O_2216,N_40367,N_46055);
xnor UO_2217 (O_2217,N_48339,N_47143);
nor UO_2218 (O_2218,N_42896,N_48787);
or UO_2219 (O_2219,N_44435,N_41972);
nor UO_2220 (O_2220,N_43326,N_48413);
and UO_2221 (O_2221,N_46039,N_47818);
or UO_2222 (O_2222,N_45347,N_43056);
nor UO_2223 (O_2223,N_44815,N_47604);
nor UO_2224 (O_2224,N_42683,N_48113);
xnor UO_2225 (O_2225,N_40625,N_40247);
nor UO_2226 (O_2226,N_47552,N_46151);
nor UO_2227 (O_2227,N_46302,N_47563);
xor UO_2228 (O_2228,N_44131,N_45071);
nand UO_2229 (O_2229,N_46821,N_40634);
xor UO_2230 (O_2230,N_40436,N_46608);
xnor UO_2231 (O_2231,N_42867,N_41216);
and UO_2232 (O_2232,N_45659,N_43250);
or UO_2233 (O_2233,N_47289,N_45185);
nand UO_2234 (O_2234,N_46814,N_43345);
xnor UO_2235 (O_2235,N_42516,N_48157);
and UO_2236 (O_2236,N_43565,N_41527);
nand UO_2237 (O_2237,N_43020,N_40042);
and UO_2238 (O_2238,N_48814,N_40315);
and UO_2239 (O_2239,N_40477,N_45559);
and UO_2240 (O_2240,N_43214,N_48474);
nand UO_2241 (O_2241,N_48885,N_43035);
nor UO_2242 (O_2242,N_46155,N_47150);
nor UO_2243 (O_2243,N_43514,N_42468);
and UO_2244 (O_2244,N_45718,N_48145);
and UO_2245 (O_2245,N_44788,N_49663);
and UO_2246 (O_2246,N_44880,N_47037);
and UO_2247 (O_2247,N_40369,N_41483);
xnor UO_2248 (O_2248,N_47983,N_46881);
and UO_2249 (O_2249,N_48006,N_48195);
nor UO_2250 (O_2250,N_40591,N_46054);
or UO_2251 (O_2251,N_42327,N_46425);
or UO_2252 (O_2252,N_49883,N_45482);
and UO_2253 (O_2253,N_41255,N_48116);
xnor UO_2254 (O_2254,N_46554,N_45810);
and UO_2255 (O_2255,N_48609,N_40985);
xor UO_2256 (O_2256,N_40491,N_46871);
and UO_2257 (O_2257,N_40760,N_46857);
xnor UO_2258 (O_2258,N_43273,N_48985);
nor UO_2259 (O_2259,N_41667,N_45032);
or UO_2260 (O_2260,N_41805,N_49474);
nor UO_2261 (O_2261,N_41352,N_42157);
or UO_2262 (O_2262,N_42028,N_41304);
and UO_2263 (O_2263,N_44594,N_44443);
and UO_2264 (O_2264,N_44313,N_48601);
or UO_2265 (O_2265,N_42563,N_47929);
and UO_2266 (O_2266,N_41152,N_42850);
or UO_2267 (O_2267,N_45012,N_48140);
and UO_2268 (O_2268,N_49409,N_44776);
and UO_2269 (O_2269,N_42733,N_49808);
nor UO_2270 (O_2270,N_46470,N_43626);
xnor UO_2271 (O_2271,N_46757,N_47661);
and UO_2272 (O_2272,N_47771,N_40245);
xnor UO_2273 (O_2273,N_49137,N_42533);
xnor UO_2274 (O_2274,N_42261,N_41142);
and UO_2275 (O_2275,N_42367,N_44014);
xor UO_2276 (O_2276,N_41323,N_45815);
or UO_2277 (O_2277,N_47596,N_44652);
nand UO_2278 (O_2278,N_48556,N_43976);
or UO_2279 (O_2279,N_42536,N_49216);
and UO_2280 (O_2280,N_41515,N_45568);
nor UO_2281 (O_2281,N_41994,N_44918);
xnor UO_2282 (O_2282,N_43158,N_49803);
or UO_2283 (O_2283,N_44989,N_48698);
or UO_2284 (O_2284,N_48706,N_42103);
xnor UO_2285 (O_2285,N_44224,N_42129);
xnor UO_2286 (O_2286,N_42797,N_42517);
xnor UO_2287 (O_2287,N_40015,N_40414);
and UO_2288 (O_2288,N_46259,N_43493);
or UO_2289 (O_2289,N_41450,N_44112);
nor UO_2290 (O_2290,N_41012,N_49573);
nand UO_2291 (O_2291,N_43917,N_44726);
nand UO_2292 (O_2292,N_45181,N_41547);
or UO_2293 (O_2293,N_48830,N_46019);
or UO_2294 (O_2294,N_49691,N_48489);
nand UO_2295 (O_2295,N_41318,N_42785);
nor UO_2296 (O_2296,N_44808,N_40800);
xor UO_2297 (O_2297,N_42543,N_49807);
nand UO_2298 (O_2298,N_43132,N_46103);
and UO_2299 (O_2299,N_42121,N_40311);
or UO_2300 (O_2300,N_40171,N_45908);
or UO_2301 (O_2301,N_48747,N_46911);
xor UO_2302 (O_2302,N_47078,N_41185);
and UO_2303 (O_2303,N_48158,N_49541);
or UO_2304 (O_2304,N_46086,N_44272);
and UO_2305 (O_2305,N_40819,N_40336);
xnor UO_2306 (O_2306,N_43462,N_40628);
or UO_2307 (O_2307,N_41985,N_40966);
xor UO_2308 (O_2308,N_41609,N_46737);
or UO_2309 (O_2309,N_43355,N_41377);
nor UO_2310 (O_2310,N_40260,N_47569);
or UO_2311 (O_2311,N_49861,N_40600);
nor UO_2312 (O_2312,N_49080,N_48197);
and UO_2313 (O_2313,N_46121,N_40373);
and UO_2314 (O_2314,N_48125,N_43136);
and UO_2315 (O_2315,N_44502,N_43844);
nand UO_2316 (O_2316,N_48950,N_44077);
or UO_2317 (O_2317,N_43032,N_43729);
xor UO_2318 (O_2318,N_41562,N_48425);
and UO_2319 (O_2319,N_42566,N_43556);
nor UO_2320 (O_2320,N_43215,N_45967);
or UO_2321 (O_2321,N_47275,N_45296);
nand UO_2322 (O_2322,N_46165,N_40639);
nor UO_2323 (O_2323,N_46586,N_43076);
and UO_2324 (O_2324,N_43518,N_41626);
nor UO_2325 (O_2325,N_40538,N_46483);
nand UO_2326 (O_2326,N_41646,N_48289);
or UO_2327 (O_2327,N_49686,N_40257);
nand UO_2328 (O_2328,N_43503,N_41201);
xor UO_2329 (O_2329,N_43271,N_48272);
xnor UO_2330 (O_2330,N_42344,N_40251);
nor UO_2331 (O_2331,N_46539,N_43252);
and UO_2332 (O_2332,N_45394,N_45306);
or UO_2333 (O_2333,N_41366,N_49406);
nand UO_2334 (O_2334,N_43316,N_48265);
and UO_2335 (O_2335,N_40700,N_40860);
nand UO_2336 (O_2336,N_45978,N_41289);
nor UO_2337 (O_2337,N_47068,N_47589);
nand UO_2338 (O_2338,N_44327,N_42116);
xor UO_2339 (O_2339,N_40866,N_46310);
or UO_2340 (O_2340,N_47581,N_48230);
and UO_2341 (O_2341,N_42638,N_46698);
nand UO_2342 (O_2342,N_40136,N_43611);
and UO_2343 (O_2343,N_42890,N_42196);
or UO_2344 (O_2344,N_44425,N_45664);
or UO_2345 (O_2345,N_45321,N_42257);
xor UO_2346 (O_2346,N_47067,N_47265);
or UO_2347 (O_2347,N_45518,N_49110);
nand UO_2348 (O_2348,N_42779,N_43939);
xor UO_2349 (O_2349,N_45031,N_42872);
nand UO_2350 (O_2350,N_40722,N_42759);
nor UO_2351 (O_2351,N_44740,N_48417);
xnor UO_2352 (O_2352,N_48642,N_45666);
and UO_2353 (O_2353,N_47164,N_45873);
or UO_2354 (O_2354,N_41222,N_42251);
and UO_2355 (O_2355,N_42094,N_46166);
xor UO_2356 (O_2356,N_42651,N_42319);
or UO_2357 (O_2357,N_41877,N_47654);
nor UO_2358 (O_2358,N_45063,N_48976);
nand UO_2359 (O_2359,N_41958,N_45729);
and UO_2360 (O_2360,N_46401,N_40633);
nor UO_2361 (O_2361,N_46277,N_47349);
xnor UO_2362 (O_2362,N_43233,N_47534);
or UO_2363 (O_2363,N_48400,N_40360);
nand UO_2364 (O_2364,N_44998,N_40750);
and UO_2365 (O_2365,N_41788,N_48396);
nor UO_2366 (O_2366,N_45925,N_45096);
or UO_2367 (O_2367,N_43792,N_49066);
nand UO_2368 (O_2368,N_42933,N_45982);
xnor UO_2369 (O_2369,N_42965,N_44358);
nand UO_2370 (O_2370,N_49948,N_47762);
nor UO_2371 (O_2371,N_43969,N_40795);
and UO_2372 (O_2372,N_48408,N_47866);
nand UO_2373 (O_2373,N_44009,N_40284);
nand UO_2374 (O_2374,N_42330,N_47472);
xor UO_2375 (O_2375,N_45067,N_40074);
and UO_2376 (O_2376,N_43135,N_45421);
nand UO_2377 (O_2377,N_43208,N_47966);
and UO_2378 (O_2378,N_44352,N_42379);
nor UO_2379 (O_2379,N_40040,N_42869);
xnor UO_2380 (O_2380,N_40848,N_45489);
nand UO_2381 (O_2381,N_48171,N_45540);
nand UO_2382 (O_2382,N_42708,N_42190);
xor UO_2383 (O_2383,N_43765,N_46548);
xor UO_2384 (O_2384,N_45009,N_49836);
or UO_2385 (O_2385,N_43426,N_46845);
nor UO_2386 (O_2386,N_45481,N_40962);
and UO_2387 (O_2387,N_40153,N_45831);
nand UO_2388 (O_2388,N_41071,N_43329);
nand UO_2389 (O_2389,N_49044,N_46208);
nor UO_2390 (O_2390,N_43017,N_43648);
and UO_2391 (O_2391,N_48663,N_46519);
nor UO_2392 (O_2392,N_46223,N_48945);
nand UO_2393 (O_2393,N_48323,N_49521);
xnor UO_2394 (O_2394,N_49435,N_43092);
xnor UO_2395 (O_2395,N_49231,N_48689);
or UO_2396 (O_2396,N_48317,N_41381);
nand UO_2397 (O_2397,N_40462,N_49264);
nand UO_2398 (O_2398,N_46649,N_43490);
xnor UO_2399 (O_2399,N_43189,N_46803);
nand UO_2400 (O_2400,N_49802,N_43538);
and UO_2401 (O_2401,N_45378,N_43622);
xnor UO_2402 (O_2402,N_42471,N_43510);
xor UO_2403 (O_2403,N_40856,N_46303);
or UO_2404 (O_2404,N_49298,N_46028);
nor UO_2405 (O_2405,N_42045,N_45229);
and UO_2406 (O_2406,N_43073,N_47617);
or UO_2407 (O_2407,N_48898,N_47538);
nor UO_2408 (O_2408,N_45590,N_44362);
nand UO_2409 (O_2409,N_41565,N_47683);
nor UO_2410 (O_2410,N_47072,N_41358);
nand UO_2411 (O_2411,N_49052,N_49117);
xnor UO_2412 (O_2412,N_46929,N_40854);
or UO_2413 (O_2413,N_41743,N_47445);
and UO_2414 (O_2414,N_48907,N_42588);
nand UO_2415 (O_2415,N_43029,N_41795);
and UO_2416 (O_2416,N_43910,N_41529);
xnor UO_2417 (O_2417,N_49839,N_40910);
and UO_2418 (O_2418,N_46967,N_42280);
nand UO_2419 (O_2419,N_43575,N_45958);
or UO_2420 (O_2420,N_47710,N_44353);
and UO_2421 (O_2421,N_46356,N_44688);
and UO_2422 (O_2422,N_41409,N_48117);
and UO_2423 (O_2423,N_45531,N_48228);
or UO_2424 (O_2424,N_42722,N_40191);
nor UO_2425 (O_2425,N_43274,N_46622);
and UO_2426 (O_2426,N_43571,N_41087);
or UO_2427 (O_2427,N_42987,N_43784);
and UO_2428 (O_2428,N_41906,N_48776);
or UO_2429 (O_2429,N_43513,N_47451);
nor UO_2430 (O_2430,N_43871,N_47304);
nand UO_2431 (O_2431,N_44286,N_43239);
and UO_2432 (O_2432,N_49991,N_43176);
xor UO_2433 (O_2433,N_41212,N_46199);
nor UO_2434 (O_2434,N_48607,N_48891);
nor UO_2435 (O_2435,N_44198,N_49596);
nand UO_2436 (O_2436,N_48353,N_47199);
nand UO_2437 (O_2437,N_42527,N_49070);
xor UO_2438 (O_2438,N_44210,N_46189);
nor UO_2439 (O_2439,N_49774,N_49636);
nor UO_2440 (O_2440,N_45436,N_45599);
nand UO_2441 (O_2441,N_43776,N_45415);
and UO_2442 (O_2442,N_43096,N_45472);
nand UO_2443 (O_2443,N_41872,N_43822);
nand UO_2444 (O_2444,N_45040,N_44707);
xnor UO_2445 (O_2445,N_48130,N_41308);
nand UO_2446 (O_2446,N_47915,N_42473);
xnor UO_2447 (O_2447,N_46602,N_45562);
nand UO_2448 (O_2448,N_42109,N_41091);
or UO_2449 (O_2449,N_47934,N_49171);
or UO_2450 (O_2450,N_46263,N_43536);
or UO_2451 (O_2451,N_47613,N_42658);
xnor UO_2452 (O_2452,N_45285,N_40914);
or UO_2453 (O_2453,N_41324,N_49895);
nor UO_2454 (O_2454,N_41912,N_48972);
or UO_2455 (O_2455,N_40927,N_49878);
xor UO_2456 (O_2456,N_47032,N_41291);
xor UO_2457 (O_2457,N_42597,N_44393);
nor UO_2458 (O_2458,N_48597,N_44576);
or UO_2459 (O_2459,N_46973,N_41068);
and UO_2460 (O_2460,N_47109,N_44722);
or UO_2461 (O_2461,N_43540,N_45677);
xor UO_2462 (O_2462,N_49265,N_47152);
or UO_2463 (O_2463,N_49239,N_45966);
and UO_2464 (O_2464,N_43919,N_49743);
nor UO_2465 (O_2465,N_42339,N_47456);
and UO_2466 (O_2466,N_48434,N_44664);
or UO_2467 (O_2467,N_49903,N_45610);
nand UO_2468 (O_2468,N_45105,N_47659);
and UO_2469 (O_2469,N_49410,N_48290);
xor UO_2470 (O_2470,N_47370,N_44990);
or UO_2471 (O_2471,N_45171,N_43529);
and UO_2472 (O_2472,N_47404,N_48603);
xnor UO_2473 (O_2473,N_49872,N_45483);
nand UO_2474 (O_2474,N_46638,N_46397);
nor UO_2475 (O_2475,N_41218,N_41507);
nand UO_2476 (O_2476,N_40059,N_48051);
xor UO_2477 (O_2477,N_44236,N_43391);
and UO_2478 (O_2478,N_47627,N_40647);
nand UO_2479 (O_2479,N_48855,N_44702);
nor UO_2480 (O_2480,N_43961,N_44135);
or UO_2481 (O_2481,N_42375,N_42249);
nor UO_2482 (O_2482,N_48297,N_48028);
nor UO_2483 (O_2483,N_42929,N_40777);
or UO_2484 (O_2484,N_44862,N_49844);
nand UO_2485 (O_2485,N_45597,N_46333);
nand UO_2486 (O_2486,N_45444,N_43048);
and UO_2487 (O_2487,N_43140,N_46222);
and UO_2488 (O_2488,N_43340,N_45571);
or UO_2489 (O_2489,N_48817,N_44339);
or UO_2490 (O_2490,N_41131,N_47998);
nand UO_2491 (O_2491,N_49315,N_46076);
xnor UO_2492 (O_2492,N_40312,N_41236);
and UO_2493 (O_2493,N_43989,N_43369);
and UO_2494 (O_2494,N_49456,N_43899);
nand UO_2495 (O_2495,N_41616,N_44473);
nand UO_2496 (O_2496,N_48311,N_43438);
and UO_2497 (O_2497,N_49351,N_40495);
or UO_2498 (O_2498,N_41050,N_40225);
and UO_2499 (O_2499,N_42907,N_46309);
nand UO_2500 (O_2500,N_48724,N_45690);
nor UO_2501 (O_2501,N_42419,N_44803);
and UO_2502 (O_2502,N_43358,N_44881);
nor UO_2503 (O_2503,N_45627,N_46952);
nor UO_2504 (O_2504,N_44411,N_41432);
nor UO_2505 (O_2505,N_47284,N_44622);
nor UO_2506 (O_2506,N_48630,N_49773);
or UO_2507 (O_2507,N_43500,N_43382);
nor UO_2508 (O_2508,N_41712,N_49447);
or UO_2509 (O_2509,N_43196,N_40349);
or UO_2510 (O_2510,N_48557,N_40210);
xnor UO_2511 (O_2511,N_49827,N_41076);
nand UO_2512 (O_2512,N_47080,N_42784);
nand UO_2513 (O_2513,N_41058,N_48594);
and UO_2514 (O_2514,N_43279,N_45945);
xor UO_2515 (O_2515,N_49220,N_44283);
nor UO_2516 (O_2516,N_46504,N_40308);
nand UO_2517 (O_2517,N_46517,N_46960);
or UO_2518 (O_2518,N_43336,N_47333);
and UO_2519 (O_2519,N_43615,N_43617);
nor UO_2520 (O_2520,N_46148,N_41459);
or UO_2521 (O_2521,N_48503,N_44558);
and UO_2522 (O_2522,N_42691,N_48367);
and UO_2523 (O_2523,N_44265,N_40043);
or UO_2524 (O_2524,N_42663,N_45126);
nor UO_2525 (O_2525,N_48874,N_48170);
nor UO_2526 (O_2526,N_46702,N_48872);
nor UO_2527 (O_2527,N_49251,N_44867);
xnor UO_2528 (O_2528,N_47471,N_49189);
and UO_2529 (O_2529,N_42154,N_42318);
nand UO_2530 (O_2530,N_46677,N_45581);
nand UO_2531 (O_2531,N_47246,N_43773);
nor UO_2532 (O_2532,N_49893,N_45072);
nand UO_2533 (O_2533,N_44361,N_40525);
and UO_2534 (O_2534,N_47660,N_41887);
and UO_2535 (O_2535,N_42009,N_42668);
and UO_2536 (O_2536,N_40490,N_46716);
or UO_2537 (O_2537,N_43394,N_46254);
nand UO_2538 (O_2538,N_43008,N_40061);
nand UO_2539 (O_2539,N_44457,N_43762);
and UO_2540 (O_2540,N_43901,N_48153);
and UO_2541 (O_2541,N_42433,N_45327);
or UO_2542 (O_2542,N_40397,N_47460);
nand UO_2543 (O_2543,N_41383,N_41752);
nor UO_2544 (O_2544,N_45897,N_47950);
xor UO_2545 (O_2545,N_47995,N_49232);
nor UO_2546 (O_2546,N_43979,N_43950);
nand UO_2547 (O_2547,N_44888,N_40923);
and UO_2548 (O_2548,N_43456,N_49158);
nand UO_2549 (O_2549,N_42974,N_42635);
or UO_2550 (O_2550,N_46663,N_45801);
nand UO_2551 (O_2551,N_47931,N_44727);
or UO_2552 (O_2552,N_48610,N_44076);
nor UO_2553 (O_2553,N_44613,N_40140);
or UO_2554 (O_2554,N_49656,N_41976);
nor UO_2555 (O_2555,N_41368,N_43701);
nor UO_2556 (O_2556,N_40204,N_46933);
or UO_2557 (O_2557,N_46953,N_41316);
or UO_2558 (O_2558,N_49352,N_44231);
nand UO_2559 (O_2559,N_42614,N_41952);
xor UO_2560 (O_2560,N_47777,N_49695);
nand UO_2561 (O_2561,N_46695,N_46200);
nor UO_2562 (O_2562,N_41653,N_47257);
nand UO_2563 (O_2563,N_45546,N_41097);
nor UO_2564 (O_2564,N_40937,N_41679);
or UO_2565 (O_2565,N_48303,N_43098);
and UO_2566 (O_2566,N_48873,N_41691);
nand UO_2567 (O_2567,N_49344,N_49855);
or UO_2568 (O_2568,N_44239,N_45363);
nand UO_2569 (O_2569,N_49049,N_42026);
nand UO_2570 (O_2570,N_48412,N_44181);
nand UO_2571 (O_2571,N_46986,N_41968);
nor UO_2572 (O_2572,N_41004,N_44405);
xor UO_2573 (O_2573,N_43090,N_43480);
or UO_2574 (O_2574,N_44512,N_44368);
nand UO_2575 (O_2575,N_48143,N_45503);
and UO_2576 (O_2576,N_40173,N_49762);
xor UO_2577 (O_2577,N_43337,N_40209);
nor UO_2578 (O_2578,N_41243,N_44429);
and UO_2579 (O_2579,N_48832,N_46523);
and UO_2580 (O_2580,N_41779,N_40549);
or UO_2581 (O_2581,N_42520,N_48882);
or UO_2582 (O_2582,N_47773,N_41849);
and UO_2583 (O_2583,N_42899,N_41026);
or UO_2584 (O_2584,N_47894,N_40891);
or UO_2585 (O_2585,N_48430,N_42684);
nor UO_2586 (O_2586,N_42921,N_41703);
nor UO_2587 (O_2587,N_43965,N_40296);
xor UO_2588 (O_2588,N_40017,N_43984);
and UO_2589 (O_2589,N_44960,N_40744);
and UO_2590 (O_2590,N_46867,N_45151);
or UO_2591 (O_2591,N_42167,N_46492);
xor UO_2592 (O_2592,N_41762,N_43883);
nor UO_2593 (O_2593,N_49443,N_44983);
and UO_2594 (O_2594,N_49188,N_40287);
and UO_2595 (O_2595,N_45617,N_49379);
or UO_2596 (O_2596,N_45106,N_48483);
xnor UO_2597 (O_2597,N_47050,N_48606);
and UO_2598 (O_2598,N_48292,N_48736);
or UO_2599 (O_2599,N_45152,N_48418);
or UO_2600 (O_2600,N_42232,N_44102);
or UO_2601 (O_2601,N_42512,N_42852);
xor UO_2602 (O_2602,N_46879,N_40182);
nand UO_2603 (O_2603,N_49122,N_42521);
or UO_2604 (O_2604,N_40775,N_42421);
nor UO_2605 (O_2605,N_47884,N_40761);
and UO_2606 (O_2606,N_40057,N_42999);
nor UO_2607 (O_2607,N_49899,N_46621);
nor UO_2608 (O_2608,N_46159,N_48027);
nor UO_2609 (O_2609,N_42654,N_49286);
or UO_2610 (O_2610,N_46251,N_45668);
xor UO_2611 (O_2611,N_40073,N_46207);
nor UO_2612 (O_2612,N_46385,N_45567);
xor UO_2613 (O_2613,N_43341,N_44778);
nand UO_2614 (O_2614,N_48134,N_49620);
nor UO_2615 (O_2615,N_42643,N_41375);
xnor UO_2616 (O_2616,N_48808,N_47689);
and UO_2617 (O_2617,N_45028,N_46043);
nor UO_2618 (O_2618,N_47775,N_46242);
nand UO_2619 (O_2619,N_40535,N_45397);
and UO_2620 (O_2620,N_45034,N_42903);
nor UO_2621 (O_2621,N_40207,N_40773);
nand UO_2622 (O_2622,N_48794,N_41187);
nand UO_2623 (O_2623,N_48846,N_42598);
or UO_2624 (O_2624,N_49957,N_43390);
and UO_2625 (O_2625,N_41400,N_41254);
nand UO_2626 (O_2626,N_49768,N_46240);
nand UO_2627 (O_2627,N_47400,N_42914);
and UO_2628 (O_2628,N_43593,N_40534);
or UO_2629 (O_2629,N_40125,N_43258);
xnor UO_2630 (O_2630,N_48238,N_48837);
and UO_2631 (O_2631,N_41545,N_41842);
and UO_2632 (O_2632,N_45570,N_49244);
nand UO_2633 (O_2633,N_42877,N_42252);
or UO_2634 (O_2634,N_45274,N_45208);
or UO_2635 (O_2635,N_43546,N_48859);
and UO_2636 (O_2636,N_42750,N_46453);
or UO_2637 (O_2637,N_40975,N_45325);
and UO_2638 (O_2638,N_45365,N_48711);
xnor UO_2639 (O_2639,N_48919,N_48294);
xor UO_2640 (O_2640,N_48748,N_44958);
and UO_2641 (O_2641,N_49747,N_42584);
xnor UO_2642 (O_2642,N_47420,N_41911);
and UO_2643 (O_2643,N_46496,N_46672);
and UO_2644 (O_2644,N_49640,N_45375);
or UO_2645 (O_2645,N_49724,N_47645);
and UO_2646 (O_2646,N_41960,N_41654);
nor UO_2647 (O_2647,N_41224,N_43023);
or UO_2648 (O_2648,N_45460,N_49964);
or UO_2649 (O_2649,N_41933,N_43333);
or UO_2650 (O_2650,N_40508,N_44006);
nor UO_2651 (O_2651,N_43339,N_46465);
xor UO_2652 (O_2652,N_46682,N_40666);
and UO_2653 (O_2653,N_47243,N_48823);
xnor UO_2654 (O_2654,N_41946,N_42259);
and UO_2655 (O_2655,N_40427,N_48126);
nand UO_2656 (O_2656,N_48111,N_49285);
nor UO_2657 (O_2657,N_48308,N_40479);
nor UO_2658 (O_2658,N_42224,N_41355);
nand UO_2659 (O_2659,N_47557,N_42185);
and UO_2660 (O_2660,N_49621,N_45536);
and UO_2661 (O_2661,N_46044,N_41311);
nor UO_2662 (O_2662,N_45919,N_48114);
and UO_2663 (O_2663,N_49845,N_44855);
nand UO_2664 (O_2664,N_43719,N_45303);
and UO_2665 (O_2665,N_46618,N_44319);
or UO_2666 (O_2666,N_48324,N_44827);
nor UO_2667 (O_2667,N_42472,N_40814);
nor UO_2668 (O_2668,N_45385,N_42989);
nand UO_2669 (O_2669,N_45246,N_42067);
or UO_2670 (O_2670,N_44276,N_48404);
nand UO_2671 (O_2671,N_40199,N_40252);
nand UO_2672 (O_2672,N_44404,N_49039);
or UO_2673 (O_2673,N_47087,N_47133);
or UO_2674 (O_2674,N_42332,N_48783);
and UO_2675 (O_2675,N_49048,N_46283);
or UO_2676 (O_2676,N_43028,N_48927);
or UO_2677 (O_2677,N_40454,N_46439);
nor UO_2678 (O_2678,N_49717,N_41166);
nand UO_2679 (O_2679,N_46402,N_41777);
or UO_2680 (O_2680,N_42650,N_43717);
nand UO_2681 (O_2681,N_42424,N_41768);
nor UO_2682 (O_2682,N_46035,N_45777);
and UO_2683 (O_2683,N_46728,N_43952);
nor UO_2684 (O_2684,N_48875,N_43220);
or UO_2685 (O_2685,N_46773,N_47062);
nand UO_2686 (O_2686,N_43645,N_41846);
or UO_2687 (O_2687,N_44434,N_47034);
xnor UO_2688 (O_2688,N_48542,N_41268);
nand UO_2689 (O_2689,N_44328,N_40442);
or UO_2690 (O_2690,N_43267,N_46226);
xor UO_2691 (O_2691,N_40138,N_45901);
nand UO_2692 (O_2692,N_43259,N_49197);
xnor UO_2693 (O_2693,N_42886,N_44648);
and UO_2694 (O_2694,N_47081,N_49837);
nor UO_2695 (O_2695,N_46011,N_40843);
and UO_2696 (O_2696,N_43881,N_46606);
nor UO_2697 (O_2697,N_43646,N_43505);
nand UO_2698 (O_2698,N_40747,N_44591);
xnor UO_2699 (O_2699,N_43145,N_45252);
or UO_2700 (O_2700,N_43614,N_40996);
nand UO_2701 (O_2701,N_40567,N_48671);
or UO_2702 (O_2702,N_43385,N_40677);
and UO_2703 (O_2703,N_45328,N_48242);
and UO_2704 (O_2704,N_42892,N_41466);
and UO_2705 (O_2705,N_46546,N_45078);
xnor UO_2706 (O_2706,N_48152,N_45108);
or UO_2707 (O_2707,N_41750,N_44047);
and UO_2708 (O_2708,N_42680,N_44748);
nand UO_2709 (O_2709,N_41641,N_41696);
xor UO_2710 (O_2710,N_43319,N_45987);
xnor UO_2711 (O_2711,N_47215,N_40877);
or UO_2712 (O_2712,N_45487,N_43046);
or UO_2713 (O_2713,N_45697,N_48570);
nand UO_2714 (O_2714,N_42150,N_43932);
xor UO_2715 (O_2715,N_48376,N_42976);
and UO_2716 (O_2716,N_42133,N_47605);
nor UO_2717 (O_2717,N_47840,N_43996);
and UO_2718 (O_2718,N_40194,N_49566);
nand UO_2719 (O_2719,N_44221,N_48384);
or UO_2720 (O_2720,N_47852,N_47980);
and UO_2721 (O_2721,N_42409,N_40053);
or UO_2722 (O_2722,N_47493,N_42100);
nor UO_2723 (O_2723,N_44571,N_45519);
nor UO_2724 (O_2724,N_41727,N_48053);
or UO_2725 (O_2725,N_48383,N_49005);
and UO_2726 (O_2726,N_47831,N_46435);
nand UO_2727 (O_2727,N_45983,N_44459);
or UO_2728 (O_2728,N_46287,N_40291);
or UO_2729 (O_2729,N_42228,N_43099);
nand UO_2730 (O_2730,N_49829,N_43697);
or UO_2731 (O_2731,N_41711,N_40310);
xor UO_2732 (O_2732,N_45812,N_46705);
xnor UO_2733 (O_2733,N_45577,N_46657);
nor UO_2734 (O_2734,N_42895,N_46394);
and UO_2735 (O_2735,N_49532,N_47056);
nor UO_2736 (O_2736,N_43789,N_44971);
nand UO_2737 (O_2737,N_49460,N_48024);
or UO_2738 (O_2738,N_44233,N_41541);
nand UO_2739 (O_2739,N_44246,N_41618);
nand UO_2740 (O_2740,N_43249,N_41257);
nor UO_2741 (O_2741,N_44129,N_42766);
xor UO_2742 (O_2742,N_40702,N_41824);
xnor UO_2743 (O_2743,N_47741,N_40484);
and UO_2744 (O_2744,N_44797,N_41839);
xor UO_2745 (O_2745,N_49575,N_46736);
or UO_2746 (O_2746,N_46112,N_48639);
nand UO_2747 (O_2747,N_42161,N_45672);
xor UO_2748 (O_2748,N_44723,N_46408);
and UO_2749 (O_2749,N_46642,N_41095);
and UO_2750 (O_2750,N_40237,N_47147);
nand UO_2751 (O_2751,N_42400,N_43801);
nand UO_2752 (O_2752,N_42953,N_43348);
nor UO_2753 (O_2753,N_45928,N_42553);
xor UO_2754 (O_2754,N_42068,N_43014);
or UO_2755 (O_2755,N_41489,N_47142);
and UO_2756 (O_2756,N_40275,N_40576);
nand UO_2757 (O_2757,N_47746,N_44963);
or UO_2758 (O_2758,N_49604,N_43263);
or UO_2759 (O_2759,N_45164,N_46812);
and UO_2760 (O_2760,N_46566,N_48346);
or UO_2761 (O_2761,N_41306,N_42241);
and UO_2762 (O_2762,N_44628,N_45652);
xnor UO_2763 (O_2763,N_49175,N_42523);
xor UO_2764 (O_2764,N_48319,N_44305);
nand UO_2765 (O_2765,N_47279,N_45318);
xnor UO_2766 (O_2766,N_41219,N_40418);
nor UO_2767 (O_2767,N_43644,N_42369);
and UO_2768 (O_2768,N_47219,N_43620);
nor UO_2769 (O_2769,N_46530,N_47308);
and UO_2770 (O_2770,N_43433,N_44310);
nor UO_2771 (O_2771,N_41573,N_42857);
or UO_2772 (O_2772,N_46660,N_47091);
nand UO_2773 (O_2773,N_42202,N_47479);
xnor UO_2774 (O_2774,N_48082,N_46653);
nand UO_2775 (O_2775,N_45701,N_48097);
nand UO_2776 (O_2776,N_43618,N_49416);
nand UO_2777 (O_2777,N_43120,N_48568);
or UO_2778 (O_2778,N_43756,N_49176);
nand UO_2779 (O_2779,N_41736,N_42748);
and UO_2780 (O_2780,N_44595,N_47356);
xnor UO_2781 (O_2781,N_44228,N_42711);
xnor UO_2782 (O_2782,N_45868,N_41054);
xor UO_2783 (O_2783,N_44997,N_42153);
or UO_2784 (O_2784,N_45055,N_46920);
and UO_2785 (O_2785,N_44828,N_49278);
and UO_2786 (O_2786,N_47301,N_41715);
nor UO_2787 (O_2787,N_49776,N_41681);
xnor UO_2788 (O_2788,N_49858,N_46275);
nand UO_2789 (O_2789,N_43624,N_42023);
xor UO_2790 (O_2790,N_41614,N_41247);
xor UO_2791 (O_2791,N_47482,N_47519);
or UO_2792 (O_2792,N_40133,N_49814);
nor UO_2793 (O_2793,N_45214,N_44999);
xor UO_2794 (O_2794,N_40027,N_42876);
xor UO_2795 (O_2795,N_46215,N_40167);
and UO_2796 (O_2796,N_48987,N_43600);
xnor UO_2797 (O_2797,N_46932,N_44107);
and UO_2798 (O_2798,N_43199,N_43745);
or UO_2799 (O_2799,N_47377,N_43922);
xnor UO_2800 (O_2800,N_42476,N_49766);
nor UO_2801 (O_2801,N_42812,N_46156);
nor UO_2802 (O_2802,N_45992,N_45826);
nor UO_2803 (O_2803,N_42884,N_47470);
nand UO_2804 (O_2804,N_45160,N_45973);
and UO_2805 (O_2805,N_40274,N_41883);
and UO_2806 (O_2806,N_49036,N_45224);
nor UO_2807 (O_2807,N_46851,N_43698);
nand UO_2808 (O_2808,N_47430,N_48373);
and UO_2809 (O_2809,N_42586,N_48562);
and UO_2810 (O_2810,N_43072,N_44573);
xnor UO_2811 (O_2811,N_41270,N_48251);
nor UO_2812 (O_2812,N_42459,N_46289);
or UO_2813 (O_2813,N_45584,N_43577);
xnor UO_2814 (O_2814,N_41817,N_47721);
and UO_2815 (O_2815,N_45310,N_45989);
nand UO_2816 (O_2816,N_47841,N_47322);
nor UO_2817 (O_2817,N_46110,N_49909);
or UO_2818 (O_2818,N_46675,N_41938);
nor UO_2819 (O_2819,N_43649,N_45008);
or UO_2820 (O_2820,N_42661,N_46711);
nor UO_2821 (O_2821,N_43667,N_43651);
xor UO_2822 (O_2822,N_48354,N_48527);
and UO_2823 (O_2823,N_48992,N_45785);
and UO_2824 (O_2824,N_41193,N_43815);
and UO_2825 (O_2825,N_49792,N_46308);
nand UO_2826 (O_2826,N_49694,N_47837);
nor UO_2827 (O_2827,N_43109,N_45558);
nor UO_2828 (O_2828,N_41815,N_45264);
or UO_2829 (O_2829,N_49779,N_44367);
nor UO_2830 (O_2830,N_44065,N_43923);
nor UO_2831 (O_2831,N_42220,N_45761);
or UO_2832 (O_2832,N_41313,N_40705);
nor UO_2833 (O_2833,N_45856,N_46357);
nand UO_2834 (O_2834,N_46804,N_42053);
nor UO_2835 (O_2835,N_45392,N_44739);
nand UO_2836 (O_2836,N_49846,N_46789);
xor UO_2837 (O_2837,N_45976,N_41587);
nand UO_2838 (O_2838,N_43539,N_43356);
xor UO_2839 (O_2839,N_44821,N_46172);
xnor UO_2840 (O_2840,N_40862,N_49689);
or UO_2841 (O_2841,N_44766,N_49266);
and UO_2842 (O_2842,N_48678,N_46243);
and UO_2843 (O_2843,N_46758,N_43978);
nand UO_2844 (O_2844,N_40796,N_49503);
nor UO_2845 (O_2845,N_48271,N_43155);
and UO_2846 (O_2846,N_41993,N_45800);
nor UO_2847 (O_2847,N_44456,N_47715);
or UO_2848 (O_2848,N_48737,N_48713);
or UO_2849 (O_2849,N_41127,N_47882);
and UO_2850 (O_2850,N_46325,N_46568);
nor UO_2851 (O_2851,N_46842,N_47750);
nand UO_2852 (O_2852,N_41604,N_47986);
nand UO_2853 (O_2853,N_42576,N_42407);
nand UO_2854 (O_2854,N_48673,N_43833);
nor UO_2855 (O_2855,N_47410,N_49933);
nor UO_2856 (O_2856,N_40406,N_46097);
nand UO_2857 (O_2857,N_46786,N_45373);
and UO_2858 (O_2858,N_42698,N_48864);
and UO_2859 (O_2859,N_44194,N_43446);
nand UO_2860 (O_2860,N_42105,N_41907);
nand UO_2861 (O_2861,N_43805,N_48256);
xnor UO_2862 (O_2862,N_40845,N_44130);
nand UO_2863 (O_2863,N_41233,N_45114);
or UO_2864 (O_2864,N_45359,N_49462);
nand UO_2865 (O_2865,N_44988,N_41559);
and UO_2866 (O_2866,N_43443,N_41171);
or UO_2867 (O_2867,N_43460,N_45128);
and UO_2868 (O_2868,N_40624,N_45374);
or UO_2869 (O_2869,N_42127,N_48935);
xnor UO_2870 (O_2870,N_42679,N_40314);
nand UO_2871 (O_2871,N_42864,N_40326);
nand UO_2872 (O_2872,N_41589,N_42503);
or UO_2873 (O_2873,N_41882,N_40716);
and UO_2874 (O_2874,N_45615,N_48569);
nand UO_2875 (O_2875,N_49522,N_46963);
nor UO_2876 (O_2876,N_44751,N_46643);
or UO_2877 (O_2877,N_49881,N_46718);
and UO_2878 (O_2878,N_48769,N_49728);
and UO_2879 (O_2879,N_41148,N_42660);
xor UO_2880 (O_2880,N_46024,N_44099);
xnor UO_2881 (O_2881,N_40433,N_42403);
nand UO_2882 (O_2882,N_47580,N_42349);
xnor UO_2883 (O_2883,N_43559,N_46318);
nand UO_2884 (O_2884,N_49537,N_48758);
or UO_2885 (O_2885,N_43108,N_48381);
xnor UO_2886 (O_2886,N_46224,N_40517);
nor UO_2887 (O_2887,N_45555,N_45642);
xnor UO_2888 (O_2888,N_47353,N_40564);
nand UO_2889 (O_2889,N_46295,N_49797);
nor UO_2890 (O_2890,N_44643,N_42823);
nor UO_2891 (O_2891,N_45905,N_40366);
and UO_2892 (O_2892,N_41792,N_40398);
nor UO_2893 (O_2893,N_40339,N_48013);
nand UO_2894 (O_2894,N_47235,N_49648);
nor UO_2895 (O_2895,N_41863,N_43367);
and UO_2896 (O_2896,N_47230,N_47477);
or UO_2897 (O_2897,N_44912,N_46124);
nand UO_2898 (O_2898,N_49261,N_41630);
or UO_2899 (O_2899,N_47981,N_40410);
nor UO_2900 (O_2900,N_42552,N_40857);
nand UO_2901 (O_2901,N_47450,N_48704);
and UO_2902 (O_2902,N_42807,N_49740);
nor UO_2903 (O_2903,N_42137,N_45176);
or UO_2904 (O_2904,N_47547,N_48374);
or UO_2905 (O_2905,N_46820,N_40377);
nand UO_2906 (O_2906,N_40916,N_49915);
xnor UO_2907 (O_2907,N_46717,N_41228);
or UO_2908 (O_2908,N_46654,N_47726);
xnor UO_2909 (O_2909,N_42798,N_47339);
nand UO_2910 (O_2910,N_44440,N_44831);
and UO_2911 (O_2911,N_45342,N_49106);
nor UO_2912 (O_2912,N_41129,N_42366);
nand UO_2913 (O_2913,N_45278,N_47584);
or UO_2914 (O_2914,N_44372,N_44284);
xnor UO_2915 (O_2915,N_43769,N_40655);
nor UO_2916 (O_2916,N_47059,N_47952);
or UO_2917 (O_2917,N_43826,N_41979);
and UO_2918 (O_2918,N_47418,N_49758);
xor UO_2919 (O_2919,N_40934,N_48288);
xnor UO_2920 (O_2920,N_47170,N_47714);
or UO_2921 (O_2921,N_47821,N_48571);
and UO_2922 (O_2922,N_41905,N_46469);
nor UO_2923 (O_2923,N_43038,N_46306);
nand UO_2924 (O_2924,N_46260,N_47751);
nand UO_2925 (O_2925,N_41771,N_49243);
xor UO_2926 (O_2926,N_47468,N_49544);
and UO_2927 (O_2927,N_49516,N_49354);
and UO_2928 (O_2928,N_46137,N_42916);
and UO_2929 (O_2929,N_49876,N_46426);
and UO_2930 (O_2930,N_43452,N_48276);
and UO_2931 (O_2931,N_45594,N_46463);
xor UO_2932 (O_2932,N_45383,N_47146);
or UO_2933 (O_2933,N_48092,N_43364);
or UO_2934 (O_2934,N_41932,N_41532);
and UO_2935 (O_2935,N_40935,N_40156);
xnor UO_2936 (O_2936,N_43512,N_44996);
or UO_2937 (O_2937,N_46468,N_43060);
nor UO_2938 (O_2938,N_43968,N_48017);
xor UO_2939 (O_2939,N_47568,N_40405);
xor UO_2940 (O_2940,N_47249,N_46364);
nor UO_2941 (O_2941,N_49428,N_40774);
xnor UO_2942 (O_2942,N_46613,N_49786);
nand UO_2943 (O_2943,N_45037,N_47025);
xnor UO_2944 (O_2944,N_44038,N_49938);
or UO_2945 (O_2945,N_48843,N_40116);
xnor UO_2946 (O_2946,N_49753,N_48994);
nand UO_2947 (O_2947,N_47306,N_47073);
and UO_2948 (O_2948,N_44145,N_41581);
and UO_2949 (O_2949,N_44278,N_48078);
and UO_2950 (O_2950,N_40035,N_46078);
and UO_2951 (O_2951,N_47313,N_44661);
nand UO_2952 (O_2952,N_47161,N_42163);
nand UO_2953 (O_2953,N_47869,N_45121);
nor UO_2954 (O_2954,N_40597,N_49982);
and UO_2955 (O_2955,N_48910,N_41610);
nor UO_2956 (O_2956,N_47122,N_46324);
nand UO_2957 (O_2957,N_47799,N_41003);
nor UO_2958 (O_2958,N_47098,N_45210);
and UO_2959 (O_2959,N_47319,N_49426);
xor UO_2960 (O_2960,N_45170,N_47218);
xnor UO_2961 (O_2961,N_40285,N_44143);
xnor UO_2962 (O_2962,N_43481,N_49587);
xnor UO_2963 (O_2963,N_43303,N_47417);
xor UO_2964 (O_2964,N_46036,N_46678);
and UO_2965 (O_2965,N_44054,N_41083);
and UO_2966 (O_2966,N_48980,N_44426);
xnor UO_2967 (O_2967,N_41180,N_48800);
nand UO_2968 (O_2968,N_43581,N_42882);
nand UO_2969 (O_2969,N_44336,N_41687);
xor UO_2970 (O_2970,N_45538,N_41930);
and UO_2971 (O_2971,N_45695,N_46796);
and UO_2972 (O_2972,N_47624,N_43188);
xor UO_2973 (O_2973,N_41346,N_48257);
xnor UO_2974 (O_2974,N_44180,N_45566);
nor UO_2975 (O_2975,N_44066,N_45396);
xnor UO_2976 (O_2976,N_40717,N_42915);
and UO_2977 (O_2977,N_49126,N_47530);
or UO_2978 (O_2978,N_47455,N_45038);
nor UO_2979 (O_2979,N_45788,N_44615);
xnor UO_2980 (O_2980,N_44843,N_47022);
nand UO_2981 (O_2981,N_49481,N_49700);
nor UO_2982 (O_2982,N_47446,N_41591);
and UO_2983 (O_2983,N_48244,N_42634);
xnor UO_2984 (O_2984,N_41540,N_43487);
nand UO_2985 (O_2985,N_47606,N_41931);
and UO_2986 (O_2986,N_44159,N_44462);
nand UO_2987 (O_2987,N_40571,N_46844);
nor UO_2988 (O_2988,N_46142,N_44307);
xor UO_2989 (O_2989,N_40362,N_42397);
xor UO_2990 (O_2990,N_41283,N_43305);
xor UO_2991 (O_2991,N_43195,N_45713);
nand UO_2992 (O_2992,N_47523,N_45646);
and UO_2993 (O_2993,N_44132,N_48632);
xor UO_2994 (O_2994,N_48887,N_42066);
nand UO_2995 (O_2995,N_42964,N_46570);
nand UO_2996 (O_2996,N_41122,N_44936);
xnor UO_2997 (O_2997,N_49152,N_46212);
and UO_2998 (O_2998,N_44472,N_43057);
xor UO_2999 (O_2999,N_45159,N_42843);
and UO_3000 (O_3000,N_42594,N_49071);
nand UO_3001 (O_3001,N_42815,N_47168);
nor UO_3002 (O_3002,N_41709,N_44074);
nor UO_3003 (O_3003,N_47440,N_49129);
nand UO_3004 (O_3004,N_40965,N_42992);
or UO_3005 (O_3005,N_48090,N_40422);
nor UO_3006 (O_3006,N_43895,N_42765);
nand UO_3007 (O_3007,N_48895,N_48771);
or UO_3008 (O_3008,N_40055,N_49383);
or UO_3009 (O_3009,N_48973,N_45269);
nand UO_3010 (O_3010,N_49105,N_43640);
and UO_3011 (O_3011,N_45116,N_40248);
nor UO_3012 (O_3012,N_49939,N_43797);
and UO_3013 (O_3013,N_46813,N_43555);
and UO_3014 (O_3014,N_48372,N_45794);
xor UO_3015 (O_3015,N_40344,N_40683);
and UO_3016 (O_3016,N_44585,N_44083);
nand UO_3017 (O_3017,N_49469,N_49027);
and UO_3018 (O_3018,N_46412,N_41741);
nand UO_3019 (O_3019,N_44370,N_49086);
nor UO_3020 (O_3020,N_43343,N_43054);
nand UO_3021 (O_3021,N_48389,N_43024);
and UO_3022 (O_3022,N_40333,N_46891);
nand UO_3023 (O_3023,N_45271,N_45423);
or UO_3024 (O_3024,N_48213,N_46125);
nand UO_3025 (O_3025,N_44640,N_42922);
or UO_3026 (O_3026,N_45728,N_44325);
or UO_3027 (O_3027,N_48380,N_47586);
xnor UO_3028 (O_3028,N_42442,N_48336);
and UO_3029 (O_3029,N_47629,N_48640);
xor UO_3030 (O_3030,N_48291,N_48963);
nand UO_3031 (O_3031,N_43080,N_49504);
nand UO_3032 (O_3032,N_46565,N_49463);
xor UO_3033 (O_3033,N_48660,N_40370);
nor UO_3034 (O_3034,N_46680,N_45542);
and UO_3035 (O_3035,N_46464,N_42605);
xnor UO_3036 (O_3036,N_40328,N_43261);
xor UO_3037 (O_3037,N_47019,N_45475);
xor UO_3038 (O_3038,N_46913,N_48954);
or UO_3039 (O_3039,N_48647,N_41525);
nor UO_3040 (O_3040,N_48779,N_40870);
nor UO_3041 (O_3041,N_40649,N_42847);
and UO_3042 (O_3042,N_46846,N_47749);
xnor UO_3043 (O_3043,N_48501,N_49485);
nor UO_3044 (O_3044,N_42342,N_44522);
xnor UO_3045 (O_3045,N_42110,N_46670);
nor UO_3046 (O_3046,N_47758,N_46688);
nor UO_3047 (O_3047,N_41062,N_48645);
nand UO_3048 (O_3048,N_43299,N_41729);
or UO_3049 (O_3049,N_46007,N_46396);
and UO_3050 (O_3050,N_47823,N_47224);
nand UO_3051 (O_3051,N_40114,N_47850);
nor UO_3052 (O_3052,N_46320,N_43384);
or UO_3053 (O_3053,N_44665,N_42461);
nor UO_3054 (O_3054,N_48212,N_49992);
xor UO_3055 (O_3055,N_45486,N_45054);
or UO_3056 (O_3056,N_49749,N_47398);
or UO_3057 (O_3057,N_45505,N_43022);
nor UO_3058 (O_3058,N_47309,N_49672);
nor UO_3059 (O_3059,N_46673,N_47560);
xnor UO_3060 (O_3060,N_48065,N_48364);
nor UO_3061 (O_3061,N_45052,N_47669);
nor UO_3062 (O_3062,N_48466,N_48349);
or UO_3063 (O_3063,N_46236,N_42244);
nor UO_3064 (O_3064,N_46082,N_47447);
nor UO_3065 (O_3065,N_42874,N_45109);
nand UO_3066 (O_3066,N_47029,N_48780);
or UO_3067 (O_3067,N_47517,N_44938);
and UO_3068 (O_3068,N_40180,N_47149);
or UO_3069 (O_3069,N_49124,N_40811);
nor UO_3070 (O_3070,N_49421,N_41039);
nand UO_3071 (O_3071,N_44824,N_44921);
nand UO_3072 (O_3072,N_40494,N_45473);
xor UO_3073 (O_3073,N_43206,N_45228);
nand UO_3074 (O_3074,N_40161,N_44270);
and UO_3075 (O_3075,N_40146,N_47548);
and UO_3076 (O_3076,N_47763,N_45884);
nand UO_3077 (O_3077,N_41498,N_40062);
nand UO_3078 (O_3078,N_47987,N_48592);
nand UO_3079 (O_3079,N_47206,N_44584);
or UO_3080 (O_3080,N_40177,N_45353);
nor UO_3081 (O_3081,N_42749,N_46855);
or UO_3082 (O_3082,N_40792,N_41376);
xor UO_3083 (O_3083,N_43696,N_41176);
or UO_3084 (O_3084,N_45003,N_40048);
and UO_3085 (O_3085,N_49015,N_44668);
nand UO_3086 (O_3086,N_41675,N_42970);
nand UO_3087 (O_3087,N_46708,N_46383);
or UO_3088 (O_3088,N_45215,N_45188);
nand UO_3089 (O_3089,N_46127,N_46456);
nor UO_3090 (O_3090,N_45941,N_48159);
or UO_3091 (O_3091,N_44818,N_43380);
or UO_3092 (O_3092,N_44439,N_44597);
nor UO_3093 (O_3093,N_44206,N_41182);
nor UO_3094 (O_3094,N_46373,N_49929);
nand UO_3095 (O_3095,N_43050,N_42377);
xor UO_3096 (O_3096,N_48583,N_49465);
nor UO_3097 (O_3097,N_45909,N_48703);
and UO_3098 (O_3098,N_49021,N_49514);
nor UO_3099 (O_3099,N_48009,N_43723);
nor UO_3100 (O_3100,N_47501,N_42919);
and UO_3101 (O_3101,N_46120,N_41106);
and UO_3102 (O_3102,N_46077,N_41823);
xnor UO_3103 (O_3103,N_43908,N_40473);
and UO_3104 (O_3104,N_49350,N_40596);
and UO_3105 (O_3105,N_40986,N_43689);
and UO_3106 (O_3106,N_47954,N_44497);
or UO_3107 (O_3107,N_46046,N_40389);
nand UO_3108 (O_3108,N_45931,N_48611);
or UO_3109 (O_3109,N_41197,N_47524);
and UO_3110 (O_3110,N_41203,N_47559);
and UO_3111 (O_3111,N_49625,N_40246);
or UO_3112 (O_3112,N_40537,N_41974);
xor UO_3113 (O_3113,N_41025,N_41935);
nand UO_3114 (O_3114,N_41423,N_40790);
xnor UO_3115 (O_3115,N_41086,N_40487);
nand UO_3116 (O_3116,N_48730,N_44891);
nor UO_3117 (O_3117,N_40955,N_42781);
or UO_3118 (O_3118,N_41786,N_48285);
nand UO_3119 (O_3119,N_40813,N_45372);
or UO_3120 (O_3120,N_42537,N_45549);
or UO_3121 (O_3121,N_40723,N_43985);
xor UO_3122 (O_3122,N_47812,N_48498);
and UO_3123 (O_3123,N_46228,N_40013);
and UO_3124 (O_3124,N_49598,N_42996);
and UO_3125 (O_3125,N_40342,N_49257);
or UO_3126 (O_3126,N_43741,N_46134);
nor UO_3127 (O_3127,N_47975,N_45804);
or UO_3128 (O_3128,N_41758,N_40115);
and UO_3129 (O_3129,N_49919,N_42292);
and UO_3130 (O_3130,N_47241,N_49714);
xnor UO_3131 (O_3131,N_44705,N_41061);
xnor UO_3132 (O_3132,N_48091,N_48765);
nand UO_3133 (O_3133,N_47511,N_45453);
nand UO_3134 (O_3134,N_47919,N_49509);
or UO_3135 (O_3135,N_46403,N_47590);
xor UO_3136 (O_3136,N_42619,N_47083);
nor UO_3137 (O_3137,N_44050,N_42814);
or UO_3138 (O_3138,N_44572,N_48385);
nor UO_3139 (O_3139,N_48147,N_44464);
nor UO_3140 (O_3140,N_49348,N_48585);
nor UO_3141 (O_3141,N_49337,N_40828);
xor UO_3142 (O_3142,N_49627,N_49611);
xnor UO_3143 (O_3143,N_49862,N_49472);
nand UO_3144 (O_3144,N_49812,N_43811);
nand UO_3145 (O_3145,N_48714,N_45331);
and UO_3146 (O_3146,N_47892,N_43795);
or UO_3147 (O_3147,N_45449,N_47186);
xnor UO_3148 (O_3148,N_40028,N_49000);
xnor UO_3149 (O_3149,N_44973,N_42540);
and UO_3150 (O_3150,N_47713,N_47776);
xor UO_3151 (O_3151,N_44747,N_45543);
xnor UO_3152 (O_3152,N_40426,N_40933);
nand UO_3153 (O_3153,N_41811,N_46001);
or UO_3154 (O_3154,N_47203,N_43913);
and UO_3155 (O_3155,N_45239,N_42878);
or UO_3156 (O_3156,N_49372,N_40769);
nand UO_3157 (O_3157,N_45060,N_42256);
nor UO_3158 (O_3158,N_45377,N_42038);
xor UO_3159 (O_3159,N_42667,N_45077);
nor UO_3160 (O_3160,N_44403,N_44965);
and UO_3161 (O_3161,N_45474,N_43231);
and UO_3162 (O_3162,N_45139,N_45758);
nand UO_3163 (O_3163,N_41598,N_43839);
nor UO_3164 (O_3164,N_49798,N_49401);
xor UO_3165 (O_3165,N_44317,N_42937);
nor UO_3166 (O_3166,N_45402,N_41737);
and UO_3167 (O_3167,N_49607,N_44503);
xnor UO_3168 (O_3168,N_46659,N_43378);
and UO_3169 (O_3169,N_48173,N_46805);
nand UO_3170 (O_3170,N_47704,N_46000);
and UO_3171 (O_3171,N_44489,N_43227);
xor UO_3172 (O_3172,N_43506,N_45058);
nand UO_3173 (O_3173,N_49042,N_46056);
nor UO_3174 (O_3174,N_46219,N_46458);
nand UO_3175 (O_3175,N_46756,N_40545);
and UO_3176 (O_3176,N_47274,N_45050);
xnor UO_3177 (O_3177,N_45276,N_40122);
or UO_3178 (O_3178,N_45349,N_43652);
nand UO_3179 (O_3179,N_47856,N_42647);
xnor UO_3180 (O_3180,N_40332,N_44894);
xor UO_3181 (O_3181,N_44031,N_45462);
xnor UO_3182 (O_3182,N_47324,N_47874);
xnor UO_3183 (O_3183,N_40741,N_49332);
and UO_3184 (O_3184,N_43449,N_45192);
or UO_3185 (O_3185,N_47239,N_42335);
or UO_3186 (O_3186,N_41454,N_46877);
xor UO_3187 (O_3187,N_49630,N_41300);
xor UO_3188 (O_3188,N_47453,N_47185);
and UO_3189 (O_3189,N_42695,N_41975);
nor UO_3190 (O_3190,N_44865,N_47525);
nand UO_3191 (O_3191,N_47040,N_45272);
or UO_3192 (O_3192,N_43283,N_41305);
xor UO_3193 (O_3193,N_40911,N_40957);
nor UO_3194 (O_3194,N_46808,N_42037);
and UO_3195 (O_3195,N_46662,N_45878);
and UO_3196 (O_3196,N_47003,N_44749);
nand UO_3197 (O_3197,N_49342,N_42354);
and UO_3198 (O_3198,N_49033,N_46249);
xnor UO_3199 (O_3199,N_41640,N_49918);
and UO_3200 (O_3200,N_42325,N_45456);
or UO_3201 (O_3201,N_45001,N_46916);
xnor UO_3202 (O_3202,N_42022,N_42997);
xor UO_3203 (O_3203,N_46490,N_40203);
xnor UO_3204 (O_3204,N_45887,N_43065);
xnor UO_3205 (O_3205,N_46304,N_47058);
or UO_3206 (O_3206,N_43678,N_49571);
xnor UO_3207 (O_3207,N_41868,N_48214);
and UO_3208 (O_3208,N_40918,N_40143);
and UO_3209 (O_3209,N_43353,N_49058);
and UO_3210 (O_3210,N_45523,N_42793);
or UO_3211 (O_3211,N_46830,N_40988);
xor UO_3212 (O_3212,N_48614,N_47811);
xnor UO_3213 (O_3213,N_47125,N_43331);
nand UO_3214 (O_3214,N_48422,N_40323);
or UO_3215 (O_3215,N_41259,N_45350);
and UO_3216 (O_3216,N_46290,N_45608);
or UO_3217 (O_3217,N_42778,N_40520);
xor UO_3218 (O_3218,N_49931,N_43612);
nand UO_3219 (O_3219,N_40330,N_45455);
or UO_3220 (O_3220,N_45696,N_49470);
and UO_3221 (O_3221,N_44450,N_45307);
and UO_3222 (O_3222,N_41439,N_40885);
or UO_3223 (O_3223,N_41462,N_49811);
xor UO_3224 (O_3224,N_42120,N_41296);
and UO_3225 (O_3225,N_47288,N_45660);
nor UO_3226 (O_3226,N_40764,N_41981);
xor UO_3227 (O_3227,N_41344,N_41512);
or UO_3228 (O_3228,N_45755,N_41126);
or UO_3229 (O_3229,N_46921,N_43796);
nor UO_3230 (O_3230,N_45671,N_45656);
xor UO_3231 (O_3231,N_49206,N_42322);
xor UO_3232 (O_3232,N_40945,N_47844);
and UO_3233 (O_3233,N_45655,N_41723);
and UO_3234 (O_3234,N_47838,N_46797);
or UO_3235 (O_3235,N_44663,N_43843);
xnor UO_3236 (O_3236,N_41413,N_40890);
xor UO_3237 (O_3237,N_45734,N_48893);
and UO_3238 (O_3238,N_42825,N_47674);
xor UO_3239 (O_3239,N_45962,N_45533);
and UO_3240 (O_3240,N_42526,N_45371);
xnor UO_3241 (O_3241,N_47829,N_45235);
nor UO_3242 (O_3242,N_49222,N_47598);
xnor UO_3243 (O_3243,N_46405,N_47815);
nand UO_3244 (O_3244,N_49794,N_46866);
nand UO_3245 (O_3245,N_42905,N_46559);
or UO_3246 (O_3246,N_44694,N_43642);
or UO_3247 (O_3247,N_42490,N_48492);
or UO_3248 (O_3248,N_45764,N_42329);
nor UO_3249 (O_3249,N_42229,N_49674);
nor UO_3250 (O_3250,N_47116,N_48160);
and UO_3251 (O_3251,N_49098,N_44691);
nor UO_3252 (O_3252,N_49132,N_47171);
or UO_3253 (O_3253,N_47858,N_40443);
xnor UO_3254 (O_3254,N_46700,N_45168);
and UO_3255 (O_3255,N_47824,N_47805);
and UO_3256 (O_3256,N_47434,N_44586);
nand UO_3257 (O_3257,N_41720,N_42076);
and UO_3258 (O_3258,N_41234,N_44444);
and UO_3259 (O_3259,N_45517,N_47208);
nor UO_3260 (O_3260,N_49392,N_40288);
or UO_3261 (O_3261,N_46579,N_48889);
and UO_3262 (O_3262,N_48796,N_40733);
nor UO_3263 (O_3263,N_42013,N_49449);
or UO_3264 (O_3264,N_44507,N_48738);
nand UO_3265 (O_3265,N_40574,N_48879);
or UO_3266 (O_3266,N_44167,N_41336);
or UO_3267 (O_3267,N_46181,N_42821);
and UO_3268 (O_3268,N_47814,N_46297);
and UO_3269 (O_3269,N_45740,N_47543);
nand UO_3270 (O_3270,N_40045,N_46080);
or UO_3271 (O_3271,N_48119,N_48750);
or UO_3272 (O_3272,N_45544,N_46334);
or UO_3273 (O_3273,N_43799,N_48435);
nor UO_3274 (O_3274,N_40316,N_45914);
nor UO_3275 (O_3275,N_46720,N_43212);
nor UO_3276 (O_3276,N_46389,N_49491);
nand UO_3277 (O_3277,N_46671,N_45957);
and UO_3278 (O_3278,N_47251,N_42404);
nor UO_3279 (O_3279,N_48681,N_42033);
or UO_3280 (O_3280,N_41755,N_40187);
xnor UO_3281 (O_3281,N_48469,N_45611);
nand UO_3282 (O_3282,N_40570,N_48139);
or UO_3283 (O_3283,N_40675,N_42357);
xor UO_3284 (O_3284,N_48920,N_41482);
and UO_3285 (O_3285,N_49397,N_46774);
and UO_3286 (O_3286,N_40731,N_44520);
xor UO_3287 (O_3287,N_46030,N_48558);
nor UO_3288 (O_3288,N_49880,N_40821);
nand UO_3289 (O_3289,N_46934,N_46182);
and UO_3290 (O_3290,N_43314,N_40691);
or UO_3291 (O_3291,N_44455,N_45283);
xor UO_3292 (O_3292,N_42449,N_43226);
xnor UO_3293 (O_3293,N_45731,N_49088);
or UO_3294 (O_3294,N_48651,N_47664);
nand UO_3295 (O_3295,N_48749,N_40404);
nand UO_3296 (O_3296,N_45930,N_43591);
xnor UO_3297 (O_3297,N_49828,N_40496);
nor UO_3298 (O_3298,N_41918,N_42392);
xnor UO_3299 (O_3299,N_45081,N_44540);
or UO_3300 (O_3300,N_41855,N_47644);
nor UO_3301 (O_3301,N_43663,N_41657);
and UO_3302 (O_3302,N_42752,N_48026);
xnor UO_3303 (O_3303,N_46841,N_43953);
xor UO_3304 (O_3304,N_49697,N_47094);
nor UO_3305 (O_3305,N_41042,N_45924);
nor UO_3306 (O_3306,N_48415,N_47140);
nand UO_3307 (O_3307,N_42860,N_49325);
nand UO_3308 (O_3308,N_49666,N_40307);
and UO_3309 (O_3309,N_44446,N_42191);
xor UO_3310 (O_3310,N_44465,N_40713);
and UO_3311 (O_3311,N_43270,N_44379);
nor UO_3312 (O_3312,N_42287,N_49160);
xor UO_3313 (O_3313,N_46937,N_45816);
nor UO_3314 (O_3314,N_46571,N_42180);
and UO_3315 (O_3315,N_44969,N_40990);
nand UO_3316 (O_3316,N_43880,N_48019);
nand UO_3317 (O_3317,N_47442,N_45497);
and UO_3318 (O_3318,N_41487,N_44924);
xor UO_3319 (O_3319,N_49411,N_42234);
nor UO_3320 (O_3320,N_47935,N_45154);
or UO_3321 (O_3321,N_46370,N_44979);
xnor UO_3322 (O_3322,N_40145,N_45243);
or UO_3323 (O_3323,N_42531,N_47583);
xnor UO_3324 (O_3324,N_46578,N_49143);
or UO_3325 (O_3325,N_40029,N_47668);
nor UO_3326 (O_3326,N_46615,N_45177);
or UO_3327 (O_3327,N_44618,N_49505);
and UO_3328 (O_3328,N_48682,N_43916);
xor UO_3329 (O_3329,N_43714,N_46847);
nor UO_3330 (O_3330,N_47074,N_44701);
and UO_3331 (O_3331,N_43404,N_49289);
nor UO_3332 (O_3332,N_42108,N_46138);
nand UO_3333 (O_3333,N_41751,N_47315);
and UO_3334 (O_3334,N_49194,N_48652);
and UO_3335 (O_3335,N_44499,N_45935);
or UO_3336 (O_3336,N_42943,N_47637);
xor UO_3337 (O_3337,N_44375,N_47038);
or UO_3338 (O_3338,N_45739,N_48064);
nand UO_3339 (O_3339,N_42316,N_42305);
xnor UO_3340 (O_3340,N_40817,N_47141);
xnor UO_3341 (O_3341,N_42730,N_43000);
and UO_3342 (O_3342,N_43668,N_42267);
nor UO_3343 (O_3343,N_47064,N_47444);
or UO_3344 (O_3344,N_45916,N_48896);
or UO_3345 (O_3345,N_45379,N_43876);
and UO_3346 (O_3346,N_40575,N_45079);
nor UO_3347 (O_3347,N_48938,N_46398);
xor UO_3348 (O_3348,N_41680,N_44438);
or UO_3349 (O_3349,N_42639,N_49647);
or UO_3350 (O_3350,N_48490,N_40024);
nor UO_3351 (O_3351,N_45412,N_48360);
or UO_3352 (O_3352,N_42906,N_44062);
or UO_3353 (O_3353,N_45305,N_43890);
xor UO_3354 (O_3354,N_43184,N_46941);
or UO_3355 (O_3355,N_47183,N_42718);
or UO_3356 (O_3356,N_49083,N_45409);
nor UO_3357 (O_3357,N_47443,N_45834);
nor UO_3358 (O_3358,N_48282,N_44752);
or UO_3359 (O_3359,N_48989,N_43524);
xor UO_3360 (O_3360,N_45478,N_41633);
and UO_3361 (O_3361,N_44301,N_48825);
xnor UO_3362 (O_3362,N_45025,N_45835);
nand UO_3363 (O_3363,N_46331,N_43613);
or UO_3364 (O_3364,N_49139,N_44734);
or UO_3365 (O_3365,N_42304,N_47976);
and UO_3366 (O_3366,N_45906,N_49997);
xor UO_3367 (O_3367,N_43584,N_48983);
nor UO_3368 (O_3368,N_42855,N_46045);
or UO_3369 (O_3369,N_46244,N_43920);
nor UO_3370 (O_3370,N_41188,N_43472);
and UO_3371 (O_3371,N_42792,N_47553);
and UO_3372 (O_3372,N_44631,N_40313);
or UO_3373 (O_3373,N_41414,N_46518);
xnor UO_3374 (O_3374,N_41619,N_47772);
nor UO_3375 (O_3375,N_44779,N_46141);
nor UO_3376 (O_3376,N_43144,N_40726);
nand UO_3377 (O_3377,N_42426,N_48653);
and UO_3378 (O_3378,N_43677,N_40823);
xor UO_3379 (O_3379,N_40542,N_40930);
xor UO_3380 (O_3380,N_40383,N_45912);
nand UO_3381 (O_3381,N_44235,N_42848);
and UO_3382 (O_3382,N_46196,N_44285);
xor UO_3383 (O_3383,N_42284,N_44218);
nor UO_3384 (O_3384,N_45972,N_48761);
xnor UO_3385 (O_3385,N_49497,N_48936);
nand UO_3386 (O_3386,N_40601,N_45311);
nand UO_3387 (O_3387,N_41363,N_40205);
and UO_3388 (O_3388,N_43710,N_44200);
nor UO_3389 (O_3389,N_46430,N_48050);
and UO_3390 (O_3390,N_46987,N_43733);
and UO_3391 (O_3391,N_40805,N_47694);
xnor UO_3392 (O_3392,N_48166,N_49121);
xnor UO_3393 (O_3393,N_46008,N_43960);
and UO_3394 (O_3394,N_45119,N_46775);
and UO_3395 (O_3395,N_43544,N_44482);
nand UO_3396 (O_3396,N_42504,N_44728);
nor UO_3397 (O_3397,N_47978,N_48138);
nand UO_3398 (O_3398,N_49296,N_43892);
and UO_3399 (O_3399,N_40375,N_42270);
nand UO_3400 (O_3400,N_43970,N_40186);
nand UO_3401 (O_3401,N_42170,N_45725);
xnor UO_3402 (O_3402,N_47781,N_40190);
or UO_3403 (O_3403,N_41678,N_47779);
xor UO_3404 (O_3404,N_49423,N_46428);
nor UO_3405 (O_3405,N_48163,N_49825);
nor UO_3406 (O_3406,N_44553,N_42370);
nor UO_3407 (O_3407,N_49010,N_40619);
and UO_3408 (O_3408,N_49871,N_43841);
or UO_3409 (O_3409,N_40492,N_41684);
or UO_3410 (O_3410,N_45948,N_40939);
xnor UO_3411 (O_3411,N_47745,N_44422);
and UO_3412 (O_3412,N_42642,N_48328);
nor UO_3413 (O_3413,N_46452,N_40483);
xor UO_3414 (O_3414,N_40825,N_44267);
nor UO_3415 (O_3415,N_41808,N_44384);
or UO_3416 (O_3416,N_43129,N_40960);
and UO_3417 (O_3417,N_45490,N_44616);
nor UO_3418 (O_3418,N_45399,N_43997);
nand UO_3419 (O_3419,N_45005,N_43842);
and UO_3420 (O_3420,N_45620,N_42386);
and UO_3421 (O_3421,N_44256,N_45833);
nor UO_3422 (O_3422,N_48405,N_41427);
xnor UO_3423 (O_3423,N_49218,N_44492);
nor UO_3424 (O_3424,N_47255,N_40648);
xor UO_3425 (O_3425,N_42744,N_48543);
nor UO_3426 (O_3426,N_40439,N_41513);
nand UO_3427 (O_3427,N_49940,N_42832);
or UO_3428 (O_3428,N_43570,N_42511);
nor UO_3429 (O_3429,N_41897,N_46532);
nand UO_3430 (O_3430,N_45993,N_42767);
nor UO_3431 (O_3431,N_45454,N_45092);
and UO_3432 (O_3432,N_42277,N_44390);
nor UO_3433 (O_3433,N_42551,N_44991);
nor UO_3434 (O_3434,N_40230,N_49346);
and UO_3435 (O_3435,N_44442,N_40942);
nor UO_3436 (O_3436,N_47955,N_40374);
and UO_3437 (O_3437,N_47435,N_43324);
and UO_3438 (O_3438,N_41903,N_44743);
xor UO_3439 (O_3439,N_48624,N_43988);
or UO_3440 (O_3440,N_42542,N_44849);
nand UO_3441 (O_3441,N_47119,N_48559);
and UO_3442 (O_3442,N_49785,N_42350);
or UO_3443 (O_3443,N_42788,N_46587);
xor UO_3444 (O_3444,N_49791,N_41901);
nor UO_3445 (O_3445,N_48079,N_45960);
or UO_3446 (O_3446,N_45442,N_48581);
xor UO_3447 (O_3447,N_46901,N_42717);
nand UO_3448 (O_3448,N_45678,N_48496);
and UO_3449 (O_3449,N_49511,N_45765);
nand UO_3450 (O_3450,N_43295,N_44780);
and UO_3451 (O_3451,N_48020,N_41453);
nor UO_3452 (O_3452,N_45193,N_46460);
and UO_3453 (O_3453,N_45744,N_49681);
nor UO_3454 (O_3454,N_41929,N_47520);
xnor UO_3455 (O_3455,N_49764,N_41536);
and UO_3456 (O_3456,N_46282,N_42940);
nor UO_3457 (O_3457,N_42374,N_41360);
nand UO_3458 (O_3458,N_45809,N_44022);
and UO_3459 (O_3459,N_41372,N_45427);
and UO_3460 (O_3460,N_46925,N_44645);
nand UO_3461 (O_3461,N_44096,N_43455);
and UO_3462 (O_3462,N_44898,N_43783);
nand UO_3463 (O_3463,N_44059,N_45940);
and UO_3464 (O_3464,N_44768,N_45361);
nor UO_3465 (O_3465,N_49582,N_49680);
xor UO_3466 (O_3466,N_46583,N_49981);
xnor UO_3467 (O_3467,N_47826,N_42112);
and UO_3468 (O_3468,N_47427,N_47933);
nand UO_3469 (O_3469,N_45545,N_41638);
nand UO_3470 (O_3470,N_44399,N_47092);
and UO_3471 (O_3471,N_48348,N_42963);
or UO_3472 (O_3472,N_49103,N_49476);
or UO_3473 (O_3473,N_40144,N_41704);
nor UO_3474 (O_3474,N_47759,N_45645);
and UO_3475 (O_3475,N_48545,N_45882);
xor UO_3476 (O_3476,N_42961,N_44500);
nor UO_3477 (O_3477,N_40168,N_48391);
nand UO_3478 (O_3478,N_47350,N_46341);
or UO_3479 (O_3479,N_44509,N_48390);
and UO_3480 (O_3480,N_46231,N_44165);
xnor UO_3481 (O_3481,N_46447,N_41252);
nand UO_3482 (O_3482,N_44770,N_44337);
and UO_3483 (O_3483,N_43847,N_48548);
xor UO_3484 (O_3484,N_40755,N_47341);
nor UO_3485 (O_3485,N_47614,N_45781);
and UO_3486 (O_3486,N_40032,N_45845);
and UO_3487 (O_3487,N_41576,N_40152);
or UO_3488 (O_3488,N_42687,N_41275);
nor UO_3489 (O_3489,N_49280,N_40038);
nor UO_3490 (O_3490,N_43047,N_42729);
or UO_3491 (O_3491,N_49459,N_47205);
and UO_3492 (O_3492,N_46202,N_49684);
or UO_3493 (O_3493,N_46489,N_42746);
or UO_3494 (O_3494,N_41464,N_49061);
nand UO_3495 (O_3495,N_49507,N_43458);
or UO_3496 (O_3496,N_45242,N_42338);
nor UO_3497 (O_3497,N_42618,N_43877);
xor UO_3498 (O_3498,N_43816,N_44491);
nand UO_3499 (O_3499,N_45495,N_47227);
and UO_3500 (O_3500,N_49806,N_42697);
xor UO_3501 (O_3501,N_40786,N_46723);
xnor UO_3502 (O_3502,N_41020,N_44587);
nor UO_3503 (O_3503,N_42144,N_41034);
or UO_3504 (O_3504,N_43859,N_49644);
or UO_3505 (O_3505,N_44575,N_47262);
nor UO_3506 (O_3506,N_49874,N_45089);
nor UO_3507 (O_3507,N_43193,N_43255);
nand UO_3508 (O_3508,N_47163,N_42790);
or UO_3509 (O_3509,N_48918,N_45841);
xnor UO_3510 (O_3510,N_42982,N_47045);
nor UO_3511 (O_3511,N_42950,N_40893);
and UO_3512 (O_3512,N_48547,N_43175);
nor UO_3513 (O_3513,N_47992,N_40039);
xnor UO_3514 (O_3514,N_41374,N_41258);
or UO_3515 (O_3515,N_48094,N_43725);
nand UO_3516 (O_3516,N_48431,N_44859);
and UO_3517 (O_3517,N_46950,N_40514);
and UO_3518 (O_3518,N_45245,N_44879);
and UO_3519 (O_3519,N_41497,N_41322);
xor UO_3520 (O_3520,N_43253,N_49227);
nand UO_3521 (O_3521,N_47687,N_41232);
nand UO_3522 (O_3522,N_46616,N_48948);
and UO_3523 (O_3523,N_48368,N_43338);
or UO_3524 (O_3524,N_45514,N_41871);
or UO_3525 (O_3525,N_48278,N_46811);
and UO_3526 (O_3526,N_42073,N_44801);
nor UO_3527 (O_3527,N_43183,N_45334);
or UO_3528 (O_3528,N_44073,N_48770);
nor UO_3529 (O_3529,N_44909,N_41348);
xnor UO_3530 (O_3530,N_44578,N_43172);
and UO_3531 (O_3531,N_46798,N_48521);
or UO_3532 (O_3532,N_48613,N_45051);
and UO_3533 (O_3533,N_49787,N_43125);
nor UO_3534 (O_3534,N_45551,N_46843);
or UO_3535 (O_3535,N_43681,N_49084);
and UO_3536 (O_3536,N_46158,N_44196);
xor UO_3537 (O_3537,N_48752,N_42145);
nand UO_3538 (O_3538,N_41605,N_46131);
nand UO_3539 (O_3539,N_40263,N_49353);
nor UO_3540 (O_3540,N_45142,N_48264);
xor UO_3541 (O_3541,N_42831,N_42308);
and UO_3542 (O_3542,N_42693,N_41493);
nand UO_3543 (O_3543,N_44796,N_49661);
and UO_3544 (O_3544,N_41449,N_47454);
nand UO_3545 (O_3545,N_41007,N_41418);
nor UO_3546 (O_3546,N_43804,N_46576);
xnor UO_3547 (O_3547,N_49482,N_44926);
nand UO_3548 (O_3548,N_41231,N_45526);
xnor UO_3549 (O_3549,N_46194,N_46610);
nor UO_3550 (O_3550,N_46422,N_48332);
and UO_3551 (O_3551,N_42352,N_48397);
xnor UO_3552 (O_3552,N_42072,N_47011);
and UO_3553 (O_3553,N_49770,N_45784);
xnor UO_3554 (O_3554,N_43893,N_44139);
nand UO_3555 (O_3555,N_42694,N_45471);
nor UO_3556 (O_3556,N_43414,N_42050);
nand UO_3557 (O_3557,N_48600,N_40052);
and UO_3558 (O_3558,N_47925,N_40324);
or UO_3559 (O_3559,N_45277,N_45260);
xor UO_3560 (O_3560,N_40594,N_42258);
or UO_3561 (O_3561,N_49012,N_47314);
and UO_3562 (O_3562,N_48307,N_46140);
or UO_3563 (O_3563,N_48792,N_40448);
xnor UO_3564 (O_3564,N_47991,N_47464);
nand UO_3565 (O_3565,N_42165,N_48513);
nand UO_3566 (O_3566,N_47145,N_49072);
or UO_3567 (O_3567,N_42800,N_41548);
and UO_3568 (O_3568,N_47727,N_46233);
and UO_3569 (O_3569,N_46060,N_47437);
xnor UO_3570 (O_3570,N_40912,N_47086);
or UO_3571 (O_3571,N_46374,N_49583);
nor UO_3572 (O_3572,N_44948,N_45295);
and UO_3573 (O_3573,N_44637,N_42178);
xnor UO_3574 (O_3574,N_46074,N_42420);
xor UO_3575 (O_3575,N_43951,N_48685);
nor UO_3576 (O_3576,N_44274,N_43447);
and UO_3577 (O_3577,N_47906,N_46599);
or UO_3578 (O_3578,N_42430,N_40264);
xnor UO_3579 (O_3579,N_46511,N_40970);
or UO_3580 (O_3580,N_40302,N_47200);
xor UO_3581 (O_3581,N_40415,N_42689);
and UO_3582 (O_3582,N_40036,N_47028);
nor UO_3583 (O_3583,N_49467,N_42833);
nor UO_3584 (O_3584,N_43553,N_41307);
or UO_3585 (O_3585,N_46459,N_45732);
xor UO_3586 (O_3586,N_44341,N_43093);
xor UO_3587 (O_3587,N_45991,N_42176);
or UO_3588 (O_3588,N_44042,N_41467);
or UO_3589 (O_3589,N_42993,N_41134);
and UO_3590 (O_3590,N_46279,N_46766);
or UO_3591 (O_3591,N_43086,N_41387);
nor UO_3592 (O_3592,N_40737,N_49419);
nand UO_3593 (O_3593,N_48274,N_44199);
nor UO_3594 (O_3594,N_44536,N_46521);
and UO_3595 (O_3595,N_42816,N_45267);
nor UO_3596 (O_3596,N_47936,N_45778);
nor UO_3597 (O_3597,N_43375,N_41655);
nand UO_3598 (O_3598,N_44978,N_44529);
or UO_3599 (O_3599,N_40265,N_49249);
nand UO_3600 (O_3600,N_43091,N_49294);
nor UO_3601 (O_3601,N_48969,N_44333);
nor UO_3602 (O_3602,N_47439,N_47252);
xnor UO_3603 (O_3603,N_44790,N_40756);
xnor UO_3604 (O_3604,N_47287,N_41159);
nor UO_3605 (O_3605,N_44029,N_47234);
and UO_3606 (O_3606,N_46119,N_44738);
xnor UO_3607 (O_3607,N_46256,N_43453);
nor UO_3608 (O_3608,N_41149,N_41103);
or UO_3609 (O_3609,N_44304,N_48224);
nor UO_3610 (O_3610,N_44935,N_41663);
or UO_3611 (O_3611,N_48446,N_46574);
and UO_3612 (O_3612,N_42574,N_45162);
or UO_3613 (O_3613,N_46090,N_47394);
nor UO_3614 (O_3614,N_43256,N_49676);
nor UO_3615 (O_3615,N_46413,N_44085);
or UO_3616 (O_3616,N_46557,N_48978);
and UO_3617 (O_3617,N_41393,N_43562);
nand UO_3618 (O_3618,N_49366,N_46872);
nor UO_3619 (O_3619,N_46710,N_41325);
and UO_3620 (O_3620,N_48161,N_43527);
nand UO_3621 (O_3621,N_48836,N_43311);
nand UO_3622 (O_3622,N_41505,N_49868);
nand UO_3623 (O_3623,N_43545,N_45256);
xnor UO_3624 (O_3624,N_43264,N_46475);
nor UO_3625 (O_3625,N_47137,N_46051);
xor UO_3626 (O_3626,N_40553,N_44134);
xnor UO_3627 (O_3627,N_47280,N_44183);
and UO_3628 (O_3628,N_44581,N_49003);
nand UO_3629 (O_3629,N_42528,N_44136);
nor UO_3630 (O_3630,N_44266,N_45808);
and UO_3631 (O_3631,N_45138,N_47026);
and UO_3632 (O_3632,N_47876,N_41632);
nor UO_3633 (O_3633,N_47703,N_40071);
xor UO_3634 (O_3634,N_45135,N_40583);
nand UO_3635 (O_3635,N_44383,N_48942);
and UO_3636 (O_3636,N_48200,N_45867);
nor UO_3637 (O_3637,N_44711,N_42715);
or UO_3638 (O_3638,N_41138,N_49041);
xor UO_3639 (O_3639,N_45464,N_47932);
and UO_3640 (O_3640,N_40703,N_47338);
and UO_3641 (O_3641,N_43477,N_40178);
nand UO_3642 (O_3642,N_43122,N_46099);
and UO_3643 (O_3643,N_49664,N_44506);
and UO_3644 (O_3644,N_44458,N_41522);
nor UO_3645 (O_3645,N_43933,N_46023);
xor UO_3646 (O_3646,N_46029,N_41170);
nand UO_3647 (O_3647,N_45319,N_47900);
nand UO_3648 (O_3648,N_43926,N_43166);
or UO_3649 (O_3649,N_44579,N_40000);
or UO_3650 (O_3650,N_47813,N_44841);
and UO_3651 (O_3651,N_48183,N_44857);
or UO_3652 (O_3652,N_42980,N_41783);
nand UO_3653 (O_3653,N_46346,N_42482);
xnor UO_3654 (O_3654,N_43647,N_48784);
nor UO_3655 (O_3655,N_49155,N_45705);
xor UO_3656 (O_3656,N_44245,N_49319);
nand UO_3657 (O_3657,N_45424,N_47807);
and UO_3658 (O_3658,N_49626,N_47023);
or UO_3659 (O_3659,N_44467,N_43040);
or UO_3660 (O_3660,N_46528,N_42057);
nand UO_3661 (O_3661,N_42310,N_41662);
xnor UO_3662 (O_3662,N_40096,N_44431);
nand UO_3663 (O_3663,N_43832,N_48826);
xor UO_3664 (O_3664,N_44568,N_48785);
or UO_3665 (O_3665,N_46047,N_45299);
nor UO_3666 (O_3666,N_46545,N_41519);
and UO_3667 (O_3667,N_41029,N_45448);
or UO_3668 (O_3668,N_44322,N_40192);
nand UO_3669 (O_3669,N_41864,N_45163);
and UO_3670 (O_3670,N_49952,N_42581);
or UO_3671 (O_3671,N_48802,N_45984);
nor UO_3672 (O_3672,N_41692,N_46118);
xnor UO_3673 (O_3673,N_46938,N_41179);
or UO_3674 (O_3674,N_48810,N_49159);
nand UO_3675 (O_3675,N_42192,N_42908);
and UO_3676 (O_3676,N_41326,N_47226);
xnor UO_3677 (O_3677,N_43856,N_44538);
nand UO_3678 (O_3678,N_40501,N_41390);
nand UO_3679 (O_3679,N_45724,N_40759);
and UO_3680 (O_3680,N_45408,N_42769);
xor UO_3681 (O_3681,N_40023,N_40938);
nor UO_3682 (O_3682,N_40993,N_48254);
xor UO_3683 (O_3683,N_43052,N_44312);
nor UO_3684 (O_3684,N_44374,N_40286);
nor UO_3685 (O_3685,N_49413,N_41588);
nor UO_3686 (O_3686,N_47977,N_46763);
nand UO_3687 (O_3687,N_48286,N_40582);
or UO_3688 (O_3688,N_46861,N_43727);
and UO_3689 (O_3689,N_48767,N_43987);
and UO_3690 (O_3690,N_44049,N_47070);
nand UO_3691 (O_3691,N_43021,N_49297);
xnor UO_3692 (O_3692,N_41891,N_45553);
nor UO_3693 (O_3693,N_45860,N_45297);
nand UO_3694 (O_3694,N_44002,N_44052);
nor UO_3695 (O_3695,N_48359,N_42622);
or UO_3696 (O_3696,N_43235,N_47107);
and UO_3697 (O_3697,N_41564,N_48162);
xor UO_3698 (O_3698,N_41853,N_47663);
xor UO_3699 (O_3699,N_44816,N_46467);
nand UO_3700 (O_3700,N_48788,N_42629);
nor UO_3701 (O_3701,N_45292,N_46940);
nand UO_3702 (O_3702,N_48146,N_44925);
xor UO_3703 (O_3703,N_47510,N_47692);
nor UO_3704 (O_3704,N_46087,N_49591);
and UO_3705 (O_3705,N_47940,N_48076);
nor UO_3706 (O_3706,N_49127,N_43786);
xnor UO_3707 (O_3707,N_41223,N_43837);
or UO_3708 (O_3708,N_47007,N_40668);
xor UO_3709 (O_3709,N_47217,N_46697);
nand UO_3710 (O_3710,N_42844,N_40170);
nor UO_3711 (O_3711,N_42233,N_45631);
nor UO_3712 (O_3712,N_41998,N_45595);
or UO_3713 (O_3713,N_40322,N_40395);
and UO_3714 (O_3714,N_47110,N_43278);
or UO_3715 (O_3715,N_47756,N_42481);
or UO_3716 (O_3716,N_47939,N_44094);
xor UO_3717 (O_3717,N_40357,N_48729);
and UO_3718 (O_3718,N_48720,N_44329);
or UO_3719 (O_3719,N_42005,N_49750);
nand UO_3720 (O_3720,N_44667,N_48851);
and UO_3721 (O_3721,N_48633,N_49492);
xor UO_3722 (O_3722,N_48127,N_42529);
or UO_3723 (O_3723,N_48060,N_43654);
and UO_3724 (O_3724,N_46596,N_45733);
and UO_3725 (O_3725,N_48047,N_47825);
xor UO_3726 (O_3726,N_47621,N_43168);
or UO_3727 (O_3727,N_49212,N_45918);
and UO_3728 (O_3728,N_48393,N_49120);
and UO_3729 (O_3729,N_44157,N_46516);
xor UO_3730 (O_3730,N_40126,N_48427);
and UO_3731 (O_3731,N_46286,N_46169);
xnor UO_3732 (O_3732,N_45265,N_49235);
xor UO_3733 (O_3733,N_49210,N_48656);
nor UO_3734 (O_3734,N_42959,N_48960);
nand UO_3735 (O_3735,N_42246,N_41118);
nand UO_3736 (O_3736,N_49430,N_49001);
or UO_3737 (O_3737,N_45286,N_45434);
nand UO_3738 (O_3738,N_47521,N_44563);
xor UO_3739 (O_3739,N_47412,N_41622);
xnor UO_3740 (O_3740,N_41613,N_49558);
nor UO_3741 (O_3741,N_46996,N_48433);
or UO_3742 (O_3742,N_42858,N_44754);
nand UO_3743 (O_3743,N_45694,N_44255);
nor UO_3744 (O_3744,N_42960,N_40524);
or UO_3745 (O_3745,N_42602,N_41828);
nand UO_3746 (O_3746,N_43887,N_49230);
and UO_3747 (O_3747,N_46291,N_40148);
and UO_3748 (O_3748,N_42589,N_47902);
nand UO_3749 (O_3749,N_40160,N_44433);
or UO_3750 (O_3750,N_46053,N_42263);
xnor UO_3751 (O_3751,N_41396,N_41925);
and UO_3752 (O_3752,N_49382,N_40320);
nor UO_3753 (O_3753,N_43445,N_49341);
and UO_3754 (O_3754,N_45115,N_43947);
or UO_3755 (O_3755,N_44041,N_47988);
and UO_3756 (O_3756,N_44149,N_47748);
nand UO_3757 (O_3757,N_40104,N_40556);
nor UO_3758 (O_3758,N_48186,N_40886);
or UO_3759 (O_3759,N_47344,N_44687);
and UO_3760 (O_3760,N_45354,N_42041);
xnor UO_3761 (O_3761,N_43973,N_49045);
and UO_3762 (O_3762,N_44122,N_47436);
and UO_3763 (O_3763,N_42827,N_42897);
nand UO_3764 (O_3764,N_48622,N_48561);
xor UO_3765 (O_3765,N_48456,N_44033);
and UO_3766 (O_3766,N_43867,N_44783);
or UO_3767 (O_3767,N_49288,N_45682);
xor UO_3768 (O_3768,N_44635,N_44530);
xor UO_3769 (O_3769,N_43711,N_44452);
and UO_3770 (O_3770,N_43576,N_42664);
or UO_3771 (O_3771,N_40915,N_45279);
xnor UO_3772 (O_3772,N_40088,N_47769);
nand UO_3773 (O_3773,N_40707,N_48229);
or UO_3774 (O_3774,N_43397,N_42741);
nor UO_3775 (O_3775,N_49519,N_47402);
nand UO_3776 (O_3776,N_41558,N_44437);
and UO_3777 (O_3777,N_47539,N_48974);
or UO_3778 (O_3778,N_49184,N_47475);
or UO_3779 (O_3779,N_45959,N_42312);
and UO_3780 (O_3780,N_41898,N_44717);
nand UO_3781 (O_3781,N_43327,N_49564);
xor UO_3782 (O_3782,N_44675,N_42466);
or UO_3783 (O_3783,N_46069,N_40789);
nor UO_3784 (O_3784,N_44168,N_43485);
and UO_3785 (O_3785,N_45687,N_49252);
nor UO_3786 (O_3786,N_40977,N_40478);
and UO_3787 (O_3787,N_49303,N_41642);
nor UO_3788 (O_3788,N_47202,N_47188);
and UO_3789 (O_3789,N_46828,N_48644);
and UO_3790 (O_3790,N_45157,N_47974);
xor UO_3791 (O_3791,N_40932,N_43934);
nand UO_3792 (O_3792,N_40012,N_44323);
nand UO_3793 (O_3793,N_44554,N_40765);
and UO_3794 (O_3794,N_45556,N_48700);
or UO_3795 (O_3795,N_40746,N_46626);
or UO_3796 (O_3796,N_46555,N_45662);
or UO_3797 (O_3797,N_48772,N_44496);
xor UO_3798 (O_3798,N_46958,N_42242);
nor UO_3799 (O_3799,N_48553,N_42182);
or UO_3800 (O_3800,N_40044,N_44417);
nand UO_3801 (O_3801,N_43990,N_45900);
or UO_3802 (O_3802,N_49035,N_41643);
or UO_3803 (O_3803,N_43044,N_45915);
nand UO_3804 (O_3804,N_44176,N_46560);
xnor UO_3805 (O_3805,N_45798,N_48343);
nor UO_3806 (O_3806,N_42559,N_49347);
nand UO_3807 (O_3807,N_42448,N_43318);
and UO_3808 (O_3808,N_47238,N_47957);
nor UO_3809 (O_3809,N_42171,N_43351);
nand UO_3810 (O_3810,N_43809,N_43238);
nor UO_3811 (O_3811,N_40468,N_41299);
nor UO_3812 (O_3812,N_42212,N_42365);
or UO_3813 (O_3813,N_40403,N_43650);
nor UO_3814 (O_3814,N_43633,N_40393);
xor UO_3815 (O_3815,N_48000,N_45074);
or UO_3816 (O_3816,N_44204,N_43975);
nor UO_3817 (O_3817,N_48225,N_46268);
and UO_3818 (O_3818,N_49506,N_43301);
nand UO_3819 (O_3819,N_49215,N_46968);
nor UO_3820 (O_3820,N_40944,N_47123);
xor UO_3821 (O_3821,N_44851,N_44408);
xnor UO_3822 (O_3822,N_48444,N_44832);
or UO_3823 (O_3823,N_44380,N_43686);
and UO_3824 (O_3824,N_44044,N_42393);
xnor UO_3825 (O_3825,N_47615,N_47993);
and UO_3826 (O_3826,N_49996,N_40653);
or UO_3827 (O_3827,N_47008,N_48494);
or UO_3828 (O_3828,N_40054,N_44532);
xnor UO_3829 (O_3829,N_47496,N_49030);
xor UO_3830 (O_3830,N_46065,N_47250);
or UO_3831 (O_3831,N_49941,N_45281);
nand UO_3832 (O_3832,N_45861,N_44003);
nand UO_3833 (O_3833,N_45000,N_46542);
nand UO_3834 (O_3834,N_45187,N_41446);
or UO_3835 (O_3835,N_42736,N_44708);
or UO_3836 (O_3836,N_45679,N_48745);
or UO_3837 (O_3837,N_42863,N_48217);
and UO_3838 (O_3838,N_41014,N_46210);
xnor UO_3839 (O_3839,N_43352,N_44992);
or UO_3840 (O_3840,N_49804,N_47055);
nand UO_3841 (O_3841,N_40515,N_43085);
or UO_3842 (O_3842,N_45995,N_41399);
xnor UO_3843 (O_3843,N_46944,N_41733);
and UO_3844 (O_3844,N_45017,N_45097);
nor UO_3845 (O_3845,N_48440,N_40630);
or UO_3846 (O_3846,N_42592,N_47578);
nand UO_3847 (O_3847,N_45742,N_41410);
nor UO_3848 (O_3848,N_45122,N_43817);
or UO_3849 (O_3849,N_47639,N_45703);
xnor UO_3850 (O_3850,N_46505,N_45322);
xnor UO_3851 (O_3851,N_47405,N_45977);
xnor UO_3852 (O_3852,N_40480,N_46192);
or UO_3853 (O_3853,N_47697,N_47641);
xor UO_3854 (O_3854,N_44813,N_40235);
nor UO_3855 (O_3855,N_41078,N_44672);
xnor UO_3856 (O_3856,N_42115,N_49466);
nor UO_3857 (O_3857,N_49739,N_46058);
or UO_3858 (O_3858,N_49138,N_44654);
or UO_3859 (O_3859,N_44930,N_40218);
or UO_3860 (O_3860,N_49905,N_40162);
nand UO_3861 (O_3861,N_45030,N_49461);
or UO_3862 (O_3862,N_47740,N_41292);
nand UO_3863 (O_3863,N_43755,N_48753);
nor UO_3864 (O_3864,N_43639,N_41053);
or UO_3865 (O_3865,N_43004,N_44657);
and UO_3866 (O_3866,N_45147,N_49822);
or UO_3867 (O_3867,N_44430,N_40020);
and UO_3868 (O_3868,N_45626,N_46972);
nand UO_3869 (O_3869,N_46073,N_44670);
and UO_3870 (O_3870,N_42238,N_46535);
nand UO_3871 (O_3871,N_46441,N_45753);
or UO_3872 (O_3872,N_41321,N_49282);
nand UO_3873 (O_3873,N_41753,N_42346);
nor UO_3874 (O_3874,N_48155,N_41361);
xnor UO_3875 (O_3875,N_43873,N_47269);
xnor UO_3876 (O_3876,N_48599,N_45604);
and UO_3877 (O_3877,N_43690,N_46358);
nor UO_3878 (O_3878,N_45211,N_42671);
nor UO_3879 (O_3879,N_43669,N_46067);
nand UO_3880 (O_3880,N_46267,N_40165);
and UO_3881 (O_3881,N_42972,N_42055);
or UO_3882 (O_3882,N_42032,N_40217);
and UO_3883 (O_3883,N_49361,N_48202);
xor UO_3884 (O_3884,N_48522,N_40987);
or UO_3885 (O_3885,N_42567,N_42010);
or UO_3886 (O_3886,N_47956,N_46501);
and UO_3887 (O_3887,N_43197,N_46410);
nand UO_3888 (O_3888,N_43280,N_47859);
xor UO_3889 (O_3889,N_47551,N_43595);
nand UO_3890 (O_3890,N_47638,N_41022);
and UO_3891 (O_3891,N_45127,N_40835);
or UO_3892 (O_3892,N_42117,N_43942);
or UO_3893 (O_3893,N_42302,N_42507);
and UO_3894 (O_3894,N_49147,N_41492);
nor UO_3895 (O_3895,N_46816,N_45352);
and UO_3896 (O_3896,N_49146,N_45248);
nor UO_3897 (O_3897,N_47885,N_45700);
or UO_3898 (O_3898,N_41173,N_46776);
xnor UO_3899 (O_3899,N_42530,N_43335);
and UO_3900 (O_3900,N_49795,N_41893);
and UO_3901 (O_3901,N_46645,N_43858);
xnor UO_3902 (O_3902,N_44292,N_40354);
and UO_3903 (O_3903,N_42978,N_43423);
and UO_3904 (O_3904,N_46597,N_48240);
xor UO_3905 (O_3905,N_42128,N_41221);
or UO_3906 (O_3906,N_49830,N_41623);
nand UO_3907 (O_3907,N_40810,N_42747);
nor UO_3908 (O_3908,N_47296,N_44932);
or UO_3909 (O_3909,N_49339,N_47677);
nor UO_3910 (O_3910,N_49310,N_42783);
nand UO_3911 (O_3911,N_44977,N_42856);
and UO_3912 (O_3912,N_40682,N_46624);
and UO_3913 (O_3913,N_45747,N_46646);
nor UO_3914 (O_3914,N_43361,N_41333);
xor UO_3915 (O_3915,N_40341,N_44010);
xor UO_3916 (O_3916,N_47861,N_49592);
and UO_3917 (O_3917,N_45346,N_47371);
nand UO_3918 (O_3918,N_40270,N_46976);
xor UO_3919 (O_3919,N_41431,N_40358);
xnor UO_3920 (O_3920,N_43019,N_46648);
and UO_3921 (O_3921,N_49898,N_40609);
nand UO_3922 (O_3922,N_46969,N_45827);
nor UO_3923 (O_3923,N_46882,N_41085);
nor UO_3924 (O_3924,N_40555,N_48419);
or UO_3925 (O_3925,N_47335,N_45870);
xor UO_3926 (O_3926,N_43580,N_45382);
or UO_3927 (O_3927,N_47778,N_42060);
nand UO_3928 (O_3928,N_43205,N_40280);
and UO_3929 (O_3929,N_40888,N_43006);
and UO_3930 (O_3930,N_48330,N_45776);
xnor UO_3931 (O_3931,N_42912,N_46878);
or UO_3932 (O_3932,N_41554,N_42535);
and UO_3933 (O_3933,N_46605,N_45837);
xor UO_3934 (O_3934,N_47414,N_40384);
xnor UO_3935 (O_3935,N_40865,N_43317);
nor UO_3936 (O_3936,N_47266,N_42739);
nand UO_3937 (O_3937,N_45792,N_44961);
nand UO_3938 (O_3938,N_48773,N_41141);
nor UO_3939 (O_3939,N_46593,N_44397);
nor UO_3940 (O_3940,N_43627,N_42677);
nand UO_3941 (O_3941,N_45874,N_48208);
xnor UO_3942 (O_3942,N_45605,N_49163);
or UO_3943 (O_3943,N_40696,N_41302);
nor UO_3944 (O_3944,N_49870,N_41982);
and UO_3945 (O_3945,N_43362,N_46849);
nand UO_3946 (O_3946,N_44244,N_44868);
or UO_3947 (O_3947,N_41761,N_42134);
xor UO_3948 (O_3948,N_42464,N_47690);
xor UO_3949 (O_3949,N_41961,N_49882);
xnor UO_3950 (O_3950,N_43425,N_49796);
and UO_3951 (O_3951,N_45287,N_45942);
xnor UO_3952 (O_3952,N_40111,N_42948);
or UO_3953 (O_3953,N_48732,N_45113);
nor UO_3954 (O_3954,N_41634,N_48886);
xor UO_3955 (O_3955,N_42927,N_49994);
nor UO_3956 (O_3956,N_44820,N_46062);
or UO_3957 (O_3957,N_45975,N_47481);
and UO_3958 (O_3958,N_43039,N_47709);
nand UO_3959 (O_3959,N_40094,N_45515);
nand UO_3960 (O_3960,N_41627,N_48012);
nor UO_3961 (O_3961,N_48122,N_47323);
and UO_3962 (O_3962,N_48314,N_44919);
and UO_3963 (O_3963,N_42949,N_48366);
or UO_3964 (O_3964,N_40121,N_48301);
and UO_3965 (O_3965,N_43049,N_47159);
nand UO_3966 (O_3966,N_47722,N_42824);
nand UO_3967 (O_3967,N_41631,N_44424);
nor UO_3968 (O_3968,N_46419,N_47099);
or UO_3969 (O_3969,N_40614,N_49053);
and UO_3970 (O_3970,N_41728,N_43011);
xor UO_3971 (O_3971,N_46100,N_45560);
or UO_3972 (O_3972,N_49763,N_44545);
nor UO_3973 (O_3973,N_40229,N_48420);
xnor UO_3974 (O_3974,N_40745,N_42696);
nand UO_3975 (O_3975,N_47809,N_41884);
or UO_3976 (O_3976,N_46512,N_46136);
nand UO_3977 (O_3977,N_46311,N_45301);
nor UO_3978 (O_3978,N_42222,N_49248);
nor UO_3979 (O_3979,N_47194,N_44590);
or UO_3980 (O_3980,N_41601,N_46168);
nand UO_3981 (O_3981,N_44943,N_41878);
and UO_3982 (O_3982,N_48123,N_42462);
xnor UO_3983 (O_3983,N_49983,N_48925);
nor UO_3984 (O_3984,N_43604,N_44981);
and UO_3985 (O_3985,N_49960,N_47281);
nor UO_3986 (O_3986,N_48849,N_49642);
and UO_3987 (O_3987,N_47533,N_46020);
or UO_3988 (O_3988,N_40920,N_48388);
nand UO_3989 (O_3989,N_48567,N_43879);
xor UO_3990 (O_3990,N_46461,N_45355);
or UO_3991 (O_3991,N_40476,N_40293);
nor UO_3992 (O_3992,N_49047,N_45598);
and UO_3993 (O_3993,N_41615,N_45086);
or UO_3994 (O_3994,N_45338,N_44975);
and UO_3995 (O_3995,N_47944,N_42146);
or UO_3996 (O_3996,N_43444,N_49972);
xor UO_3997 (O_3997,N_47582,N_40577);
and UO_3998 (O_3998,N_49553,N_47595);
nor UO_3999 (O_3999,N_42917,N_45288);
and UO_4000 (O_4000,N_48937,N_40095);
nand UO_4001 (O_4001,N_47719,N_43499);
xor UO_4002 (O_4002,N_44345,N_41246);
or UO_4003 (O_4003,N_48789,N_49385);
nor UO_4004 (O_4004,N_42499,N_44469);
nor UO_4005 (O_4005,N_43930,N_49008);
or UO_4006 (O_4006,N_47705,N_43421);
xor UO_4007 (O_4007,N_46092,N_47278);
nor UO_4008 (O_4008,N_44043,N_44463);
nand UO_4009 (O_4009,N_44387,N_48718);
nand UO_4010 (O_4010,N_48044,N_47305);
nand UO_4011 (O_4011,N_47725,N_45380);
and UO_4012 (O_4012,N_48475,N_40868);
or UO_4013 (O_4013,N_43728,N_42143);
xor UO_4014 (O_4014,N_46529,N_43862);
nor UO_4015 (O_4015,N_44185,N_47272);
nand UO_4016 (O_4016,N_48819,N_40654);
or UO_4017 (O_4017,N_49259,N_48344);
and UO_4018 (O_4018,N_48479,N_41331);
nor UO_4019 (O_4019,N_49704,N_47652);
and UO_4020 (O_4020,N_48149,N_47425);
nor UO_4021 (O_4021,N_44321,N_41241);
xor UO_4022 (O_4022,N_46818,N_48941);
or UO_4023 (O_4023,N_44658,N_47134);
nand UO_4024 (O_4024,N_41683,N_42568);
xnor UO_4025 (O_4025,N_44360,N_46990);
and UO_4026 (O_4026,N_41701,N_44175);
or UO_4027 (O_4027,N_49615,N_45643);
nor UO_4028 (O_4028,N_43635,N_44147);
and UO_4029 (O_4029,N_44427,N_42740);
or UO_4030 (O_4030,N_42550,N_45639);
xnor UO_4031 (O_4031,N_46221,N_40518);
nand UO_4032 (O_4032,N_48302,N_49065);
nand UO_4033 (O_4033,N_43037,N_42331);
xor UO_4034 (O_4034,N_49273,N_47701);
nand UO_4035 (O_4035,N_48136,N_40909);
nor UO_4036 (O_4036,N_45259,N_42806);
nand UO_4037 (O_4037,N_45418,N_43373);
xnor UO_4038 (O_4038,N_43631,N_47177);
or UO_4039 (O_4039,N_45280,N_47365);
nand UO_4040 (O_4040,N_46884,N_46367);
and UO_4041 (O_4041,N_48866,N_42538);
nand UO_4042 (O_4042,N_49906,N_40636);
and UO_4043 (O_4043,N_49820,N_44644);
or UO_4044 (O_4044,N_42690,N_48478);
and UO_4045 (O_4045,N_44173,N_47047);
or UO_4046 (O_4046,N_42682,N_43332);
or UO_4047 (O_4047,N_49453,N_44356);
or UO_4048 (O_4048,N_42981,N_47973);
nand UO_4049 (O_4049,N_49488,N_49276);
or UO_4050 (O_4050,N_42616,N_48852);
nand UO_4051 (O_4051,N_43802,N_41177);
and UO_4052 (O_4052,N_49034,N_49225);
and UO_4053 (O_4053,N_47867,N_40808);
xnor UO_4054 (O_4054,N_49546,N_47063);
or UO_4055 (O_4055,N_44720,N_41767);
xor UO_4056 (O_4056,N_43322,N_49593);
xnor UO_4057 (O_4057,N_40898,N_47717);
and UO_4058 (O_4058,N_44662,N_41816);
or UO_4059 (O_4059,N_48970,N_44060);
nor UO_4060 (O_4060,N_40958,N_40142);
and UO_4061 (O_4061,N_41702,N_40757);
nand UO_4062 (O_4062,N_40878,N_46834);
nor UO_4063 (O_4063,N_47039,N_49236);
nor UO_4064 (O_4064,N_45218,N_40728);
xnor UO_4065 (O_4065,N_40037,N_49568);
or UO_4066 (O_4066,N_40033,N_40743);
nor UO_4067 (O_4067,N_43582,N_46133);
or UO_4068 (O_4068,N_47343,N_41290);
nor UO_4069 (O_4069,N_43289,N_42131);
nor UO_4070 (O_4070,N_40572,N_41469);
nor UO_4071 (O_4071,N_48654,N_42439);
xor UO_4072 (O_4072,N_45179,N_46160);
xnor UO_4073 (O_4073,N_49690,N_41557);
or UO_4074 (O_4074,N_42082,N_48683);
nor UO_4075 (O_4075,N_46255,N_41124);
nor UO_4076 (O_4076,N_44781,N_47385);
nor UO_4077 (O_4077,N_41570,N_47755);
or UO_4078 (O_4078,N_43419,N_40430);
nor UO_4079 (O_4079,N_42168,N_47642);
and UO_4080 (O_4080,N_43778,N_46307);
nand UO_4081 (O_4081,N_43619,N_48341);
or UO_4082 (O_4082,N_49944,N_45955);
and UO_4083 (O_4083,N_44908,N_40271);
xnor UO_4084 (O_4084,N_41426,N_41092);
nor UO_4085 (O_4085,N_48432,N_49605);
nor UO_4086 (O_4086,N_42106,N_40489);
or UO_4087 (O_4087,N_47077,N_46070);
xor UO_4088 (O_4088,N_49927,N_48326);
and UO_4089 (O_4089,N_41575,N_47594);
nand UO_4090 (O_4090,N_44746,N_48834);
nand UO_4091 (O_4091,N_45268,N_47802);
nand UO_4092 (O_4092,N_47724,N_46288);
and UO_4093 (O_4093,N_48731,N_45688);
and UO_4094 (O_4094,N_47731,N_41199);
xnor UO_4095 (O_4095,N_44518,N_42678);
nand UO_4096 (O_4096,N_43752,N_45291);
nand UO_4097 (O_4097,N_41280,N_47057);
xnor UO_4098 (O_4098,N_48759,N_43171);
nor UO_4099 (O_4099,N_43392,N_40011);
nor UO_4100 (O_4100,N_40581,N_44205);
or UO_4101 (O_4101,N_45021,N_44249);
and UO_4102 (O_4102,N_40461,N_44106);
nor UO_4103 (O_4103,N_49077,N_49358);
or UO_4104 (O_4104,N_48218,N_48867);
nand UO_4105 (O_4105,N_45863,N_41962);
nor UO_4106 (O_4106,N_45509,N_45511);
and UO_4107 (O_4107,N_40672,N_43875);
xor UO_4108 (O_4108,N_41671,N_40688);
nor UO_4109 (O_4109,N_41806,N_45843);
and UO_4110 (O_4110,N_41354,N_45825);
nand UO_4111 (O_4111,N_43516,N_46235);
xor UO_4112 (O_4112,N_46713,N_41273);
and UO_4113 (O_4113,N_45250,N_48997);
or UO_4114 (O_4114,N_48809,N_42417);
and UO_4115 (O_4115,N_43230,N_48829);
nand UO_4116 (O_4116,N_46391,N_43848);
xnor UO_4117 (O_4117,N_41496,N_42838);
and UO_4118 (O_4118,N_41405,N_43567);
and UO_4119 (O_4119,N_42273,N_40135);
nor UO_4120 (O_4120,N_45806,N_42295);
or UO_4121 (O_4121,N_46919,N_41965);
or UO_4122 (O_4122,N_48520,N_49398);
nand UO_4123 (O_4123,N_40928,N_41890);
or UO_4124 (O_4124,N_44605,N_49190);
xor UO_4125 (O_4125,N_41698,N_45819);
nor UO_4126 (O_4126,N_40046,N_47699);
xor UO_4127 (O_4127,N_46213,N_40876);
and UO_4128 (O_4128,N_44061,N_43735);
and UO_4129 (O_4129,N_43914,N_48658);
and UO_4130 (O_4130,N_41009,N_40749);
xnor UO_4131 (O_4131,N_44679,N_44254);
or UO_4132 (O_4132,N_49682,N_45952);
nand UO_4133 (O_4133,N_40770,N_41286);
or UO_4134 (O_4134,N_46176,N_41419);
nor UO_4135 (O_4135,N_45343,N_47914);
nor UO_4136 (O_4136,N_41211,N_47556);
nor UO_4137 (O_4137,N_43396,N_41433);
nor UO_4138 (O_4138,N_43105,N_40816);
and UO_4139 (O_4139,N_44282,N_49468);
nor UO_4140 (O_4140,N_46917,N_43511);
and UO_4141 (O_4141,N_49515,N_44092);
nand UO_4142 (O_4142,N_45537,N_46033);
or UO_4143 (O_4143,N_43154,N_47292);
or UO_4144 (O_4144,N_48820,N_47299);
nand UO_4145 (O_4145,N_48443,N_49725);
xor UO_4146 (O_4146,N_47282,N_41448);
nor UO_4147 (O_4147,N_42363,N_48719);
and UO_4148 (O_4148,N_48411,N_42644);
nor UO_4149 (O_4149,N_47089,N_43434);
or UO_4150 (O_4150,N_40290,N_46974);
xnor UO_4151 (O_4151,N_43911,N_43119);
nor UO_4152 (O_4152,N_41269,N_43653);
and UO_4153 (O_4153,N_42132,N_40371);
nand UO_4154 (O_4154,N_49202,N_47985);
or UO_4155 (O_4155,N_40463,N_47181);
nand UO_4156 (O_4156,N_47330,N_41010);
nand UO_4157 (O_4157,N_44287,N_42030);
nor UO_4158 (O_4158,N_40729,N_49569);
xnor UO_4159 (O_4159,N_46838,N_44250);
xnor UO_4160 (O_4160,N_49517,N_43228);
and UO_4161 (O_4161,N_45492,N_44289);
nand UO_4162 (O_4162,N_42035,N_42429);
nand UO_4163 (O_4163,N_42371,N_45275);
or UO_4164 (O_4164,N_40892,N_48618);
nor UO_4165 (O_4165,N_42098,N_48375);
nand UO_4166 (O_4166,N_43416,N_41386);
nor UO_4167 (O_4167,N_46725,N_44799);
or UO_4168 (O_4168,N_45100,N_48387);
nor UO_4169 (O_4169,N_47768,N_46791);
nand UO_4170 (O_4170,N_44582,N_48057);
nand UO_4171 (O_4171,N_41625,N_48072);
or UO_4172 (O_4172,N_49865,N_43025);
and UO_4173 (O_4173,N_46266,N_47105);
nor UO_4174 (O_4174,N_46211,N_40106);
and UO_4175 (O_4175,N_44762,N_43835);
xnor UO_4176 (O_4176,N_42061,N_46025);
nand UO_4177 (O_4177,N_40214,N_46048);
xnor UO_4178 (O_4178,N_47622,N_43411);
and UO_4179 (O_4179,N_47507,N_48184);
nand UO_4180 (O_4180,N_46094,N_42786);
nand UO_4181 (O_4181,N_48144,N_43897);
nor UO_4182 (O_4182,N_47770,N_41059);
nand UO_4183 (O_4183,N_40568,N_42931);
or UO_4184 (O_4184,N_40034,N_40429);
nor UO_4185 (O_4185,N_43257,N_45842);
nor UO_4186 (O_4186,N_49063,N_44609);
nor UO_4187 (O_4187,N_49412,N_48510);
or UO_4188 (O_4188,N_40334,N_45902);
nor UO_4189 (O_4189,N_40329,N_46623);
nor UO_4190 (O_4190,N_49318,N_42865);
xor UO_4191 (O_4191,N_41951,N_47245);
xnor UO_4192 (O_4192,N_49761,N_43517);
or UO_4193 (O_4193,N_42795,N_42051);
and UO_4194 (O_4194,N_43687,N_46157);
or UO_4195 (O_4195,N_40824,N_47706);
nor UO_4196 (O_4196,N_41438,N_49020);
xnor UO_4197 (O_4197,N_42460,N_40353);
nand UO_4198 (O_4198,N_40787,N_42652);
and UO_4199 (O_4199,N_49452,N_40376);
and UO_4200 (O_4200,N_48902,N_44346);
nor UO_4201 (O_4201,N_49819,N_40721);
xnor UO_4202 (O_4202,N_48845,N_44693);
xnor UO_4203 (O_4203,N_47567,N_43084);
and UO_4204 (O_4204,N_47696,N_48499);
and UO_4205 (O_4205,N_48514,N_49115);
nor UO_4206 (O_4206,N_47428,N_47782);
xnor UO_4207 (O_4207,N_45498,N_44551);
nand UO_4208 (O_4208,N_42712,N_46253);
xor UO_4209 (O_4209,N_43276,N_41773);
nor UO_4210 (O_4210,N_49380,N_43552);
and UO_4211 (O_4211,N_41082,N_48458);
nor UO_4212 (O_4212,N_47640,N_46966);
nand UO_4213 (O_4213,N_49192,N_41060);
or UO_4214 (O_4214,N_49374,N_40536);
or UO_4215 (O_4215,N_42452,N_47573);
and UO_4216 (O_4216,N_43177,N_48096);
and UO_4217 (O_4217,N_41919,N_45065);
or UO_4218 (O_4218,N_40164,N_47860);
and UO_4219 (O_4219,N_44611,N_43541);
nor UO_4220 (O_4220,N_47729,N_40840);
and UO_4221 (O_4221,N_43306,N_42920);
and UO_4222 (O_4222,N_42015,N_47348);
or UO_4223 (O_4223,N_40098,N_43260);
nor UO_4224 (O_4224,N_46640,N_40361);
or UO_4225 (O_4225,N_49974,N_42450);
xor UO_4226 (O_4226,N_46220,N_41553);
xor UO_4227 (O_4227,N_49432,N_41602);
nor UO_4228 (O_4228,N_41310,N_40530);
and UO_4229 (O_4229,N_46980,N_44019);
xnor UO_4230 (O_4230,N_49277,N_49653);
nor UO_4231 (O_4231,N_49096,N_45053);
nor UO_4232 (O_4232,N_42969,N_45704);
and UO_4233 (O_4233,N_42756,N_45996);
nand UO_4234 (O_4234,N_43977,N_45658);
nand UO_4235 (O_4235,N_49087,N_42086);
and UO_4236 (O_4236,N_48988,N_45313);
nand UO_4237 (O_4237,N_44775,N_40879);
and UO_4238 (O_4238,N_49834,N_41130);
xnor UO_4239 (O_4239,N_42456,N_45143);
nor UO_4240 (O_4240,N_41937,N_40558);
and UO_4241 (O_4241,N_48247,N_45337);
xnor UO_4242 (O_4242,N_40276,N_48182);
or UO_4243 (O_4243,N_42620,N_46922);
or UO_4244 (O_4244,N_42029,N_40869);
or UO_4245 (O_4245,N_47994,N_41481);
xnor UO_4246 (O_4246,N_47571,N_40736);
xnor UO_4247 (O_4247,N_42918,N_42975);
or UO_4248 (O_4248,N_40432,N_44334);
nand UO_4249 (O_4249,N_40189,N_47577);
xor UO_4250 (O_4250,N_42612,N_49464);
xor UO_4251 (O_4251,N_41997,N_41574);
and UO_4252 (O_4252,N_41836,N_40202);
nand UO_4253 (O_4253,N_41285,N_47949);
xor UO_4254 (O_4254,N_40785,N_47832);
and UO_4255 (O_4255,N_46298,N_46050);
or UO_4256 (O_4256,N_48180,N_40120);
and UO_4257 (O_4257,N_45290,N_40130);
nor UO_4258 (O_4258,N_42444,N_42649);
xor UO_4259 (O_4259,N_40179,N_44230);
xor UO_4260 (O_4260,N_44829,N_44959);
nor UO_4261 (O_4261,N_46232,N_48194);
nand UO_4262 (O_4262,N_49241,N_41689);
nor UO_4263 (O_4263,N_48287,N_47959);
and UO_4264 (O_4264,N_45770,N_45929);
nand UO_4265 (O_4265,N_45866,N_45033);
nor UO_4266 (O_4266,N_40003,N_41388);
or UO_4267 (O_4267,N_48842,N_44454);
nor UO_4268 (O_4268,N_40616,N_49300);
nand UO_4269 (O_4269,N_41030,N_49333);
xnor UO_4270 (O_4270,N_46703,N_43767);
nor UO_4271 (O_4271,N_45123,N_44649);
nand UO_4272 (O_4272,N_44852,N_49473);
and UO_4273 (O_4273,N_40351,N_40363);
nor UO_4274 (O_4274,N_48934,N_43371);
or UO_4275 (O_4275,N_44604,N_45936);
or UO_4276 (O_4276,N_49888,N_48591);
or UO_4277 (O_4277,N_45986,N_48502);
nand UO_4278 (O_4278,N_49313,N_45789);
xor UO_4279 (O_4279,N_44528,N_41677);
nor UO_4280 (O_4280,N_46262,N_48791);
and UO_4281 (O_4281,N_42742,N_43609);
or UO_4282 (O_4282,N_41174,N_44114);
and UO_4283 (O_4283,N_46369,N_43944);
xor UO_4284 (O_4284,N_40294,N_41599);
and UO_4285 (O_4285,N_46784,N_41123);
xnor UO_4286 (O_4286,N_46948,N_41382);
xnor UO_4287 (O_4287,N_41984,N_48551);
and UO_4288 (O_4288,N_48693,N_44121);
or UO_4289 (O_4289,N_43163,N_43774);
and UO_4290 (O_4290,N_43053,N_48279);
or UO_4291 (O_4291,N_47795,N_47135);
and UO_4292 (O_4292,N_48093,N_43236);
and UO_4293 (O_4293,N_40224,N_49090);
nand UO_4294 (O_4294,N_49377,N_44823);
or UO_4295 (O_4295,N_45814,N_44896);
or UO_4296 (O_4296,N_45954,N_40254);
xnor UO_4297 (O_4297,N_42632,N_40438);
and UO_4298 (O_4298,N_49089,N_47597);
xnor UO_4299 (O_4299,N_43509,N_46411);
and UO_4300 (O_4300,N_47685,N_44993);
or UO_4301 (O_4301,N_41239,N_48587);
xor UO_4302 (O_4302,N_45184,N_43846);
xnor UO_4303 (O_4303,N_44845,N_42463);
nor UO_4304 (O_4304,N_49589,N_42383);
nor UO_4305 (O_4305,N_42268,N_43995);
nor UO_4306 (O_4306,N_42952,N_43002);
or UO_4307 (O_4307,N_49400,N_43209);
or UO_4308 (O_4308,N_45335,N_44261);
nor UO_4309 (O_4309,N_41389,N_43033);
xnor UO_4310 (O_4310,N_45461,N_45426);
or UO_4311 (O_4311,N_45681,N_48015);
nand UO_4312 (O_4312,N_47666,N_47458);
and UO_4313 (O_4313,N_44523,N_40626);
nor UO_4314 (O_4314,N_40724,N_44838);
or UO_4315 (O_4315,N_43399,N_43632);
xnor UO_4316 (O_4316,N_45563,N_42525);
nor UO_4317 (O_4317,N_45249,N_43266);
or UO_4318 (O_4318,N_44090,N_46595);
nor UO_4319 (O_4319,N_40158,N_41008);
xor UO_4320 (O_4320,N_44927,N_43440);
nor UO_4321 (O_4321,N_43683,N_45899);
or UO_4322 (O_4322,N_46107,N_41089);
xnor UO_4323 (O_4323,N_43222,N_45876);
nor UO_4324 (O_4324,N_41764,N_44546);
and UO_4325 (O_4325,N_49457,N_44494);
and UO_4326 (O_4326,N_40385,N_45362);
nor UO_4327 (O_4327,N_47864,N_45980);
xor UO_4328 (O_4328,N_42745,N_45332);
nand UO_4329 (O_4329,N_44115,N_44178);
nor UO_4330 (O_4330,N_47192,N_48519);
nor UO_4331 (O_4331,N_47329,N_42988);
and UO_4332 (O_4332,N_47889,N_41294);
xnor UO_4333 (O_4333,N_47516,N_44068);
and UO_4334 (O_4334,N_41732,N_42885);
or UO_4335 (O_4335,N_47896,N_40450);
nor UO_4336 (O_4336,N_43418,N_44216);
nor UO_4337 (O_4337,N_45251,N_41829);
and UO_4338 (O_4338,N_40049,N_41458);
nor UO_4339 (O_4339,N_46421,N_41859);
or UO_4340 (O_4340,N_47473,N_46767);
nand UO_4341 (O_4341,N_49778,N_42500);
xor UO_4342 (O_4342,N_40295,N_41186);
nand UO_4343 (O_4343,N_40740,N_42591);
or UO_4344 (O_4344,N_46218,N_46438);
nor UO_4345 (O_4345,N_48634,N_49028);
xor UO_4346 (O_4346,N_48667,N_46637);
nand UO_4347 (O_4347,N_42819,N_47128);
and UO_4348 (O_4348,N_48068,N_42492);
or UO_4349 (O_4349,N_41265,N_45111);
nor UO_4350 (O_4350,N_48575,N_41488);
and UO_4351 (O_4351,N_48998,N_42353);
nand UO_4352 (O_4352,N_42513,N_43464);
nor UO_4353 (O_4353,N_43685,N_47421);
nand UO_4354 (O_4354,N_42973,N_47112);
or UO_4355 (O_4355,N_47386,N_45166);
and UO_4356 (O_4356,N_45197,N_46466);
xnor UO_4357 (O_4357,N_40947,N_49102);
nand UO_4358 (O_4358,N_41365,N_40699);
and UO_4359 (O_4359,N_45389,N_41790);
or UO_4360 (O_4360,N_48320,N_44945);
nor UO_4361 (O_4361,N_44308,N_43764);
xnor UO_4362 (O_4362,N_44844,N_46081);
or UO_4363 (O_4363,N_42764,N_49651);
or UO_4364 (O_4364,N_44381,N_43294);
nand UO_4365 (O_4365,N_47498,N_43219);
xor UO_4366 (O_4366,N_48085,N_47236);
xnor UO_4367 (O_4367,N_45534,N_48831);
xnor UO_4368 (O_4368,N_40498,N_40279);
nor UO_4369 (O_4369,N_41567,N_46105);
xnor UO_4370 (O_4370,N_40346,N_46899);
nor UO_4371 (O_4371,N_40693,N_45148);
and UO_4372 (O_4372,N_42909,N_41063);
nand UO_4373 (O_4373,N_42483,N_49173);
nand UO_4374 (O_4374,N_48620,N_46336);
and UO_4375 (O_4375,N_44082,N_40382);
and UO_4376 (O_4376,N_49224,N_47989);
xor UO_4377 (O_4377,N_43141,N_46431);
and UO_4378 (O_4378,N_41518,N_49111);
and UO_4379 (O_4379,N_44550,N_48550);
xor UO_4380 (O_4380,N_47730,N_46252);
nand UO_4381 (O_4381,N_41668,N_43395);
and UO_4382 (O_4382,N_40867,N_48777);
nor UO_4383 (O_4383,N_49850,N_46191);
nand UO_4384 (O_4384,N_40797,N_41421);
nor UO_4385 (O_4385,N_45623,N_44124);
nand UO_4386 (O_4386,N_42428,N_43365);
or UO_4387 (O_4387,N_48944,N_43089);
xnor UO_4388 (O_4388,N_44732,N_42358);
or UO_4389 (O_4389,N_41178,N_44606);
nand UO_4390 (O_4390,N_40097,N_42990);
nand UO_4391 (O_4391,N_43623,N_49094);
or UO_4392 (O_4392,N_45880,N_48953);
and UO_4393 (O_4393,N_45255,N_45333);
xnor UO_4394 (O_4394,N_42757,N_43523);
xnor UO_4395 (O_4395,N_46683,N_41953);
or UO_4396 (O_4396,N_41335,N_41116);
and UO_4397 (O_4397,N_47187,N_40424);
xor UO_4398 (O_4398,N_40951,N_43991);
nor UO_4399 (O_4399,N_44448,N_41436);
or UO_4400 (O_4400,N_49293,N_42701);
and UO_4401 (O_4401,N_41271,N_45314);
and UO_4402 (O_4402,N_46342,N_47052);
nor UO_4403 (O_4403,N_43088,N_43982);
or UO_4404 (O_4404,N_48853,N_41018);
or UO_4405 (O_4405,N_44184,N_41818);
and UO_4406 (O_4406,N_44045,N_49458);
nor UO_4407 (O_4407,N_41240,N_45198);
or UO_4408 (O_4408,N_49343,N_43955);
and UO_4409 (O_4409,N_45990,N_46694);
and UO_4410 (O_4410,N_48892,N_41600);
xor UO_4411 (O_4411,N_42040,N_44682);
and UO_4412 (O_4412,N_42179,N_49857);
nor UO_4413 (O_4413,N_42445,N_49389);
or UO_4414 (O_4414,N_46497,N_44650);
or UO_4415 (O_4415,N_46895,N_41747);
and UO_4416 (O_4416,N_44007,N_42519);
and UO_4417 (O_4417,N_42487,N_45779);
xnor UO_4418 (O_4418,N_41484,N_49545);
or UO_4419 (O_4419,N_44769,N_47267);
nand UO_4420 (O_4420,N_43526,N_47862);
xnor UO_4421 (O_4421,N_48894,N_49675);
nor UO_4422 (O_4422,N_45433,N_49520);
xor UO_4423 (O_4423,N_48069,N_48361);
xnor UO_4424 (O_4424,N_45315,N_40752);
nand UO_4425 (O_4425,N_49840,N_49754);
xor UO_4426 (O_4426,N_45042,N_47489);
xor UO_4427 (O_4427,N_46203,N_45877);
nand UO_4428 (O_4428,N_46139,N_49713);
nand UO_4429 (O_4429,N_45883,N_40277);
and UO_4430 (O_4430,N_46741,N_47129);
nand UO_4431 (O_4431,N_46924,N_43566);
xor UO_4432 (O_4432,N_44692,N_43560);
xor UO_4433 (O_4433,N_42303,N_44974);
nor UO_4434 (O_4434,N_45622,N_49720);
xor UO_4435 (O_4435,N_43420,N_48018);
nor UO_4436 (O_4436,N_47817,N_44760);
nor UO_4437 (O_4437,N_42802,N_42768);
or UO_4438 (O_4438,N_47536,N_44392);
nand UO_4439 (O_4439,N_40784,N_49616);
or UO_4440 (O_4440,N_48315,N_44293);
nand UO_4441 (O_4441,N_48345,N_41278);
nand UO_4442 (O_4442,N_43655,N_41819);
nor UO_4443 (O_4443,N_41028,N_48529);
and UO_4444 (O_4444,N_40631,N_45356);
nor UO_4445 (O_4445,N_40802,N_43001);
nor UO_4446 (O_4446,N_42822,N_42645);
xnor UO_4447 (O_4447,N_46742,N_44436);
or UO_4448 (O_4448,N_46174,N_46591);
xnor UO_4449 (O_4449,N_48929,N_44839);
and UO_4450 (O_4450,N_48106,N_47839);
xor UO_4451 (O_4451,N_40635,N_44548);
nand UO_4452 (O_4452,N_49258,N_41401);
xor UO_4453 (O_4453,N_47311,N_49956);
nor UO_4454 (O_4454,N_48602,N_40234);
xor UO_4455 (O_4455,N_44288,N_49775);
and UO_4456 (O_4456,N_48312,N_45104);
nand UO_4457 (O_4457,N_44011,N_48207);
and UO_4458 (O_4458,N_46577,N_49329);
nor UO_4459 (O_4459,N_47500,N_40249);
or UO_4460 (O_4460,N_47540,N_43699);
xor UO_4461 (O_4461,N_40849,N_44712);
xor UO_4462 (O_4462,N_48715,N_43393);
nand UO_4463 (O_4463,N_47651,N_43937);
or UO_4464 (O_4464,N_40573,N_46353);
nand UO_4465 (O_4465,N_43313,N_49314);
nand UO_4466 (O_4466,N_41620,N_41157);
or UO_4467 (O_4467,N_43016,N_46759);
or UO_4468 (O_4468,N_49128,N_42962);
nand UO_4469 (O_4469,N_47383,N_45997);
xnor UO_4470 (O_4470,N_42837,N_47558);
nor UO_4471 (O_4471,N_42138,N_44669);
and UO_4472 (O_4472,N_43780,N_48966);
or UO_4473 (O_4473,N_41971,N_41047);
nor UO_4474 (O_4474,N_41120,N_43147);
xor UO_4475 (O_4475,N_48495,N_44478);
xnor UO_4476 (O_4476,N_49017,N_40147);
nor UO_4477 (O_4477,N_40301,N_41056);
nand UO_4478 (O_4478,N_43198,N_45266);
xor UO_4479 (O_4479,N_46476,N_40124);
xnor UO_4480 (O_4480,N_47228,N_44101);
xnor UO_4481 (O_4481,N_48268,N_41314);
nand UO_4482 (O_4482,N_46380,N_45585);
nand UO_4483 (O_4483,N_46722,N_43791);
nor UO_4484 (O_4484,N_47967,N_45613);
xor UO_4485 (O_4485,N_45922,N_47422);
and UO_4486 (O_4486,N_42986,N_42274);
nor UO_4487 (O_4487,N_48222,N_46729);
nand UO_4488 (O_4488,N_49099,N_41566);
xnor UO_4489 (O_4489,N_47494,N_47093);
nand UO_4490 (O_4490,N_40337,N_40940);
xnor UO_4491 (O_4491,N_46770,N_41309);
or UO_4492 (O_4492,N_43673,N_42436);
nor UO_4493 (O_4493,N_42541,N_40009);
and UO_4494 (O_4494,N_41583,N_45943);
or UO_4495 (O_4495,N_49186,N_47223);
nand UO_4496 (O_4496,N_48176,N_41207);
nor UO_4497 (O_4497,N_42156,N_41100);
xnor UO_4498 (O_4498,N_42498,N_44642);
nor UO_4499 (O_4499,N_44758,N_42924);
nand UO_4500 (O_4500,N_48995,N_49894);
and UO_4501 (O_4501,N_42173,N_40541);
nor UO_4502 (O_4502,N_45934,N_49327);
nor UO_4503 (O_4503,N_40386,N_40250);
nand UO_4504 (O_4504,N_49479,N_42042);
xnor UO_4505 (O_4505,N_44028,N_47276);
xnor UO_4506 (O_4506,N_46327,N_47767);
nand UO_4507 (O_4507,N_49535,N_44026);
nand UO_4508 (O_4508,N_41651,N_46563);
or UO_4509 (O_4509,N_48690,N_42328);
nor UO_4510 (O_4510,N_48463,N_41534);
xnor UO_4511 (O_4511,N_48947,N_49790);
xnor UO_4512 (O_4512,N_48650,N_48540);
xnor UO_4513 (O_4513,N_45601,N_47114);
xor UO_4514 (O_4514,N_41740,N_47201);
nor UO_4515 (O_4515,N_46170,N_48398);
or UO_4516 (O_4516,N_47229,N_41889);
nand UO_4517 (O_4517,N_43863,N_43840);
nor UO_4518 (O_4518,N_48841,N_47665);
xor UO_4519 (O_4519,N_49013,N_49200);
or UO_4520 (O_4520,N_49693,N_40847);
nand UO_4521 (O_4521,N_40640,N_41044);
or UO_4522 (O_4522,N_40586,N_46009);
nand UO_4523 (O_4523,N_40772,N_44729);
nor UO_4524 (O_4524,N_45999,N_42345);
nand UO_4525 (O_4525,N_43522,N_46531);
nor UO_4526 (O_4526,N_49835,N_46636);
xnor UO_4527 (O_4527,N_48588,N_44761);
nor UO_4528 (O_4528,N_45616,N_49976);
or UO_4529 (O_4529,N_48023,N_45002);
nor UO_4530 (O_4530,N_46072,N_41215);
or UO_4531 (O_4531,N_45654,N_48426);
xnor UO_4532 (O_4532,N_47562,N_41700);
nand UO_4533 (O_4533,N_47836,N_40081);
nor UO_4534 (O_4534,N_49381,N_42934);
xor UO_4535 (O_4535,N_47576,N_45420);
or UO_4536 (O_4536,N_41163,N_47132);
nor UO_4537 (O_4537,N_48203,N_45233);
or UO_4538 (O_4538,N_45969,N_40714);
or UO_4539 (O_4539,N_45308,N_48584);
nand UO_4540 (O_4540,N_43427,N_46117);
nor UO_4541 (O_4541,N_41332,N_44242);
xor UO_4542 (O_4542,N_46162,N_47736);
nor UO_4543 (O_4543,N_45888,N_40579);
xor UO_4544 (O_4544,N_45970,N_47340);
and UO_4545 (O_4545,N_42705,N_48835);
nand UO_4546 (O_4546,N_41927,N_43657);
nor UO_4547 (O_4547,N_47680,N_49394);
nor UO_4548 (O_4548,N_42148,N_43221);
and UO_4549 (O_4549,N_40447,N_48429);
or UO_4550 (O_4550,N_44295,N_46135);
nor UO_4551 (O_4551,N_40995,N_41551);
nor UO_4552 (O_4552,N_42024,N_47528);
and UO_4553 (O_4553,N_43790,N_47115);
and UO_4554 (O_4554,N_48379,N_41986);
nand UO_4555 (O_4555,N_44561,N_46898);
nand UO_4556 (O_4556,N_40895,N_47819);
xnor UO_4557 (O_4557,N_47766,N_40566);
xor UO_4558 (O_4558,N_49483,N_43692);
nor UO_4559 (O_4559,N_42096,N_42382);
and UO_4560 (O_4560,N_43589,N_49287);
nand UO_4561 (O_4561,N_49493,N_43872);
or UO_4562 (O_4562,N_45304,N_46635);
xnor UO_4563 (O_4563,N_48098,N_46300);
nor UO_4564 (O_4564,N_46627,N_44021);
and UO_4565 (O_4565,N_48590,N_42700);
nor UO_4566 (O_4566,N_40359,N_43726);
or UO_4567 (O_4567,N_44091,N_41710);
or UO_4568 (O_4568,N_42205,N_49692);
or UO_4569 (O_4569,N_45685,N_40093);
nand UO_4570 (O_4570,N_42773,N_42434);
or UO_4571 (O_4571,N_49669,N_43588);
or UO_4572 (O_4572,N_46472,N_45230);
and UO_4573 (O_4573,N_48263,N_47374);
or UO_4574 (O_4574,N_48441,N_43807);
nand UO_4575 (O_4575,N_49082,N_43240);
or UO_4576 (O_4576,N_43245,N_40259);
or UO_4577 (O_4577,N_45624,N_44549);
nor UO_4578 (O_4578,N_49985,N_48211);
xnor UO_4579 (O_4579,N_41514,N_49655);
nand UO_4580 (O_4580,N_40959,N_46726);
and UO_4581 (O_4581,N_47881,N_42675);
nand UO_4582 (O_4582,N_49848,N_40917);
or UO_4583 (O_4583,N_48196,N_49500);
nand UO_4584 (O_4584,N_48546,N_45849);
or UO_4585 (O_4585,N_46387,N_49723);
xnor UO_4586 (O_4586,N_44777,N_42298);
nor UO_4587 (O_4587,N_40212,N_42255);
nand UO_4588 (O_4588,N_40222,N_41988);
xnor UO_4589 (O_4589,N_44075,N_46806);
or UO_4590 (O_4590,N_45493,N_41105);
or UO_4591 (O_4591,N_45772,N_43665);
or UO_4592 (O_4592,N_40004,N_48454);
or UO_4593 (O_4593,N_48573,N_43628);
or UO_4594 (O_4594,N_47529,N_44453);
nor UO_4595 (O_4595,N_45360,N_45257);
nand UO_4596 (O_4596,N_40441,N_46632);
xor UO_4597 (O_4597,N_40875,N_46964);
or UO_4598 (O_4598,N_47816,N_46093);
nand UO_4599 (O_4599,N_47650,N_46594);
xor UO_4600 (O_4600,N_48734,N_44577);
nand UO_4601 (O_4601,N_44785,N_47017);
nor UO_4602 (O_4602,N_42704,N_42199);
nor UO_4603 (O_4603,N_48234,N_48016);
xnor UO_4604 (O_4604,N_46956,N_47901);
nor UO_4605 (O_4605,N_47628,N_41995);
nor UO_4606 (O_4606,N_44903,N_40278);
and UO_4607 (O_4607,N_45463,N_47625);
nor UO_4608 (O_4608,N_47695,N_44209);
and UO_4609 (O_4609,N_46101,N_48847);
nand UO_4610 (O_4610,N_49006,N_48582);
nand UO_4611 (O_4611,N_49925,N_40513);
or UO_4612 (O_4612,N_41503,N_46870);
nor UO_4613 (O_4613,N_40547,N_46153);
or UO_4614 (O_4614,N_40543,N_44186);
nand UO_4615 (O_4615,N_49307,N_46752);
xnor UO_4616 (O_4616,N_41032,N_47240);
nor UO_4617 (O_4617,N_43463,N_44348);
and UO_4618 (O_4618,N_45039,N_46799);
or UO_4619 (O_4619,N_41923,N_41649);
or UO_4620 (O_4620,N_48436,N_47893);
or UO_4621 (O_4621,N_49984,N_41312);
and UO_4622 (O_4622,N_49268,N_46188);
xor UO_4623 (O_4623,N_49302,N_49712);
xor UO_4624 (O_4624,N_43972,N_42510);
and UO_4625 (O_4625,N_42231,N_49789);
nor UO_4626 (O_4626,N_40272,N_47774);
nor UO_4627 (O_4627,N_44833,N_42791);
nor UO_4628 (O_4628,N_46721,N_45093);
nor UO_4629 (O_4629,N_43312,N_47337);
and UO_4630 (O_4630,N_49118,N_48221);
nor UO_4631 (O_4631,N_40735,N_46238);
xnor UO_4632 (O_4632,N_43173,N_48331);
nor UO_4633 (O_4633,N_40219,N_43800);
nor UO_4634 (O_4634,N_44485,N_40022);
and UO_4635 (O_4635,N_43110,N_49180);
xor UO_4636 (O_4636,N_47478,N_43525);
or UO_4637 (O_4637,N_42001,N_41845);
and UO_4638 (O_4638,N_49934,N_42313);
or UO_4639 (O_4639,N_49279,N_42183);
and UO_4640 (O_4640,N_42485,N_47082);
and UO_4641 (O_4641,N_41350,N_41579);
and UO_4642 (O_4642,N_46184,N_47220);
nand UO_4643 (O_4643,N_48982,N_49301);
or UO_4644 (O_4644,N_41023,N_46997);
and UO_4645 (O_4645,N_43139,N_43304);
and UO_4646 (O_4646,N_44144,N_46988);
nor UO_4647 (O_4647,N_42875,N_41682);
or UO_4648 (O_4648,N_48687,N_41843);
or UO_4649 (O_4649,N_46198,N_47204);
nand UO_4650 (O_4650,N_40268,N_46936);
xnor UO_4651 (O_4651,N_40110,N_49973);
nand UO_4652 (O_4652,N_48778,N_46785);
nand UO_4653 (O_4653,N_49513,N_47912);
xor UO_4654 (O_4654,N_47211,N_41885);
and UO_4655 (O_4655,N_47891,N_40644);
nand UO_4656 (O_4656,N_41798,N_46993);
nand UO_4657 (O_4657,N_44850,N_40921);
or UO_4658 (O_4658,N_40255,N_41040);
nand UO_4659 (O_4659,N_45858,N_41096);
or UO_4660 (O_4660,N_47051,N_47139);
or UO_4661 (O_4661,N_45364,N_49877);
nor UO_4662 (O_4662,N_48608,N_47834);
and UO_4663 (O_4663,N_49617,N_49328);
nor UO_4664 (O_4664,N_41826,N_48083);
xor UO_4665 (O_4665,N_46644,N_48531);
nor UO_4666 (O_4666,N_42572,N_49549);
or UO_4667 (O_4667,N_43605,N_46163);
nor UO_4668 (O_4668,N_45336,N_46109);
and UO_4669 (O_4669,N_45026,N_45565);
nor UO_4670 (O_4670,N_44201,N_40064);
nand UO_4671 (O_4671,N_43055,N_41552);
and UO_4672 (O_4672,N_40826,N_43272);
nand UO_4673 (O_4673,N_42044,N_45194);
and UO_4674 (O_4674,N_44876,N_41749);
or UO_4675 (O_4675,N_47635,N_49932);
or UO_4676 (O_4676,N_42582,N_48816);
nor UO_4677 (O_4677,N_49349,N_44449);
nand UO_4678 (O_4678,N_40421,N_49062);
nor UO_4679 (O_4679,N_44000,N_42206);
nor UO_4680 (O_4680,N_40692,N_42299);
and UO_4681 (O_4681,N_45994,N_45196);
or UO_4682 (O_4682,N_41338,N_44197);
nor UO_4683 (O_4683,N_41714,N_40089);
or UO_4684 (O_4684,N_48041,N_40176);
nand UO_4685 (O_4685,N_42787,N_45398);
or UO_4686 (O_4686,N_49873,N_49854);
nor UO_4687 (O_4687,N_45090,N_44432);
and UO_4688 (O_4688,N_46874,N_43127);
or UO_4689 (O_4689,N_45411,N_45637);
nor UO_4690 (O_4690,N_44447,N_43170);
nor UO_4691 (O_4691,N_40469,N_44970);
and UO_4692 (O_4692,N_43354,N_40973);
or UO_4693 (O_4693,N_45358,N_43213);
nor UO_4694 (O_4694,N_48803,N_43940);
nor UO_4695 (O_4695,N_47648,N_47151);
xor UO_4696 (O_4696,N_41392,N_40401);
nand UO_4697 (O_4697,N_41117,N_43010);
xor UO_4698 (O_4698,N_44756,N_44893);
nand UO_4699 (O_4699,N_49254,N_42213);
nand UO_4700 (O_4700,N_43574,N_49860);
nand UO_4701 (O_4701,N_47671,N_47505);
and UO_4702 (O_4702,N_47698,N_43730);
nor UO_4703 (O_4703,N_40318,N_47632);
and UO_4704 (O_4704,N_43441,N_41516);
xor UO_4705 (O_4705,N_47148,N_47742);
nand UO_4706 (O_4706,N_47541,N_49771);
or UO_4707 (O_4707,N_41145,N_47788);
or UO_4708 (O_4708,N_42994,N_47048);
or UO_4709 (O_4709,N_41852,N_43296);
and UO_4710 (O_4710,N_48468,N_40188);
nand UO_4711 (O_4711,N_44371,N_42226);
and UO_4712 (O_4712,N_46537,N_46393);
xnor UO_4713 (O_4713,N_43417,N_41267);
xnor UO_4714 (O_4714,N_45561,N_42641);
xor UO_4715 (O_4715,N_42447,N_40220);
and UO_4716 (O_4716,N_44389,N_46979);
nor UO_4717 (O_4717,N_41550,N_43586);
nor UO_4718 (O_4718,N_46178,N_40070);
xnor UO_4719 (O_4719,N_40982,N_41739);
xor UO_4720 (O_4720,N_44034,N_44342);
nand UO_4721 (O_4721,N_40150,N_40684);
or UO_4722 (O_4722,N_41899,N_47835);
and UO_4723 (O_4723,N_46704,N_45780);
nor UO_4724 (O_4724,N_40529,N_45757);
and UO_4725 (O_4725,N_44848,N_49029);
xnor UO_4726 (O_4726,N_49729,N_47395);
nor UO_4727 (O_4727,N_42083,N_43954);
nand UO_4728 (O_4728,N_45790,N_43543);
or UO_4729 (O_4729,N_41876,N_45938);
and UO_4730 (O_4730,N_42372,N_43328);
xor UO_4731 (O_4731,N_41766,N_41841);
nor UO_4732 (O_4732,N_47100,N_46273);
xnor UO_4733 (O_4733,N_46462,N_40185);
xor UO_4734 (O_4734,N_43265,N_48858);
nor UO_4735 (O_4735,N_49292,N_47865);
and UO_4736 (O_4736,N_47672,N_43927);
nor UO_4737 (O_4737,N_47794,N_48061);
nor UO_4738 (O_4738,N_46400,N_47618);
nor UO_4739 (O_4739,N_46888,N_40908);
nor UO_4740 (O_4740,N_43439,N_41652);
xnor UO_4741 (O_4741,N_48209,N_49168);
or UO_4742 (O_4742,N_40379,N_41685);
nor UO_4743 (O_4743,N_42290,N_49914);
or UO_4744 (O_4744,N_42218,N_49321);
nand UO_4745 (O_4745,N_47947,N_44950);
or UO_4746 (O_4746,N_48897,N_43929);
nor UO_4747 (O_4747,N_44316,N_45629);
or UO_4748 (O_4748,N_45430,N_46102);
xor UO_4749 (O_4749,N_48999,N_44227);
and UO_4750 (O_4750,N_41590,N_48909);
nor UO_4751 (O_4751,N_45241,N_44569);
and UO_4752 (O_4752,N_43237,N_44817);
or UO_4753 (O_4753,N_40221,N_48708);
and UO_4754 (O_4754,N_49291,N_45085);
and UO_4755 (O_4755,N_46179,N_43853);
xor UO_4756 (O_4756,N_40471,N_43070);
xor UO_4757 (O_4757,N_42122,N_41524);
or UO_4758 (O_4758,N_45202,N_49577);
nand UO_4759 (O_4759,N_45405,N_45189);
nor UO_4760 (O_4760,N_40016,N_46975);
or UO_4761 (O_4761,N_49454,N_46656);
nor UO_4762 (O_4762,N_42971,N_40812);
or UO_4763 (O_4763,N_43659,N_44480);
and UO_4764 (O_4764,N_40086,N_45840);
nand UO_4765 (O_4765,N_49817,N_43638);
xnor UO_4766 (O_4766,N_45149,N_41495);
xnor UO_4767 (O_4767,N_48621,N_45069);
nand UO_4768 (O_4768,N_43782,N_49852);
nor UO_4769 (O_4769,N_47502,N_41041);
xnor UO_4770 (O_4770,N_49097,N_43707);
xnor UO_4771 (O_4771,N_46588,N_44698);
xnor UO_4772 (O_4772,N_45879,N_41748);
and UO_4773 (O_4773,N_48877,N_46350);
xor UO_4774 (O_4774,N_49446,N_43224);
xor UO_4775 (O_4775,N_43829,N_46669);
nand UO_4776 (O_4776,N_48526,N_40047);
nor UO_4777 (O_4777,N_46827,N_43461);
nand UO_4778 (O_4778,N_43966,N_42294);
and UO_4779 (O_4779,N_40521,N_46258);
xor UO_4780 (O_4780,N_48220,N_41437);
and UO_4781 (O_4781,N_47382,N_42054);
nor UO_4782 (O_4782,N_42754,N_45129);
or UO_4783 (O_4783,N_42254,N_48445);
nor UO_4784 (O_4784,N_45419,N_41560);
nor UO_4785 (O_4785,N_40698,N_46865);
nor UO_4786 (O_4786,N_46915,N_43721);
nor UO_4787 (O_4787,N_42706,N_43744);
nand UO_4788 (O_4788,N_40131,N_45047);
xor UO_4789 (O_4789,N_49673,N_42402);
nand UO_4790 (O_4790,N_47830,N_43946);
or UO_4791 (O_4791,N_41206,N_40831);
or UO_4792 (O_4792,N_45787,N_46510);
or UO_4793 (O_4793,N_46507,N_43861);
xor UO_4794 (O_4794,N_44483,N_46010);
or UO_4795 (O_4795,N_46589,N_47647);
nor UO_4796 (O_4796,N_44666,N_47043);
nand UO_4797 (O_4797,N_48070,N_45981);
or UO_4798 (O_4798,N_46061,N_45525);
xnor UO_4799 (O_4799,N_40267,N_44382);
nor UO_4800 (O_4800,N_43287,N_41031);
nor UO_4801 (O_4801,N_42763,N_49639);
and UO_4802 (O_4802,N_47392,N_49234);
nor UO_4803 (O_4803,N_40497,N_41052);
and UO_4804 (O_4804,N_42782,N_45368);
or UO_4805 (O_4805,N_46321,N_48080);
nand UO_4806 (O_4806,N_40201,N_47355);
and UO_4807 (O_4807,N_48721,N_40273);
nor UO_4808 (O_4808,N_41870,N_49977);
and UO_4809 (O_4809,N_47764,N_41708);
nand UO_4810 (O_4810,N_40063,N_47014);
or UO_4811 (O_4811,N_42508,N_43476);
xor UO_4812 (O_4812,N_43754,N_49590);
or UO_4813 (O_4813,N_40458,N_48295);
xnor UO_4814 (O_4814,N_48735,N_44736);
or UO_4815 (O_4815,N_42384,N_46800);
xor UO_4816 (O_4816,N_47566,N_42951);
nor UO_4817 (O_4817,N_42008,N_48169);
nand UO_4818 (O_4818,N_42737,N_41328);
xor UO_4819 (O_4819,N_42666,N_48199);
and UO_4820 (O_4820,N_48595,N_48046);
or UO_4821 (O_4821,N_49886,N_45458);
nand UO_4822 (O_4822,N_40031,N_41881);
and UO_4823 (O_4823,N_49439,N_43041);
nor UO_4824 (O_4824,N_44080,N_49623);
nand UO_4825 (O_4825,N_49896,N_46436);
nand UO_4826 (O_4826,N_49496,N_46801);
nor UO_4827 (O_4827,N_48717,N_41341);
and UO_4828 (O_4828,N_42142,N_46002);
nor UO_4829 (O_4829,N_49752,N_42724);
xor UO_4830 (O_4830,N_47911,N_47013);
and UO_4831 (O_4831,N_43282,N_45832);
or UO_4832 (O_4832,N_49420,N_41384);
or UO_4833 (O_4833,N_47393,N_46493);
xnor UO_4834 (O_4834,N_46362,N_43492);
nor UO_4835 (O_4835,N_45618,N_48403);
nor UO_4836 (O_4836,N_42515,N_40751);
and UO_4837 (O_4837,N_41837,N_44987);
xnor UO_4838 (O_4838,N_47526,N_47316);
and UO_4839 (O_4839,N_44566,N_40309);
nor UO_4840 (O_4840,N_48177,N_45263);
and UO_4841 (O_4841,N_46312,N_42946);
or UO_4842 (O_4842,N_43216,N_44309);
nor UO_4843 (O_4843,N_46617,N_42360);
and UO_4844 (O_4844,N_40539,N_40557);
xnor UO_4845 (O_4845,N_47784,N_48662);
nor UO_4846 (O_4846,N_49702,N_44493);
and UO_4847 (O_4847,N_42716,N_49744);
nand UO_4848 (O_4848,N_48876,N_41140);
nor UO_4849 (O_4849,N_44763,N_46790);
nand UO_4850 (O_4850,N_41319,N_49951);
or UO_4851 (O_4851,N_46488,N_42036);
or UO_4852 (O_4852,N_44299,N_45174);
or UO_4853 (O_4853,N_41936,N_42388);
or UO_4854 (O_4854,N_41073,N_41295);
nand UO_4855 (O_4855,N_40069,N_40632);
nor UO_4856 (O_4856,N_49993,N_40378);
xor UO_4857 (O_4857,N_43162,N_48039);
nand UO_4858 (O_4858,N_42601,N_43130);
or UO_4859 (O_4859,N_40550,N_49056);
nand UO_4860 (O_4860,N_40771,N_44161);
nand UO_4861 (O_4861,N_49455,N_43018);
nor UO_4862 (O_4862,N_43884,N_48979);
nand UO_4863 (O_4863,N_43468,N_45889);
xnor UO_4864 (O_4864,N_44414,N_45095);
xor UO_4865 (O_4865,N_45048,N_47718);
or UO_4866 (O_4866,N_44786,N_41250);
nor UO_4867 (O_4867,N_42151,N_47069);
nor UO_4868 (O_4868,N_42265,N_42547);
or UO_4869 (O_4869,N_47997,N_49164);
or UO_4870 (O_4870,N_40159,N_43634);
nor UO_4871 (O_4871,N_40506,N_47879);
xor UO_4872 (O_4872,N_45813,N_49633);
nand UO_4873 (O_4873,N_45006,N_48193);
xor UO_4874 (O_4874,N_40434,N_48811);
xnor UO_4875 (O_4875,N_44172,N_43431);
and UO_4876 (O_4876,N_41104,N_41744);
nor UO_4877 (O_4877,N_41301,N_49495);
or UO_4878 (O_4878,N_42714,N_42394);
xnor UO_4879 (O_4879,N_45018,N_41135);
and UO_4880 (O_4880,N_48544,N_48243);
xor UO_4881 (O_4881,N_49815,N_40068);
or UO_4882 (O_4882,N_40500,N_44673);
xor UO_4883 (O_4883,N_42901,N_49156);
xnor UO_4884 (O_4884,N_49884,N_42613);
nor UO_4885 (O_4885,N_43573,N_49116);
or UO_4886 (O_4886,N_45120,N_45752);
xnor UO_4887 (O_4887,N_47285,N_44952);
nor UO_4888 (O_4888,N_44087,N_41867);
nor UO_4889 (O_4889,N_41996,N_49004);
or UO_4890 (O_4890,N_45799,N_42936);
and UO_4891 (O_4891,N_42587,N_40669);
nor UO_4892 (O_4892,N_46777,N_48821);
xnor UO_4893 (O_4893,N_40502,N_45145);
or UO_4894 (O_4894,N_45963,N_48369);
and UO_4895 (O_4895,N_46679,N_41067);
and UO_4896 (O_4896,N_45738,N_40078);
nor UO_4897 (O_4897,N_46180,N_44552);
nand UO_4898 (O_4898,N_46315,N_47854);
nand UO_4899 (O_4899,N_41160,N_44984);
or UO_4900 (O_4900,N_43436,N_48900);
or UO_4901 (O_4901,N_48179,N_41151);
xnor UO_4902 (O_4902,N_42871,N_45852);
xor UO_4903 (O_4903,N_47754,N_45390);
nor UO_4904 (O_4904,N_48509,N_42558);
and UO_4905 (O_4905,N_40419,N_43483);
nand UO_4906 (O_4906,N_41718,N_42497);
or UO_4907 (O_4907,N_48491,N_47887);
and UO_4908 (O_4908,N_41330,N_47303);
nor UO_4909 (O_4909,N_40107,N_40906);
xor UO_4910 (O_4910,N_41248,N_40605);
nor UO_4911 (O_4911,N_42031,N_46687);
xnor UO_4912 (O_4912,N_45702,N_41345);
nor UO_4913 (O_4913,N_45818,N_46013);
or UO_4914 (O_4914,N_49393,N_48701);
and UO_4915 (O_4915,N_43608,N_45432);
nor UO_4916 (O_4916,N_47449,N_48668);
xnor UO_4917 (O_4917,N_40512,N_40331);
or UO_4918 (O_4918,N_42446,N_48726);
and UO_4919 (O_4919,N_41214,N_42702);
xnor UO_4920 (O_4920,N_47169,N_42390);
and UO_4921 (O_4921,N_44320,N_45578);
nand UO_4922 (O_4922,N_42873,N_44058);
nand UO_4923 (O_4923,N_43602,N_45131);
xor UO_4924 (O_4924,N_49928,N_41756);
or UO_4925 (O_4925,N_46217,N_46323);
and UO_4926 (O_4926,N_49290,N_43528);
xor UO_4927 (O_4927,N_41190,N_45330);
nand UO_4928 (O_4928,N_41978,N_44461);
nand UO_4929 (O_4929,N_48917,N_49445);
or UO_4930 (O_4930,N_44355,N_48911);
nor UO_4931 (O_4931,N_40883,N_40839);
nand UO_4932 (O_4932,N_43083,N_42904);
and UO_4933 (O_4933,N_47210,N_44907);
nor UO_4934 (O_4934,N_41693,N_43234);
nand UO_4935 (O_4935,N_47071,N_42957);
nor UO_4936 (O_4936,N_46792,N_40621);
xor UO_4937 (O_4937,N_41217,N_42881);
nand UO_4938 (O_4938,N_42571,N_47295);
and UO_4939 (O_4939,N_43941,N_42422);
nor UO_4940 (O_4940,N_41500,N_41144);
or UO_4941 (O_4941,N_43254,N_42720);
nor UO_4942 (O_4942,N_49851,N_44291);
nor UO_4943 (O_4943,N_42983,N_44715);
nor UO_4944 (O_4944,N_43898,N_41969);
or UO_4945 (O_4945,N_46701,N_46779);
xnor UO_4946 (O_4946,N_43201,N_48340);
or UO_4947 (O_4947,N_46732,N_46543);
or UO_4948 (O_4948,N_49525,N_43309);
or UO_4949 (O_4949,N_49100,N_40132);
nand UO_4950 (O_4950,N_46343,N_48322);
nand UO_4951 (O_4951,N_49018,N_42203);
and UO_4952 (O_4952,N_47191,N_43550);
or UO_4953 (O_4953,N_48088,N_43160);
xor UO_4954 (O_4954,N_41797,N_49431);
xnor UO_4955 (O_4955,N_41920,N_41394);
or UO_4956 (O_4956,N_49863,N_41896);
xnor UO_4957 (O_4957,N_44412,N_42282);
and UO_4958 (O_4958,N_47843,N_40457);
xor UO_4959 (O_4959,N_44314,N_44158);
xor UO_4960 (O_4960,N_41380,N_45220);
nor UO_4961 (O_4961,N_45270,N_43297);
nand UO_4962 (O_4962,N_46508,N_42761);
nand UO_4963 (O_4963,N_41865,N_41941);
and UO_4964 (O_4964,N_47570,N_48605);
nand UO_4965 (O_4965,N_40994,N_41057);
nand UO_4966 (O_4966,N_43357,N_46299);
nand UO_4967 (O_4967,N_40505,N_44273);
nor UO_4968 (O_4968,N_49359,N_47061);
nor UO_4969 (O_4969,N_47342,N_42413);
nand UO_4970 (O_4970,N_47984,N_49574);
or UO_4971 (O_4971,N_48480,N_46382);
and UO_4972 (O_4972,N_44441,N_41264);
nand UO_4973 (O_4973,N_45548,N_49751);
xor UO_4974 (O_4974,N_44886,N_45369);
and UO_4975 (O_4975,N_48505,N_48774);
nor UO_4976 (O_4976,N_47890,N_44737);
xor UO_4977 (O_4977,N_43232,N_40963);
nand UO_4978 (O_4978,N_44565,N_42415);
nand UO_4979 (O_4979,N_42135,N_44505);
and UO_4980 (O_4980,N_49709,N_45439);
xnor UO_4981 (O_4981,N_48124,N_40976);
and UO_4982 (O_4982,N_49726,N_42967);
and UO_4983 (O_4983,N_49619,N_43597);
and UO_4984 (O_4984,N_49154,N_47946);
nand UO_4985 (O_4985,N_46750,N_41334);
nor UO_4986 (O_4986,N_47716,N_43737);
and UO_4987 (O_4987,N_47369,N_47165);
or UO_4988 (O_4988,N_43410,N_40981);
nor UO_4989 (O_4989,N_46601,N_46826);
nor UO_4990 (O_4990,N_43915,N_45699);
nor UO_4991 (O_4991,N_48025,N_49107);
and UO_4992 (O_4992,N_49978,N_41612);
nor UO_4993 (O_4993,N_41229,N_46502);
and UO_4994 (O_4994,N_48266,N_43451);
or UO_4995 (O_4995,N_45329,N_44481);
nand UO_4996 (O_4996,N_40058,N_49856);
nor UO_4997 (O_4997,N_49247,N_46322);
xnor UO_4998 (O_4998,N_40815,N_45673);
nand UO_4999 (O_4999,N_40887,N_40989);
endmodule