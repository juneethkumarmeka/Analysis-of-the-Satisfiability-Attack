module basic_2500_25000_3000_8_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_153,In_1537);
xnor U1 (N_1,In_1210,In_640);
and U2 (N_2,In_2362,In_370);
xor U3 (N_3,In_1971,In_1133);
nand U4 (N_4,In_1858,In_41);
nor U5 (N_5,In_2045,In_499);
xnor U6 (N_6,In_1279,In_1068);
nand U7 (N_7,In_553,In_20);
or U8 (N_8,In_134,In_1415);
nand U9 (N_9,In_1373,In_118);
or U10 (N_10,In_1643,In_2289);
nor U11 (N_11,In_149,In_1556);
nand U12 (N_12,In_1466,In_2429);
nor U13 (N_13,In_1735,In_29);
xor U14 (N_14,In_1629,In_1314);
or U15 (N_15,In_732,In_424);
or U16 (N_16,In_457,In_855);
nand U17 (N_17,In_1663,In_1396);
or U18 (N_18,In_616,In_1368);
nand U19 (N_19,In_1533,In_696);
xnor U20 (N_20,In_878,In_1823);
nor U21 (N_21,In_22,In_2);
nor U22 (N_22,In_1132,In_1265);
or U23 (N_23,In_633,In_915);
nor U24 (N_24,In_668,In_1728);
or U25 (N_25,In_1755,In_290);
xnor U26 (N_26,In_48,In_1341);
or U27 (N_27,In_1790,In_903);
xor U28 (N_28,In_1019,In_2485);
xnor U29 (N_29,In_1099,In_493);
xnor U30 (N_30,In_1912,In_1953);
and U31 (N_31,In_156,In_219);
or U32 (N_32,In_526,In_842);
or U33 (N_33,In_1304,In_1448);
or U34 (N_34,In_598,In_433);
xor U35 (N_35,In_7,In_1468);
nor U36 (N_36,In_1390,In_1369);
and U37 (N_37,In_2334,In_185);
and U38 (N_38,In_1416,In_1159);
and U39 (N_39,In_1921,In_250);
nor U40 (N_40,In_2379,In_1385);
nand U41 (N_41,In_154,In_1753);
xnor U42 (N_42,In_1324,In_2342);
and U43 (N_43,In_913,In_1577);
and U44 (N_44,In_2156,In_2399);
xor U45 (N_45,In_438,In_2455);
and U46 (N_46,In_2041,In_308);
and U47 (N_47,In_1425,In_170);
nand U48 (N_48,In_2110,In_2099);
and U49 (N_49,In_267,In_1748);
and U50 (N_50,In_994,In_2032);
xor U51 (N_51,In_2471,In_2422);
nor U52 (N_52,In_284,In_2168);
xor U53 (N_53,In_343,In_1870);
or U54 (N_54,In_396,In_1072);
nand U55 (N_55,In_248,In_2354);
or U56 (N_56,In_548,In_751);
or U57 (N_57,In_722,In_958);
nor U58 (N_58,In_2194,In_1006);
or U59 (N_59,In_1609,In_1082);
or U60 (N_60,In_2076,In_1137);
or U61 (N_61,In_1836,In_675);
xnor U62 (N_62,In_2237,In_2199);
nand U63 (N_63,In_2358,In_1933);
nand U64 (N_64,In_737,In_1796);
nor U65 (N_65,In_1786,In_2177);
xnor U66 (N_66,In_157,In_2019);
or U67 (N_67,In_560,In_1856);
and U68 (N_68,In_1597,In_1482);
and U69 (N_69,In_2190,In_115);
and U70 (N_70,In_1538,In_479);
nand U71 (N_71,In_2267,In_1372);
nor U72 (N_72,In_1767,In_1391);
xnor U73 (N_73,In_1920,In_1807);
nand U74 (N_74,In_410,In_1325);
and U75 (N_75,In_1282,In_851);
xnor U76 (N_76,In_2273,In_533);
and U77 (N_77,In_1426,In_1861);
or U78 (N_78,In_2486,In_1816);
nand U79 (N_79,In_1370,In_1128);
nor U80 (N_80,In_1393,In_949);
nand U81 (N_81,In_2068,In_1305);
nand U82 (N_82,In_1860,In_801);
or U83 (N_83,In_1313,In_2048);
nand U84 (N_84,In_2424,In_2265);
and U85 (N_85,In_1129,In_376);
or U86 (N_86,In_2108,In_838);
and U87 (N_87,In_2003,In_1526);
and U88 (N_88,In_2166,In_1378);
or U89 (N_89,In_2097,In_2414);
nand U90 (N_90,In_872,In_1020);
nand U91 (N_91,In_2274,In_670);
xor U92 (N_92,In_247,In_993);
xnor U93 (N_93,In_991,In_2347);
nor U94 (N_94,In_2320,In_275);
nor U95 (N_95,In_2253,In_1736);
nand U96 (N_96,In_368,In_1881);
xor U97 (N_97,In_1238,In_719);
nor U98 (N_98,In_46,In_920);
xnor U99 (N_99,In_1605,In_1254);
nand U100 (N_100,In_918,In_2114);
xor U101 (N_101,In_681,In_362);
and U102 (N_102,In_459,In_1443);
and U103 (N_103,In_324,In_1607);
nor U104 (N_104,In_179,In_217);
or U105 (N_105,In_1659,In_1316);
xor U106 (N_106,In_2390,In_2409);
nand U107 (N_107,In_1059,In_1996);
nand U108 (N_108,In_1959,In_2262);
xor U109 (N_109,In_2492,In_518);
xnor U110 (N_110,In_705,In_1015);
nand U111 (N_111,In_371,In_1563);
and U112 (N_112,In_1321,In_1772);
nor U113 (N_113,In_2346,In_1938);
and U114 (N_114,In_1768,In_1797);
xnor U115 (N_115,In_1815,In_956);
nand U116 (N_116,In_1242,In_1653);
xnor U117 (N_117,In_1449,In_58);
and U118 (N_118,In_184,In_2195);
or U119 (N_119,In_590,In_2119);
or U120 (N_120,In_114,In_1584);
and U121 (N_121,In_861,In_849);
xnor U122 (N_122,In_1199,In_1096);
or U123 (N_123,In_1939,In_1339);
nand U124 (N_124,In_565,In_1734);
and U125 (N_125,In_1061,In_662);
or U126 (N_126,In_916,In_1338);
nand U127 (N_127,In_1866,In_1724);
nor U128 (N_128,In_2152,In_151);
xnor U129 (N_129,In_2225,In_1170);
nand U130 (N_130,In_1360,In_1737);
or U131 (N_131,In_572,In_191);
and U132 (N_132,In_2078,In_1923);
and U133 (N_133,In_1271,In_1947);
xor U134 (N_134,In_2123,In_2293);
xor U135 (N_135,In_1520,In_1917);
nand U136 (N_136,In_1037,In_1453);
and U137 (N_137,In_1273,In_1214);
or U138 (N_138,In_615,In_912);
nand U139 (N_139,In_1495,In_1299);
nor U140 (N_140,In_305,In_1875);
nor U141 (N_141,In_144,In_1165);
nand U142 (N_142,In_531,In_1596);
and U143 (N_143,In_1804,In_1429);
nor U144 (N_144,In_2440,In_1149);
or U145 (N_145,In_2472,In_887);
nor U146 (N_146,In_741,In_1490);
nand U147 (N_147,In_1513,In_661);
or U148 (N_148,In_815,In_885);
nand U149 (N_149,In_784,In_655);
nand U150 (N_150,In_2474,In_2007);
nand U151 (N_151,In_713,In_1435);
or U152 (N_152,In_523,In_954);
xor U153 (N_153,In_847,In_1806);
and U154 (N_154,In_657,In_2477);
and U155 (N_155,In_972,In_1264);
and U156 (N_156,In_116,In_299);
xor U157 (N_157,In_852,In_871);
or U158 (N_158,In_1418,In_1451);
and U159 (N_159,In_1579,In_2340);
or U160 (N_160,In_2407,In_778);
xnor U161 (N_161,In_1410,In_1855);
nand U162 (N_162,In_365,In_1898);
xnor U163 (N_163,In_987,In_419);
and U164 (N_164,In_1144,In_552);
and U165 (N_165,In_1913,In_388);
nor U166 (N_166,In_1446,In_2155);
or U167 (N_167,In_1140,In_1180);
and U168 (N_168,In_2404,In_1585);
xnor U169 (N_169,In_2174,In_605);
and U170 (N_170,In_1143,In_2268);
or U171 (N_171,In_1723,In_1460);
nor U172 (N_172,In_864,In_1572);
or U173 (N_173,In_937,In_2207);
nand U174 (N_174,In_409,In_168);
and U175 (N_175,In_1141,In_59);
xnor U176 (N_176,In_1750,In_820);
xor U177 (N_177,In_2088,In_1261);
xnor U178 (N_178,In_599,In_1280);
and U179 (N_179,In_2396,In_1039);
xor U180 (N_180,In_2109,In_233);
or U181 (N_181,In_102,In_1903);
and U182 (N_182,In_919,In_2370);
xnor U183 (N_183,In_1908,In_265);
and U184 (N_184,In_1207,In_2256);
nor U185 (N_185,In_1820,In_1948);
nor U186 (N_186,In_550,In_1877);
nor U187 (N_187,In_1650,In_829);
and U188 (N_188,In_1709,In_2187);
xnor U189 (N_189,In_1127,In_1094);
xor U190 (N_190,In_1691,In_844);
xor U191 (N_191,In_1887,In_2116);
or U192 (N_192,In_1553,In_1949);
nor U193 (N_193,In_1978,In_812);
and U194 (N_194,In_2304,In_47);
nor U195 (N_195,In_418,In_1827);
xnor U196 (N_196,In_1671,In_1116);
nand U197 (N_197,In_425,In_930);
or U198 (N_198,In_873,In_2022);
nor U199 (N_199,In_1555,In_360);
and U200 (N_200,In_2463,In_692);
nand U201 (N_201,In_2427,In_728);
nand U202 (N_202,In_1999,In_1994);
nor U203 (N_203,In_1102,In_1479);
nor U204 (N_204,In_2281,In_1248);
and U205 (N_205,In_860,In_8);
and U206 (N_206,In_458,In_75);
and U207 (N_207,In_2292,In_16);
nor U208 (N_208,In_2460,In_1894);
or U209 (N_209,In_1480,In_2306);
nand U210 (N_210,In_122,In_543);
or U211 (N_211,In_1439,In_1486);
nand U212 (N_212,In_28,In_799);
nand U213 (N_213,In_2352,In_165);
xor U214 (N_214,In_2013,In_462);
xnor U215 (N_215,In_1871,In_924);
nand U216 (N_216,In_2009,In_1067);
and U217 (N_217,In_2481,In_1963);
or U218 (N_218,In_223,In_752);
nand U219 (N_219,In_630,In_1950);
nor U220 (N_220,In_2498,In_1168);
and U221 (N_221,In_465,In_619);
and U222 (N_222,In_902,In_1529);
nand U223 (N_223,In_2196,In_271);
nand U224 (N_224,In_310,In_708);
xnor U225 (N_225,In_883,In_487);
nand U226 (N_226,In_1358,In_1157);
and U227 (N_227,In_1547,In_1590);
and U228 (N_228,In_1826,In_1665);
nor U229 (N_229,In_2121,In_868);
nor U230 (N_230,In_2066,In_515);
nor U231 (N_231,In_610,In_2435);
and U232 (N_232,In_1632,In_1198);
nor U233 (N_233,In_2457,In_2375);
xor U234 (N_234,In_1893,In_1303);
and U235 (N_235,In_338,In_266);
and U236 (N_236,In_1295,In_146);
nor U237 (N_237,In_745,In_824);
nand U238 (N_238,In_227,In_1186);
xnor U239 (N_239,In_1326,In_1668);
xor U240 (N_240,In_648,In_2303);
xnor U241 (N_241,In_2489,In_42);
xor U242 (N_242,In_166,In_774);
and U243 (N_243,In_2131,In_392);
nand U244 (N_244,In_975,In_2201);
or U245 (N_245,In_431,In_1405);
or U246 (N_246,In_967,In_2033);
xor U247 (N_247,In_1621,In_359);
xor U248 (N_248,In_2077,In_323);
or U249 (N_249,In_1987,In_637);
and U250 (N_250,In_2333,In_879);
or U251 (N_251,In_316,In_612);
or U252 (N_252,In_914,In_21);
nor U253 (N_253,In_693,In_813);
nand U254 (N_254,In_990,In_1746);
xnor U255 (N_255,In_161,In_2251);
and U256 (N_256,In_772,In_2192);
nand U257 (N_257,In_1614,In_743);
xnor U258 (N_258,In_672,In_143);
nand U259 (N_259,In_2193,In_2208);
or U260 (N_260,In_2327,In_1840);
xnor U261 (N_261,In_1452,In_817);
or U262 (N_262,In_1383,In_1337);
and U263 (N_263,In_298,In_581);
and U264 (N_264,In_5,In_1525);
xor U265 (N_265,In_1883,In_1260);
xnor U266 (N_266,In_2247,In_2428);
and U267 (N_267,In_1689,In_0);
or U268 (N_268,In_2025,In_2072);
and U269 (N_269,In_1275,In_2316);
nor U270 (N_270,In_241,In_1064);
or U271 (N_271,In_196,In_768);
xnor U272 (N_272,In_1110,In_1907);
and U273 (N_273,In_1192,In_1161);
nand U274 (N_274,In_900,In_1681);
nor U275 (N_275,In_1459,In_120);
xnor U276 (N_276,In_1002,In_1450);
or U277 (N_277,In_1436,In_1009);
and U278 (N_278,In_322,In_839);
nand U279 (N_279,In_2240,In_2243);
or U280 (N_280,In_2000,In_2015);
xor U281 (N_281,In_1212,In_72);
nand U282 (N_282,In_43,In_1989);
and U283 (N_283,In_2408,In_1524);
or U284 (N_284,In_329,In_910);
xor U285 (N_285,In_1889,In_272);
and U286 (N_286,In_1980,In_1362);
xnor U287 (N_287,In_1763,In_1612);
nor U288 (N_288,In_1702,In_1924);
nand U289 (N_289,In_158,In_1708);
nor U290 (N_290,In_653,In_2439);
nor U291 (N_291,In_1536,In_1813);
and U292 (N_292,In_2146,In_625);
xor U293 (N_293,In_632,In_1489);
or U294 (N_294,In_595,In_353);
nor U295 (N_295,In_1592,In_1773);
xnor U296 (N_296,In_1139,In_755);
nor U297 (N_297,In_1431,In_2220);
or U298 (N_298,In_629,In_1550);
and U299 (N_299,In_1035,In_73);
or U300 (N_300,In_1070,In_344);
nand U301 (N_301,In_470,In_1003);
nor U302 (N_302,In_2211,In_2248);
nor U303 (N_303,In_1432,In_69);
and U304 (N_304,In_592,In_1058);
nand U305 (N_305,In_702,In_2028);
and U306 (N_306,In_45,In_2266);
nand U307 (N_307,In_330,In_1902);
or U308 (N_308,In_1849,In_1005);
and U309 (N_309,In_2223,In_1501);
or U310 (N_310,In_969,In_56);
or U311 (N_311,In_1069,In_82);
xnor U312 (N_312,In_1098,In_1718);
or U313 (N_313,In_210,In_1473);
nor U314 (N_314,In_391,In_2239);
nand U315 (N_315,In_525,In_2126);
xor U316 (N_316,In_1943,In_2449);
nor U317 (N_317,In_1984,In_2314);
nor U318 (N_318,In_1222,In_1052);
or U319 (N_319,In_757,In_769);
or U320 (N_320,In_224,In_2117);
and U321 (N_321,In_571,In_881);
or U322 (N_322,In_1328,In_1784);
or U323 (N_323,In_1623,In_1729);
nor U324 (N_324,In_2005,In_489);
nand U325 (N_325,In_2210,In_608);
nor U326 (N_326,In_382,In_31);
nand U327 (N_327,In_289,In_1043);
xor U328 (N_328,In_2487,In_1589);
xnor U329 (N_329,In_108,In_1617);
nand U330 (N_330,In_907,In_1941);
xnor U331 (N_331,In_213,In_2483);
nor U332 (N_332,In_1483,In_1906);
nand U333 (N_333,In_2325,In_1666);
xor U334 (N_334,In_78,In_1915);
nor U335 (N_335,In_2016,In_1174);
xor U336 (N_336,In_1056,In_2444);
or U337 (N_337,In_1970,In_1371);
xnor U338 (N_338,In_1101,In_393);
nand U339 (N_339,In_1895,In_1673);
xor U340 (N_340,In_2468,In_2291);
xor U341 (N_341,In_1071,In_1720);
or U342 (N_342,In_1825,In_1966);
nand U343 (N_343,In_1967,In_2226);
nor U344 (N_344,In_1437,In_1365);
nand U345 (N_345,In_495,In_83);
and U346 (N_346,In_160,In_351);
xor U347 (N_347,In_1669,In_446);
and U348 (N_348,In_2259,In_1769);
xor U349 (N_349,In_1231,In_203);
xor U350 (N_350,In_1352,In_68);
nand U351 (N_351,In_1511,In_23);
nor U352 (N_352,In_2158,In_1350);
or U353 (N_353,In_1879,In_422);
nand U354 (N_354,In_206,In_1188);
or U355 (N_355,In_201,In_911);
nand U356 (N_356,In_1626,In_2418);
nand U357 (N_357,In_2360,In_2105);
nor U358 (N_358,In_112,In_1808);
nand U359 (N_359,In_2386,In_138);
and U360 (N_360,In_2214,In_1692);
or U361 (N_361,In_2172,In_997);
nand U362 (N_362,In_1685,In_482);
xor U363 (N_363,In_231,In_906);
xor U364 (N_364,In_1089,In_889);
and U365 (N_365,In_398,In_1677);
xor U366 (N_366,In_593,In_1843);
and U367 (N_367,In_1134,In_1738);
nand U368 (N_368,In_1042,In_2298);
xor U369 (N_369,In_390,In_944);
or U370 (N_370,In_2153,In_2496);
and U371 (N_371,In_1310,In_2217);
nor U372 (N_372,In_1249,In_726);
nand U373 (N_373,In_1945,In_2389);
xor U374 (N_374,In_2378,In_1988);
xnor U375 (N_375,In_1688,In_1591);
xor U376 (N_376,In_1095,In_1497);
nor U377 (N_377,In_291,In_1931);
xor U378 (N_378,In_1029,In_1789);
nand U379 (N_379,In_420,In_567);
nor U380 (N_380,In_894,In_837);
nand U381 (N_381,In_1674,In_2335);
or U382 (N_382,In_643,In_1751);
nand U383 (N_383,In_586,In_254);
or U384 (N_384,In_2415,In_237);
and U385 (N_385,In_205,In_614);
nor U386 (N_386,In_1884,In_955);
nand U387 (N_387,In_962,In_1266);
and U388 (N_388,In_507,In_1055);
and U389 (N_389,In_1256,In_2343);
nor U390 (N_390,In_415,In_2283);
nor U391 (N_391,In_1298,In_1929);
nor U392 (N_392,In_1509,In_1783);
nand U393 (N_393,In_946,In_1166);
nand U394 (N_394,In_428,In_270);
and U395 (N_395,In_803,In_355);
nand U396 (N_396,In_1441,In_113);
or U397 (N_397,In_321,In_1108);
nand U398 (N_398,In_1834,In_1657);
nand U399 (N_399,In_1874,In_983);
nand U400 (N_400,In_1031,In_337);
or U401 (N_401,In_600,In_498);
nor U402 (N_402,In_2018,In_357);
nor U403 (N_403,In_1492,In_1232);
or U404 (N_404,In_1976,In_226);
or U405 (N_405,In_1974,In_574);
nor U406 (N_406,In_2493,In_1175);
and U407 (N_407,In_2055,In_1900);
nand U408 (N_408,In_55,In_1594);
or U409 (N_409,In_1184,In_1507);
nand U410 (N_410,In_1474,In_235);
and U411 (N_411,In_1284,In_1481);
nor U412 (N_412,In_327,In_2456);
nor U413 (N_413,In_2398,In_1331);
xor U414 (N_414,In_1580,In_819);
nor U415 (N_415,In_1956,In_2180);
nand U416 (N_416,In_840,In_2170);
and U417 (N_417,In_301,In_1540);
nor U418 (N_418,In_2056,In_230);
nand U419 (N_419,In_1206,In_1754);
nor U420 (N_420,In_256,In_1183);
nor U421 (N_421,In_1701,In_1091);
xnor U422 (N_422,In_806,In_1560);
nor U423 (N_423,In_426,In_1575);
and U424 (N_424,In_2138,In_1027);
xnor U425 (N_425,In_1595,In_1542);
nand U426 (N_426,In_2495,In_2423);
nand U427 (N_427,In_1106,In_1711);
nor U428 (N_428,In_623,In_37);
nand U429 (N_429,In_1998,In_1257);
nand U430 (N_430,In_2085,In_239);
nor U431 (N_431,In_94,In_1152);
or U432 (N_432,In_14,In_935);
xnor U433 (N_433,In_486,In_1211);
nor U434 (N_434,In_472,In_1100);
and U435 (N_435,In_874,In_1777);
or U436 (N_436,In_859,In_843);
xnor U437 (N_437,In_826,In_1641);
xnor U438 (N_438,In_2059,In_1011);
and U439 (N_439,In_609,In_2042);
and U440 (N_440,In_1686,In_995);
nand U441 (N_441,In_897,In_501);
or U442 (N_442,In_2447,In_1347);
and U443 (N_443,In_1440,In_1225);
and U444 (N_444,In_1964,In_24);
xor U445 (N_445,In_278,In_805);
nor U446 (N_446,In_17,In_1794);
xor U447 (N_447,In_945,In_2332);
or U448 (N_448,In_286,In_1610);
nand U449 (N_449,In_1319,In_703);
and U450 (N_450,In_188,In_809);
and U451 (N_451,In_658,In_1234);
xnor U452 (N_452,In_334,In_2206);
xor U453 (N_453,In_1076,In_2252);
nand U454 (N_454,In_1512,In_374);
and U455 (N_455,In_700,In_1690);
xnor U456 (N_456,In_939,In_1196);
nor U457 (N_457,In_2165,In_2075);
and U458 (N_458,In_1714,In_1354);
xor U459 (N_459,In_1705,In_1812);
or U460 (N_460,In_1146,In_448);
or U461 (N_461,In_80,In_1646);
xnor U462 (N_462,In_1467,In_1733);
xnor U463 (N_463,In_1169,In_91);
nor U464 (N_464,In_1892,In_1545);
or U465 (N_465,In_1910,In_546);
or U466 (N_466,In_148,In_578);
nor U467 (N_467,In_1469,In_287);
nor U468 (N_468,In_1394,In_1219);
xor U469 (N_469,In_1664,In_669);
or U470 (N_470,In_452,In_2096);
nand U471 (N_471,In_765,In_1873);
or U472 (N_472,In_1658,In_475);
or U473 (N_473,In_342,In_141);
or U474 (N_474,In_2421,In_2244);
xor U475 (N_475,In_39,In_208);
nand U476 (N_476,In_863,In_1115);
and U477 (N_477,In_92,In_1022);
or U478 (N_478,In_356,In_1821);
nand U479 (N_479,In_4,In_621);
nor U480 (N_480,In_597,In_1539);
and U481 (N_481,In_1290,In_110);
xnor U482 (N_482,In_957,In_800);
and U483 (N_483,In_787,In_57);
and U484 (N_484,In_1119,In_690);
and U485 (N_485,In_1496,In_1670);
or U486 (N_486,In_2143,In_1471);
nor U487 (N_487,In_1601,In_2425);
xnor U488 (N_488,In_684,In_1402);
xnor U489 (N_489,In_1905,In_1619);
nor U490 (N_490,In_19,In_1302);
and U491 (N_491,In_2371,In_1228);
or U492 (N_492,In_2275,In_2465);
nand U493 (N_493,In_1158,In_496);
or U494 (N_494,In_1600,In_1163);
or U495 (N_495,In_1935,In_63);
nand U496 (N_496,In_1819,In_1851);
or U497 (N_497,In_367,In_776);
xor U498 (N_498,In_2232,In_2010);
and U499 (N_499,In_2027,In_214);
and U500 (N_500,In_1333,In_746);
xor U501 (N_501,In_1981,In_2338);
nand U502 (N_502,In_1220,In_255);
nor U503 (N_503,In_1230,In_1640);
and U504 (N_504,In_2312,In_180);
nand U505 (N_505,In_1090,In_971);
or U506 (N_506,In_383,In_2090);
nand U507 (N_507,In_1445,In_1417);
nand U508 (N_508,In_2348,In_1156);
nand U509 (N_509,In_779,In_2063);
nand U510 (N_510,In_1925,In_2141);
or U511 (N_511,In_2426,In_710);
xor U512 (N_512,In_279,In_1616);
and U513 (N_513,In_2081,In_1381);
and U514 (N_514,In_238,In_64);
nor U515 (N_515,In_2024,In_97);
nor U516 (N_516,In_1203,In_2441);
xnor U517 (N_517,In_2419,In_539);
nand U518 (N_518,In_848,In_727);
and U519 (N_519,In_2285,In_2301);
nand U520 (N_520,In_162,In_1424);
nor U521 (N_521,In_2036,In_1630);
nand U522 (N_522,In_875,In_311);
and U523 (N_523,In_2140,In_1167);
nand U524 (N_524,In_2035,In_401);
xnor U525 (N_525,In_1859,In_617);
and U526 (N_526,In_2459,In_2458);
xnor U527 (N_527,In_1239,In_1032);
nor U528 (N_528,In_1791,In_1025);
and U529 (N_529,In_1345,In_2282);
or U530 (N_530,In_717,In_2271);
xnor U531 (N_531,In_1522,In_218);
and U532 (N_532,In_1086,In_2246);
nand U533 (N_533,In_220,In_1036);
or U534 (N_534,In_682,In_268);
or U535 (N_535,In_601,In_1824);
nand U536 (N_536,In_1916,In_2176);
or U537 (N_537,In_627,In_790);
and U538 (N_538,In_2228,In_361);
nand U539 (N_539,In_246,In_1624);
nor U540 (N_540,In_502,In_909);
xor U541 (N_541,In_1904,In_2488);
or U542 (N_542,In_85,In_602);
nor U543 (N_543,In_782,In_1491);
or U544 (N_544,In_676,In_61);
nand U545 (N_545,In_51,In_2391);
xnor U546 (N_546,In_1803,In_2008);
or U547 (N_547,In_1869,In_1693);
or U548 (N_548,In_200,In_1576);
xor U549 (N_549,In_926,In_1710);
or U550 (N_550,In_1837,In_2071);
or U551 (N_551,In_1444,In_163);
nand U552 (N_552,In_2050,In_2204);
xnor U553 (N_553,In_2183,In_2494);
and U554 (N_554,In_899,In_1918);
nor U555 (N_555,In_445,In_2230);
xnor U556 (N_556,In_182,In_1464);
and U557 (N_557,In_1764,In_2082);
nor U558 (N_558,In_2162,In_1406);
nor U559 (N_559,In_2401,In_1770);
nor U560 (N_560,In_1955,In_1063);
nand U561 (N_561,In_1543,In_1756);
nand U562 (N_562,In_2436,In_1034);
or U563 (N_563,In_2329,In_99);
nand U564 (N_564,In_147,In_1972);
nand U565 (N_565,In_2083,In_202);
xor U566 (N_566,In_10,In_1081);
xor U567 (N_567,In_1079,In_1363);
xnor U568 (N_568,In_2305,In_1485);
xor U569 (N_569,In_1991,In_100);
and U570 (N_570,In_483,In_846);
or U571 (N_571,In_666,In_651);
and U572 (N_572,In_155,In_1236);
nand U573 (N_573,In_2467,In_1523);
or U574 (N_574,In_194,In_547);
nor U575 (N_575,In_209,In_1779);
or U576 (N_576,In_832,In_435);
xor U577 (N_577,In_867,In_981);
xor U578 (N_578,In_1244,In_2442);
nand U579 (N_579,In_2261,In_1528);
nor U580 (N_580,In_2450,In_934);
nand U581 (N_581,In_888,In_77);
nor U582 (N_582,In_288,In_789);
and U583 (N_583,In_90,In_551);
or U584 (N_584,In_1201,In_229);
nor U585 (N_585,In_1147,In_1250);
nand U586 (N_586,In_594,In_1461);
or U587 (N_587,In_959,In_1546);
or U588 (N_588,In_908,In_1123);
nand U589 (N_589,In_67,In_1901);
nor U590 (N_590,In_282,In_1622);
xnor U591 (N_591,In_2434,In_1296);
or U592 (N_592,In_44,In_1798);
nor U593 (N_593,In_1336,In_734);
nor U594 (N_594,In_49,In_933);
nor U595 (N_595,In_2091,In_455);
nor U596 (N_596,In_1077,In_86);
xnor U597 (N_597,In_1030,In_1795);
and U598 (N_598,In_891,In_1678);
xnor U599 (N_599,In_2344,In_1004);
and U600 (N_600,In_52,In_827);
nand U601 (N_601,In_1349,In_2387);
nor U602 (N_602,In_1716,In_456);
and U603 (N_603,In_1977,In_260);
nor U604 (N_604,In_1343,In_1570);
or U605 (N_605,In_432,In_2355);
xor U606 (N_606,In_807,In_1835);
or U607 (N_607,In_101,In_2242);
and U608 (N_608,In_173,In_709);
xnor U609 (N_609,In_2129,In_505);
and U610 (N_610,In_104,In_575);
and U611 (N_611,In_348,In_2432);
nor U612 (N_612,In_654,In_1356);
nand U613 (N_613,In_922,In_2235);
and U614 (N_614,In_3,In_1914);
and U615 (N_615,In_1558,In_1787);
or U616 (N_616,In_177,In_369);
and U617 (N_617,In_1662,In_211);
xnor U618 (N_618,In_607,In_1599);
xnor U619 (N_619,In_2476,In_1878);
nand U620 (N_620,In_1882,In_399);
xor U621 (N_621,In_1744,In_1130);
or U622 (N_622,In_1131,In_866);
or U623 (N_623,In_2349,In_2029);
and U624 (N_624,In_1897,In_167);
or U625 (N_625,In_429,In_1992);
nand U626 (N_626,In_1766,In_973);
nand U627 (N_627,In_1017,In_898);
and U628 (N_628,In_1329,In_841);
and U629 (N_629,In_1427,In_2451);
nand U630 (N_630,In_2188,In_679);
or U631 (N_631,In_1909,In_414);
nor U632 (N_632,In_2067,In_1694);
nor U633 (N_633,In_347,In_1348);
and U634 (N_634,In_412,In_2443);
nand U635 (N_635,In_2317,In_2257);
nand U636 (N_636,In_106,In_1745);
xnor U637 (N_637,In_798,In_2186);
or U638 (N_638,In_335,In_1934);
and U639 (N_639,In_1252,In_1311);
xnor U640 (N_640,In_541,In_1508);
and U641 (N_641,In_2361,In_1010);
nand U642 (N_642,In_504,In_1320);
xnor U643 (N_643,In_2134,In_2279);
nor U644 (N_644,In_1162,In_1246);
or U645 (N_645,In_2098,In_917);
and U646 (N_646,In_2269,In_1706);
xor U647 (N_647,In_1604,In_754);
xor U648 (N_648,In_1229,In_364);
xnor U649 (N_649,In_1454,In_1582);
and U650 (N_650,In_2218,In_1765);
or U651 (N_651,In_797,In_931);
nand U652 (N_652,In_536,In_346);
or U653 (N_653,In_2026,In_777);
xor U654 (N_654,In_2260,In_1046);
xnor U655 (N_655,In_1105,In_1936);
nand U656 (N_656,In_2086,In_759);
xor U657 (N_657,In_1182,In_1442);
or U658 (N_658,In_2417,In_882);
xnor U659 (N_659,In_1253,In_1611);
xor U660 (N_660,In_1151,In_1154);
xor U661 (N_661,In_1309,In_936);
xnor U662 (N_662,In_478,In_277);
and U663 (N_663,In_352,In_749);
nand U664 (N_664,In_1732,In_1726);
or U665 (N_665,In_1559,In_1503);
xnor U666 (N_666,In_1937,In_1684);
and U667 (N_667,In_2249,In_979);
or U668 (N_668,In_212,In_2278);
nand U669 (N_669,In_1476,In_89);
nand U670 (N_670,In_1185,In_1506);
nor U671 (N_671,In_836,In_2139);
and U672 (N_672,In_1270,In_928);
nor U673 (N_673,In_1255,In_1499);
nand U674 (N_674,In_835,In_480);
or U675 (N_675,In_2127,In_1644);
or U676 (N_676,In_1026,In_1190);
xor U677 (N_677,In_733,In_296);
and U678 (N_678,In_1863,In_1308);
xor U679 (N_679,In_542,In_1038);
xor U680 (N_680,In_1625,In_2490);
nor U681 (N_681,In_974,In_1514);
nor U682 (N_682,In_136,In_1548);
nand U683 (N_683,In_1505,In_2175);
xor U684 (N_684,In_2357,In_2065);
nor U685 (N_685,In_976,In_785);
nor U686 (N_686,In_1549,In_698);
and U687 (N_687,In_65,In_109);
or U688 (N_688,In_126,In_1160);
nor U689 (N_689,In_2229,In_687);
and U690 (N_690,In_2324,In_986);
nand U691 (N_691,In_509,In_312);
nand U692 (N_692,In_204,In_1288);
and U693 (N_693,In_1535,In_2064);
nor U694 (N_694,In_831,In_1922);
nor U695 (N_695,In_760,In_304);
or U696 (N_696,In_2216,In_1477);
nand U697 (N_697,In_468,In_2073);
nand U698 (N_698,In_1951,In_2368);
and U699 (N_699,In_665,In_2080);
xor U700 (N_700,In_1330,In_1944);
xnor U701 (N_701,In_968,In_130);
xnor U702 (N_702,In_2054,In_303);
or U703 (N_703,In_2150,In_1120);
and U704 (N_704,In_1890,In_1521);
and U705 (N_705,In_175,In_822);
xnor U706 (N_706,In_18,In_1060);
xnor U707 (N_707,In_492,In_336);
nor U708 (N_708,In_1986,In_1074);
xnor U709 (N_709,In_2236,In_2053);
nand U710 (N_710,In_2411,In_1698);
nor U711 (N_711,In_1969,In_701);
nor U712 (N_712,In_1865,In_454);
xor U713 (N_713,In_169,In_1602);
nand U714 (N_714,In_358,In_880);
and U715 (N_715,In_2359,In_940);
xor U716 (N_716,In_1263,In_1195);
xor U717 (N_717,In_1713,In_121);
or U718 (N_718,In_262,In_996);
xnor U719 (N_719,In_2128,In_1109);
xor U720 (N_720,In_1457,In_30);
nand U721 (N_721,In_932,In_1850);
nor U722 (N_722,In_2037,In_1760);
and U723 (N_723,In_76,In_927);
nor U724 (N_724,In_1946,In_81);
nor U725 (N_725,In_1317,In_2167);
or U726 (N_726,In_186,In_2482);
and U727 (N_727,In_738,In_720);
or U728 (N_728,In_1757,In_2462);
or U729 (N_729,In_960,In_354);
or U730 (N_730,In_642,In_556);
nor U731 (N_731,In_1114,In_1300);
xnor U732 (N_732,In_460,In_2393);
and U733 (N_733,In_2070,In_2322);
nand U734 (N_734,In_2164,In_1065);
and U735 (N_735,In_477,In_481);
or U736 (N_736,In_780,In_1541);
and U737 (N_737,In_306,In_763);
nor U738 (N_738,In_2205,In_1752);
xnor U739 (N_739,In_36,In_554);
or U740 (N_740,In_1118,In_2363);
and U741 (N_741,In_1351,In_124);
xor U742 (N_742,In_1741,In_1126);
or U743 (N_743,In_1155,In_2299);
or U744 (N_744,In_88,In_856);
or U745 (N_745,In_2203,In_1717);
nand U746 (N_746,In_1725,In_263);
nor U747 (N_747,In_307,In_2094);
and U748 (N_748,In_1374,In_862);
or U749 (N_749,In_591,In_1940);
or U750 (N_750,In_389,In_961);
or U751 (N_751,In_796,In_965);
or U752 (N_752,In_269,In_2339);
xor U753 (N_753,In_510,In_2120);
and U754 (N_754,In_503,In_2280);
or U755 (N_755,In_802,In_1066);
xor U756 (N_756,In_1564,In_1399);
nor U757 (N_757,In_1012,In_667);
nor U758 (N_758,In_1785,In_1240);
or U759 (N_759,In_1927,In_1312);
and U760 (N_760,In_98,In_386);
nand U761 (N_761,In_1051,In_297);
nand U762 (N_762,In_2185,In_127);
and U763 (N_763,In_2160,In_634);
nand U764 (N_764,In_833,In_756);
and U765 (N_765,In_2011,In_33);
and U766 (N_766,In_1715,In_792);
xnor U767 (N_767,In_1247,In_724);
nand U768 (N_768,In_1899,In_1958);
xnor U769 (N_769,In_2294,In_1422);
or U770 (N_770,In_1649,In_2093);
nand U771 (N_771,In_1566,In_372);
or U772 (N_772,In_133,In_1872);
or U773 (N_773,In_2133,In_1306);
nand U774 (N_774,In_2058,In_484);
xor U775 (N_775,In_1654,In_569);
xnor U776 (N_776,In_402,In_2137);
xnor U777 (N_777,In_1023,In_473);
or U778 (N_778,In_988,In_171);
nor U779 (N_779,In_884,In_292);
nor U780 (N_780,In_1104,In_1519);
xor U781 (N_781,In_2497,In_535);
nand U782 (N_782,In_1008,In_411);
nor U783 (N_783,In_1502,In_529);
nand U784 (N_784,In_1743,In_1651);
nor U785 (N_785,In_1259,In_989);
nor U786 (N_786,In_638,In_406);
or U787 (N_787,In_925,In_1687);
or U788 (N_788,In_561,In_2403);
xor U789 (N_789,In_1886,In_2052);
nand U790 (N_790,In_1982,In_2330);
or U791 (N_791,In_1205,In_1961);
and U792 (N_792,In_1455,In_2234);
nor U793 (N_793,In_620,In_1802);
xor U794 (N_794,In_1857,In_139);
nor U795 (N_795,In_688,In_1854);
xor U796 (N_796,In_2031,In_2410);
and U797 (N_797,In_340,In_1583);
nor U798 (N_798,In_1138,In_1565);
and U799 (N_799,In_1567,In_2149);
nand U800 (N_800,In_2189,In_1660);
xor U801 (N_801,In_1224,In_430);
and U802 (N_802,In_1213,In_742);
nor U803 (N_803,In_938,In_1189);
and U804 (N_804,In_707,In_2191);
nor U805 (N_805,In_1021,In_1990);
and U806 (N_806,In_320,In_403);
nor U807 (N_807,In_2184,In_1033);
xnor U808 (N_808,In_530,In_537);
xor U809 (N_809,In_1551,In_766);
and U810 (N_810,In_964,In_2264);
nor U811 (N_811,In_416,In_332);
or U812 (N_812,In_1245,In_40);
nand U813 (N_813,In_1355,In_2373);
xnor U814 (N_814,In_2323,In_1407);
xnor U815 (N_815,In_1050,In_1739);
nand U816 (N_816,In_2163,In_1831);
xor U817 (N_817,In_2309,In_714);
nand U818 (N_818,In_384,In_953);
xnor U819 (N_819,In_512,In_1194);
and U820 (N_820,In_54,In_317);
nand U821 (N_821,In_2351,In_1817);
and U822 (N_822,In_1712,In_1973);
nand U823 (N_823,In_923,In_195);
xnor U824 (N_824,In_2100,In_1327);
nand U825 (N_825,In_2161,In_1761);
xor U826 (N_826,In_1588,In_300);
xnor U827 (N_827,In_519,In_2241);
nand U828 (N_828,In_439,In_264);
nand U829 (N_829,In_93,In_2295);
xor U830 (N_830,In_442,In_886);
nor U831 (N_831,In_1661,In_443);
nor U832 (N_832,In_1699,In_739);
nand U833 (N_833,In_747,In_673);
or U834 (N_834,In_251,In_1301);
nand U835 (N_835,In_453,In_1985);
nand U836 (N_836,In_152,In_2284);
xnor U837 (N_837,In_1993,In_1771);
and U838 (N_838,In_1667,In_857);
and U839 (N_839,In_775,In_1080);
xor U840 (N_840,In_228,In_748);
or U841 (N_841,In_318,In_544);
or U842 (N_842,In_145,In_466);
or U843 (N_843,In_373,In_639);
nand U844 (N_844,In_1384,In_2473);
nand U845 (N_845,In_2326,In_397);
xor U846 (N_846,In_527,In_1434);
xnor U847 (N_847,In_1178,In_2148);
nor U848 (N_848,In_1382,In_450);
nand U849 (N_849,In_1430,In_2124);
xor U850 (N_850,In_1136,In_1083);
or U851 (N_851,In_2382,In_1111);
and U852 (N_852,In_74,In_731);
and U853 (N_853,In_773,In_1862);
xor U854 (N_854,In_2397,In_740);
nand U855 (N_855,In_2130,In_1846);
xnor U856 (N_856,In_434,In_1647);
xnor U857 (N_857,In_1680,In_15);
nor U858 (N_858,In_375,In_2336);
nand U859 (N_859,In_1209,In_671);
xnor U860 (N_860,In_689,In_234);
nand U861 (N_861,In_236,In_1801);
or U862 (N_862,In_2321,In_2350);
xnor U863 (N_863,In_84,In_613);
nor U864 (N_864,In_2151,In_2366);
or U865 (N_865,In_1000,In_1518);
or U866 (N_866,In_1504,In_1470);
xnor U867 (N_867,In_1593,In_564);
or U868 (N_868,In_854,In_1618);
xnor U869 (N_869,In_199,In_2113);
nand U870 (N_870,In_222,In_767);
nand U871 (N_871,In_735,In_1084);
or U872 (N_872,In_1731,In_1124);
or U873 (N_873,In_506,In_1125);
and U874 (N_874,In_2328,In_580);
nand U875 (N_875,In_1179,In_1811);
xnor U876 (N_876,In_107,In_1278);
xor U877 (N_877,In_1013,In_2365);
and U878 (N_878,In_408,In_2238);
and U879 (N_879,In_1634,In_2297);
or U880 (N_880,In_2142,In_1400);
nand U881 (N_881,In_1891,In_1527);
nor U882 (N_882,In_1932,In_1223);
and U883 (N_883,In_2179,In_999);
xor U884 (N_884,In_2345,In_2420);
and U885 (N_885,In_941,In_1226);
nor U886 (N_886,In_2079,In_2095);
nor U887 (N_887,In_1838,In_952);
nand U888 (N_888,In_921,In_808);
and U889 (N_889,In_2038,In_1387);
nor U890 (N_890,In_1277,In_1842);
nand U891 (N_891,In_1919,In_441);
and U892 (N_892,In_712,In_1353);
and U893 (N_893,In_197,In_577);
xor U894 (N_894,In_1049,In_71);
and U895 (N_895,In_2331,In_781);
nand U896 (N_896,In_2157,In_2388);
nand U897 (N_897,In_2062,In_1758);
nor U898 (N_898,In_1268,In_589);
nor U899 (N_899,In_2380,In_770);
xor U900 (N_900,In_2454,In_193);
nor U901 (N_901,In_1332,In_579);
nor U902 (N_902,In_1620,In_1075);
nand U903 (N_903,In_845,In_1809);
nand U904 (N_904,In_1177,In_1573);
or U905 (N_905,In_723,In_904);
or U906 (N_906,In_2385,In_2039);
nor U907 (N_907,In_697,In_1014);
nor U908 (N_908,In_95,In_1587);
nor U909 (N_909,In_2272,In_378);
and U910 (N_910,In_1704,In_1243);
nor U911 (N_911,In_558,In_869);
and U912 (N_912,In_691,In_2112);
nor U913 (N_913,In_285,In_405);
or U914 (N_914,In_2061,In_699);
or U915 (N_915,In_463,In_1975);
and U916 (N_916,In_1204,In_2310);
and U917 (N_917,In_1433,In_582);
nand U918 (N_918,In_2212,In_1868);
nand U919 (N_919,In_1557,In_984);
xnor U920 (N_920,In_1928,In_1438);
or U921 (N_921,In_1380,In_2044);
and U922 (N_922,In_659,In_319);
nor U923 (N_923,In_522,In_1463);
and U924 (N_924,In_471,In_302);
and U925 (N_925,In_2069,In_13);
or U926 (N_926,In_520,In_1960);
or U927 (N_927,In_1404,In_2466);
nor U928 (N_928,In_584,In_2448);
xor U929 (N_929,In_563,In_1414);
nand U930 (N_930,In_1639,In_1346);
nor U931 (N_931,In_823,In_32);
nand U932 (N_932,In_1829,In_2227);
nand U933 (N_933,In_1293,In_142);
or U934 (N_934,In_2145,In_105);
xor U935 (N_935,In_943,In_1844);
nor U936 (N_936,In_183,In_2107);
nor U937 (N_937,In_1016,In_1581);
nor U938 (N_938,In_2047,In_566);
or U939 (N_939,In_1645,In_1235);
xor U940 (N_940,In_363,In_2258);
nor U941 (N_941,In_540,In_2341);
xor U942 (N_942,In_1361,In_804);
nand U943 (N_943,In_159,In_240);
xor U944 (N_944,In_1833,In_694);
or U945 (N_945,In_1880,In_257);
nor U946 (N_946,In_2101,In_721);
nand U947 (N_947,In_1420,In_137);
or U948 (N_948,In_1047,In_2034);
or U949 (N_949,In_1983,In_641);
xnor U950 (N_950,In_331,In_1458);
and U951 (N_951,In_664,In_1342);
xnor U952 (N_952,In_50,In_1062);
and U953 (N_953,In_178,In_1832);
or U954 (N_954,In_12,In_1571);
or U955 (N_955,In_215,In_328);
nor U956 (N_956,In_2182,In_1087);
and U957 (N_957,In_870,In_2089);
or U958 (N_958,In_750,In_1814);
xnor U959 (N_959,In_1428,In_1251);
and U960 (N_960,In_1456,In_980);
nand U961 (N_961,In_2276,In_534);
nand U962 (N_962,In_2296,In_2337);
and U963 (N_963,In_345,In_339);
xor U964 (N_964,In_1078,In_1041);
or U965 (N_965,In_1633,In_27);
and U966 (N_966,In_771,In_685);
nor U967 (N_967,In_604,In_1995);
or U968 (N_968,In_253,In_1805);
nor U969 (N_969,In_447,In_606);
nor U970 (N_970,In_192,In_929);
nand U971 (N_971,In_660,In_2374);
and U972 (N_972,In_1267,In_1403);
nand U973 (N_973,In_1048,In_2270);
and U974 (N_974,In_2051,In_1112);
or U975 (N_975,In_1997,In_858);
xnor U976 (N_976,In_341,In_876);
xnor U977 (N_977,In_557,In_2395);
xor U978 (N_978,In_1447,In_1274);
nor U979 (N_979,In_830,In_508);
xnor U980 (N_980,In_70,In_652);
and U981 (N_981,In_1412,In_1297);
or U982 (N_982,In_1648,In_1762);
xor U983 (N_983,In_131,In_585);
nor U984 (N_984,In_1419,In_764);
xnor U985 (N_985,In_350,In_1389);
nor U986 (N_986,In_1218,In_1318);
nor U987 (N_987,In_2464,In_2231);
xnor U988 (N_988,In_514,In_1494);
or U989 (N_989,In_715,In_1462);
and U990 (N_990,In_216,In_992);
or U991 (N_991,In_1531,In_1544);
nor U992 (N_992,In_315,In_2383);
nand U993 (N_993,In_1830,In_677);
nor U994 (N_994,In_649,In_1028);
nor U995 (N_995,In_440,In_788);
and U996 (N_996,In_1379,In_79);
nand U997 (N_997,In_1472,In_711);
and U998 (N_998,In_1652,In_2311);
xor U999 (N_999,In_1122,In_1852);
xnor U1000 (N_1000,In_1148,In_1979);
xor U1001 (N_1001,In_243,In_273);
xor U1002 (N_1002,In_2308,In_1776);
nand U1003 (N_1003,In_1885,In_1366);
xnor U1004 (N_1004,In_795,In_1793);
xor U1005 (N_1005,In_293,In_2197);
nor U1006 (N_1006,In_1053,In_2215);
nor U1007 (N_1007,In_2125,In_125);
nand U1008 (N_1008,In_164,In_622);
and U1009 (N_1009,In_1292,In_816);
nor U1010 (N_1010,In_2221,In_1672);
xor U1011 (N_1011,In_2377,In_150);
or U1012 (N_1012,In_2416,In_1682);
xnor U1013 (N_1013,In_791,In_1586);
nand U1014 (N_1014,In_66,In_476);
or U1015 (N_1015,In_451,In_1774);
and U1016 (N_1016,In_1315,In_2290);
nand U1017 (N_1017,In_1954,In_2092);
nand U1018 (N_1018,In_686,In_1121);
and U1019 (N_1019,In_2144,In_1287);
or U1020 (N_1020,In_421,In_2318);
and U1021 (N_1021,In_427,In_877);
nor U1022 (N_1022,In_1237,In_225);
or U1023 (N_1023,In_718,In_1465);
or U1024 (N_1024,In_1818,In_644);
xnor U1025 (N_1025,In_1258,In_1103);
nand U1026 (N_1026,In_1635,In_865);
and U1027 (N_1027,In_834,In_1272);
or U1028 (N_1028,In_404,In_174);
or U1029 (N_1029,In_313,In_413);
or U1030 (N_1030,In_762,In_568);
or U1031 (N_1031,In_2115,In_2200);
xnor U1032 (N_1032,In_490,In_467);
nor U1033 (N_1033,In_513,In_1085);
xnor U1034 (N_1034,In_725,In_1675);
nand U1035 (N_1035,In_645,In_1810);
or U1036 (N_1036,In_494,In_1775);
and U1037 (N_1037,In_62,In_221);
xor U1038 (N_1038,In_2400,In_1241);
or U1039 (N_1039,In_2154,In_1782);
xor U1040 (N_1040,In_1574,In_1552);
xnor U1041 (N_1041,In_626,In_249);
nand U1042 (N_1042,In_1864,In_129);
nor U1043 (N_1043,In_244,In_1516);
or U1044 (N_1044,In_1598,In_1627);
and U1045 (N_1045,In_1578,In_128);
nand U1046 (N_1046,In_2406,In_1276);
or U1047 (N_1047,In_950,In_1695);
and U1048 (N_1048,In_2178,In_511);
nor U1049 (N_1049,In_729,In_761);
nand U1050 (N_1050,In_736,In_232);
or U1051 (N_1051,In_2021,In_2224);
nand U1052 (N_1052,In_258,In_2159);
nand U1053 (N_1053,In_1221,In_794);
nand U1054 (N_1054,In_2245,In_1322);
or U1055 (N_1055,In_1397,In_2319);
and U1056 (N_1056,In_1510,In_559);
nor U1057 (N_1057,In_2198,In_1294);
nand U1058 (N_1058,In_951,In_2480);
xor U1059 (N_1059,In_683,In_2049);
xnor U1060 (N_1060,In_2430,In_2255);
xor U1061 (N_1061,In_825,In_1562);
nor U1062 (N_1062,In_2002,In_636);
nor U1063 (N_1063,In_2453,In_295);
nand U1064 (N_1064,In_1018,In_1853);
and U1065 (N_1065,In_978,In_261);
nor U1066 (N_1066,In_2147,In_674);
nand U1067 (N_1067,In_1291,In_1386);
and U1068 (N_1068,In_1554,In_2102);
nand U1069 (N_1069,In_380,In_1117);
nand U1070 (N_1070,In_2499,In_786);
xnor U1071 (N_1071,In_1839,In_1911);
xor U1072 (N_1072,In_1696,In_1747);
or U1073 (N_1073,In_1364,In_333);
xnor U1074 (N_1074,In_1093,In_1057);
nand U1075 (N_1075,In_283,In_890);
nor U1076 (N_1076,In_1845,In_678);
or U1077 (N_1077,In_2017,In_485);
xor U1078 (N_1078,In_1375,In_1215);
nor U1079 (N_1079,In_1216,In_1040);
and U1080 (N_1080,In_2001,In_2219);
and U1081 (N_1081,In_60,In_1730);
nor U1082 (N_1082,In_1413,In_1);
nand U1083 (N_1083,In_1262,In_1193);
xor U1084 (N_1084,In_618,In_280);
and U1085 (N_1085,In_377,In_1045);
nor U1086 (N_1086,In_394,In_646);
and U1087 (N_1087,In_252,In_1289);
xor U1088 (N_1088,In_26,In_366);
and U1089 (N_1089,In_1421,In_635);
xor U1090 (N_1090,In_1679,In_1778);
nand U1091 (N_1091,In_2209,In_656);
xor U1092 (N_1092,In_538,In_1344);
nand U1093 (N_1093,In_2392,In_716);
xor U1094 (N_1094,In_497,In_948);
and U1095 (N_1095,In_245,In_2431);
or U1096 (N_1096,In_611,In_34);
nand U1097 (N_1097,In_1307,In_1636);
nand U1098 (N_1098,In_242,In_977);
or U1099 (N_1099,In_1283,In_1227);
nand U1100 (N_1100,In_1749,In_1926);
nand U1101 (N_1101,In_1475,In_2478);
and U1102 (N_1102,In_294,In_2014);
nand U1103 (N_1103,In_2254,In_449);
nor U1104 (N_1104,In_516,In_1930);
xnor U1105 (N_1105,In_281,In_407);
nand U1106 (N_1106,In_555,In_893);
nor U1107 (N_1107,In_1568,In_111);
or U1108 (N_1108,In_1153,In_437);
or U1109 (N_1109,In_1700,In_1822);
xor U1110 (N_1110,In_2288,In_814);
nand U1111 (N_1111,In_521,In_2384);
nand U1112 (N_1112,In_1792,In_2202);
or U1113 (N_1113,In_1942,In_1631);
and U1114 (N_1114,In_524,In_2043);
nand U1115 (N_1115,In_2084,In_1642);
or U1116 (N_1116,In_2023,In_811);
xnor U1117 (N_1117,In_2479,In_1001);
or U1118 (N_1118,In_1719,In_942);
nor U1119 (N_1119,In_2169,In_1569);
xnor U1120 (N_1120,In_1638,In_2087);
nand U1121 (N_1121,In_1788,In_1615);
nor U1122 (N_1122,In_2181,In_123);
xor U1123 (N_1123,In_2484,In_2287);
xor U1124 (N_1124,In_1888,In_140);
and U1125 (N_1125,In_1335,In_821);
nor U1126 (N_1126,In_532,In_103);
and U1127 (N_1127,In_1828,In_1488);
and U1128 (N_1128,In_2020,In_1376);
and U1129 (N_1129,In_423,In_2364);
nor U1130 (N_1130,In_2491,In_259);
or U1131 (N_1131,In_11,In_1401);
xnor U1132 (N_1132,In_2445,In_1408);
and U1133 (N_1133,In_2118,In_1197);
xor U1134 (N_1134,In_549,In_2222);
xor U1135 (N_1135,In_444,In_758);
nor U1136 (N_1136,In_562,In_1281);
or U1137 (N_1137,In_2173,In_38);
and U1138 (N_1138,In_1493,In_2171);
xnor U1139 (N_1139,In_1340,In_1703);
or U1140 (N_1140,In_753,In_385);
xor U1141 (N_1141,In_947,In_309);
xor U1142 (N_1142,In_400,In_810);
nand U1143 (N_1143,In_1423,In_1359);
xnor U1144 (N_1144,In_1487,In_1707);
nor U1145 (N_1145,In_2104,In_2213);
nand U1146 (N_1146,In_2040,In_1740);
nor U1147 (N_1147,In_1721,In_1478);
or U1148 (N_1148,In_2012,In_1097);
nand U1149 (N_1149,In_570,In_1655);
nor U1150 (N_1150,In_1007,In_2136);
nand U1151 (N_1151,In_1142,In_1377);
xor U1152 (N_1152,In_1334,In_96);
xor U1153 (N_1153,In_189,In_1395);
and U1154 (N_1154,In_695,In_704);
nand U1155 (N_1155,In_1637,In_1799);
or U1156 (N_1156,In_1044,In_1357);
and U1157 (N_1157,In_2405,In_1088);
nor U1158 (N_1158,In_181,In_1145);
nand U1159 (N_1159,In_1952,In_2433);
xnor U1160 (N_1160,In_706,In_2302);
nor U1161 (N_1161,In_2030,In_87);
or U1162 (N_1162,In_2004,In_1208);
or U1163 (N_1163,In_1603,In_436);
nand U1164 (N_1164,In_1676,In_982);
or U1165 (N_1165,In_985,In_176);
and U1166 (N_1166,In_1867,In_2300);
and U1167 (N_1167,In_744,In_892);
xor U1168 (N_1168,In_1968,In_2438);
or U1169 (N_1169,In_1107,In_117);
nor U1170 (N_1170,In_545,In_1092);
or U1171 (N_1171,In_2122,In_1957);
xor U1172 (N_1172,In_1411,In_1517);
nor U1173 (N_1173,In_325,In_349);
nor U1174 (N_1174,In_1608,In_2277);
nand U1175 (N_1175,In_381,In_647);
nand U1176 (N_1176,In_1113,In_783);
nand U1177 (N_1177,In_132,In_1781);
xnor U1178 (N_1178,In_2452,In_1515);
nand U1179 (N_1179,In_1367,In_187);
nor U1180 (N_1180,In_1896,In_1392);
and U1181 (N_1181,In_35,In_1285);
xor U1182 (N_1182,In_474,In_2313);
nand U1183 (N_1183,In_2315,In_2286);
nand U1184 (N_1184,In_488,In_314);
nor U1185 (N_1185,In_1054,In_1181);
and U1186 (N_1186,In_1172,In_2437);
xnor U1187 (N_1187,In_2060,In_1800);
and U1188 (N_1188,In_1388,In_2046);
nor U1189 (N_1189,In_2263,In_528);
nand U1190 (N_1190,In_2103,In_2132);
nand U1191 (N_1191,In_1286,In_119);
xnor U1192 (N_1192,In_2469,In_172);
nor U1193 (N_1193,In_469,In_680);
nand U1194 (N_1194,In_517,In_379);
and U1195 (N_1195,In_631,In_1848);
and U1196 (N_1196,In_905,In_2353);
nand U1197 (N_1197,In_850,In_1202);
or U1198 (N_1198,In_9,In_901);
and U1199 (N_1199,In_491,In_2402);
nor U1200 (N_1200,In_395,In_2381);
or U1201 (N_1201,In_1269,In_1024);
xnor U1202 (N_1202,In_1164,In_2367);
nor U1203 (N_1203,In_417,In_793);
or U1204 (N_1204,In_6,In_603);
and U1205 (N_1205,In_963,In_2376);
xor U1206 (N_1206,In_2356,In_1200);
xnor U1207 (N_1207,In_2394,In_650);
and U1208 (N_1208,In_1534,In_2372);
and U1209 (N_1209,In_1847,In_2074);
or U1210 (N_1210,In_1233,In_853);
xor U1211 (N_1211,In_1606,In_1722);
and U1212 (N_1212,In_2446,In_1561);
xnor U1213 (N_1213,In_1150,In_2369);
or U1214 (N_1214,In_730,In_1409);
nor U1215 (N_1215,In_1727,In_1323);
and U1216 (N_1216,In_573,In_461);
nand U1217 (N_1217,In_53,In_588);
nor U1218 (N_1218,In_1965,In_818);
xor U1219 (N_1219,In_583,In_276);
and U1220 (N_1220,In_1498,In_1187);
or U1221 (N_1221,In_1530,In_2250);
xor U1222 (N_1222,In_25,In_1841);
or U1223 (N_1223,In_2461,In_1173);
nor U1224 (N_1224,In_2111,In_1759);
and U1225 (N_1225,In_596,In_1191);
nand U1226 (N_1226,In_970,In_190);
nor U1227 (N_1227,In_207,In_2233);
xor U1228 (N_1228,In_1135,In_1613);
and U1229 (N_1229,In_2412,In_663);
nor U1230 (N_1230,In_1532,In_500);
and U1231 (N_1231,In_2135,In_326);
or U1232 (N_1232,In_587,In_895);
nor U1233 (N_1233,In_1500,In_1176);
xnor U1234 (N_1234,In_1073,In_2307);
or U1235 (N_1235,In_896,In_2057);
xnor U1236 (N_1236,In_1398,In_1962);
and U1237 (N_1237,In_628,In_2106);
nor U1238 (N_1238,In_2475,In_1217);
nor U1239 (N_1239,In_1628,In_464);
xnor U1240 (N_1240,In_966,In_387);
and U1241 (N_1241,In_2413,In_624);
and U1242 (N_1242,In_998,In_2006);
nor U1243 (N_1243,In_1697,In_1742);
or U1244 (N_1244,In_1484,In_1656);
or U1245 (N_1245,In_828,In_576);
nor U1246 (N_1246,In_198,In_1876);
and U1247 (N_1247,In_1171,In_274);
and U1248 (N_1248,In_135,In_1683);
and U1249 (N_1249,In_2470,In_1780);
nand U1250 (N_1250,In_1328,In_202);
xor U1251 (N_1251,In_1305,In_1545);
xor U1252 (N_1252,In_943,In_158);
nor U1253 (N_1253,In_132,In_462);
nor U1254 (N_1254,In_1304,In_143);
or U1255 (N_1255,In_2408,In_312);
nor U1256 (N_1256,In_135,In_608);
or U1257 (N_1257,In_1441,In_57);
and U1258 (N_1258,In_746,In_2247);
xor U1259 (N_1259,In_166,In_1223);
nand U1260 (N_1260,In_623,In_428);
nand U1261 (N_1261,In_2383,In_951);
nor U1262 (N_1262,In_1474,In_1887);
xor U1263 (N_1263,In_1571,In_2343);
or U1264 (N_1264,In_946,In_1266);
xor U1265 (N_1265,In_723,In_1173);
xnor U1266 (N_1266,In_1859,In_1624);
and U1267 (N_1267,In_642,In_2018);
nor U1268 (N_1268,In_135,In_290);
or U1269 (N_1269,In_1847,In_2097);
nor U1270 (N_1270,In_2443,In_1508);
and U1271 (N_1271,In_940,In_584);
nand U1272 (N_1272,In_61,In_2375);
xnor U1273 (N_1273,In_1742,In_1466);
or U1274 (N_1274,In_1459,In_1420);
nand U1275 (N_1275,In_175,In_29);
nor U1276 (N_1276,In_1237,In_1692);
and U1277 (N_1277,In_2134,In_951);
and U1278 (N_1278,In_2188,In_1467);
nand U1279 (N_1279,In_1347,In_698);
or U1280 (N_1280,In_2376,In_2023);
or U1281 (N_1281,In_1708,In_1666);
nor U1282 (N_1282,In_1115,In_60);
or U1283 (N_1283,In_1897,In_1680);
xnor U1284 (N_1284,In_1726,In_2244);
or U1285 (N_1285,In_1449,In_1975);
xor U1286 (N_1286,In_1512,In_1994);
and U1287 (N_1287,In_75,In_323);
and U1288 (N_1288,In_1245,In_1986);
nand U1289 (N_1289,In_458,In_2075);
and U1290 (N_1290,In_1245,In_35);
nand U1291 (N_1291,In_1561,In_143);
nor U1292 (N_1292,In_486,In_539);
or U1293 (N_1293,In_2337,In_2288);
xnor U1294 (N_1294,In_656,In_2245);
or U1295 (N_1295,In_2166,In_154);
nand U1296 (N_1296,In_1818,In_1279);
and U1297 (N_1297,In_803,In_667);
and U1298 (N_1298,In_660,In_1647);
nor U1299 (N_1299,In_636,In_2266);
nor U1300 (N_1300,In_344,In_1665);
nand U1301 (N_1301,In_2240,In_1767);
or U1302 (N_1302,In_591,In_365);
nand U1303 (N_1303,In_901,In_21);
or U1304 (N_1304,In_2428,In_992);
nand U1305 (N_1305,In_1389,In_2266);
and U1306 (N_1306,In_275,In_2279);
nand U1307 (N_1307,In_2093,In_1029);
nand U1308 (N_1308,In_1764,In_1125);
nor U1309 (N_1309,In_20,In_1258);
nand U1310 (N_1310,In_31,In_694);
nor U1311 (N_1311,In_252,In_1172);
and U1312 (N_1312,In_1536,In_113);
or U1313 (N_1313,In_2012,In_1346);
nor U1314 (N_1314,In_1193,In_1298);
nor U1315 (N_1315,In_2166,In_1920);
xnor U1316 (N_1316,In_2381,In_1692);
xor U1317 (N_1317,In_1483,In_2160);
xor U1318 (N_1318,In_1758,In_693);
nor U1319 (N_1319,In_1866,In_354);
xnor U1320 (N_1320,In_1234,In_1719);
xnor U1321 (N_1321,In_2072,In_1859);
nor U1322 (N_1322,In_2153,In_1831);
nor U1323 (N_1323,In_1448,In_2382);
xnor U1324 (N_1324,In_948,In_1246);
xnor U1325 (N_1325,In_964,In_304);
or U1326 (N_1326,In_2019,In_1382);
xnor U1327 (N_1327,In_2423,In_662);
and U1328 (N_1328,In_2184,In_1409);
nand U1329 (N_1329,In_497,In_337);
or U1330 (N_1330,In_797,In_730);
xnor U1331 (N_1331,In_2418,In_330);
nand U1332 (N_1332,In_705,In_1288);
nand U1333 (N_1333,In_275,In_1277);
nand U1334 (N_1334,In_502,In_1354);
xor U1335 (N_1335,In_586,In_1951);
xor U1336 (N_1336,In_1279,In_2156);
xor U1337 (N_1337,In_1191,In_1004);
and U1338 (N_1338,In_2256,In_158);
nor U1339 (N_1339,In_24,In_1427);
nor U1340 (N_1340,In_1417,In_2445);
or U1341 (N_1341,In_1630,In_2351);
or U1342 (N_1342,In_1556,In_700);
xnor U1343 (N_1343,In_562,In_1163);
nor U1344 (N_1344,In_1777,In_2275);
or U1345 (N_1345,In_2487,In_2439);
nand U1346 (N_1346,In_622,In_1596);
nor U1347 (N_1347,In_2435,In_524);
nor U1348 (N_1348,In_738,In_596);
and U1349 (N_1349,In_440,In_2369);
nor U1350 (N_1350,In_84,In_1141);
nor U1351 (N_1351,In_1537,In_88);
or U1352 (N_1352,In_1189,In_234);
or U1353 (N_1353,In_1886,In_540);
nor U1354 (N_1354,In_1807,In_164);
nor U1355 (N_1355,In_1544,In_1312);
or U1356 (N_1356,In_580,In_1891);
or U1357 (N_1357,In_2164,In_1050);
and U1358 (N_1358,In_2323,In_825);
or U1359 (N_1359,In_210,In_340);
and U1360 (N_1360,In_914,In_801);
nor U1361 (N_1361,In_1544,In_1168);
or U1362 (N_1362,In_1238,In_144);
xor U1363 (N_1363,In_2336,In_1740);
and U1364 (N_1364,In_1339,In_558);
and U1365 (N_1365,In_945,In_1198);
xor U1366 (N_1366,In_319,In_203);
nand U1367 (N_1367,In_1450,In_1133);
and U1368 (N_1368,In_15,In_1363);
nor U1369 (N_1369,In_1666,In_1867);
nor U1370 (N_1370,In_2314,In_1171);
and U1371 (N_1371,In_368,In_2377);
nand U1372 (N_1372,In_1681,In_1615);
nor U1373 (N_1373,In_979,In_602);
and U1374 (N_1374,In_670,In_1345);
nor U1375 (N_1375,In_533,In_181);
xor U1376 (N_1376,In_536,In_2471);
and U1377 (N_1377,In_1040,In_82);
nand U1378 (N_1378,In_2187,In_1404);
nand U1379 (N_1379,In_1009,In_1502);
or U1380 (N_1380,In_2261,In_2448);
xor U1381 (N_1381,In_303,In_757);
nor U1382 (N_1382,In_303,In_1009);
nor U1383 (N_1383,In_2110,In_516);
nand U1384 (N_1384,In_1861,In_1583);
xnor U1385 (N_1385,In_1929,In_1221);
xnor U1386 (N_1386,In_563,In_209);
nor U1387 (N_1387,In_730,In_708);
and U1388 (N_1388,In_2408,In_2495);
xnor U1389 (N_1389,In_236,In_81);
nor U1390 (N_1390,In_2141,In_2111);
and U1391 (N_1391,In_2224,In_836);
nor U1392 (N_1392,In_1377,In_323);
xnor U1393 (N_1393,In_74,In_2072);
nand U1394 (N_1394,In_416,In_600);
nor U1395 (N_1395,In_976,In_965);
and U1396 (N_1396,In_59,In_735);
nand U1397 (N_1397,In_531,In_439);
and U1398 (N_1398,In_1275,In_2393);
nand U1399 (N_1399,In_2029,In_739);
nand U1400 (N_1400,In_78,In_1931);
nand U1401 (N_1401,In_913,In_649);
and U1402 (N_1402,In_603,In_32);
or U1403 (N_1403,In_2471,In_1370);
xnor U1404 (N_1404,In_486,In_2436);
or U1405 (N_1405,In_1605,In_606);
xor U1406 (N_1406,In_544,In_1029);
xnor U1407 (N_1407,In_1623,In_266);
xnor U1408 (N_1408,In_1619,In_928);
nor U1409 (N_1409,In_2300,In_1150);
xor U1410 (N_1410,In_1585,In_577);
xor U1411 (N_1411,In_1931,In_46);
or U1412 (N_1412,In_735,In_48);
nor U1413 (N_1413,In_477,In_959);
nand U1414 (N_1414,In_2081,In_892);
xnor U1415 (N_1415,In_1510,In_1045);
nor U1416 (N_1416,In_48,In_142);
xnor U1417 (N_1417,In_1487,In_1195);
or U1418 (N_1418,In_1284,In_499);
or U1419 (N_1419,In_293,In_8);
and U1420 (N_1420,In_2340,In_1927);
xnor U1421 (N_1421,In_1521,In_1647);
xor U1422 (N_1422,In_2374,In_1601);
or U1423 (N_1423,In_2342,In_902);
xnor U1424 (N_1424,In_1906,In_1283);
nand U1425 (N_1425,In_1725,In_644);
nand U1426 (N_1426,In_2398,In_2273);
xnor U1427 (N_1427,In_811,In_826);
or U1428 (N_1428,In_383,In_1276);
nand U1429 (N_1429,In_446,In_540);
nand U1430 (N_1430,In_1688,In_1067);
xor U1431 (N_1431,In_922,In_1801);
and U1432 (N_1432,In_221,In_1328);
xnor U1433 (N_1433,In_2034,In_1334);
or U1434 (N_1434,In_2362,In_2247);
xnor U1435 (N_1435,In_1852,In_2101);
nor U1436 (N_1436,In_857,In_1663);
and U1437 (N_1437,In_888,In_980);
and U1438 (N_1438,In_1845,In_80);
nor U1439 (N_1439,In_1586,In_701);
nand U1440 (N_1440,In_1736,In_2133);
and U1441 (N_1441,In_1911,In_1930);
and U1442 (N_1442,In_1020,In_746);
and U1443 (N_1443,In_1615,In_2354);
nand U1444 (N_1444,In_1809,In_651);
or U1445 (N_1445,In_1280,In_464);
nor U1446 (N_1446,In_1503,In_1996);
xor U1447 (N_1447,In_2096,In_211);
or U1448 (N_1448,In_1371,In_416);
and U1449 (N_1449,In_2078,In_183);
nor U1450 (N_1450,In_2093,In_633);
xor U1451 (N_1451,In_1199,In_2017);
nor U1452 (N_1452,In_2437,In_1405);
xor U1453 (N_1453,In_1465,In_1346);
and U1454 (N_1454,In_1726,In_1569);
or U1455 (N_1455,In_835,In_1281);
and U1456 (N_1456,In_2299,In_265);
or U1457 (N_1457,In_2081,In_2332);
and U1458 (N_1458,In_1123,In_2464);
or U1459 (N_1459,In_2035,In_124);
and U1460 (N_1460,In_1639,In_1676);
and U1461 (N_1461,In_896,In_2419);
xor U1462 (N_1462,In_2390,In_1189);
and U1463 (N_1463,In_1617,In_950);
nand U1464 (N_1464,In_2482,In_2403);
and U1465 (N_1465,In_1931,In_1226);
xor U1466 (N_1466,In_531,In_90);
nor U1467 (N_1467,In_844,In_577);
and U1468 (N_1468,In_1611,In_1131);
xnor U1469 (N_1469,In_1809,In_1262);
and U1470 (N_1470,In_1690,In_1483);
nor U1471 (N_1471,In_2340,In_816);
or U1472 (N_1472,In_258,In_1247);
and U1473 (N_1473,In_2341,In_311);
or U1474 (N_1474,In_1690,In_282);
and U1475 (N_1475,In_1984,In_1167);
nor U1476 (N_1476,In_2414,In_1572);
nand U1477 (N_1477,In_1473,In_767);
and U1478 (N_1478,In_2175,In_1214);
nand U1479 (N_1479,In_2418,In_1643);
nand U1480 (N_1480,In_481,In_1506);
or U1481 (N_1481,In_1597,In_252);
and U1482 (N_1482,In_2060,In_2013);
nor U1483 (N_1483,In_950,In_1326);
and U1484 (N_1484,In_2316,In_2412);
xor U1485 (N_1485,In_2464,In_1094);
xnor U1486 (N_1486,In_835,In_48);
or U1487 (N_1487,In_268,In_1716);
and U1488 (N_1488,In_861,In_1603);
xnor U1489 (N_1489,In_2208,In_41);
or U1490 (N_1490,In_1670,In_2225);
nor U1491 (N_1491,In_1957,In_1586);
xnor U1492 (N_1492,In_1580,In_2336);
nor U1493 (N_1493,In_60,In_536);
nand U1494 (N_1494,In_655,In_1167);
and U1495 (N_1495,In_2194,In_295);
and U1496 (N_1496,In_1389,In_2314);
or U1497 (N_1497,In_1602,In_160);
and U1498 (N_1498,In_1376,In_2437);
xnor U1499 (N_1499,In_429,In_1433);
nor U1500 (N_1500,In_1913,In_2143);
nor U1501 (N_1501,In_859,In_2152);
or U1502 (N_1502,In_1024,In_1240);
xnor U1503 (N_1503,In_800,In_221);
nor U1504 (N_1504,In_224,In_592);
nand U1505 (N_1505,In_1319,In_569);
xor U1506 (N_1506,In_2097,In_502);
xnor U1507 (N_1507,In_1531,In_569);
or U1508 (N_1508,In_545,In_230);
xor U1509 (N_1509,In_2003,In_422);
and U1510 (N_1510,In_613,In_347);
and U1511 (N_1511,In_564,In_2309);
and U1512 (N_1512,In_1032,In_1475);
and U1513 (N_1513,In_253,In_1972);
and U1514 (N_1514,In_2353,In_942);
nand U1515 (N_1515,In_13,In_1524);
nor U1516 (N_1516,In_168,In_36);
xor U1517 (N_1517,In_1624,In_15);
and U1518 (N_1518,In_667,In_185);
nor U1519 (N_1519,In_1080,In_1077);
nand U1520 (N_1520,In_2018,In_2350);
nand U1521 (N_1521,In_2264,In_1982);
nand U1522 (N_1522,In_2277,In_1641);
and U1523 (N_1523,In_1048,In_376);
nor U1524 (N_1524,In_701,In_236);
or U1525 (N_1525,In_1866,In_2446);
or U1526 (N_1526,In_1161,In_743);
nand U1527 (N_1527,In_1580,In_859);
nor U1528 (N_1528,In_749,In_1653);
xnor U1529 (N_1529,In_1795,In_2244);
and U1530 (N_1530,In_2046,In_2192);
nand U1531 (N_1531,In_962,In_106);
xnor U1532 (N_1532,In_900,In_803);
or U1533 (N_1533,In_199,In_1937);
nand U1534 (N_1534,In_67,In_1915);
or U1535 (N_1535,In_2149,In_1225);
nor U1536 (N_1536,In_2378,In_907);
or U1537 (N_1537,In_732,In_2185);
nand U1538 (N_1538,In_1577,In_372);
and U1539 (N_1539,In_2125,In_2064);
nand U1540 (N_1540,In_1494,In_647);
or U1541 (N_1541,In_1444,In_2362);
xor U1542 (N_1542,In_946,In_1424);
or U1543 (N_1543,In_91,In_1541);
and U1544 (N_1544,In_1890,In_2442);
or U1545 (N_1545,In_1027,In_1235);
xnor U1546 (N_1546,In_2012,In_141);
xnor U1547 (N_1547,In_920,In_2384);
nand U1548 (N_1548,In_1037,In_837);
xnor U1549 (N_1549,In_2174,In_286);
or U1550 (N_1550,In_115,In_2235);
or U1551 (N_1551,In_1215,In_1832);
xnor U1552 (N_1552,In_1731,In_1378);
nand U1553 (N_1553,In_132,In_2483);
nor U1554 (N_1554,In_1845,In_1681);
or U1555 (N_1555,In_604,In_1992);
nor U1556 (N_1556,In_1634,In_243);
nor U1557 (N_1557,In_940,In_265);
nand U1558 (N_1558,In_1175,In_961);
xnor U1559 (N_1559,In_1702,In_1150);
or U1560 (N_1560,In_223,In_1834);
or U1561 (N_1561,In_1181,In_1912);
or U1562 (N_1562,In_2405,In_1417);
nand U1563 (N_1563,In_1603,In_12);
nor U1564 (N_1564,In_1267,In_851);
xnor U1565 (N_1565,In_2123,In_737);
and U1566 (N_1566,In_2434,In_1364);
nor U1567 (N_1567,In_564,In_1371);
xnor U1568 (N_1568,In_1399,In_361);
xor U1569 (N_1569,In_1222,In_1701);
or U1570 (N_1570,In_2207,In_2141);
xnor U1571 (N_1571,In_1152,In_1839);
or U1572 (N_1572,In_2110,In_1605);
or U1573 (N_1573,In_1387,In_2053);
and U1574 (N_1574,In_957,In_1422);
nor U1575 (N_1575,In_893,In_1213);
xor U1576 (N_1576,In_2082,In_1066);
or U1577 (N_1577,In_2212,In_981);
xnor U1578 (N_1578,In_996,In_2485);
nand U1579 (N_1579,In_2264,In_2208);
xnor U1580 (N_1580,In_1949,In_1477);
and U1581 (N_1581,In_260,In_2363);
or U1582 (N_1582,In_91,In_2144);
or U1583 (N_1583,In_775,In_938);
and U1584 (N_1584,In_1454,In_723);
nand U1585 (N_1585,In_1389,In_488);
xor U1586 (N_1586,In_283,In_2263);
nor U1587 (N_1587,In_2168,In_1309);
nand U1588 (N_1588,In_1152,In_1127);
nor U1589 (N_1589,In_1808,In_1106);
nor U1590 (N_1590,In_1304,In_2133);
nand U1591 (N_1591,In_1807,In_1634);
nand U1592 (N_1592,In_1833,In_40);
nor U1593 (N_1593,In_2171,In_132);
or U1594 (N_1594,In_1421,In_264);
and U1595 (N_1595,In_1731,In_1782);
nor U1596 (N_1596,In_33,In_939);
nand U1597 (N_1597,In_1128,In_2427);
nor U1598 (N_1598,In_312,In_1335);
nor U1599 (N_1599,In_2490,In_1923);
nor U1600 (N_1600,In_373,In_1908);
xnor U1601 (N_1601,In_65,In_16);
xnor U1602 (N_1602,In_1853,In_1384);
xnor U1603 (N_1603,In_627,In_84);
xor U1604 (N_1604,In_1497,In_701);
xor U1605 (N_1605,In_836,In_2455);
or U1606 (N_1606,In_504,In_391);
nand U1607 (N_1607,In_82,In_1750);
nand U1608 (N_1608,In_347,In_251);
xor U1609 (N_1609,In_1812,In_640);
xnor U1610 (N_1610,In_972,In_2478);
xor U1611 (N_1611,In_1319,In_2327);
and U1612 (N_1612,In_1347,In_272);
or U1613 (N_1613,In_929,In_2081);
nor U1614 (N_1614,In_1704,In_1282);
or U1615 (N_1615,In_512,In_1500);
and U1616 (N_1616,In_837,In_2399);
or U1617 (N_1617,In_2242,In_755);
nand U1618 (N_1618,In_2253,In_1098);
or U1619 (N_1619,In_1038,In_788);
xor U1620 (N_1620,In_753,In_857);
or U1621 (N_1621,In_452,In_2141);
or U1622 (N_1622,In_2243,In_9);
xor U1623 (N_1623,In_1691,In_1315);
nand U1624 (N_1624,In_205,In_60);
and U1625 (N_1625,In_1446,In_837);
xnor U1626 (N_1626,In_1011,In_1490);
nand U1627 (N_1627,In_2245,In_8);
nand U1628 (N_1628,In_1237,In_2094);
or U1629 (N_1629,In_1387,In_1107);
xor U1630 (N_1630,In_794,In_144);
nor U1631 (N_1631,In_1732,In_1498);
nor U1632 (N_1632,In_420,In_2309);
nand U1633 (N_1633,In_2239,In_198);
xnor U1634 (N_1634,In_26,In_1574);
nor U1635 (N_1635,In_1873,In_2277);
and U1636 (N_1636,In_413,In_1757);
or U1637 (N_1637,In_1230,In_1831);
xor U1638 (N_1638,In_1047,In_85);
and U1639 (N_1639,In_2159,In_1199);
and U1640 (N_1640,In_951,In_2351);
nor U1641 (N_1641,In_1529,In_1722);
or U1642 (N_1642,In_2066,In_1702);
and U1643 (N_1643,In_1277,In_38);
nor U1644 (N_1644,In_41,In_347);
nor U1645 (N_1645,In_1212,In_2455);
nand U1646 (N_1646,In_1590,In_2361);
and U1647 (N_1647,In_1594,In_2138);
and U1648 (N_1648,In_1180,In_1138);
or U1649 (N_1649,In_1720,In_1106);
xnor U1650 (N_1650,In_38,In_1814);
nor U1651 (N_1651,In_566,In_482);
and U1652 (N_1652,In_703,In_398);
nor U1653 (N_1653,In_272,In_698);
or U1654 (N_1654,In_572,In_1690);
xor U1655 (N_1655,In_973,In_1099);
and U1656 (N_1656,In_1244,In_1532);
nand U1657 (N_1657,In_1051,In_1909);
or U1658 (N_1658,In_1205,In_2222);
xnor U1659 (N_1659,In_2157,In_2057);
xnor U1660 (N_1660,In_2098,In_1049);
nor U1661 (N_1661,In_1586,In_2004);
nor U1662 (N_1662,In_1064,In_1995);
nor U1663 (N_1663,In_647,In_193);
nor U1664 (N_1664,In_1261,In_857);
nor U1665 (N_1665,In_30,In_27);
nand U1666 (N_1666,In_948,In_1051);
nor U1667 (N_1667,In_1562,In_1986);
nand U1668 (N_1668,In_1157,In_1654);
and U1669 (N_1669,In_1920,In_485);
nor U1670 (N_1670,In_125,In_632);
nand U1671 (N_1671,In_69,In_188);
or U1672 (N_1672,In_1645,In_796);
nor U1673 (N_1673,In_929,In_889);
nor U1674 (N_1674,In_1927,In_2158);
nand U1675 (N_1675,In_1732,In_618);
nand U1676 (N_1676,In_1538,In_1913);
nor U1677 (N_1677,In_1332,In_279);
or U1678 (N_1678,In_1350,In_1703);
xnor U1679 (N_1679,In_2050,In_1375);
and U1680 (N_1680,In_334,In_1367);
nor U1681 (N_1681,In_1167,In_230);
or U1682 (N_1682,In_1619,In_2448);
and U1683 (N_1683,In_1861,In_638);
nor U1684 (N_1684,In_62,In_214);
or U1685 (N_1685,In_1793,In_1494);
nand U1686 (N_1686,In_533,In_2406);
or U1687 (N_1687,In_19,In_618);
nand U1688 (N_1688,In_527,In_2495);
or U1689 (N_1689,In_1931,In_1581);
xnor U1690 (N_1690,In_330,In_1943);
nor U1691 (N_1691,In_560,In_2130);
or U1692 (N_1692,In_915,In_825);
nor U1693 (N_1693,In_1587,In_251);
nand U1694 (N_1694,In_194,In_1248);
xor U1695 (N_1695,In_866,In_611);
nor U1696 (N_1696,In_691,In_496);
and U1697 (N_1697,In_1356,In_451);
and U1698 (N_1698,In_2296,In_1083);
xor U1699 (N_1699,In_1146,In_228);
and U1700 (N_1700,In_1945,In_2133);
nand U1701 (N_1701,In_2434,In_2175);
and U1702 (N_1702,In_1379,In_441);
and U1703 (N_1703,In_1870,In_2318);
or U1704 (N_1704,In_658,In_2053);
nand U1705 (N_1705,In_766,In_60);
nand U1706 (N_1706,In_2142,In_1218);
nor U1707 (N_1707,In_1421,In_2316);
nor U1708 (N_1708,In_1432,In_1189);
nor U1709 (N_1709,In_284,In_2062);
nand U1710 (N_1710,In_40,In_906);
or U1711 (N_1711,In_1776,In_1124);
nand U1712 (N_1712,In_878,In_1422);
or U1713 (N_1713,In_901,In_1908);
or U1714 (N_1714,In_1990,In_2187);
or U1715 (N_1715,In_215,In_2362);
nor U1716 (N_1716,In_1497,In_945);
and U1717 (N_1717,In_1462,In_628);
nand U1718 (N_1718,In_636,In_235);
or U1719 (N_1719,In_1045,In_239);
nand U1720 (N_1720,In_1635,In_782);
nand U1721 (N_1721,In_11,In_1059);
nand U1722 (N_1722,In_1073,In_1021);
or U1723 (N_1723,In_695,In_517);
nand U1724 (N_1724,In_2479,In_1098);
nor U1725 (N_1725,In_1552,In_1190);
xor U1726 (N_1726,In_1297,In_2396);
or U1727 (N_1727,In_1876,In_667);
and U1728 (N_1728,In_2099,In_1355);
and U1729 (N_1729,In_1386,In_273);
nand U1730 (N_1730,In_468,In_2383);
xor U1731 (N_1731,In_537,In_428);
nand U1732 (N_1732,In_1953,In_2272);
nand U1733 (N_1733,In_663,In_144);
and U1734 (N_1734,In_1227,In_2310);
nand U1735 (N_1735,In_796,In_1160);
nor U1736 (N_1736,In_1819,In_1233);
or U1737 (N_1737,In_638,In_1225);
or U1738 (N_1738,In_2410,In_685);
nor U1739 (N_1739,In_845,In_840);
xor U1740 (N_1740,In_490,In_1388);
nor U1741 (N_1741,In_553,In_1112);
nand U1742 (N_1742,In_285,In_2437);
xor U1743 (N_1743,In_1233,In_2227);
or U1744 (N_1744,In_1015,In_753);
and U1745 (N_1745,In_1109,In_1744);
nor U1746 (N_1746,In_16,In_2138);
xnor U1747 (N_1747,In_2443,In_2006);
nor U1748 (N_1748,In_1823,In_1323);
or U1749 (N_1749,In_1969,In_1664);
or U1750 (N_1750,In_2308,In_1283);
nor U1751 (N_1751,In_129,In_1650);
nand U1752 (N_1752,In_1690,In_2008);
xnor U1753 (N_1753,In_877,In_938);
nor U1754 (N_1754,In_1685,In_1927);
nor U1755 (N_1755,In_1622,In_1404);
or U1756 (N_1756,In_198,In_367);
and U1757 (N_1757,In_2192,In_1414);
or U1758 (N_1758,In_1713,In_1118);
and U1759 (N_1759,In_2382,In_124);
xor U1760 (N_1760,In_1177,In_517);
nor U1761 (N_1761,In_1859,In_491);
and U1762 (N_1762,In_1335,In_2481);
nand U1763 (N_1763,In_38,In_148);
xnor U1764 (N_1764,In_2422,In_1274);
xnor U1765 (N_1765,In_781,In_2250);
or U1766 (N_1766,In_2499,In_124);
xor U1767 (N_1767,In_2120,In_2124);
or U1768 (N_1768,In_700,In_2172);
or U1769 (N_1769,In_711,In_2489);
xor U1770 (N_1770,In_1496,In_2040);
or U1771 (N_1771,In_288,In_1774);
nor U1772 (N_1772,In_480,In_1849);
and U1773 (N_1773,In_1126,In_1911);
nor U1774 (N_1774,In_149,In_553);
xor U1775 (N_1775,In_616,In_1805);
and U1776 (N_1776,In_4,In_12);
or U1777 (N_1777,In_1706,In_1024);
nand U1778 (N_1778,In_952,In_2008);
nor U1779 (N_1779,In_48,In_1319);
or U1780 (N_1780,In_1060,In_1961);
xnor U1781 (N_1781,In_260,In_1441);
nand U1782 (N_1782,In_466,In_2453);
or U1783 (N_1783,In_1019,In_907);
nor U1784 (N_1784,In_1809,In_968);
xnor U1785 (N_1785,In_710,In_1502);
nand U1786 (N_1786,In_2034,In_14);
and U1787 (N_1787,In_2361,In_1004);
or U1788 (N_1788,In_649,In_2302);
xnor U1789 (N_1789,In_1658,In_2407);
and U1790 (N_1790,In_751,In_1933);
or U1791 (N_1791,In_2410,In_2329);
nor U1792 (N_1792,In_410,In_1019);
nand U1793 (N_1793,In_1847,In_1927);
and U1794 (N_1794,In_31,In_489);
nor U1795 (N_1795,In_708,In_203);
nor U1796 (N_1796,In_2394,In_602);
xor U1797 (N_1797,In_1355,In_1973);
nand U1798 (N_1798,In_1903,In_1411);
or U1799 (N_1799,In_1688,In_611);
nor U1800 (N_1800,In_2241,In_549);
xnor U1801 (N_1801,In_68,In_640);
or U1802 (N_1802,In_938,In_1124);
nand U1803 (N_1803,In_2044,In_2083);
or U1804 (N_1804,In_1598,In_555);
and U1805 (N_1805,In_932,In_1350);
or U1806 (N_1806,In_1014,In_2394);
xnor U1807 (N_1807,In_343,In_373);
and U1808 (N_1808,In_78,In_1143);
and U1809 (N_1809,In_383,In_1495);
and U1810 (N_1810,In_1879,In_1309);
nor U1811 (N_1811,In_1381,In_2298);
nor U1812 (N_1812,In_381,In_1088);
or U1813 (N_1813,In_666,In_1630);
or U1814 (N_1814,In_1714,In_1373);
nor U1815 (N_1815,In_1021,In_454);
nand U1816 (N_1816,In_1046,In_1657);
and U1817 (N_1817,In_1767,In_2117);
nor U1818 (N_1818,In_1533,In_958);
or U1819 (N_1819,In_1640,In_1183);
or U1820 (N_1820,In_1604,In_2353);
xnor U1821 (N_1821,In_676,In_1276);
and U1822 (N_1822,In_303,In_1984);
nand U1823 (N_1823,In_1436,In_741);
nand U1824 (N_1824,In_111,In_2368);
and U1825 (N_1825,In_1306,In_1521);
nor U1826 (N_1826,In_1190,In_1390);
and U1827 (N_1827,In_2329,In_1562);
and U1828 (N_1828,In_440,In_1290);
and U1829 (N_1829,In_2254,In_55);
xor U1830 (N_1830,In_160,In_1192);
and U1831 (N_1831,In_1156,In_61);
or U1832 (N_1832,In_1322,In_388);
nand U1833 (N_1833,In_1122,In_2272);
or U1834 (N_1834,In_149,In_878);
nor U1835 (N_1835,In_234,In_677);
or U1836 (N_1836,In_410,In_2002);
nand U1837 (N_1837,In_67,In_1753);
or U1838 (N_1838,In_1367,In_873);
or U1839 (N_1839,In_35,In_210);
and U1840 (N_1840,In_26,In_746);
nor U1841 (N_1841,In_1767,In_2457);
nand U1842 (N_1842,In_0,In_2002);
nor U1843 (N_1843,In_289,In_791);
and U1844 (N_1844,In_2414,In_830);
nor U1845 (N_1845,In_94,In_1480);
nand U1846 (N_1846,In_2088,In_2412);
nor U1847 (N_1847,In_1917,In_1151);
nand U1848 (N_1848,In_1587,In_2263);
and U1849 (N_1849,In_1043,In_937);
xnor U1850 (N_1850,In_767,In_1628);
nand U1851 (N_1851,In_1677,In_1720);
nand U1852 (N_1852,In_886,In_2136);
nor U1853 (N_1853,In_1001,In_2054);
nor U1854 (N_1854,In_1423,In_2097);
xnor U1855 (N_1855,In_2060,In_2469);
nand U1856 (N_1856,In_1918,In_1075);
or U1857 (N_1857,In_2018,In_1425);
nand U1858 (N_1858,In_2118,In_916);
and U1859 (N_1859,In_636,In_739);
nand U1860 (N_1860,In_1033,In_1542);
nor U1861 (N_1861,In_1225,In_752);
nand U1862 (N_1862,In_1143,In_678);
and U1863 (N_1863,In_2288,In_2059);
xor U1864 (N_1864,In_2081,In_1620);
and U1865 (N_1865,In_273,In_647);
and U1866 (N_1866,In_740,In_936);
nand U1867 (N_1867,In_1334,In_554);
nand U1868 (N_1868,In_26,In_1737);
or U1869 (N_1869,In_1369,In_1823);
or U1870 (N_1870,In_2256,In_1222);
nand U1871 (N_1871,In_133,In_2294);
nand U1872 (N_1872,In_1423,In_1687);
nor U1873 (N_1873,In_737,In_1976);
and U1874 (N_1874,In_1643,In_1999);
and U1875 (N_1875,In_2158,In_922);
xor U1876 (N_1876,In_2242,In_1975);
or U1877 (N_1877,In_1491,In_727);
and U1878 (N_1878,In_1929,In_525);
nor U1879 (N_1879,In_1347,In_1380);
nand U1880 (N_1880,In_1984,In_519);
nor U1881 (N_1881,In_515,In_1604);
nand U1882 (N_1882,In_279,In_1624);
nor U1883 (N_1883,In_231,In_1385);
or U1884 (N_1884,In_2106,In_2120);
nor U1885 (N_1885,In_844,In_749);
nand U1886 (N_1886,In_2154,In_380);
nor U1887 (N_1887,In_366,In_1624);
xor U1888 (N_1888,In_909,In_1415);
nor U1889 (N_1889,In_1676,In_51);
and U1890 (N_1890,In_179,In_2337);
nor U1891 (N_1891,In_1137,In_1088);
nor U1892 (N_1892,In_921,In_1403);
or U1893 (N_1893,In_19,In_1307);
nor U1894 (N_1894,In_2038,In_1368);
nand U1895 (N_1895,In_648,In_2369);
nor U1896 (N_1896,In_1203,In_887);
or U1897 (N_1897,In_1152,In_639);
and U1898 (N_1898,In_1568,In_1664);
or U1899 (N_1899,In_1416,In_175);
and U1900 (N_1900,In_1561,In_1443);
and U1901 (N_1901,In_1073,In_1342);
or U1902 (N_1902,In_1251,In_710);
or U1903 (N_1903,In_1067,In_1765);
xnor U1904 (N_1904,In_2320,In_1011);
or U1905 (N_1905,In_1279,In_2474);
nor U1906 (N_1906,In_2008,In_2258);
nand U1907 (N_1907,In_1632,In_2324);
or U1908 (N_1908,In_214,In_382);
and U1909 (N_1909,In_1342,In_2015);
nor U1910 (N_1910,In_2355,In_2366);
xnor U1911 (N_1911,In_932,In_1634);
xnor U1912 (N_1912,In_0,In_1366);
nand U1913 (N_1913,In_1801,In_1334);
xnor U1914 (N_1914,In_1309,In_2197);
xor U1915 (N_1915,In_336,In_2264);
or U1916 (N_1916,In_1591,In_981);
and U1917 (N_1917,In_234,In_269);
xor U1918 (N_1918,In_2448,In_2325);
nor U1919 (N_1919,In_149,In_1068);
and U1920 (N_1920,In_2390,In_1828);
nand U1921 (N_1921,In_1884,In_392);
nor U1922 (N_1922,In_1216,In_2061);
xor U1923 (N_1923,In_459,In_66);
nor U1924 (N_1924,In_808,In_756);
and U1925 (N_1925,In_501,In_2434);
and U1926 (N_1926,In_1583,In_83);
nor U1927 (N_1927,In_1712,In_171);
nand U1928 (N_1928,In_1355,In_1950);
and U1929 (N_1929,In_266,In_1626);
nor U1930 (N_1930,In_77,In_919);
nand U1931 (N_1931,In_2326,In_674);
xnor U1932 (N_1932,In_987,In_2186);
nor U1933 (N_1933,In_572,In_2365);
nand U1934 (N_1934,In_1585,In_1096);
nand U1935 (N_1935,In_1321,In_59);
and U1936 (N_1936,In_1276,In_987);
or U1937 (N_1937,In_249,In_1525);
xor U1938 (N_1938,In_1610,In_1354);
nor U1939 (N_1939,In_1237,In_2142);
nand U1940 (N_1940,In_1255,In_1021);
nor U1941 (N_1941,In_732,In_190);
or U1942 (N_1942,In_1610,In_2307);
or U1943 (N_1943,In_2417,In_2223);
xnor U1944 (N_1944,In_1124,In_1198);
xor U1945 (N_1945,In_953,In_1736);
nand U1946 (N_1946,In_1850,In_270);
or U1947 (N_1947,In_1839,In_1113);
or U1948 (N_1948,In_908,In_1957);
nor U1949 (N_1949,In_1751,In_814);
and U1950 (N_1950,In_398,In_1263);
nor U1951 (N_1951,In_13,In_1700);
or U1952 (N_1952,In_588,In_916);
or U1953 (N_1953,In_445,In_1332);
and U1954 (N_1954,In_1847,In_314);
nor U1955 (N_1955,In_2351,In_1833);
xnor U1956 (N_1956,In_42,In_597);
xnor U1957 (N_1957,In_559,In_2399);
nor U1958 (N_1958,In_2431,In_986);
nand U1959 (N_1959,In_1741,In_1285);
and U1960 (N_1960,In_890,In_826);
xnor U1961 (N_1961,In_2427,In_791);
and U1962 (N_1962,In_2250,In_1042);
or U1963 (N_1963,In_2196,In_1783);
nand U1964 (N_1964,In_51,In_1606);
nand U1965 (N_1965,In_2310,In_2005);
nand U1966 (N_1966,In_334,In_820);
or U1967 (N_1967,In_1056,In_1346);
nor U1968 (N_1968,In_8,In_1452);
xor U1969 (N_1969,In_1204,In_1828);
and U1970 (N_1970,In_2495,In_1140);
or U1971 (N_1971,In_1252,In_1151);
nand U1972 (N_1972,In_297,In_2148);
xnor U1973 (N_1973,In_1309,In_491);
or U1974 (N_1974,In_1823,In_481);
or U1975 (N_1975,In_349,In_296);
and U1976 (N_1976,In_333,In_2473);
or U1977 (N_1977,In_1002,In_893);
xnor U1978 (N_1978,In_109,In_287);
or U1979 (N_1979,In_1079,In_699);
xor U1980 (N_1980,In_1539,In_1368);
or U1981 (N_1981,In_1827,In_2072);
xor U1982 (N_1982,In_680,In_1611);
nor U1983 (N_1983,In_570,In_239);
and U1984 (N_1984,In_541,In_2020);
or U1985 (N_1985,In_1175,In_1288);
or U1986 (N_1986,In_1078,In_474);
nor U1987 (N_1987,In_1026,In_779);
nand U1988 (N_1988,In_2461,In_323);
and U1989 (N_1989,In_702,In_503);
xor U1990 (N_1990,In_1357,In_1897);
nor U1991 (N_1991,In_2440,In_1432);
and U1992 (N_1992,In_95,In_1355);
or U1993 (N_1993,In_1045,In_916);
xor U1994 (N_1994,In_2063,In_555);
xnor U1995 (N_1995,In_135,In_1262);
or U1996 (N_1996,In_2227,In_1035);
nor U1997 (N_1997,In_1936,In_743);
nor U1998 (N_1998,In_1231,In_1287);
nor U1999 (N_1999,In_1961,In_1476);
nor U2000 (N_2000,In_341,In_1063);
nor U2001 (N_2001,In_93,In_605);
xor U2002 (N_2002,In_1559,In_1778);
nor U2003 (N_2003,In_2038,In_1326);
or U2004 (N_2004,In_1787,In_1279);
nor U2005 (N_2005,In_818,In_1655);
xnor U2006 (N_2006,In_1650,In_1225);
and U2007 (N_2007,In_1572,In_1558);
xor U2008 (N_2008,In_16,In_1084);
xnor U2009 (N_2009,In_263,In_98);
and U2010 (N_2010,In_992,In_1754);
and U2011 (N_2011,In_1268,In_1533);
nor U2012 (N_2012,In_554,In_1433);
xnor U2013 (N_2013,In_1616,In_284);
xnor U2014 (N_2014,In_1924,In_2469);
or U2015 (N_2015,In_1940,In_1864);
xor U2016 (N_2016,In_825,In_1780);
xor U2017 (N_2017,In_394,In_1538);
and U2018 (N_2018,In_2314,In_616);
and U2019 (N_2019,In_652,In_2011);
nor U2020 (N_2020,In_1413,In_1485);
and U2021 (N_2021,In_1842,In_378);
or U2022 (N_2022,In_1758,In_128);
or U2023 (N_2023,In_1337,In_2018);
nor U2024 (N_2024,In_1613,In_1713);
nor U2025 (N_2025,In_1250,In_2221);
nor U2026 (N_2026,In_1583,In_421);
or U2027 (N_2027,In_2158,In_1749);
xnor U2028 (N_2028,In_129,In_2210);
nand U2029 (N_2029,In_270,In_2456);
and U2030 (N_2030,In_1767,In_1070);
or U2031 (N_2031,In_703,In_1951);
or U2032 (N_2032,In_1168,In_300);
or U2033 (N_2033,In_1050,In_231);
nand U2034 (N_2034,In_1430,In_2210);
or U2035 (N_2035,In_2348,In_2463);
or U2036 (N_2036,In_1362,In_1056);
and U2037 (N_2037,In_1984,In_1879);
xor U2038 (N_2038,In_1149,In_809);
nor U2039 (N_2039,In_2417,In_128);
nand U2040 (N_2040,In_2310,In_2094);
nand U2041 (N_2041,In_2265,In_1828);
or U2042 (N_2042,In_1052,In_2334);
and U2043 (N_2043,In_835,In_1701);
nand U2044 (N_2044,In_1201,In_2401);
and U2045 (N_2045,In_2325,In_1631);
or U2046 (N_2046,In_702,In_2431);
nand U2047 (N_2047,In_263,In_945);
or U2048 (N_2048,In_403,In_1862);
nor U2049 (N_2049,In_649,In_1162);
or U2050 (N_2050,In_1875,In_360);
nand U2051 (N_2051,In_1241,In_1619);
xnor U2052 (N_2052,In_52,In_321);
and U2053 (N_2053,In_1278,In_850);
nand U2054 (N_2054,In_1679,In_1447);
xnor U2055 (N_2055,In_1678,In_577);
nor U2056 (N_2056,In_2170,In_2131);
nor U2057 (N_2057,In_2275,In_2073);
xor U2058 (N_2058,In_965,In_983);
nand U2059 (N_2059,In_944,In_336);
xnor U2060 (N_2060,In_1544,In_928);
nand U2061 (N_2061,In_815,In_2212);
nor U2062 (N_2062,In_548,In_558);
and U2063 (N_2063,In_1425,In_765);
xor U2064 (N_2064,In_48,In_1493);
xnor U2065 (N_2065,In_1765,In_1709);
and U2066 (N_2066,In_1794,In_1536);
xor U2067 (N_2067,In_1403,In_1439);
and U2068 (N_2068,In_595,In_1517);
xnor U2069 (N_2069,In_1708,In_2303);
nand U2070 (N_2070,In_825,In_708);
nor U2071 (N_2071,In_52,In_585);
and U2072 (N_2072,In_1312,In_1647);
nor U2073 (N_2073,In_940,In_1078);
and U2074 (N_2074,In_2444,In_302);
nor U2075 (N_2075,In_505,In_853);
xor U2076 (N_2076,In_1388,In_167);
xnor U2077 (N_2077,In_2250,In_1232);
nand U2078 (N_2078,In_1218,In_2402);
nor U2079 (N_2079,In_2445,In_293);
xnor U2080 (N_2080,In_981,In_992);
and U2081 (N_2081,In_2395,In_1991);
or U2082 (N_2082,In_979,In_745);
or U2083 (N_2083,In_2292,In_1759);
nand U2084 (N_2084,In_2427,In_263);
and U2085 (N_2085,In_701,In_1413);
xor U2086 (N_2086,In_424,In_326);
or U2087 (N_2087,In_797,In_1577);
or U2088 (N_2088,In_2440,In_944);
and U2089 (N_2089,In_1944,In_1398);
and U2090 (N_2090,In_1258,In_980);
and U2091 (N_2091,In_1578,In_927);
nand U2092 (N_2092,In_966,In_1279);
nand U2093 (N_2093,In_1484,In_879);
and U2094 (N_2094,In_1907,In_977);
nand U2095 (N_2095,In_1737,In_929);
xor U2096 (N_2096,In_218,In_1374);
nand U2097 (N_2097,In_2065,In_157);
nor U2098 (N_2098,In_1430,In_1873);
or U2099 (N_2099,In_1968,In_248);
xor U2100 (N_2100,In_990,In_2193);
and U2101 (N_2101,In_2371,In_2471);
nor U2102 (N_2102,In_767,In_2240);
and U2103 (N_2103,In_1758,In_444);
xor U2104 (N_2104,In_872,In_659);
nand U2105 (N_2105,In_2410,In_1543);
nor U2106 (N_2106,In_1671,In_1694);
or U2107 (N_2107,In_2258,In_856);
and U2108 (N_2108,In_1006,In_1547);
and U2109 (N_2109,In_1299,In_666);
xnor U2110 (N_2110,In_2187,In_1199);
or U2111 (N_2111,In_1498,In_1055);
or U2112 (N_2112,In_2191,In_826);
nor U2113 (N_2113,In_2272,In_1611);
nor U2114 (N_2114,In_1825,In_1249);
nand U2115 (N_2115,In_686,In_1763);
and U2116 (N_2116,In_829,In_1448);
or U2117 (N_2117,In_391,In_2179);
nand U2118 (N_2118,In_2026,In_1380);
nor U2119 (N_2119,In_647,In_94);
or U2120 (N_2120,In_1488,In_1345);
nor U2121 (N_2121,In_2052,In_1719);
or U2122 (N_2122,In_237,In_2473);
nor U2123 (N_2123,In_923,In_567);
xnor U2124 (N_2124,In_1602,In_1009);
xnor U2125 (N_2125,In_583,In_967);
and U2126 (N_2126,In_927,In_1760);
and U2127 (N_2127,In_700,In_637);
or U2128 (N_2128,In_560,In_826);
or U2129 (N_2129,In_1676,In_2255);
nor U2130 (N_2130,In_266,In_1135);
nand U2131 (N_2131,In_606,In_1694);
xor U2132 (N_2132,In_1872,In_2440);
nand U2133 (N_2133,In_890,In_1055);
nand U2134 (N_2134,In_544,In_392);
and U2135 (N_2135,In_127,In_947);
and U2136 (N_2136,In_1078,In_224);
and U2137 (N_2137,In_1879,In_1176);
xor U2138 (N_2138,In_2118,In_840);
nand U2139 (N_2139,In_1406,In_2480);
xnor U2140 (N_2140,In_2170,In_2107);
and U2141 (N_2141,In_1823,In_2073);
and U2142 (N_2142,In_1803,In_445);
nor U2143 (N_2143,In_2292,In_1789);
xnor U2144 (N_2144,In_1461,In_2262);
xnor U2145 (N_2145,In_866,In_1133);
and U2146 (N_2146,In_2145,In_464);
or U2147 (N_2147,In_1142,In_1792);
and U2148 (N_2148,In_958,In_408);
nor U2149 (N_2149,In_1207,In_2181);
xor U2150 (N_2150,In_176,In_822);
nor U2151 (N_2151,In_469,In_2308);
xnor U2152 (N_2152,In_1897,In_2010);
or U2153 (N_2153,In_1892,In_1962);
xnor U2154 (N_2154,In_545,In_267);
and U2155 (N_2155,In_428,In_547);
and U2156 (N_2156,In_1194,In_1897);
or U2157 (N_2157,In_239,In_1491);
or U2158 (N_2158,In_2094,In_335);
xor U2159 (N_2159,In_2462,In_1094);
or U2160 (N_2160,In_1113,In_2308);
or U2161 (N_2161,In_2274,In_842);
nand U2162 (N_2162,In_2375,In_2244);
or U2163 (N_2163,In_67,In_2382);
nand U2164 (N_2164,In_1354,In_2049);
and U2165 (N_2165,In_1852,In_1210);
xor U2166 (N_2166,In_1045,In_2244);
and U2167 (N_2167,In_814,In_1243);
nand U2168 (N_2168,In_2386,In_2151);
nor U2169 (N_2169,In_2106,In_1854);
xor U2170 (N_2170,In_599,In_464);
and U2171 (N_2171,In_267,In_435);
or U2172 (N_2172,In_12,In_142);
nor U2173 (N_2173,In_869,In_295);
xnor U2174 (N_2174,In_1902,In_1515);
nor U2175 (N_2175,In_34,In_42);
nand U2176 (N_2176,In_294,In_88);
nor U2177 (N_2177,In_2142,In_1439);
and U2178 (N_2178,In_1377,In_1595);
nand U2179 (N_2179,In_1817,In_1689);
nor U2180 (N_2180,In_2402,In_1515);
and U2181 (N_2181,In_223,In_1217);
xnor U2182 (N_2182,In_626,In_224);
or U2183 (N_2183,In_1292,In_1073);
nor U2184 (N_2184,In_1313,In_2164);
nor U2185 (N_2185,In_1381,In_527);
nor U2186 (N_2186,In_891,In_811);
or U2187 (N_2187,In_811,In_2035);
or U2188 (N_2188,In_2143,In_749);
and U2189 (N_2189,In_2197,In_2490);
or U2190 (N_2190,In_2066,In_1916);
nor U2191 (N_2191,In_1500,In_249);
or U2192 (N_2192,In_1163,In_2408);
nand U2193 (N_2193,In_1524,In_543);
nand U2194 (N_2194,In_2293,In_1847);
nor U2195 (N_2195,In_978,In_1551);
nor U2196 (N_2196,In_682,In_1488);
and U2197 (N_2197,In_1672,In_2290);
and U2198 (N_2198,In_2477,In_1685);
xor U2199 (N_2199,In_953,In_73);
and U2200 (N_2200,In_663,In_39);
and U2201 (N_2201,In_1548,In_2120);
nor U2202 (N_2202,In_2412,In_1932);
or U2203 (N_2203,In_2267,In_1474);
nand U2204 (N_2204,In_1052,In_744);
xor U2205 (N_2205,In_1758,In_2206);
and U2206 (N_2206,In_2249,In_1512);
and U2207 (N_2207,In_2025,In_883);
xnor U2208 (N_2208,In_1795,In_979);
or U2209 (N_2209,In_2465,In_1212);
or U2210 (N_2210,In_1759,In_796);
and U2211 (N_2211,In_834,In_912);
nor U2212 (N_2212,In_355,In_32);
nand U2213 (N_2213,In_870,In_453);
or U2214 (N_2214,In_1600,In_782);
nor U2215 (N_2215,In_124,In_997);
nand U2216 (N_2216,In_1441,In_2374);
and U2217 (N_2217,In_1574,In_1496);
xor U2218 (N_2218,In_294,In_359);
nand U2219 (N_2219,In_2026,In_1491);
nand U2220 (N_2220,In_1299,In_2158);
or U2221 (N_2221,In_1801,In_645);
xnor U2222 (N_2222,In_108,In_1270);
xor U2223 (N_2223,In_342,In_508);
xor U2224 (N_2224,In_2041,In_1882);
nand U2225 (N_2225,In_2064,In_479);
xor U2226 (N_2226,In_1187,In_1966);
nand U2227 (N_2227,In_1408,In_888);
nand U2228 (N_2228,In_1972,In_650);
xnor U2229 (N_2229,In_894,In_1258);
nand U2230 (N_2230,In_2119,In_2405);
or U2231 (N_2231,In_167,In_199);
nand U2232 (N_2232,In_1745,In_1287);
xor U2233 (N_2233,In_2083,In_493);
or U2234 (N_2234,In_1430,In_843);
nand U2235 (N_2235,In_219,In_1395);
and U2236 (N_2236,In_1228,In_1987);
and U2237 (N_2237,In_171,In_1505);
or U2238 (N_2238,In_1001,In_1745);
nor U2239 (N_2239,In_1159,In_85);
nor U2240 (N_2240,In_603,In_699);
xnor U2241 (N_2241,In_1622,In_1076);
nand U2242 (N_2242,In_1905,In_290);
nor U2243 (N_2243,In_1864,In_783);
nand U2244 (N_2244,In_233,In_367);
xnor U2245 (N_2245,In_2299,In_80);
nor U2246 (N_2246,In_1719,In_59);
nand U2247 (N_2247,In_1596,In_2201);
nand U2248 (N_2248,In_2204,In_790);
or U2249 (N_2249,In_280,In_406);
or U2250 (N_2250,In_28,In_1735);
nand U2251 (N_2251,In_1418,In_256);
nand U2252 (N_2252,In_811,In_83);
or U2253 (N_2253,In_1268,In_998);
xor U2254 (N_2254,In_1548,In_93);
nor U2255 (N_2255,In_1385,In_1488);
xnor U2256 (N_2256,In_914,In_1208);
xor U2257 (N_2257,In_851,In_881);
nand U2258 (N_2258,In_2122,In_985);
or U2259 (N_2259,In_335,In_570);
nor U2260 (N_2260,In_1557,In_308);
and U2261 (N_2261,In_695,In_2437);
xnor U2262 (N_2262,In_794,In_2169);
and U2263 (N_2263,In_843,In_1869);
xor U2264 (N_2264,In_1879,In_922);
or U2265 (N_2265,In_2239,In_141);
and U2266 (N_2266,In_519,In_815);
nand U2267 (N_2267,In_2396,In_1323);
nor U2268 (N_2268,In_1513,In_608);
nor U2269 (N_2269,In_2161,In_1986);
and U2270 (N_2270,In_834,In_2098);
nand U2271 (N_2271,In_975,In_2455);
nand U2272 (N_2272,In_649,In_557);
or U2273 (N_2273,In_455,In_1994);
nand U2274 (N_2274,In_237,In_2077);
and U2275 (N_2275,In_927,In_2083);
nor U2276 (N_2276,In_1117,In_1246);
nand U2277 (N_2277,In_1431,In_628);
nor U2278 (N_2278,In_198,In_976);
or U2279 (N_2279,In_1250,In_1744);
nand U2280 (N_2280,In_1751,In_65);
xnor U2281 (N_2281,In_1411,In_879);
or U2282 (N_2282,In_1869,In_1724);
and U2283 (N_2283,In_2134,In_1941);
or U2284 (N_2284,In_1309,In_1724);
nand U2285 (N_2285,In_2464,In_1584);
or U2286 (N_2286,In_474,In_1336);
or U2287 (N_2287,In_1452,In_957);
or U2288 (N_2288,In_770,In_312);
or U2289 (N_2289,In_461,In_238);
xnor U2290 (N_2290,In_2016,In_2167);
nand U2291 (N_2291,In_2219,In_908);
or U2292 (N_2292,In_1221,In_2224);
xor U2293 (N_2293,In_1522,In_1007);
nand U2294 (N_2294,In_705,In_589);
and U2295 (N_2295,In_1419,In_520);
and U2296 (N_2296,In_69,In_1353);
nor U2297 (N_2297,In_234,In_25);
nor U2298 (N_2298,In_954,In_2);
nand U2299 (N_2299,In_2214,In_1865);
nand U2300 (N_2300,In_265,In_239);
and U2301 (N_2301,In_444,In_1618);
and U2302 (N_2302,In_1947,In_674);
and U2303 (N_2303,In_2277,In_1110);
nand U2304 (N_2304,In_834,In_1110);
nor U2305 (N_2305,In_1334,In_992);
and U2306 (N_2306,In_811,In_1970);
or U2307 (N_2307,In_573,In_590);
nor U2308 (N_2308,In_2474,In_914);
nor U2309 (N_2309,In_650,In_2286);
xnor U2310 (N_2310,In_1848,In_1147);
and U2311 (N_2311,In_1902,In_1236);
nor U2312 (N_2312,In_1728,In_2381);
nor U2313 (N_2313,In_1932,In_487);
nand U2314 (N_2314,In_14,In_1839);
or U2315 (N_2315,In_2340,In_1132);
and U2316 (N_2316,In_1319,In_2018);
xor U2317 (N_2317,In_2426,In_430);
xor U2318 (N_2318,In_699,In_1421);
nand U2319 (N_2319,In_128,In_1769);
nand U2320 (N_2320,In_285,In_495);
and U2321 (N_2321,In_752,In_47);
nor U2322 (N_2322,In_1230,In_2411);
nand U2323 (N_2323,In_2017,In_1833);
or U2324 (N_2324,In_2493,In_2013);
nand U2325 (N_2325,In_1860,In_492);
or U2326 (N_2326,In_1742,In_1404);
nand U2327 (N_2327,In_1759,In_271);
nor U2328 (N_2328,In_1945,In_391);
and U2329 (N_2329,In_1760,In_359);
nor U2330 (N_2330,In_1895,In_1645);
and U2331 (N_2331,In_577,In_1962);
xor U2332 (N_2332,In_2153,In_1015);
or U2333 (N_2333,In_1311,In_1891);
and U2334 (N_2334,In_1829,In_1713);
xnor U2335 (N_2335,In_2363,In_1961);
or U2336 (N_2336,In_1371,In_1605);
or U2337 (N_2337,In_331,In_2062);
or U2338 (N_2338,In_1854,In_1511);
nand U2339 (N_2339,In_371,In_1702);
xnor U2340 (N_2340,In_1007,In_2157);
and U2341 (N_2341,In_1226,In_1042);
nor U2342 (N_2342,In_2454,In_445);
xor U2343 (N_2343,In_1819,In_1265);
and U2344 (N_2344,In_2217,In_2140);
or U2345 (N_2345,In_2309,In_2081);
and U2346 (N_2346,In_100,In_871);
nand U2347 (N_2347,In_1286,In_2015);
and U2348 (N_2348,In_1049,In_473);
nand U2349 (N_2349,In_1118,In_1505);
xnor U2350 (N_2350,In_1069,In_368);
nand U2351 (N_2351,In_818,In_1440);
nand U2352 (N_2352,In_2481,In_1406);
nand U2353 (N_2353,In_61,In_1019);
nand U2354 (N_2354,In_1034,In_1971);
nand U2355 (N_2355,In_237,In_841);
and U2356 (N_2356,In_754,In_235);
nor U2357 (N_2357,In_419,In_167);
xnor U2358 (N_2358,In_755,In_1197);
nor U2359 (N_2359,In_374,In_1505);
nand U2360 (N_2360,In_1465,In_1910);
nand U2361 (N_2361,In_1693,In_1195);
nor U2362 (N_2362,In_1802,In_841);
and U2363 (N_2363,In_434,In_1556);
and U2364 (N_2364,In_404,In_957);
and U2365 (N_2365,In_2291,In_1776);
xor U2366 (N_2366,In_2378,In_2198);
and U2367 (N_2367,In_1208,In_1690);
and U2368 (N_2368,In_2042,In_431);
or U2369 (N_2369,In_1047,In_2254);
and U2370 (N_2370,In_2197,In_1210);
xnor U2371 (N_2371,In_1891,In_774);
and U2372 (N_2372,In_485,In_501);
nand U2373 (N_2373,In_1459,In_171);
xor U2374 (N_2374,In_1815,In_825);
or U2375 (N_2375,In_2363,In_963);
nand U2376 (N_2376,In_614,In_1908);
nand U2377 (N_2377,In_779,In_1404);
and U2378 (N_2378,In_1313,In_2341);
nand U2379 (N_2379,In_1398,In_1137);
nand U2380 (N_2380,In_1441,In_878);
xnor U2381 (N_2381,In_1692,In_15);
nor U2382 (N_2382,In_2123,In_704);
nand U2383 (N_2383,In_1031,In_1310);
nor U2384 (N_2384,In_417,In_1952);
nand U2385 (N_2385,In_1846,In_1624);
and U2386 (N_2386,In_401,In_320);
nor U2387 (N_2387,In_2088,In_2041);
xnor U2388 (N_2388,In_360,In_2298);
and U2389 (N_2389,In_1303,In_170);
nor U2390 (N_2390,In_2494,In_385);
nand U2391 (N_2391,In_1161,In_1337);
or U2392 (N_2392,In_969,In_933);
nor U2393 (N_2393,In_627,In_919);
xnor U2394 (N_2394,In_1293,In_2411);
xor U2395 (N_2395,In_792,In_587);
and U2396 (N_2396,In_2180,In_1099);
and U2397 (N_2397,In_323,In_1167);
nand U2398 (N_2398,In_280,In_2379);
nand U2399 (N_2399,In_774,In_2353);
nand U2400 (N_2400,In_1950,In_2284);
nand U2401 (N_2401,In_1590,In_2080);
nor U2402 (N_2402,In_984,In_1193);
or U2403 (N_2403,In_1023,In_785);
and U2404 (N_2404,In_1552,In_80);
nand U2405 (N_2405,In_1445,In_991);
nand U2406 (N_2406,In_1290,In_2197);
xnor U2407 (N_2407,In_29,In_1039);
and U2408 (N_2408,In_1011,In_116);
nor U2409 (N_2409,In_2122,In_1242);
xnor U2410 (N_2410,In_721,In_2179);
and U2411 (N_2411,In_306,In_1389);
nand U2412 (N_2412,In_1141,In_1653);
and U2413 (N_2413,In_510,In_1751);
nor U2414 (N_2414,In_2105,In_841);
xnor U2415 (N_2415,In_452,In_456);
or U2416 (N_2416,In_1348,In_2311);
xnor U2417 (N_2417,In_1030,In_1475);
xor U2418 (N_2418,In_1956,In_436);
nor U2419 (N_2419,In_1900,In_456);
nand U2420 (N_2420,In_376,In_886);
and U2421 (N_2421,In_2316,In_611);
and U2422 (N_2422,In_2251,In_502);
nand U2423 (N_2423,In_543,In_1159);
nand U2424 (N_2424,In_2274,In_897);
nand U2425 (N_2425,In_1946,In_1342);
nand U2426 (N_2426,In_2204,In_1337);
xnor U2427 (N_2427,In_953,In_1710);
or U2428 (N_2428,In_2107,In_2377);
xor U2429 (N_2429,In_1911,In_1998);
xnor U2430 (N_2430,In_2458,In_75);
and U2431 (N_2431,In_1861,In_413);
and U2432 (N_2432,In_1856,In_2192);
xnor U2433 (N_2433,In_251,In_1078);
nor U2434 (N_2434,In_1162,In_1419);
or U2435 (N_2435,In_2068,In_1871);
or U2436 (N_2436,In_1572,In_2041);
and U2437 (N_2437,In_704,In_146);
nand U2438 (N_2438,In_1997,In_1008);
nor U2439 (N_2439,In_2412,In_1808);
or U2440 (N_2440,In_1685,In_1120);
xnor U2441 (N_2441,In_105,In_316);
nand U2442 (N_2442,In_1660,In_730);
or U2443 (N_2443,In_784,In_626);
and U2444 (N_2444,In_0,In_476);
and U2445 (N_2445,In_1250,In_1028);
nand U2446 (N_2446,In_1170,In_1915);
nand U2447 (N_2447,In_149,In_1010);
nor U2448 (N_2448,In_353,In_1155);
nor U2449 (N_2449,In_2492,In_1651);
and U2450 (N_2450,In_2326,In_291);
or U2451 (N_2451,In_2382,In_852);
nand U2452 (N_2452,In_481,In_915);
nand U2453 (N_2453,In_1500,In_1588);
or U2454 (N_2454,In_707,In_1326);
nor U2455 (N_2455,In_45,In_743);
nand U2456 (N_2456,In_191,In_1171);
nor U2457 (N_2457,In_1712,In_727);
and U2458 (N_2458,In_1318,In_277);
nand U2459 (N_2459,In_1298,In_1037);
and U2460 (N_2460,In_1384,In_2025);
or U2461 (N_2461,In_1779,In_1892);
nand U2462 (N_2462,In_180,In_2316);
or U2463 (N_2463,In_1293,In_364);
nand U2464 (N_2464,In_1461,In_1079);
xnor U2465 (N_2465,In_804,In_549);
and U2466 (N_2466,In_2243,In_2005);
nand U2467 (N_2467,In_1110,In_2408);
nand U2468 (N_2468,In_2105,In_34);
xnor U2469 (N_2469,In_247,In_808);
xnor U2470 (N_2470,In_812,In_922);
or U2471 (N_2471,In_124,In_1076);
nor U2472 (N_2472,In_2144,In_144);
nand U2473 (N_2473,In_766,In_1928);
and U2474 (N_2474,In_2327,In_2021);
nand U2475 (N_2475,In_158,In_2096);
or U2476 (N_2476,In_1592,In_694);
nor U2477 (N_2477,In_489,In_1098);
or U2478 (N_2478,In_569,In_1673);
and U2479 (N_2479,In_1822,In_1140);
or U2480 (N_2480,In_1368,In_822);
nor U2481 (N_2481,In_161,In_522);
nor U2482 (N_2482,In_1899,In_1341);
xnor U2483 (N_2483,In_1611,In_1246);
or U2484 (N_2484,In_1874,In_1643);
nand U2485 (N_2485,In_1179,In_1758);
nand U2486 (N_2486,In_461,In_1325);
or U2487 (N_2487,In_780,In_474);
or U2488 (N_2488,In_1759,In_1615);
nor U2489 (N_2489,In_1508,In_829);
and U2490 (N_2490,In_663,In_796);
or U2491 (N_2491,In_507,In_1135);
nor U2492 (N_2492,In_1605,In_483);
and U2493 (N_2493,In_814,In_623);
or U2494 (N_2494,In_768,In_908);
and U2495 (N_2495,In_397,In_1606);
and U2496 (N_2496,In_1047,In_1476);
or U2497 (N_2497,In_143,In_217);
and U2498 (N_2498,In_486,In_1294);
nand U2499 (N_2499,In_690,In_1745);
nand U2500 (N_2500,In_832,In_2025);
nor U2501 (N_2501,In_2082,In_2451);
xor U2502 (N_2502,In_620,In_2068);
nor U2503 (N_2503,In_1144,In_1662);
nand U2504 (N_2504,In_518,In_1674);
and U2505 (N_2505,In_319,In_357);
nor U2506 (N_2506,In_2161,In_2437);
and U2507 (N_2507,In_2364,In_1712);
xnor U2508 (N_2508,In_1004,In_1501);
xor U2509 (N_2509,In_2362,In_1185);
xnor U2510 (N_2510,In_127,In_1156);
nor U2511 (N_2511,In_1873,In_570);
xnor U2512 (N_2512,In_1249,In_1671);
xor U2513 (N_2513,In_810,In_2088);
nand U2514 (N_2514,In_25,In_104);
nor U2515 (N_2515,In_858,In_1739);
nand U2516 (N_2516,In_222,In_1574);
nand U2517 (N_2517,In_2086,In_385);
xnor U2518 (N_2518,In_2238,In_843);
and U2519 (N_2519,In_1156,In_187);
xnor U2520 (N_2520,In_725,In_2053);
or U2521 (N_2521,In_113,In_93);
nor U2522 (N_2522,In_1196,In_1792);
nor U2523 (N_2523,In_729,In_1885);
nor U2524 (N_2524,In_251,In_1118);
xor U2525 (N_2525,In_2133,In_1623);
and U2526 (N_2526,In_909,In_1312);
xor U2527 (N_2527,In_426,In_2383);
or U2528 (N_2528,In_1094,In_1276);
and U2529 (N_2529,In_1714,In_1835);
and U2530 (N_2530,In_2226,In_370);
nand U2531 (N_2531,In_1634,In_846);
or U2532 (N_2532,In_1548,In_2470);
nor U2533 (N_2533,In_1254,In_2338);
xnor U2534 (N_2534,In_683,In_1128);
and U2535 (N_2535,In_1556,In_1290);
xor U2536 (N_2536,In_777,In_1402);
or U2537 (N_2537,In_2032,In_1929);
nor U2538 (N_2538,In_2184,In_2117);
nand U2539 (N_2539,In_571,In_998);
and U2540 (N_2540,In_1054,In_619);
nand U2541 (N_2541,In_2136,In_2391);
or U2542 (N_2542,In_2139,In_2195);
nand U2543 (N_2543,In_878,In_1810);
or U2544 (N_2544,In_1787,In_872);
nor U2545 (N_2545,In_959,In_1175);
nor U2546 (N_2546,In_2169,In_1305);
xor U2547 (N_2547,In_1474,In_1071);
and U2548 (N_2548,In_496,In_702);
nand U2549 (N_2549,In_1743,In_1824);
nor U2550 (N_2550,In_1128,In_209);
xnor U2551 (N_2551,In_678,In_176);
nor U2552 (N_2552,In_36,In_1166);
nor U2553 (N_2553,In_1703,In_702);
and U2554 (N_2554,In_510,In_306);
nand U2555 (N_2555,In_901,In_1421);
or U2556 (N_2556,In_183,In_1644);
nand U2557 (N_2557,In_452,In_1855);
nand U2558 (N_2558,In_462,In_1202);
or U2559 (N_2559,In_1366,In_267);
xnor U2560 (N_2560,In_1585,In_1233);
xor U2561 (N_2561,In_1972,In_134);
nor U2562 (N_2562,In_1978,In_689);
nand U2563 (N_2563,In_699,In_2010);
or U2564 (N_2564,In_2378,In_1606);
xor U2565 (N_2565,In_386,In_1798);
and U2566 (N_2566,In_501,In_635);
or U2567 (N_2567,In_1513,In_1186);
nand U2568 (N_2568,In_91,In_1031);
xnor U2569 (N_2569,In_2472,In_498);
or U2570 (N_2570,In_2056,In_574);
and U2571 (N_2571,In_1500,In_400);
or U2572 (N_2572,In_1108,In_2214);
nand U2573 (N_2573,In_1746,In_1384);
and U2574 (N_2574,In_2397,In_2105);
and U2575 (N_2575,In_1781,In_267);
nor U2576 (N_2576,In_1160,In_1715);
or U2577 (N_2577,In_799,In_2155);
nor U2578 (N_2578,In_1234,In_1928);
and U2579 (N_2579,In_2238,In_270);
nand U2580 (N_2580,In_672,In_287);
nand U2581 (N_2581,In_408,In_1360);
and U2582 (N_2582,In_122,In_1486);
nor U2583 (N_2583,In_2089,In_629);
nand U2584 (N_2584,In_1148,In_1992);
and U2585 (N_2585,In_1766,In_1710);
and U2586 (N_2586,In_1770,In_1206);
xnor U2587 (N_2587,In_462,In_1980);
and U2588 (N_2588,In_597,In_1351);
xnor U2589 (N_2589,In_1223,In_1218);
nand U2590 (N_2590,In_2318,In_480);
nor U2591 (N_2591,In_100,In_2422);
or U2592 (N_2592,In_1073,In_448);
and U2593 (N_2593,In_1677,In_1965);
or U2594 (N_2594,In_2171,In_541);
xor U2595 (N_2595,In_849,In_1917);
and U2596 (N_2596,In_205,In_1729);
nor U2597 (N_2597,In_1561,In_798);
and U2598 (N_2598,In_1176,In_2136);
or U2599 (N_2599,In_1573,In_1220);
xor U2600 (N_2600,In_78,In_1117);
or U2601 (N_2601,In_309,In_1058);
or U2602 (N_2602,In_2286,In_462);
nor U2603 (N_2603,In_527,In_1071);
nand U2604 (N_2604,In_636,In_2405);
and U2605 (N_2605,In_1427,In_2140);
nor U2606 (N_2606,In_1715,In_2477);
or U2607 (N_2607,In_2250,In_201);
nor U2608 (N_2608,In_382,In_1837);
and U2609 (N_2609,In_790,In_1965);
and U2610 (N_2610,In_2127,In_1398);
xor U2611 (N_2611,In_233,In_408);
nor U2612 (N_2612,In_453,In_2096);
or U2613 (N_2613,In_462,In_152);
or U2614 (N_2614,In_253,In_2305);
xnor U2615 (N_2615,In_1699,In_2222);
nor U2616 (N_2616,In_467,In_484);
xor U2617 (N_2617,In_191,In_561);
nor U2618 (N_2618,In_844,In_1328);
and U2619 (N_2619,In_776,In_2091);
and U2620 (N_2620,In_1676,In_529);
and U2621 (N_2621,In_29,In_686);
nand U2622 (N_2622,In_1306,In_1030);
nand U2623 (N_2623,In_154,In_2211);
and U2624 (N_2624,In_708,In_163);
nand U2625 (N_2625,In_148,In_120);
xor U2626 (N_2626,In_1380,In_1166);
nor U2627 (N_2627,In_1875,In_361);
or U2628 (N_2628,In_1863,In_1893);
nand U2629 (N_2629,In_1614,In_2315);
and U2630 (N_2630,In_1754,In_462);
nor U2631 (N_2631,In_54,In_1728);
and U2632 (N_2632,In_375,In_1352);
nor U2633 (N_2633,In_1802,In_2153);
and U2634 (N_2634,In_2398,In_870);
nor U2635 (N_2635,In_274,In_262);
xor U2636 (N_2636,In_1677,In_2430);
or U2637 (N_2637,In_2064,In_2093);
and U2638 (N_2638,In_1344,In_1587);
xnor U2639 (N_2639,In_536,In_111);
and U2640 (N_2640,In_45,In_1477);
nand U2641 (N_2641,In_122,In_1716);
and U2642 (N_2642,In_132,In_2335);
and U2643 (N_2643,In_1374,In_589);
xnor U2644 (N_2644,In_1829,In_426);
xnor U2645 (N_2645,In_357,In_946);
nand U2646 (N_2646,In_2255,In_442);
and U2647 (N_2647,In_543,In_2239);
nor U2648 (N_2648,In_186,In_2325);
nor U2649 (N_2649,In_385,In_1961);
nor U2650 (N_2650,In_2399,In_1513);
nor U2651 (N_2651,In_1956,In_1036);
nand U2652 (N_2652,In_1015,In_2485);
and U2653 (N_2653,In_1146,In_576);
xor U2654 (N_2654,In_1327,In_2433);
nand U2655 (N_2655,In_203,In_469);
nor U2656 (N_2656,In_1146,In_1505);
xor U2657 (N_2657,In_2202,In_1592);
nand U2658 (N_2658,In_2414,In_433);
nand U2659 (N_2659,In_136,In_726);
or U2660 (N_2660,In_1761,In_1887);
nand U2661 (N_2661,In_54,In_1206);
nand U2662 (N_2662,In_1761,In_2419);
nor U2663 (N_2663,In_1500,In_735);
xnor U2664 (N_2664,In_141,In_2473);
nand U2665 (N_2665,In_2421,In_502);
and U2666 (N_2666,In_264,In_302);
and U2667 (N_2667,In_1430,In_2400);
nor U2668 (N_2668,In_2368,In_1626);
nor U2669 (N_2669,In_72,In_2483);
xnor U2670 (N_2670,In_1798,In_427);
nand U2671 (N_2671,In_843,In_603);
xor U2672 (N_2672,In_1849,In_526);
xnor U2673 (N_2673,In_2316,In_1252);
and U2674 (N_2674,In_1513,In_197);
nand U2675 (N_2675,In_1780,In_771);
nor U2676 (N_2676,In_2048,In_90);
nand U2677 (N_2677,In_411,In_683);
or U2678 (N_2678,In_1335,In_179);
nand U2679 (N_2679,In_1862,In_191);
or U2680 (N_2680,In_209,In_1303);
nor U2681 (N_2681,In_618,In_1722);
xnor U2682 (N_2682,In_2187,In_1816);
nand U2683 (N_2683,In_1440,In_340);
and U2684 (N_2684,In_228,In_1808);
or U2685 (N_2685,In_1679,In_1903);
nand U2686 (N_2686,In_2402,In_1710);
and U2687 (N_2687,In_51,In_2488);
nor U2688 (N_2688,In_1004,In_855);
or U2689 (N_2689,In_2409,In_2346);
nor U2690 (N_2690,In_1621,In_1564);
nor U2691 (N_2691,In_891,In_1054);
xor U2692 (N_2692,In_2254,In_1777);
or U2693 (N_2693,In_2301,In_1865);
xor U2694 (N_2694,In_2361,In_171);
xor U2695 (N_2695,In_930,In_992);
nand U2696 (N_2696,In_1396,In_901);
nor U2697 (N_2697,In_864,In_1901);
and U2698 (N_2698,In_586,In_720);
nand U2699 (N_2699,In_1362,In_230);
and U2700 (N_2700,In_1274,In_2396);
nand U2701 (N_2701,In_2270,In_2050);
or U2702 (N_2702,In_1126,In_1731);
xnor U2703 (N_2703,In_1201,In_1683);
nand U2704 (N_2704,In_1514,In_2462);
or U2705 (N_2705,In_2062,In_452);
nand U2706 (N_2706,In_1603,In_323);
or U2707 (N_2707,In_593,In_661);
or U2708 (N_2708,In_876,In_671);
nand U2709 (N_2709,In_1053,In_1697);
nand U2710 (N_2710,In_1291,In_2025);
xor U2711 (N_2711,In_1974,In_1180);
nor U2712 (N_2712,In_1253,In_1315);
nor U2713 (N_2713,In_1189,In_1810);
and U2714 (N_2714,In_2374,In_525);
and U2715 (N_2715,In_1534,In_447);
or U2716 (N_2716,In_832,In_1217);
and U2717 (N_2717,In_1805,In_127);
or U2718 (N_2718,In_1948,In_50);
xnor U2719 (N_2719,In_870,In_1546);
nor U2720 (N_2720,In_852,In_2415);
nor U2721 (N_2721,In_416,In_2074);
and U2722 (N_2722,In_1845,In_660);
and U2723 (N_2723,In_10,In_613);
xor U2724 (N_2724,In_1255,In_1524);
or U2725 (N_2725,In_411,In_184);
xor U2726 (N_2726,In_320,In_1424);
or U2727 (N_2727,In_309,In_737);
nor U2728 (N_2728,In_638,In_2209);
nor U2729 (N_2729,In_174,In_1453);
nand U2730 (N_2730,In_259,In_516);
nand U2731 (N_2731,In_2425,In_1433);
or U2732 (N_2732,In_1211,In_272);
nor U2733 (N_2733,In_1595,In_597);
or U2734 (N_2734,In_441,In_1898);
xor U2735 (N_2735,In_351,In_1274);
xor U2736 (N_2736,In_698,In_318);
xnor U2737 (N_2737,In_2175,In_1267);
xnor U2738 (N_2738,In_1280,In_2225);
or U2739 (N_2739,In_1649,In_1052);
nand U2740 (N_2740,In_1561,In_236);
nand U2741 (N_2741,In_390,In_2165);
xnor U2742 (N_2742,In_2230,In_1930);
xnor U2743 (N_2743,In_608,In_1633);
nand U2744 (N_2744,In_889,In_2355);
nor U2745 (N_2745,In_316,In_1616);
nor U2746 (N_2746,In_572,In_715);
nand U2747 (N_2747,In_2054,In_203);
nand U2748 (N_2748,In_1230,In_1428);
nand U2749 (N_2749,In_1627,In_621);
nand U2750 (N_2750,In_2400,In_68);
xnor U2751 (N_2751,In_2092,In_1847);
nor U2752 (N_2752,In_592,In_1544);
nor U2753 (N_2753,In_602,In_1082);
and U2754 (N_2754,In_2011,In_445);
nand U2755 (N_2755,In_1152,In_2273);
nor U2756 (N_2756,In_1588,In_2093);
nor U2757 (N_2757,In_1759,In_276);
nor U2758 (N_2758,In_243,In_1864);
nand U2759 (N_2759,In_2126,In_797);
nor U2760 (N_2760,In_472,In_245);
and U2761 (N_2761,In_1868,In_1552);
and U2762 (N_2762,In_2412,In_367);
xnor U2763 (N_2763,In_1017,In_1770);
xnor U2764 (N_2764,In_1387,In_2001);
nor U2765 (N_2765,In_242,In_1950);
nor U2766 (N_2766,In_547,In_2286);
nand U2767 (N_2767,In_1117,In_386);
or U2768 (N_2768,In_925,In_530);
nor U2769 (N_2769,In_791,In_1403);
and U2770 (N_2770,In_852,In_1809);
nor U2771 (N_2771,In_1891,In_1169);
nand U2772 (N_2772,In_1093,In_1956);
xnor U2773 (N_2773,In_2082,In_1925);
nand U2774 (N_2774,In_661,In_1914);
xor U2775 (N_2775,In_381,In_1769);
nor U2776 (N_2776,In_616,In_790);
and U2777 (N_2777,In_2118,In_237);
and U2778 (N_2778,In_1587,In_1581);
xor U2779 (N_2779,In_2029,In_2331);
or U2780 (N_2780,In_1253,In_296);
nor U2781 (N_2781,In_1311,In_1652);
or U2782 (N_2782,In_417,In_1564);
xor U2783 (N_2783,In_1595,In_1024);
or U2784 (N_2784,In_556,In_2001);
xor U2785 (N_2785,In_1731,In_146);
or U2786 (N_2786,In_78,In_2448);
nand U2787 (N_2787,In_350,In_277);
xnor U2788 (N_2788,In_592,In_1317);
and U2789 (N_2789,In_1898,In_838);
xor U2790 (N_2790,In_2274,In_1789);
nor U2791 (N_2791,In_1981,In_1047);
nor U2792 (N_2792,In_159,In_665);
xor U2793 (N_2793,In_1067,In_1347);
and U2794 (N_2794,In_1939,In_1215);
xor U2795 (N_2795,In_2241,In_2268);
nor U2796 (N_2796,In_2022,In_267);
nor U2797 (N_2797,In_2281,In_681);
nor U2798 (N_2798,In_36,In_2402);
or U2799 (N_2799,In_1457,In_355);
nand U2800 (N_2800,In_2294,In_1222);
nand U2801 (N_2801,In_1130,In_1406);
or U2802 (N_2802,In_378,In_832);
and U2803 (N_2803,In_2120,In_2047);
and U2804 (N_2804,In_1335,In_1092);
xnor U2805 (N_2805,In_2398,In_1500);
and U2806 (N_2806,In_1804,In_1581);
nand U2807 (N_2807,In_528,In_1430);
or U2808 (N_2808,In_1305,In_2441);
xnor U2809 (N_2809,In_105,In_2373);
nor U2810 (N_2810,In_290,In_2110);
nor U2811 (N_2811,In_1206,In_51);
nor U2812 (N_2812,In_32,In_156);
and U2813 (N_2813,In_1403,In_2103);
xor U2814 (N_2814,In_2088,In_1927);
xnor U2815 (N_2815,In_2274,In_2280);
xor U2816 (N_2816,In_1921,In_38);
and U2817 (N_2817,In_154,In_2432);
and U2818 (N_2818,In_2178,In_2426);
or U2819 (N_2819,In_1007,In_1349);
nand U2820 (N_2820,In_1839,In_1428);
nand U2821 (N_2821,In_812,In_9);
nand U2822 (N_2822,In_1969,In_197);
or U2823 (N_2823,In_2438,In_449);
and U2824 (N_2824,In_1044,In_2365);
xnor U2825 (N_2825,In_1431,In_892);
and U2826 (N_2826,In_1430,In_2021);
xnor U2827 (N_2827,In_1838,In_26);
nand U2828 (N_2828,In_641,In_223);
or U2829 (N_2829,In_697,In_76);
nand U2830 (N_2830,In_1465,In_1336);
xnor U2831 (N_2831,In_789,In_1087);
nor U2832 (N_2832,In_1062,In_1308);
nor U2833 (N_2833,In_877,In_1294);
nand U2834 (N_2834,In_2213,In_431);
or U2835 (N_2835,In_1955,In_1317);
and U2836 (N_2836,In_368,In_478);
nand U2837 (N_2837,In_1136,In_1463);
xnor U2838 (N_2838,In_2005,In_964);
nand U2839 (N_2839,In_1579,In_2425);
and U2840 (N_2840,In_1890,In_643);
or U2841 (N_2841,In_1607,In_988);
or U2842 (N_2842,In_554,In_189);
and U2843 (N_2843,In_1228,In_2038);
nor U2844 (N_2844,In_222,In_858);
or U2845 (N_2845,In_353,In_423);
xor U2846 (N_2846,In_542,In_282);
or U2847 (N_2847,In_1645,In_613);
xor U2848 (N_2848,In_1722,In_2376);
or U2849 (N_2849,In_848,In_545);
xor U2850 (N_2850,In_1514,In_288);
or U2851 (N_2851,In_104,In_366);
and U2852 (N_2852,In_2498,In_939);
xor U2853 (N_2853,In_2262,In_1202);
nand U2854 (N_2854,In_1001,In_695);
xor U2855 (N_2855,In_2092,In_1675);
nor U2856 (N_2856,In_898,In_1023);
xnor U2857 (N_2857,In_239,In_891);
and U2858 (N_2858,In_1874,In_1130);
nor U2859 (N_2859,In_2458,In_799);
or U2860 (N_2860,In_2403,In_1824);
xor U2861 (N_2861,In_90,In_656);
nand U2862 (N_2862,In_1934,In_1227);
and U2863 (N_2863,In_12,In_202);
and U2864 (N_2864,In_2221,In_1244);
xnor U2865 (N_2865,In_1777,In_1075);
nor U2866 (N_2866,In_1715,In_1679);
and U2867 (N_2867,In_2230,In_2465);
nor U2868 (N_2868,In_1167,In_1519);
nand U2869 (N_2869,In_1403,In_1475);
or U2870 (N_2870,In_2428,In_1295);
nand U2871 (N_2871,In_1645,In_219);
or U2872 (N_2872,In_1957,In_2146);
and U2873 (N_2873,In_2493,In_723);
or U2874 (N_2874,In_2071,In_2349);
or U2875 (N_2875,In_264,In_18);
nor U2876 (N_2876,In_1450,In_1046);
nand U2877 (N_2877,In_1985,In_774);
and U2878 (N_2878,In_1095,In_1867);
or U2879 (N_2879,In_491,In_980);
or U2880 (N_2880,In_1780,In_772);
nor U2881 (N_2881,In_330,In_147);
or U2882 (N_2882,In_1887,In_675);
xnor U2883 (N_2883,In_1817,In_195);
nand U2884 (N_2884,In_1437,In_2098);
nor U2885 (N_2885,In_2244,In_2120);
nand U2886 (N_2886,In_2192,In_523);
nand U2887 (N_2887,In_1537,In_85);
or U2888 (N_2888,In_1897,In_2328);
or U2889 (N_2889,In_150,In_1605);
nand U2890 (N_2890,In_2209,In_1861);
nor U2891 (N_2891,In_61,In_928);
or U2892 (N_2892,In_1109,In_1913);
xnor U2893 (N_2893,In_53,In_2347);
or U2894 (N_2894,In_2250,In_1210);
nor U2895 (N_2895,In_811,In_589);
nand U2896 (N_2896,In_1990,In_1815);
or U2897 (N_2897,In_1495,In_525);
nand U2898 (N_2898,In_1205,In_1704);
nor U2899 (N_2899,In_672,In_2469);
and U2900 (N_2900,In_1203,In_227);
nor U2901 (N_2901,In_1750,In_2448);
nand U2902 (N_2902,In_2435,In_598);
or U2903 (N_2903,In_1208,In_2178);
xnor U2904 (N_2904,In_1348,In_1468);
nor U2905 (N_2905,In_241,In_2288);
xnor U2906 (N_2906,In_1980,In_2011);
nor U2907 (N_2907,In_192,In_2175);
nand U2908 (N_2908,In_324,In_1519);
nand U2909 (N_2909,In_431,In_1308);
nor U2910 (N_2910,In_1260,In_819);
or U2911 (N_2911,In_2388,In_1158);
nand U2912 (N_2912,In_2452,In_2119);
xnor U2913 (N_2913,In_2268,In_1663);
xor U2914 (N_2914,In_986,In_1083);
nand U2915 (N_2915,In_1852,In_354);
xnor U2916 (N_2916,In_1841,In_1106);
xnor U2917 (N_2917,In_1171,In_1162);
nand U2918 (N_2918,In_860,In_1366);
nor U2919 (N_2919,In_1176,In_982);
and U2920 (N_2920,In_1630,In_2198);
nor U2921 (N_2921,In_758,In_415);
and U2922 (N_2922,In_2262,In_95);
or U2923 (N_2923,In_2102,In_1386);
xnor U2924 (N_2924,In_2020,In_1478);
and U2925 (N_2925,In_1891,In_1667);
xnor U2926 (N_2926,In_1336,In_2361);
nor U2927 (N_2927,In_1259,In_216);
xor U2928 (N_2928,In_1912,In_1951);
xor U2929 (N_2929,In_1975,In_922);
nand U2930 (N_2930,In_756,In_426);
nor U2931 (N_2931,In_350,In_1476);
and U2932 (N_2932,In_321,In_1995);
xnor U2933 (N_2933,In_1318,In_2145);
xnor U2934 (N_2934,In_512,In_1572);
xor U2935 (N_2935,In_2232,In_2068);
nor U2936 (N_2936,In_1299,In_1484);
nand U2937 (N_2937,In_1748,In_2226);
and U2938 (N_2938,In_587,In_2076);
xnor U2939 (N_2939,In_1138,In_1494);
or U2940 (N_2940,In_89,In_1324);
xnor U2941 (N_2941,In_1655,In_2345);
and U2942 (N_2942,In_2167,In_564);
nand U2943 (N_2943,In_2041,In_767);
xnor U2944 (N_2944,In_2153,In_225);
nand U2945 (N_2945,In_1373,In_1471);
and U2946 (N_2946,In_2467,In_564);
and U2947 (N_2947,In_1463,In_714);
xor U2948 (N_2948,In_2120,In_1600);
nor U2949 (N_2949,In_1519,In_37);
nor U2950 (N_2950,In_1682,In_2286);
nor U2951 (N_2951,In_793,In_1198);
nor U2952 (N_2952,In_945,In_2133);
or U2953 (N_2953,In_211,In_2130);
or U2954 (N_2954,In_1530,In_522);
nand U2955 (N_2955,In_55,In_633);
nand U2956 (N_2956,In_1049,In_1458);
nand U2957 (N_2957,In_1728,In_1524);
xnor U2958 (N_2958,In_2204,In_615);
and U2959 (N_2959,In_1998,In_525);
xnor U2960 (N_2960,In_699,In_925);
or U2961 (N_2961,In_1387,In_912);
xnor U2962 (N_2962,In_210,In_2034);
xnor U2963 (N_2963,In_2223,In_885);
and U2964 (N_2964,In_576,In_1556);
and U2965 (N_2965,In_103,In_1231);
nand U2966 (N_2966,In_515,In_504);
nor U2967 (N_2967,In_793,In_2426);
nand U2968 (N_2968,In_1961,In_32);
nand U2969 (N_2969,In_83,In_1399);
or U2970 (N_2970,In_2155,In_2239);
nor U2971 (N_2971,In_1444,In_235);
nand U2972 (N_2972,In_519,In_1647);
nand U2973 (N_2973,In_549,In_2110);
nand U2974 (N_2974,In_660,In_1185);
or U2975 (N_2975,In_1735,In_1660);
or U2976 (N_2976,In_1854,In_1547);
or U2977 (N_2977,In_1953,In_736);
nand U2978 (N_2978,In_708,In_814);
nand U2979 (N_2979,In_2422,In_643);
xor U2980 (N_2980,In_1042,In_288);
or U2981 (N_2981,In_401,In_948);
or U2982 (N_2982,In_2185,In_1454);
xor U2983 (N_2983,In_63,In_2280);
or U2984 (N_2984,In_1138,In_1029);
or U2985 (N_2985,In_1940,In_31);
or U2986 (N_2986,In_981,In_662);
xnor U2987 (N_2987,In_1015,In_2125);
or U2988 (N_2988,In_2076,In_1266);
nand U2989 (N_2989,In_1896,In_1699);
and U2990 (N_2990,In_897,In_992);
or U2991 (N_2991,In_446,In_1847);
nor U2992 (N_2992,In_334,In_2437);
nand U2993 (N_2993,In_801,In_661);
nand U2994 (N_2994,In_931,In_1221);
and U2995 (N_2995,In_2101,In_1416);
xor U2996 (N_2996,In_1879,In_2254);
xor U2997 (N_2997,In_1269,In_1066);
nor U2998 (N_2998,In_936,In_1312);
nand U2999 (N_2999,In_1224,In_2347);
xnor U3000 (N_3000,In_1595,In_1927);
or U3001 (N_3001,In_2304,In_833);
and U3002 (N_3002,In_2091,In_1907);
and U3003 (N_3003,In_478,In_1835);
nand U3004 (N_3004,In_2229,In_781);
and U3005 (N_3005,In_548,In_1953);
nand U3006 (N_3006,In_415,In_2084);
or U3007 (N_3007,In_778,In_1199);
nor U3008 (N_3008,In_1227,In_215);
and U3009 (N_3009,In_411,In_953);
nor U3010 (N_3010,In_154,In_768);
xor U3011 (N_3011,In_1118,In_2020);
or U3012 (N_3012,In_2479,In_640);
and U3013 (N_3013,In_2141,In_2070);
or U3014 (N_3014,In_457,In_343);
and U3015 (N_3015,In_2270,In_622);
or U3016 (N_3016,In_97,In_1568);
nand U3017 (N_3017,In_1088,In_2297);
and U3018 (N_3018,In_1255,In_1404);
nand U3019 (N_3019,In_1114,In_2111);
nor U3020 (N_3020,In_831,In_1687);
nand U3021 (N_3021,In_2066,In_709);
and U3022 (N_3022,In_1040,In_2416);
nand U3023 (N_3023,In_1573,In_563);
xnor U3024 (N_3024,In_1131,In_2338);
and U3025 (N_3025,In_689,In_785);
or U3026 (N_3026,In_581,In_885);
nand U3027 (N_3027,In_2333,In_585);
xor U3028 (N_3028,In_129,In_1283);
xor U3029 (N_3029,In_1757,In_988);
xnor U3030 (N_3030,In_1791,In_1627);
xnor U3031 (N_3031,In_1160,In_1865);
xnor U3032 (N_3032,In_2496,In_1440);
nand U3033 (N_3033,In_754,In_1507);
xnor U3034 (N_3034,In_2063,In_2044);
nand U3035 (N_3035,In_168,In_2265);
and U3036 (N_3036,In_877,In_1415);
xnor U3037 (N_3037,In_1754,In_2317);
nor U3038 (N_3038,In_1999,In_1521);
nor U3039 (N_3039,In_908,In_721);
nand U3040 (N_3040,In_727,In_2216);
and U3041 (N_3041,In_1475,In_1940);
and U3042 (N_3042,In_268,In_2214);
nand U3043 (N_3043,In_1009,In_1361);
nor U3044 (N_3044,In_53,In_240);
nand U3045 (N_3045,In_122,In_1239);
and U3046 (N_3046,In_1132,In_1541);
nand U3047 (N_3047,In_1506,In_1809);
nand U3048 (N_3048,In_2224,In_1335);
nor U3049 (N_3049,In_1332,In_1041);
nor U3050 (N_3050,In_560,In_628);
nand U3051 (N_3051,In_225,In_1950);
nor U3052 (N_3052,In_779,In_1466);
and U3053 (N_3053,In_871,In_2338);
nor U3054 (N_3054,In_1273,In_226);
xor U3055 (N_3055,In_1339,In_255);
or U3056 (N_3056,In_2320,In_2151);
nor U3057 (N_3057,In_1298,In_2191);
and U3058 (N_3058,In_594,In_1125);
nor U3059 (N_3059,In_82,In_100);
or U3060 (N_3060,In_1588,In_57);
nand U3061 (N_3061,In_1350,In_453);
nand U3062 (N_3062,In_1114,In_1147);
xor U3063 (N_3063,In_1664,In_835);
and U3064 (N_3064,In_23,In_1536);
nand U3065 (N_3065,In_848,In_1595);
and U3066 (N_3066,In_687,In_828);
nand U3067 (N_3067,In_388,In_299);
nor U3068 (N_3068,In_451,In_196);
xnor U3069 (N_3069,In_2149,In_2004);
nand U3070 (N_3070,In_857,In_1658);
nand U3071 (N_3071,In_1450,In_772);
xnor U3072 (N_3072,In_1692,In_1955);
or U3073 (N_3073,In_971,In_1205);
xnor U3074 (N_3074,In_508,In_2382);
and U3075 (N_3075,In_67,In_117);
nand U3076 (N_3076,In_1702,In_1802);
or U3077 (N_3077,In_1416,In_1816);
xor U3078 (N_3078,In_632,In_2191);
and U3079 (N_3079,In_447,In_2269);
nor U3080 (N_3080,In_710,In_2084);
and U3081 (N_3081,In_1526,In_1963);
xor U3082 (N_3082,In_1085,In_105);
and U3083 (N_3083,In_925,In_630);
and U3084 (N_3084,In_1705,In_2249);
nor U3085 (N_3085,In_1597,In_1018);
nand U3086 (N_3086,In_1223,In_840);
or U3087 (N_3087,In_1046,In_839);
nor U3088 (N_3088,In_1460,In_462);
nand U3089 (N_3089,In_636,In_1432);
xor U3090 (N_3090,In_1867,In_427);
nor U3091 (N_3091,In_2381,In_10);
xnor U3092 (N_3092,In_1734,In_316);
and U3093 (N_3093,In_1041,In_1541);
or U3094 (N_3094,In_1445,In_673);
nor U3095 (N_3095,In_1207,In_1279);
nor U3096 (N_3096,In_118,In_127);
nand U3097 (N_3097,In_1954,In_1403);
or U3098 (N_3098,In_84,In_146);
xor U3099 (N_3099,In_773,In_1286);
xor U3100 (N_3100,In_2433,In_265);
xnor U3101 (N_3101,In_623,In_2206);
nor U3102 (N_3102,In_1919,In_1735);
or U3103 (N_3103,In_1083,In_21);
or U3104 (N_3104,In_399,In_768);
and U3105 (N_3105,In_2415,In_1177);
and U3106 (N_3106,In_2485,In_1490);
nand U3107 (N_3107,In_1263,In_2085);
and U3108 (N_3108,In_2031,In_260);
xor U3109 (N_3109,In_1835,In_856);
nand U3110 (N_3110,In_1497,In_148);
and U3111 (N_3111,In_813,In_2319);
xnor U3112 (N_3112,In_2085,In_1404);
xor U3113 (N_3113,In_2372,In_1256);
and U3114 (N_3114,In_2326,In_1397);
and U3115 (N_3115,In_239,In_1087);
and U3116 (N_3116,In_1839,In_2433);
nand U3117 (N_3117,In_1912,In_60);
nand U3118 (N_3118,In_1801,In_1939);
xor U3119 (N_3119,In_10,In_2372);
and U3120 (N_3120,In_1828,In_1542);
and U3121 (N_3121,In_196,In_1417);
or U3122 (N_3122,In_1458,In_1595);
nor U3123 (N_3123,In_492,In_808);
nand U3124 (N_3124,In_1344,In_330);
nor U3125 (N_3125,N_2033,N_1013);
and U3126 (N_3126,N_2061,N_2665);
nor U3127 (N_3127,N_1525,N_1511);
nor U3128 (N_3128,N_1022,N_2511);
xnor U3129 (N_3129,N_826,N_2763);
nor U3130 (N_3130,N_2747,N_1236);
nand U3131 (N_3131,N_730,N_2266);
nor U3132 (N_3132,N_805,N_848);
xnor U3133 (N_3133,N_450,N_1614);
or U3134 (N_3134,N_3068,N_2437);
nand U3135 (N_3135,N_1556,N_2406);
xor U3136 (N_3136,N_471,N_396);
xnor U3137 (N_3137,N_1093,N_2713);
nand U3138 (N_3138,N_598,N_1935);
nor U3139 (N_3139,N_2753,N_806);
and U3140 (N_3140,N_892,N_376);
or U3141 (N_3141,N_223,N_2557);
and U3142 (N_3142,N_1131,N_2021);
xor U3143 (N_3143,N_1851,N_1517);
xnor U3144 (N_3144,N_350,N_1967);
xnor U3145 (N_3145,N_1626,N_1750);
or U3146 (N_3146,N_1086,N_2923);
xor U3147 (N_3147,N_868,N_1780);
nand U3148 (N_3148,N_365,N_2931);
nor U3149 (N_3149,N_1520,N_2322);
xor U3150 (N_3150,N_2653,N_1095);
nor U3151 (N_3151,N_1049,N_1152);
nand U3152 (N_3152,N_1716,N_1384);
nor U3153 (N_3153,N_1515,N_372);
nand U3154 (N_3154,N_1749,N_225);
xnor U3155 (N_3155,N_171,N_3043);
nand U3156 (N_3156,N_3053,N_1690);
nor U3157 (N_3157,N_1184,N_26);
or U3158 (N_3158,N_2843,N_2860);
or U3159 (N_3159,N_2586,N_2217);
and U3160 (N_3160,N_1121,N_2508);
or U3161 (N_3161,N_1688,N_525);
nor U3162 (N_3162,N_2925,N_2764);
or U3163 (N_3163,N_2244,N_2034);
nor U3164 (N_3164,N_832,N_2769);
xor U3165 (N_3165,N_2131,N_1718);
or U3166 (N_3166,N_2699,N_10);
and U3167 (N_3167,N_668,N_883);
nand U3168 (N_3168,N_3022,N_722);
nor U3169 (N_3169,N_1312,N_1113);
and U3170 (N_3170,N_1106,N_2646);
and U3171 (N_3171,N_205,N_763);
nor U3172 (N_3172,N_2195,N_3001);
and U3173 (N_3173,N_2041,N_775);
xnor U3174 (N_3174,N_1559,N_1466);
nand U3175 (N_3175,N_198,N_2527);
and U3176 (N_3176,N_2086,N_418);
and U3177 (N_3177,N_857,N_229);
nor U3178 (N_3178,N_2804,N_2569);
nand U3179 (N_3179,N_1276,N_1392);
xor U3180 (N_3180,N_329,N_125);
and U3181 (N_3181,N_403,N_2015);
nor U3182 (N_3182,N_1205,N_801);
nand U3183 (N_3183,N_628,N_264);
nor U3184 (N_3184,N_603,N_687);
nor U3185 (N_3185,N_1543,N_2615);
xor U3186 (N_3186,N_2016,N_1292);
and U3187 (N_3187,N_273,N_1732);
and U3188 (N_3188,N_2897,N_3077);
nor U3189 (N_3189,N_1598,N_924);
nor U3190 (N_3190,N_191,N_1344);
xnor U3191 (N_3191,N_130,N_1270);
or U3192 (N_3192,N_633,N_2855);
or U3193 (N_3193,N_1711,N_1553);
nand U3194 (N_3194,N_2844,N_2497);
xor U3195 (N_3195,N_1035,N_2768);
or U3196 (N_3196,N_1783,N_246);
nor U3197 (N_3197,N_1209,N_2515);
nand U3198 (N_3198,N_2255,N_1786);
xor U3199 (N_3199,N_1720,N_511);
nor U3200 (N_3200,N_2666,N_908);
or U3201 (N_3201,N_944,N_2649);
or U3202 (N_3202,N_2474,N_2120);
nor U3203 (N_3203,N_2671,N_2473);
or U3204 (N_3204,N_48,N_375);
nor U3205 (N_3205,N_440,N_1029);
and U3206 (N_3206,N_2270,N_1074);
xor U3207 (N_3207,N_2353,N_677);
nand U3208 (N_3208,N_2701,N_254);
nor U3209 (N_3209,N_1552,N_1172);
nand U3210 (N_3210,N_2415,N_662);
and U3211 (N_3211,N_2959,N_1162);
nor U3212 (N_3212,N_946,N_720);
xnor U3213 (N_3213,N_240,N_1171);
or U3214 (N_3214,N_255,N_2992);
nand U3215 (N_3215,N_887,N_1341);
nand U3216 (N_3216,N_1643,N_2731);
nand U3217 (N_3217,N_129,N_45);
and U3218 (N_3218,N_2096,N_599);
xor U3219 (N_3219,N_955,N_88);
nor U3220 (N_3220,N_371,N_3070);
nand U3221 (N_3221,N_2155,N_1413);
and U3222 (N_3222,N_2674,N_190);
or U3223 (N_3223,N_425,N_2501);
and U3224 (N_3224,N_1289,N_1141);
and U3225 (N_3225,N_1275,N_1211);
and U3226 (N_3226,N_2981,N_1377);
xor U3227 (N_3227,N_2877,N_299);
or U3228 (N_3228,N_1400,N_2933);
nand U3229 (N_3229,N_204,N_2519);
or U3230 (N_3230,N_127,N_2012);
or U3231 (N_3231,N_520,N_701);
or U3232 (N_3232,N_684,N_2572);
nand U3233 (N_3233,N_2559,N_1260);
xnor U3234 (N_3234,N_920,N_1134);
nor U3235 (N_3235,N_1539,N_1862);
nor U3236 (N_3236,N_2737,N_1503);
and U3237 (N_3237,N_517,N_2551);
or U3238 (N_3238,N_1507,N_2281);
or U3239 (N_3239,N_302,N_636);
nand U3240 (N_3240,N_776,N_2370);
or U3241 (N_3241,N_608,N_2967);
or U3242 (N_3242,N_2889,N_2818);
xnor U3243 (N_3243,N_550,N_1871);
or U3244 (N_3244,N_623,N_1118);
and U3245 (N_3245,N_998,N_2004);
xor U3246 (N_3246,N_723,N_2469);
nand U3247 (N_3247,N_1941,N_2374);
and U3248 (N_3248,N_747,N_1537);
or U3249 (N_3249,N_1476,N_1789);
xor U3250 (N_3250,N_2640,N_556);
or U3251 (N_3251,N_2518,N_2529);
and U3252 (N_3252,N_359,N_117);
or U3253 (N_3253,N_1526,N_1970);
or U3254 (N_3254,N_2715,N_1482);
or U3255 (N_3255,N_2777,N_354);
nor U3256 (N_3256,N_1811,N_1165);
xnor U3257 (N_3257,N_854,N_2725);
xor U3258 (N_3258,N_962,N_781);
and U3259 (N_3259,N_1681,N_1226);
and U3260 (N_3260,N_1046,N_2611);
and U3261 (N_3261,N_3123,N_2320);
nand U3262 (N_3262,N_3012,N_1306);
xnor U3263 (N_3263,N_1683,N_670);
nor U3264 (N_3264,N_1194,N_1560);
nand U3265 (N_3265,N_577,N_2929);
nor U3266 (N_3266,N_2533,N_1446);
nor U3267 (N_3267,N_1833,N_2790);
or U3268 (N_3268,N_1168,N_3023);
and U3269 (N_3269,N_700,N_1300);
nor U3270 (N_3270,N_1792,N_1521);
xnor U3271 (N_3271,N_164,N_2341);
xnor U3272 (N_3272,N_1704,N_2150);
and U3273 (N_3273,N_1529,N_1747);
or U3274 (N_3274,N_67,N_2346);
nor U3275 (N_3275,N_706,N_2347);
nor U3276 (N_3276,N_2687,N_1338);
nor U3277 (N_3277,N_332,N_338);
nand U3278 (N_3278,N_218,N_767);
nand U3279 (N_3279,N_2328,N_2167);
nand U3280 (N_3280,N_289,N_2812);
nor U3281 (N_3281,N_1116,N_347);
xor U3282 (N_3282,N_2007,N_2607);
nand U3283 (N_3283,N_3014,N_2118);
nor U3284 (N_3284,N_1942,N_966);
nand U3285 (N_3285,N_2418,N_2040);
nor U3286 (N_3286,N_957,N_2896);
xnor U3287 (N_3287,N_1990,N_2985);
and U3288 (N_3288,N_37,N_2813);
nor U3289 (N_3289,N_2214,N_2090);
xor U3290 (N_3290,N_705,N_1557);
nand U3291 (N_3291,N_953,N_2207);
xnor U3292 (N_3292,N_2265,N_1848);
nor U3293 (N_3293,N_1272,N_1702);
nand U3294 (N_3294,N_2165,N_1650);
nor U3295 (N_3295,N_2471,N_241);
and U3296 (N_3296,N_1000,N_1047);
or U3297 (N_3297,N_2956,N_1354);
and U3298 (N_3298,N_1422,N_2539);
or U3299 (N_3299,N_206,N_2754);
and U3300 (N_3300,N_708,N_2302);
nand U3301 (N_3301,N_1411,N_1769);
nor U3302 (N_3302,N_2157,N_2606);
nand U3303 (N_3303,N_116,N_33);
or U3304 (N_3304,N_2655,N_2290);
nor U3305 (N_3305,N_385,N_2957);
and U3306 (N_3306,N_1613,N_2130);
or U3307 (N_3307,N_2888,N_1889);
xnor U3308 (N_3308,N_1902,N_1578);
xnor U3309 (N_3309,N_1549,N_138);
and U3310 (N_3310,N_3028,N_180);
xnor U3311 (N_3311,N_968,N_3118);
nand U3312 (N_3312,N_843,N_1555);
nand U3313 (N_3313,N_2367,N_2476);
nand U3314 (N_3314,N_1495,N_856);
and U3315 (N_3315,N_2111,N_136);
and U3316 (N_3316,N_1691,N_569);
or U3317 (N_3317,N_1577,N_894);
nor U3318 (N_3318,N_147,N_2898);
or U3319 (N_3319,N_934,N_1264);
and U3320 (N_3320,N_2548,N_2078);
or U3321 (N_3321,N_2512,N_1137);
or U3322 (N_3322,N_2117,N_31);
or U3323 (N_3323,N_1542,N_2354);
nand U3324 (N_3324,N_2387,N_1887);
or U3325 (N_3325,N_1831,N_211);
xnor U3326 (N_3326,N_459,N_1877);
and U3327 (N_3327,N_1311,N_1310);
xor U3328 (N_3328,N_2991,N_3092);
nor U3329 (N_3329,N_2892,N_3031);
xor U3330 (N_3330,N_1208,N_2462);
nand U3331 (N_3331,N_2261,N_1016);
and U3332 (N_3332,N_1096,N_1498);
and U3333 (N_3333,N_552,N_159);
and U3334 (N_3334,N_551,N_483);
nand U3335 (N_3335,N_793,N_2383);
or U3336 (N_3336,N_247,N_2988);
nand U3337 (N_3337,N_1320,N_2802);
or U3338 (N_3338,N_1684,N_2884);
and U3339 (N_3339,N_792,N_2116);
xor U3340 (N_3340,N_3105,N_1661);
nor U3341 (N_3341,N_852,N_1977);
and U3342 (N_3342,N_395,N_1269);
nor U3343 (N_3343,N_1144,N_1605);
xnor U3344 (N_3344,N_527,N_72);
nor U3345 (N_3345,N_1087,N_1782);
and U3346 (N_3346,N_3062,N_769);
nor U3347 (N_3347,N_1174,N_2407);
or U3348 (N_3348,N_678,N_2576);
xor U3349 (N_3349,N_1898,N_213);
or U3350 (N_3350,N_2570,N_2102);
or U3351 (N_3351,N_2596,N_2202);
nor U3352 (N_3352,N_1535,N_847);
xor U3353 (N_3353,N_1706,N_1908);
nand U3354 (N_3354,N_658,N_2759);
xnor U3355 (N_3355,N_461,N_3084);
or U3356 (N_3356,N_2068,N_3027);
nand U3357 (N_3357,N_992,N_1781);
or U3358 (N_3358,N_1623,N_2975);
nor U3359 (N_3359,N_1389,N_2592);
xor U3360 (N_3360,N_2736,N_1216);
and U3361 (N_3361,N_671,N_1234);
or U3362 (N_3362,N_1123,N_497);
and U3363 (N_3363,N_518,N_726);
and U3364 (N_3364,N_581,N_1301);
nor U3365 (N_3365,N_493,N_2986);
xnor U3366 (N_3366,N_1610,N_745);
nand U3367 (N_3367,N_2779,N_3114);
xnor U3368 (N_3368,N_2093,N_782);
and U3369 (N_3369,N_1998,N_1985);
nor U3370 (N_3370,N_975,N_1630);
and U3371 (N_3371,N_224,N_1659);
nand U3372 (N_3372,N_736,N_1745);
or U3373 (N_3373,N_914,N_195);
and U3374 (N_3374,N_1945,N_2463);
or U3375 (N_3375,N_73,N_2184);
or U3376 (N_3376,N_2216,N_2796);
and U3377 (N_3377,N_2807,N_269);
or U3378 (N_3378,N_2075,N_521);
nand U3379 (N_3379,N_2751,N_280);
and U3380 (N_3380,N_1426,N_2932);
nand U3381 (N_3381,N_1464,N_135);
nor U3382 (N_3382,N_2386,N_2417);
xor U3383 (N_3383,N_1654,N_484);
nand U3384 (N_3384,N_2242,N_653);
nor U3385 (N_3385,N_77,N_566);
nand U3386 (N_3386,N_2791,N_1401);
nor U3387 (N_3387,N_2561,N_785);
nand U3388 (N_3388,N_988,N_896);
and U3389 (N_3389,N_999,N_1081);
nor U3390 (N_3390,N_2361,N_2404);
or U3391 (N_3391,N_93,N_2679);
or U3392 (N_3392,N_1425,N_2924);
and U3393 (N_3393,N_2849,N_1759);
nor U3394 (N_3394,N_1816,N_2708);
nor U3395 (N_3395,N_2050,N_1891);
xor U3396 (N_3396,N_833,N_336);
and U3397 (N_3397,N_1380,N_2369);
xor U3398 (N_3398,N_1304,N_1996);
xor U3399 (N_3399,N_3002,N_1054);
and U3400 (N_3400,N_2144,N_275);
or U3401 (N_3401,N_2663,N_2803);
nor U3402 (N_3402,N_1766,N_393);
nor U3403 (N_3403,N_2724,N_1394);
nand U3404 (N_3404,N_1274,N_1128);
nor U3405 (N_3405,N_2252,N_1764);
xnor U3406 (N_3406,N_106,N_305);
xnor U3407 (N_3407,N_1008,N_312);
nor U3408 (N_3408,N_1876,N_912);
nand U3409 (N_3409,N_853,N_1060);
xnor U3410 (N_3410,N_2444,N_2336);
xor U3411 (N_3411,N_739,N_1391);
nand U3412 (N_3412,N_1360,N_1378);
or U3413 (N_3413,N_1470,N_1760);
or U3414 (N_3414,N_2026,N_891);
and U3415 (N_3415,N_2797,N_2647);
or U3416 (N_3416,N_1925,N_1736);
nor U3417 (N_3417,N_54,N_313);
nand U3418 (N_3418,N_2492,N_3078);
and U3419 (N_3419,N_2965,N_2089);
xor U3420 (N_3420,N_1059,N_470);
nand U3421 (N_3421,N_2142,N_410);
nor U3422 (N_3422,N_869,N_1175);
and U3423 (N_3423,N_2421,N_1776);
and U3424 (N_3424,N_424,N_2123);
and U3425 (N_3425,N_2656,N_554);
and U3426 (N_3426,N_2590,N_717);
nor U3427 (N_3427,N_1268,N_1944);
nand U3428 (N_3428,N_1913,N_1149);
nand U3429 (N_3429,N_771,N_688);
and U3430 (N_3430,N_1682,N_1761);
and U3431 (N_3431,N_1890,N_613);
and U3432 (N_3432,N_2056,N_460);
or U3433 (N_3433,N_62,N_1561);
and U3434 (N_3434,N_1739,N_310);
nor U3435 (N_3435,N_2171,N_746);
or U3436 (N_3436,N_2830,N_573);
nand U3437 (N_3437,N_2219,N_252);
xor U3438 (N_3438,N_2499,N_983);
nand U3439 (N_3439,N_86,N_2429);
xnor U3440 (N_3440,N_337,N_1397);
or U3441 (N_3441,N_2178,N_2189);
and U3442 (N_3442,N_1359,N_1078);
xnor U3443 (N_3443,N_3071,N_2648);
nand U3444 (N_3444,N_1412,N_2236);
xor U3445 (N_3445,N_2467,N_1617);
xor U3446 (N_3446,N_1758,N_3046);
and U3447 (N_3447,N_2943,N_1827);
xnor U3448 (N_3448,N_2300,N_1697);
and U3449 (N_3449,N_2478,N_1488);
nor U3450 (N_3450,N_2629,N_2749);
and U3451 (N_3451,N_1893,N_2274);
nor U3452 (N_3452,N_812,N_2864);
xor U3453 (N_3453,N_2293,N_849);
and U3454 (N_3454,N_1416,N_226);
and U3455 (N_3455,N_535,N_2465);
nor U3456 (N_3456,N_786,N_3061);
and U3457 (N_3457,N_544,N_829);
nor U3458 (N_3458,N_1901,N_987);
and U3459 (N_3459,N_523,N_81);
nor U3460 (N_3460,N_1325,N_1738);
xor U3461 (N_3461,N_850,N_788);
xnor U3462 (N_3462,N_539,N_107);
nor U3463 (N_3463,N_360,N_2173);
and U3464 (N_3464,N_2454,N_91);
nand U3465 (N_3465,N_364,N_2310);
nand U3466 (N_3466,N_2201,N_1546);
xor U3467 (N_3467,N_2876,N_165);
nand U3468 (N_3468,N_1991,N_2064);
nor U3469 (N_3469,N_537,N_1186);
xor U3470 (N_3470,N_2968,N_1319);
and U3471 (N_3471,N_1248,N_208);
and U3472 (N_3472,N_2416,N_1136);
nand U3473 (N_3473,N_1082,N_666);
xnor U3474 (N_3474,N_285,N_2024);
xor U3475 (N_3475,N_835,N_1091);
or U3476 (N_3476,N_2453,N_1179);
and U3477 (N_3477,N_2275,N_1536);
nand U3478 (N_3478,N_1263,N_2490);
xnor U3479 (N_3479,N_737,N_993);
or U3480 (N_3480,N_1563,N_2487);
nand U3481 (N_3481,N_889,N_1487);
nand U3482 (N_3482,N_2890,N_2937);
nor U3483 (N_3483,N_1918,N_2822);
nand U3484 (N_3484,N_1259,N_2958);
nand U3485 (N_3485,N_1953,N_1012);
nand U3486 (N_3486,N_1345,N_1204);
xor U3487 (N_3487,N_3102,N_1757);
and U3488 (N_3488,N_1130,N_2598);
or U3489 (N_3489,N_1424,N_2887);
nand U3490 (N_3490,N_1227,N_2719);
nor U3491 (N_3491,N_811,N_2294);
or U3492 (N_3492,N_110,N_1243);
and U3493 (N_3493,N_2970,N_1139);
and U3494 (N_3494,N_256,N_2690);
xnor U3495 (N_3495,N_1971,N_268);
and U3496 (N_3496,N_1068,N_214);
nand U3497 (N_3497,N_842,N_2199);
or U3498 (N_3498,N_2066,N_825);
nand U3499 (N_3499,N_433,N_1662);
nor U3500 (N_3500,N_1596,N_773);
or U3501 (N_3501,N_1142,N_2865);
nor U3502 (N_3502,N_2593,N_2554);
and U3503 (N_3503,N_47,N_2788);
and U3504 (N_3504,N_201,N_7);
nor U3505 (N_3505,N_2976,N_2254);
nor U3506 (N_3506,N_1646,N_2603);
xor U3507 (N_3507,N_1932,N_349);
xor U3508 (N_3508,N_2745,N_1580);
nor U3509 (N_3509,N_494,N_1011);
xor U3510 (N_3510,N_1177,N_2678);
nor U3511 (N_3511,N_187,N_3025);
nand U3512 (N_3512,N_2776,N_2119);
and U3513 (N_3513,N_945,N_1057);
nand U3514 (N_3514,N_2185,N_168);
nand U3515 (N_3515,N_2778,N_634);
or U3516 (N_3516,N_2074,N_239);
and U3517 (N_3517,N_2532,N_1885);
and U3518 (N_3518,N_1850,N_647);
xnor U3519 (N_3519,N_1027,N_1829);
and U3520 (N_3520,N_2857,N_3042);
or U3521 (N_3521,N_770,N_1314);
or U3522 (N_3522,N_2609,N_2963);
or U3523 (N_3523,N_272,N_713);
and U3524 (N_3524,N_2289,N_2179);
xnor U3525 (N_3525,N_140,N_2748);
xnor U3526 (N_3526,N_3055,N_1317);
and U3527 (N_3527,N_2152,N_432);
xnor U3528 (N_3528,N_202,N_1727);
nand U3529 (N_3529,N_614,N_950);
nor U3530 (N_3530,N_694,N_2269);
or U3531 (N_3531,N_609,N_616);
and U3532 (N_3532,N_2296,N_1109);
and U3533 (N_3533,N_1722,N_2838);
xor U3534 (N_3534,N_78,N_2315);
and U3535 (N_3535,N_143,N_2685);
nor U3536 (N_3536,N_1079,N_2659);
or U3537 (N_3537,N_1245,N_582);
nand U3538 (N_3538,N_2885,N_1493);
nor U3539 (N_3539,N_1694,N_2732);
and U3540 (N_3540,N_1419,N_984);
nor U3541 (N_3541,N_1153,N_2610);
and U3542 (N_3542,N_1562,N_538);
or U3543 (N_3543,N_2409,N_2560);
nand U3544 (N_3544,N_437,N_464);
and U3545 (N_3545,N_1966,N_954);
or U3546 (N_3546,N_2460,N_427);
and U3547 (N_3547,N_796,N_1604);
xor U3548 (N_3548,N_704,N_230);
or U3549 (N_3549,N_2516,N_949);
xor U3550 (N_3550,N_1176,N_1280);
nand U3551 (N_3551,N_1864,N_1403);
and U3552 (N_3552,N_1147,N_1937);
and U3553 (N_3553,N_2626,N_2716);
or U3554 (N_3554,N_1938,N_1454);
xor U3555 (N_3555,N_532,N_738);
xor U3556 (N_3556,N_2673,N_2573);
and U3557 (N_3557,N_2839,N_676);
and U3558 (N_3558,N_2808,N_1804);
nand U3559 (N_3559,N_1069,N_804);
or U3560 (N_3560,N_2447,N_3006);
or U3561 (N_3561,N_2231,N_817);
xnor U3562 (N_3562,N_373,N_681);
nand U3563 (N_3563,N_2886,N_1242);
xnor U3564 (N_3564,N_1585,N_1808);
or U3565 (N_3565,N_452,N_469);
and U3566 (N_3566,N_1009,N_618);
and U3567 (N_3567,N_2352,N_3091);
nand U3568 (N_3568,N_711,N_1313);
xnor U3569 (N_3569,N_2348,N_731);
and U3570 (N_3570,N_867,N_1406);
or U3571 (N_3571,N_1039,N_1163);
and U3572 (N_3572,N_870,N_2455);
and U3573 (N_3573,N_543,N_2681);
xnor U3574 (N_3574,N_1,N_1231);
and U3575 (N_3575,N_1185,N_1538);
nand U3576 (N_3576,N_2509,N_1730);
nor U3577 (N_3577,N_1066,N_79);
or U3578 (N_3578,N_790,N_1615);
and U3579 (N_3579,N_392,N_271);
and U3580 (N_3580,N_644,N_2750);
and U3581 (N_3581,N_1958,N_466);
and U3582 (N_3582,N_818,N_1713);
or U3583 (N_3583,N_621,N_3047);
nor U3584 (N_3584,N_1407,N_2795);
xnor U3585 (N_3585,N_2196,N_188);
xor U3586 (N_3586,N_2625,N_1133);
nor U3587 (N_3587,N_1672,N_657);
xnor U3588 (N_3588,N_1374,N_148);
or U3589 (N_3589,N_43,N_38);
xor U3590 (N_3590,N_174,N_1169);
nand U3591 (N_3591,N_2203,N_1903);
nand U3592 (N_3592,N_3085,N_2919);
and U3593 (N_3593,N_2556,N_2613);
xor U3594 (N_3594,N_2264,N_1888);
and U3595 (N_3595,N_249,N_1190);
and U3596 (N_3596,N_16,N_1492);
nand U3597 (N_3597,N_1220,N_1459);
xnor U3598 (N_3598,N_703,N_2316);
or U3599 (N_3599,N_1428,N_68);
nand U3600 (N_3600,N_415,N_2106);
nand U3601 (N_3601,N_2032,N_186);
or U3602 (N_3602,N_2000,N_595);
or U3603 (N_3603,N_591,N_570);
and U3604 (N_3604,N_815,N_2342);
nand U3605 (N_3605,N_5,N_2926);
nand U3606 (N_3606,N_772,N_3067);
xor U3607 (N_3607,N_986,N_1652);
nor U3608 (N_3608,N_3020,N_2321);
or U3609 (N_3609,N_1221,N_1496);
nor U3610 (N_3610,N_1599,N_721);
and U3611 (N_3611,N_3007,N_142);
nand U3612 (N_3612,N_1326,N_789);
and U3613 (N_3613,N_495,N_1989);
xnor U3614 (N_3614,N_1239,N_1540);
nor U3615 (N_3615,N_2019,N_1915);
nand U3616 (N_3616,N_1440,N_3080);
nor U3617 (N_3617,N_389,N_2436);
nor U3618 (N_3618,N_504,N_58);
nor U3619 (N_3619,N_2905,N_343);
and U3620 (N_3620,N_1628,N_1909);
or U3621 (N_3621,N_1752,N_1950);
xor U3622 (N_3622,N_2451,N_132);
xor U3623 (N_3623,N_488,N_197);
nand U3624 (N_3624,N_87,N_2755);
xnor U3625 (N_3625,N_2027,N_2558);
nand U3626 (N_3626,N_1667,N_542);
or U3627 (N_3627,N_2491,N_2771);
xnor U3628 (N_3628,N_1436,N_2368);
and U3629 (N_3629,N_2974,N_560);
xor U3630 (N_3630,N_370,N_2841);
and U3631 (N_3631,N_185,N_1348);
nor U3632 (N_3632,N_451,N_938);
nand U3633 (N_3633,N_547,N_27);
nand U3634 (N_3634,N_1393,N_923);
nand U3635 (N_3635,N_698,N_683);
and U3636 (N_3636,N_565,N_231);
or U3637 (N_3637,N_293,N_2503);
nor U3638 (N_3638,N_1504,N_383);
or U3639 (N_3639,N_757,N_2457);
xor U3640 (N_3640,N_473,N_1399);
or U3641 (N_3641,N_1339,N_2267);
xor U3642 (N_3642,N_648,N_2912);
or U3643 (N_3643,N_758,N_61);
or U3644 (N_3644,N_2502,N_2644);
and U3645 (N_3645,N_1132,N_2263);
xor U3646 (N_3646,N_1215,N_367);
nand U3647 (N_3647,N_3013,N_2978);
and U3648 (N_3648,N_1547,N_19);
or U3649 (N_3649,N_2466,N_1058);
and U3650 (N_3650,N_699,N_2400);
xnor U3651 (N_3651,N_1611,N_2009);
or U3652 (N_3652,N_308,N_2098);
and U3653 (N_3653,N_2223,N_209);
nor U3654 (N_3654,N_1728,N_2917);
or U3655 (N_3655,N_2543,N_3075);
or U3656 (N_3656,N_189,N_724);
nor U3657 (N_3657,N_2017,N_2544);
and U3658 (N_3658,N_1787,N_932);
xnor U3659 (N_3659,N_642,N_791);
nor U3660 (N_3660,N_1930,N_266);
nor U3661 (N_3661,N_2530,N_1427);
nand U3662 (N_3662,N_1701,N_2129);
and U3663 (N_3663,N_342,N_2835);
and U3664 (N_3664,N_1420,N_1969);
and U3665 (N_3665,N_2304,N_1516);
nor U3666 (N_3666,N_1125,N_2278);
xor U3667 (N_3667,N_2706,N_1298);
nor U3668 (N_3668,N_3099,N_2405);
or U3669 (N_3669,N_951,N_530);
and U3670 (N_3670,N_1279,N_2760);
nand U3671 (N_3671,N_2836,N_1648);
and U3672 (N_3672,N_1641,N_2136);
or U3673 (N_3673,N_480,N_834);
nand U3674 (N_3674,N_514,N_882);
nand U3675 (N_3675,N_2398,N_1527);
nand U3676 (N_3676,N_1978,N_1213);
and U3677 (N_3677,N_402,N_2866);
nand U3678 (N_3678,N_115,N_1045);
and U3679 (N_3679,N_2209,N_2134);
or U3680 (N_3680,N_1886,N_442);
and U3681 (N_3681,N_2043,N_435);
nand U3682 (N_3682,N_2848,N_1845);
and U3683 (N_3683,N_1545,N_1920);
and U3684 (N_3684,N_2935,N_1405);
or U3685 (N_3685,N_982,N_2882);
or U3686 (N_3686,N_777,N_1444);
nor U3687 (N_3687,N_1452,N_1921);
and U3688 (N_3688,N_2397,N_1509);
or U3689 (N_3689,N_3107,N_1387);
and U3690 (N_3690,N_1385,N_3066);
nor U3691 (N_3691,N_3117,N_3060);
xor U3692 (N_3692,N_1791,N_2365);
or U3693 (N_3693,N_587,N_2709);
or U3694 (N_3694,N_1104,N_2226);
nor U3695 (N_3695,N_1018,N_1825);
xnor U3696 (N_3696,N_2928,N_1505);
and U3697 (N_3697,N_328,N_2262);
xnor U3698 (N_3698,N_1853,N_1056);
nand U3699 (N_3699,N_2698,N_1192);
nand U3700 (N_3700,N_1836,N_2962);
nor U3701 (N_3701,N_2862,N_323);
xor U3702 (N_3702,N_1622,N_2099);
and U3703 (N_3703,N_1140,N_2200);
and U3704 (N_3704,N_1731,N_2045);
nand U3705 (N_3705,N_836,N_679);
or U3706 (N_3706,N_1010,N_640);
nand U3707 (N_3707,N_1575,N_2627);
and U3708 (N_3708,N_1129,N_487);
and U3709 (N_3709,N_2292,N_2094);
xnor U3710 (N_3710,N_1432,N_541);
nor U3711 (N_3711,N_794,N_99);
nand U3712 (N_3712,N_1777,N_1218);
nand U3713 (N_3713,N_2441,N_3057);
nor U3714 (N_3714,N_477,N_2941);
or U3715 (N_3715,N_1840,N_421);
xnor U3716 (N_3716,N_1026,N_851);
or U3717 (N_3717,N_1352,N_2594);
or U3718 (N_3718,N_1987,N_718);
and U3719 (N_3719,N_1303,N_669);
and U3720 (N_3720,N_430,N_813);
nor U3721 (N_3721,N_162,N_1193);
xnor U3722 (N_3722,N_263,N_2789);
nor U3723 (N_3723,N_1647,N_2082);
nor U3724 (N_3724,N_2233,N_1830);
nand U3725 (N_3725,N_203,N_734);
xor U3726 (N_3726,N_1621,N_1986);
xnor U3727 (N_3727,N_909,N_6);
and U3728 (N_3728,N_612,N_1675);
or U3729 (N_3729,N_1788,N_2637);
and U3730 (N_3730,N_751,N_685);
or U3731 (N_3731,N_1594,N_2095);
nand U3732 (N_3732,N_444,N_1308);
nor U3733 (N_3733,N_2938,N_2675);
and U3734 (N_3734,N_1094,N_2081);
xnor U3735 (N_3735,N_674,N_314);
nor U3736 (N_3736,N_2856,N_1124);
nor U3737 (N_3737,N_2850,N_2946);
or U3738 (N_3738,N_611,N_2504);
nor U3739 (N_3739,N_157,N_915);
or U3740 (N_3740,N_1098,N_2723);
nand U3741 (N_3741,N_1017,N_1601);
or U3742 (N_3742,N_1566,N_105);
nand U3743 (N_3743,N_2811,N_2430);
and U3744 (N_3744,N_496,N_910);
xnor U3745 (N_3745,N_1460,N_1285);
nor U3746 (N_3746,N_238,N_1768);
nor U3747 (N_3747,N_572,N_42);
or U3748 (N_3748,N_1995,N_405);
nor U3749 (N_3749,N_1572,N_1210);
nor U3750 (N_3750,N_1609,N_1588);
or U3751 (N_3751,N_2373,N_467);
xnor U3752 (N_3752,N_1437,N_1821);
xnor U3753 (N_3753,N_563,N_318);
and U3754 (N_3754,N_1302,N_2158);
or U3755 (N_3755,N_904,N_2224);
or U3756 (N_3756,N_1734,N_2305);
nor U3757 (N_3757,N_2055,N_637);
nand U3758 (N_3758,N_1674,N_274);
nor U3759 (N_3759,N_3058,N_1286);
nor U3760 (N_3760,N_1774,N_2618);
and U3761 (N_3761,N_114,N_1595);
or U3762 (N_3762,N_498,N_1376);
or U3763 (N_3763,N_927,N_2443);
nand U3764 (N_3764,N_1222,N_619);
nor U3765 (N_3765,N_1826,N_732);
nor U3766 (N_3766,N_1858,N_1315);
nand U3767 (N_3767,N_400,N_2020);
xor U3768 (N_3768,N_235,N_2364);
and U3769 (N_3769,N_2143,N_2340);
nand U3770 (N_3770,N_348,N_2221);
nor U3771 (N_3771,N_1865,N_877);
and U3772 (N_3772,N_150,N_36);
or U3773 (N_3773,N_149,N_1415);
xor U3774 (N_3774,N_3019,N_445);
or U3775 (N_3775,N_2918,N_996);
or U3776 (N_3776,N_1361,N_2210);
and U3777 (N_3777,N_2084,N_406);
and U3778 (N_3778,N_167,N_2104);
and U3779 (N_3779,N_2670,N_2258);
or U3780 (N_3780,N_1015,N_844);
or U3781 (N_3781,N_2357,N_766);
or U3782 (N_3782,N_8,N_3072);
nor U3783 (N_3783,N_1202,N_956);
nor U3784 (N_3784,N_885,N_462);
nor U3785 (N_3785,N_193,N_3056);
nand U3786 (N_3786,N_2794,N_431);
nand U3787 (N_3787,N_1894,N_3029);
nand U3788 (N_3788,N_2535,N_2410);
nor U3789 (N_3789,N_2459,N_562);
or U3790 (N_3790,N_3051,N_3011);
and U3791 (N_3791,N_423,N_1678);
nor U3792 (N_3792,N_1258,N_1102);
nor U3793 (N_3793,N_352,N_729);
nand U3794 (N_3794,N_380,N_2044);
nand U3795 (N_3795,N_2622,N_1997);
nor U3796 (N_3796,N_304,N_1228);
and U3797 (N_3797,N_2765,N_1763);
xnor U3798 (N_3798,N_808,N_2805);
and U3799 (N_3799,N_733,N_1692);
nand U3800 (N_3800,N_1157,N_2168);
nor U3801 (N_3801,N_2029,N_75);
or U3802 (N_3802,N_141,N_888);
nand U3803 (N_3803,N_1441,N_2781);
or U3804 (N_3804,N_2907,N_622);
nand U3805 (N_3805,N_3096,N_172);
or U3806 (N_3806,N_1838,N_2854);
and U3807 (N_3807,N_2072,N_822);
or U3808 (N_3808,N_2494,N_2472);
or U3809 (N_3809,N_1271,N_2893);
nand U3810 (N_3810,N_643,N_2010);
and U3811 (N_3811,N_260,N_490);
and U3812 (N_3812,N_84,N_2138);
and U3813 (N_3813,N_1367,N_2419);
xor U3814 (N_3814,N_2528,N_913);
and U3815 (N_3815,N_1358,N_3088);
nand U3816 (N_3816,N_2661,N_2025);
nor U3817 (N_3817,N_2696,N_1892);
nand U3818 (N_3818,N_49,N_1981);
nor U3819 (N_3819,N_2608,N_1849);
xnor U3820 (N_3820,N_2580,N_2983);
xnor U3821 (N_3821,N_340,N_2883);
or U3822 (N_3822,N_40,N_2578);
and U3823 (N_3823,N_1988,N_903);
and U3824 (N_3824,N_222,N_1043);
xor U3825 (N_3825,N_1055,N_1126);
nand U3826 (N_3826,N_1246,N_2775);
or U3827 (N_3827,N_2058,N_2282);
nand U3828 (N_3828,N_936,N_740);
and U3829 (N_3829,N_1625,N_1658);
xor U3830 (N_3830,N_2235,N_837);
xnor U3831 (N_3831,N_2088,N_1772);
nor U3832 (N_3832,N_561,N_3103);
nor U3833 (N_3833,N_973,N_1351);
and U3834 (N_3834,N_620,N_2700);
and U3835 (N_3835,N_1322,N_2867);
xnor U3836 (N_3836,N_2014,N_1805);
xnor U3837 (N_3837,N_2694,N_2344);
and U3838 (N_3838,N_2939,N_3120);
or U3839 (N_3839,N_1486,N_1832);
nor U3840 (N_3840,N_1188,N_1719);
nand U3841 (N_3841,N_3044,N_1873);
xnor U3842 (N_3842,N_1417,N_1143);
or U3843 (N_3843,N_236,N_1244);
xor U3844 (N_3844,N_1743,N_1700);
or U3845 (N_3845,N_1735,N_327);
nand U3846 (N_3846,N_3093,N_3039);
nor U3847 (N_3847,N_2003,N_2109);
nor U3848 (N_3848,N_257,N_2980);
or U3849 (N_3849,N_1755,N_3079);
and U3850 (N_3850,N_606,N_2858);
and U3851 (N_3851,N_1340,N_377);
xnor U3852 (N_3852,N_1061,N_237);
nor U3853 (N_3853,N_2564,N_1813);
and U3854 (N_3854,N_1815,N_1725);
xor U3855 (N_3855,N_1999,N_2523);
nand U3856 (N_3856,N_1240,N_1295);
nand U3857 (N_3857,N_2208,N_2955);
xnor U3858 (N_3858,N_702,N_1696);
nand U3859 (N_3859,N_2450,N_2013);
and U3860 (N_3860,N_859,N_624);
nor U3861 (N_3861,N_20,N_991);
nand U3862 (N_3862,N_1741,N_971);
and U3863 (N_3863,N_66,N_14);
xor U3864 (N_3864,N_1923,N_1897);
xnor U3865 (N_3865,N_605,N_227);
nor U3866 (N_3866,N_2076,N_2565);
or U3867 (N_3867,N_2065,N_2568);
or U3868 (N_3868,N_3121,N_333);
and U3869 (N_3869,N_2914,N_3052);
nor U3870 (N_3870,N_2911,N_2424);
nor U3871 (N_3871,N_1824,N_2334);
nor U3872 (N_3872,N_2011,N_2636);
and U3873 (N_3873,N_32,N_1954);
xor U3874 (N_3874,N_1431,N_714);
nand U3875 (N_3875,N_2018,N_265);
or U3876 (N_3876,N_2641,N_2420);
xnor U3877 (N_3877,N_890,N_2704);
xnor U3878 (N_3878,N_2339,N_1687);
nor U3879 (N_3879,N_576,N_948);
nor U3880 (N_3880,N_2966,N_1518);
nor U3881 (N_3881,N_331,N_980);
nor U3882 (N_3882,N_1483,N_3004);
nand U3883 (N_3883,N_2902,N_2739);
xor U3884 (N_3884,N_1032,N_196);
or U3885 (N_3885,N_902,N_1324);
nand U3886 (N_3886,N_2291,N_2900);
or U3887 (N_3887,N_2934,N_898);
nand U3888 (N_3888,N_2936,N_2826);
nand U3889 (N_3889,N_696,N_2445);
xor U3890 (N_3890,N_366,N_2180);
and U3891 (N_3891,N_947,N_2449);
nand U3892 (N_3892,N_589,N_334);
and U3893 (N_3893,N_2693,N_2360);
xnor U3894 (N_3894,N_1573,N_2680);
and U3895 (N_3895,N_2634,N_2829);
and U3896 (N_3896,N_2960,N_768);
or U3897 (N_3897,N_660,N_2163);
xnor U3898 (N_3898,N_220,N_3034);
nand U3899 (N_3899,N_839,N_2401);
nor U3900 (N_3900,N_823,N_1533);
xor U3901 (N_3901,N_146,N_1567);
and U3902 (N_3902,N_1841,N_1155);
xor U3903 (N_3903,N_1963,N_546);
xor U3904 (N_3904,N_96,N_1508);
and U3905 (N_3905,N_1146,N_761);
nor U3906 (N_3906,N_2232,N_1726);
nand U3907 (N_3907,N_64,N_1695);
xnor U3908 (N_3908,N_9,N_515);
xnor U3909 (N_3909,N_2510,N_262);
nand U3910 (N_3910,N_315,N_838);
nor U3911 (N_3911,N_2046,N_1232);
or U3912 (N_3912,N_2121,N_356);
or U3913 (N_3913,N_2628,N_2356);
or U3914 (N_3914,N_97,N_1497);
xor U3915 (N_3915,N_320,N_1984);
nor U3916 (N_3916,N_919,N_940);
xor U3917 (N_3917,N_3009,N_3048);
nand U3918 (N_3918,N_1589,N_192);
and U3919 (N_3919,N_557,N_2349);
nand U3920 (N_3920,N_3015,N_604);
or U3921 (N_3921,N_1767,N_2743);
or U3922 (N_3922,N_574,N_1586);
nor U3923 (N_3923,N_250,N_2650);
nor U3924 (N_3924,N_952,N_558);
and U3925 (N_3925,N_1072,N_2176);
xor U3926 (N_3926,N_691,N_2243);
xnor U3927 (N_3927,N_2891,N_2425);
nand U3928 (N_3928,N_351,N_2351);
nand U3929 (N_3929,N_122,N_2692);
or U3930 (N_3930,N_69,N_2916);
nand U3931 (N_3931,N_593,N_2059);
nor U3932 (N_3932,N_298,N_2689);
nand U3933 (N_3933,N_579,N_759);
nor U3934 (N_3934,N_1637,N_2880);
nand U3935 (N_3935,N_2464,N_2114);
and U3936 (N_3936,N_2772,N_1423);
or U3937 (N_3937,N_2873,N_667);
nor U3938 (N_3938,N_434,N_1707);
or U3939 (N_3939,N_2950,N_3024);
xor U3940 (N_3940,N_1689,N_800);
xor U3941 (N_3941,N_1006,N_30);
nand U3942 (N_3942,N_1434,N_1251);
nand U3943 (N_3943,N_181,N_3073);
nor U3944 (N_3944,N_872,N_2821);
and U3945 (N_3945,N_1429,N_1866);
or U3946 (N_3946,N_1657,N_2279);
nor U3947 (N_3947,N_2396,N_545);
or U3948 (N_3948,N_1007,N_2851);
xor U3949 (N_3949,N_1120,N_2899);
nand U3950 (N_3950,N_56,N_1372);
nor U3951 (N_3951,N_860,N_1564);
and U3952 (N_3952,N_1834,N_399);
or U3953 (N_3953,N_3021,N_881);
and U3954 (N_3954,N_1023,N_1523);
or U3955 (N_3955,N_2358,N_1224);
xnor U3956 (N_3956,N_2584,N_412);
nor U3957 (N_3957,N_2571,N_2695);
nor U3958 (N_3958,N_2913,N_1281);
or U3959 (N_3959,N_1653,N_2534);
xnor U3960 (N_3960,N_1600,N_1291);
or U3961 (N_3961,N_2697,N_2575);
and U3962 (N_3962,N_1854,N_2782);
nand U3963 (N_3963,N_378,N_2198);
xnor U3964 (N_3964,N_2122,N_2714);
nor U3965 (N_3965,N_1334,N_590);
nor U3966 (N_3966,N_692,N_754);
and U3967 (N_3967,N_2206,N_2154);
xnor U3968 (N_3968,N_625,N_1491);
nor U3969 (N_3969,N_326,N_646);
xnor U3970 (N_3970,N_1448,N_134);
xnor U3971 (N_3971,N_309,N_1952);
and U3972 (N_3972,N_1512,N_2313);
or U3973 (N_3973,N_407,N_712);
nand U3974 (N_3974,N_635,N_1331);
nand U3975 (N_3975,N_1257,N_2403);
xnor U3976 (N_3976,N_3016,N_2427);
or U3977 (N_3977,N_2868,N_1668);
and U3978 (N_3978,N_1602,N_2175);
nor U3979 (N_3979,N_154,N_2809);
or U3980 (N_3980,N_1238,N_2479);
nor U3981 (N_3981,N_457,N_580);
xor U3982 (N_3982,N_2645,N_1449);
nor U3983 (N_3983,N_22,N_652);
and U3984 (N_3984,N_1307,N_1881);
and U3985 (N_3985,N_1900,N_2722);
nand U3986 (N_3986,N_1478,N_458);
and U3987 (N_3987,N_1028,N_2260);
and U3988 (N_3988,N_865,N_2677);
xnor U3989 (N_3989,N_2140,N_874);
xor U3990 (N_3990,N_2757,N_1842);
xor U3991 (N_3991,N_626,N_176);
nor U3992 (N_3992,N_1673,N_1531);
and U3993 (N_3993,N_1031,N_2828);
or U3994 (N_3994,N_1105,N_465);
and U3995 (N_3995,N_510,N_361);
or U3996 (N_3996,N_802,N_1402);
or U3997 (N_3997,N_111,N_819);
xnor U3998 (N_3998,N_109,N_522);
xor U3999 (N_3999,N_108,N_25);
and U4000 (N_4000,N_426,N_937);
and U4001 (N_4001,N_2652,N_1671);
or U4002 (N_4002,N_1265,N_2906);
nor U4003 (N_4003,N_404,N_1223);
nor U4004 (N_4004,N_592,N_985);
and U4005 (N_4005,N_1994,N_689);
nand U4006 (N_4006,N_2712,N_1443);
nor U4007 (N_4007,N_283,N_232);
or U4008 (N_4008,N_1337,N_2513);
nand U4009 (N_4009,N_1679,N_1979);
and U4010 (N_4010,N_1975,N_939);
xor U4011 (N_4011,N_1631,N_322);
and U4012 (N_4012,N_2408,N_2752);
xor U4013 (N_4013,N_583,N_1565);
and U4014 (N_4014,N_2054,N_2092);
or U4015 (N_4015,N_28,N_1127);
nand U4016 (N_4016,N_387,N_1408);
xnor U4017 (N_4017,N_2721,N_1203);
xnor U4018 (N_4018,N_2488,N_492);
or U4019 (N_4019,N_1467,N_118);
and U4020 (N_4020,N_468,N_1070);
xnor U4021 (N_4021,N_2052,N_1225);
xor U4022 (N_4022,N_2842,N_2079);
and U4023 (N_4023,N_103,N_1063);
xor U4024 (N_4024,N_2792,N_1005);
or U4025 (N_4025,N_507,N_2847);
nand U4026 (N_4026,N_2588,N_930);
or U4027 (N_4027,N_2547,N_516);
and U4028 (N_4028,N_1550,N_158);
nand U4029 (N_4029,N_357,N_964);
nand U4030 (N_4030,N_3108,N_686);
or U4031 (N_4031,N_294,N_661);
or U4032 (N_4032,N_2521,N_1252);
nor U4033 (N_4033,N_200,N_2947);
and U4034 (N_4034,N_1065,N_2920);
nor U4035 (N_4035,N_2507,N_1649);
and U4036 (N_4036,N_2814,N_1636);
and U4037 (N_4037,N_1949,N_2399);
nor U4038 (N_4038,N_2234,N_1632);
nand U4039 (N_4039,N_1558,N_2070);
nand U4040 (N_4040,N_911,N_2388);
nor U4041 (N_4041,N_2524,N_1810);
nor U4042 (N_4042,N_2785,N_325);
and U4043 (N_4043,N_2228,N_1173);
nor U4044 (N_4044,N_548,N_384);
and U4045 (N_4045,N_2579,N_1199);
or U4046 (N_4046,N_1762,N_2688);
nand U4047 (N_4047,N_1597,N_1992);
or U4048 (N_4048,N_2182,N_2686);
nor U4049 (N_4049,N_1445,N_133);
nand U4050 (N_4050,N_233,N_1316);
or U4051 (N_4051,N_2555,N_1475);
nor U4052 (N_4052,N_629,N_2668);
nor U4053 (N_4053,N_2621,N_481);
and U4054 (N_4054,N_2125,N_2391);
or U4055 (N_4055,N_2080,N_2498);
nor U4056 (N_4056,N_1514,N_1869);
nor U4057 (N_4057,N_2823,N_1906);
nor U4058 (N_4058,N_1929,N_990);
nand U4059 (N_4059,N_1619,N_1201);
and U4060 (N_4060,N_128,N_1773);
and U4061 (N_4061,N_1771,N_2930);
xnor U4062 (N_4062,N_2633,N_2738);
and U4063 (N_4063,N_1135,N_177);
xnor U4064 (N_4064,N_972,N_799);
nor U4065 (N_4065,N_871,N_1882);
nand U4066 (N_4066,N_1180,N_478);
and U4067 (N_4067,N_2100,N_2506);
xnor U4068 (N_4068,N_1278,N_529);
or U4069 (N_4069,N_2624,N_2662);
or U4070 (N_4070,N_974,N_1582);
or U4071 (N_4071,N_2005,N_1148);
nor U4072 (N_4072,N_2038,N_2030);
and U4073 (N_4073,N_1305,N_2971);
nand U4074 (N_4074,N_2485,N_2113);
nor U4075 (N_4075,N_2248,N_1576);
xnor U4076 (N_4076,N_1960,N_2664);
nand U4077 (N_4077,N_1481,N_2128);
or U4078 (N_4078,N_1846,N_436);
xor U4079 (N_4079,N_391,N_284);
or U4080 (N_4080,N_50,N_443);
or U4081 (N_4081,N_2483,N_1680);
xnor U4082 (N_4082,N_650,N_1323);
nand U4083 (N_4083,N_1386,N_2286);
nor U4084 (N_4084,N_1161,N_2869);
and U4085 (N_4085,N_286,N_3074);
nor U4086 (N_4086,N_2859,N_502);
nand U4087 (N_4087,N_1198,N_2733);
and U4088 (N_4088,N_2259,N_1318);
nor U4089 (N_4089,N_2325,N_2703);
and U4090 (N_4090,N_1254,N_2227);
nand U4091 (N_4091,N_2077,N_2600);
or U4092 (N_4092,N_743,N_2793);
nor U4093 (N_4093,N_1784,N_1266);
xnor U4094 (N_4094,N_2177,N_1980);
xor U4095 (N_4095,N_2901,N_2414);
nor U4096 (N_4096,N_18,N_166);
nor U4097 (N_4097,N_1051,N_169);
and U4098 (N_4098,N_2595,N_680);
xor U4099 (N_4099,N_1471,N_659);
xnor U4100 (N_4100,N_3,N_3082);
xor U4101 (N_4101,N_98,N_417);
or U4102 (N_4102,N_803,N_2964);
xor U4103 (N_4103,N_2323,N_564);
or U4104 (N_4104,N_976,N_163);
or U4105 (N_4105,N_649,N_178);
xor U4106 (N_4106,N_1398,N_1052);
nand U4107 (N_4107,N_755,N_3086);
xor U4108 (N_4108,N_880,N_981);
nor U4109 (N_4109,N_2999,N_1910);
or U4110 (N_4110,N_1080,N_2073);
xnor U4111 (N_4111,N_1895,N_1592);
nor U4112 (N_4112,N_1859,N_1603);
xor U4113 (N_4113,N_2063,N_1927);
or U4114 (N_4114,N_2164,N_2277);
nand U4115 (N_4115,N_155,N_1532);
nand U4116 (N_4116,N_2135,N_59);
nor U4117 (N_4117,N_2439,N_2314);
or U4118 (N_4118,N_2585,N_368);
and U4119 (N_4119,N_682,N_2806);
or U4120 (N_4120,N_831,N_1383);
nand U4121 (N_4121,N_1293,N_2537);
and U4122 (N_4122,N_2422,N_2087);
nor U4123 (N_4123,N_1669,N_756);
nand U4124 (N_4124,N_2145,N_2022);
xnor U4125 (N_4125,N_2434,N_989);
nand U4126 (N_4126,N_1857,N_2863);
xor U4127 (N_4127,N_1014,N_3124);
and U4128 (N_4128,N_306,N_645);
and U4129 (N_4129,N_2423,N_145);
xor U4130 (N_4130,N_21,N_845);
or U4131 (N_4131,N_783,N_1794);
or U4132 (N_4132,N_1948,N_3064);
xor U4133 (N_4133,N_1729,N_90);
and U4134 (N_4134,N_632,N_2550);
or U4135 (N_4135,N_1439,N_997);
or U4136 (N_4136,N_210,N_2);
and U4137 (N_4137,N_1024,N_2525);
nor U4138 (N_4138,N_2008,N_1544);
and U4139 (N_4139,N_2577,N_2389);
and U4140 (N_4140,N_3000,N_1342);
xor U4141 (N_4141,N_1993,N_291);
nor U4142 (N_4142,N_2249,N_12);
or U4143 (N_4143,N_453,N_821);
or U4144 (N_4144,N_324,N_3065);
xor U4145 (N_4145,N_2318,N_2740);
nand U4146 (N_4146,N_2720,N_2241);
nor U4147 (N_4147,N_182,N_160);
or U4148 (N_4148,N_2448,N_2761);
and U4149 (N_4149,N_1250,N_184);
nor U4150 (N_4150,N_2707,N_296);
and U4151 (N_4151,N_1798,N_1048);
and U4152 (N_4152,N_2500,N_3109);
or U4153 (N_4153,N_2514,N_1474);
and U4154 (N_4154,N_3054,N_1122);
and U4155 (N_4155,N_1447,N_1458);
or U4156 (N_4156,N_1839,N_1607);
and U4157 (N_4157,N_1583,N_615);
nand U4158 (N_4158,N_567,N_1414);
nor U4159 (N_4159,N_1119,N_1002);
and U4160 (N_4160,N_472,N_1004);
nand U4161 (N_4161,N_1801,N_2875);
nor U4162 (N_4162,N_1450,N_1333);
xnor U4163 (N_4163,N_977,N_11);
and U4164 (N_4164,N_1710,N_1050);
xnor U4165 (N_4165,N_1612,N_916);
xor U4166 (N_4166,N_1961,N_1705);
and U4167 (N_4167,N_1917,N_39);
or U4168 (N_4168,N_449,N_979);
nand U4169 (N_4169,N_2819,N_531);
nor U4170 (N_4170,N_65,N_2705);
nand U4171 (N_4171,N_398,N_2921);
and U4172 (N_4172,N_762,N_113);
nor U4173 (N_4173,N_2908,N_929);
xor U4174 (N_4174,N_2741,N_355);
and U4175 (N_4175,N_2597,N_2332);
nand U4176 (N_4176,N_1579,N_1703);
nand U4177 (N_4177,N_76,N_2133);
nor U4178 (N_4178,N_1290,N_1660);
nor U4179 (N_4179,N_1214,N_1581);
nor U4180 (N_4180,N_2989,N_1629);
and U4181 (N_4181,N_2984,N_2308);
nand U4182 (N_4182,N_1796,N_1020);
nor U4183 (N_4183,N_2238,N_282);
nor U4184 (N_4184,N_553,N_508);
nand U4185 (N_4185,N_1751,N_1754);
or U4186 (N_4186,N_1951,N_907);
nand U4187 (N_4187,N_500,N_2824);
nand U4188 (N_4188,N_2051,N_3122);
or U4189 (N_4189,N_693,N_1003);
xnor U4190 (N_4190,N_2319,N_1926);
nand U4191 (N_4191,N_3050,N_2619);
or U4192 (N_4192,N_300,N_70);
nand U4193 (N_4193,N_1097,N_1084);
or U4194 (N_4194,N_2744,N_95);
nor U4195 (N_4195,N_1828,N_2742);
xor U4196 (N_4196,N_2160,N_3037);
xor U4197 (N_4197,N_559,N_2091);
nor U4198 (N_4198,N_1297,N_2345);
nand U4199 (N_4199,N_13,N_863);
and U4200 (N_4200,N_2942,N_651);
nand U4201 (N_4201,N_234,N_840);
nand U4202 (N_4202,N_82,N_369);
nand U4203 (N_4203,N_3090,N_1721);
or U4204 (N_4204,N_1947,N_512);
nand U4205 (N_4205,N_2193,N_2927);
nor U4206 (N_4206,N_876,N_816);
or U4207 (N_4207,N_394,N_2230);
nor U4208 (N_4208,N_2042,N_1196);
and U4209 (N_4209,N_978,N_2390);
nand U4210 (N_4210,N_2801,N_1666);
and U4211 (N_4211,N_2520,N_1241);
nor U4212 (N_4212,N_741,N_1207);
nor U4213 (N_4213,N_303,N_2172);
and U4214 (N_4214,N_2979,N_1896);
or U4215 (N_4215,N_2711,N_3017);
nor U4216 (N_4216,N_2540,N_2285);
nand U4217 (N_4217,N_764,N_46);
or U4218 (N_4218,N_57,N_446);
nand U4219 (N_4219,N_2734,N_455);
or U4220 (N_4220,N_1327,N_1435);
nor U4221 (N_4221,N_2057,N_475);
or U4222 (N_4222,N_2350,N_2654);
nand U4223 (N_4223,N_1640,N_600);
xnor U4224 (N_4224,N_926,N_1807);
or U4225 (N_4225,N_2623,N_1101);
or U4226 (N_4226,N_1934,N_447);
nor U4227 (N_4227,N_1785,N_3003);
and U4228 (N_4228,N_2101,N_1092);
nor U4229 (N_4229,N_1584,N_2482);
xor U4230 (N_4230,N_1463,N_1753);
nand U4231 (N_4231,N_2237,N_1645);
nand U4232 (N_4232,N_886,N_1455);
and U4233 (N_4233,N_297,N_513);
xnor U4234 (N_4234,N_1965,N_1714);
and U4235 (N_4235,N_278,N_1156);
nand U4236 (N_4236,N_2338,N_279);
nand U4237 (N_4237,N_2324,N_935);
or U4238 (N_4238,N_123,N_267);
nor U4239 (N_4239,N_918,N_827);
and U4240 (N_4240,N_2973,N_765);
and U4241 (N_4241,N_1309,N_1353);
and U4242 (N_4242,N_1819,N_2433);
xor U4243 (N_4243,N_933,N_1778);
and U4244 (N_4244,N_1356,N_2229);
xnor U4245 (N_4245,N_2105,N_1843);
nor U4246 (N_4246,N_2151,N_709);
nand U4247 (N_4247,N_1712,N_2730);
and U4248 (N_4248,N_3030,N_476);
xnor U4249 (N_4249,N_1502,N_1907);
and U4250 (N_4250,N_1332,N_2944);
nand U4251 (N_4251,N_2307,N_243);
nand U4252 (N_4252,N_2337,N_2475);
and U4253 (N_4253,N_4,N_277);
xor U4254 (N_4254,N_524,N_2276);
nand U4255 (N_4255,N_778,N_2987);
or U4256 (N_4256,N_2169,N_1860);
nor U4257 (N_4257,N_92,N_2702);
nand U4258 (N_4258,N_1294,N_1606);
nor U4259 (N_4259,N_1379,N_2379);
nor U4260 (N_4260,N_2669,N_311);
or U4261 (N_4261,N_102,N_3049);
nor U4262 (N_4262,N_3101,N_1042);
nand U4263 (N_4263,N_479,N_1364);
and U4264 (N_4264,N_795,N_2187);
xnor U4265 (N_4265,N_943,N_153);
and U4266 (N_4266,N_607,N_2834);
and U4267 (N_4267,N_1715,N_3041);
or U4268 (N_4268,N_2783,N_346);
xnor U4269 (N_4269,N_533,N_3033);
or U4270 (N_4270,N_784,N_1528);
xnor U4271 (N_4271,N_2298,N_2538);
or U4272 (N_4272,N_2395,N_654);
or U4273 (N_4273,N_2212,N_1217);
xor U4274 (N_4274,N_2181,N_760);
or U4275 (N_4275,N_2542,N_89);
and U4276 (N_4276,N_173,N_1390);
xor U4277 (N_4277,N_416,N_2949);
and U4278 (N_4278,N_2631,N_1574);
and U4279 (N_4279,N_3040,N_2148);
and U4280 (N_4280,N_941,N_2363);
and U4281 (N_4281,N_2380,N_408);
or U4282 (N_4282,N_2413,N_1939);
and U4283 (N_4283,N_124,N_1479);
xor U4284 (N_4284,N_474,N_1328);
xor U4285 (N_4285,N_748,N_3115);
nand U4286 (N_4286,N_52,N_663);
and U4287 (N_4287,N_2132,N_1855);
nor U4288 (N_4288,N_228,N_2257);
xnor U4289 (N_4289,N_1433,N_301);
or U4290 (N_4290,N_1077,N_744);
xnor U4291 (N_4291,N_1928,N_1075);
or U4292 (N_4292,N_2359,N_2620);
or U4293 (N_4293,N_1187,N_2190);
nand U4294 (N_4294,N_2727,N_2954);
or U4295 (N_4295,N_2994,N_2299);
nand U4296 (N_4296,N_893,N_1685);
or U4297 (N_4297,N_489,N_1670);
and U4298 (N_4298,N_119,N_2371);
xnor U4299 (N_4299,N_1388,N_429);
nand U4300 (N_4300,N_1370,N_1797);
nand U4301 (N_4301,N_2833,N_3026);
nor U4302 (N_4302,N_1040,N_3081);
nor U4303 (N_4303,N_2922,N_2083);
nand U4304 (N_4304,N_1107,N_878);
nand U4305 (N_4305,N_3063,N_390);
nor U4306 (N_4306,N_2283,N_2787);
nor U4307 (N_4307,N_281,N_1693);
and U4308 (N_4308,N_1737,N_63);
nand U4309 (N_4309,N_2879,N_1145);
or U4310 (N_4310,N_1219,N_1083);
nand U4311 (N_4311,N_506,N_3097);
xnor U4312 (N_4312,N_1964,N_2601);
xnor U4313 (N_4313,N_1150,N_1490);
and U4314 (N_4314,N_1709,N_1473);
and U4315 (N_4315,N_2541,N_2799);
nand U4316 (N_4316,N_1404,N_2997);
nor U4317 (N_4317,N_319,N_2071);
xnor U4318 (N_4318,N_2211,N_809);
xnor U4319 (N_4319,N_1822,N_639);
and U4320 (N_4320,N_2428,N_212);
nand U4321 (N_4321,N_2642,N_1946);
xnor U4322 (N_4322,N_2103,N_1793);
nor U4323 (N_4323,N_1090,N_242);
xnor U4324 (N_4324,N_1972,N_287);
or U4325 (N_4325,N_1099,N_1494);
xnor U4326 (N_4326,N_1914,N_2362);
and U4327 (N_4327,N_2635,N_1933);
and U4328 (N_4328,N_1299,N_1748);
and U4329 (N_4329,N_1861,N_630);
or U4330 (N_4330,N_1038,N_1362);
xnor U4331 (N_4331,N_1790,N_2784);
and U4332 (N_4332,N_100,N_1733);
and U4333 (N_4333,N_1608,N_2309);
and U4334 (N_4334,N_1233,N_2329);
nor U4335 (N_4335,N_1976,N_85);
or U4336 (N_4336,N_23,N_258);
xnor U4337 (N_4337,N_1756,N_2141);
or U4338 (N_4338,N_2952,N_2426);
and U4339 (N_4339,N_2297,N_317);
nor U4340 (N_4340,N_1638,N_1395);
nor U4341 (N_4341,N_2194,N_41);
nand U4342 (N_4342,N_2377,N_1806);
nor U4343 (N_4343,N_2852,N_55);
or U4344 (N_4344,N_321,N_2126);
and U4345 (N_4345,N_454,N_2735);
xnor U4346 (N_4346,N_1111,N_586);
nor U4347 (N_4347,N_568,N_2496);
or U4348 (N_4348,N_94,N_1277);
nand U4349 (N_4349,N_270,N_505);
or U4350 (N_4350,N_83,N_617);
nand U4351 (N_4351,N_1551,N_1418);
nand U4352 (N_4352,N_362,N_855);
or U4353 (N_4353,N_597,N_1618);
or U4354 (N_4354,N_862,N_1524);
or U4355 (N_4355,N_959,N_80);
or U4356 (N_4356,N_3112,N_1067);
xnor U4357 (N_4357,N_2682,N_672);
xnor U4358 (N_4358,N_1795,N_1814);
or U4359 (N_4359,N_307,N_1365);
and U4360 (N_4360,N_1856,N_1570);
or U4361 (N_4361,N_627,N_2107);
or U4362 (N_4362,N_1197,N_1151);
nor U4363 (N_4363,N_2250,N_1802);
nor U4364 (N_4364,N_719,N_2295);
nand U4365 (N_4365,N_1453,N_1874);
nor U4366 (N_4366,N_2583,N_2728);
nand U4367 (N_4367,N_374,N_1206);
nor U4368 (N_4368,N_1103,N_1438);
xnor U4369 (N_4369,N_2432,N_3010);
xor U4370 (N_4370,N_1593,N_2023);
or U4371 (N_4371,N_2431,N_2326);
and U4372 (N_4372,N_15,N_2904);
or U4373 (N_4373,N_221,N_2589);
xnor U4374 (N_4374,N_1373,N_1462);
and U4375 (N_4375,N_2612,N_2036);
and U4376 (N_4376,N_3087,N_2853);
nor U4377 (N_4377,N_1655,N_967);
nand U4378 (N_4378,N_1468,N_2456);
and U4379 (N_4379,N_1818,N_2031);
and U4380 (N_4380,N_1273,N_503);
xnor U4381 (N_4381,N_217,N_2562);
or U4382 (N_4382,N_2484,N_1283);
xnor U4383 (N_4383,N_1870,N_456);
nand U4384 (N_4384,N_2840,N_151);
xnor U4385 (N_4385,N_101,N_2251);
nand U4386 (N_4386,N_1335,N_170);
nor U4387 (N_4387,N_3008,N_1868);
or U4388 (N_4388,N_1037,N_2166);
or U4389 (N_4389,N_1820,N_2271);
and U4390 (N_4390,N_509,N_35);
xor U4391 (N_4391,N_1837,N_448);
and U4392 (N_4392,N_2067,N_53);
xnor U4393 (N_4393,N_1510,N_1936);
nand U4394 (N_4394,N_1282,N_2767);
or U4395 (N_4395,N_1457,N_1288);
xor U4396 (N_4396,N_1740,N_2657);
and U4397 (N_4397,N_1001,N_2381);
xnor U4398 (N_4398,N_1656,N_3116);
nand U4399 (N_4399,N_1019,N_2392);
nand U4400 (N_4400,N_2773,N_2915);
nor U4401 (N_4401,N_752,N_428);
and U4402 (N_4402,N_2762,N_1073);
nor U4403 (N_4403,N_3119,N_74);
and U4404 (N_4404,N_2284,N_1541);
or U4405 (N_4405,N_931,N_1633);
nand U4406 (N_4406,N_71,N_875);
or U4407 (N_4407,N_2780,N_2006);
xnor U4408 (N_4408,N_144,N_1717);
nand U4409 (N_4409,N_1164,N_2470);
nor U4410 (N_4410,N_363,N_1642);
or U4411 (N_4411,N_2375,N_2097);
or U4412 (N_4412,N_199,N_1357);
or U4413 (N_4413,N_1742,N_675);
and U4414 (N_4414,N_1501,N_1062);
nor U4415 (N_4415,N_2587,N_2599);
nand U4416 (N_4416,N_2870,N_585);
or U4417 (N_4417,N_401,N_29);
or U4418 (N_4418,N_1287,N_486);
or U4419 (N_4419,N_248,N_601);
or U4420 (N_4420,N_2489,N_2137);
or U4421 (N_4421,N_382,N_2758);
nand U4422 (N_4422,N_1676,N_2684);
nor U4423 (N_4423,N_774,N_463);
nor U4424 (N_4424,N_1021,N_413);
nand U4425 (N_4425,N_1033,N_2552);
nand U4426 (N_4426,N_1330,N_3089);
xor U4427 (N_4427,N_2366,N_2481);
xor U4428 (N_4428,N_2085,N_1904);
or U4429 (N_4429,N_2411,N_386);
or U4430 (N_4430,N_1181,N_2446);
and U4431 (N_4431,N_1569,N_1456);
or U4432 (N_4432,N_2486,N_2312);
nand U4433 (N_4433,N_602,N_2522);
and U4434 (N_4434,N_353,N_1677);
xnor U4435 (N_4435,N_3036,N_1355);
nand U4436 (N_4436,N_2139,N_861);
nand U4437 (N_4437,N_1229,N_1115);
or U4438 (N_4438,N_2330,N_482);
and U4439 (N_4439,N_1905,N_549);
and U4440 (N_4440,N_1183,N_2205);
and U4441 (N_4441,N_2438,N_2402);
and U4442 (N_4442,N_3104,N_2048);
xor U4443 (N_4443,N_2800,N_2162);
or U4444 (N_4444,N_2894,N_3076);
and U4445 (N_4445,N_2909,N_2149);
and U4446 (N_4446,N_2049,N_1108);
and U4447 (N_4447,N_2306,N_1982);
xnor U4448 (N_4448,N_728,N_1053);
nor U4449 (N_4449,N_716,N_963);
nand U4450 (N_4450,N_438,N_422);
nand U4451 (N_4451,N_2874,N_1382);
xor U4452 (N_4452,N_864,N_2817);
and U4453 (N_4453,N_1880,N_1624);
nor U4454 (N_4454,N_1744,N_379);
or U4455 (N_4455,N_244,N_288);
or U4456 (N_4456,N_2878,N_2213);
xor U4457 (N_4457,N_1085,N_1159);
nor U4458 (N_4458,N_2977,N_2378);
nand U4459 (N_4459,N_17,N_1366);
nor U4460 (N_4460,N_1158,N_2273);
nand U4461 (N_4461,N_2972,N_536);
and U4462 (N_4462,N_2774,N_51);
and U4463 (N_4463,N_2002,N_1371);
xor U4464 (N_4464,N_873,N_2037);
and U4465 (N_4465,N_2115,N_2639);
nand U4466 (N_4466,N_1878,N_921);
or U4467 (N_4467,N_697,N_779);
or U4468 (N_4468,N_707,N_571);
or U4469 (N_4469,N_846,N_1472);
and U4470 (N_4470,N_2440,N_2153);
or U4471 (N_4471,N_824,N_3035);
or U4472 (N_4472,N_797,N_596);
and U4473 (N_4473,N_2591,N_2186);
and U4474 (N_4474,N_2825,N_1112);
xnor U4475 (N_4475,N_2159,N_897);
nand U4476 (N_4476,N_2990,N_958);
or U4477 (N_4477,N_2385,N_2343);
or U4478 (N_4478,N_2574,N_1256);
xnor U4479 (N_4479,N_1189,N_925);
nor U4480 (N_4480,N_1644,N_2047);
and U4481 (N_4481,N_215,N_656);
nand U4482 (N_4482,N_1916,N_2170);
and U4483 (N_4483,N_519,N_1025);
or U4484 (N_4484,N_1170,N_2317);
nor U4485 (N_4485,N_858,N_2053);
nand U4486 (N_4486,N_814,N_183);
xnor U4487 (N_4487,N_1034,N_2910);
and U4488 (N_4488,N_121,N_1852);
xor U4489 (N_4489,N_2110,N_1943);
xnor U4490 (N_4490,N_749,N_2192);
xnor U4491 (N_4491,N_899,N_1922);
and U4492 (N_4492,N_2881,N_1195);
or U4493 (N_4493,N_2493,N_2382);
and U4494 (N_4494,N_2039,N_588);
and U4495 (N_4495,N_2845,N_526);
and U4496 (N_4496,N_884,N_1369);
nor U4497 (N_4497,N_1267,N_2161);
and U4498 (N_4498,N_2183,N_2871);
nor U4499 (N_4499,N_339,N_1519);
xor U4500 (N_4500,N_2816,N_1591);
or U4501 (N_4501,N_960,N_1974);
xnor U4502 (N_4502,N_2632,N_1421);
nand U4503 (N_4503,N_2940,N_2461);
and U4504 (N_4504,N_194,N_1847);
xor U4505 (N_4505,N_895,N_1620);
nor U4506 (N_4506,N_1191,N_2651);
nand U4507 (N_4507,N_2846,N_828);
and U4508 (N_4508,N_1765,N_1803);
xor U4509 (N_4509,N_24,N_1160);
or U4510 (N_4510,N_942,N_584);
nand U4511 (N_4511,N_295,N_810);
or U4512 (N_4512,N_216,N_3100);
or U4513 (N_4513,N_1616,N_2028);
xor U4514 (N_4514,N_1973,N_179);
or U4515 (N_4515,N_381,N_1779);
or U4516 (N_4516,N_753,N_1506);
and U4517 (N_4517,N_2953,N_126);
and U4518 (N_4518,N_655,N_251);
and U4519 (N_4519,N_1178,N_1442);
xor U4520 (N_4520,N_120,N_540);
and U4521 (N_4521,N_1076,N_1329);
or U4522 (N_4522,N_1883,N_1983);
and U4523 (N_4523,N_1255,N_965);
xnor U4524 (N_4524,N_3032,N_1775);
and U4525 (N_4525,N_1698,N_2245);
nand U4526 (N_4526,N_1513,N_841);
or U4527 (N_4527,N_1100,N_2710);
and U4528 (N_4528,N_3045,N_1708);
and U4529 (N_4529,N_1430,N_2832);
nor U4530 (N_4530,N_3111,N_1499);
xor U4531 (N_4531,N_3098,N_1723);
xnor U4532 (N_4532,N_139,N_1044);
or U4533 (N_4533,N_1911,N_695);
nor U4534 (N_4534,N_594,N_1296);
nor U4535 (N_4535,N_2815,N_2546);
and U4536 (N_4536,N_1381,N_3106);
nor U4537 (N_4537,N_104,N_1212);
or U4538 (N_4538,N_2372,N_1912);
nor U4539 (N_4539,N_638,N_555);
nand U4540 (N_4540,N_2951,N_1182);
nand U4541 (N_4541,N_1639,N_900);
nor U4542 (N_4542,N_866,N_2301);
and U4543 (N_4543,N_1477,N_1746);
nand U4544 (N_4544,N_1812,N_2452);
or U4545 (N_4545,N_2786,N_2553);
or U4546 (N_4546,N_441,N_491);
nand U4547 (N_4547,N_2435,N_485);
nand U4548 (N_4548,N_673,N_787);
xor U4549 (N_4549,N_727,N_2069);
nand U4550 (N_4550,N_2303,N_3018);
and U4551 (N_4551,N_259,N_1571);
and U4552 (N_4552,N_1089,N_1663);
nand U4553 (N_4553,N_710,N_2355);
or U4554 (N_4554,N_969,N_905);
nand U4555 (N_4555,N_994,N_1940);
xor U4556 (N_4556,N_2147,N_1699);
or U4557 (N_4557,N_917,N_3094);
nand U4558 (N_4558,N_2961,N_3005);
xnor U4559 (N_4559,N_742,N_316);
xnor U4560 (N_4560,N_2246,N_2672);
nor U4561 (N_4561,N_1347,N_2995);
nand U4562 (N_4562,N_830,N_1167);
and U4563 (N_4563,N_1627,N_161);
and U4564 (N_4564,N_2468,N_388);
and U4565 (N_4565,N_528,N_1724);
nor U4566 (N_4566,N_735,N_2667);
or U4567 (N_4567,N_2218,N_420);
or U4568 (N_4568,N_2225,N_1409);
or U4569 (N_4569,N_2729,N_715);
nor U4570 (N_4570,N_1823,N_725);
nand U4571 (N_4571,N_1522,N_60);
nand U4572 (N_4572,N_2156,N_2982);
nor U4573 (N_4573,N_2993,N_820);
and U4574 (N_4574,N_2872,N_2458);
xor U4575 (N_4575,N_276,N_1114);
or U4576 (N_4576,N_1071,N_261);
nand U4577 (N_4577,N_2394,N_2280);
or U4578 (N_4578,N_2272,N_175);
nand U4579 (N_4579,N_1350,N_1955);
nand U4580 (N_4580,N_2333,N_2327);
and U4581 (N_4581,N_3069,N_1590);
and U4582 (N_4582,N_2256,N_1651);
and U4583 (N_4583,N_2831,N_2756);
nand U4584 (N_4584,N_2247,N_2660);
nand U4585 (N_4585,N_1863,N_2770);
nor U4586 (N_4586,N_1346,N_2197);
or U4587 (N_4587,N_1261,N_1872);
xor U4588 (N_4588,N_1800,N_1247);
nor U4589 (N_4589,N_1064,N_137);
or U4590 (N_4590,N_439,N_1410);
nand U4591 (N_4591,N_2630,N_397);
nand U4592 (N_4592,N_2239,N_1530);
or U4593 (N_4593,N_1485,N_1036);
nand U4594 (N_4594,N_928,N_1375);
nor U4595 (N_4595,N_1396,N_341);
xor U4596 (N_4596,N_995,N_2810);
nor U4597 (N_4597,N_290,N_2549);
xnor U4598 (N_4598,N_1635,N_1110);
nor U4599 (N_4599,N_1962,N_1587);
or U4600 (N_4600,N_2174,N_411);
xor U4601 (N_4601,N_2442,N_807);
nor U4602 (N_4602,N_780,N_2691);
xnor U4603 (N_4603,N_2616,N_2393);
xnor U4604 (N_4604,N_1879,N_34);
xnor U4605 (N_4605,N_2717,N_1284);
xor U4606 (N_4606,N_2412,N_2718);
xnor U4607 (N_4607,N_2545,N_1817);
nor U4608 (N_4608,N_2948,N_1634);
nand U4609 (N_4609,N_2820,N_1844);
nand U4610 (N_4610,N_3083,N_2124);
xor U4611 (N_4611,N_1899,N_2567);
and U4612 (N_4612,N_2287,N_330);
or U4613 (N_4613,N_2253,N_922);
nand U4614 (N_4614,N_1500,N_2477);
and U4615 (N_4615,N_2127,N_2001);
or U4616 (N_4616,N_344,N_610);
xor U4617 (N_4617,N_2335,N_1343);
and U4618 (N_4618,N_1154,N_906);
nor U4619 (N_4619,N_1230,N_3113);
nand U4620 (N_4620,N_152,N_219);
nand U4621 (N_4621,N_665,N_2146);
or U4622 (N_4622,N_501,N_2563);
or U4623 (N_4623,N_414,N_2998);
nor U4624 (N_4624,N_419,N_1959);
or U4625 (N_4625,N_879,N_2566);
nor U4626 (N_4626,N_970,N_1200);
xor U4627 (N_4627,N_2726,N_1349);
xor U4628 (N_4628,N_2060,N_1249);
and U4629 (N_4629,N_2602,N_2638);
and U4630 (N_4630,N_2188,N_1237);
or U4631 (N_4631,N_253,N_2746);
xor U4632 (N_4632,N_2108,N_156);
nor U4633 (N_4633,N_2895,N_750);
xor U4634 (N_4634,N_3110,N_1924);
or U4635 (N_4635,N_2614,N_798);
or U4636 (N_4636,N_2204,N_1321);
nand U4637 (N_4637,N_1957,N_1484);
or U4638 (N_4638,N_641,N_1235);
and U4639 (N_4639,N_2903,N_44);
and U4640 (N_4640,N_1088,N_1117);
or U4641 (N_4641,N_2240,N_1534);
nor U4642 (N_4642,N_2604,N_1884);
nor U4643 (N_4643,N_901,N_2288);
xnor U4644 (N_4644,N_1919,N_112);
xor U4645 (N_4645,N_207,N_2220);
and U4646 (N_4646,N_409,N_1665);
nor U4647 (N_4647,N_2582,N_961);
and U4648 (N_4648,N_1469,N_2517);
nor U4649 (N_4649,N_2331,N_2945);
or U4650 (N_4650,N_1041,N_131);
or U4651 (N_4651,N_2658,N_2495);
nor U4652 (N_4652,N_2376,N_358);
nand U4653 (N_4653,N_1968,N_2798);
xnor U4654 (N_4654,N_2112,N_3059);
nor U4655 (N_4655,N_2683,N_0);
xnor U4656 (N_4656,N_2531,N_2996);
nor U4657 (N_4657,N_3095,N_631);
and U4658 (N_4658,N_2222,N_2643);
nand U4659 (N_4659,N_2605,N_1568);
xor U4660 (N_4660,N_1461,N_2062);
nor U4661 (N_4661,N_534,N_345);
and U4662 (N_4662,N_1664,N_2827);
nor U4663 (N_4663,N_2766,N_2268);
xnor U4664 (N_4664,N_2617,N_1875);
and U4665 (N_4665,N_2536,N_664);
or U4666 (N_4666,N_1956,N_578);
or U4667 (N_4667,N_1030,N_292);
and U4668 (N_4668,N_2311,N_1262);
nor U4669 (N_4669,N_2526,N_1166);
xnor U4670 (N_4670,N_1770,N_1489);
and U4671 (N_4671,N_245,N_1451);
nor U4672 (N_4672,N_1336,N_1554);
nand U4673 (N_4673,N_1368,N_690);
xor U4674 (N_4674,N_2191,N_1465);
and U4675 (N_4675,N_1253,N_1809);
nand U4676 (N_4676,N_1686,N_2969);
nor U4677 (N_4677,N_499,N_2837);
nand U4678 (N_4678,N_1799,N_2384);
and U4679 (N_4679,N_1363,N_335);
nor U4680 (N_4680,N_1931,N_1867);
nand U4681 (N_4681,N_2505,N_1835);
xor U4682 (N_4682,N_1138,N_2215);
and U4683 (N_4683,N_1548,N_575);
xnor U4684 (N_4684,N_3038,N_2480);
and U4685 (N_4685,N_2861,N_2676);
xor U4686 (N_4686,N_1480,N_2035);
or U4687 (N_4687,N_2581,N_1771);
xor U4688 (N_4688,N_1548,N_2675);
or U4689 (N_4689,N_975,N_2867);
xnor U4690 (N_4690,N_864,N_1603);
xnor U4691 (N_4691,N_627,N_2830);
and U4692 (N_4692,N_512,N_1037);
nor U4693 (N_4693,N_2488,N_1882);
nand U4694 (N_4694,N_1658,N_2358);
nand U4695 (N_4695,N_699,N_1864);
nor U4696 (N_4696,N_1322,N_2403);
or U4697 (N_4697,N_2885,N_2098);
or U4698 (N_4698,N_1806,N_1679);
and U4699 (N_4699,N_938,N_1945);
xnor U4700 (N_4700,N_1154,N_2830);
xnor U4701 (N_4701,N_2019,N_314);
nand U4702 (N_4702,N_327,N_1763);
nor U4703 (N_4703,N_509,N_1945);
and U4704 (N_4704,N_684,N_158);
and U4705 (N_4705,N_1148,N_2652);
or U4706 (N_4706,N_2267,N_1192);
or U4707 (N_4707,N_1208,N_2855);
and U4708 (N_4708,N_929,N_243);
nand U4709 (N_4709,N_2654,N_2346);
and U4710 (N_4710,N_2729,N_2762);
and U4711 (N_4711,N_1596,N_2078);
xnor U4712 (N_4712,N_2915,N_1140);
and U4713 (N_4713,N_2101,N_2047);
nand U4714 (N_4714,N_479,N_1674);
xnor U4715 (N_4715,N_1961,N_1035);
nand U4716 (N_4716,N_1443,N_1532);
xor U4717 (N_4717,N_1003,N_1926);
or U4718 (N_4718,N_1046,N_787);
xnor U4719 (N_4719,N_50,N_1207);
nand U4720 (N_4720,N_696,N_444);
and U4721 (N_4721,N_1284,N_2042);
or U4722 (N_4722,N_2444,N_1748);
nor U4723 (N_4723,N_244,N_2563);
nor U4724 (N_4724,N_2001,N_767);
nand U4725 (N_4725,N_116,N_1542);
nor U4726 (N_4726,N_1179,N_1681);
nand U4727 (N_4727,N_3064,N_2676);
nand U4728 (N_4728,N_1074,N_1444);
nor U4729 (N_4729,N_188,N_2040);
nor U4730 (N_4730,N_314,N_2507);
or U4731 (N_4731,N_1612,N_2130);
and U4732 (N_4732,N_160,N_317);
nand U4733 (N_4733,N_727,N_1891);
and U4734 (N_4734,N_2467,N_90);
and U4735 (N_4735,N_1738,N_2067);
xor U4736 (N_4736,N_358,N_2966);
nand U4737 (N_4737,N_1339,N_146);
nor U4738 (N_4738,N_2216,N_2169);
nor U4739 (N_4739,N_934,N_2254);
or U4740 (N_4740,N_291,N_3001);
nand U4741 (N_4741,N_1208,N_2372);
xor U4742 (N_4742,N_955,N_154);
or U4743 (N_4743,N_1205,N_2908);
nand U4744 (N_4744,N_1902,N_512);
xnor U4745 (N_4745,N_1880,N_2159);
and U4746 (N_4746,N_96,N_783);
nor U4747 (N_4747,N_1802,N_1926);
xnor U4748 (N_4748,N_2939,N_434);
nand U4749 (N_4749,N_946,N_2276);
nor U4750 (N_4750,N_1317,N_683);
or U4751 (N_4751,N_998,N_326);
xnor U4752 (N_4752,N_920,N_2005);
or U4753 (N_4753,N_1263,N_2224);
or U4754 (N_4754,N_1154,N_2383);
and U4755 (N_4755,N_3010,N_1671);
nor U4756 (N_4756,N_197,N_2151);
and U4757 (N_4757,N_2605,N_2287);
and U4758 (N_4758,N_2261,N_500);
nand U4759 (N_4759,N_397,N_1690);
or U4760 (N_4760,N_2727,N_1481);
or U4761 (N_4761,N_2667,N_2432);
xnor U4762 (N_4762,N_1962,N_2356);
nor U4763 (N_4763,N_288,N_1853);
nand U4764 (N_4764,N_956,N_2499);
xnor U4765 (N_4765,N_785,N_174);
and U4766 (N_4766,N_0,N_543);
or U4767 (N_4767,N_1152,N_1961);
nand U4768 (N_4768,N_571,N_2866);
nand U4769 (N_4769,N_1291,N_384);
nand U4770 (N_4770,N_731,N_2280);
or U4771 (N_4771,N_2345,N_2515);
and U4772 (N_4772,N_2336,N_1991);
nor U4773 (N_4773,N_1358,N_2359);
xnor U4774 (N_4774,N_1136,N_696);
nand U4775 (N_4775,N_1571,N_1449);
nand U4776 (N_4776,N_1557,N_2301);
nand U4777 (N_4777,N_2442,N_776);
nor U4778 (N_4778,N_1424,N_1637);
nor U4779 (N_4779,N_419,N_1452);
nand U4780 (N_4780,N_822,N_2776);
and U4781 (N_4781,N_246,N_2095);
and U4782 (N_4782,N_2394,N_2954);
nor U4783 (N_4783,N_2024,N_671);
nor U4784 (N_4784,N_3095,N_2816);
and U4785 (N_4785,N_592,N_2);
nor U4786 (N_4786,N_1184,N_3109);
xnor U4787 (N_4787,N_366,N_1354);
and U4788 (N_4788,N_2704,N_200);
or U4789 (N_4789,N_2237,N_2380);
nor U4790 (N_4790,N_1280,N_868);
xnor U4791 (N_4791,N_2746,N_2832);
nor U4792 (N_4792,N_1373,N_650);
xor U4793 (N_4793,N_1345,N_2593);
and U4794 (N_4794,N_2969,N_1985);
or U4795 (N_4795,N_138,N_1783);
nand U4796 (N_4796,N_3114,N_1388);
and U4797 (N_4797,N_2697,N_2489);
and U4798 (N_4798,N_306,N_1166);
nand U4799 (N_4799,N_2995,N_2788);
xor U4800 (N_4800,N_2255,N_238);
nor U4801 (N_4801,N_1752,N_2446);
or U4802 (N_4802,N_1570,N_1145);
and U4803 (N_4803,N_1875,N_2023);
or U4804 (N_4804,N_538,N_1180);
or U4805 (N_4805,N_1845,N_2);
xnor U4806 (N_4806,N_2573,N_2962);
or U4807 (N_4807,N_1429,N_146);
xnor U4808 (N_4808,N_60,N_3098);
nand U4809 (N_4809,N_1742,N_2742);
nor U4810 (N_4810,N_894,N_559);
or U4811 (N_4811,N_53,N_1906);
and U4812 (N_4812,N_569,N_1466);
nor U4813 (N_4813,N_2365,N_1815);
and U4814 (N_4814,N_1371,N_305);
xor U4815 (N_4815,N_1311,N_1201);
nand U4816 (N_4816,N_537,N_3033);
or U4817 (N_4817,N_349,N_341);
or U4818 (N_4818,N_1278,N_1647);
and U4819 (N_4819,N_1500,N_468);
xor U4820 (N_4820,N_399,N_761);
xnor U4821 (N_4821,N_2513,N_1322);
nand U4822 (N_4822,N_2120,N_399);
and U4823 (N_4823,N_1587,N_1231);
xor U4824 (N_4824,N_2969,N_2223);
or U4825 (N_4825,N_12,N_2706);
xor U4826 (N_4826,N_1748,N_1771);
nand U4827 (N_4827,N_1620,N_2276);
nor U4828 (N_4828,N_1502,N_1040);
and U4829 (N_4829,N_1637,N_783);
and U4830 (N_4830,N_1935,N_1939);
nand U4831 (N_4831,N_1769,N_1228);
nand U4832 (N_4832,N_2856,N_1690);
nor U4833 (N_4833,N_2100,N_2401);
xnor U4834 (N_4834,N_2442,N_33);
nand U4835 (N_4835,N_2876,N_2594);
and U4836 (N_4836,N_1385,N_2061);
xor U4837 (N_4837,N_15,N_655);
or U4838 (N_4838,N_377,N_978);
or U4839 (N_4839,N_2117,N_1150);
nor U4840 (N_4840,N_7,N_2875);
nand U4841 (N_4841,N_1225,N_2639);
and U4842 (N_4842,N_2307,N_2738);
nor U4843 (N_4843,N_184,N_2306);
nor U4844 (N_4844,N_428,N_1250);
nor U4845 (N_4845,N_165,N_224);
nor U4846 (N_4846,N_2159,N_2390);
or U4847 (N_4847,N_390,N_1794);
xnor U4848 (N_4848,N_1382,N_1423);
nand U4849 (N_4849,N_1602,N_327);
nor U4850 (N_4850,N_880,N_2060);
xnor U4851 (N_4851,N_611,N_664);
xnor U4852 (N_4852,N_2646,N_434);
xnor U4853 (N_4853,N_2820,N_438);
nand U4854 (N_4854,N_1662,N_2789);
nand U4855 (N_4855,N_2068,N_1353);
or U4856 (N_4856,N_2477,N_2733);
and U4857 (N_4857,N_2187,N_154);
nor U4858 (N_4858,N_1130,N_1190);
and U4859 (N_4859,N_882,N_74);
nand U4860 (N_4860,N_2041,N_1987);
nor U4861 (N_4861,N_2220,N_958);
xnor U4862 (N_4862,N_1586,N_1398);
nand U4863 (N_4863,N_1291,N_2940);
and U4864 (N_4864,N_2259,N_464);
nor U4865 (N_4865,N_1422,N_761);
xnor U4866 (N_4866,N_2527,N_252);
and U4867 (N_4867,N_2212,N_1945);
nand U4868 (N_4868,N_1667,N_155);
nand U4869 (N_4869,N_1996,N_1357);
nor U4870 (N_4870,N_1849,N_951);
or U4871 (N_4871,N_2588,N_2225);
xor U4872 (N_4872,N_758,N_2);
or U4873 (N_4873,N_823,N_1867);
or U4874 (N_4874,N_1140,N_1872);
nor U4875 (N_4875,N_1183,N_593);
or U4876 (N_4876,N_61,N_1418);
nand U4877 (N_4877,N_340,N_1163);
nor U4878 (N_4878,N_1127,N_722);
xor U4879 (N_4879,N_1869,N_47);
nand U4880 (N_4880,N_462,N_1868);
or U4881 (N_4881,N_2522,N_1868);
nor U4882 (N_4882,N_183,N_207);
nor U4883 (N_4883,N_2022,N_2859);
and U4884 (N_4884,N_2381,N_2958);
nand U4885 (N_4885,N_841,N_835);
nand U4886 (N_4886,N_2127,N_2209);
xnor U4887 (N_4887,N_2379,N_1191);
xnor U4888 (N_4888,N_706,N_1908);
nor U4889 (N_4889,N_2814,N_1004);
nor U4890 (N_4890,N_1088,N_1320);
xor U4891 (N_4891,N_170,N_2619);
or U4892 (N_4892,N_1084,N_1378);
xor U4893 (N_4893,N_1685,N_1639);
nor U4894 (N_4894,N_1294,N_2882);
xnor U4895 (N_4895,N_419,N_2672);
and U4896 (N_4896,N_1693,N_2990);
nor U4897 (N_4897,N_1143,N_3069);
nand U4898 (N_4898,N_2567,N_2262);
and U4899 (N_4899,N_1847,N_2200);
or U4900 (N_4900,N_1913,N_2985);
or U4901 (N_4901,N_2181,N_1284);
xor U4902 (N_4902,N_1165,N_2308);
xnor U4903 (N_4903,N_2776,N_544);
nor U4904 (N_4904,N_341,N_1184);
nand U4905 (N_4905,N_3094,N_79);
xnor U4906 (N_4906,N_2871,N_1003);
nand U4907 (N_4907,N_1319,N_425);
nand U4908 (N_4908,N_267,N_626);
xnor U4909 (N_4909,N_1772,N_1424);
nand U4910 (N_4910,N_761,N_2432);
and U4911 (N_4911,N_158,N_555);
nand U4912 (N_4912,N_1652,N_2671);
and U4913 (N_4913,N_2293,N_1905);
nand U4914 (N_4914,N_1471,N_3114);
or U4915 (N_4915,N_1052,N_1068);
xor U4916 (N_4916,N_3062,N_1872);
and U4917 (N_4917,N_1539,N_2969);
nand U4918 (N_4918,N_2420,N_2994);
or U4919 (N_4919,N_1190,N_1919);
xnor U4920 (N_4920,N_2998,N_1070);
xor U4921 (N_4921,N_1480,N_1637);
nand U4922 (N_4922,N_2283,N_2873);
or U4923 (N_4923,N_1939,N_1100);
and U4924 (N_4924,N_503,N_1218);
or U4925 (N_4925,N_684,N_69);
xnor U4926 (N_4926,N_1664,N_1161);
and U4927 (N_4927,N_2618,N_2447);
xor U4928 (N_4928,N_2142,N_2169);
xor U4929 (N_4929,N_1531,N_2028);
nand U4930 (N_4930,N_324,N_2432);
xnor U4931 (N_4931,N_2605,N_1779);
nor U4932 (N_4932,N_570,N_1887);
nor U4933 (N_4933,N_1493,N_1485);
or U4934 (N_4934,N_2179,N_2215);
xnor U4935 (N_4935,N_1081,N_2141);
and U4936 (N_4936,N_1641,N_1643);
nor U4937 (N_4937,N_1031,N_800);
nand U4938 (N_4938,N_1244,N_256);
and U4939 (N_4939,N_2413,N_1790);
nor U4940 (N_4940,N_2109,N_1505);
and U4941 (N_4941,N_370,N_473);
and U4942 (N_4942,N_2512,N_1644);
nand U4943 (N_4943,N_2734,N_311);
nor U4944 (N_4944,N_2873,N_2145);
xor U4945 (N_4945,N_3006,N_1476);
or U4946 (N_4946,N_1578,N_500);
xor U4947 (N_4947,N_2633,N_2774);
and U4948 (N_4948,N_1539,N_1086);
xnor U4949 (N_4949,N_2911,N_2886);
nor U4950 (N_4950,N_135,N_733);
and U4951 (N_4951,N_1118,N_2858);
nor U4952 (N_4952,N_3062,N_1656);
or U4953 (N_4953,N_838,N_2905);
xnor U4954 (N_4954,N_2545,N_903);
xor U4955 (N_4955,N_1143,N_2765);
xnor U4956 (N_4956,N_2541,N_852);
xor U4957 (N_4957,N_806,N_71);
xnor U4958 (N_4958,N_1379,N_2609);
nor U4959 (N_4959,N_302,N_1216);
nand U4960 (N_4960,N_2867,N_2373);
nand U4961 (N_4961,N_517,N_1756);
nand U4962 (N_4962,N_2219,N_280);
or U4963 (N_4963,N_2548,N_1171);
and U4964 (N_4964,N_483,N_2290);
and U4965 (N_4965,N_1768,N_37);
nand U4966 (N_4966,N_1277,N_1329);
nor U4967 (N_4967,N_1181,N_28);
or U4968 (N_4968,N_137,N_574);
nor U4969 (N_4969,N_548,N_2069);
nor U4970 (N_4970,N_493,N_189);
nand U4971 (N_4971,N_269,N_786);
xnor U4972 (N_4972,N_620,N_1687);
or U4973 (N_4973,N_1968,N_2810);
or U4974 (N_4974,N_601,N_1572);
or U4975 (N_4975,N_1293,N_1054);
and U4976 (N_4976,N_1449,N_1168);
and U4977 (N_4977,N_1138,N_698);
or U4978 (N_4978,N_1109,N_509);
or U4979 (N_4979,N_422,N_314);
xnor U4980 (N_4980,N_3094,N_442);
xnor U4981 (N_4981,N_989,N_1902);
or U4982 (N_4982,N_1937,N_244);
nand U4983 (N_4983,N_1459,N_2492);
xnor U4984 (N_4984,N_1471,N_407);
or U4985 (N_4985,N_2847,N_181);
xor U4986 (N_4986,N_2506,N_3069);
and U4987 (N_4987,N_1235,N_309);
xor U4988 (N_4988,N_1284,N_3062);
nor U4989 (N_4989,N_1632,N_1735);
xor U4990 (N_4990,N_998,N_256);
and U4991 (N_4991,N_2350,N_693);
xnor U4992 (N_4992,N_2325,N_2054);
or U4993 (N_4993,N_220,N_2575);
xnor U4994 (N_4994,N_453,N_572);
or U4995 (N_4995,N_2130,N_2525);
nor U4996 (N_4996,N_1121,N_2174);
and U4997 (N_4997,N_1322,N_272);
nor U4998 (N_4998,N_2218,N_1177);
or U4999 (N_4999,N_1574,N_2287);
nand U5000 (N_5000,N_775,N_1800);
or U5001 (N_5001,N_1222,N_1243);
or U5002 (N_5002,N_1142,N_2972);
or U5003 (N_5003,N_1152,N_2563);
nand U5004 (N_5004,N_2404,N_2895);
xnor U5005 (N_5005,N_1129,N_3001);
nand U5006 (N_5006,N_2557,N_2463);
or U5007 (N_5007,N_2631,N_1020);
or U5008 (N_5008,N_848,N_418);
xnor U5009 (N_5009,N_2125,N_87);
and U5010 (N_5010,N_57,N_999);
or U5011 (N_5011,N_1933,N_2554);
nand U5012 (N_5012,N_1277,N_554);
or U5013 (N_5013,N_1216,N_2487);
or U5014 (N_5014,N_199,N_1271);
or U5015 (N_5015,N_1542,N_1978);
or U5016 (N_5016,N_377,N_1572);
nand U5017 (N_5017,N_734,N_1293);
xor U5018 (N_5018,N_2553,N_1122);
xor U5019 (N_5019,N_1309,N_1658);
nor U5020 (N_5020,N_2116,N_2348);
nor U5021 (N_5021,N_2497,N_2268);
and U5022 (N_5022,N_1839,N_1351);
nand U5023 (N_5023,N_1135,N_1235);
and U5024 (N_5024,N_1156,N_1998);
xor U5025 (N_5025,N_1196,N_2709);
nand U5026 (N_5026,N_2211,N_2468);
nor U5027 (N_5027,N_1935,N_1840);
or U5028 (N_5028,N_2195,N_422);
xor U5029 (N_5029,N_50,N_1627);
and U5030 (N_5030,N_496,N_1053);
or U5031 (N_5031,N_1738,N_769);
xor U5032 (N_5032,N_1411,N_1649);
nor U5033 (N_5033,N_90,N_2288);
nor U5034 (N_5034,N_1507,N_2071);
or U5035 (N_5035,N_2881,N_1041);
nor U5036 (N_5036,N_1543,N_1131);
xnor U5037 (N_5037,N_1348,N_422);
or U5038 (N_5038,N_1485,N_1434);
xnor U5039 (N_5039,N_2773,N_2073);
and U5040 (N_5040,N_2823,N_679);
nand U5041 (N_5041,N_980,N_1780);
or U5042 (N_5042,N_1621,N_2608);
xor U5043 (N_5043,N_1136,N_1045);
and U5044 (N_5044,N_1416,N_672);
nor U5045 (N_5045,N_2850,N_1503);
nor U5046 (N_5046,N_1461,N_2814);
xor U5047 (N_5047,N_2212,N_2022);
or U5048 (N_5048,N_2752,N_2051);
and U5049 (N_5049,N_2217,N_563);
or U5050 (N_5050,N_245,N_734);
and U5051 (N_5051,N_259,N_2143);
nand U5052 (N_5052,N_1419,N_1259);
nor U5053 (N_5053,N_2349,N_135);
nor U5054 (N_5054,N_2761,N_2092);
xor U5055 (N_5055,N_908,N_279);
nand U5056 (N_5056,N_2510,N_929);
nor U5057 (N_5057,N_1882,N_1291);
nand U5058 (N_5058,N_2049,N_1679);
or U5059 (N_5059,N_2183,N_1874);
xnor U5060 (N_5060,N_1408,N_1696);
nand U5061 (N_5061,N_2402,N_327);
nand U5062 (N_5062,N_1691,N_254);
or U5063 (N_5063,N_1220,N_2691);
xor U5064 (N_5064,N_2916,N_29);
or U5065 (N_5065,N_2064,N_1196);
nand U5066 (N_5066,N_1574,N_1209);
and U5067 (N_5067,N_2286,N_1090);
or U5068 (N_5068,N_935,N_1691);
nor U5069 (N_5069,N_237,N_864);
xnor U5070 (N_5070,N_14,N_924);
nor U5071 (N_5071,N_3075,N_2804);
and U5072 (N_5072,N_354,N_1281);
and U5073 (N_5073,N_636,N_2331);
nand U5074 (N_5074,N_1952,N_1739);
or U5075 (N_5075,N_285,N_2190);
xor U5076 (N_5076,N_1411,N_2912);
or U5077 (N_5077,N_1597,N_124);
nor U5078 (N_5078,N_2508,N_2410);
nand U5079 (N_5079,N_887,N_2739);
nand U5080 (N_5080,N_316,N_2115);
xor U5081 (N_5081,N_1807,N_3049);
and U5082 (N_5082,N_2287,N_854);
nor U5083 (N_5083,N_1233,N_2064);
xnor U5084 (N_5084,N_627,N_1823);
nor U5085 (N_5085,N_596,N_604);
or U5086 (N_5086,N_2134,N_2871);
nand U5087 (N_5087,N_1304,N_542);
nor U5088 (N_5088,N_1032,N_1955);
nor U5089 (N_5089,N_1730,N_769);
and U5090 (N_5090,N_1999,N_617);
and U5091 (N_5091,N_234,N_1421);
xnor U5092 (N_5092,N_1427,N_747);
or U5093 (N_5093,N_2590,N_2146);
nand U5094 (N_5094,N_675,N_2994);
nor U5095 (N_5095,N_344,N_1065);
and U5096 (N_5096,N_2755,N_579);
nor U5097 (N_5097,N_1265,N_1177);
nand U5098 (N_5098,N_1029,N_2385);
and U5099 (N_5099,N_2898,N_1839);
and U5100 (N_5100,N_324,N_656);
and U5101 (N_5101,N_194,N_767);
xor U5102 (N_5102,N_2175,N_2274);
nor U5103 (N_5103,N_28,N_3081);
xnor U5104 (N_5104,N_454,N_2163);
nor U5105 (N_5105,N_230,N_2549);
and U5106 (N_5106,N_2878,N_1702);
nand U5107 (N_5107,N_1400,N_216);
or U5108 (N_5108,N_159,N_2779);
nor U5109 (N_5109,N_1272,N_2103);
and U5110 (N_5110,N_1168,N_1525);
and U5111 (N_5111,N_2510,N_235);
nor U5112 (N_5112,N_837,N_2499);
nand U5113 (N_5113,N_2138,N_2735);
and U5114 (N_5114,N_211,N_184);
or U5115 (N_5115,N_2815,N_2450);
xnor U5116 (N_5116,N_2855,N_1615);
or U5117 (N_5117,N_1061,N_2032);
xnor U5118 (N_5118,N_2978,N_1178);
nand U5119 (N_5119,N_2101,N_1089);
nand U5120 (N_5120,N_1832,N_295);
nor U5121 (N_5121,N_923,N_2277);
and U5122 (N_5122,N_257,N_919);
and U5123 (N_5123,N_634,N_1534);
xor U5124 (N_5124,N_421,N_2555);
nand U5125 (N_5125,N_2228,N_1603);
or U5126 (N_5126,N_1621,N_870);
nor U5127 (N_5127,N_1499,N_2691);
nor U5128 (N_5128,N_1469,N_1048);
or U5129 (N_5129,N_1878,N_1271);
nand U5130 (N_5130,N_2581,N_2972);
nor U5131 (N_5131,N_2890,N_2745);
xor U5132 (N_5132,N_1586,N_2119);
and U5133 (N_5133,N_753,N_2500);
xnor U5134 (N_5134,N_1220,N_793);
nand U5135 (N_5135,N_2881,N_2851);
nand U5136 (N_5136,N_2716,N_98);
nand U5137 (N_5137,N_457,N_2594);
and U5138 (N_5138,N_1832,N_562);
and U5139 (N_5139,N_2568,N_1464);
nor U5140 (N_5140,N_2851,N_1990);
nand U5141 (N_5141,N_1559,N_199);
or U5142 (N_5142,N_2832,N_1600);
xnor U5143 (N_5143,N_2065,N_1728);
nor U5144 (N_5144,N_2221,N_299);
or U5145 (N_5145,N_1946,N_1855);
and U5146 (N_5146,N_167,N_2227);
nor U5147 (N_5147,N_973,N_711);
xnor U5148 (N_5148,N_965,N_346);
or U5149 (N_5149,N_557,N_489);
or U5150 (N_5150,N_2303,N_2775);
and U5151 (N_5151,N_1722,N_102);
and U5152 (N_5152,N_269,N_1005);
or U5153 (N_5153,N_2427,N_1419);
xnor U5154 (N_5154,N_488,N_1701);
xnor U5155 (N_5155,N_2226,N_356);
nand U5156 (N_5156,N_2250,N_1979);
nor U5157 (N_5157,N_1132,N_74);
nand U5158 (N_5158,N_2853,N_2594);
nand U5159 (N_5159,N_1165,N_2519);
xor U5160 (N_5160,N_2656,N_412);
or U5161 (N_5161,N_1771,N_2681);
or U5162 (N_5162,N_2458,N_2018);
nor U5163 (N_5163,N_2630,N_455);
xor U5164 (N_5164,N_1707,N_2723);
nor U5165 (N_5165,N_2404,N_2134);
or U5166 (N_5166,N_2643,N_595);
nand U5167 (N_5167,N_2099,N_1120);
xor U5168 (N_5168,N_2605,N_856);
nand U5169 (N_5169,N_3093,N_2785);
nor U5170 (N_5170,N_2202,N_3110);
nand U5171 (N_5171,N_2738,N_3085);
nor U5172 (N_5172,N_1805,N_2609);
and U5173 (N_5173,N_1060,N_875);
and U5174 (N_5174,N_2620,N_1557);
and U5175 (N_5175,N_1998,N_2194);
or U5176 (N_5176,N_2032,N_1914);
nor U5177 (N_5177,N_2289,N_2696);
nand U5178 (N_5178,N_218,N_2721);
or U5179 (N_5179,N_2650,N_177);
nand U5180 (N_5180,N_674,N_2047);
nand U5181 (N_5181,N_2070,N_2414);
nand U5182 (N_5182,N_2018,N_1056);
and U5183 (N_5183,N_2400,N_1659);
xnor U5184 (N_5184,N_2118,N_2396);
and U5185 (N_5185,N_1758,N_2030);
nand U5186 (N_5186,N_1151,N_2302);
nor U5187 (N_5187,N_618,N_1767);
and U5188 (N_5188,N_1957,N_2321);
and U5189 (N_5189,N_59,N_830);
and U5190 (N_5190,N_619,N_2772);
nor U5191 (N_5191,N_2920,N_3055);
or U5192 (N_5192,N_2600,N_1661);
xor U5193 (N_5193,N_1208,N_2246);
nor U5194 (N_5194,N_587,N_140);
nor U5195 (N_5195,N_169,N_1692);
xor U5196 (N_5196,N_1202,N_934);
or U5197 (N_5197,N_2485,N_784);
nor U5198 (N_5198,N_3053,N_2387);
nor U5199 (N_5199,N_2653,N_405);
xor U5200 (N_5200,N_1876,N_1213);
nor U5201 (N_5201,N_356,N_1275);
or U5202 (N_5202,N_3115,N_2316);
xnor U5203 (N_5203,N_2703,N_2922);
nor U5204 (N_5204,N_1949,N_219);
nand U5205 (N_5205,N_1225,N_1705);
xor U5206 (N_5206,N_3013,N_842);
xor U5207 (N_5207,N_1803,N_219);
nand U5208 (N_5208,N_2117,N_977);
and U5209 (N_5209,N_82,N_2661);
and U5210 (N_5210,N_1724,N_207);
and U5211 (N_5211,N_2193,N_1899);
xor U5212 (N_5212,N_1163,N_2790);
and U5213 (N_5213,N_2949,N_901);
nand U5214 (N_5214,N_2840,N_1822);
and U5215 (N_5215,N_2697,N_1303);
and U5216 (N_5216,N_2176,N_2393);
nand U5217 (N_5217,N_1821,N_1184);
xnor U5218 (N_5218,N_1295,N_2796);
nor U5219 (N_5219,N_344,N_1379);
or U5220 (N_5220,N_1057,N_2797);
nor U5221 (N_5221,N_1079,N_1450);
nor U5222 (N_5222,N_618,N_2795);
nand U5223 (N_5223,N_921,N_2987);
xnor U5224 (N_5224,N_2703,N_840);
xnor U5225 (N_5225,N_2134,N_790);
nand U5226 (N_5226,N_1678,N_1758);
xor U5227 (N_5227,N_24,N_1767);
nor U5228 (N_5228,N_2535,N_2236);
and U5229 (N_5229,N_3028,N_2912);
nor U5230 (N_5230,N_309,N_2590);
nor U5231 (N_5231,N_2696,N_1096);
xor U5232 (N_5232,N_2014,N_2574);
or U5233 (N_5233,N_379,N_2214);
and U5234 (N_5234,N_1279,N_310);
nand U5235 (N_5235,N_1320,N_2255);
nor U5236 (N_5236,N_1337,N_428);
and U5237 (N_5237,N_1710,N_1574);
or U5238 (N_5238,N_360,N_2418);
or U5239 (N_5239,N_1532,N_877);
or U5240 (N_5240,N_2287,N_2325);
or U5241 (N_5241,N_2192,N_681);
nor U5242 (N_5242,N_1885,N_2434);
xor U5243 (N_5243,N_3011,N_1490);
xnor U5244 (N_5244,N_2036,N_1536);
xor U5245 (N_5245,N_243,N_167);
nor U5246 (N_5246,N_1222,N_18);
nand U5247 (N_5247,N_2660,N_1194);
xnor U5248 (N_5248,N_1852,N_1319);
nor U5249 (N_5249,N_686,N_120);
nand U5250 (N_5250,N_1183,N_2351);
and U5251 (N_5251,N_1864,N_956);
and U5252 (N_5252,N_1523,N_2147);
nor U5253 (N_5253,N_732,N_1894);
nand U5254 (N_5254,N_2808,N_1279);
nor U5255 (N_5255,N_2866,N_798);
and U5256 (N_5256,N_1611,N_2318);
nand U5257 (N_5257,N_2378,N_3112);
xnor U5258 (N_5258,N_1414,N_1754);
xor U5259 (N_5259,N_1466,N_1795);
and U5260 (N_5260,N_514,N_1401);
nand U5261 (N_5261,N_506,N_176);
nor U5262 (N_5262,N_1975,N_44);
nand U5263 (N_5263,N_2066,N_281);
and U5264 (N_5264,N_2978,N_1759);
or U5265 (N_5265,N_1856,N_2396);
and U5266 (N_5266,N_2158,N_2514);
or U5267 (N_5267,N_1950,N_1886);
nor U5268 (N_5268,N_1524,N_629);
or U5269 (N_5269,N_2662,N_1278);
xor U5270 (N_5270,N_580,N_1819);
nand U5271 (N_5271,N_2927,N_639);
nor U5272 (N_5272,N_341,N_3124);
nor U5273 (N_5273,N_2769,N_967);
nand U5274 (N_5274,N_1575,N_2402);
or U5275 (N_5275,N_776,N_797);
nor U5276 (N_5276,N_745,N_1271);
nand U5277 (N_5277,N_1824,N_2857);
nand U5278 (N_5278,N_1078,N_2817);
or U5279 (N_5279,N_447,N_542);
nand U5280 (N_5280,N_1223,N_549);
and U5281 (N_5281,N_946,N_1192);
xor U5282 (N_5282,N_146,N_2983);
xor U5283 (N_5283,N_641,N_355);
and U5284 (N_5284,N_2954,N_1806);
nand U5285 (N_5285,N_2604,N_640);
nor U5286 (N_5286,N_2540,N_837);
and U5287 (N_5287,N_607,N_1031);
or U5288 (N_5288,N_145,N_122);
nor U5289 (N_5289,N_1329,N_826);
or U5290 (N_5290,N_1450,N_1662);
and U5291 (N_5291,N_1662,N_478);
and U5292 (N_5292,N_720,N_1193);
and U5293 (N_5293,N_2958,N_1572);
and U5294 (N_5294,N_2477,N_2395);
or U5295 (N_5295,N_2822,N_2729);
or U5296 (N_5296,N_1891,N_1227);
and U5297 (N_5297,N_1932,N_61);
nand U5298 (N_5298,N_2852,N_1932);
nor U5299 (N_5299,N_1918,N_364);
nor U5300 (N_5300,N_1139,N_1576);
nand U5301 (N_5301,N_1518,N_281);
xnor U5302 (N_5302,N_2979,N_18);
nor U5303 (N_5303,N_2026,N_2970);
xnor U5304 (N_5304,N_2387,N_1463);
nand U5305 (N_5305,N_836,N_1149);
xor U5306 (N_5306,N_499,N_435);
nand U5307 (N_5307,N_1605,N_1533);
nor U5308 (N_5308,N_2764,N_2117);
nand U5309 (N_5309,N_2479,N_2078);
and U5310 (N_5310,N_2053,N_1081);
nand U5311 (N_5311,N_442,N_558);
nand U5312 (N_5312,N_2059,N_2174);
and U5313 (N_5313,N_339,N_2031);
and U5314 (N_5314,N_1064,N_2460);
xor U5315 (N_5315,N_1429,N_2783);
xor U5316 (N_5316,N_1747,N_995);
xnor U5317 (N_5317,N_1995,N_1530);
or U5318 (N_5318,N_1039,N_113);
and U5319 (N_5319,N_2554,N_1);
and U5320 (N_5320,N_2291,N_645);
or U5321 (N_5321,N_69,N_2468);
and U5322 (N_5322,N_1337,N_1768);
nor U5323 (N_5323,N_863,N_1554);
nor U5324 (N_5324,N_1249,N_2729);
nand U5325 (N_5325,N_301,N_308);
xor U5326 (N_5326,N_140,N_736);
xnor U5327 (N_5327,N_1553,N_1322);
and U5328 (N_5328,N_1839,N_1088);
or U5329 (N_5329,N_1302,N_285);
nand U5330 (N_5330,N_2272,N_713);
and U5331 (N_5331,N_2770,N_2719);
nor U5332 (N_5332,N_2045,N_2637);
xor U5333 (N_5333,N_2023,N_2665);
nand U5334 (N_5334,N_1033,N_2181);
nor U5335 (N_5335,N_2153,N_1665);
or U5336 (N_5336,N_2031,N_2050);
and U5337 (N_5337,N_2172,N_2551);
and U5338 (N_5338,N_1170,N_3077);
and U5339 (N_5339,N_1939,N_1056);
and U5340 (N_5340,N_1226,N_272);
xnor U5341 (N_5341,N_2302,N_1355);
and U5342 (N_5342,N_1586,N_2343);
nand U5343 (N_5343,N_644,N_468);
nor U5344 (N_5344,N_1310,N_2358);
xnor U5345 (N_5345,N_55,N_2811);
or U5346 (N_5346,N_2028,N_1180);
nand U5347 (N_5347,N_591,N_2137);
nand U5348 (N_5348,N_239,N_2521);
or U5349 (N_5349,N_1688,N_218);
xnor U5350 (N_5350,N_2697,N_2940);
nor U5351 (N_5351,N_1783,N_776);
and U5352 (N_5352,N_2202,N_2055);
nand U5353 (N_5353,N_2300,N_1053);
or U5354 (N_5354,N_1103,N_541);
nor U5355 (N_5355,N_841,N_380);
nand U5356 (N_5356,N_2506,N_1550);
xor U5357 (N_5357,N_883,N_1686);
xnor U5358 (N_5358,N_952,N_2028);
and U5359 (N_5359,N_1191,N_2123);
and U5360 (N_5360,N_2163,N_750);
and U5361 (N_5361,N_2362,N_651);
nand U5362 (N_5362,N_605,N_833);
and U5363 (N_5363,N_2003,N_2140);
and U5364 (N_5364,N_2817,N_209);
and U5365 (N_5365,N_2124,N_40);
or U5366 (N_5366,N_1696,N_942);
or U5367 (N_5367,N_1460,N_2861);
and U5368 (N_5368,N_357,N_1557);
or U5369 (N_5369,N_1414,N_352);
xor U5370 (N_5370,N_313,N_2234);
xnor U5371 (N_5371,N_383,N_2934);
nand U5372 (N_5372,N_2894,N_241);
and U5373 (N_5373,N_73,N_2986);
nor U5374 (N_5374,N_1955,N_2513);
or U5375 (N_5375,N_1614,N_1411);
and U5376 (N_5376,N_1076,N_2929);
or U5377 (N_5377,N_358,N_522);
nor U5378 (N_5378,N_2200,N_934);
or U5379 (N_5379,N_1965,N_368);
and U5380 (N_5380,N_906,N_1368);
nor U5381 (N_5381,N_2959,N_2833);
nand U5382 (N_5382,N_177,N_1924);
or U5383 (N_5383,N_2755,N_1158);
and U5384 (N_5384,N_1029,N_1515);
and U5385 (N_5385,N_2513,N_3100);
nor U5386 (N_5386,N_2857,N_2901);
nand U5387 (N_5387,N_192,N_2870);
or U5388 (N_5388,N_2074,N_2140);
or U5389 (N_5389,N_2342,N_1254);
xnor U5390 (N_5390,N_2198,N_2711);
nor U5391 (N_5391,N_785,N_2187);
nand U5392 (N_5392,N_1497,N_487);
or U5393 (N_5393,N_704,N_504);
nor U5394 (N_5394,N_1780,N_464);
xor U5395 (N_5395,N_2627,N_1923);
and U5396 (N_5396,N_2690,N_253);
nor U5397 (N_5397,N_2048,N_1126);
and U5398 (N_5398,N_2209,N_1993);
or U5399 (N_5399,N_2319,N_2955);
xor U5400 (N_5400,N_770,N_2011);
and U5401 (N_5401,N_1123,N_2671);
nand U5402 (N_5402,N_2997,N_332);
xnor U5403 (N_5403,N_443,N_267);
nor U5404 (N_5404,N_257,N_1758);
nand U5405 (N_5405,N_1532,N_2274);
nand U5406 (N_5406,N_33,N_49);
xnor U5407 (N_5407,N_316,N_1657);
and U5408 (N_5408,N_1318,N_2074);
nor U5409 (N_5409,N_1030,N_2514);
xor U5410 (N_5410,N_2666,N_2619);
nor U5411 (N_5411,N_75,N_22);
nand U5412 (N_5412,N_2496,N_2645);
nor U5413 (N_5413,N_3058,N_2378);
nor U5414 (N_5414,N_2465,N_1459);
or U5415 (N_5415,N_1002,N_1601);
nand U5416 (N_5416,N_765,N_3097);
xnor U5417 (N_5417,N_68,N_113);
and U5418 (N_5418,N_2119,N_557);
and U5419 (N_5419,N_1783,N_2039);
nor U5420 (N_5420,N_2403,N_2797);
and U5421 (N_5421,N_2654,N_14);
xnor U5422 (N_5422,N_678,N_2243);
xnor U5423 (N_5423,N_2728,N_1121);
nor U5424 (N_5424,N_1668,N_2801);
or U5425 (N_5425,N_186,N_692);
and U5426 (N_5426,N_2503,N_2634);
or U5427 (N_5427,N_2354,N_1242);
nor U5428 (N_5428,N_1551,N_1603);
or U5429 (N_5429,N_2786,N_1066);
or U5430 (N_5430,N_2215,N_1616);
or U5431 (N_5431,N_1084,N_216);
nor U5432 (N_5432,N_1753,N_217);
or U5433 (N_5433,N_1376,N_421);
xnor U5434 (N_5434,N_2687,N_3077);
nand U5435 (N_5435,N_2747,N_876);
nor U5436 (N_5436,N_470,N_1328);
or U5437 (N_5437,N_456,N_383);
nor U5438 (N_5438,N_2444,N_1384);
or U5439 (N_5439,N_923,N_2193);
xnor U5440 (N_5440,N_1685,N_2618);
or U5441 (N_5441,N_1969,N_630);
nand U5442 (N_5442,N_3043,N_955);
xnor U5443 (N_5443,N_2114,N_3027);
and U5444 (N_5444,N_1633,N_1536);
nor U5445 (N_5445,N_2249,N_2847);
and U5446 (N_5446,N_2259,N_2942);
xnor U5447 (N_5447,N_2188,N_3043);
or U5448 (N_5448,N_1215,N_771);
or U5449 (N_5449,N_1592,N_400);
nand U5450 (N_5450,N_613,N_1624);
nor U5451 (N_5451,N_1832,N_369);
xnor U5452 (N_5452,N_800,N_2750);
and U5453 (N_5453,N_1930,N_561);
or U5454 (N_5454,N_2390,N_2222);
xnor U5455 (N_5455,N_1144,N_2423);
or U5456 (N_5456,N_3037,N_2153);
xor U5457 (N_5457,N_1621,N_256);
or U5458 (N_5458,N_2194,N_1230);
nor U5459 (N_5459,N_767,N_2988);
nor U5460 (N_5460,N_1790,N_2970);
or U5461 (N_5461,N_1406,N_3044);
nand U5462 (N_5462,N_1116,N_665);
and U5463 (N_5463,N_2062,N_2521);
or U5464 (N_5464,N_1258,N_2813);
nor U5465 (N_5465,N_2251,N_1833);
nor U5466 (N_5466,N_2666,N_2564);
nor U5467 (N_5467,N_566,N_842);
or U5468 (N_5468,N_2736,N_511);
or U5469 (N_5469,N_1117,N_2648);
nand U5470 (N_5470,N_2839,N_1670);
or U5471 (N_5471,N_1560,N_496);
and U5472 (N_5472,N_2836,N_2572);
nand U5473 (N_5473,N_2984,N_610);
nand U5474 (N_5474,N_770,N_2171);
xor U5475 (N_5475,N_369,N_2043);
xnor U5476 (N_5476,N_2231,N_1089);
and U5477 (N_5477,N_2905,N_292);
nand U5478 (N_5478,N_2866,N_1659);
nor U5479 (N_5479,N_816,N_2862);
or U5480 (N_5480,N_1382,N_1705);
and U5481 (N_5481,N_390,N_2627);
or U5482 (N_5482,N_2513,N_345);
xor U5483 (N_5483,N_1329,N_1002);
or U5484 (N_5484,N_556,N_2897);
xnor U5485 (N_5485,N_1121,N_2925);
or U5486 (N_5486,N_1247,N_2790);
nand U5487 (N_5487,N_2487,N_979);
and U5488 (N_5488,N_1515,N_172);
nand U5489 (N_5489,N_1354,N_492);
and U5490 (N_5490,N_1734,N_457);
nand U5491 (N_5491,N_2650,N_162);
xnor U5492 (N_5492,N_1885,N_806);
nor U5493 (N_5493,N_1847,N_2053);
xor U5494 (N_5494,N_2869,N_1807);
and U5495 (N_5495,N_2985,N_14);
or U5496 (N_5496,N_2595,N_2896);
xor U5497 (N_5497,N_521,N_1889);
nand U5498 (N_5498,N_1643,N_249);
or U5499 (N_5499,N_1702,N_1922);
nand U5500 (N_5500,N_2367,N_1858);
nor U5501 (N_5501,N_29,N_1550);
nor U5502 (N_5502,N_737,N_2615);
nand U5503 (N_5503,N_1124,N_99);
nand U5504 (N_5504,N_2814,N_1357);
nor U5505 (N_5505,N_1632,N_2291);
nand U5506 (N_5506,N_415,N_102);
and U5507 (N_5507,N_2937,N_1274);
xnor U5508 (N_5508,N_1657,N_2896);
nand U5509 (N_5509,N_952,N_204);
nand U5510 (N_5510,N_577,N_1724);
nand U5511 (N_5511,N_836,N_2259);
or U5512 (N_5512,N_1810,N_265);
and U5513 (N_5513,N_1105,N_2018);
or U5514 (N_5514,N_992,N_457);
nand U5515 (N_5515,N_377,N_2147);
and U5516 (N_5516,N_1486,N_661);
and U5517 (N_5517,N_213,N_570);
xor U5518 (N_5518,N_1562,N_691);
and U5519 (N_5519,N_2836,N_827);
or U5520 (N_5520,N_896,N_2353);
nor U5521 (N_5521,N_2904,N_2199);
nor U5522 (N_5522,N_1777,N_1920);
nor U5523 (N_5523,N_2094,N_359);
nor U5524 (N_5524,N_1584,N_1437);
nand U5525 (N_5525,N_143,N_926);
and U5526 (N_5526,N_102,N_2707);
nor U5527 (N_5527,N_792,N_2886);
xnor U5528 (N_5528,N_427,N_831);
and U5529 (N_5529,N_1202,N_2947);
and U5530 (N_5530,N_1530,N_2036);
and U5531 (N_5531,N_638,N_1507);
or U5532 (N_5532,N_1540,N_972);
nor U5533 (N_5533,N_1649,N_740);
and U5534 (N_5534,N_3124,N_1646);
and U5535 (N_5535,N_1728,N_1002);
nand U5536 (N_5536,N_3013,N_2897);
and U5537 (N_5537,N_1538,N_2532);
nor U5538 (N_5538,N_1837,N_1409);
nor U5539 (N_5539,N_1085,N_1079);
or U5540 (N_5540,N_3009,N_2449);
and U5541 (N_5541,N_1430,N_1561);
nor U5542 (N_5542,N_2425,N_913);
nor U5543 (N_5543,N_2144,N_2270);
and U5544 (N_5544,N_2107,N_228);
nor U5545 (N_5545,N_760,N_515);
xor U5546 (N_5546,N_350,N_1246);
nor U5547 (N_5547,N_2620,N_1842);
and U5548 (N_5548,N_277,N_1698);
nor U5549 (N_5549,N_2692,N_441);
nor U5550 (N_5550,N_1446,N_1750);
xnor U5551 (N_5551,N_1565,N_1239);
and U5552 (N_5552,N_1006,N_1362);
and U5553 (N_5553,N_2912,N_807);
nand U5554 (N_5554,N_490,N_2304);
xnor U5555 (N_5555,N_1735,N_171);
or U5556 (N_5556,N_173,N_2176);
and U5557 (N_5557,N_1939,N_3032);
and U5558 (N_5558,N_2676,N_2946);
nor U5559 (N_5559,N_1495,N_2334);
nor U5560 (N_5560,N_2046,N_1361);
xnor U5561 (N_5561,N_2440,N_22);
and U5562 (N_5562,N_42,N_2360);
or U5563 (N_5563,N_2282,N_996);
xor U5564 (N_5564,N_1517,N_1762);
or U5565 (N_5565,N_1267,N_1018);
or U5566 (N_5566,N_2494,N_2969);
nand U5567 (N_5567,N_2340,N_2816);
or U5568 (N_5568,N_2530,N_1658);
or U5569 (N_5569,N_534,N_1512);
nor U5570 (N_5570,N_2794,N_60);
and U5571 (N_5571,N_1791,N_2329);
nor U5572 (N_5572,N_1038,N_587);
nand U5573 (N_5573,N_2164,N_1295);
nand U5574 (N_5574,N_2572,N_2187);
nor U5575 (N_5575,N_2800,N_1540);
and U5576 (N_5576,N_1958,N_2155);
xor U5577 (N_5577,N_2299,N_430);
nor U5578 (N_5578,N_1998,N_1199);
or U5579 (N_5579,N_837,N_1274);
or U5580 (N_5580,N_1813,N_145);
nand U5581 (N_5581,N_2743,N_2054);
or U5582 (N_5582,N_2862,N_1327);
nand U5583 (N_5583,N_2597,N_1376);
or U5584 (N_5584,N_2496,N_2828);
or U5585 (N_5585,N_3044,N_2416);
or U5586 (N_5586,N_1103,N_1856);
nand U5587 (N_5587,N_186,N_1079);
and U5588 (N_5588,N_782,N_3023);
or U5589 (N_5589,N_1957,N_1712);
xnor U5590 (N_5590,N_1813,N_1315);
nor U5591 (N_5591,N_255,N_706);
xnor U5592 (N_5592,N_789,N_977);
nor U5593 (N_5593,N_1308,N_354);
nand U5594 (N_5594,N_2762,N_2428);
nand U5595 (N_5595,N_307,N_1225);
nand U5596 (N_5596,N_1011,N_170);
nand U5597 (N_5597,N_2983,N_3109);
xnor U5598 (N_5598,N_416,N_1820);
nand U5599 (N_5599,N_2244,N_994);
nor U5600 (N_5600,N_1532,N_1368);
xnor U5601 (N_5601,N_178,N_3069);
or U5602 (N_5602,N_240,N_1562);
and U5603 (N_5603,N_3027,N_1727);
and U5604 (N_5604,N_3034,N_2948);
and U5605 (N_5605,N_580,N_2225);
or U5606 (N_5606,N_2416,N_1339);
xor U5607 (N_5607,N_997,N_2805);
nor U5608 (N_5608,N_530,N_1253);
nor U5609 (N_5609,N_944,N_84);
xnor U5610 (N_5610,N_1023,N_1307);
and U5611 (N_5611,N_1034,N_2582);
nor U5612 (N_5612,N_1794,N_2283);
xor U5613 (N_5613,N_1559,N_1764);
nand U5614 (N_5614,N_1774,N_813);
nor U5615 (N_5615,N_2823,N_590);
and U5616 (N_5616,N_1774,N_1886);
and U5617 (N_5617,N_249,N_3037);
and U5618 (N_5618,N_178,N_1133);
and U5619 (N_5619,N_202,N_1340);
nand U5620 (N_5620,N_893,N_2568);
or U5621 (N_5621,N_3028,N_2987);
nor U5622 (N_5622,N_2103,N_2235);
or U5623 (N_5623,N_2883,N_2232);
xor U5624 (N_5624,N_2403,N_2740);
nor U5625 (N_5625,N_2810,N_2949);
nand U5626 (N_5626,N_2814,N_2653);
nand U5627 (N_5627,N_1225,N_2766);
xnor U5628 (N_5628,N_193,N_2841);
xor U5629 (N_5629,N_219,N_2866);
or U5630 (N_5630,N_23,N_1337);
and U5631 (N_5631,N_2605,N_1029);
or U5632 (N_5632,N_645,N_586);
xnor U5633 (N_5633,N_2305,N_87);
xor U5634 (N_5634,N_2665,N_750);
or U5635 (N_5635,N_2784,N_396);
nor U5636 (N_5636,N_1926,N_241);
or U5637 (N_5637,N_45,N_1624);
nand U5638 (N_5638,N_2600,N_185);
xor U5639 (N_5639,N_2946,N_1910);
and U5640 (N_5640,N_251,N_2896);
and U5641 (N_5641,N_635,N_1650);
and U5642 (N_5642,N_2423,N_3087);
xor U5643 (N_5643,N_1777,N_3095);
and U5644 (N_5644,N_2465,N_734);
nand U5645 (N_5645,N_336,N_559);
xnor U5646 (N_5646,N_3061,N_2840);
nand U5647 (N_5647,N_1961,N_2397);
nor U5648 (N_5648,N_160,N_2478);
xor U5649 (N_5649,N_1607,N_2070);
or U5650 (N_5650,N_964,N_2658);
and U5651 (N_5651,N_84,N_324);
xor U5652 (N_5652,N_705,N_42);
nor U5653 (N_5653,N_2466,N_1985);
xnor U5654 (N_5654,N_672,N_362);
nor U5655 (N_5655,N_2307,N_3053);
xor U5656 (N_5656,N_889,N_2021);
nor U5657 (N_5657,N_1381,N_1820);
and U5658 (N_5658,N_1020,N_2036);
and U5659 (N_5659,N_1642,N_1976);
xnor U5660 (N_5660,N_2871,N_534);
or U5661 (N_5661,N_2780,N_1344);
nand U5662 (N_5662,N_462,N_2995);
xnor U5663 (N_5663,N_184,N_447);
nand U5664 (N_5664,N_1419,N_509);
and U5665 (N_5665,N_2470,N_2304);
nor U5666 (N_5666,N_2142,N_2603);
nand U5667 (N_5667,N_2560,N_2128);
xor U5668 (N_5668,N_501,N_504);
xnor U5669 (N_5669,N_108,N_2792);
and U5670 (N_5670,N_51,N_760);
nand U5671 (N_5671,N_1491,N_902);
nor U5672 (N_5672,N_302,N_2180);
nand U5673 (N_5673,N_767,N_2066);
xor U5674 (N_5674,N_3022,N_2573);
or U5675 (N_5675,N_3057,N_1965);
or U5676 (N_5676,N_118,N_319);
nor U5677 (N_5677,N_460,N_2943);
nand U5678 (N_5678,N_2616,N_1165);
and U5679 (N_5679,N_3114,N_2892);
and U5680 (N_5680,N_2283,N_665);
nor U5681 (N_5681,N_1813,N_344);
xnor U5682 (N_5682,N_2868,N_180);
and U5683 (N_5683,N_2700,N_2864);
nand U5684 (N_5684,N_2754,N_2294);
and U5685 (N_5685,N_1278,N_93);
nor U5686 (N_5686,N_122,N_823);
or U5687 (N_5687,N_2986,N_920);
and U5688 (N_5688,N_1669,N_214);
or U5689 (N_5689,N_2509,N_2901);
nor U5690 (N_5690,N_304,N_1448);
nand U5691 (N_5691,N_2809,N_579);
xnor U5692 (N_5692,N_2260,N_1788);
or U5693 (N_5693,N_932,N_2265);
nor U5694 (N_5694,N_1276,N_2686);
nand U5695 (N_5695,N_1241,N_185);
or U5696 (N_5696,N_1146,N_990);
and U5697 (N_5697,N_1840,N_1836);
and U5698 (N_5698,N_2014,N_1303);
nand U5699 (N_5699,N_46,N_367);
or U5700 (N_5700,N_917,N_136);
or U5701 (N_5701,N_2241,N_497);
xnor U5702 (N_5702,N_1707,N_2215);
xor U5703 (N_5703,N_1074,N_2950);
nand U5704 (N_5704,N_2069,N_1288);
xor U5705 (N_5705,N_920,N_2482);
and U5706 (N_5706,N_447,N_2510);
nand U5707 (N_5707,N_438,N_495);
nor U5708 (N_5708,N_2936,N_1653);
or U5709 (N_5709,N_1941,N_1233);
nor U5710 (N_5710,N_1554,N_514);
and U5711 (N_5711,N_107,N_435);
or U5712 (N_5712,N_748,N_369);
nor U5713 (N_5713,N_2893,N_2111);
or U5714 (N_5714,N_448,N_2337);
nor U5715 (N_5715,N_726,N_625);
nand U5716 (N_5716,N_743,N_1632);
or U5717 (N_5717,N_421,N_24);
or U5718 (N_5718,N_899,N_464);
xor U5719 (N_5719,N_142,N_2339);
nor U5720 (N_5720,N_2628,N_2893);
nand U5721 (N_5721,N_1266,N_1143);
or U5722 (N_5722,N_955,N_22);
and U5723 (N_5723,N_2986,N_69);
nor U5724 (N_5724,N_1635,N_951);
xnor U5725 (N_5725,N_2939,N_1669);
or U5726 (N_5726,N_571,N_2900);
nor U5727 (N_5727,N_2812,N_1519);
and U5728 (N_5728,N_1433,N_692);
nor U5729 (N_5729,N_2699,N_718);
or U5730 (N_5730,N_1841,N_68);
xor U5731 (N_5731,N_1927,N_1785);
xor U5732 (N_5732,N_1329,N_1046);
xnor U5733 (N_5733,N_2812,N_442);
or U5734 (N_5734,N_1966,N_846);
nor U5735 (N_5735,N_2794,N_3052);
and U5736 (N_5736,N_1138,N_448);
or U5737 (N_5737,N_2614,N_453);
and U5738 (N_5738,N_1004,N_2841);
xnor U5739 (N_5739,N_282,N_367);
or U5740 (N_5740,N_3027,N_2347);
xor U5741 (N_5741,N_515,N_1434);
nand U5742 (N_5742,N_1543,N_1642);
nand U5743 (N_5743,N_2608,N_2374);
and U5744 (N_5744,N_2577,N_2007);
or U5745 (N_5745,N_2154,N_1876);
nor U5746 (N_5746,N_602,N_847);
nand U5747 (N_5747,N_98,N_1385);
and U5748 (N_5748,N_1398,N_743);
nor U5749 (N_5749,N_2322,N_1001);
nand U5750 (N_5750,N_7,N_2329);
and U5751 (N_5751,N_1667,N_795);
and U5752 (N_5752,N_3091,N_229);
and U5753 (N_5753,N_836,N_1013);
xor U5754 (N_5754,N_1373,N_2708);
nor U5755 (N_5755,N_1240,N_473);
nand U5756 (N_5756,N_226,N_1884);
or U5757 (N_5757,N_434,N_2472);
nand U5758 (N_5758,N_1291,N_2255);
nand U5759 (N_5759,N_1414,N_1774);
nand U5760 (N_5760,N_226,N_1056);
nor U5761 (N_5761,N_263,N_2529);
nor U5762 (N_5762,N_915,N_474);
nand U5763 (N_5763,N_697,N_1438);
and U5764 (N_5764,N_1156,N_1905);
nor U5765 (N_5765,N_2246,N_2416);
and U5766 (N_5766,N_1052,N_544);
xor U5767 (N_5767,N_2851,N_830);
nand U5768 (N_5768,N_2164,N_237);
nand U5769 (N_5769,N_2170,N_836);
xor U5770 (N_5770,N_1291,N_1607);
or U5771 (N_5771,N_2317,N_2405);
or U5772 (N_5772,N_2128,N_161);
and U5773 (N_5773,N_2273,N_3035);
xnor U5774 (N_5774,N_304,N_2078);
xor U5775 (N_5775,N_517,N_2337);
or U5776 (N_5776,N_1577,N_1757);
xnor U5777 (N_5777,N_2426,N_2123);
xnor U5778 (N_5778,N_533,N_18);
xnor U5779 (N_5779,N_1684,N_21);
nor U5780 (N_5780,N_278,N_1728);
xnor U5781 (N_5781,N_148,N_2998);
nand U5782 (N_5782,N_498,N_2648);
nor U5783 (N_5783,N_1970,N_1133);
nand U5784 (N_5784,N_185,N_912);
or U5785 (N_5785,N_571,N_752);
nor U5786 (N_5786,N_353,N_2608);
nand U5787 (N_5787,N_1096,N_1015);
and U5788 (N_5788,N_2778,N_2061);
and U5789 (N_5789,N_1902,N_762);
or U5790 (N_5790,N_229,N_1689);
and U5791 (N_5791,N_1641,N_1023);
nor U5792 (N_5792,N_2512,N_2375);
nand U5793 (N_5793,N_1522,N_560);
nor U5794 (N_5794,N_468,N_1284);
xor U5795 (N_5795,N_1435,N_573);
nor U5796 (N_5796,N_2230,N_766);
xor U5797 (N_5797,N_367,N_677);
and U5798 (N_5798,N_506,N_752);
nor U5799 (N_5799,N_1159,N_80);
xnor U5800 (N_5800,N_2952,N_1701);
nor U5801 (N_5801,N_2511,N_837);
nand U5802 (N_5802,N_685,N_3108);
or U5803 (N_5803,N_811,N_2695);
or U5804 (N_5804,N_2818,N_2148);
nand U5805 (N_5805,N_884,N_52);
and U5806 (N_5806,N_2609,N_1834);
or U5807 (N_5807,N_1424,N_2000);
nor U5808 (N_5808,N_1784,N_1918);
nand U5809 (N_5809,N_140,N_882);
xor U5810 (N_5810,N_2382,N_1649);
nand U5811 (N_5811,N_12,N_1089);
xor U5812 (N_5812,N_2924,N_3026);
xnor U5813 (N_5813,N_1901,N_1264);
nand U5814 (N_5814,N_1840,N_1203);
xnor U5815 (N_5815,N_1949,N_3007);
nand U5816 (N_5816,N_1758,N_2111);
or U5817 (N_5817,N_42,N_727);
nand U5818 (N_5818,N_1137,N_1937);
nor U5819 (N_5819,N_2267,N_1824);
nor U5820 (N_5820,N_507,N_1547);
nor U5821 (N_5821,N_512,N_2834);
or U5822 (N_5822,N_1483,N_1125);
nand U5823 (N_5823,N_3031,N_1149);
or U5824 (N_5824,N_325,N_985);
or U5825 (N_5825,N_2064,N_1621);
or U5826 (N_5826,N_1606,N_1636);
or U5827 (N_5827,N_2917,N_452);
nand U5828 (N_5828,N_313,N_2931);
and U5829 (N_5829,N_859,N_2301);
nand U5830 (N_5830,N_1086,N_1243);
xor U5831 (N_5831,N_1424,N_1357);
or U5832 (N_5832,N_1342,N_2051);
or U5833 (N_5833,N_710,N_321);
or U5834 (N_5834,N_2985,N_1755);
or U5835 (N_5835,N_2014,N_851);
and U5836 (N_5836,N_1368,N_1981);
or U5837 (N_5837,N_122,N_413);
or U5838 (N_5838,N_230,N_1668);
xnor U5839 (N_5839,N_2633,N_1080);
or U5840 (N_5840,N_3118,N_785);
or U5841 (N_5841,N_3016,N_523);
nand U5842 (N_5842,N_994,N_435);
nor U5843 (N_5843,N_2890,N_800);
nand U5844 (N_5844,N_1898,N_1989);
and U5845 (N_5845,N_1493,N_141);
and U5846 (N_5846,N_534,N_3049);
nor U5847 (N_5847,N_2425,N_676);
nor U5848 (N_5848,N_2133,N_1143);
nand U5849 (N_5849,N_2682,N_1043);
nor U5850 (N_5850,N_2611,N_2677);
nor U5851 (N_5851,N_2300,N_2825);
nand U5852 (N_5852,N_1416,N_76);
or U5853 (N_5853,N_2238,N_168);
and U5854 (N_5854,N_267,N_2959);
nor U5855 (N_5855,N_56,N_1045);
xor U5856 (N_5856,N_2525,N_2783);
and U5857 (N_5857,N_1839,N_1536);
or U5858 (N_5858,N_1110,N_143);
or U5859 (N_5859,N_2602,N_2546);
nor U5860 (N_5860,N_917,N_3062);
or U5861 (N_5861,N_3080,N_800);
or U5862 (N_5862,N_2386,N_1900);
and U5863 (N_5863,N_25,N_483);
or U5864 (N_5864,N_2028,N_25);
or U5865 (N_5865,N_485,N_1252);
or U5866 (N_5866,N_2960,N_651);
and U5867 (N_5867,N_767,N_1609);
xor U5868 (N_5868,N_2369,N_15);
xnor U5869 (N_5869,N_1180,N_37);
or U5870 (N_5870,N_3066,N_879);
nor U5871 (N_5871,N_2745,N_1322);
nor U5872 (N_5872,N_595,N_2570);
and U5873 (N_5873,N_1574,N_2079);
xnor U5874 (N_5874,N_2852,N_1722);
nand U5875 (N_5875,N_601,N_2483);
and U5876 (N_5876,N_2973,N_599);
or U5877 (N_5877,N_514,N_1654);
and U5878 (N_5878,N_1955,N_2872);
nand U5879 (N_5879,N_424,N_835);
nor U5880 (N_5880,N_363,N_2383);
and U5881 (N_5881,N_1411,N_2035);
or U5882 (N_5882,N_1050,N_680);
and U5883 (N_5883,N_656,N_2085);
nor U5884 (N_5884,N_1263,N_3084);
or U5885 (N_5885,N_147,N_2694);
and U5886 (N_5886,N_1034,N_413);
and U5887 (N_5887,N_1275,N_1985);
nand U5888 (N_5888,N_1033,N_2934);
or U5889 (N_5889,N_1117,N_1460);
and U5890 (N_5890,N_78,N_1852);
nor U5891 (N_5891,N_274,N_2424);
nand U5892 (N_5892,N_1442,N_1613);
or U5893 (N_5893,N_2281,N_2731);
or U5894 (N_5894,N_175,N_847);
xor U5895 (N_5895,N_1755,N_136);
nor U5896 (N_5896,N_1280,N_94);
nor U5897 (N_5897,N_2768,N_1146);
or U5898 (N_5898,N_2711,N_1672);
and U5899 (N_5899,N_2697,N_674);
nand U5900 (N_5900,N_2800,N_2304);
xor U5901 (N_5901,N_2296,N_587);
or U5902 (N_5902,N_1819,N_2178);
or U5903 (N_5903,N_2803,N_2139);
or U5904 (N_5904,N_2790,N_999);
or U5905 (N_5905,N_7,N_465);
and U5906 (N_5906,N_2873,N_113);
xor U5907 (N_5907,N_1148,N_1338);
or U5908 (N_5908,N_2503,N_483);
nand U5909 (N_5909,N_1235,N_3050);
nor U5910 (N_5910,N_1828,N_2135);
and U5911 (N_5911,N_40,N_1982);
nor U5912 (N_5912,N_2711,N_2120);
nor U5913 (N_5913,N_2425,N_1520);
and U5914 (N_5914,N_1461,N_2820);
nand U5915 (N_5915,N_1109,N_2527);
or U5916 (N_5916,N_417,N_550);
xnor U5917 (N_5917,N_1932,N_2800);
xnor U5918 (N_5918,N_1912,N_2511);
nand U5919 (N_5919,N_56,N_1510);
nor U5920 (N_5920,N_1173,N_1082);
and U5921 (N_5921,N_2414,N_606);
nand U5922 (N_5922,N_730,N_2883);
and U5923 (N_5923,N_1343,N_2132);
or U5924 (N_5924,N_230,N_1748);
or U5925 (N_5925,N_2036,N_206);
and U5926 (N_5926,N_1471,N_675);
nor U5927 (N_5927,N_40,N_1825);
or U5928 (N_5928,N_2907,N_2880);
and U5929 (N_5929,N_89,N_2927);
and U5930 (N_5930,N_663,N_2737);
and U5931 (N_5931,N_2676,N_3054);
nand U5932 (N_5932,N_2046,N_1137);
xnor U5933 (N_5933,N_1328,N_3123);
nor U5934 (N_5934,N_514,N_2657);
nor U5935 (N_5935,N_1699,N_2394);
nor U5936 (N_5936,N_2628,N_2746);
or U5937 (N_5937,N_2509,N_2720);
nor U5938 (N_5938,N_1529,N_2977);
or U5939 (N_5939,N_2932,N_1944);
xor U5940 (N_5940,N_188,N_3049);
nand U5941 (N_5941,N_2422,N_1701);
nor U5942 (N_5942,N_599,N_2842);
nand U5943 (N_5943,N_1730,N_240);
nand U5944 (N_5944,N_2035,N_1543);
xor U5945 (N_5945,N_1462,N_3021);
and U5946 (N_5946,N_3054,N_1956);
xnor U5947 (N_5947,N_2398,N_488);
xnor U5948 (N_5948,N_2244,N_1858);
or U5949 (N_5949,N_961,N_332);
and U5950 (N_5950,N_1398,N_1772);
nor U5951 (N_5951,N_509,N_2539);
nor U5952 (N_5952,N_1050,N_682);
nand U5953 (N_5953,N_518,N_942);
nor U5954 (N_5954,N_3054,N_243);
nand U5955 (N_5955,N_1830,N_1509);
and U5956 (N_5956,N_1889,N_104);
nor U5957 (N_5957,N_1839,N_2645);
nand U5958 (N_5958,N_85,N_2473);
and U5959 (N_5959,N_1841,N_2252);
or U5960 (N_5960,N_2092,N_783);
nand U5961 (N_5961,N_1023,N_3084);
nor U5962 (N_5962,N_1900,N_1125);
and U5963 (N_5963,N_1675,N_2340);
and U5964 (N_5964,N_2350,N_638);
xnor U5965 (N_5965,N_813,N_824);
xnor U5966 (N_5966,N_2546,N_2666);
or U5967 (N_5967,N_838,N_1132);
and U5968 (N_5968,N_2765,N_913);
xnor U5969 (N_5969,N_415,N_22);
xnor U5970 (N_5970,N_1019,N_607);
and U5971 (N_5971,N_1309,N_1337);
nor U5972 (N_5972,N_983,N_3081);
nand U5973 (N_5973,N_18,N_2574);
nor U5974 (N_5974,N_1961,N_730);
nor U5975 (N_5975,N_633,N_486);
or U5976 (N_5976,N_2381,N_805);
or U5977 (N_5977,N_3110,N_3047);
and U5978 (N_5978,N_309,N_1640);
xor U5979 (N_5979,N_2621,N_881);
xnor U5980 (N_5980,N_253,N_689);
nand U5981 (N_5981,N_873,N_2017);
xor U5982 (N_5982,N_768,N_3010);
xor U5983 (N_5983,N_1584,N_243);
or U5984 (N_5984,N_2181,N_2031);
xor U5985 (N_5985,N_2651,N_117);
xnor U5986 (N_5986,N_1984,N_464);
xnor U5987 (N_5987,N_1488,N_75);
xnor U5988 (N_5988,N_2803,N_1943);
or U5989 (N_5989,N_546,N_1188);
xnor U5990 (N_5990,N_132,N_2918);
nor U5991 (N_5991,N_2822,N_2714);
nand U5992 (N_5992,N_1503,N_1075);
nor U5993 (N_5993,N_380,N_574);
and U5994 (N_5994,N_2670,N_239);
and U5995 (N_5995,N_555,N_2986);
nor U5996 (N_5996,N_116,N_245);
nor U5997 (N_5997,N_1234,N_2669);
or U5998 (N_5998,N_1083,N_2272);
nor U5999 (N_5999,N_2909,N_2892);
nand U6000 (N_6000,N_635,N_1536);
or U6001 (N_6001,N_2116,N_355);
and U6002 (N_6002,N_989,N_2116);
xor U6003 (N_6003,N_813,N_3069);
or U6004 (N_6004,N_1824,N_116);
xor U6005 (N_6005,N_912,N_2050);
nor U6006 (N_6006,N_1047,N_2823);
xor U6007 (N_6007,N_1245,N_2868);
nor U6008 (N_6008,N_36,N_3042);
or U6009 (N_6009,N_1676,N_1843);
nor U6010 (N_6010,N_159,N_2630);
xor U6011 (N_6011,N_2350,N_3071);
nor U6012 (N_6012,N_2652,N_2117);
and U6013 (N_6013,N_1942,N_627);
and U6014 (N_6014,N_2939,N_267);
or U6015 (N_6015,N_1985,N_882);
or U6016 (N_6016,N_1803,N_71);
nor U6017 (N_6017,N_2242,N_1401);
xor U6018 (N_6018,N_1482,N_2525);
nand U6019 (N_6019,N_2888,N_412);
and U6020 (N_6020,N_1934,N_2954);
xor U6021 (N_6021,N_1407,N_1423);
and U6022 (N_6022,N_1979,N_2174);
xor U6023 (N_6023,N_138,N_1749);
or U6024 (N_6024,N_234,N_2354);
nand U6025 (N_6025,N_2260,N_170);
or U6026 (N_6026,N_858,N_561);
and U6027 (N_6027,N_1128,N_1427);
and U6028 (N_6028,N_2045,N_624);
nor U6029 (N_6029,N_1065,N_365);
xor U6030 (N_6030,N_8,N_2489);
xnor U6031 (N_6031,N_1124,N_1881);
nor U6032 (N_6032,N_1653,N_2303);
or U6033 (N_6033,N_1833,N_1553);
nand U6034 (N_6034,N_2981,N_118);
or U6035 (N_6035,N_1717,N_1986);
and U6036 (N_6036,N_1266,N_954);
nand U6037 (N_6037,N_413,N_95);
nand U6038 (N_6038,N_2782,N_2306);
nand U6039 (N_6039,N_2973,N_254);
nand U6040 (N_6040,N_912,N_2453);
xor U6041 (N_6041,N_1744,N_271);
nand U6042 (N_6042,N_1025,N_139);
xnor U6043 (N_6043,N_1337,N_981);
xor U6044 (N_6044,N_720,N_76);
nand U6045 (N_6045,N_157,N_1252);
nand U6046 (N_6046,N_2220,N_2910);
nor U6047 (N_6047,N_1109,N_495);
or U6048 (N_6048,N_1355,N_12);
nor U6049 (N_6049,N_1249,N_2606);
or U6050 (N_6050,N_1251,N_169);
or U6051 (N_6051,N_382,N_43);
and U6052 (N_6052,N_1776,N_829);
and U6053 (N_6053,N_2051,N_2352);
or U6054 (N_6054,N_177,N_1506);
or U6055 (N_6055,N_2594,N_506);
xor U6056 (N_6056,N_681,N_677);
nand U6057 (N_6057,N_2567,N_2119);
xnor U6058 (N_6058,N_563,N_1754);
and U6059 (N_6059,N_889,N_1900);
nand U6060 (N_6060,N_1536,N_2235);
and U6061 (N_6061,N_1329,N_3040);
or U6062 (N_6062,N_1175,N_2610);
and U6063 (N_6063,N_238,N_1043);
xnor U6064 (N_6064,N_325,N_1012);
nor U6065 (N_6065,N_123,N_2661);
nor U6066 (N_6066,N_1726,N_2023);
nor U6067 (N_6067,N_1309,N_3018);
nor U6068 (N_6068,N_2496,N_1181);
or U6069 (N_6069,N_2841,N_1213);
nand U6070 (N_6070,N_2620,N_1283);
or U6071 (N_6071,N_2371,N_999);
and U6072 (N_6072,N_1120,N_2171);
xnor U6073 (N_6073,N_1379,N_1928);
nand U6074 (N_6074,N_648,N_2922);
nor U6075 (N_6075,N_2534,N_1248);
and U6076 (N_6076,N_877,N_1085);
or U6077 (N_6077,N_873,N_1897);
nor U6078 (N_6078,N_1695,N_3119);
nor U6079 (N_6079,N_750,N_2329);
nand U6080 (N_6080,N_966,N_1537);
nor U6081 (N_6081,N_657,N_1680);
xor U6082 (N_6082,N_3104,N_2488);
and U6083 (N_6083,N_1046,N_2823);
and U6084 (N_6084,N_2000,N_1839);
nor U6085 (N_6085,N_1501,N_1555);
and U6086 (N_6086,N_2252,N_2289);
nand U6087 (N_6087,N_2855,N_892);
and U6088 (N_6088,N_366,N_327);
xor U6089 (N_6089,N_1740,N_1453);
and U6090 (N_6090,N_117,N_2206);
nand U6091 (N_6091,N_21,N_37);
or U6092 (N_6092,N_2066,N_2097);
or U6093 (N_6093,N_1427,N_2365);
or U6094 (N_6094,N_1154,N_1815);
nand U6095 (N_6095,N_1803,N_1120);
nor U6096 (N_6096,N_151,N_2559);
nand U6097 (N_6097,N_2287,N_884);
and U6098 (N_6098,N_1749,N_426);
or U6099 (N_6099,N_929,N_2627);
nand U6100 (N_6100,N_1364,N_271);
and U6101 (N_6101,N_868,N_1429);
and U6102 (N_6102,N_2833,N_1383);
xnor U6103 (N_6103,N_2973,N_784);
or U6104 (N_6104,N_2829,N_3021);
nor U6105 (N_6105,N_2362,N_1294);
or U6106 (N_6106,N_190,N_919);
nor U6107 (N_6107,N_580,N_2344);
xor U6108 (N_6108,N_747,N_2021);
xor U6109 (N_6109,N_1800,N_1137);
xor U6110 (N_6110,N_77,N_786);
xor U6111 (N_6111,N_664,N_1010);
and U6112 (N_6112,N_2616,N_2231);
xnor U6113 (N_6113,N_1752,N_163);
nor U6114 (N_6114,N_152,N_3075);
xor U6115 (N_6115,N_1228,N_2294);
or U6116 (N_6116,N_2530,N_16);
nand U6117 (N_6117,N_20,N_609);
or U6118 (N_6118,N_2799,N_2731);
xnor U6119 (N_6119,N_43,N_2633);
nand U6120 (N_6120,N_393,N_369);
nor U6121 (N_6121,N_2181,N_1819);
nor U6122 (N_6122,N_1339,N_981);
and U6123 (N_6123,N_1950,N_1717);
and U6124 (N_6124,N_1954,N_1691);
nand U6125 (N_6125,N_1363,N_1906);
or U6126 (N_6126,N_2920,N_2095);
and U6127 (N_6127,N_18,N_1474);
xnor U6128 (N_6128,N_2538,N_1834);
xnor U6129 (N_6129,N_2442,N_1727);
or U6130 (N_6130,N_2869,N_1181);
or U6131 (N_6131,N_865,N_2582);
or U6132 (N_6132,N_3096,N_1483);
and U6133 (N_6133,N_2283,N_19);
nand U6134 (N_6134,N_1077,N_221);
or U6135 (N_6135,N_3001,N_904);
and U6136 (N_6136,N_1794,N_97);
xor U6137 (N_6137,N_92,N_60);
xor U6138 (N_6138,N_382,N_1184);
and U6139 (N_6139,N_416,N_1954);
or U6140 (N_6140,N_780,N_2734);
xor U6141 (N_6141,N_1437,N_2681);
xnor U6142 (N_6142,N_1242,N_11);
and U6143 (N_6143,N_2314,N_3117);
and U6144 (N_6144,N_2185,N_496);
xor U6145 (N_6145,N_314,N_677);
and U6146 (N_6146,N_26,N_834);
and U6147 (N_6147,N_370,N_357);
nor U6148 (N_6148,N_2330,N_381);
or U6149 (N_6149,N_768,N_2888);
nor U6150 (N_6150,N_3055,N_1587);
and U6151 (N_6151,N_2149,N_2468);
nand U6152 (N_6152,N_2680,N_2708);
or U6153 (N_6153,N_2557,N_1837);
nand U6154 (N_6154,N_2388,N_1384);
or U6155 (N_6155,N_2690,N_2453);
nor U6156 (N_6156,N_1828,N_1279);
nor U6157 (N_6157,N_290,N_1186);
and U6158 (N_6158,N_1212,N_752);
or U6159 (N_6159,N_359,N_1986);
or U6160 (N_6160,N_2354,N_532);
nand U6161 (N_6161,N_919,N_2619);
or U6162 (N_6162,N_441,N_24);
and U6163 (N_6163,N_2706,N_2392);
and U6164 (N_6164,N_1017,N_1277);
xnor U6165 (N_6165,N_2509,N_2734);
xor U6166 (N_6166,N_2540,N_1383);
nor U6167 (N_6167,N_407,N_1932);
nand U6168 (N_6168,N_1682,N_335);
and U6169 (N_6169,N_184,N_173);
xor U6170 (N_6170,N_2329,N_3074);
nor U6171 (N_6171,N_1237,N_2599);
or U6172 (N_6172,N_2433,N_141);
and U6173 (N_6173,N_148,N_312);
and U6174 (N_6174,N_566,N_400);
xor U6175 (N_6175,N_1552,N_2036);
nand U6176 (N_6176,N_2907,N_1383);
nand U6177 (N_6177,N_2254,N_778);
or U6178 (N_6178,N_1034,N_1819);
nand U6179 (N_6179,N_236,N_62);
or U6180 (N_6180,N_176,N_968);
xor U6181 (N_6181,N_1900,N_617);
or U6182 (N_6182,N_2827,N_227);
or U6183 (N_6183,N_1197,N_2733);
xor U6184 (N_6184,N_1827,N_2829);
or U6185 (N_6185,N_1526,N_2009);
nand U6186 (N_6186,N_3109,N_1369);
xor U6187 (N_6187,N_2071,N_768);
nand U6188 (N_6188,N_1474,N_1898);
nor U6189 (N_6189,N_3122,N_364);
and U6190 (N_6190,N_1957,N_2092);
nand U6191 (N_6191,N_2828,N_2501);
nor U6192 (N_6192,N_2923,N_464);
xnor U6193 (N_6193,N_2402,N_2382);
nor U6194 (N_6194,N_2569,N_194);
xnor U6195 (N_6195,N_2003,N_2627);
nand U6196 (N_6196,N_2079,N_445);
and U6197 (N_6197,N_1469,N_2788);
nor U6198 (N_6198,N_608,N_60);
nand U6199 (N_6199,N_1276,N_759);
xor U6200 (N_6200,N_1976,N_109);
xor U6201 (N_6201,N_783,N_654);
nand U6202 (N_6202,N_432,N_2494);
or U6203 (N_6203,N_702,N_535);
nor U6204 (N_6204,N_2205,N_1610);
or U6205 (N_6205,N_2649,N_2310);
xnor U6206 (N_6206,N_2760,N_3022);
nor U6207 (N_6207,N_2397,N_2551);
and U6208 (N_6208,N_1457,N_296);
or U6209 (N_6209,N_1925,N_1197);
nor U6210 (N_6210,N_2805,N_1027);
nor U6211 (N_6211,N_981,N_2817);
nor U6212 (N_6212,N_2849,N_1976);
or U6213 (N_6213,N_3116,N_584);
xnor U6214 (N_6214,N_1715,N_947);
nand U6215 (N_6215,N_2212,N_1148);
and U6216 (N_6216,N_2218,N_1406);
xnor U6217 (N_6217,N_2879,N_1182);
or U6218 (N_6218,N_2073,N_649);
nand U6219 (N_6219,N_1964,N_1469);
or U6220 (N_6220,N_1469,N_1009);
xnor U6221 (N_6221,N_125,N_2185);
nand U6222 (N_6222,N_1688,N_1424);
nand U6223 (N_6223,N_751,N_2640);
xnor U6224 (N_6224,N_1775,N_1509);
or U6225 (N_6225,N_582,N_1567);
nand U6226 (N_6226,N_6,N_2175);
nor U6227 (N_6227,N_759,N_106);
or U6228 (N_6228,N_1328,N_2247);
nor U6229 (N_6229,N_2367,N_2216);
nor U6230 (N_6230,N_2560,N_1440);
nor U6231 (N_6231,N_2220,N_653);
nor U6232 (N_6232,N_2948,N_2697);
nand U6233 (N_6233,N_2199,N_507);
nor U6234 (N_6234,N_264,N_2291);
nand U6235 (N_6235,N_927,N_2071);
nand U6236 (N_6236,N_1899,N_1621);
or U6237 (N_6237,N_350,N_1170);
or U6238 (N_6238,N_587,N_1497);
nor U6239 (N_6239,N_1361,N_1850);
or U6240 (N_6240,N_2665,N_1770);
nand U6241 (N_6241,N_1491,N_2093);
nor U6242 (N_6242,N_1152,N_874);
xor U6243 (N_6243,N_1578,N_2777);
xnor U6244 (N_6244,N_2405,N_1984);
nand U6245 (N_6245,N_622,N_2867);
nor U6246 (N_6246,N_436,N_2057);
and U6247 (N_6247,N_1732,N_2403);
or U6248 (N_6248,N_1833,N_1929);
nor U6249 (N_6249,N_1192,N_900);
nor U6250 (N_6250,N_5890,N_3464);
xor U6251 (N_6251,N_6193,N_3970);
xor U6252 (N_6252,N_6148,N_4338);
nor U6253 (N_6253,N_3597,N_3956);
nor U6254 (N_6254,N_5512,N_4327);
or U6255 (N_6255,N_5760,N_5852);
nand U6256 (N_6256,N_5561,N_4901);
and U6257 (N_6257,N_4244,N_3548);
or U6258 (N_6258,N_4121,N_3552);
and U6259 (N_6259,N_5099,N_4020);
nand U6260 (N_6260,N_3163,N_5148);
or U6261 (N_6261,N_4213,N_4273);
xnor U6262 (N_6262,N_5865,N_4237);
or U6263 (N_6263,N_5984,N_4366);
nor U6264 (N_6264,N_5569,N_3647);
xnor U6265 (N_6265,N_5291,N_5572);
xnor U6266 (N_6266,N_3499,N_5018);
xnor U6267 (N_6267,N_3798,N_3431);
nand U6268 (N_6268,N_5767,N_3869);
or U6269 (N_6269,N_6137,N_5120);
and U6270 (N_6270,N_4629,N_3878);
and U6271 (N_6271,N_3158,N_3157);
nor U6272 (N_6272,N_3831,N_6054);
xnor U6273 (N_6273,N_4181,N_4625);
and U6274 (N_6274,N_3215,N_3188);
nor U6275 (N_6275,N_3770,N_3493);
xnor U6276 (N_6276,N_3489,N_5769);
nand U6277 (N_6277,N_6123,N_3361);
or U6278 (N_6278,N_4240,N_3775);
xor U6279 (N_6279,N_6026,N_3646);
nor U6280 (N_6280,N_6167,N_4175);
nand U6281 (N_6281,N_3717,N_5160);
or U6282 (N_6282,N_4365,N_3708);
nor U6283 (N_6283,N_6049,N_5388);
nand U6284 (N_6284,N_4420,N_3274);
xnor U6285 (N_6285,N_4956,N_5960);
or U6286 (N_6286,N_4130,N_5445);
nand U6287 (N_6287,N_5700,N_5834);
nor U6288 (N_6288,N_5024,N_3253);
xor U6289 (N_6289,N_3758,N_4569);
xnor U6290 (N_6290,N_5458,N_5638);
nor U6291 (N_6291,N_5823,N_3351);
and U6292 (N_6292,N_5224,N_5434);
xnor U6293 (N_6293,N_6055,N_5393);
xnor U6294 (N_6294,N_3306,N_3425);
nor U6295 (N_6295,N_3655,N_5109);
nor U6296 (N_6296,N_5545,N_4056);
nor U6297 (N_6297,N_4634,N_5106);
nand U6298 (N_6298,N_3358,N_4219);
and U6299 (N_6299,N_4789,N_4941);
xnor U6300 (N_6300,N_4149,N_5176);
or U6301 (N_6301,N_3964,N_6012);
xor U6302 (N_6302,N_5350,N_3266);
nor U6303 (N_6303,N_5399,N_5808);
xnor U6304 (N_6304,N_3927,N_5802);
and U6305 (N_6305,N_5619,N_6128);
and U6306 (N_6306,N_4844,N_4387);
xnor U6307 (N_6307,N_4684,N_4484);
and U6308 (N_6308,N_3461,N_5617);
or U6309 (N_6309,N_5085,N_5990);
nor U6310 (N_6310,N_5908,N_4514);
nor U6311 (N_6311,N_6221,N_5416);
xor U6312 (N_6312,N_5341,N_5989);
xor U6313 (N_6313,N_5365,N_4544);
nand U6314 (N_6314,N_6130,N_6230);
nor U6315 (N_6315,N_3901,N_4057);
or U6316 (N_6316,N_3560,N_4722);
and U6317 (N_6317,N_5742,N_4876);
xor U6318 (N_6318,N_4389,N_5433);
and U6319 (N_6319,N_3214,N_6249);
and U6320 (N_6320,N_3134,N_5052);
and U6321 (N_6321,N_5666,N_5389);
and U6322 (N_6322,N_6206,N_3734);
xor U6323 (N_6323,N_5415,N_5611);
and U6324 (N_6324,N_6182,N_4969);
nand U6325 (N_6325,N_4934,N_6090);
xnor U6326 (N_6326,N_6170,N_4643);
and U6327 (N_6327,N_4803,N_3935);
and U6328 (N_6328,N_5845,N_3842);
xor U6329 (N_6329,N_4356,N_4177);
or U6330 (N_6330,N_5849,N_4767);
xor U6331 (N_6331,N_4314,N_5750);
or U6332 (N_6332,N_3514,N_4352);
or U6333 (N_6333,N_4779,N_3380);
nand U6334 (N_6334,N_4704,N_5991);
or U6335 (N_6335,N_4670,N_4041);
nor U6336 (N_6336,N_3776,N_4978);
and U6337 (N_6337,N_6073,N_4375);
nor U6338 (N_6338,N_5038,N_3558);
nor U6339 (N_6339,N_5154,N_4695);
or U6340 (N_6340,N_4716,N_3382);
or U6341 (N_6341,N_5609,N_4824);
or U6342 (N_6342,N_4033,N_5161);
xor U6343 (N_6343,N_5999,N_3246);
and U6344 (N_6344,N_5735,N_4842);
xnor U6345 (N_6345,N_5444,N_6025);
nor U6346 (N_6346,N_5368,N_5044);
nor U6347 (N_6347,N_5843,N_3572);
nand U6348 (N_6348,N_3746,N_4667);
xor U6349 (N_6349,N_3581,N_5352);
or U6350 (N_6350,N_6177,N_4432);
nor U6351 (N_6351,N_4720,N_3853);
and U6352 (N_6352,N_5199,N_4532);
xor U6353 (N_6353,N_4859,N_3230);
xnor U6354 (N_6354,N_5556,N_4599);
nor U6355 (N_6355,N_5016,N_5259);
xnor U6356 (N_6356,N_3377,N_5382);
xor U6357 (N_6357,N_4621,N_3446);
nor U6358 (N_6358,N_5061,N_4833);
and U6359 (N_6359,N_3139,N_3143);
and U6360 (N_6360,N_4879,N_4315);
nand U6361 (N_6361,N_5169,N_5779);
or U6362 (N_6362,N_5534,N_4129);
xor U6363 (N_6363,N_3828,N_5130);
and U6364 (N_6364,N_6009,N_5475);
and U6365 (N_6365,N_5039,N_3966);
and U6366 (N_6366,N_5510,N_5807);
and U6367 (N_6367,N_5643,N_6071);
nand U6368 (N_6368,N_4084,N_3763);
and U6369 (N_6369,N_4191,N_5210);
or U6370 (N_6370,N_4466,N_3934);
or U6371 (N_6371,N_4571,N_4782);
nand U6372 (N_6372,N_3883,N_3862);
or U6373 (N_6373,N_5172,N_5765);
nor U6374 (N_6374,N_4769,N_5268);
and U6375 (N_6375,N_3528,N_5000);
and U6376 (N_6376,N_6135,N_5439);
and U6377 (N_6377,N_4301,N_5763);
nor U6378 (N_6378,N_3444,N_5205);
xor U6379 (N_6379,N_5491,N_5860);
xnor U6380 (N_6380,N_4417,N_5518);
nand U6381 (N_6381,N_5926,N_4322);
nor U6382 (N_6382,N_4049,N_5963);
nor U6383 (N_6383,N_3661,N_3456);
nor U6384 (N_6384,N_5895,N_5567);
and U6385 (N_6385,N_3559,N_5201);
and U6386 (N_6386,N_3908,N_3880);
nand U6387 (N_6387,N_3692,N_4689);
xor U6388 (N_6388,N_4924,N_5806);
and U6389 (N_6389,N_5403,N_5134);
nand U6390 (N_6390,N_4421,N_3971);
or U6391 (N_6391,N_3921,N_5628);
nand U6392 (N_6392,N_3307,N_4019);
and U6393 (N_6393,N_4671,N_3886);
nor U6394 (N_6394,N_5898,N_4410);
or U6395 (N_6395,N_3327,N_4402);
nor U6396 (N_6396,N_3443,N_5065);
xor U6397 (N_6397,N_4040,N_4717);
nor U6398 (N_6398,N_5012,N_3940);
nor U6399 (N_6399,N_4369,N_4307);
or U6400 (N_6400,N_5427,N_6102);
nand U6401 (N_6401,N_5840,N_4561);
or U6402 (N_6402,N_5237,N_3529);
nand U6403 (N_6403,N_3626,N_5559);
and U6404 (N_6404,N_4528,N_3600);
or U6405 (N_6405,N_3939,N_3974);
nand U6406 (N_6406,N_5253,N_3884);
xor U6407 (N_6407,N_4986,N_3374);
or U6408 (N_6408,N_4989,N_3636);
or U6409 (N_6409,N_5528,N_6243);
and U6410 (N_6410,N_5479,N_5198);
or U6411 (N_6411,N_4266,N_4027);
nor U6412 (N_6412,N_3453,N_4498);
nor U6413 (N_6413,N_4666,N_3249);
and U6414 (N_6414,N_3863,N_6060);
nor U6415 (N_6415,N_3495,N_6212);
xnor U6416 (N_6416,N_5620,N_5300);
or U6417 (N_6417,N_6231,N_3543);
and U6418 (N_6418,N_3978,N_3891);
and U6419 (N_6419,N_3843,N_3930);
and U6420 (N_6420,N_4274,N_4101);
nor U6421 (N_6421,N_4535,N_5305);
nand U6422 (N_6422,N_4503,N_4463);
and U6423 (N_6423,N_3609,N_5948);
nand U6424 (N_6424,N_3813,N_3824);
or U6425 (N_6425,N_6142,N_3743);
and U6426 (N_6426,N_3440,N_5836);
xnor U6427 (N_6427,N_5679,N_4642);
nand U6428 (N_6428,N_5599,N_3232);
or U6429 (N_6429,N_4423,N_5233);
and U6430 (N_6430,N_5805,N_4234);
and U6431 (N_6431,N_3565,N_4874);
and U6432 (N_6432,N_5452,N_3194);
and U6433 (N_6433,N_5287,N_4891);
and U6434 (N_6434,N_5293,N_6104);
nor U6435 (N_6435,N_4756,N_3496);
and U6436 (N_6436,N_3989,N_4857);
xor U6437 (N_6437,N_5047,N_5958);
xnor U6438 (N_6438,N_5404,N_4665);
xor U6439 (N_6439,N_5332,N_5207);
xnor U6440 (N_6440,N_3521,N_4267);
and U6441 (N_6441,N_5451,N_5068);
or U6442 (N_6442,N_4930,N_4167);
and U6443 (N_6443,N_3149,N_3318);
and U6444 (N_6444,N_3788,N_5232);
or U6445 (N_6445,N_5928,N_3730);
xnor U6446 (N_6446,N_5630,N_4697);
xor U6447 (N_6447,N_4805,N_4898);
nand U6448 (N_6448,N_4091,N_5992);
or U6449 (N_6449,N_4964,N_4164);
nand U6450 (N_6450,N_3926,N_3791);
xnor U6451 (N_6451,N_4415,N_3397);
and U6452 (N_6452,N_3129,N_5829);
nor U6453 (N_6453,N_4312,N_6066);
nor U6454 (N_6454,N_4127,N_6214);
nor U6455 (N_6455,N_4940,N_4058);
and U6456 (N_6456,N_5498,N_4124);
nand U6457 (N_6457,N_4038,N_3986);
nor U6458 (N_6458,N_5457,N_4126);
nor U6459 (N_6459,N_5973,N_4031);
or U6460 (N_6460,N_3724,N_5480);
nor U6461 (N_6461,N_4462,N_5733);
and U6462 (N_6462,N_3447,N_4194);
xor U6463 (N_6463,N_4636,N_4723);
nor U6464 (N_6464,N_4497,N_4743);
or U6465 (N_6465,N_5318,N_4468);
xnor U6466 (N_6466,N_4587,N_4386);
or U6467 (N_6467,N_4192,N_5896);
xor U6468 (N_6468,N_5657,N_3202);
nand U6469 (N_6469,N_4975,N_4652);
nand U6470 (N_6470,N_5764,N_5554);
or U6471 (N_6471,N_5037,N_4783);
xnor U6472 (N_6472,N_5003,N_5429);
nor U6473 (N_6473,N_3478,N_4631);
nand U6474 (N_6474,N_4712,N_3160);
xnor U6475 (N_6475,N_4479,N_4646);
nand U6476 (N_6476,N_4458,N_5606);
or U6477 (N_6477,N_5351,N_4355);
nand U6478 (N_6478,N_3535,N_4418);
or U6479 (N_6479,N_3281,N_4039);
xnor U6480 (N_6480,N_3710,N_3270);
nor U6481 (N_6481,N_6028,N_4525);
nand U6482 (N_6482,N_6046,N_5927);
xor U6483 (N_6483,N_4226,N_4353);
and U6484 (N_6484,N_5951,N_5124);
xor U6485 (N_6485,N_5661,N_3268);
nor U6486 (N_6486,N_6196,N_3303);
or U6487 (N_6487,N_3211,N_5241);
and U6488 (N_6488,N_6183,N_4155);
nand U6489 (N_6489,N_4762,N_5041);
nand U6490 (N_6490,N_6179,N_5437);
nor U6491 (N_6491,N_3797,N_3342);
and U6492 (N_6492,N_3326,N_4095);
nand U6493 (N_6493,N_4638,N_3635);
or U6494 (N_6494,N_4097,N_4131);
or U6495 (N_6495,N_4845,N_6217);
xor U6496 (N_6496,N_5833,N_4028);
xor U6497 (N_6497,N_3866,N_4046);
and U6498 (N_6498,N_4557,N_6087);
xor U6499 (N_6499,N_5922,N_3375);
and U6500 (N_6500,N_3563,N_3819);
nor U6501 (N_6501,N_5127,N_4885);
xnor U6502 (N_6502,N_3859,N_4291);
nand U6503 (N_6503,N_3553,N_4431);
and U6504 (N_6504,N_6097,N_3618);
or U6505 (N_6505,N_4921,N_3678);
and U6506 (N_6506,N_3295,N_5731);
nor U6507 (N_6507,N_4054,N_4311);
or U6508 (N_6508,N_5162,N_3670);
and U6509 (N_6509,N_4635,N_3718);
nand U6510 (N_6510,N_3686,N_4972);
and U6511 (N_6511,N_4796,N_5118);
nor U6512 (N_6512,N_5604,N_4905);
nand U6513 (N_6513,N_5692,N_5637);
nand U6514 (N_6514,N_4559,N_5804);
xnor U6515 (N_6515,N_3821,N_5174);
nand U6516 (N_6516,N_5209,N_3871);
and U6517 (N_6517,N_6072,N_5838);
xor U6518 (N_6518,N_6129,N_6110);
and U6519 (N_6519,N_4118,N_4009);
xnor U6520 (N_6520,N_4651,N_4718);
or U6521 (N_6521,N_4527,N_4235);
and U6522 (N_6522,N_4611,N_5740);
and U6523 (N_6523,N_5191,N_4087);
nor U6524 (N_6524,N_4572,N_4427);
and U6525 (N_6525,N_5060,N_5917);
nand U6526 (N_6526,N_5593,N_4128);
nor U6527 (N_6527,N_3448,N_3159);
xnor U6528 (N_6528,N_5976,N_3879);
xor U6529 (N_6529,N_4005,N_5255);
nand U6530 (N_6530,N_3737,N_5705);
nand U6531 (N_6531,N_4560,N_3515);
nor U6532 (N_6532,N_5281,N_5527);
xor U6533 (N_6533,N_4688,N_4145);
or U6534 (N_6534,N_4563,N_5348);
and U6535 (N_6535,N_3765,N_4659);
xor U6536 (N_6536,N_5777,N_5781);
nand U6537 (N_6537,N_3186,N_4531);
nand U6538 (N_6538,N_5677,N_5858);
or U6539 (N_6539,N_4345,N_3641);
xor U6540 (N_6540,N_5030,N_4304);
or U6541 (N_6541,N_4915,N_4802);
nand U6542 (N_6542,N_4872,N_4052);
or U6543 (N_6543,N_4440,N_4048);
xor U6544 (N_6544,N_5048,N_3851);
xor U6545 (N_6545,N_5844,N_5385);
or U6546 (N_6546,N_3755,N_3167);
xor U6547 (N_6547,N_5871,N_5193);
and U6548 (N_6548,N_3392,N_5508);
or U6549 (N_6549,N_3373,N_4606);
and U6550 (N_6550,N_4250,N_5234);
or U6551 (N_6551,N_4663,N_3704);
nor U6552 (N_6552,N_3338,N_4061);
and U6553 (N_6553,N_5734,N_4770);
and U6554 (N_6554,N_5246,N_5675);
nor U6555 (N_6555,N_5655,N_3679);
or U6556 (N_6556,N_4008,N_5962);
xor U6557 (N_6557,N_3191,N_4910);
and U6558 (N_6558,N_5141,N_4324);
nand U6559 (N_6559,N_3504,N_6248);
nand U6560 (N_6560,N_4758,N_4021);
and U6561 (N_6561,N_5980,N_5854);
and U6562 (N_6562,N_5035,N_3996);
and U6563 (N_6563,N_5949,N_5827);
nand U6564 (N_6564,N_5126,N_6098);
or U6565 (N_6565,N_3205,N_3227);
nor U6566 (N_6566,N_3296,N_4137);
xor U6567 (N_6567,N_5329,N_3463);
nor U6568 (N_6568,N_4995,N_3881);
xnor U6569 (N_6569,N_5585,N_3950);
nor U6570 (N_6570,N_4412,N_5652);
nand U6571 (N_6571,N_4255,N_5603);
and U6572 (N_6572,N_3457,N_5330);
nand U6573 (N_6573,N_4071,N_4271);
and U6574 (N_6574,N_5098,N_4690);
nand U6575 (N_6575,N_5227,N_3352);
xnor U6576 (N_6576,N_4216,N_4552);
nor U6577 (N_6577,N_4618,N_3182);
or U6578 (N_6578,N_5155,N_3534);
xor U6579 (N_6579,N_3252,N_3490);
xnor U6580 (N_6580,N_3823,N_5482);
and U6581 (N_6581,N_6024,N_4657);
xnor U6582 (N_6582,N_5634,N_5851);
xnor U6583 (N_6583,N_5054,N_5537);
nor U6584 (N_6584,N_4554,N_3217);
or U6585 (N_6585,N_5421,N_4515);
and U6586 (N_6586,N_4407,N_5629);
nand U6587 (N_6587,N_4203,N_5678);
nand U6588 (N_6588,N_3822,N_4007);
and U6589 (N_6589,N_4523,N_3816);
xnor U6590 (N_6590,N_6045,N_5624);
nor U6591 (N_6591,N_4063,N_3222);
nand U6592 (N_6592,N_3519,N_3261);
or U6593 (N_6593,N_4826,N_5424);
nor U6594 (N_6594,N_5290,N_3394);
xor U6595 (N_6595,N_5495,N_3507);
nor U6596 (N_6596,N_3719,N_4493);
nor U6597 (N_6597,N_5633,N_4681);
nand U6598 (N_6598,N_4067,N_5813);
and U6599 (N_6599,N_4214,N_3216);
nand U6600 (N_6600,N_4329,N_6075);
or U6601 (N_6601,N_3968,N_4086);
and U6602 (N_6602,N_5682,N_5073);
xor U6603 (N_6603,N_3805,N_5815);
xor U6604 (N_6604,N_4753,N_4974);
nand U6605 (N_6605,N_4729,N_3691);
and U6606 (N_6606,N_3287,N_3850);
nor U6607 (N_6607,N_3497,N_5817);
nand U6608 (N_6608,N_3740,N_4456);
xor U6609 (N_6609,N_4825,N_4812);
or U6610 (N_6610,N_4676,N_5934);
nor U6611 (N_6611,N_3840,N_4481);
and U6612 (N_6612,N_3613,N_3723);
nand U6613 (N_6613,N_4724,N_3573);
or U6614 (N_6614,N_5430,N_5409);
nor U6615 (N_6615,N_4607,N_4383);
xor U6616 (N_6616,N_4763,N_6229);
nor U6617 (N_6617,N_4558,N_4740);
nor U6618 (N_6618,N_4895,N_3757);
nand U6619 (N_6619,N_6062,N_3633);
xnor U6620 (N_6620,N_3315,N_5058);
xnor U6621 (N_6621,N_3505,N_5114);
nor U6622 (N_6622,N_3162,N_5203);
and U6623 (N_6623,N_4373,N_5235);
and U6624 (N_6624,N_3694,N_6078);
xnor U6625 (N_6625,N_4516,N_3402);
or U6626 (N_6626,N_3128,N_4927);
or U6627 (N_6627,N_5213,N_4169);
nor U6628 (N_6628,N_4254,N_3698);
nand U6629 (N_6629,N_5143,N_3961);
xnor U6630 (N_6630,N_5333,N_5251);
or U6631 (N_6631,N_4438,N_5472);
nor U6632 (N_6632,N_3774,N_5596);
or U6633 (N_6633,N_3432,N_5449);
or U6634 (N_6634,N_4798,N_3283);
nand U6635 (N_6635,N_3907,N_5204);
xnor U6636 (N_6636,N_6089,N_5078);
nand U6637 (N_6637,N_4959,N_4566);
xor U6638 (N_6638,N_3174,N_3471);
nor U6639 (N_6639,N_5031,N_4994);
nand U6640 (N_6640,N_4776,N_5803);
nand U6641 (N_6641,N_4174,N_4694);
nor U6642 (N_6642,N_3229,N_3712);
xor U6643 (N_6643,N_5214,N_4201);
nor U6644 (N_6644,N_4630,N_4212);
and U6645 (N_6645,N_5615,N_3937);
nand U6646 (N_6646,N_3984,N_4728);
nor U6647 (N_6647,N_6068,N_5089);
nand U6648 (N_6648,N_6122,N_3759);
or U6649 (N_6649,N_5323,N_6127);
nor U6650 (N_6650,N_3672,N_5243);
nand U6651 (N_6651,N_5525,N_3736);
and U6652 (N_6652,N_3451,N_5668);
nor U6653 (N_6653,N_5131,N_4397);
and U6654 (N_6654,N_4434,N_5891);
nor U6655 (N_6655,N_4894,N_5343);
nor U6656 (N_6656,N_5959,N_5257);
nor U6657 (N_6657,N_4744,N_6033);
xor U6658 (N_6658,N_6157,N_4828);
and U6659 (N_6659,N_4483,N_4245);
or U6660 (N_6660,N_5056,N_6011);
nor U6661 (N_6661,N_3731,N_5889);
or U6662 (N_6662,N_5878,N_3860);
nand U6663 (N_6663,N_5342,N_3333);
xor U6664 (N_6664,N_3892,N_3153);
xnor U6665 (N_6665,N_5171,N_3218);
nor U6666 (N_6666,N_5288,N_4188);
nor U6667 (N_6667,N_4496,N_3265);
nand U6668 (N_6668,N_3356,N_3664);
or U6669 (N_6669,N_5185,N_3876);
or U6670 (N_6670,N_3399,N_4911);
nor U6671 (N_6671,N_3301,N_3258);
xor U6672 (N_6672,N_5656,N_4877);
xor U6673 (N_6673,N_4268,N_3951);
or U6674 (N_6674,N_4938,N_3508);
or U6675 (N_6675,N_4284,N_4435);
nand U6676 (N_6676,N_3225,N_4928);
xnor U6677 (N_6677,N_6223,N_3629);
nor U6678 (N_6678,N_3417,N_3437);
nand U6679 (N_6679,N_6180,N_6165);
nand U6680 (N_6680,N_6070,N_5790);
xnor U6681 (N_6681,N_5866,N_4449);
nor U6682 (N_6682,N_3165,N_5536);
and U6683 (N_6683,N_4912,N_5286);
and U6684 (N_6684,N_5483,N_6092);
xor U6685 (N_6685,N_3711,N_5184);
nor U6686 (N_6686,N_3137,N_4977);
xnor U6687 (N_6687,N_4870,N_4734);
nand U6688 (N_6688,N_3419,N_3952);
and U6689 (N_6689,N_4069,N_5576);
or U6690 (N_6690,N_5419,N_6084);
xnor U6691 (N_6691,N_4965,N_3349);
and U6692 (N_6692,N_3674,N_5759);
or U6693 (N_6693,N_6003,N_3304);
or U6694 (N_6694,N_6086,N_4453);
and U6695 (N_6695,N_5654,N_4070);
nand U6696 (N_6696,N_4840,N_4173);
or U6697 (N_6697,N_3802,N_4967);
or U6698 (N_6698,N_3663,N_4036);
or U6699 (N_6699,N_3709,N_4372);
nand U6700 (N_6700,N_4597,N_3720);
xor U6701 (N_6701,N_4025,N_3236);
or U6702 (N_6702,N_5816,N_3854);
xnor U6703 (N_6703,N_5762,N_4550);
xnor U6704 (N_6704,N_5021,N_4820);
nand U6705 (N_6705,N_3127,N_4178);
nand U6706 (N_6706,N_3485,N_4248);
and U6707 (N_6707,N_5441,N_4116);
or U6708 (N_6708,N_3993,N_5886);
nor U6709 (N_6709,N_5880,N_4096);
nand U6710 (N_6710,N_4180,N_3815);
nor U6711 (N_6711,N_5316,N_3834);
xor U6712 (N_6712,N_5943,N_5571);
nor U6713 (N_6713,N_4448,N_3282);
xnor U6714 (N_6714,N_5163,N_4018);
nand U6715 (N_6715,N_3796,N_5448);
or U6716 (N_6716,N_5704,N_4055);
or U6717 (N_6717,N_4752,N_6147);
and U6718 (N_6718,N_4494,N_5256);
nor U6719 (N_6719,N_3297,N_4939);
or U6720 (N_6720,N_5888,N_4342);
nand U6721 (N_6721,N_4391,N_3339);
xnor U6722 (N_6722,N_5244,N_6111);
nand U6723 (N_6723,N_4968,N_5746);
and U6724 (N_6724,N_6168,N_5828);
nand U6725 (N_6725,N_5837,N_3347);
nand U6726 (N_6726,N_4923,N_5747);
nor U6727 (N_6727,N_3389,N_3739);
nand U6728 (N_6728,N_4401,N_6094);
nor U6729 (N_6729,N_3412,N_3538);
and U6730 (N_6730,N_5123,N_4029);
nor U6731 (N_6731,N_4962,N_3381);
nor U6732 (N_6732,N_4991,N_3969);
and U6733 (N_6733,N_5524,N_4822);
nand U6734 (N_6734,N_3762,N_3790);
or U6735 (N_6735,N_3605,N_5489);
nor U6736 (N_6736,N_5726,N_3914);
or U6737 (N_6737,N_5090,N_5195);
or U6738 (N_6738,N_5460,N_3684);
nor U6739 (N_6739,N_4733,N_5453);
xnor U6740 (N_6740,N_5664,N_3346);
and U6741 (N_6741,N_3179,N_5181);
or U6742 (N_6742,N_5520,N_4976);
nand U6743 (N_6743,N_6041,N_4034);
nand U6744 (N_6744,N_5432,N_6224);
nor U6745 (N_6745,N_3826,N_5360);
and U6746 (N_6746,N_3491,N_4658);
or U6747 (N_6747,N_5771,N_5551);
xor U6748 (N_6748,N_6056,N_5622);
nand U6749 (N_6749,N_4231,N_3360);
or U6750 (N_6750,N_5824,N_5050);
nor U6751 (N_6751,N_3290,N_5487);
and U6752 (N_6752,N_5902,N_5674);
and U6753 (N_6753,N_5294,N_3271);
xor U6754 (N_6754,N_3324,N_3248);
or U6755 (N_6755,N_4500,N_4112);
nand U6756 (N_6756,N_3537,N_4211);
nor U6757 (N_6757,N_5435,N_4290);
xor U6758 (N_6758,N_3806,N_5349);
and U6759 (N_6759,N_5770,N_5942);
nand U6760 (N_6760,N_5685,N_5605);
and U6761 (N_6761,N_5321,N_4799);
or U6762 (N_6762,N_3903,N_4661);
nand U6763 (N_6763,N_4220,N_5947);
or U6764 (N_6764,N_3820,N_4882);
nand U6765 (N_6765,N_4141,N_3973);
xnor U6766 (N_6766,N_5159,N_3606);
or U6767 (N_6767,N_5987,N_6238);
nor U6768 (N_6768,N_3354,N_4371);
nand U6769 (N_6769,N_4142,N_4970);
or U6770 (N_6770,N_4474,N_4205);
or U6771 (N_6771,N_3187,N_4590);
or U6772 (N_6772,N_5069,N_5775);
and U6773 (N_6773,N_6225,N_3503);
or U6774 (N_6774,N_5669,N_6178);
or U6775 (N_6775,N_5049,N_5901);
xnor U6776 (N_6776,N_5340,N_4202);
or U6777 (N_6777,N_5364,N_5977);
and U6778 (N_6778,N_5749,N_3200);
and U6779 (N_6779,N_5530,N_3846);
nor U6780 (N_6780,N_3308,N_5855);
or U6781 (N_6781,N_6043,N_4470);
nor U6782 (N_6782,N_5784,N_4251);
or U6783 (N_6783,N_3598,N_4992);
xnor U6784 (N_6784,N_3450,N_5904);
or U6785 (N_6785,N_4296,N_3423);
nand U6786 (N_6786,N_4906,N_4513);
nor U6787 (N_6787,N_3501,N_4595);
nand U6788 (N_6788,N_3243,N_5548);
or U6789 (N_6789,N_5104,N_5391);
and U6790 (N_6790,N_3658,N_3226);
or U6791 (N_6791,N_3900,N_4596);
nor U6792 (N_6792,N_5786,N_3329);
and U6793 (N_6793,N_4012,N_3941);
xnor U6794 (N_6794,N_5346,N_3735);
and U6795 (N_6795,N_5707,N_3277);
or U6796 (N_6796,N_5296,N_6064);
nor U6797 (N_6797,N_3317,N_5706);
and U6798 (N_6798,N_4351,N_3627);
xor U6799 (N_6799,N_4090,N_4719);
nor U6800 (N_6800,N_5932,N_3192);
nand U6801 (N_6801,N_4319,N_5553);
nand U6802 (N_6802,N_5312,N_3569);
xor U6803 (N_6803,N_5295,N_6205);
and U6804 (N_6804,N_3982,N_5418);
xnor U6805 (N_6805,N_3751,N_3716);
xor U6806 (N_6806,N_3979,N_5226);
nand U6807 (N_6807,N_3588,N_4679);
xor U6808 (N_6808,N_4754,N_3809);
and U6809 (N_6809,N_5149,N_3906);
nand U6810 (N_6810,N_4949,N_4576);
and U6811 (N_6811,N_3204,N_3722);
nor U6812 (N_6812,N_3555,N_3152);
nand U6813 (N_6813,N_5107,N_4476);
nand U6814 (N_6814,N_3785,N_3807);
xnor U6815 (N_6815,N_5857,N_6216);
and U6816 (N_6816,N_5334,N_6042);
nor U6817 (N_6817,N_5376,N_4958);
and U6818 (N_6818,N_4836,N_5179);
and U6819 (N_6819,N_4287,N_5507);
xnor U6820 (N_6820,N_5575,N_4265);
nand U6821 (N_6821,N_4261,N_6010);
nand U6822 (N_6822,N_5954,N_5988);
nor U6823 (N_6823,N_3337,N_3156);
nor U6824 (N_6824,N_4477,N_4806);
and U6825 (N_6825,N_3267,N_3779);
or U6826 (N_6826,N_4888,N_6039);
or U6827 (N_6827,N_5190,N_5477);
nor U6828 (N_6828,N_4305,N_5550);
nor U6829 (N_6829,N_4152,N_4542);
xor U6830 (N_6830,N_6096,N_6126);
nor U6831 (N_6831,N_4567,N_6004);
nor U6832 (N_6832,N_6153,N_5412);
xnor U6833 (N_6833,N_6228,N_3488);
and U6834 (N_6834,N_4858,N_3240);
or U6835 (N_6835,N_4793,N_5470);
xnor U6836 (N_6836,N_5088,N_4253);
nand U6837 (N_6837,N_3781,N_5466);
and U6838 (N_6838,N_3164,N_5910);
nand U6839 (N_6839,N_4416,N_5027);
xnor U6840 (N_6840,N_4760,N_6051);
xnor U6841 (N_6841,N_5681,N_4868);
and U6842 (N_6842,N_3780,N_4721);
xnor U6843 (N_6843,N_4639,N_4687);
or U6844 (N_6844,N_4908,N_5975);
xnor U6845 (N_6845,N_4134,N_5062);
nand U6846 (N_6846,N_4381,N_5223);
xor U6847 (N_6847,N_3279,N_3673);
or U6848 (N_6848,N_6031,N_4884);
xnor U6849 (N_6849,N_3237,N_4843);
and U6850 (N_6850,N_4818,N_4487);
and U6851 (N_6851,N_3517,N_3455);
nor U6852 (N_6852,N_4993,N_5953);
or U6853 (N_6853,N_6175,N_4419);
or U6854 (N_6854,N_4374,N_4699);
nor U6855 (N_6855,N_4680,N_5138);
nand U6856 (N_6856,N_5588,N_4002);
xnor U6857 (N_6857,N_5355,N_3172);
nand U6858 (N_6858,N_3278,N_5454);
xnor U6859 (N_6859,N_3577,N_4551);
or U6860 (N_6860,N_3390,N_6121);
and U6861 (N_6861,N_4832,N_4577);
nand U6862 (N_6862,N_4983,N_4589);
nor U6863 (N_6863,N_4239,N_3213);
nand U6864 (N_6864,N_5578,N_3938);
nand U6865 (N_6865,N_4282,N_4368);
nand U6866 (N_6866,N_4869,N_5903);
xor U6867 (N_6867,N_6226,N_4749);
and U6868 (N_6868,N_4672,N_4568);
xor U6869 (N_6869,N_4102,N_6242);
xnor U6870 (N_6870,N_3865,N_4546);
nand U6871 (N_6871,N_4283,N_5405);
nor U6872 (N_6872,N_3408,N_3255);
or U6873 (N_6873,N_6063,N_6209);
or U6874 (N_6874,N_6176,N_5568);
or U6875 (N_6875,N_4306,N_4960);
and U6876 (N_6876,N_3888,N_3430);
and U6877 (N_6877,N_4321,N_4179);
nand U6878 (N_6878,N_5011,N_3299);
and U6879 (N_6879,N_5228,N_4308);
nand U6880 (N_6880,N_3147,N_4800);
and U6881 (N_6881,N_4713,N_4429);
nor U6882 (N_6882,N_5401,N_5499);
or U6883 (N_6883,N_5462,N_5595);
nand U6884 (N_6884,N_4083,N_3895);
nor U6885 (N_6885,N_5046,N_5598);
and U6886 (N_6886,N_3753,N_3449);
xor U6887 (N_6887,N_6067,N_4883);
nand U6888 (N_6888,N_4339,N_4098);
nand U6889 (N_6889,N_4010,N_5727);
nand U6890 (N_6890,N_4409,N_3524);
or U6891 (N_6891,N_4706,N_5133);
or U6892 (N_6892,N_5320,N_4451);
xnor U6893 (N_6893,N_3818,N_4472);
xor U6894 (N_6894,N_3944,N_4162);
xor U6895 (N_6895,N_3379,N_4147);
nand U6896 (N_6896,N_3725,N_3835);
nor U6897 (N_6897,N_3936,N_5465);
or U6898 (N_6898,N_6186,N_5280);
nor U6899 (N_6899,N_3610,N_3445);
nand U6900 (N_6900,N_4032,N_4787);
nor U6901 (N_6901,N_3983,N_4582);
xnor U6902 (N_6902,N_3395,N_4925);
xor U6903 (N_6903,N_6053,N_4075);
xnor U6904 (N_6904,N_3335,N_4814);
xnor U6905 (N_6905,N_4725,N_6233);
xor U6906 (N_6906,N_3144,N_3942);
xnor U6907 (N_6907,N_4450,N_5438);
or U6908 (N_6908,N_5885,N_5408);
or U6909 (N_6909,N_3212,N_3949);
nand U6910 (N_6910,N_3438,N_5319);
and U6911 (N_6911,N_3987,N_4317);
and U6912 (N_6912,N_3312,N_5208);
xor U6913 (N_6913,N_4570,N_3371);
nor U6914 (N_6914,N_3472,N_5982);
nand U6915 (N_6915,N_3889,N_4241);
nor U6916 (N_6916,N_4043,N_4064);
nor U6917 (N_6917,N_4115,N_4648);
or U6918 (N_6918,N_4653,N_5032);
nand U6919 (N_6919,N_4598,N_3911);
xnor U6920 (N_6920,N_5730,N_5506);
xor U6921 (N_6921,N_4863,N_4157);
nor U6922 (N_6922,N_5969,N_6220);
nand U6923 (N_6923,N_4540,N_4236);
nor U6924 (N_6924,N_4185,N_5995);
and U6925 (N_6925,N_5215,N_3428);
or U6926 (N_6926,N_3284,N_4821);
or U6927 (N_6927,N_5874,N_4459);
nand U6928 (N_6928,N_6174,N_5712);
or U6929 (N_6929,N_4580,N_5381);
nand U6930 (N_6930,N_3208,N_5292);
or U6931 (N_6931,N_4981,N_4333);
nor U6932 (N_6932,N_6093,N_3799);
or U6933 (N_6933,N_4328,N_5612);
nor U6934 (N_6934,N_3829,N_3310);
or U6935 (N_6935,N_6246,N_6140);
and U6936 (N_6936,N_3131,N_4445);
nor U6937 (N_6937,N_4955,N_4637);
xor U6938 (N_6938,N_4813,N_5684);
nor U6939 (N_6939,N_3706,N_4015);
nor U6940 (N_6940,N_5879,N_4755);
nand U6941 (N_6941,N_3474,N_6138);
nor U6942 (N_6942,N_4139,N_5239);
and U6943 (N_6943,N_3150,N_3420);
xnor U6944 (N_6944,N_4750,N_3873);
xnor U6945 (N_6945,N_4517,N_3557);
xnor U6946 (N_6946,N_4781,N_3833);
and U6947 (N_6947,N_4602,N_3651);
nand U6948 (N_6948,N_6037,N_3264);
nand U6949 (N_6949,N_4318,N_6236);
and U6950 (N_6950,N_5378,N_3749);
and U6951 (N_6951,N_3772,N_5103);
and U6952 (N_6952,N_4693,N_5663);
and U6953 (N_6953,N_4172,N_3808);
xor U6954 (N_6954,N_5220,N_5070);
nor U6955 (N_6955,N_3468,N_5269);
and U6956 (N_6956,N_4259,N_4708);
or U6957 (N_6957,N_4746,N_5384);
and U6958 (N_6958,N_4217,N_4228);
xor U6959 (N_6959,N_4299,N_6059);
xor U6960 (N_6960,N_3562,N_4641);
and U6961 (N_6961,N_3933,N_3680);
nor U6962 (N_6962,N_4171,N_5277);
nor U6963 (N_6963,N_3203,N_5887);
xnor U6964 (N_6964,N_6077,N_5564);
xnor U6965 (N_6965,N_3166,N_5345);
nor U6966 (N_6966,N_6150,N_5137);
or U6967 (N_6967,N_4951,N_4624);
xor U6968 (N_6968,N_5117,N_4616);
or U6969 (N_6969,N_4024,N_3407);
or U6970 (N_6970,N_5249,N_5868);
xnor U6971 (N_6971,N_3502,N_5356);
and U6972 (N_6972,N_4668,N_4791);
and U6973 (N_6973,N_5597,N_4136);
nor U6974 (N_6974,N_4303,N_4850);
xnor U6975 (N_6975,N_3434,N_4819);
xor U6976 (N_6976,N_3498,N_5414);
or U6977 (N_6977,N_5076,N_3396);
xnor U6978 (N_6978,N_4873,N_4944);
xor U6979 (N_6979,N_4471,N_3990);
nor U6980 (N_6980,N_3632,N_5830);
and U6981 (N_6981,N_6082,N_4200);
and U6982 (N_6982,N_4062,N_4683);
xor U6983 (N_6983,N_5513,N_3738);
nor U6984 (N_6984,N_4144,N_3976);
nor U6985 (N_6985,N_4685,N_5410);
xor U6986 (N_6986,N_6163,N_3322);
and U6987 (N_6987,N_5486,N_6112);
xnor U6988 (N_6988,N_5847,N_4380);
or U6989 (N_6989,N_5423,N_5756);
nand U6990 (N_6990,N_4736,N_6188);
or U6991 (N_6991,N_5467,N_4614);
and U6992 (N_6992,N_4889,N_4610);
xor U6993 (N_6993,N_3477,N_4547);
or U6994 (N_6994,N_5785,N_5067);
xnor U6995 (N_6995,N_4436,N_4533);
nor U6996 (N_6996,N_5484,N_3624);
and U6997 (N_6997,N_4654,N_5583);
or U6998 (N_6998,N_4957,N_3611);
nand U6999 (N_6999,N_3804,N_4001);
or U7000 (N_7000,N_4094,N_5042);
or U7001 (N_7001,N_5822,N_5129);
xor U7002 (N_7002,N_4196,N_4336);
or U7003 (N_7003,N_4044,N_4817);
nor U7004 (N_7004,N_4601,N_5150);
or U7005 (N_7005,N_3916,N_4555);
and U7006 (N_7006,N_3168,N_5387);
xor U7007 (N_7007,N_4093,N_4378);
and U7008 (N_7008,N_5002,N_3241);
and U7009 (N_7009,N_5956,N_4076);
nor U7010 (N_7010,N_4778,N_5013);
or U7011 (N_7011,N_3677,N_5059);
xnor U7012 (N_7012,N_4110,N_4346);
nor U7013 (N_7013,N_5170,N_3533);
nand U7014 (N_7014,N_4461,N_4709);
and U7015 (N_7015,N_4229,N_3958);
nand U7016 (N_7016,N_3803,N_3904);
nor U7017 (N_7017,N_3233,N_6065);
nand U7018 (N_7018,N_5864,N_5379);
nand U7019 (N_7019,N_4792,N_4979);
xnor U7020 (N_7020,N_6021,N_6149);
nand U7021 (N_7021,N_4332,N_5468);
nand U7022 (N_7022,N_3848,N_3954);
and U7023 (N_7023,N_4715,N_3578);
nand U7024 (N_7024,N_3292,N_5950);
nand U7025 (N_7025,N_4140,N_3697);
xnor U7026 (N_7026,N_4156,N_5711);
xor U7027 (N_7027,N_3587,N_5610);
nand U7028 (N_7028,N_4289,N_3959);
nor U7029 (N_7029,N_3741,N_4506);
and U7030 (N_7030,N_5591,N_5736);
nor U7031 (N_7031,N_4135,N_4952);
xor U7032 (N_7032,N_5640,N_3378);
or U7033 (N_7033,N_4620,N_6113);
and U7034 (N_7034,N_5761,N_6105);
or U7035 (N_7035,N_5231,N_5665);
or U7036 (N_7036,N_5336,N_6085);
and U7037 (N_7037,N_3414,N_3701);
nor U7038 (N_7038,N_5289,N_4082);
or U7039 (N_7039,N_3416,N_5225);
xnor U7040 (N_7040,N_6076,N_4565);
nor U7041 (N_7041,N_5307,N_6000);
xor U7042 (N_7042,N_5426,N_4475);
nand U7043 (N_7043,N_6044,N_4232);
or U7044 (N_7044,N_3387,N_4504);
or U7045 (N_7045,N_4748,N_5094);
nand U7046 (N_7046,N_5347,N_3403);
and U7047 (N_7047,N_3800,N_4838);
or U7048 (N_7048,N_6134,N_5646);
or U7049 (N_7049,N_4151,N_4727);
nor U7050 (N_7050,N_5315,N_5112);
or U7051 (N_7051,N_4835,N_4574);
and U7052 (N_7052,N_5377,N_5946);
nor U7053 (N_7053,N_5282,N_4060);
or U7054 (N_7054,N_4741,N_3516);
nor U7055 (N_7055,N_5850,N_5407);
or U7056 (N_7056,N_4811,N_4388);
or U7057 (N_7057,N_3582,N_4065);
and U7058 (N_7058,N_3699,N_3832);
and U7059 (N_7059,N_5997,N_4447);
nand U7060 (N_7060,N_5254,N_3897);
or U7061 (N_7061,N_5580,N_4081);
or U7062 (N_7062,N_4186,N_4913);
nand U7063 (N_7063,N_3845,N_5635);
nor U7064 (N_7064,N_3909,N_5916);
xor U7065 (N_7065,N_5218,N_4737);
and U7066 (N_7066,N_3583,N_5648);
and U7067 (N_7067,N_3839,N_3196);
nand U7068 (N_7068,N_5972,N_5463);
and U7069 (N_7069,N_3874,N_4330);
nand U7070 (N_7070,N_5728,N_3707);
and U7071 (N_7071,N_3180,N_6109);
xor U7072 (N_7072,N_4732,N_5252);
and U7073 (N_7073,N_5128,N_3348);
xnor U7074 (N_7074,N_3693,N_3593);
xor U7075 (N_7075,N_5546,N_5521);
nor U7076 (N_7076,N_6197,N_3640);
or U7077 (N_7077,N_3817,N_4337);
nor U7078 (N_7078,N_4183,N_4059);
nor U7079 (N_7079,N_5841,N_5001);
nor U7080 (N_7080,N_3340,N_5189);
nor U7081 (N_7081,N_3325,N_4242);
nor U7082 (N_7082,N_6203,N_4340);
nor U7083 (N_7083,N_5930,N_3844);
xor U7084 (N_7084,N_4195,N_5776);
nor U7085 (N_7085,N_5194,N_5832);
nand U7086 (N_7086,N_3721,N_5600);
and U7087 (N_7087,N_3784,N_3235);
nand U7088 (N_7088,N_5029,N_4691);
and U7089 (N_7089,N_5380,N_5780);
nor U7090 (N_7090,N_3619,N_4320);
nand U7091 (N_7091,N_3837,N_5022);
and U7092 (N_7092,N_3219,N_5178);
nand U7093 (N_7093,N_3750,N_4105);
and U7094 (N_7094,N_4892,N_3286);
xor U7095 (N_7095,N_5614,N_5799);
and U7096 (N_7096,N_3135,N_4066);
nand U7097 (N_7097,N_3177,N_6120);
and U7098 (N_7098,N_4243,N_6100);
xnor U7099 (N_7099,N_4022,N_5751);
and U7100 (N_7100,N_4961,N_3475);
nand U7101 (N_7101,N_5846,N_4692);
and U7102 (N_7102,N_5248,N_4221);
nor U7103 (N_7103,N_4455,N_4543);
xor U7104 (N_7104,N_3199,N_3169);
nand U7105 (N_7105,N_4165,N_4808);
or U7106 (N_7106,N_4673,N_4398);
nor U7107 (N_7107,N_3201,N_5339);
nand U7108 (N_7108,N_3141,N_6029);
xnor U7109 (N_7109,N_6020,N_4119);
xnor U7110 (N_7110,N_5897,N_5503);
nor U7111 (N_7111,N_3195,N_5659);
xnor U7112 (N_7112,N_4424,N_3997);
and U7113 (N_7113,N_4640,N_6162);
or U7114 (N_7114,N_4023,N_3247);
xor U7115 (N_7115,N_4696,N_6119);
xnor U7116 (N_7116,N_3171,N_4016);
nor U7117 (N_7117,N_4897,N_5873);
nand U7118 (N_7118,N_5768,N_4644);
nor U7119 (N_7119,N_4534,N_4847);
and U7120 (N_7120,N_5461,N_4591);
nand U7121 (N_7121,N_5373,N_3353);
or U7122 (N_7122,N_5601,N_4933);
xor U7123 (N_7123,N_3476,N_5111);
nand U7124 (N_7124,N_5122,N_5362);
nor U7125 (N_7125,N_4600,N_4252);
nor U7126 (N_7126,N_3946,N_3170);
and U7127 (N_7127,N_5582,N_5045);
or U7128 (N_7128,N_5842,N_6107);
and U7129 (N_7129,N_5722,N_4711);
nor U7130 (N_7130,N_3852,N_4584);
nand U7131 (N_7131,N_5375,N_6032);
or U7132 (N_7132,N_3523,N_4390);
and U7133 (N_7133,N_5558,N_4488);
and U7134 (N_7134,N_3442,N_5641);
xor U7135 (N_7135,N_5788,N_5566);
xnor U7136 (N_7136,N_3789,N_4950);
nor U7137 (N_7137,N_3929,N_5132);
and U7138 (N_7138,N_3305,N_6237);
and U7139 (N_7139,N_6058,N_4918);
or U7140 (N_7140,N_4334,N_3486);
nor U7141 (N_7141,N_3924,N_4206);
xor U7142 (N_7142,N_3594,N_3948);
nor U7143 (N_7143,N_5936,N_5981);
or U7144 (N_7144,N_4478,N_5795);
xor U7145 (N_7145,N_5607,N_5702);
xnor U7146 (N_7146,N_5219,N_4909);
and U7147 (N_7147,N_5714,N_5631);
nor U7148 (N_7148,N_5724,N_5298);
nand U7149 (N_7149,N_3649,N_6169);
and U7150 (N_7150,N_4223,N_5651);
nand U7151 (N_7151,N_3280,N_4745);
nand U7152 (N_7152,N_6115,N_3638);
or U7153 (N_7153,N_5136,N_5676);
nand U7154 (N_7154,N_6116,N_4499);
nor U7155 (N_7155,N_5743,N_4893);
xnor U7156 (N_7156,N_3130,N_4106);
or U7157 (N_7157,N_3998,N_5519);
and U7158 (N_7158,N_3454,N_4771);
nand U7159 (N_7159,N_4399,N_5812);
and U7160 (N_7160,N_3967,N_3263);
nor U7161 (N_7161,N_6202,N_3849);
xnor U7162 (N_7162,N_5589,N_3269);
and U7163 (N_7163,N_6245,N_5872);
nand U7164 (N_7164,N_5778,N_4774);
and U7165 (N_7165,N_5425,N_3580);
or U7166 (N_7166,N_5302,N_5279);
nand U7167 (N_7167,N_3681,N_3890);
nand U7168 (N_7168,N_3370,N_5344);
xor U7169 (N_7169,N_4537,N_5820);
and U7170 (N_7170,N_4275,N_4839);
or U7171 (N_7171,N_3513,N_3919);
and U7172 (N_7172,N_5034,N_4247);
and U7173 (N_7173,N_4224,N_5687);
xnor U7174 (N_7174,N_5247,N_3473);
or U7175 (N_7175,N_5271,N_5758);
nor U7176 (N_7176,N_6189,N_3359);
and U7177 (N_7177,N_3905,N_4189);
nand U7178 (N_7178,N_3539,N_3668);
nand U7179 (N_7179,N_5400,N_4604);
nor U7180 (N_7180,N_5180,N_3466);
and U7181 (N_7181,N_5019,N_5542);
nand U7182 (N_7182,N_3793,N_3554);
nor U7183 (N_7183,N_4867,N_4764);
and U7184 (N_7184,N_5142,N_3574);
xnor U7185 (N_7185,N_3511,N_3857);
xnor U7186 (N_7186,N_4218,N_5825);
xor U7187 (N_7187,N_5080,N_5297);
xnor U7188 (N_7188,N_3509,N_3259);
or U7189 (N_7189,N_3136,N_6048);
xor U7190 (N_7190,N_4773,N_4425);
nor U7191 (N_7191,N_3391,N_3867);
and U7192 (N_7192,N_5101,N_4608);
nor U7193 (N_7193,N_5028,N_4457);
or U7194 (N_7194,N_6018,N_5359);
nand U7195 (N_7195,N_5517,N_3603);
or U7196 (N_7196,N_5586,N_5970);
nand U7197 (N_7197,N_5772,N_5121);
nand U7198 (N_7198,N_5192,N_5853);
and U7199 (N_7199,N_5709,N_5892);
nand U7200 (N_7200,N_4660,N_4276);
or U7201 (N_7201,N_5370,N_5055);
nand U7202 (N_7202,N_4170,N_4855);
nand U7203 (N_7203,N_4522,N_4358);
or U7204 (N_7204,N_4208,N_5986);
xnor U7205 (N_7205,N_4354,N_3570);
and U7206 (N_7206,N_3426,N_5945);
xor U7207 (N_7207,N_5691,N_5650);
or U7208 (N_7208,N_3481,N_4104);
or U7209 (N_7209,N_4700,N_5053);
xor U7210 (N_7210,N_4107,N_5238);
and U7211 (N_7211,N_4932,N_4347);
or U7212 (N_7212,N_6139,N_5680);
nor U7213 (N_7213,N_5818,N_3330);
or U7214 (N_7214,N_4460,N_4117);
nand U7215 (N_7215,N_4433,N_3607);
nand U7216 (N_7216,N_4539,N_5275);
xor U7217 (N_7217,N_4085,N_4617);
xnor U7218 (N_7218,N_4103,N_4361);
and U7219 (N_7219,N_5870,N_6081);
or U7220 (N_7220,N_5396,N_3207);
nand U7221 (N_7221,N_3250,N_4230);
and U7222 (N_7222,N_3732,N_5560);
or U7223 (N_7223,N_5485,N_6079);
and U7224 (N_7224,N_5216,N_4603);
or U7225 (N_7225,N_5911,N_5590);
xor U7226 (N_7226,N_4160,N_3920);
and U7227 (N_7227,N_4536,N_5082);
or U7228 (N_7228,N_6117,N_5800);
or U7229 (N_7229,N_4650,N_5636);
nand U7230 (N_7230,N_3760,N_4880);
or U7231 (N_7231,N_6007,N_5971);
nand U7232 (N_7232,N_5869,N_5794);
nand U7233 (N_7233,N_5264,N_5744);
and U7234 (N_7234,N_6143,N_3769);
nand U7235 (N_7235,N_5694,N_4444);
or U7236 (N_7236,N_3616,N_5383);
nand U7237 (N_7237,N_3436,N_4491);
and U7238 (N_7238,N_3133,N_5108);
nor U7239 (N_7239,N_4946,N_4829);
nor U7240 (N_7240,N_3896,N_5789);
or U7241 (N_7241,N_6172,N_3650);
and U7242 (N_7242,N_5957,N_5005);
and U7243 (N_7243,N_3571,N_4074);
nor U7244 (N_7244,N_5721,N_5417);
and U7245 (N_7245,N_6005,N_4899);
nor U7246 (N_7246,N_4518,N_5071);
nor U7247 (N_7247,N_4207,N_4827);
or U7248 (N_7248,N_4887,N_6036);
and U7249 (N_7249,N_5471,N_3189);
nor U7250 (N_7250,N_4966,N_3579);
xnor U7251 (N_7251,N_4313,N_5925);
nand U7252 (N_7252,N_6099,N_4519);
and U7253 (N_7253,N_4045,N_5442);
nor U7254 (N_7254,N_4866,N_5811);
nor U7255 (N_7255,N_3314,N_3689);
or U7256 (N_7256,N_5592,N_4612);
and U7257 (N_7257,N_4878,N_4530);
or U7258 (N_7258,N_4260,N_4865);
and U7259 (N_7259,N_4586,N_4846);
nand U7260 (N_7260,N_3801,N_5436);
xor U7261 (N_7261,N_5274,N_6211);
or U7262 (N_7262,N_5563,N_5814);
or U7263 (N_7263,N_4233,N_4509);
and U7264 (N_7264,N_5523,N_5683);
or U7265 (N_7265,N_5882,N_4256);
xnor U7266 (N_7266,N_5266,N_5328);
or U7267 (N_7267,N_5915,N_6125);
or U7268 (N_7268,N_4816,N_3604);
nand U7269 (N_7269,N_3512,N_5539);
nand U7270 (N_7270,N_4987,N_4187);
and U7271 (N_7271,N_5608,N_3980);
and U7272 (N_7272,N_3275,N_3487);
and U7273 (N_7273,N_3696,N_6155);
xor U7274 (N_7274,N_5540,N_4931);
nor U7275 (N_7275,N_5145,N_5125);
nand U7276 (N_7276,N_6080,N_3198);
nand U7277 (N_7277,N_5086,N_3590);
and U7278 (N_7278,N_4006,N_3546);
nor U7279 (N_7279,N_4400,N_3885);
and U7280 (N_7280,N_5732,N_6232);
and U7281 (N_7281,N_5369,N_6208);
nand U7282 (N_7282,N_4331,N_6069);
and U7283 (N_7283,N_5710,N_5533);
and U7284 (N_7284,N_6001,N_5935);
nand U7285 (N_7285,N_4592,N_4914);
nor U7286 (N_7286,N_3917,N_4943);
xor U7287 (N_7287,N_3999,N_4298);
and U7288 (N_7288,N_6088,N_6013);
or U7289 (N_7289,N_4286,N_4875);
and U7290 (N_7290,N_4649,N_3656);
or U7291 (N_7291,N_3931,N_3733);
nor U7292 (N_7292,N_4406,N_3341);
xor U7293 (N_7293,N_4726,N_3228);
nor U7294 (N_7294,N_5616,N_3810);
or U7295 (N_7295,N_5066,N_6108);
and U7296 (N_7296,N_4548,N_5168);
xnor U7297 (N_7297,N_5993,N_3623);
nand U7298 (N_7298,N_4073,N_5757);
nor U7299 (N_7299,N_4113,N_4485);
or U7300 (N_7300,N_3323,N_5357);
nand U7301 (N_7301,N_5723,N_5964);
nand U7302 (N_7302,N_6015,N_3981);
xor U7303 (N_7303,N_5626,N_6052);
and U7304 (N_7304,N_3742,N_4759);
and U7305 (N_7305,N_3154,N_5202);
or U7306 (N_7306,N_4579,N_5921);
nand U7307 (N_7307,N_5303,N_5481);
nor U7308 (N_7308,N_4615,N_3363);
and U7309 (N_7309,N_5164,N_5562);
and U7310 (N_7310,N_4480,N_3612);
nor U7311 (N_7311,N_3288,N_3794);
xnor U7312 (N_7312,N_5552,N_4633);
and U7313 (N_7313,N_5265,N_5797);
and U7314 (N_7314,N_4645,N_3257);
nor U7315 (N_7315,N_3321,N_3847);
and U7316 (N_7316,N_4520,N_3556);
nor U7317 (N_7317,N_4176,N_4896);
and U7318 (N_7318,N_3467,N_5326);
nor U7319 (N_7319,N_5952,N_5544);
or U7320 (N_7320,N_4916,N_5787);
xnor U7321 (N_7321,N_6181,N_3666);
xor U7322 (N_7322,N_5547,N_5998);
and U7323 (N_7323,N_3500,N_5673);
xor U7324 (N_7324,N_3703,N_6016);
nor U7325 (N_7325,N_5083,N_4050);
nand U7326 (N_7326,N_3811,N_3435);
and U7327 (N_7327,N_4000,N_5358);
nand U7328 (N_7328,N_3644,N_5906);
or U7329 (N_7329,N_5893,N_4080);
nand U7330 (N_7330,N_3953,N_3506);
xnor U7331 (N_7331,N_4797,N_3928);
xnor U7332 (N_7332,N_5618,N_5660);
nor U7333 (N_7333,N_4508,N_4998);
and U7334 (N_7334,N_3918,N_3424);
and U7335 (N_7335,N_4788,N_4403);
or U7336 (N_7336,N_5322,N_3183);
nand U7337 (N_7337,N_3393,N_3536);
nand U7338 (N_7338,N_3386,N_3433);
nand U7339 (N_7339,N_5324,N_5907);
xnor U7340 (N_7340,N_4929,N_4982);
nor U7341 (N_7341,N_3294,N_4795);
nor U7342 (N_7342,N_6234,N_5140);
nor U7343 (N_7343,N_5317,N_5116);
nand U7344 (N_7344,N_3510,N_6047);
nor U7345 (N_7345,N_3825,N_5175);
xnor U7346 (N_7346,N_5040,N_5745);
nand U7347 (N_7347,N_4831,N_5912);
and U7348 (N_7348,N_3596,N_3957);
or U7349 (N_7349,N_5514,N_6190);
and U7350 (N_7350,N_3669,N_4984);
xor U7351 (N_7351,N_4441,N_5644);
nor U7352 (N_7352,N_4861,N_3328);
and U7353 (N_7353,N_4761,N_5165);
nand U7354 (N_7354,N_6215,N_5526);
nor U7355 (N_7355,N_5538,N_3357);
and U7356 (N_7356,N_3631,N_3923);
nand U7357 (N_7357,N_3355,N_6034);
or U7358 (N_7358,N_4656,N_4490);
and U7359 (N_7359,N_4853,N_5459);
and U7360 (N_7360,N_4215,N_6194);
nor U7361 (N_7361,N_5719,N_5270);
xnor U7362 (N_7362,N_4197,N_4114);
nor U7363 (N_7363,N_3932,N_4714);
nor U7364 (N_7364,N_3814,N_5914);
or U7365 (N_7365,N_3460,N_4937);
and U7366 (N_7366,N_5642,N_6035);
xor U7367 (N_7367,N_3599,N_5455);
nor U7368 (N_7368,N_3963,N_6244);
nand U7369 (N_7369,N_5166,N_4766);
xnor U7370 (N_7370,N_5532,N_3766);
and U7371 (N_7371,N_4111,N_4851);
xor U7372 (N_7372,N_4272,N_4735);
xnor U7373 (N_7373,N_5699,N_3589);
nor U7374 (N_7374,N_4469,N_4810);
or U7375 (N_7375,N_6195,N_4281);
xnor U7376 (N_7376,N_6022,N_3875);
nor U7377 (N_7377,N_3540,N_3309);
or U7378 (N_7378,N_3245,N_4158);
nor U7379 (N_7379,N_3602,N_5717);
nand U7380 (N_7380,N_5693,N_5974);
and U7381 (N_7381,N_4849,N_3332);
nor U7382 (N_7382,N_6159,N_4988);
and U7383 (N_7383,N_3452,N_3915);
and U7384 (N_7384,N_5918,N_3870);
xnor U7385 (N_7385,N_5978,N_3175);
nor U7386 (N_7386,N_3782,N_4739);
and U7387 (N_7387,N_3761,N_4627);
nand U7388 (N_7388,N_4053,N_5443);
nor U7389 (N_7389,N_6222,N_3220);
and U7390 (N_7390,N_5020,N_5701);
and U7391 (N_7391,N_3401,N_5284);
and U7392 (N_7392,N_5877,N_6160);
or U7393 (N_7393,N_3561,N_4360);
or U7394 (N_7394,N_4593,N_4919);
or U7395 (N_7395,N_4302,N_4837);
nand U7396 (N_7396,N_3526,N_5690);
and U7397 (N_7397,N_5938,N_5397);
and U7398 (N_7398,N_4830,N_4655);
xor U7399 (N_7399,N_3827,N_3404);
or U7400 (N_7400,N_4780,N_3652);
xnor U7401 (N_7401,N_5197,N_3988);
or U7402 (N_7402,N_4973,N_5647);
nor U7403 (N_7403,N_3595,N_5309);
nand U7404 (N_7404,N_6247,N_3547);
nor U7405 (N_7405,N_4948,N_4678);
and U7406 (N_7406,N_4166,N_5084);
nand U7407 (N_7407,N_4258,N_5671);
nand U7408 (N_7408,N_4350,N_3756);
or U7409 (N_7409,N_3877,N_4382);
xnor U7410 (N_7410,N_6158,N_3994);
nand U7411 (N_7411,N_5703,N_5394);
nor U7412 (N_7412,N_4936,N_5574);
xor U7413 (N_7413,N_5516,N_6156);
nor U7414 (N_7414,N_6240,N_3662);
xor U7415 (N_7415,N_4902,N_4072);
nor U7416 (N_7416,N_4473,N_3576);
and U7417 (N_7417,N_3364,N_4146);
or U7418 (N_7418,N_5658,N_3527);
or U7419 (N_7419,N_5494,N_3173);
or U7420 (N_7420,N_4225,N_4294);
and U7421 (N_7421,N_3244,N_4293);
xor U7422 (N_7422,N_3645,N_3985);
nand U7423 (N_7423,N_3372,N_5188);
nand U7424 (N_7424,N_4507,N_5696);
xor U7425 (N_7425,N_3418,N_4854);
nor U7426 (N_7426,N_5531,N_5267);
nand U7427 (N_7427,N_5557,N_3955);
or U7428 (N_7428,N_5688,N_3922);
or U7429 (N_7429,N_4512,N_3140);
xor U7430 (N_7430,N_5372,N_4619);
xnor U7431 (N_7431,N_4947,N_5217);
xor U7432 (N_7432,N_4385,N_5773);
nand U7433 (N_7433,N_5753,N_6152);
nor U7434 (N_7434,N_6095,N_5151);
nor U7435 (N_7435,N_4583,N_3343);
xor U7436 (N_7436,N_3238,N_3682);
nand U7437 (N_7437,N_3836,N_4454);
nor U7438 (N_7438,N_3925,N_5697);
nor U7439 (N_7439,N_3887,N_3126);
xnor U7440 (N_7440,N_4148,N_6083);
xnor U7441 (N_7441,N_3184,N_5924);
xor U7442 (N_7442,N_5398,N_6103);
nor U7443 (N_7443,N_4077,N_3992);
nor U7444 (N_7444,N_3586,N_6091);
xor U7445 (N_7445,N_5801,N_5392);
and U7446 (N_7446,N_3812,N_5478);
nor U7447 (N_7447,N_3962,N_5308);
or U7448 (N_7448,N_4526,N_5081);
nor U7449 (N_7449,N_4605,N_4562);
nor U7450 (N_7450,N_5541,N_5156);
or U7451 (N_7451,N_4359,N_6171);
and U7452 (N_7452,N_6141,N_4047);
xnor U7453 (N_7453,N_6199,N_3311);
or U7454 (N_7454,N_4890,N_4277);
xor U7455 (N_7455,N_5859,N_6136);
nor U7456 (N_7456,N_5230,N_3530);
nand U7457 (N_7457,N_5361,N_5278);
or U7458 (N_7458,N_4794,N_5422);
xnor U7459 (N_7459,N_4751,N_3855);
nand U7460 (N_7460,N_3439,N_5496);
xnor U7461 (N_7461,N_5004,N_5577);
or U7462 (N_7462,N_4193,N_5325);
nor U7463 (N_7463,N_4626,N_5720);
xnor U7464 (N_7464,N_4343,N_5933);
or U7465 (N_7465,N_4702,N_3947);
and U7466 (N_7466,N_5782,N_6187);
and U7467 (N_7467,N_3482,N_3422);
and U7468 (N_7468,N_5968,N_3617);
and U7469 (N_7469,N_3376,N_5940);
nand U7470 (N_7470,N_5152,N_4446);
or U7471 (N_7471,N_3771,N_4100);
and U7472 (N_7472,N_4682,N_4807);
and U7473 (N_7473,N_3713,N_3768);
and U7474 (N_7474,N_5979,N_5077);
or U7475 (N_7475,N_5791,N_5996);
xor U7476 (N_7476,N_4190,N_3398);
xnor U7477 (N_7477,N_4996,N_4564);
xor U7478 (N_7478,N_5335,N_3368);
nor U7479 (N_7479,N_5985,N_5810);
and U7480 (N_7480,N_4920,N_4292);
nor U7481 (N_7481,N_6204,N_3575);
nor U7482 (N_7482,N_3648,N_4405);
nand U7483 (N_7483,N_4150,N_5653);
and U7484 (N_7484,N_3316,N_3858);
nand U7485 (N_7485,N_3239,N_4848);
nor U7486 (N_7486,N_5505,N_6184);
nor U7487 (N_7487,N_5876,N_3161);
xor U7488 (N_7488,N_4677,N_5672);
xor U7489 (N_7489,N_3525,N_5115);
nor U7490 (N_7490,N_5587,N_3429);
nor U7491 (N_7491,N_3700,N_5920);
or U7492 (N_7492,N_3551,N_3480);
nand U7493 (N_7493,N_6239,N_4442);
nor U7494 (N_7494,N_5725,N_3178);
and U7495 (N_7495,N_5402,N_4521);
or U7496 (N_7496,N_5250,N_3410);
and U7497 (N_7497,N_4553,N_3676);
and U7498 (N_7498,N_4900,N_5766);
nor U7499 (N_7499,N_4731,N_5602);
nand U7500 (N_7500,N_5200,N_3748);
xor U7501 (N_7501,N_4309,N_3462);
or U7502 (N_7502,N_5263,N_4376);
nor U7503 (N_7503,N_3726,N_5798);
or U7504 (N_7504,N_4465,N_5476);
or U7505 (N_7505,N_4344,N_3362);
xnor U7506 (N_7506,N_5095,N_3210);
or U7507 (N_7507,N_6144,N_3385);
and U7508 (N_7508,N_4089,N_5075);
xor U7509 (N_7509,N_4078,N_4632);
and U7510 (N_7510,N_3893,N_3369);
nor U7511 (N_7511,N_3251,N_4585);
nand U7512 (N_7512,N_5406,N_4182);
nand U7513 (N_7513,N_5187,N_5100);
xnor U7514 (N_7514,N_3899,N_5862);
nor U7515 (N_7515,N_5261,N_3841);
and U7516 (N_7516,N_3773,N_3685);
and U7517 (N_7517,N_3972,N_4204);
nor U7518 (N_7518,N_4377,N_5446);
or U7519 (N_7519,N_4262,N_6040);
nor U7520 (N_7520,N_5139,N_4871);
nor U7521 (N_7521,N_3151,N_3608);
xnor U7522 (N_7522,N_5584,N_5570);
or U7523 (N_7523,N_5057,N_3415);
xor U7524 (N_7524,N_3620,N_3872);
nand U7525 (N_7525,N_3336,N_5390);
or U7526 (N_7526,N_5748,N_3405);
xor U7527 (N_7527,N_5863,N_4511);
or U7528 (N_7528,N_4042,N_6161);
nand U7529 (N_7529,N_6118,N_4980);
and U7530 (N_7530,N_5983,N_5183);
and U7531 (N_7531,N_5965,N_3366);
and U7532 (N_7532,N_5632,N_5955);
xor U7533 (N_7533,N_3687,N_3792);
nand U7534 (N_7534,N_3643,N_3206);
nand U7535 (N_7535,N_3272,N_4310);
and U7536 (N_7536,N_4529,N_4917);
xor U7537 (N_7537,N_3688,N_4954);
nand U7538 (N_7538,N_3465,N_6201);
nand U7539 (N_7539,N_4123,N_4017);
nand U7540 (N_7540,N_5905,N_5093);
nor U7541 (N_7541,N_4864,N_3234);
and U7542 (N_7542,N_3777,N_4886);
or U7543 (N_7543,N_3260,N_5431);
xnor U7544 (N_7544,N_4404,N_4133);
nand U7545 (N_7545,N_5072,N_6006);
or U7546 (N_7546,N_3254,N_5306);
xnor U7547 (N_7547,N_3787,N_5272);
or U7548 (N_7548,N_5835,N_4775);
and U7549 (N_7549,N_5221,N_6198);
or U7550 (N_7550,N_4971,N_3690);
and U7551 (N_7551,N_5900,N_4662);
or U7552 (N_7552,N_4392,N_3209);
nor U7553 (N_7553,N_3441,N_3193);
nand U7554 (N_7554,N_4295,N_3856);
xor U7555 (N_7555,N_3421,N_4742);
nand U7556 (N_7556,N_4297,N_3714);
nor U7557 (N_7557,N_5783,N_5488);
and U7558 (N_7558,N_5276,N_4664);
nand U7559 (N_7559,N_4768,N_3413);
nor U7560 (N_7560,N_4222,N_4026);
nor U7561 (N_7561,N_3531,N_5310);
or U7562 (N_7562,N_5796,N_3541);
or U7563 (N_7563,N_4999,N_5555);
and U7564 (N_7564,N_3197,N_3293);
and U7565 (N_7565,N_4384,N_3400);
xnor U7566 (N_7566,N_5741,N_5792);
nor U7567 (N_7567,N_3427,N_6114);
or U7568 (N_7568,N_5173,N_4004);
and U7569 (N_7569,N_5967,N_5509);
xor U7570 (N_7570,N_5861,N_4288);
nor U7571 (N_7571,N_3273,N_4109);
or U7572 (N_7572,N_5074,N_5338);
and U7573 (N_7573,N_5440,N_3630);
nand U7574 (N_7574,N_5051,N_3276);
and U7575 (N_7575,N_3614,N_4482);
xor U7576 (N_7576,N_4823,N_3659);
and U7577 (N_7577,N_4443,N_5755);
or U7578 (N_7578,N_4138,N_4395);
xnor U7579 (N_7579,N_4505,N_4784);
and U7580 (N_7580,N_3830,N_4489);
and U7581 (N_7581,N_4945,N_5314);
or U7582 (N_7582,N_4068,N_3715);
and U7583 (N_7583,N_4092,N_4963);
xnor U7584 (N_7584,N_6213,N_4370);
nor U7585 (N_7585,N_4647,N_5469);
nand U7586 (N_7586,N_3568,N_5374);
xor U7587 (N_7587,N_4108,N_3786);
and U7588 (N_7588,N_5420,N_5262);
nand U7589 (N_7589,N_5371,N_3654);
nor U7590 (N_7590,N_3665,N_3868);
or U7591 (N_7591,N_4348,N_3705);
xor U7592 (N_7592,N_5549,N_5501);
nand U7593 (N_7593,N_3132,N_3300);
and U7594 (N_7594,N_4997,N_4452);
nor U7595 (N_7595,N_5063,N_4364);
nor U7596 (N_7596,N_6166,N_3458);
nor U7597 (N_7597,N_5581,N_3256);
nand U7598 (N_7598,N_5708,N_4051);
xnor U7599 (N_7599,N_4394,N_5931);
nand U7600 (N_7600,N_4014,N_4594);
nor U7601 (N_7601,N_5273,N_4464);
nor U7602 (N_7602,N_6145,N_3345);
nor U7603 (N_7603,N_4279,N_4501);
and U7604 (N_7604,N_4159,N_5497);
and U7605 (N_7605,N_5313,N_4926);
or U7606 (N_7606,N_4161,N_5196);
nand U7607 (N_7607,N_4030,N_3795);
or U7608 (N_7608,N_5311,N_5492);
and U7609 (N_7609,N_5821,N_4037);
nand U7610 (N_7610,N_4227,N_3459);
or U7611 (N_7611,N_3991,N_6210);
or U7612 (N_7612,N_5464,N_5147);
and U7613 (N_7613,N_5043,N_5017);
xnor U7614 (N_7614,N_6019,N_3291);
xor U7615 (N_7615,N_6146,N_5937);
and U7616 (N_7616,N_5363,N_3653);
xor U7617 (N_7617,N_6200,N_3639);
nor U7618 (N_7618,N_3383,N_5625);
xnor U7619 (N_7619,N_4154,N_6173);
xnor U7620 (N_7620,N_3542,N_5354);
nand U7621 (N_7621,N_5097,N_3592);
xor U7622 (N_7622,N_5008,N_6002);
or U7623 (N_7623,N_6132,N_3894);
or U7624 (N_7624,N_3625,N_4285);
nand U7625 (N_7625,N_3622,N_5023);
and U7626 (N_7626,N_3671,N_4953);
and U7627 (N_7627,N_5848,N_5738);
and U7628 (N_7628,N_5222,N_4379);
nor U7629 (N_7629,N_3727,N_5515);
xnor U7630 (N_7630,N_4467,N_5092);
nand U7631 (N_7631,N_4349,N_5211);
xnor U7632 (N_7632,N_5867,N_4437);
and U7633 (N_7633,N_5242,N_5474);
nand U7634 (N_7634,N_3223,N_5157);
nand U7635 (N_7635,N_4495,N_3520);
xor U7636 (N_7636,N_3591,N_4168);
nand U7637 (N_7637,N_3675,N_3185);
and U7638 (N_7638,N_5623,N_5327);
nand U7639 (N_7639,N_4804,N_4738);
nand U7640 (N_7640,N_3388,N_4125);
nor U7641 (N_7641,N_4316,N_5686);
and U7642 (N_7642,N_4703,N_3484);
xnor U7643 (N_7643,N_6124,N_5649);
and U7644 (N_7644,N_5579,N_4430);
or U7645 (N_7645,N_6164,N_3319);
nand U7646 (N_7646,N_5939,N_5158);
or U7647 (N_7647,N_4246,N_4132);
or U7648 (N_7648,N_4815,N_4362);
xor U7649 (N_7649,N_5473,N_4669);
and U7650 (N_7650,N_5944,N_4545);
or U7651 (N_7651,N_3125,N_3479);
or U7652 (N_7652,N_5007,N_3728);
nand U7653 (N_7653,N_6133,N_4357);
and U7654 (N_7654,N_4199,N_5826);
nand U7655 (N_7655,N_6008,N_4907);
xor U7656 (N_7656,N_3470,N_3902);
or U7657 (N_7657,N_3190,N_4935);
and U7658 (N_7658,N_3601,N_5033);
nand U7659 (N_7659,N_5565,N_3910);
xnor U7660 (N_7660,N_3176,N_3864);
and U7661 (N_7661,N_4510,N_6101);
xnor U7662 (N_7662,N_3945,N_5774);
or U7663 (N_7663,N_3767,N_6057);
nor U7664 (N_7664,N_4904,N_4707);
nand U7665 (N_7665,N_5411,N_5206);
and U7666 (N_7666,N_5456,N_6241);
nor U7667 (N_7667,N_3752,N_5366);
or U7668 (N_7668,N_6074,N_4088);
nor U7669 (N_7669,N_5337,N_4184);
or U7670 (N_7670,N_5113,N_4834);
xor U7671 (N_7671,N_4573,N_4790);
or U7672 (N_7672,N_6154,N_5831);
or U7673 (N_7673,N_3744,N_4079);
nand U7674 (N_7674,N_4903,N_5285);
nor U7675 (N_7675,N_4674,N_5135);
nor U7676 (N_7676,N_4326,N_5729);
xor U7677 (N_7677,N_3615,N_5413);
and U7678 (N_7678,N_4628,N_3409);
nand U7679 (N_7679,N_3313,N_5177);
nor U7680 (N_7680,N_3898,N_5529);
and U7681 (N_7681,N_3285,N_4772);
xnor U7682 (N_7682,N_4325,N_4198);
nor U7683 (N_7683,N_3754,N_5716);
nand U7684 (N_7684,N_5884,N_4765);
nor U7685 (N_7685,N_4852,N_5236);
xnor U7686 (N_7686,N_4502,N_4556);
or U7687 (N_7687,N_5809,N_5913);
nand U7688 (N_7688,N_6131,N_5504);
nand U7689 (N_7689,N_3657,N_4011);
nor U7690 (N_7690,N_3549,N_3550);
or U7691 (N_7691,N_5522,N_4786);
and U7692 (N_7692,N_5739,N_4264);
xnor U7693 (N_7693,N_5573,N_4922);
nor U7694 (N_7694,N_4747,N_4414);
xnor U7695 (N_7695,N_5819,N_5793);
nor U7696 (N_7696,N_5621,N_4541);
and U7697 (N_7697,N_4860,N_3146);
nor U7698 (N_7698,N_5919,N_4578);
xnor U7699 (N_7699,N_5146,N_5839);
and U7700 (N_7700,N_4396,N_3334);
or U7701 (N_7701,N_5260,N_4841);
or U7702 (N_7702,N_3492,N_3912);
xor U7703 (N_7703,N_3344,N_4581);
or U7704 (N_7704,N_6030,N_5752);
xor U7705 (N_7705,N_5662,N_4801);
and U7706 (N_7706,N_5698,N_4701);
xor U7707 (N_7707,N_5229,N_5535);
nand U7708 (N_7708,N_3567,N_5186);
nor U7709 (N_7709,N_3331,N_4942);
nor U7710 (N_7710,N_4163,N_4486);
nor U7711 (N_7711,N_4705,N_4985);
xnor U7712 (N_7712,N_4575,N_4013);
and U7713 (N_7713,N_5923,N_4856);
nand U7714 (N_7714,N_5493,N_4003);
nor U7715 (N_7715,N_5015,N_5212);
and U7716 (N_7716,N_3584,N_4426);
nand U7717 (N_7717,N_4422,N_4990);
nor U7718 (N_7718,N_3660,N_5428);
nor U7719 (N_7719,N_4439,N_3242);
or U7720 (N_7720,N_5064,N_5258);
nor U7721 (N_7721,N_3145,N_3838);
or U7722 (N_7722,N_4492,N_3642);
nor U7723 (N_7723,N_3585,N_4623);
and U7724 (N_7724,N_5713,N_4280);
xnor U7725 (N_7725,N_3320,N_5395);
nor U7726 (N_7726,N_4367,N_3365);
nor U7727 (N_7727,N_3783,N_5331);
and U7728 (N_7728,N_5091,N_4698);
nor U7729 (N_7729,N_3975,N_6185);
xor U7730 (N_7730,N_6191,N_5490);
or U7731 (N_7731,N_3231,N_3882);
and U7732 (N_7732,N_4363,N_3181);
nand U7733 (N_7733,N_4413,N_3913);
xor U7734 (N_7734,N_5966,N_5627);
nand U7735 (N_7735,N_3747,N_5881);
nor U7736 (N_7736,N_3965,N_4710);
nor U7737 (N_7737,N_3142,N_6017);
and U7738 (N_7738,N_5153,N_6014);
nand U7739 (N_7739,N_3494,N_3628);
and U7740 (N_7740,N_5010,N_4099);
xnor U7741 (N_7741,N_5096,N_5006);
nand U7742 (N_7742,N_5875,N_5301);
and U7743 (N_7743,N_3411,N_3861);
xnor U7744 (N_7744,N_5715,N_3469);
nand U7745 (N_7745,N_4881,N_6038);
nor U7746 (N_7746,N_3138,N_4323);
nor U7747 (N_7747,N_5036,N_5511);
nand U7748 (N_7748,N_5299,N_6227);
xnor U7749 (N_7749,N_3302,N_4777);
and U7750 (N_7750,N_5667,N_6050);
nor U7751 (N_7751,N_4862,N_5961);
nor U7752 (N_7752,N_4538,N_5087);
xor U7753 (N_7753,N_3148,N_3564);
xor U7754 (N_7754,N_5941,N_3224);
nand U7755 (N_7755,N_4035,N_3977);
and U7756 (N_7756,N_4300,N_5883);
and U7757 (N_7757,N_5909,N_5718);
nor U7758 (N_7758,N_3566,N_5899);
nand U7759 (N_7759,N_4411,N_6218);
and U7760 (N_7760,N_3350,N_3298);
xnor U7761 (N_7761,N_4120,N_4757);
or U7762 (N_7762,N_4524,N_6106);
xor U7763 (N_7763,N_6192,N_5500);
and U7764 (N_7764,N_3532,N_3262);
nand U7765 (N_7765,N_4588,N_6023);
nor U7766 (N_7766,N_4335,N_5119);
and U7767 (N_7767,N_3764,N_5009);
nand U7768 (N_7768,N_3544,N_4249);
xor U7769 (N_7769,N_5737,N_4270);
nand U7770 (N_7770,N_5543,N_3545);
nor U7771 (N_7771,N_5447,N_5167);
nor U7772 (N_7772,N_4785,N_5367);
nand U7773 (N_7773,N_5386,N_3745);
xnor U7774 (N_7774,N_3634,N_4393);
or U7775 (N_7775,N_4549,N_4122);
or U7776 (N_7776,N_3637,N_6219);
or U7777 (N_7777,N_6151,N_5929);
nand U7778 (N_7778,N_5025,N_4675);
nor U7779 (N_7779,N_3667,N_5182);
nor U7780 (N_7780,N_5079,N_5450);
nand U7781 (N_7781,N_6027,N_5695);
nor U7782 (N_7782,N_5994,N_5613);
xor U7783 (N_7783,N_5110,N_5670);
nand U7784 (N_7784,N_3483,N_4408);
and U7785 (N_7785,N_3367,N_3778);
xnor U7786 (N_7786,N_5689,N_4341);
xor U7787 (N_7787,N_5240,N_5105);
and U7788 (N_7788,N_3522,N_4263);
xor U7789 (N_7789,N_4428,N_3384);
and U7790 (N_7790,N_5754,N_4622);
xor U7791 (N_7791,N_5144,N_4153);
xnor U7792 (N_7792,N_4269,N_4278);
and U7793 (N_7793,N_6207,N_3406);
nand U7794 (N_7794,N_5283,N_5594);
xor U7795 (N_7795,N_6061,N_3995);
xnor U7796 (N_7796,N_4143,N_5894);
nor U7797 (N_7797,N_5026,N_3702);
and U7798 (N_7798,N_5102,N_3155);
nand U7799 (N_7799,N_5639,N_3518);
nor U7800 (N_7800,N_3221,N_4613);
xor U7801 (N_7801,N_3960,N_4210);
xnor U7802 (N_7802,N_4209,N_5245);
or U7803 (N_7803,N_5502,N_5014);
xnor U7804 (N_7804,N_4238,N_4809);
nor U7805 (N_7805,N_5856,N_5645);
and U7806 (N_7806,N_4730,N_4609);
and U7807 (N_7807,N_3729,N_4686);
nor U7808 (N_7808,N_3943,N_4257);
or U7809 (N_7809,N_3695,N_3289);
and U7810 (N_7810,N_6235,N_3621);
nor U7811 (N_7811,N_3683,N_5353);
xnor U7812 (N_7812,N_5304,N_3208);
xnor U7813 (N_7813,N_4724,N_3356);
nor U7814 (N_7814,N_4249,N_4536);
nand U7815 (N_7815,N_5296,N_4811);
and U7816 (N_7816,N_4085,N_5038);
or U7817 (N_7817,N_4942,N_3657);
xor U7818 (N_7818,N_4217,N_5855);
nor U7819 (N_7819,N_5313,N_4394);
or U7820 (N_7820,N_4686,N_5762);
and U7821 (N_7821,N_3297,N_6245);
nand U7822 (N_7822,N_5108,N_3413);
xor U7823 (N_7823,N_4774,N_5345);
or U7824 (N_7824,N_3246,N_5992);
nand U7825 (N_7825,N_3460,N_5642);
xnor U7826 (N_7826,N_3770,N_5382);
or U7827 (N_7827,N_4793,N_4092);
and U7828 (N_7828,N_6127,N_4456);
nor U7829 (N_7829,N_5404,N_4852);
xnor U7830 (N_7830,N_5232,N_4887);
nand U7831 (N_7831,N_5057,N_5390);
xor U7832 (N_7832,N_3445,N_3570);
and U7833 (N_7833,N_5330,N_3676);
xor U7834 (N_7834,N_4976,N_4347);
nor U7835 (N_7835,N_5493,N_5375);
and U7836 (N_7836,N_5834,N_4949);
xor U7837 (N_7837,N_5341,N_3247);
nand U7838 (N_7838,N_4530,N_3397);
or U7839 (N_7839,N_4309,N_4625);
nor U7840 (N_7840,N_6156,N_3960);
nand U7841 (N_7841,N_5496,N_4612);
or U7842 (N_7842,N_3878,N_4288);
xnor U7843 (N_7843,N_4357,N_4433);
nand U7844 (N_7844,N_4952,N_3570);
xor U7845 (N_7845,N_4768,N_5091);
and U7846 (N_7846,N_3715,N_5374);
nor U7847 (N_7847,N_3665,N_4053);
nor U7848 (N_7848,N_5692,N_4903);
nor U7849 (N_7849,N_3154,N_5521);
or U7850 (N_7850,N_4123,N_3681);
and U7851 (N_7851,N_4527,N_6087);
and U7852 (N_7852,N_3583,N_3419);
xor U7853 (N_7853,N_5142,N_3141);
nor U7854 (N_7854,N_5937,N_5099);
xor U7855 (N_7855,N_5954,N_4209);
or U7856 (N_7856,N_3715,N_3203);
nand U7857 (N_7857,N_3764,N_3684);
nand U7858 (N_7858,N_5998,N_6125);
and U7859 (N_7859,N_5164,N_5619);
nand U7860 (N_7860,N_5670,N_5933);
nor U7861 (N_7861,N_3923,N_3151);
nor U7862 (N_7862,N_4849,N_4560);
nor U7863 (N_7863,N_4133,N_4202);
or U7864 (N_7864,N_4817,N_3683);
xnor U7865 (N_7865,N_5281,N_3970);
or U7866 (N_7866,N_3822,N_3985);
and U7867 (N_7867,N_5372,N_4417);
or U7868 (N_7868,N_4723,N_5740);
or U7869 (N_7869,N_4676,N_5408);
and U7870 (N_7870,N_4512,N_5777);
xnor U7871 (N_7871,N_4153,N_4240);
nor U7872 (N_7872,N_4284,N_6177);
xor U7873 (N_7873,N_5677,N_4943);
nor U7874 (N_7874,N_5471,N_4417);
or U7875 (N_7875,N_5374,N_4029);
and U7876 (N_7876,N_5068,N_4105);
nand U7877 (N_7877,N_6081,N_5090);
nor U7878 (N_7878,N_4503,N_6109);
xnor U7879 (N_7879,N_5023,N_6209);
nor U7880 (N_7880,N_4790,N_5492);
nand U7881 (N_7881,N_5988,N_6093);
and U7882 (N_7882,N_3996,N_5859);
nor U7883 (N_7883,N_6119,N_3763);
and U7884 (N_7884,N_4277,N_6082);
nor U7885 (N_7885,N_4338,N_3562);
or U7886 (N_7886,N_3488,N_5310);
or U7887 (N_7887,N_6123,N_4953);
xor U7888 (N_7888,N_3869,N_4425);
nand U7889 (N_7889,N_4829,N_4345);
nand U7890 (N_7890,N_3285,N_4822);
or U7891 (N_7891,N_4993,N_3792);
and U7892 (N_7892,N_4406,N_4201);
nand U7893 (N_7893,N_6033,N_3743);
nand U7894 (N_7894,N_5899,N_4678);
and U7895 (N_7895,N_5478,N_5061);
nand U7896 (N_7896,N_5621,N_5850);
and U7897 (N_7897,N_4496,N_4627);
nand U7898 (N_7898,N_4128,N_5971);
xor U7899 (N_7899,N_3791,N_3949);
xnor U7900 (N_7900,N_3527,N_3616);
or U7901 (N_7901,N_5052,N_3844);
or U7902 (N_7902,N_3700,N_3913);
and U7903 (N_7903,N_3341,N_6214);
nand U7904 (N_7904,N_3289,N_5654);
or U7905 (N_7905,N_4013,N_4429);
nand U7906 (N_7906,N_5789,N_3401);
xnor U7907 (N_7907,N_5061,N_4505);
or U7908 (N_7908,N_4940,N_4869);
xor U7909 (N_7909,N_5502,N_3230);
and U7910 (N_7910,N_4247,N_3853);
nor U7911 (N_7911,N_4191,N_3384);
nand U7912 (N_7912,N_3842,N_4971);
or U7913 (N_7913,N_4687,N_4067);
and U7914 (N_7914,N_3395,N_4349);
xor U7915 (N_7915,N_4884,N_3624);
xor U7916 (N_7916,N_4856,N_6124);
nand U7917 (N_7917,N_4228,N_5111);
xnor U7918 (N_7918,N_5738,N_4994);
or U7919 (N_7919,N_4998,N_4683);
or U7920 (N_7920,N_4945,N_4814);
nand U7921 (N_7921,N_6151,N_6124);
xor U7922 (N_7922,N_3189,N_6145);
xor U7923 (N_7923,N_6208,N_5850);
nand U7924 (N_7924,N_5685,N_5968);
xor U7925 (N_7925,N_6010,N_5874);
xnor U7926 (N_7926,N_4865,N_4816);
or U7927 (N_7927,N_4134,N_5561);
nand U7928 (N_7928,N_4565,N_4520);
nor U7929 (N_7929,N_5633,N_4940);
nor U7930 (N_7930,N_4799,N_4868);
xor U7931 (N_7931,N_5076,N_3975);
xnor U7932 (N_7932,N_5242,N_4318);
nand U7933 (N_7933,N_4709,N_3733);
nor U7934 (N_7934,N_3137,N_3943);
xnor U7935 (N_7935,N_4732,N_5253);
xor U7936 (N_7936,N_4422,N_5931);
xnor U7937 (N_7937,N_5132,N_4749);
and U7938 (N_7938,N_5882,N_4607);
and U7939 (N_7939,N_4068,N_5834);
nand U7940 (N_7940,N_3334,N_5813);
xnor U7941 (N_7941,N_3853,N_3742);
xnor U7942 (N_7942,N_3506,N_4953);
or U7943 (N_7943,N_5619,N_4384);
nor U7944 (N_7944,N_5154,N_3412);
and U7945 (N_7945,N_5266,N_4909);
xnor U7946 (N_7946,N_4973,N_3682);
and U7947 (N_7947,N_4822,N_3828);
xor U7948 (N_7948,N_3930,N_4994);
or U7949 (N_7949,N_3210,N_4334);
and U7950 (N_7950,N_4684,N_5449);
nand U7951 (N_7951,N_5634,N_4530);
or U7952 (N_7952,N_5043,N_6216);
xor U7953 (N_7953,N_5160,N_5344);
and U7954 (N_7954,N_3501,N_3464);
xnor U7955 (N_7955,N_5308,N_5489);
or U7956 (N_7956,N_3316,N_5621);
xor U7957 (N_7957,N_4623,N_5006);
or U7958 (N_7958,N_5853,N_3786);
and U7959 (N_7959,N_3480,N_3310);
nor U7960 (N_7960,N_6052,N_5899);
and U7961 (N_7961,N_6046,N_5323);
nand U7962 (N_7962,N_4248,N_3452);
nand U7963 (N_7963,N_5007,N_4420);
xnor U7964 (N_7964,N_3762,N_4816);
xnor U7965 (N_7965,N_3345,N_4864);
nand U7966 (N_7966,N_6114,N_5702);
xor U7967 (N_7967,N_4869,N_5680);
xor U7968 (N_7968,N_5665,N_4755);
and U7969 (N_7969,N_4460,N_3390);
nand U7970 (N_7970,N_4673,N_3249);
xor U7971 (N_7971,N_3477,N_4877);
nand U7972 (N_7972,N_4231,N_3825);
xnor U7973 (N_7973,N_5202,N_4120);
and U7974 (N_7974,N_6112,N_6160);
xnor U7975 (N_7975,N_3295,N_3950);
and U7976 (N_7976,N_4123,N_3401);
xor U7977 (N_7977,N_4772,N_3594);
or U7978 (N_7978,N_3573,N_5672);
nor U7979 (N_7979,N_5174,N_3198);
and U7980 (N_7980,N_3558,N_5859);
and U7981 (N_7981,N_3367,N_3490);
or U7982 (N_7982,N_5808,N_3656);
nor U7983 (N_7983,N_5071,N_5074);
nand U7984 (N_7984,N_3721,N_5306);
nand U7985 (N_7985,N_4551,N_3925);
xnor U7986 (N_7986,N_3476,N_3308);
xnor U7987 (N_7987,N_5067,N_3976);
xnor U7988 (N_7988,N_5437,N_4401);
nand U7989 (N_7989,N_4011,N_5291);
xnor U7990 (N_7990,N_3999,N_4570);
xnor U7991 (N_7991,N_5091,N_4452);
and U7992 (N_7992,N_6184,N_3638);
or U7993 (N_7993,N_3468,N_4704);
nand U7994 (N_7994,N_6128,N_4777);
and U7995 (N_7995,N_6004,N_3579);
nand U7996 (N_7996,N_4085,N_5640);
xor U7997 (N_7997,N_3211,N_4082);
and U7998 (N_7998,N_4369,N_5727);
nor U7999 (N_7999,N_5407,N_5029);
nand U8000 (N_8000,N_3943,N_3951);
nor U8001 (N_8001,N_5502,N_4212);
nand U8002 (N_8002,N_5803,N_5297);
nand U8003 (N_8003,N_3495,N_3823);
xnor U8004 (N_8004,N_4573,N_4944);
and U8005 (N_8005,N_5250,N_4866);
and U8006 (N_8006,N_5937,N_3268);
xnor U8007 (N_8007,N_4956,N_5387);
or U8008 (N_8008,N_3963,N_3243);
or U8009 (N_8009,N_5417,N_3491);
xnor U8010 (N_8010,N_5234,N_5132);
nor U8011 (N_8011,N_5394,N_4927);
xnor U8012 (N_8012,N_3239,N_3429);
xnor U8013 (N_8013,N_3831,N_3649);
and U8014 (N_8014,N_5629,N_3320);
nor U8015 (N_8015,N_3247,N_4732);
xor U8016 (N_8016,N_5667,N_5729);
or U8017 (N_8017,N_5413,N_6155);
nand U8018 (N_8018,N_3450,N_5602);
xnor U8019 (N_8019,N_5888,N_5906);
xnor U8020 (N_8020,N_3209,N_4128);
and U8021 (N_8021,N_3391,N_5546);
and U8022 (N_8022,N_4195,N_5438);
or U8023 (N_8023,N_3948,N_4440);
or U8024 (N_8024,N_3673,N_5959);
nor U8025 (N_8025,N_5762,N_4645);
xnor U8026 (N_8026,N_4693,N_3457);
xnor U8027 (N_8027,N_4100,N_5675);
nand U8028 (N_8028,N_5117,N_4887);
or U8029 (N_8029,N_5343,N_6127);
and U8030 (N_8030,N_5855,N_5595);
xnor U8031 (N_8031,N_5870,N_5222);
nor U8032 (N_8032,N_3483,N_3158);
xor U8033 (N_8033,N_4270,N_6165);
nand U8034 (N_8034,N_5485,N_3448);
xnor U8035 (N_8035,N_6111,N_3281);
and U8036 (N_8036,N_4788,N_5482);
or U8037 (N_8037,N_3575,N_3336);
and U8038 (N_8038,N_5470,N_4486);
nand U8039 (N_8039,N_4662,N_6222);
nand U8040 (N_8040,N_4300,N_3216);
nand U8041 (N_8041,N_4618,N_4639);
xnor U8042 (N_8042,N_3695,N_5601);
or U8043 (N_8043,N_3932,N_5636);
xnor U8044 (N_8044,N_3359,N_4417);
or U8045 (N_8045,N_5540,N_3361);
nor U8046 (N_8046,N_3669,N_5185);
and U8047 (N_8047,N_6160,N_5490);
nor U8048 (N_8048,N_3611,N_4249);
nor U8049 (N_8049,N_4468,N_5356);
or U8050 (N_8050,N_6231,N_5692);
and U8051 (N_8051,N_5625,N_4165);
xor U8052 (N_8052,N_4230,N_3262);
and U8053 (N_8053,N_4022,N_4290);
or U8054 (N_8054,N_5709,N_5540);
nand U8055 (N_8055,N_5289,N_5746);
or U8056 (N_8056,N_3947,N_4202);
or U8057 (N_8057,N_5149,N_5479);
nand U8058 (N_8058,N_3315,N_3870);
nor U8059 (N_8059,N_4128,N_4145);
nor U8060 (N_8060,N_3978,N_4868);
xor U8061 (N_8061,N_3656,N_4473);
nor U8062 (N_8062,N_4920,N_5127);
nor U8063 (N_8063,N_5258,N_3696);
nor U8064 (N_8064,N_3648,N_4866);
nand U8065 (N_8065,N_6213,N_6157);
and U8066 (N_8066,N_5285,N_4573);
nor U8067 (N_8067,N_5096,N_5112);
nor U8068 (N_8068,N_4857,N_3126);
and U8069 (N_8069,N_5521,N_6179);
xnor U8070 (N_8070,N_4354,N_4951);
xor U8071 (N_8071,N_5301,N_3810);
and U8072 (N_8072,N_4579,N_3810);
xnor U8073 (N_8073,N_3227,N_3310);
and U8074 (N_8074,N_5929,N_4398);
nand U8075 (N_8075,N_3736,N_5838);
xnor U8076 (N_8076,N_5739,N_5669);
nor U8077 (N_8077,N_3274,N_4801);
nor U8078 (N_8078,N_4811,N_5956);
or U8079 (N_8079,N_5813,N_5615);
or U8080 (N_8080,N_3589,N_5402);
or U8081 (N_8081,N_3279,N_3502);
xor U8082 (N_8082,N_3625,N_4779);
or U8083 (N_8083,N_4337,N_4290);
xnor U8084 (N_8084,N_3171,N_6204);
and U8085 (N_8085,N_4003,N_3594);
or U8086 (N_8086,N_3234,N_4129);
and U8087 (N_8087,N_3422,N_4334);
xnor U8088 (N_8088,N_5870,N_4133);
or U8089 (N_8089,N_3788,N_3739);
xnor U8090 (N_8090,N_4153,N_5472);
xnor U8091 (N_8091,N_4913,N_4459);
nand U8092 (N_8092,N_3140,N_3377);
and U8093 (N_8093,N_5893,N_4969);
nor U8094 (N_8094,N_4705,N_4223);
and U8095 (N_8095,N_4769,N_3375);
or U8096 (N_8096,N_4091,N_5777);
and U8097 (N_8097,N_3923,N_5303);
nor U8098 (N_8098,N_6117,N_3408);
nand U8099 (N_8099,N_3442,N_3289);
or U8100 (N_8100,N_4379,N_5856);
nor U8101 (N_8101,N_4994,N_4835);
nor U8102 (N_8102,N_5741,N_5613);
nor U8103 (N_8103,N_5935,N_3998);
nor U8104 (N_8104,N_4562,N_5309);
and U8105 (N_8105,N_3184,N_3812);
or U8106 (N_8106,N_3682,N_3779);
or U8107 (N_8107,N_4499,N_5182);
or U8108 (N_8108,N_4790,N_4412);
or U8109 (N_8109,N_5530,N_4219);
or U8110 (N_8110,N_4727,N_5195);
nand U8111 (N_8111,N_5283,N_6123);
and U8112 (N_8112,N_5403,N_3855);
nand U8113 (N_8113,N_5677,N_5662);
xor U8114 (N_8114,N_3168,N_5863);
and U8115 (N_8115,N_4276,N_3264);
or U8116 (N_8116,N_6004,N_5541);
xor U8117 (N_8117,N_6187,N_3590);
or U8118 (N_8118,N_4765,N_3561);
and U8119 (N_8119,N_4614,N_5258);
nand U8120 (N_8120,N_3474,N_5718);
nor U8121 (N_8121,N_5514,N_4290);
nor U8122 (N_8122,N_3743,N_3195);
xnor U8123 (N_8123,N_6157,N_4794);
or U8124 (N_8124,N_3315,N_3837);
or U8125 (N_8125,N_3175,N_4602);
and U8126 (N_8126,N_4028,N_4694);
or U8127 (N_8127,N_3818,N_5092);
nor U8128 (N_8128,N_5221,N_3439);
and U8129 (N_8129,N_5751,N_3159);
nand U8130 (N_8130,N_3392,N_4243);
or U8131 (N_8131,N_3945,N_4502);
xor U8132 (N_8132,N_3643,N_5443);
nor U8133 (N_8133,N_3188,N_4644);
nor U8134 (N_8134,N_3171,N_5611);
nor U8135 (N_8135,N_6093,N_4318);
or U8136 (N_8136,N_4403,N_4743);
and U8137 (N_8137,N_3479,N_3523);
xor U8138 (N_8138,N_3276,N_5096);
nand U8139 (N_8139,N_6111,N_4116);
nor U8140 (N_8140,N_4449,N_4103);
nand U8141 (N_8141,N_6035,N_4732);
nand U8142 (N_8142,N_3431,N_4117);
and U8143 (N_8143,N_5497,N_3782);
nand U8144 (N_8144,N_4208,N_3314);
nor U8145 (N_8145,N_5158,N_6079);
xnor U8146 (N_8146,N_3195,N_3710);
or U8147 (N_8147,N_4973,N_5329);
and U8148 (N_8148,N_3310,N_5875);
nand U8149 (N_8149,N_3529,N_3795);
or U8150 (N_8150,N_5088,N_3899);
nor U8151 (N_8151,N_3598,N_5861);
nor U8152 (N_8152,N_5473,N_5813);
or U8153 (N_8153,N_5595,N_4906);
and U8154 (N_8154,N_4458,N_3514);
nor U8155 (N_8155,N_4083,N_4177);
xnor U8156 (N_8156,N_5799,N_5159);
and U8157 (N_8157,N_3264,N_5307);
xnor U8158 (N_8158,N_3571,N_6036);
nor U8159 (N_8159,N_6132,N_3216);
xor U8160 (N_8160,N_3344,N_3476);
nor U8161 (N_8161,N_4783,N_5786);
or U8162 (N_8162,N_3307,N_5152);
nor U8163 (N_8163,N_6086,N_5837);
and U8164 (N_8164,N_5871,N_3158);
nand U8165 (N_8165,N_3253,N_5026);
or U8166 (N_8166,N_4964,N_5169);
xnor U8167 (N_8167,N_5677,N_4726);
nor U8168 (N_8168,N_3279,N_3338);
or U8169 (N_8169,N_6132,N_4738);
nand U8170 (N_8170,N_4141,N_4064);
xnor U8171 (N_8171,N_3839,N_5293);
xor U8172 (N_8172,N_6163,N_6090);
or U8173 (N_8173,N_4424,N_4947);
or U8174 (N_8174,N_3366,N_5578);
and U8175 (N_8175,N_3426,N_5992);
xnor U8176 (N_8176,N_4861,N_4421);
and U8177 (N_8177,N_5967,N_3435);
xor U8178 (N_8178,N_5706,N_3751);
xnor U8179 (N_8179,N_3762,N_5991);
or U8180 (N_8180,N_3953,N_4386);
nor U8181 (N_8181,N_5930,N_4815);
xor U8182 (N_8182,N_6032,N_5846);
nor U8183 (N_8183,N_5097,N_3617);
xnor U8184 (N_8184,N_5686,N_4270);
nor U8185 (N_8185,N_3222,N_5749);
nor U8186 (N_8186,N_5191,N_4233);
xor U8187 (N_8187,N_4669,N_3256);
xor U8188 (N_8188,N_5727,N_5112);
nand U8189 (N_8189,N_5251,N_4947);
xnor U8190 (N_8190,N_5435,N_5994);
or U8191 (N_8191,N_3274,N_3451);
or U8192 (N_8192,N_6118,N_4706);
or U8193 (N_8193,N_5496,N_4615);
nor U8194 (N_8194,N_3981,N_4972);
and U8195 (N_8195,N_6022,N_3306);
and U8196 (N_8196,N_4686,N_5635);
xor U8197 (N_8197,N_5734,N_3154);
or U8198 (N_8198,N_4239,N_5755);
xor U8199 (N_8199,N_3930,N_6024);
nor U8200 (N_8200,N_5809,N_6243);
nor U8201 (N_8201,N_5451,N_5230);
and U8202 (N_8202,N_6245,N_3670);
xnor U8203 (N_8203,N_3129,N_4998);
nor U8204 (N_8204,N_5349,N_4319);
and U8205 (N_8205,N_5276,N_5526);
or U8206 (N_8206,N_3639,N_4212);
and U8207 (N_8207,N_6141,N_4425);
or U8208 (N_8208,N_3735,N_3967);
and U8209 (N_8209,N_3915,N_4455);
xnor U8210 (N_8210,N_5919,N_4885);
or U8211 (N_8211,N_4233,N_4619);
xnor U8212 (N_8212,N_4978,N_3146);
or U8213 (N_8213,N_5443,N_5966);
nand U8214 (N_8214,N_5782,N_3715);
nand U8215 (N_8215,N_4833,N_3197);
nor U8216 (N_8216,N_3833,N_5133);
nand U8217 (N_8217,N_5347,N_5650);
nand U8218 (N_8218,N_6015,N_4380);
and U8219 (N_8219,N_5498,N_3827);
and U8220 (N_8220,N_3459,N_4071);
or U8221 (N_8221,N_3424,N_6243);
or U8222 (N_8222,N_5297,N_3405);
nor U8223 (N_8223,N_5863,N_4363);
nand U8224 (N_8224,N_5719,N_4836);
and U8225 (N_8225,N_3432,N_4683);
nand U8226 (N_8226,N_5142,N_5906);
nand U8227 (N_8227,N_4962,N_5817);
and U8228 (N_8228,N_6045,N_5722);
or U8229 (N_8229,N_3771,N_4512);
xor U8230 (N_8230,N_3287,N_3732);
and U8231 (N_8231,N_3534,N_4747);
or U8232 (N_8232,N_5608,N_3317);
or U8233 (N_8233,N_3290,N_3309);
or U8234 (N_8234,N_5824,N_5898);
and U8235 (N_8235,N_4323,N_5570);
and U8236 (N_8236,N_4070,N_5752);
xor U8237 (N_8237,N_3983,N_5401);
or U8238 (N_8238,N_4340,N_3925);
xor U8239 (N_8239,N_3460,N_3349);
nand U8240 (N_8240,N_5179,N_6246);
or U8241 (N_8241,N_5241,N_4615);
and U8242 (N_8242,N_4609,N_3499);
nor U8243 (N_8243,N_5357,N_3189);
nor U8244 (N_8244,N_5061,N_5089);
nor U8245 (N_8245,N_3844,N_4144);
xnor U8246 (N_8246,N_4951,N_5120);
nand U8247 (N_8247,N_3879,N_4603);
xnor U8248 (N_8248,N_4470,N_4469);
nand U8249 (N_8249,N_4064,N_4449);
and U8250 (N_8250,N_3887,N_5621);
nand U8251 (N_8251,N_3129,N_4999);
nor U8252 (N_8252,N_3595,N_5492);
and U8253 (N_8253,N_3323,N_4818);
and U8254 (N_8254,N_4152,N_3305);
and U8255 (N_8255,N_3414,N_5941);
or U8256 (N_8256,N_4533,N_5042);
and U8257 (N_8257,N_5294,N_5469);
or U8258 (N_8258,N_4731,N_6150);
nand U8259 (N_8259,N_5412,N_4447);
nor U8260 (N_8260,N_5093,N_3207);
xor U8261 (N_8261,N_5731,N_5880);
and U8262 (N_8262,N_4438,N_5501);
xor U8263 (N_8263,N_5980,N_3365);
nand U8264 (N_8264,N_5647,N_3889);
nor U8265 (N_8265,N_3685,N_5249);
and U8266 (N_8266,N_4250,N_3528);
nand U8267 (N_8267,N_5080,N_4988);
xnor U8268 (N_8268,N_6048,N_3577);
xor U8269 (N_8269,N_5672,N_4865);
and U8270 (N_8270,N_4333,N_3801);
or U8271 (N_8271,N_5149,N_3134);
nor U8272 (N_8272,N_3202,N_3401);
nand U8273 (N_8273,N_4228,N_6218);
xor U8274 (N_8274,N_6164,N_3999);
xnor U8275 (N_8275,N_4667,N_6061);
nor U8276 (N_8276,N_4823,N_3132);
xnor U8277 (N_8277,N_3868,N_5732);
xnor U8278 (N_8278,N_4148,N_3456);
or U8279 (N_8279,N_5535,N_4340);
nor U8280 (N_8280,N_5837,N_5722);
xnor U8281 (N_8281,N_5488,N_4902);
and U8282 (N_8282,N_6010,N_3505);
nand U8283 (N_8283,N_6032,N_3844);
and U8284 (N_8284,N_5229,N_4166);
nand U8285 (N_8285,N_4118,N_3307);
or U8286 (N_8286,N_5348,N_3909);
nand U8287 (N_8287,N_5937,N_4310);
xor U8288 (N_8288,N_4561,N_5180);
nor U8289 (N_8289,N_3363,N_5745);
and U8290 (N_8290,N_5750,N_5947);
or U8291 (N_8291,N_5769,N_5118);
xor U8292 (N_8292,N_3252,N_5621);
nor U8293 (N_8293,N_6032,N_5619);
xor U8294 (N_8294,N_4506,N_3583);
or U8295 (N_8295,N_3778,N_3479);
or U8296 (N_8296,N_4252,N_5776);
nor U8297 (N_8297,N_4062,N_3754);
nor U8298 (N_8298,N_4071,N_5170);
nor U8299 (N_8299,N_5010,N_4643);
nor U8300 (N_8300,N_4831,N_4278);
and U8301 (N_8301,N_5123,N_3175);
or U8302 (N_8302,N_4111,N_6030);
xor U8303 (N_8303,N_6106,N_5396);
and U8304 (N_8304,N_4745,N_4051);
nand U8305 (N_8305,N_4055,N_4242);
and U8306 (N_8306,N_4678,N_5344);
xor U8307 (N_8307,N_3477,N_5104);
and U8308 (N_8308,N_4295,N_6109);
or U8309 (N_8309,N_5540,N_5090);
and U8310 (N_8310,N_3574,N_4744);
or U8311 (N_8311,N_5681,N_6163);
and U8312 (N_8312,N_4947,N_3311);
nor U8313 (N_8313,N_6039,N_4420);
nor U8314 (N_8314,N_5207,N_5468);
nor U8315 (N_8315,N_3813,N_3463);
xor U8316 (N_8316,N_5668,N_5903);
and U8317 (N_8317,N_3814,N_4070);
nor U8318 (N_8318,N_3501,N_4832);
nor U8319 (N_8319,N_3217,N_4109);
or U8320 (N_8320,N_5393,N_6236);
xor U8321 (N_8321,N_4885,N_4607);
or U8322 (N_8322,N_5945,N_5940);
or U8323 (N_8323,N_6220,N_5296);
nor U8324 (N_8324,N_5288,N_3885);
nand U8325 (N_8325,N_6131,N_3378);
nor U8326 (N_8326,N_3603,N_5389);
and U8327 (N_8327,N_5862,N_6201);
xor U8328 (N_8328,N_3759,N_3427);
or U8329 (N_8329,N_4298,N_4420);
nand U8330 (N_8330,N_5292,N_5316);
and U8331 (N_8331,N_6078,N_4925);
and U8332 (N_8332,N_4689,N_3193);
xor U8333 (N_8333,N_4169,N_3179);
or U8334 (N_8334,N_3579,N_3974);
nand U8335 (N_8335,N_3219,N_3349);
or U8336 (N_8336,N_6099,N_5701);
and U8337 (N_8337,N_4781,N_6197);
or U8338 (N_8338,N_5801,N_4567);
xor U8339 (N_8339,N_5398,N_5149);
nor U8340 (N_8340,N_5556,N_5252);
nand U8341 (N_8341,N_5593,N_3890);
xor U8342 (N_8342,N_5681,N_4366);
xnor U8343 (N_8343,N_4764,N_3780);
xor U8344 (N_8344,N_4444,N_3598);
or U8345 (N_8345,N_5853,N_6072);
nand U8346 (N_8346,N_4000,N_3157);
nor U8347 (N_8347,N_5235,N_3300);
and U8348 (N_8348,N_4064,N_4771);
or U8349 (N_8349,N_3922,N_6043);
nand U8350 (N_8350,N_4169,N_3407);
and U8351 (N_8351,N_4558,N_5989);
nand U8352 (N_8352,N_6008,N_3169);
and U8353 (N_8353,N_5397,N_4920);
and U8354 (N_8354,N_5646,N_3896);
or U8355 (N_8355,N_5367,N_5055);
and U8356 (N_8356,N_3633,N_3441);
or U8357 (N_8357,N_3499,N_4867);
nand U8358 (N_8358,N_4609,N_3503);
and U8359 (N_8359,N_5601,N_3214);
nand U8360 (N_8360,N_3643,N_3384);
nand U8361 (N_8361,N_3365,N_3613);
and U8362 (N_8362,N_3333,N_4665);
xor U8363 (N_8363,N_3393,N_4927);
and U8364 (N_8364,N_4357,N_4606);
or U8365 (N_8365,N_5047,N_3570);
and U8366 (N_8366,N_5556,N_4274);
nand U8367 (N_8367,N_4524,N_5672);
and U8368 (N_8368,N_5183,N_3893);
and U8369 (N_8369,N_3744,N_4232);
or U8370 (N_8370,N_3170,N_3819);
xor U8371 (N_8371,N_5742,N_4864);
xor U8372 (N_8372,N_3402,N_5177);
and U8373 (N_8373,N_5324,N_4312);
nor U8374 (N_8374,N_4624,N_4405);
xnor U8375 (N_8375,N_6149,N_5520);
nor U8376 (N_8376,N_6234,N_6048);
xor U8377 (N_8377,N_4335,N_3188);
nand U8378 (N_8378,N_5666,N_4544);
and U8379 (N_8379,N_5249,N_3920);
and U8380 (N_8380,N_4944,N_3572);
and U8381 (N_8381,N_4312,N_5477);
xnor U8382 (N_8382,N_3888,N_4058);
nor U8383 (N_8383,N_5026,N_3496);
nor U8384 (N_8384,N_3204,N_5068);
and U8385 (N_8385,N_4360,N_5839);
or U8386 (N_8386,N_6106,N_3753);
xor U8387 (N_8387,N_4586,N_4280);
nor U8388 (N_8388,N_3517,N_6137);
and U8389 (N_8389,N_6116,N_3949);
and U8390 (N_8390,N_5215,N_4326);
nand U8391 (N_8391,N_5688,N_4870);
or U8392 (N_8392,N_4365,N_5126);
nor U8393 (N_8393,N_4117,N_5371);
xnor U8394 (N_8394,N_5296,N_3217);
nand U8395 (N_8395,N_5011,N_3448);
and U8396 (N_8396,N_5859,N_3786);
nor U8397 (N_8397,N_5291,N_5461);
and U8398 (N_8398,N_6186,N_5822);
or U8399 (N_8399,N_5064,N_5644);
nand U8400 (N_8400,N_3876,N_5589);
nor U8401 (N_8401,N_5718,N_3958);
nor U8402 (N_8402,N_5224,N_3743);
nor U8403 (N_8403,N_5698,N_6092);
xor U8404 (N_8404,N_3793,N_4472);
xor U8405 (N_8405,N_5576,N_5560);
nand U8406 (N_8406,N_4658,N_6194);
nor U8407 (N_8407,N_5574,N_3835);
and U8408 (N_8408,N_6126,N_3151);
xnor U8409 (N_8409,N_3745,N_5803);
or U8410 (N_8410,N_5348,N_4405);
or U8411 (N_8411,N_4460,N_3353);
xnor U8412 (N_8412,N_4292,N_4745);
nor U8413 (N_8413,N_3291,N_3491);
and U8414 (N_8414,N_5202,N_3549);
and U8415 (N_8415,N_4586,N_4554);
nand U8416 (N_8416,N_5035,N_5274);
or U8417 (N_8417,N_4123,N_5290);
xor U8418 (N_8418,N_5340,N_4558);
nor U8419 (N_8419,N_5829,N_3815);
nand U8420 (N_8420,N_3943,N_4291);
or U8421 (N_8421,N_3955,N_4128);
or U8422 (N_8422,N_5358,N_6023);
nor U8423 (N_8423,N_4100,N_5951);
nand U8424 (N_8424,N_4605,N_5896);
nor U8425 (N_8425,N_5232,N_4418);
xor U8426 (N_8426,N_5339,N_3328);
nand U8427 (N_8427,N_5185,N_5258);
or U8428 (N_8428,N_4585,N_5728);
xnor U8429 (N_8429,N_4088,N_4238);
nand U8430 (N_8430,N_5081,N_4426);
and U8431 (N_8431,N_4116,N_3208);
nor U8432 (N_8432,N_5915,N_3409);
and U8433 (N_8433,N_5566,N_5214);
or U8434 (N_8434,N_6227,N_4084);
or U8435 (N_8435,N_4570,N_4005);
or U8436 (N_8436,N_6101,N_4596);
nand U8437 (N_8437,N_3553,N_3875);
nand U8438 (N_8438,N_5541,N_4454);
xor U8439 (N_8439,N_3420,N_5142);
and U8440 (N_8440,N_5199,N_3236);
nor U8441 (N_8441,N_3146,N_6047);
nor U8442 (N_8442,N_3863,N_5534);
nor U8443 (N_8443,N_4984,N_4110);
or U8444 (N_8444,N_3865,N_3524);
xnor U8445 (N_8445,N_5065,N_5009);
xnor U8446 (N_8446,N_3242,N_4969);
nor U8447 (N_8447,N_5516,N_5943);
or U8448 (N_8448,N_5206,N_3989);
nand U8449 (N_8449,N_3480,N_4041);
xor U8450 (N_8450,N_5139,N_3975);
nand U8451 (N_8451,N_3587,N_5179);
and U8452 (N_8452,N_3298,N_5705);
nand U8453 (N_8453,N_4388,N_5583);
or U8454 (N_8454,N_4013,N_5278);
nand U8455 (N_8455,N_3801,N_6015);
and U8456 (N_8456,N_3577,N_4370);
and U8457 (N_8457,N_4044,N_5709);
nand U8458 (N_8458,N_5412,N_3780);
or U8459 (N_8459,N_5979,N_4924);
xnor U8460 (N_8460,N_5141,N_4653);
xor U8461 (N_8461,N_5774,N_3189);
nand U8462 (N_8462,N_4279,N_4139);
and U8463 (N_8463,N_3127,N_5913);
xnor U8464 (N_8464,N_3335,N_5276);
or U8465 (N_8465,N_5394,N_3614);
or U8466 (N_8466,N_4750,N_4818);
nor U8467 (N_8467,N_5701,N_5548);
nor U8468 (N_8468,N_6031,N_3207);
and U8469 (N_8469,N_5146,N_3929);
or U8470 (N_8470,N_4977,N_5601);
or U8471 (N_8471,N_5437,N_6111);
and U8472 (N_8472,N_6040,N_4987);
nor U8473 (N_8473,N_4281,N_3656);
xor U8474 (N_8474,N_4398,N_5153);
nor U8475 (N_8475,N_4121,N_5338);
nand U8476 (N_8476,N_4166,N_5077);
nand U8477 (N_8477,N_5111,N_4832);
xnor U8478 (N_8478,N_5317,N_5527);
and U8479 (N_8479,N_5791,N_4583);
nor U8480 (N_8480,N_4136,N_4549);
nand U8481 (N_8481,N_5985,N_4136);
xor U8482 (N_8482,N_5916,N_4034);
and U8483 (N_8483,N_3980,N_3807);
and U8484 (N_8484,N_3375,N_4030);
or U8485 (N_8485,N_3744,N_3253);
or U8486 (N_8486,N_3684,N_5024);
or U8487 (N_8487,N_3405,N_5530);
and U8488 (N_8488,N_6210,N_5987);
nand U8489 (N_8489,N_5260,N_3848);
and U8490 (N_8490,N_3520,N_4847);
nor U8491 (N_8491,N_4615,N_3946);
nor U8492 (N_8492,N_3213,N_4257);
nor U8493 (N_8493,N_4857,N_4127);
nand U8494 (N_8494,N_3445,N_5076);
or U8495 (N_8495,N_3503,N_4076);
and U8496 (N_8496,N_5028,N_5962);
or U8497 (N_8497,N_5379,N_4741);
nand U8498 (N_8498,N_4296,N_4580);
xnor U8499 (N_8499,N_3530,N_5661);
or U8500 (N_8500,N_4458,N_3989);
and U8501 (N_8501,N_3962,N_3939);
nor U8502 (N_8502,N_5408,N_5445);
or U8503 (N_8503,N_6174,N_5397);
or U8504 (N_8504,N_4149,N_4825);
nand U8505 (N_8505,N_4317,N_5686);
xor U8506 (N_8506,N_5824,N_4563);
nor U8507 (N_8507,N_3294,N_4499);
and U8508 (N_8508,N_4282,N_5909);
nand U8509 (N_8509,N_4090,N_3497);
nand U8510 (N_8510,N_5944,N_3584);
xnor U8511 (N_8511,N_4874,N_5597);
or U8512 (N_8512,N_6035,N_3619);
and U8513 (N_8513,N_6073,N_5518);
nor U8514 (N_8514,N_4935,N_3823);
nand U8515 (N_8515,N_6100,N_5851);
and U8516 (N_8516,N_4726,N_5339);
nand U8517 (N_8517,N_3184,N_6169);
xor U8518 (N_8518,N_5898,N_4727);
nand U8519 (N_8519,N_5277,N_4228);
and U8520 (N_8520,N_3320,N_6085);
xor U8521 (N_8521,N_5340,N_3344);
and U8522 (N_8522,N_3950,N_4010);
xnor U8523 (N_8523,N_5593,N_6179);
nor U8524 (N_8524,N_3772,N_5568);
nand U8525 (N_8525,N_6043,N_3664);
nor U8526 (N_8526,N_4163,N_4263);
nand U8527 (N_8527,N_4900,N_5776);
and U8528 (N_8528,N_6003,N_3325);
xor U8529 (N_8529,N_4865,N_3870);
or U8530 (N_8530,N_3361,N_4583);
or U8531 (N_8531,N_5721,N_4860);
nand U8532 (N_8532,N_6213,N_6085);
xor U8533 (N_8533,N_4026,N_5571);
and U8534 (N_8534,N_5292,N_6046);
xnor U8535 (N_8535,N_4641,N_5688);
or U8536 (N_8536,N_6224,N_3648);
nor U8537 (N_8537,N_5366,N_5153);
nand U8538 (N_8538,N_5880,N_5794);
nor U8539 (N_8539,N_3413,N_3619);
nand U8540 (N_8540,N_5543,N_6059);
and U8541 (N_8541,N_3228,N_4813);
nand U8542 (N_8542,N_4440,N_3572);
nand U8543 (N_8543,N_3921,N_4412);
and U8544 (N_8544,N_3450,N_3500);
nand U8545 (N_8545,N_5759,N_5998);
xnor U8546 (N_8546,N_5330,N_3783);
nand U8547 (N_8547,N_4311,N_5264);
xnor U8548 (N_8548,N_5881,N_6099);
nor U8549 (N_8549,N_6222,N_5348);
or U8550 (N_8550,N_6032,N_5544);
and U8551 (N_8551,N_3624,N_3873);
nand U8552 (N_8552,N_5004,N_5114);
or U8553 (N_8553,N_5356,N_6132);
xnor U8554 (N_8554,N_3376,N_3450);
or U8555 (N_8555,N_6103,N_5700);
nand U8556 (N_8556,N_4062,N_5991);
nor U8557 (N_8557,N_6096,N_5569);
or U8558 (N_8558,N_5236,N_5971);
xor U8559 (N_8559,N_3772,N_3348);
and U8560 (N_8560,N_3968,N_4973);
or U8561 (N_8561,N_5928,N_5937);
nand U8562 (N_8562,N_3461,N_4973);
nor U8563 (N_8563,N_6143,N_4392);
nor U8564 (N_8564,N_3943,N_5233);
nand U8565 (N_8565,N_5798,N_6023);
or U8566 (N_8566,N_5290,N_3295);
and U8567 (N_8567,N_5602,N_4391);
xnor U8568 (N_8568,N_5168,N_4946);
and U8569 (N_8569,N_5485,N_4796);
and U8570 (N_8570,N_3502,N_4489);
or U8571 (N_8571,N_3604,N_3140);
xor U8572 (N_8572,N_5337,N_3487);
and U8573 (N_8573,N_4465,N_5342);
nand U8574 (N_8574,N_3689,N_6103);
nor U8575 (N_8575,N_6204,N_5961);
nor U8576 (N_8576,N_3693,N_5213);
or U8577 (N_8577,N_5653,N_3955);
nor U8578 (N_8578,N_6094,N_3566);
and U8579 (N_8579,N_3347,N_4582);
xor U8580 (N_8580,N_4800,N_5860);
nand U8581 (N_8581,N_4741,N_6112);
xnor U8582 (N_8582,N_6247,N_3870);
nand U8583 (N_8583,N_5012,N_3653);
and U8584 (N_8584,N_3882,N_5817);
xnor U8585 (N_8585,N_3257,N_3961);
nand U8586 (N_8586,N_4492,N_5136);
nand U8587 (N_8587,N_6124,N_5844);
and U8588 (N_8588,N_5219,N_6170);
xor U8589 (N_8589,N_3783,N_3648);
and U8590 (N_8590,N_5829,N_5661);
nand U8591 (N_8591,N_3804,N_5674);
xnor U8592 (N_8592,N_3356,N_5378);
nand U8593 (N_8593,N_4394,N_3484);
and U8594 (N_8594,N_6144,N_3510);
nor U8595 (N_8595,N_5754,N_5675);
and U8596 (N_8596,N_4369,N_4966);
nor U8597 (N_8597,N_4079,N_4758);
and U8598 (N_8598,N_3295,N_3892);
nor U8599 (N_8599,N_4589,N_4586);
nand U8600 (N_8600,N_5480,N_3570);
nand U8601 (N_8601,N_4793,N_5121);
and U8602 (N_8602,N_5304,N_4777);
nand U8603 (N_8603,N_3641,N_5875);
nand U8604 (N_8604,N_4190,N_4699);
xnor U8605 (N_8605,N_3609,N_4977);
nor U8606 (N_8606,N_4297,N_4678);
xnor U8607 (N_8607,N_5435,N_4093);
and U8608 (N_8608,N_5963,N_5783);
nor U8609 (N_8609,N_3824,N_4135);
or U8610 (N_8610,N_5129,N_3888);
and U8611 (N_8611,N_5562,N_6176);
or U8612 (N_8612,N_4173,N_5380);
xnor U8613 (N_8613,N_4317,N_5847);
nor U8614 (N_8614,N_4313,N_4275);
nor U8615 (N_8615,N_4261,N_3919);
nand U8616 (N_8616,N_5524,N_4610);
nand U8617 (N_8617,N_4619,N_4948);
or U8618 (N_8618,N_3724,N_4225);
xnor U8619 (N_8619,N_4276,N_5496);
and U8620 (N_8620,N_4841,N_4983);
or U8621 (N_8621,N_5004,N_5918);
nand U8622 (N_8622,N_5647,N_4894);
nor U8623 (N_8623,N_5983,N_4862);
nand U8624 (N_8624,N_4637,N_3894);
nor U8625 (N_8625,N_3324,N_3262);
or U8626 (N_8626,N_3547,N_4286);
and U8627 (N_8627,N_5583,N_5671);
nand U8628 (N_8628,N_4739,N_5355);
and U8629 (N_8629,N_3550,N_5520);
nand U8630 (N_8630,N_5125,N_3888);
xor U8631 (N_8631,N_4910,N_4495);
xnor U8632 (N_8632,N_5320,N_3536);
nor U8633 (N_8633,N_4701,N_5444);
and U8634 (N_8634,N_4502,N_4409);
nand U8635 (N_8635,N_5352,N_4793);
xor U8636 (N_8636,N_5139,N_6174);
xor U8637 (N_8637,N_3523,N_5176);
nor U8638 (N_8638,N_4113,N_4099);
and U8639 (N_8639,N_3232,N_5528);
nor U8640 (N_8640,N_5906,N_4529);
nand U8641 (N_8641,N_4695,N_5919);
nor U8642 (N_8642,N_3748,N_5587);
or U8643 (N_8643,N_3833,N_4530);
and U8644 (N_8644,N_4898,N_3774);
xnor U8645 (N_8645,N_4300,N_3197);
or U8646 (N_8646,N_3502,N_3539);
and U8647 (N_8647,N_5182,N_4933);
and U8648 (N_8648,N_5374,N_4873);
or U8649 (N_8649,N_5314,N_4377);
or U8650 (N_8650,N_3228,N_6209);
and U8651 (N_8651,N_5933,N_5388);
nand U8652 (N_8652,N_4067,N_4111);
or U8653 (N_8653,N_4810,N_5939);
nor U8654 (N_8654,N_3998,N_5415);
or U8655 (N_8655,N_4040,N_5558);
and U8656 (N_8656,N_3616,N_4910);
and U8657 (N_8657,N_4558,N_3445);
or U8658 (N_8658,N_5598,N_4968);
and U8659 (N_8659,N_5259,N_3713);
and U8660 (N_8660,N_5873,N_5318);
and U8661 (N_8661,N_3518,N_3487);
or U8662 (N_8662,N_3917,N_5554);
xnor U8663 (N_8663,N_4728,N_3462);
or U8664 (N_8664,N_5176,N_5439);
and U8665 (N_8665,N_4621,N_3295);
nand U8666 (N_8666,N_3442,N_6106);
or U8667 (N_8667,N_4357,N_4809);
xor U8668 (N_8668,N_5471,N_4488);
nor U8669 (N_8669,N_5343,N_3278);
and U8670 (N_8670,N_5533,N_3247);
or U8671 (N_8671,N_4351,N_5692);
nor U8672 (N_8672,N_5871,N_3175);
and U8673 (N_8673,N_3184,N_4930);
and U8674 (N_8674,N_3966,N_3294);
nand U8675 (N_8675,N_5372,N_4748);
or U8676 (N_8676,N_5508,N_5685);
nand U8677 (N_8677,N_4736,N_4165);
nand U8678 (N_8678,N_4155,N_3335);
and U8679 (N_8679,N_3133,N_4058);
xnor U8680 (N_8680,N_5802,N_3837);
xor U8681 (N_8681,N_4752,N_4968);
nor U8682 (N_8682,N_5384,N_5568);
xnor U8683 (N_8683,N_3827,N_3880);
or U8684 (N_8684,N_4067,N_3524);
nor U8685 (N_8685,N_4249,N_4606);
nand U8686 (N_8686,N_3772,N_3360);
and U8687 (N_8687,N_6148,N_3910);
nand U8688 (N_8688,N_4366,N_4145);
or U8689 (N_8689,N_5707,N_4209);
or U8690 (N_8690,N_5042,N_3595);
and U8691 (N_8691,N_5707,N_6022);
nor U8692 (N_8692,N_4895,N_3858);
or U8693 (N_8693,N_3273,N_5462);
nand U8694 (N_8694,N_4691,N_3958);
nor U8695 (N_8695,N_3705,N_3795);
nor U8696 (N_8696,N_3689,N_5202);
xnor U8697 (N_8697,N_3813,N_3561);
and U8698 (N_8698,N_5797,N_5431);
nand U8699 (N_8699,N_5302,N_4881);
and U8700 (N_8700,N_4548,N_5222);
and U8701 (N_8701,N_4431,N_3902);
nand U8702 (N_8702,N_4354,N_5151);
nand U8703 (N_8703,N_5198,N_5170);
xor U8704 (N_8704,N_6200,N_4799);
and U8705 (N_8705,N_4999,N_3401);
nor U8706 (N_8706,N_3386,N_3702);
nor U8707 (N_8707,N_4341,N_4948);
nand U8708 (N_8708,N_4966,N_4327);
xor U8709 (N_8709,N_3961,N_3288);
xor U8710 (N_8710,N_3927,N_3246);
xor U8711 (N_8711,N_5921,N_4191);
nand U8712 (N_8712,N_4979,N_4213);
xor U8713 (N_8713,N_5628,N_5509);
nor U8714 (N_8714,N_4945,N_5298);
or U8715 (N_8715,N_3877,N_4136);
nand U8716 (N_8716,N_4126,N_5315);
xnor U8717 (N_8717,N_5590,N_3264);
or U8718 (N_8718,N_4309,N_5776);
or U8719 (N_8719,N_5355,N_3737);
or U8720 (N_8720,N_3225,N_4942);
and U8721 (N_8721,N_4100,N_5696);
and U8722 (N_8722,N_5021,N_5104);
or U8723 (N_8723,N_6119,N_4371);
nor U8724 (N_8724,N_6234,N_3568);
or U8725 (N_8725,N_5343,N_4776);
or U8726 (N_8726,N_3641,N_4064);
xnor U8727 (N_8727,N_6125,N_3282);
xnor U8728 (N_8728,N_5355,N_5785);
or U8729 (N_8729,N_5912,N_5058);
or U8730 (N_8730,N_5754,N_6140);
and U8731 (N_8731,N_4686,N_5997);
and U8732 (N_8732,N_5952,N_4536);
or U8733 (N_8733,N_5028,N_3468);
xnor U8734 (N_8734,N_5816,N_3137);
xor U8735 (N_8735,N_3153,N_4398);
and U8736 (N_8736,N_5862,N_5322);
nor U8737 (N_8737,N_6035,N_4306);
nand U8738 (N_8738,N_3700,N_5439);
nand U8739 (N_8739,N_4363,N_4615);
and U8740 (N_8740,N_6142,N_5820);
nor U8741 (N_8741,N_4643,N_5627);
and U8742 (N_8742,N_5917,N_5997);
and U8743 (N_8743,N_5414,N_4792);
nor U8744 (N_8744,N_5447,N_5431);
nand U8745 (N_8745,N_5456,N_3848);
nor U8746 (N_8746,N_3524,N_4332);
nor U8747 (N_8747,N_5279,N_6006);
nand U8748 (N_8748,N_5574,N_4002);
nand U8749 (N_8749,N_3661,N_3448);
nor U8750 (N_8750,N_5975,N_3746);
xor U8751 (N_8751,N_4078,N_4008);
nor U8752 (N_8752,N_5264,N_5903);
or U8753 (N_8753,N_4383,N_4759);
xnor U8754 (N_8754,N_5656,N_3622);
xor U8755 (N_8755,N_3404,N_4571);
xnor U8756 (N_8756,N_3738,N_5647);
or U8757 (N_8757,N_3617,N_5447);
nand U8758 (N_8758,N_4675,N_5436);
xnor U8759 (N_8759,N_3368,N_6240);
nor U8760 (N_8760,N_5840,N_4984);
xor U8761 (N_8761,N_4326,N_4245);
or U8762 (N_8762,N_4548,N_4802);
nor U8763 (N_8763,N_3641,N_5030);
and U8764 (N_8764,N_3884,N_5736);
xnor U8765 (N_8765,N_6223,N_4447);
xor U8766 (N_8766,N_3545,N_5113);
nand U8767 (N_8767,N_4029,N_5050);
nor U8768 (N_8768,N_3951,N_3931);
nand U8769 (N_8769,N_5466,N_4192);
xor U8770 (N_8770,N_3600,N_5739);
nand U8771 (N_8771,N_4713,N_3723);
nand U8772 (N_8772,N_5769,N_6044);
nand U8773 (N_8773,N_4427,N_5696);
and U8774 (N_8774,N_5016,N_5191);
xor U8775 (N_8775,N_4594,N_4578);
nand U8776 (N_8776,N_6124,N_5307);
or U8777 (N_8777,N_5705,N_5790);
and U8778 (N_8778,N_6077,N_5965);
nor U8779 (N_8779,N_4957,N_6069);
nor U8780 (N_8780,N_5621,N_5574);
and U8781 (N_8781,N_3531,N_5942);
and U8782 (N_8782,N_4087,N_3155);
xor U8783 (N_8783,N_6129,N_5584);
nor U8784 (N_8784,N_3307,N_5347);
and U8785 (N_8785,N_3564,N_4685);
xnor U8786 (N_8786,N_4148,N_4633);
nand U8787 (N_8787,N_6056,N_6219);
nor U8788 (N_8788,N_5739,N_3462);
xor U8789 (N_8789,N_4073,N_3974);
xnor U8790 (N_8790,N_3840,N_5757);
xnor U8791 (N_8791,N_5715,N_5814);
nor U8792 (N_8792,N_3902,N_5905);
nor U8793 (N_8793,N_3367,N_5375);
and U8794 (N_8794,N_5840,N_3644);
or U8795 (N_8795,N_5024,N_4965);
nor U8796 (N_8796,N_3147,N_5368);
nand U8797 (N_8797,N_5340,N_4958);
nor U8798 (N_8798,N_5549,N_4783);
nor U8799 (N_8799,N_3734,N_5112);
or U8800 (N_8800,N_4577,N_4311);
xor U8801 (N_8801,N_3232,N_5754);
and U8802 (N_8802,N_4875,N_5241);
nand U8803 (N_8803,N_6166,N_4721);
xor U8804 (N_8804,N_6196,N_3906);
or U8805 (N_8805,N_3478,N_3189);
nor U8806 (N_8806,N_5174,N_5129);
xnor U8807 (N_8807,N_5588,N_3802);
and U8808 (N_8808,N_3178,N_3541);
nand U8809 (N_8809,N_3302,N_5931);
or U8810 (N_8810,N_5973,N_3784);
xor U8811 (N_8811,N_5696,N_5074);
or U8812 (N_8812,N_6133,N_5265);
and U8813 (N_8813,N_3538,N_3301);
xor U8814 (N_8814,N_6207,N_4318);
nor U8815 (N_8815,N_4675,N_5927);
nand U8816 (N_8816,N_4238,N_3708);
xor U8817 (N_8817,N_3984,N_4658);
xor U8818 (N_8818,N_4448,N_5523);
nand U8819 (N_8819,N_5829,N_5651);
or U8820 (N_8820,N_3699,N_4647);
or U8821 (N_8821,N_6010,N_5369);
nand U8822 (N_8822,N_4081,N_4170);
or U8823 (N_8823,N_4987,N_5188);
nand U8824 (N_8824,N_5315,N_4170);
or U8825 (N_8825,N_4426,N_5949);
and U8826 (N_8826,N_4833,N_5218);
or U8827 (N_8827,N_4454,N_3726);
nor U8828 (N_8828,N_4118,N_6164);
nand U8829 (N_8829,N_3442,N_6145);
xor U8830 (N_8830,N_3561,N_5437);
xor U8831 (N_8831,N_6042,N_3909);
nor U8832 (N_8832,N_4248,N_3925);
or U8833 (N_8833,N_4274,N_5349);
nor U8834 (N_8834,N_5672,N_5289);
and U8835 (N_8835,N_3662,N_5919);
xor U8836 (N_8836,N_5900,N_3785);
and U8837 (N_8837,N_3985,N_5817);
and U8838 (N_8838,N_5198,N_5260);
xor U8839 (N_8839,N_5924,N_5531);
nor U8840 (N_8840,N_4620,N_3869);
nor U8841 (N_8841,N_5407,N_5680);
xnor U8842 (N_8842,N_4128,N_3144);
and U8843 (N_8843,N_4063,N_5572);
nand U8844 (N_8844,N_5534,N_6188);
and U8845 (N_8845,N_6225,N_3901);
and U8846 (N_8846,N_3380,N_3790);
nand U8847 (N_8847,N_3636,N_3393);
nor U8848 (N_8848,N_5614,N_4134);
and U8849 (N_8849,N_5006,N_5529);
nor U8850 (N_8850,N_5856,N_3275);
nor U8851 (N_8851,N_5703,N_4359);
xnor U8852 (N_8852,N_5156,N_5041);
and U8853 (N_8853,N_4398,N_6220);
nor U8854 (N_8854,N_4878,N_3215);
nand U8855 (N_8855,N_3601,N_5662);
and U8856 (N_8856,N_6135,N_3493);
and U8857 (N_8857,N_6119,N_4638);
nand U8858 (N_8858,N_5129,N_3843);
nand U8859 (N_8859,N_4398,N_3451);
nand U8860 (N_8860,N_4770,N_3295);
xnor U8861 (N_8861,N_4486,N_4044);
nand U8862 (N_8862,N_3918,N_5975);
xor U8863 (N_8863,N_5686,N_4572);
nand U8864 (N_8864,N_5966,N_5364);
xnor U8865 (N_8865,N_5227,N_5521);
nor U8866 (N_8866,N_5960,N_4130);
xor U8867 (N_8867,N_5664,N_3322);
nand U8868 (N_8868,N_6162,N_5709);
nand U8869 (N_8869,N_4395,N_4386);
and U8870 (N_8870,N_3448,N_4673);
nand U8871 (N_8871,N_4356,N_3211);
xor U8872 (N_8872,N_3128,N_6120);
nor U8873 (N_8873,N_5912,N_4530);
and U8874 (N_8874,N_4019,N_3932);
xnor U8875 (N_8875,N_4156,N_4268);
or U8876 (N_8876,N_4330,N_5119);
and U8877 (N_8877,N_3450,N_6240);
or U8878 (N_8878,N_5697,N_3735);
xnor U8879 (N_8879,N_6152,N_4844);
and U8880 (N_8880,N_4761,N_4981);
and U8881 (N_8881,N_3832,N_3478);
nor U8882 (N_8882,N_3807,N_3651);
xnor U8883 (N_8883,N_5563,N_3844);
nand U8884 (N_8884,N_3426,N_5481);
nor U8885 (N_8885,N_6012,N_3943);
xnor U8886 (N_8886,N_6197,N_3217);
or U8887 (N_8887,N_3885,N_5677);
xor U8888 (N_8888,N_5204,N_3494);
or U8889 (N_8889,N_5070,N_4986);
nor U8890 (N_8890,N_4311,N_3910);
and U8891 (N_8891,N_5113,N_4032);
nand U8892 (N_8892,N_3621,N_5887);
nor U8893 (N_8893,N_3193,N_5491);
and U8894 (N_8894,N_4581,N_4609);
xnor U8895 (N_8895,N_5685,N_3920);
xor U8896 (N_8896,N_4401,N_5844);
xnor U8897 (N_8897,N_4189,N_4778);
xnor U8898 (N_8898,N_3309,N_5497);
xnor U8899 (N_8899,N_3935,N_4181);
nor U8900 (N_8900,N_6213,N_5792);
nand U8901 (N_8901,N_3602,N_5935);
xor U8902 (N_8902,N_5919,N_5420);
nor U8903 (N_8903,N_4831,N_4152);
and U8904 (N_8904,N_4130,N_3370);
or U8905 (N_8905,N_5083,N_6064);
or U8906 (N_8906,N_3347,N_3577);
or U8907 (N_8907,N_4529,N_3525);
or U8908 (N_8908,N_3145,N_4007);
xnor U8909 (N_8909,N_4080,N_4045);
nor U8910 (N_8910,N_4825,N_4273);
nor U8911 (N_8911,N_5020,N_4840);
nand U8912 (N_8912,N_4376,N_4379);
nand U8913 (N_8913,N_4684,N_4768);
nor U8914 (N_8914,N_6037,N_5414);
xor U8915 (N_8915,N_4938,N_3801);
or U8916 (N_8916,N_4283,N_4377);
nand U8917 (N_8917,N_4165,N_5883);
nand U8918 (N_8918,N_5243,N_4869);
nand U8919 (N_8919,N_3868,N_5890);
and U8920 (N_8920,N_5323,N_4518);
and U8921 (N_8921,N_5746,N_3275);
and U8922 (N_8922,N_3601,N_3466);
or U8923 (N_8923,N_5058,N_4102);
and U8924 (N_8924,N_4045,N_6244);
or U8925 (N_8925,N_4067,N_4798);
or U8926 (N_8926,N_3846,N_4652);
and U8927 (N_8927,N_3785,N_4219);
and U8928 (N_8928,N_4708,N_5663);
xor U8929 (N_8929,N_3563,N_3285);
xnor U8930 (N_8930,N_5432,N_5729);
nor U8931 (N_8931,N_5091,N_4877);
or U8932 (N_8932,N_5133,N_5950);
nand U8933 (N_8933,N_4666,N_3758);
and U8934 (N_8934,N_5978,N_5713);
nor U8935 (N_8935,N_6118,N_5984);
nor U8936 (N_8936,N_4134,N_3516);
or U8937 (N_8937,N_3929,N_3258);
nand U8938 (N_8938,N_3637,N_3752);
nand U8939 (N_8939,N_5687,N_3996);
nor U8940 (N_8940,N_4431,N_4012);
nand U8941 (N_8941,N_5804,N_4067);
xor U8942 (N_8942,N_4014,N_4047);
xnor U8943 (N_8943,N_4965,N_4692);
or U8944 (N_8944,N_3978,N_5535);
xor U8945 (N_8945,N_3742,N_3469);
xnor U8946 (N_8946,N_3671,N_4372);
or U8947 (N_8947,N_6086,N_3373);
nand U8948 (N_8948,N_6212,N_4704);
and U8949 (N_8949,N_3681,N_3452);
xor U8950 (N_8950,N_3767,N_4867);
nor U8951 (N_8951,N_3985,N_3968);
nand U8952 (N_8952,N_3537,N_3756);
nor U8953 (N_8953,N_4020,N_6012);
or U8954 (N_8954,N_5772,N_5723);
nor U8955 (N_8955,N_5513,N_4680);
nand U8956 (N_8956,N_5125,N_3395);
and U8957 (N_8957,N_4628,N_3695);
nor U8958 (N_8958,N_5772,N_3731);
xor U8959 (N_8959,N_6238,N_3537);
nor U8960 (N_8960,N_5127,N_5022);
nor U8961 (N_8961,N_4890,N_4531);
and U8962 (N_8962,N_3924,N_4987);
xor U8963 (N_8963,N_5057,N_5145);
xnor U8964 (N_8964,N_4350,N_6157);
and U8965 (N_8965,N_4353,N_5862);
nor U8966 (N_8966,N_5242,N_4027);
and U8967 (N_8967,N_3372,N_4133);
or U8968 (N_8968,N_4450,N_4411);
xnor U8969 (N_8969,N_3536,N_3293);
xor U8970 (N_8970,N_3268,N_3562);
nor U8971 (N_8971,N_4289,N_4347);
xor U8972 (N_8972,N_5028,N_5557);
nor U8973 (N_8973,N_3531,N_3525);
or U8974 (N_8974,N_3635,N_5112);
nand U8975 (N_8975,N_4956,N_3757);
nand U8976 (N_8976,N_4950,N_3366);
and U8977 (N_8977,N_3629,N_3748);
or U8978 (N_8978,N_4811,N_4419);
xnor U8979 (N_8979,N_6132,N_3192);
and U8980 (N_8980,N_3647,N_3465);
nand U8981 (N_8981,N_4736,N_4742);
nand U8982 (N_8982,N_4088,N_4586);
and U8983 (N_8983,N_6153,N_4234);
xnor U8984 (N_8984,N_4529,N_3582);
and U8985 (N_8985,N_5548,N_3397);
xor U8986 (N_8986,N_5960,N_5124);
xor U8987 (N_8987,N_6015,N_5346);
xor U8988 (N_8988,N_5832,N_4610);
xor U8989 (N_8989,N_4251,N_4724);
or U8990 (N_8990,N_4943,N_4814);
or U8991 (N_8991,N_3149,N_4963);
or U8992 (N_8992,N_4460,N_6166);
or U8993 (N_8993,N_4217,N_6076);
and U8994 (N_8994,N_4073,N_6084);
and U8995 (N_8995,N_5188,N_3128);
and U8996 (N_8996,N_3807,N_5304);
xnor U8997 (N_8997,N_3503,N_4128);
xnor U8998 (N_8998,N_4730,N_4183);
nor U8999 (N_8999,N_6020,N_5737);
nand U9000 (N_9000,N_4330,N_4610);
or U9001 (N_9001,N_4787,N_4801);
xor U9002 (N_9002,N_5929,N_3905);
nor U9003 (N_9003,N_4456,N_5113);
and U9004 (N_9004,N_4491,N_4519);
nor U9005 (N_9005,N_4229,N_4135);
xor U9006 (N_9006,N_5011,N_3634);
and U9007 (N_9007,N_5260,N_3307);
nand U9008 (N_9008,N_5745,N_6163);
xor U9009 (N_9009,N_4062,N_4776);
xor U9010 (N_9010,N_3938,N_3639);
xor U9011 (N_9011,N_5381,N_5107);
nor U9012 (N_9012,N_5755,N_3558);
nand U9013 (N_9013,N_5264,N_5072);
xor U9014 (N_9014,N_5328,N_5886);
nor U9015 (N_9015,N_5459,N_3427);
nor U9016 (N_9016,N_4628,N_5629);
nand U9017 (N_9017,N_4482,N_3133);
nand U9018 (N_9018,N_3799,N_4403);
and U9019 (N_9019,N_3973,N_5700);
and U9020 (N_9020,N_4562,N_3493);
or U9021 (N_9021,N_4064,N_4855);
or U9022 (N_9022,N_3528,N_4268);
xor U9023 (N_9023,N_4051,N_3746);
nand U9024 (N_9024,N_5560,N_3872);
xor U9025 (N_9025,N_3311,N_5879);
nand U9026 (N_9026,N_4226,N_4913);
nor U9027 (N_9027,N_3243,N_5819);
nor U9028 (N_9028,N_4256,N_5603);
or U9029 (N_9029,N_3411,N_5440);
and U9030 (N_9030,N_6009,N_4813);
nand U9031 (N_9031,N_5322,N_3697);
xnor U9032 (N_9032,N_4775,N_5249);
nor U9033 (N_9033,N_5781,N_3810);
nor U9034 (N_9034,N_3845,N_5636);
xor U9035 (N_9035,N_3627,N_3355);
nor U9036 (N_9036,N_6076,N_3891);
nor U9037 (N_9037,N_5542,N_4618);
and U9038 (N_9038,N_3225,N_3540);
nor U9039 (N_9039,N_3927,N_4265);
nor U9040 (N_9040,N_5155,N_5194);
xor U9041 (N_9041,N_4397,N_4165);
nor U9042 (N_9042,N_6097,N_5002);
and U9043 (N_9043,N_4641,N_3612);
nand U9044 (N_9044,N_5169,N_3126);
nor U9045 (N_9045,N_3380,N_6002);
xor U9046 (N_9046,N_5649,N_4008);
xnor U9047 (N_9047,N_5039,N_3803);
xor U9048 (N_9048,N_5899,N_6157);
nor U9049 (N_9049,N_5552,N_5848);
xnor U9050 (N_9050,N_5487,N_4379);
xnor U9051 (N_9051,N_4139,N_4025);
xor U9052 (N_9052,N_5077,N_3155);
and U9053 (N_9053,N_6070,N_3864);
xnor U9054 (N_9054,N_4494,N_5338);
xnor U9055 (N_9055,N_5101,N_4011);
xor U9056 (N_9056,N_6141,N_5105);
and U9057 (N_9057,N_4586,N_4344);
and U9058 (N_9058,N_5265,N_4996);
nor U9059 (N_9059,N_6122,N_6209);
nand U9060 (N_9060,N_5286,N_4542);
nor U9061 (N_9061,N_5537,N_5677);
and U9062 (N_9062,N_5783,N_5889);
nor U9063 (N_9063,N_5768,N_3621);
nand U9064 (N_9064,N_5546,N_3268);
or U9065 (N_9065,N_5104,N_3815);
xor U9066 (N_9066,N_4320,N_4673);
and U9067 (N_9067,N_5323,N_3796);
nor U9068 (N_9068,N_5358,N_3202);
xnor U9069 (N_9069,N_3596,N_3608);
or U9070 (N_9070,N_4389,N_6016);
nand U9071 (N_9071,N_6042,N_5646);
xnor U9072 (N_9072,N_4972,N_6246);
xor U9073 (N_9073,N_4806,N_5865);
nor U9074 (N_9074,N_3502,N_4499);
nor U9075 (N_9075,N_3476,N_6027);
nand U9076 (N_9076,N_3186,N_3172);
and U9077 (N_9077,N_4108,N_3148);
xnor U9078 (N_9078,N_4275,N_5127);
nand U9079 (N_9079,N_4053,N_3357);
or U9080 (N_9080,N_5852,N_4836);
nand U9081 (N_9081,N_5797,N_4174);
nor U9082 (N_9082,N_5327,N_6242);
nand U9083 (N_9083,N_4858,N_5146);
nor U9084 (N_9084,N_5098,N_4559);
nor U9085 (N_9085,N_3130,N_5961);
or U9086 (N_9086,N_3678,N_4511);
nand U9087 (N_9087,N_3304,N_4640);
xnor U9088 (N_9088,N_4917,N_4725);
and U9089 (N_9089,N_4146,N_3377);
xor U9090 (N_9090,N_3258,N_3319);
or U9091 (N_9091,N_5759,N_4755);
nor U9092 (N_9092,N_5978,N_3286);
nand U9093 (N_9093,N_5503,N_4697);
nand U9094 (N_9094,N_5661,N_5708);
and U9095 (N_9095,N_5015,N_4888);
nand U9096 (N_9096,N_6114,N_4998);
and U9097 (N_9097,N_3129,N_3438);
nor U9098 (N_9098,N_4221,N_3881);
nand U9099 (N_9099,N_5968,N_5889);
xor U9100 (N_9100,N_4531,N_4768);
xnor U9101 (N_9101,N_3264,N_4533);
xor U9102 (N_9102,N_5741,N_6088);
nand U9103 (N_9103,N_5090,N_4689);
or U9104 (N_9104,N_3442,N_5883);
nor U9105 (N_9105,N_6135,N_6241);
xnor U9106 (N_9106,N_4939,N_3288);
nor U9107 (N_9107,N_4512,N_5590);
or U9108 (N_9108,N_3205,N_3565);
and U9109 (N_9109,N_4692,N_3517);
and U9110 (N_9110,N_5019,N_3901);
and U9111 (N_9111,N_4006,N_4999);
xor U9112 (N_9112,N_5137,N_4786);
nand U9113 (N_9113,N_4613,N_5313);
nand U9114 (N_9114,N_4595,N_5209);
nor U9115 (N_9115,N_3144,N_4829);
nor U9116 (N_9116,N_5708,N_4091);
or U9117 (N_9117,N_6127,N_5176);
nand U9118 (N_9118,N_4465,N_3308);
and U9119 (N_9119,N_4626,N_3946);
or U9120 (N_9120,N_3186,N_6131);
and U9121 (N_9121,N_5796,N_3454);
or U9122 (N_9122,N_5076,N_3908);
xor U9123 (N_9123,N_4055,N_3335);
nand U9124 (N_9124,N_3757,N_5182);
or U9125 (N_9125,N_5203,N_4273);
xnor U9126 (N_9126,N_5296,N_4307);
nand U9127 (N_9127,N_5733,N_3755);
nand U9128 (N_9128,N_3354,N_4007);
nor U9129 (N_9129,N_5340,N_3860);
nand U9130 (N_9130,N_3462,N_4217);
nand U9131 (N_9131,N_3444,N_3352);
xnor U9132 (N_9132,N_4518,N_4945);
nor U9133 (N_9133,N_5353,N_3834);
xnor U9134 (N_9134,N_4092,N_3985);
nor U9135 (N_9135,N_5880,N_3421);
and U9136 (N_9136,N_3704,N_3364);
or U9137 (N_9137,N_6060,N_3386);
xnor U9138 (N_9138,N_3707,N_5247);
or U9139 (N_9139,N_3186,N_3899);
and U9140 (N_9140,N_3791,N_4514);
or U9141 (N_9141,N_4043,N_5266);
and U9142 (N_9142,N_4297,N_4196);
or U9143 (N_9143,N_5851,N_5795);
and U9144 (N_9144,N_4476,N_6153);
and U9145 (N_9145,N_3437,N_5783);
nand U9146 (N_9146,N_5404,N_5384);
or U9147 (N_9147,N_5672,N_3519);
nand U9148 (N_9148,N_6086,N_3800);
and U9149 (N_9149,N_3488,N_3806);
nand U9150 (N_9150,N_5382,N_3190);
nor U9151 (N_9151,N_4574,N_3944);
nor U9152 (N_9152,N_4222,N_4259);
nor U9153 (N_9153,N_6016,N_3531);
xnor U9154 (N_9154,N_4008,N_3568);
nand U9155 (N_9155,N_4462,N_5502);
or U9156 (N_9156,N_3252,N_3444);
nand U9157 (N_9157,N_6058,N_4368);
nor U9158 (N_9158,N_5281,N_5077);
and U9159 (N_9159,N_6023,N_5682);
nand U9160 (N_9160,N_5432,N_5439);
or U9161 (N_9161,N_5214,N_4475);
and U9162 (N_9162,N_3525,N_4795);
nand U9163 (N_9163,N_4869,N_3597);
and U9164 (N_9164,N_4585,N_3517);
and U9165 (N_9165,N_4430,N_5328);
and U9166 (N_9166,N_3667,N_4790);
nor U9167 (N_9167,N_4913,N_3625);
and U9168 (N_9168,N_3281,N_4413);
nor U9169 (N_9169,N_4833,N_5773);
or U9170 (N_9170,N_4158,N_3574);
xnor U9171 (N_9171,N_4703,N_3840);
and U9172 (N_9172,N_5556,N_3918);
nor U9173 (N_9173,N_5148,N_4677);
nand U9174 (N_9174,N_3934,N_5978);
and U9175 (N_9175,N_6249,N_4041);
nor U9176 (N_9176,N_4763,N_4507);
nand U9177 (N_9177,N_3804,N_4418);
and U9178 (N_9178,N_3350,N_5178);
nand U9179 (N_9179,N_3953,N_4808);
and U9180 (N_9180,N_4205,N_5307);
or U9181 (N_9181,N_5639,N_5264);
or U9182 (N_9182,N_3958,N_5238);
and U9183 (N_9183,N_3526,N_3202);
or U9184 (N_9184,N_6145,N_4787);
and U9185 (N_9185,N_4355,N_4778);
nor U9186 (N_9186,N_5846,N_4272);
and U9187 (N_9187,N_3508,N_3545);
and U9188 (N_9188,N_5142,N_3845);
xor U9189 (N_9189,N_3867,N_5437);
nand U9190 (N_9190,N_5639,N_4834);
or U9191 (N_9191,N_4128,N_5579);
xnor U9192 (N_9192,N_4412,N_5094);
or U9193 (N_9193,N_3139,N_5175);
xnor U9194 (N_9194,N_4147,N_5793);
and U9195 (N_9195,N_5556,N_3652);
nor U9196 (N_9196,N_3423,N_5020);
and U9197 (N_9197,N_5141,N_5340);
and U9198 (N_9198,N_6035,N_5927);
nand U9199 (N_9199,N_3926,N_5315);
nor U9200 (N_9200,N_3559,N_4264);
and U9201 (N_9201,N_4118,N_5990);
nor U9202 (N_9202,N_5752,N_4304);
and U9203 (N_9203,N_6026,N_3705);
or U9204 (N_9204,N_4841,N_5929);
and U9205 (N_9205,N_5941,N_5293);
nand U9206 (N_9206,N_5015,N_5941);
and U9207 (N_9207,N_3434,N_5148);
and U9208 (N_9208,N_5918,N_3990);
and U9209 (N_9209,N_3888,N_6187);
nand U9210 (N_9210,N_3661,N_4230);
nand U9211 (N_9211,N_5449,N_3846);
or U9212 (N_9212,N_5816,N_4244);
nor U9213 (N_9213,N_3747,N_3956);
or U9214 (N_9214,N_5309,N_5735);
and U9215 (N_9215,N_3221,N_3561);
and U9216 (N_9216,N_5059,N_4124);
or U9217 (N_9217,N_3957,N_5181);
xor U9218 (N_9218,N_6069,N_3738);
nor U9219 (N_9219,N_3368,N_3464);
and U9220 (N_9220,N_4803,N_4930);
nand U9221 (N_9221,N_5218,N_5404);
nor U9222 (N_9222,N_3291,N_6059);
or U9223 (N_9223,N_3356,N_3482);
or U9224 (N_9224,N_4396,N_3464);
nand U9225 (N_9225,N_5546,N_3220);
or U9226 (N_9226,N_3564,N_4256);
or U9227 (N_9227,N_4639,N_4227);
nand U9228 (N_9228,N_3471,N_5108);
and U9229 (N_9229,N_3982,N_3874);
nand U9230 (N_9230,N_5100,N_3866);
nor U9231 (N_9231,N_3901,N_5442);
nor U9232 (N_9232,N_3466,N_3914);
nor U9233 (N_9233,N_4367,N_3621);
xor U9234 (N_9234,N_4919,N_4773);
or U9235 (N_9235,N_3174,N_5710);
nand U9236 (N_9236,N_5857,N_3192);
nor U9237 (N_9237,N_4694,N_4222);
nor U9238 (N_9238,N_4756,N_5198);
and U9239 (N_9239,N_3719,N_4816);
nand U9240 (N_9240,N_3296,N_3431);
nor U9241 (N_9241,N_5593,N_3650);
and U9242 (N_9242,N_4414,N_5769);
or U9243 (N_9243,N_3805,N_3566);
xnor U9244 (N_9244,N_5229,N_5632);
nor U9245 (N_9245,N_4171,N_4065);
xnor U9246 (N_9246,N_3697,N_6015);
and U9247 (N_9247,N_5613,N_4586);
nor U9248 (N_9248,N_5583,N_4657);
nor U9249 (N_9249,N_3629,N_4650);
nor U9250 (N_9250,N_3666,N_4812);
nand U9251 (N_9251,N_4350,N_3837);
or U9252 (N_9252,N_4735,N_4799);
and U9253 (N_9253,N_4125,N_6155);
or U9254 (N_9254,N_4656,N_3475);
nor U9255 (N_9255,N_4917,N_4135);
and U9256 (N_9256,N_3644,N_5572);
xor U9257 (N_9257,N_6201,N_5837);
nand U9258 (N_9258,N_6047,N_6224);
and U9259 (N_9259,N_5686,N_4386);
and U9260 (N_9260,N_5178,N_5037);
or U9261 (N_9261,N_3587,N_4724);
xor U9262 (N_9262,N_5272,N_4514);
xor U9263 (N_9263,N_4227,N_4020);
xor U9264 (N_9264,N_3518,N_3640);
and U9265 (N_9265,N_6228,N_4796);
xor U9266 (N_9266,N_5108,N_4045);
nand U9267 (N_9267,N_5415,N_5253);
and U9268 (N_9268,N_3816,N_5575);
and U9269 (N_9269,N_3855,N_3476);
nand U9270 (N_9270,N_3943,N_5860);
nor U9271 (N_9271,N_4330,N_4948);
and U9272 (N_9272,N_6006,N_3523);
and U9273 (N_9273,N_4412,N_5118);
or U9274 (N_9274,N_4148,N_5181);
or U9275 (N_9275,N_3470,N_3245);
nand U9276 (N_9276,N_5476,N_4565);
or U9277 (N_9277,N_5482,N_4636);
or U9278 (N_9278,N_5152,N_4650);
or U9279 (N_9279,N_5054,N_3226);
or U9280 (N_9280,N_3795,N_5666);
nor U9281 (N_9281,N_4492,N_5896);
or U9282 (N_9282,N_4171,N_5325);
xor U9283 (N_9283,N_3867,N_5119);
xor U9284 (N_9284,N_5121,N_4432);
and U9285 (N_9285,N_4508,N_3161);
nor U9286 (N_9286,N_5449,N_3293);
nor U9287 (N_9287,N_3997,N_4630);
or U9288 (N_9288,N_4597,N_3250);
or U9289 (N_9289,N_5297,N_3293);
nand U9290 (N_9290,N_4494,N_5539);
xnor U9291 (N_9291,N_5103,N_4358);
or U9292 (N_9292,N_5264,N_3285);
and U9293 (N_9293,N_5429,N_3555);
or U9294 (N_9294,N_6093,N_3940);
xnor U9295 (N_9295,N_3782,N_5864);
nor U9296 (N_9296,N_5230,N_3469);
or U9297 (N_9297,N_3136,N_5557);
nor U9298 (N_9298,N_5815,N_3399);
nand U9299 (N_9299,N_6008,N_6214);
xor U9300 (N_9300,N_5699,N_4771);
or U9301 (N_9301,N_6192,N_5562);
or U9302 (N_9302,N_3913,N_3754);
nor U9303 (N_9303,N_4120,N_5873);
xnor U9304 (N_9304,N_4246,N_5079);
and U9305 (N_9305,N_4129,N_6017);
nand U9306 (N_9306,N_4361,N_4643);
nand U9307 (N_9307,N_4062,N_5556);
xor U9308 (N_9308,N_5056,N_5711);
or U9309 (N_9309,N_6150,N_5361);
xnor U9310 (N_9310,N_5091,N_4030);
nand U9311 (N_9311,N_4162,N_4595);
xnor U9312 (N_9312,N_3593,N_3855);
xor U9313 (N_9313,N_3718,N_4429);
nand U9314 (N_9314,N_6183,N_5064);
nor U9315 (N_9315,N_4409,N_5873);
or U9316 (N_9316,N_3452,N_5809);
and U9317 (N_9317,N_4471,N_3705);
or U9318 (N_9318,N_4801,N_3628);
nor U9319 (N_9319,N_3999,N_3971);
nor U9320 (N_9320,N_5268,N_6139);
and U9321 (N_9321,N_4375,N_3412);
or U9322 (N_9322,N_3603,N_3638);
and U9323 (N_9323,N_4602,N_4274);
nor U9324 (N_9324,N_4696,N_4087);
xor U9325 (N_9325,N_4277,N_3606);
or U9326 (N_9326,N_3656,N_5786);
or U9327 (N_9327,N_5296,N_5808);
nor U9328 (N_9328,N_3912,N_3883);
or U9329 (N_9329,N_3935,N_4471);
xnor U9330 (N_9330,N_6155,N_4442);
or U9331 (N_9331,N_5769,N_6130);
nand U9332 (N_9332,N_5643,N_3712);
nand U9333 (N_9333,N_5173,N_3797);
nor U9334 (N_9334,N_4604,N_3609);
xnor U9335 (N_9335,N_4254,N_3723);
and U9336 (N_9336,N_5842,N_3860);
xor U9337 (N_9337,N_3428,N_3625);
and U9338 (N_9338,N_6100,N_6204);
nand U9339 (N_9339,N_5607,N_3534);
nand U9340 (N_9340,N_4620,N_4522);
and U9341 (N_9341,N_4920,N_5802);
nand U9342 (N_9342,N_4919,N_6130);
and U9343 (N_9343,N_3680,N_5131);
and U9344 (N_9344,N_4508,N_5588);
xor U9345 (N_9345,N_3494,N_5077);
or U9346 (N_9346,N_4939,N_5540);
nand U9347 (N_9347,N_4376,N_5975);
or U9348 (N_9348,N_5200,N_4258);
nor U9349 (N_9349,N_3487,N_5054);
or U9350 (N_9350,N_4163,N_5858);
or U9351 (N_9351,N_3182,N_3776);
and U9352 (N_9352,N_3712,N_5617);
nor U9353 (N_9353,N_4600,N_4313);
nor U9354 (N_9354,N_6225,N_5332);
xor U9355 (N_9355,N_5195,N_6046);
nand U9356 (N_9356,N_3499,N_5920);
nand U9357 (N_9357,N_5866,N_5678);
nand U9358 (N_9358,N_5302,N_4355);
or U9359 (N_9359,N_3285,N_6186);
nand U9360 (N_9360,N_5648,N_5261);
xnor U9361 (N_9361,N_4722,N_4431);
nand U9362 (N_9362,N_4448,N_4801);
and U9363 (N_9363,N_4917,N_4938);
and U9364 (N_9364,N_6041,N_5678);
nand U9365 (N_9365,N_5455,N_4980);
xnor U9366 (N_9366,N_5035,N_5864);
or U9367 (N_9367,N_4746,N_3270);
or U9368 (N_9368,N_5590,N_5373);
xor U9369 (N_9369,N_5539,N_3406);
and U9370 (N_9370,N_4780,N_4018);
xor U9371 (N_9371,N_5250,N_4565);
nor U9372 (N_9372,N_3757,N_3258);
xor U9373 (N_9373,N_5605,N_5775);
nand U9374 (N_9374,N_4626,N_3279);
xor U9375 (N_9375,N_8600,N_7007);
xnor U9376 (N_9376,N_6465,N_8738);
nor U9377 (N_9377,N_8786,N_6575);
and U9378 (N_9378,N_8461,N_7534);
or U9379 (N_9379,N_6757,N_6816);
and U9380 (N_9380,N_7511,N_7648);
or U9381 (N_9381,N_7249,N_8197);
xor U9382 (N_9382,N_9245,N_6421);
nor U9383 (N_9383,N_7581,N_6297);
xor U9384 (N_9384,N_9228,N_6485);
nor U9385 (N_9385,N_8752,N_9088);
nand U9386 (N_9386,N_6909,N_8222);
xnor U9387 (N_9387,N_9337,N_8538);
or U9388 (N_9388,N_6653,N_7848);
xor U9389 (N_9389,N_7814,N_8340);
nand U9390 (N_9390,N_8821,N_9239);
or U9391 (N_9391,N_7362,N_8321);
and U9392 (N_9392,N_6902,N_8090);
and U9393 (N_9393,N_6330,N_8355);
or U9394 (N_9394,N_9001,N_7657);
or U9395 (N_9395,N_8640,N_8417);
nand U9396 (N_9396,N_7619,N_7647);
xnor U9397 (N_9397,N_8798,N_8080);
or U9398 (N_9398,N_8587,N_6413);
and U9399 (N_9399,N_8509,N_8267);
and U9400 (N_9400,N_6803,N_7269);
and U9401 (N_9401,N_6601,N_6503);
or U9402 (N_9402,N_7646,N_6837);
xor U9403 (N_9403,N_8598,N_6321);
nor U9404 (N_9404,N_6326,N_7554);
nor U9405 (N_9405,N_8290,N_9284);
or U9406 (N_9406,N_8240,N_7055);
nand U9407 (N_9407,N_9050,N_8091);
xor U9408 (N_9408,N_8151,N_8649);
nor U9409 (N_9409,N_8545,N_7587);
and U9410 (N_9410,N_8942,N_9063);
xnor U9411 (N_9411,N_8721,N_8342);
nor U9412 (N_9412,N_7734,N_7670);
and U9413 (N_9413,N_7031,N_7401);
xnor U9414 (N_9414,N_7525,N_7805);
or U9415 (N_9415,N_6592,N_8904);
nand U9416 (N_9416,N_9373,N_8081);
xnor U9417 (N_9417,N_8794,N_8814);
xnor U9418 (N_9418,N_7029,N_7136);
or U9419 (N_9419,N_8628,N_6396);
and U9420 (N_9420,N_8854,N_7968);
xnor U9421 (N_9421,N_8140,N_6839);
nor U9422 (N_9422,N_6739,N_7412);
xor U9423 (N_9423,N_9179,N_8373);
nor U9424 (N_9424,N_7142,N_9273);
and U9425 (N_9425,N_8031,N_8122);
nand U9426 (N_9426,N_8800,N_8570);
or U9427 (N_9427,N_7825,N_8848);
nor U9428 (N_9428,N_6742,N_7440);
xnor U9429 (N_9429,N_6555,N_7230);
xor U9430 (N_9430,N_6303,N_7022);
nor U9431 (N_9431,N_7414,N_6513);
or U9432 (N_9432,N_8656,N_9352);
nor U9433 (N_9433,N_8737,N_7363);
and U9434 (N_9434,N_8776,N_9296);
nor U9435 (N_9435,N_6269,N_6346);
xnor U9436 (N_9436,N_9360,N_6529);
nand U9437 (N_9437,N_8317,N_7441);
xnor U9438 (N_9438,N_9312,N_8824);
and U9439 (N_9439,N_9027,N_8660);
nand U9440 (N_9440,N_8352,N_6604);
and U9441 (N_9441,N_6843,N_9225);
nand U9442 (N_9442,N_6649,N_8826);
nand U9443 (N_9443,N_8314,N_6500);
nand U9444 (N_9444,N_6463,N_9261);
nor U9445 (N_9445,N_7216,N_6659);
nand U9446 (N_9446,N_7350,N_6397);
or U9447 (N_9447,N_8005,N_7620);
or U9448 (N_9448,N_7429,N_8382);
nand U9449 (N_9449,N_7818,N_8168);
and U9450 (N_9450,N_8356,N_6988);
or U9451 (N_9451,N_7948,N_9194);
and U9452 (N_9452,N_8788,N_8278);
nor U9453 (N_9453,N_6899,N_8616);
or U9454 (N_9454,N_6964,N_7114);
nor U9455 (N_9455,N_6965,N_7950);
xor U9456 (N_9456,N_8387,N_7280);
and U9457 (N_9457,N_7176,N_6256);
nand U9458 (N_9458,N_7580,N_9233);
nand U9459 (N_9459,N_9060,N_7309);
nand U9460 (N_9460,N_7764,N_6911);
and U9461 (N_9461,N_7863,N_6361);
or U9462 (N_9462,N_6635,N_6260);
xor U9463 (N_9463,N_7408,N_9064);
or U9464 (N_9464,N_8049,N_7205);
nand U9465 (N_9465,N_7874,N_7681);
and U9466 (N_9466,N_8816,N_6301);
nor U9467 (N_9467,N_8929,N_7531);
or U9468 (N_9468,N_7806,N_6933);
xor U9469 (N_9469,N_7491,N_9149);
and U9470 (N_9470,N_9321,N_7726);
or U9471 (N_9471,N_7660,N_8413);
and U9472 (N_9472,N_6767,N_6275);
xor U9473 (N_9473,N_7043,N_9248);
xor U9474 (N_9474,N_8588,N_6449);
nor U9475 (N_9475,N_9271,N_9250);
or U9476 (N_9476,N_8004,N_7847);
xnor U9477 (N_9477,N_6760,N_6723);
nand U9478 (N_9478,N_8180,N_6554);
and U9479 (N_9479,N_6382,N_8316);
nand U9480 (N_9480,N_7944,N_7608);
nand U9481 (N_9481,N_8535,N_8074);
nand U9482 (N_9482,N_8099,N_8397);
xnor U9483 (N_9483,N_7211,N_8131);
and U9484 (N_9484,N_7493,N_8585);
or U9485 (N_9485,N_6709,N_8840);
nand U9486 (N_9486,N_6800,N_9128);
and U9487 (N_9487,N_7779,N_8939);
nor U9488 (N_9488,N_9317,N_6669);
nor U9489 (N_9489,N_8981,N_9085);
or U9490 (N_9490,N_7191,N_8772);
or U9491 (N_9491,N_6784,N_9025);
nand U9492 (N_9492,N_9366,N_7902);
or U9493 (N_9493,N_7633,N_7084);
or U9494 (N_9494,N_6790,N_9334);
xnor U9495 (N_9495,N_7997,N_6828);
nand U9496 (N_9496,N_6618,N_8946);
nand U9497 (N_9497,N_6733,N_8315);
xnor U9498 (N_9498,N_6793,N_8652);
or U9499 (N_9499,N_8347,N_7717);
xnor U9500 (N_9500,N_7527,N_7351);
nor U9501 (N_9501,N_7277,N_7448);
nand U9502 (N_9502,N_7182,N_7039);
and U9503 (N_9503,N_8915,N_6681);
nor U9504 (N_9504,N_7922,N_8708);
or U9505 (N_9505,N_9019,N_8119);
nor U9506 (N_9506,N_8763,N_7610);
nor U9507 (N_9507,N_7175,N_9133);
or U9508 (N_9508,N_8998,N_6830);
nand U9509 (N_9509,N_7908,N_9222);
xnor U9510 (N_9510,N_6333,N_6319);
nand U9511 (N_9511,N_6289,N_8052);
and U9512 (N_9512,N_6897,N_9276);
and U9513 (N_9513,N_6329,N_6610);
nor U9514 (N_9514,N_7128,N_7710);
nand U9515 (N_9515,N_7306,N_6582);
nor U9516 (N_9516,N_6936,N_6543);
and U9517 (N_9517,N_7385,N_8420);
or U9518 (N_9518,N_9353,N_9153);
nand U9519 (N_9519,N_7424,N_6721);
nand U9520 (N_9520,N_6293,N_8033);
or U9521 (N_9521,N_7522,N_7682);
and U9522 (N_9522,N_8166,N_7539);
nand U9523 (N_9523,N_7740,N_6626);
xor U9524 (N_9524,N_9047,N_7254);
nand U9525 (N_9525,N_6937,N_7083);
nor U9526 (N_9526,N_8928,N_8808);
nand U9527 (N_9527,N_6880,N_8692);
nand U9528 (N_9528,N_7459,N_8615);
or U9529 (N_9529,N_8014,N_8305);
xor U9530 (N_9530,N_8663,N_8112);
xor U9531 (N_9531,N_7295,N_8502);
nand U9532 (N_9532,N_7947,N_6282);
nand U9533 (N_9533,N_7209,N_8626);
or U9534 (N_9534,N_6906,N_9367);
xor U9535 (N_9535,N_6580,N_7165);
and U9536 (N_9536,N_6609,N_7426);
nand U9537 (N_9537,N_7784,N_6776);
nand U9538 (N_9538,N_7015,N_8927);
xor U9539 (N_9539,N_6469,N_6950);
nand U9540 (N_9540,N_6324,N_8921);
nor U9541 (N_9541,N_8299,N_9212);
xnor U9542 (N_9542,N_7862,N_8879);
nor U9543 (N_9543,N_6922,N_6913);
nand U9544 (N_9544,N_7122,N_6692);
nand U9545 (N_9545,N_7147,N_7904);
or U9546 (N_9546,N_8855,N_7297);
nand U9547 (N_9547,N_7566,N_6797);
nor U9548 (N_9548,N_8037,N_7437);
nand U9549 (N_9549,N_7869,N_6889);
xnor U9550 (N_9550,N_8221,N_8067);
nand U9551 (N_9551,N_8066,N_7129);
nor U9552 (N_9552,N_6527,N_8256);
nor U9553 (N_9553,N_7984,N_8284);
xnor U9554 (N_9554,N_8313,N_7932);
nor U9555 (N_9555,N_7852,N_8899);
or U9556 (N_9556,N_8212,N_6312);
and U9557 (N_9557,N_9029,N_8389);
and U9558 (N_9558,N_7739,N_7152);
nand U9559 (N_9559,N_7866,N_8133);
xnor U9560 (N_9560,N_6949,N_7072);
and U9561 (N_9561,N_9270,N_9316);
and U9562 (N_9562,N_8492,N_7312);
and U9563 (N_9563,N_6308,N_7893);
xor U9564 (N_9564,N_6758,N_6283);
nand U9565 (N_9565,N_6451,N_6679);
and U9566 (N_9566,N_8071,N_9286);
nor U9567 (N_9567,N_7415,N_7074);
or U9568 (N_9568,N_7960,N_8274);
or U9569 (N_9569,N_7000,N_7693);
and U9570 (N_9570,N_7803,N_8390);
xor U9571 (N_9571,N_7630,N_6625);
and U9572 (N_9572,N_6416,N_6300);
or U9573 (N_9573,N_8846,N_6887);
nand U9574 (N_9574,N_9100,N_6286);
nor U9575 (N_9575,N_8597,N_6515);
or U9576 (N_9576,N_7659,N_6380);
xnor U9577 (N_9577,N_7366,N_7578);
nand U9578 (N_9578,N_7314,N_8232);
nand U9579 (N_9579,N_6261,N_6518);
or U9580 (N_9580,N_9302,N_6440);
xnor U9581 (N_9581,N_9135,N_8963);
or U9582 (N_9582,N_9247,N_8760);
and U9583 (N_9583,N_7497,N_7365);
nand U9584 (N_9584,N_7841,N_6819);
xor U9585 (N_9585,N_8845,N_6438);
nor U9586 (N_9586,N_7969,N_6987);
nand U9587 (N_9587,N_8144,N_6255);
and U9588 (N_9588,N_8041,N_8766);
nor U9589 (N_9589,N_8498,N_7023);
nand U9590 (N_9590,N_6314,N_9189);
xor U9591 (N_9591,N_6944,N_8634);
and U9592 (N_9592,N_6672,N_7576);
nor U9593 (N_9593,N_7434,N_8124);
xnor U9594 (N_9594,N_6362,N_8251);
or U9595 (N_9595,N_6655,N_6848);
xnor U9596 (N_9596,N_7499,N_7971);
xnor U9597 (N_9597,N_8398,N_8697);
xor U9598 (N_9598,N_8249,N_7650);
nand U9599 (N_9599,N_7210,N_7262);
nand U9600 (N_9600,N_7669,N_8185);
and U9601 (N_9601,N_7172,N_6821);
xnor U9602 (N_9602,N_9055,N_7789);
nand U9603 (N_9603,N_6379,N_7958);
nor U9604 (N_9604,N_6611,N_8727);
nand U9605 (N_9605,N_7939,N_6586);
nor U9606 (N_9606,N_7416,N_9305);
or U9607 (N_9607,N_7882,N_8283);
or U9608 (N_9608,N_9372,N_8505);
and U9609 (N_9609,N_6869,N_6491);
nor U9610 (N_9610,N_7026,N_8730);
nor U9611 (N_9611,N_8228,N_9182);
nand U9612 (N_9612,N_6281,N_7452);
xnor U9613 (N_9613,N_9026,N_7141);
nand U9614 (N_9614,N_9127,N_7937);
nand U9615 (N_9615,N_6752,N_7180);
xnor U9616 (N_9616,N_7138,N_8764);
and U9617 (N_9617,N_6254,N_7329);
nand U9618 (N_9618,N_8474,N_8269);
or U9619 (N_9619,N_7732,N_8261);
xnor U9620 (N_9620,N_7632,N_8702);
and U9621 (N_9621,N_7318,N_9079);
xnor U9622 (N_9622,N_8436,N_8662);
nand U9623 (N_9623,N_8672,N_8380);
nand U9624 (N_9624,N_9186,N_7399);
xor U9625 (N_9625,N_9132,N_6863);
xnor U9626 (N_9626,N_9152,N_9341);
nor U9627 (N_9627,N_7342,N_9291);
and U9628 (N_9628,N_7133,N_8577);
and U9629 (N_9629,N_9184,N_7081);
or U9630 (N_9630,N_8886,N_8271);
nand U9631 (N_9631,N_7560,N_8667);
and U9632 (N_9632,N_7406,N_6411);
and U9633 (N_9633,N_9036,N_8980);
xor U9634 (N_9634,N_8837,N_8404);
nand U9635 (N_9635,N_9211,N_8345);
and U9636 (N_9636,N_7845,N_7387);
and U9637 (N_9637,N_8010,N_7905);
xor U9638 (N_9638,N_6876,N_8025);
nand U9639 (N_9639,N_7687,N_8924);
and U9640 (N_9640,N_9289,N_7676);
and U9641 (N_9641,N_6896,N_8114);
nor U9642 (N_9642,N_8869,N_9002);
nor U9643 (N_9643,N_8215,N_7384);
or U9644 (N_9644,N_8349,N_8643);
xor U9645 (N_9645,N_7132,N_7891);
xor U9646 (N_9646,N_8429,N_9150);
nand U9647 (N_9647,N_6483,N_9071);
nor U9648 (N_9648,N_8032,N_8252);
and U9649 (N_9649,N_6424,N_8956);
xor U9650 (N_9650,N_8078,N_9035);
xnor U9651 (N_9651,N_7060,N_6766);
nand U9652 (N_9652,N_7698,N_8027);
and U9653 (N_9653,N_6327,N_6557);
xor U9654 (N_9654,N_7642,N_6414);
nand U9655 (N_9655,N_9345,N_6455);
or U9656 (N_9656,N_8987,N_8742);
and U9657 (N_9657,N_8582,N_7322);
and U9658 (N_9658,N_7494,N_7671);
and U9659 (N_9659,N_9313,N_7354);
xnor U9660 (N_9660,N_9370,N_6967);
or U9661 (N_9661,N_7228,N_9160);
nor U9662 (N_9662,N_6394,N_8900);
xor U9663 (N_9663,N_9008,N_7278);
nor U9664 (N_9664,N_6799,N_6663);
and U9665 (N_9665,N_7054,N_7008);
nor U9666 (N_9666,N_7294,N_8160);
or U9667 (N_9667,N_9303,N_7773);
nand U9668 (N_9668,N_7906,N_9126);
nand U9669 (N_9669,N_8281,N_6400);
and U9670 (N_9670,N_7268,N_7643);
and U9671 (N_9671,N_6901,N_8931);
nand U9672 (N_9672,N_6794,N_7308);
or U9673 (N_9673,N_9246,N_8359);
nor U9674 (N_9674,N_7001,N_8477);
nor U9675 (N_9675,N_6629,N_8209);
nand U9676 (N_9676,N_6632,N_8045);
or U9677 (N_9677,N_8534,N_8207);
and U9678 (N_9678,N_8797,N_8830);
or U9679 (N_9679,N_6385,N_9151);
nor U9680 (N_9680,N_9299,N_8948);
nor U9681 (N_9681,N_7146,N_7327);
nand U9682 (N_9682,N_7157,N_8400);
nor U9683 (N_9683,N_8177,N_8077);
or U9684 (N_9684,N_7961,N_7034);
or U9685 (N_9685,N_8444,N_7068);
or U9686 (N_9686,N_7380,N_7339);
or U9687 (N_9687,N_6690,N_7194);
nand U9688 (N_9688,N_8792,N_9307);
xnor U9689 (N_9689,N_6363,N_8754);
or U9690 (N_9690,N_9145,N_7320);
nor U9691 (N_9691,N_6569,N_7481);
xnor U9692 (N_9692,N_8415,N_7995);
nor U9693 (N_9693,N_9265,N_7768);
and U9694 (N_9694,N_7056,N_7915);
and U9695 (N_9695,N_9269,N_6983);
or U9696 (N_9696,N_8455,N_9012);
nand U9697 (N_9697,N_6558,N_8009);
xor U9698 (N_9698,N_8453,N_6372);
xor U9699 (N_9699,N_6576,N_9213);
xnor U9700 (N_9700,N_7204,N_8109);
nor U9701 (N_9701,N_7436,N_7025);
xnor U9702 (N_9702,N_6975,N_7974);
and U9703 (N_9703,N_8482,N_8134);
and U9704 (N_9704,N_7876,N_6633);
nor U9705 (N_9705,N_6309,N_9336);
nor U9706 (N_9706,N_7011,N_7073);
xnor U9707 (N_9707,N_9268,N_8991);
and U9708 (N_9708,N_9175,N_8017);
xnor U9709 (N_9709,N_7198,N_7722);
xnor U9710 (N_9710,N_7087,N_8353);
nor U9711 (N_9711,N_8135,N_7872);
xor U9712 (N_9712,N_7767,N_7583);
nor U9713 (N_9713,N_9314,N_7530);
or U9714 (N_9714,N_8472,N_8083);
nand U9715 (N_9715,N_6867,N_6284);
or U9716 (N_9716,N_7118,N_9219);
xnor U9717 (N_9717,N_7959,N_9118);
or U9718 (N_9718,N_8546,N_6818);
and U9719 (N_9719,N_7106,N_6992);
or U9720 (N_9720,N_7467,N_6295);
nand U9721 (N_9721,N_8716,N_7067);
xor U9722 (N_9722,N_7769,N_6395);
and U9723 (N_9723,N_8497,N_7854);
and U9724 (N_9724,N_9348,N_9032);
or U9725 (N_9725,N_8152,N_9342);
and U9726 (N_9726,N_8046,N_6251);
or U9727 (N_9727,N_6972,N_8254);
nand U9728 (N_9728,N_8493,N_8676);
nand U9729 (N_9729,N_6699,N_7382);
nor U9730 (N_9730,N_7590,N_7519);
or U9731 (N_9731,N_9005,N_6587);
nand U9732 (N_9732,N_8319,N_7795);
xnor U9733 (N_9733,N_8079,N_6460);
xnor U9734 (N_9734,N_6805,N_7267);
or U9735 (N_9735,N_7163,N_7881);
and U9736 (N_9736,N_8035,N_8146);
nand U9737 (N_9737,N_7685,N_8393);
or U9738 (N_9738,N_7575,N_7045);
or U9739 (N_9739,N_8703,N_6780);
or U9740 (N_9740,N_7193,N_8793);
nand U9741 (N_9741,N_7809,N_8401);
nor U9742 (N_9742,N_7229,N_8849);
and U9743 (N_9743,N_6957,N_6963);
nor U9744 (N_9744,N_8510,N_7552);
or U9745 (N_9745,N_9130,N_8147);
or U9746 (N_9746,N_8377,N_8718);
nand U9747 (N_9747,N_6791,N_9041);
and U9748 (N_9748,N_9154,N_6928);
and U9749 (N_9749,N_7158,N_8611);
and U9750 (N_9750,N_6871,N_8007);
nor U9751 (N_9751,N_8013,N_6367);
and U9752 (N_9752,N_9287,N_8696);
nand U9753 (N_9753,N_6872,N_8308);
xnor U9754 (N_9754,N_9106,N_7462);
xor U9755 (N_9755,N_6546,N_7456);
nand U9756 (N_9756,N_6296,N_9096);
or U9757 (N_9757,N_8562,N_8142);
nor U9758 (N_9758,N_7753,N_7232);
nor U9759 (N_9759,N_9227,N_9343);
or U9760 (N_9760,N_7759,N_8011);
and U9761 (N_9761,N_8129,N_7987);
and U9762 (N_9762,N_7832,N_6774);
nor U9763 (N_9763,N_7201,N_8485);
and U9764 (N_9764,N_8481,N_7729);
nand U9765 (N_9765,N_7990,N_8118);
nor U9766 (N_9766,N_8571,N_9292);
nor U9767 (N_9767,N_9010,N_8996);
or U9768 (N_9768,N_7070,N_7340);
and U9769 (N_9769,N_6664,N_7461);
nor U9770 (N_9770,N_7392,N_8875);
nor U9771 (N_9771,N_7220,N_8426);
or U9772 (N_9772,N_8767,N_8822);
nor U9773 (N_9773,N_7367,N_8919);
nand U9774 (N_9774,N_8671,N_7256);
nand U9775 (N_9775,N_7250,N_9331);
or U9776 (N_9776,N_7970,N_6608);
or U9777 (N_9777,N_6636,N_8084);
xnor U9778 (N_9778,N_6858,N_8960);
nand U9779 (N_9779,N_7444,N_8819);
nand U9780 (N_9780,N_7121,N_6368);
nand U9781 (N_9781,N_6510,N_6813);
nand U9782 (N_9782,N_8522,N_6698);
and U9783 (N_9783,N_6998,N_8250);
xnor U9784 (N_9784,N_8969,N_6563);
nand U9785 (N_9785,N_8424,N_6695);
nand U9786 (N_9786,N_7478,N_7162);
or U9787 (N_9787,N_8823,N_6594);
xnor U9788 (N_9788,N_7235,N_6750);
nand U9789 (N_9789,N_8665,N_7875);
nor U9790 (N_9790,N_9031,N_6859);
and U9791 (N_9791,N_8661,N_7496);
and U9792 (N_9792,N_8694,N_9216);
and U9793 (N_9793,N_6792,N_9322);
and U9794 (N_9794,N_7471,N_8882);
or U9795 (N_9795,N_7701,N_7975);
xnor U9796 (N_9796,N_9134,N_8992);
and U9797 (N_9797,N_6701,N_8171);
and U9798 (N_9798,N_8691,N_8890);
xnor U9799 (N_9799,N_8555,N_6645);
or U9800 (N_9800,N_6966,N_7774);
nand U9801 (N_9801,N_8839,N_8573);
xor U9802 (N_9802,N_7833,N_9328);
nor U9803 (N_9803,N_9263,N_8548);
or U9804 (N_9804,N_6516,N_8515);
nor U9805 (N_9805,N_7108,N_6404);
nand U9806 (N_9806,N_6401,N_7064);
and U9807 (N_9807,N_6812,N_8062);
and U9808 (N_9808,N_8275,N_7186);
and U9809 (N_9809,N_8392,N_6494);
and U9810 (N_9810,N_8096,N_7510);
or U9811 (N_9811,N_6781,N_7549);
nor U9812 (N_9812,N_6487,N_6407);
or U9813 (N_9813,N_8264,N_7913);
nor U9814 (N_9814,N_8674,N_9094);
nand U9815 (N_9815,N_8954,N_7099);
or U9816 (N_9816,N_6727,N_7639);
and U9817 (N_9817,N_7185,N_7955);
and U9818 (N_9818,N_8194,N_8889);
xor U9819 (N_9819,N_8399,N_9249);
nor U9820 (N_9820,N_8543,N_6728);
nor U9821 (N_9821,N_6941,N_6985);
or U9822 (N_9822,N_7279,N_6638);
xnor U9823 (N_9823,N_8892,N_8309);
xor U9824 (N_9824,N_8076,N_6924);
xnor U9825 (N_9825,N_7187,N_6360);
nand U9826 (N_9826,N_8995,N_6864);
nand U9827 (N_9827,N_9282,N_6409);
xnor U9828 (N_9828,N_8906,N_9048);
or U9829 (N_9829,N_6622,N_9374);
nor U9830 (N_9830,N_6602,N_7747);
or U9831 (N_9831,N_8744,N_6550);
xor U9832 (N_9832,N_8881,N_8246);
nor U9833 (N_9833,N_6743,N_7719);
nand U9834 (N_9834,N_8645,N_7914);
nor U9835 (N_9835,N_6662,N_8951);
xnor U9836 (N_9836,N_7501,N_9170);
nor U9837 (N_9837,N_8876,N_7602);
nor U9838 (N_9838,N_6686,N_9200);
nor U9839 (N_9839,N_6322,N_7652);
nor U9840 (N_9840,N_7086,N_6884);
xor U9841 (N_9841,N_6802,N_7787);
xnor U9842 (N_9842,N_8864,N_8866);
xor U9843 (N_9843,N_7839,N_9371);
xnor U9844 (N_9844,N_6676,N_6665);
nand U9845 (N_9845,N_8847,N_7730);
xor U9846 (N_9846,N_7802,N_7164);
nand U9847 (N_9847,N_6375,N_6895);
xnor U9848 (N_9848,N_7219,N_8569);
nand U9849 (N_9849,N_7736,N_7896);
xnor U9850 (N_9850,N_8449,N_6731);
and U9851 (N_9851,N_7266,N_7888);
xor U9852 (N_9852,N_7047,N_8952);
and U9853 (N_9853,N_7556,N_9148);
nor U9854 (N_9854,N_6343,N_9325);
nor U9855 (N_9855,N_7791,N_8396);
and U9856 (N_9856,N_7668,N_8291);
or U9857 (N_9857,N_8181,N_9364);
nand U9858 (N_9858,N_7103,N_7075);
and U9859 (N_9859,N_9164,N_8000);
or U9860 (N_9860,N_6570,N_8302);
and U9861 (N_9861,N_7243,N_9192);
nand U9862 (N_9862,N_8105,N_8550);
nand U9863 (N_9863,N_8051,N_6999);
or U9864 (N_9864,N_6693,N_6267);
or U9865 (N_9865,N_6700,N_7479);
nand U9866 (N_9866,N_9242,N_6994);
or U9867 (N_9867,N_8631,N_8331);
and U9868 (N_9868,N_8053,N_8043);
nand U9869 (N_9869,N_6705,N_7672);
or U9870 (N_9870,N_7584,N_9021);
nand U9871 (N_9871,N_6833,N_6276);
or U9872 (N_9872,N_6268,N_6271);
or U9873 (N_9873,N_7601,N_8178);
nor U9874 (N_9874,N_6551,N_7526);
and U9875 (N_9875,N_7208,N_7615);
or U9876 (N_9876,N_8016,N_7418);
nor U9877 (N_9877,N_8050,N_8828);
nor U9878 (N_9878,N_6588,N_9335);
nor U9879 (N_9879,N_8973,N_8195);
and U9880 (N_9880,N_6369,N_6702);
and U9881 (N_9881,N_8637,N_7986);
and U9882 (N_9882,N_6724,N_7094);
nor U9883 (N_9883,N_7903,N_7282);
xor U9884 (N_9884,N_8297,N_7694);
and U9885 (N_9885,N_6893,N_7543);
xnor U9886 (N_9886,N_9156,N_6436);
nand U9887 (N_9887,N_7381,N_8741);
nor U9888 (N_9888,N_6619,N_7131);
and U9889 (N_9889,N_7628,N_7112);
xnor U9890 (N_9890,N_6671,N_6512);
or U9891 (N_9891,N_7623,N_6841);
nor U9892 (N_9892,N_7330,N_7224);
nand U9893 (N_9893,N_6755,N_8812);
nand U9894 (N_9894,N_7038,N_8769);
or U9895 (N_9895,N_7951,N_6265);
nand U9896 (N_9896,N_8095,N_8117);
nor U9897 (N_9897,N_9236,N_9272);
nand U9898 (N_9898,N_6612,N_7982);
nor U9899 (N_9899,N_7617,N_8435);
or U9900 (N_9900,N_7690,N_8476);
nor U9901 (N_9901,N_7829,N_7030);
and U9902 (N_9902,N_8907,N_6390);
nand U9903 (N_9903,N_6855,N_7231);
nand U9904 (N_9904,N_6980,N_6389);
and U9905 (N_9905,N_8438,N_8784);
nor U9906 (N_9906,N_9290,N_8423);
nand U9907 (N_9907,N_7311,N_9338);
nand U9908 (N_9908,N_8121,N_9259);
nor U9909 (N_9909,N_6938,N_7020);
nor U9910 (N_9910,N_8930,N_6579);
or U9911 (N_9911,N_8174,N_7754);
xor U9912 (N_9912,N_7972,N_6259);
nand U9913 (N_9913,N_6526,N_7475);
xor U9914 (N_9914,N_7884,N_8926);
and U9915 (N_9915,N_7259,N_7304);
nand U9916 (N_9916,N_7537,N_7731);
or U9917 (N_9917,N_8541,N_6885);
nor U9918 (N_9918,N_7313,N_9199);
xor U9919 (N_9919,N_8560,N_7196);
nor U9920 (N_9920,N_6874,N_8728);
or U9921 (N_9921,N_9190,N_6822);
or U9922 (N_9922,N_7474,N_9053);
and U9923 (N_9923,N_6703,N_8111);
or U9924 (N_9924,N_7513,N_9168);
nor U9925 (N_9925,N_8609,N_8938);
nand U9926 (N_9926,N_8686,N_8128);
nor U9927 (N_9927,N_8338,N_6849);
nor U9928 (N_9928,N_7824,N_6856);
nand U9929 (N_9929,N_8858,N_6307);
or U9930 (N_9930,N_7455,N_7514);
nand U9931 (N_9931,N_7263,N_7453);
nand U9932 (N_9932,N_8501,N_8959);
and U9933 (N_9933,N_8780,N_7801);
nand U9934 (N_9934,N_7107,N_7489);
nand U9935 (N_9935,N_7596,N_6392);
and U9936 (N_9936,N_7323,N_7857);
and U9937 (N_9937,N_7167,N_6561);
or U9938 (N_9938,N_7240,N_7473);
nor U9939 (N_9939,N_6642,N_7223);
nor U9940 (N_9940,N_8198,N_7046);
and U9941 (N_9941,N_6320,N_6623);
xnor U9942 (N_9942,N_7345,N_7430);
nand U9943 (N_9943,N_7236,N_8351);
and U9944 (N_9944,N_7161,N_6403);
nand U9945 (N_9945,N_6809,N_8638);
or U9946 (N_9946,N_6959,N_6535);
or U9947 (N_9947,N_8773,N_7341);
xnor U9948 (N_9948,N_8862,N_6870);
nor U9949 (N_9949,N_6423,N_8685);
and U9950 (N_9950,N_9244,N_6328);
nand U9951 (N_9951,N_8026,N_8057);
nor U9952 (N_9952,N_8410,N_8922);
and U9953 (N_9953,N_7895,N_6746);
or U9954 (N_9954,N_9191,N_8748);
nand U9955 (N_9955,N_9254,N_8478);
nand U9956 (N_9956,N_9176,N_7134);
nand U9957 (N_9957,N_7778,N_8789);
or U9958 (N_9958,N_8475,N_6477);
and U9959 (N_9959,N_7954,N_6501);
xnor U9960 (N_9960,N_6883,N_7355);
nor U9961 (N_9961,N_7640,N_6347);
nor U9962 (N_9962,N_9281,N_7135);
nand U9963 (N_9963,N_8213,N_6521);
nand U9964 (N_9964,N_7356,N_8130);
xnor U9965 (N_9965,N_7931,N_9349);
and U9966 (N_9966,N_7838,N_7546);
xnor U9967 (N_9967,N_8834,N_7333);
nor U9968 (N_9968,N_7195,N_6948);
nor U9969 (N_9969,N_6564,N_9052);
and U9970 (N_9970,N_8666,N_7091);
or U9971 (N_9971,N_8205,N_7512);
and U9972 (N_9972,N_8511,N_7999);
or U9973 (N_9973,N_6511,N_8580);
xnor U9974 (N_9974,N_7725,N_8912);
xor U9975 (N_9975,N_9278,N_7049);
nor U9976 (N_9976,N_8148,N_7388);
nand U9977 (N_9977,N_7174,N_6764);
nor U9978 (N_9978,N_7819,N_7979);
xor U9979 (N_9979,N_8591,N_6599);
xnor U9980 (N_9980,N_9260,N_7535);
nand U9981 (N_9981,N_7244,N_7618);
and U9982 (N_9982,N_7383,N_8669);
and U9983 (N_9983,N_7005,N_8561);
nor U9984 (N_9984,N_7909,N_6675);
or U9985 (N_9985,N_8378,N_7100);
or U9986 (N_9986,N_6926,N_8061);
nor U9987 (N_9987,N_8279,N_8329);
or U9988 (N_9988,N_7688,N_9294);
nor U9989 (N_9989,N_7447,N_8736);
nor U9990 (N_9990,N_7919,N_8235);
xor U9991 (N_9991,N_6748,N_8625);
xnor U9992 (N_9992,N_7589,N_7994);
and U9993 (N_9993,N_7721,N_7290);
and U9994 (N_9994,N_8260,N_8107);
xor U9995 (N_9995,N_8878,N_8211);
nand U9996 (N_9996,N_6433,N_6763);
nor U9997 (N_9997,N_8082,N_7260);
nor U9998 (N_9998,N_8223,N_7760);
nor U9999 (N_9999,N_9142,N_6278);
nor U10000 (N_10000,N_7533,N_8953);
xnor U10001 (N_10001,N_8272,N_7460);
or U10002 (N_10002,N_6549,N_7271);
nor U10003 (N_10003,N_6277,N_6956);
xor U10004 (N_10004,N_8072,N_7842);
and U10005 (N_10005,N_6991,N_6531);
and U10006 (N_10006,N_7684,N_7457);
xnor U10007 (N_10007,N_9185,N_7410);
xor U10008 (N_10008,N_6886,N_8778);
or U10009 (N_10009,N_7844,N_8815);
and U10010 (N_10010,N_6383,N_7941);
or U10011 (N_10011,N_7911,N_7713);
or U10012 (N_10012,N_9174,N_7930);
and U10013 (N_10013,N_7179,N_6448);
nor U10014 (N_10014,N_9221,N_8108);
and U10015 (N_10015,N_7014,N_7458);
and U10016 (N_10016,N_6507,N_8432);
and U10017 (N_10017,N_8042,N_6473);
xnor U10018 (N_10018,N_8903,N_8524);
nand U10019 (N_10019,N_9208,N_8857);
nand U10020 (N_10020,N_6921,N_7125);
and U10021 (N_10021,N_8012,N_6888);
xor U10022 (N_10022,N_7337,N_6506);
nor U10023 (N_10023,N_7358,N_8993);
xnor U10024 (N_10024,N_7503,N_7641);
or U10025 (N_10025,N_6796,N_8358);
nor U10026 (N_10026,N_8421,N_9091);
nor U10027 (N_10027,N_7302,N_6304);
and U10028 (N_10028,N_7663,N_7662);
and U10029 (N_10029,N_7445,N_6955);
and U10030 (N_10030,N_8827,N_8967);
xor U10031 (N_10031,N_6737,N_8363);
nor U10032 (N_10032,N_6597,N_6318);
nand U10033 (N_10033,N_7468,N_9363);
or U10034 (N_10034,N_9163,N_8103);
nand U10035 (N_10035,N_8255,N_9119);
nor U10036 (N_10036,N_7901,N_9095);
xnor U10037 (N_10037,N_7148,N_6850);
nand U10038 (N_10038,N_8700,N_8266);
xor U10039 (N_10039,N_6514,N_9122);
xnor U10040 (N_10040,N_8311,N_6882);
and U10041 (N_10041,N_7343,N_7894);
nor U10042 (N_10042,N_6285,N_6970);
nor U10043 (N_10043,N_7495,N_7218);
and U10044 (N_10044,N_8684,N_8293);
nand U10045 (N_10045,N_8286,N_7956);
or U10046 (N_10046,N_8070,N_8723);
or U10047 (N_10047,N_8430,N_7743);
nor U10048 (N_10048,N_7454,N_8262);
xnor U10049 (N_10049,N_9274,N_8932);
or U10050 (N_10050,N_8483,N_9167);
xnor U10051 (N_10051,N_9231,N_7206);
nand U10052 (N_10052,N_6680,N_9115);
nor U10053 (N_10053,N_8724,N_9365);
xor U10054 (N_10054,N_9086,N_6331);
nand U10055 (N_10055,N_8434,N_8999);
or U10056 (N_10056,N_9196,N_8937);
xor U10057 (N_10057,N_8162,N_8715);
xor U10058 (N_10058,N_6262,N_7592);
xor U10059 (N_10059,N_6710,N_9326);
or U10060 (N_10060,N_9125,N_9201);
or U10061 (N_10061,N_8156,N_9362);
or U10062 (N_10062,N_9000,N_8532);
nor U10063 (N_10063,N_6272,N_8802);
nor U10064 (N_10064,N_8623,N_8457);
and U10065 (N_10065,N_7212,N_8917);
and U10066 (N_10066,N_6951,N_6808);
nand U10067 (N_10067,N_8790,N_9304);
and U10068 (N_10068,N_9034,N_8182);
and U10069 (N_10069,N_7389,N_7810);
xnor U10070 (N_10070,N_6939,N_7611);
nand U10071 (N_10071,N_8528,N_6997);
nor U10072 (N_10072,N_8586,N_8354);
or U10073 (N_10073,N_7606,N_7855);
or U10074 (N_10074,N_8214,N_8579);
xor U10075 (N_10075,N_7058,N_7397);
nor U10076 (N_10076,N_9062,N_8173);
nor U10077 (N_10077,N_7785,N_8659);
nand U10078 (N_10078,N_7757,N_9124);
nand U10079 (N_10079,N_8898,N_8282);
nand U10080 (N_10080,N_9003,N_6778);
or U10081 (N_10081,N_7804,N_8094);
and U10082 (N_10082,N_7998,N_6717);
nand U10083 (N_10083,N_9043,N_6915);
xor U10084 (N_10084,N_8918,N_7949);
and U10085 (N_10085,N_9082,N_6356);
nand U10086 (N_10086,N_6398,N_7991);
nor U10087 (N_10087,N_8106,N_8158);
xor U10088 (N_10088,N_6565,N_6486);
nand U10089 (N_10089,N_9315,N_6393);
nor U10090 (N_10090,N_7667,N_8339);
or U10091 (N_10091,N_7558,N_6355);
xor U10092 (N_10092,N_7567,N_8451);
nor U10093 (N_10093,N_9089,N_6652);
xor U10094 (N_10094,N_8619,N_7661);
or U10095 (N_10095,N_9166,N_9230);
nand U10096 (N_10096,N_9102,N_6775);
or U10097 (N_10097,N_6787,N_7417);
nand U10098 (N_10098,N_6788,N_8803);
xnor U10099 (N_10099,N_6548,N_6759);
nand U10100 (N_10100,N_8564,N_8018);
or U10101 (N_10101,N_7069,N_8259);
nor U10102 (N_10102,N_8239,N_6977);
nor U10103 (N_10103,N_7101,N_8366);
nor U10104 (N_10104,N_7315,N_6958);
and U10105 (N_10105,N_8348,N_8567);
or U10106 (N_10106,N_7599,N_6696);
xor U10107 (N_10107,N_7547,N_7283);
nand U10108 (N_10108,N_6725,N_8936);
nor U10109 (N_10109,N_9147,N_7423);
xor U10110 (N_10110,N_8920,N_7925);
nand U10111 (N_10111,N_6298,N_6496);
nand U10112 (N_10112,N_7607,N_7521);
or U10113 (N_10113,N_8120,N_7178);
nor U10114 (N_10114,N_8233,N_7920);
nand U10115 (N_10115,N_7470,N_8357);
or U10116 (N_10116,N_8188,N_7727);
or U10117 (N_10117,N_9030,N_6651);
nor U10118 (N_10118,N_6722,N_7241);
nand U10119 (N_10119,N_8542,N_8055);
nor U10120 (N_10120,N_6426,N_7335);
xnor U10121 (N_10121,N_6694,N_7796);
or U10122 (N_10122,N_6835,N_8381);
nand U10123 (N_10123,N_7598,N_6325);
and U10124 (N_10124,N_8851,N_6879);
and U10125 (N_10125,N_7756,N_6358);
xor U10126 (N_10126,N_7899,N_6860);
and U10127 (N_10127,N_7821,N_7624);
xor U10128 (N_10128,N_8552,N_9098);
xor U10129 (N_10129,N_8747,N_7274);
nand U10130 (N_10130,N_8856,N_8581);
and U10131 (N_10131,N_8762,N_7202);
nand U10132 (N_10132,N_7016,N_8880);
and U10133 (N_10133,N_6410,N_9295);
nor U10134 (N_10134,N_8375,N_9172);
and U10135 (N_10135,N_6990,N_6447);
or U10136 (N_10136,N_6335,N_8088);
or U10137 (N_10137,N_8328,N_7427);
nor U10138 (N_10138,N_8295,N_6446);
xnor U10139 (N_10139,N_8132,N_7035);
nor U10140 (N_10140,N_6968,N_7472);
nand U10141 (N_10141,N_6704,N_7177);
nand U10142 (N_10142,N_9072,N_7130);
or U10143 (N_10143,N_7559,N_8885);
nor U10144 (N_10144,N_6761,N_8020);
and U10145 (N_10145,N_8394,N_7018);
and U10146 (N_10146,N_7831,N_6553);
nor U10147 (N_10147,N_9051,N_8719);
nand U10148 (N_10148,N_7963,N_8935);
xor U10149 (N_10149,N_7518,N_7080);
nand U10150 (N_10150,N_8761,N_7588);
nor U10151 (N_10151,N_8137,N_8325);
nor U10152 (N_10152,N_9356,N_7105);
nor U10153 (N_10153,N_6480,N_7189);
or U10154 (N_10154,N_8750,N_8949);
nor U10155 (N_10155,N_8098,N_8986);
nor U10156 (N_10156,N_8933,N_8572);
xnor U10157 (N_10157,N_8968,N_9024);
and U10158 (N_10158,N_7528,N_6350);
xnor U10159 (N_10159,N_8484,N_9318);
and U10160 (N_10160,N_7858,N_7369);
and U10161 (N_10161,N_8335,N_8832);
or U10162 (N_10162,N_8097,N_9066);
nand U10163 (N_10163,N_8679,N_8529);
xor U10164 (N_10164,N_6310,N_7515);
nand U10165 (N_10165,N_6453,N_6590);
and U10166 (N_10166,N_8408,N_6479);
or U10167 (N_10167,N_7656,N_8159);
nor U10168 (N_10168,N_7032,N_6646);
nor U10169 (N_10169,N_9141,N_6641);
nand U10170 (N_10170,N_9116,N_6357);
nand U10171 (N_10171,N_7199,N_8288);
xnor U10172 (N_10172,N_9301,N_8468);
and U10173 (N_10173,N_9324,N_6323);
xor U10174 (N_10174,N_8491,N_7723);
xnor U10175 (N_10175,N_8422,N_8877);
nor U10176 (N_10176,N_7849,N_7144);
or U10177 (N_10177,N_6373,N_8236);
or U10178 (N_10178,N_8307,N_8775);
nor U10179 (N_10179,N_7597,N_9046);
xnor U10180 (N_10180,N_7708,N_6782);
nor U10181 (N_10181,N_8087,N_8101);
nor U10182 (N_10182,N_7078,N_6640);
xor U10183 (N_10183,N_7036,N_6720);
nand U10184 (N_10184,N_7421,N_7517);
nor U10185 (N_10185,N_8170,N_7300);
nand U10186 (N_10186,N_7319,N_8589);
nand U10187 (N_10187,N_7758,N_7052);
nand U10188 (N_10188,N_8958,N_6419);
or U10189 (N_10189,N_6711,N_6471);
or U10190 (N_10190,N_6831,N_6729);
or U10191 (N_10191,N_6257,N_6660);
and U10192 (N_10192,N_7237,N_7867);
nor U10193 (N_10193,N_9028,N_6337);
and U10194 (N_10194,N_9323,N_8226);
nand U10195 (N_10195,N_9306,N_7993);
and U10196 (N_10196,N_7780,N_8289);
nor U10197 (N_10197,N_7321,N_8533);
and U10198 (N_10198,N_7137,N_6751);
and U10199 (N_10199,N_7276,N_8654);
and U10200 (N_10200,N_8343,N_6556);
and U10201 (N_10201,N_8405,N_6930);
nor U10202 (N_10202,N_6273,N_8150);
and U10203 (N_10203,N_9129,N_8668);
xor U10204 (N_10204,N_9288,N_8294);
xnor U10205 (N_10205,N_8632,N_8804);
nor U10206 (N_10206,N_7061,N_7487);
and U10207 (N_10207,N_9120,N_7173);
nor U10208 (N_10208,N_8425,N_6459);
and U10209 (N_10209,N_8911,N_8818);
xor U10210 (N_10210,N_9232,N_9020);
xor U10211 (N_10211,N_7557,N_6868);
or U10212 (N_10212,N_7168,N_6596);
or U10213 (N_10213,N_7181,N_8568);
nand U10214 (N_10214,N_8596,N_7257);
xor U10215 (N_10215,N_8883,N_9069);
and U10216 (N_10216,N_6943,N_6508);
nand U10217 (N_10217,N_8191,N_7490);
and U10218 (N_10218,N_9235,N_6923);
or U10219 (N_10219,N_7751,N_8496);
and U10220 (N_10220,N_6730,N_7378);
nand U10221 (N_10221,N_8731,N_8058);
nand U10222 (N_10222,N_6354,N_8220);
nor U10223 (N_10223,N_9197,N_9327);
xor U10224 (N_10224,N_7609,N_7715);
nor U10225 (N_10225,N_7936,N_6399);
xnor U10226 (N_10226,N_6756,N_9183);
xor U10227 (N_10227,N_6942,N_8751);
nand U10228 (N_10228,N_8673,N_8508);
nand U10229 (N_10229,N_6538,N_7783);
or U10230 (N_10230,N_7403,N_6525);
and U10231 (N_10231,N_7523,N_9180);
nor U10232 (N_10232,N_7090,N_8141);
nand U10233 (N_10233,N_7709,N_6735);
or U10234 (N_10234,N_7465,N_8304);
xnor U10235 (N_10235,N_9056,N_6732);
nor U10236 (N_10236,N_7402,N_6661);
nor U10237 (N_10237,N_6978,N_7123);
or U10238 (N_10238,N_8153,N_8592);
xor U10239 (N_10239,N_6517,N_9355);
and U10240 (N_10240,N_8874,N_6408);
or U10241 (N_10241,N_7404,N_8807);
or U10242 (N_10242,N_6540,N_8362);
and U10243 (N_10243,N_7310,N_6713);
xor U10244 (N_10244,N_7553,N_6544);
xnor U10245 (N_10245,N_8243,N_6630);
nor U10246 (N_10246,N_8850,N_6683);
or U10247 (N_10247,N_8441,N_7328);
or U10248 (N_10248,N_8977,N_9339);
and U10249 (N_10249,N_7871,N_7066);
and U10250 (N_10250,N_8563,N_6658);
xnor U10251 (N_10251,N_8164,N_8479);
nand U10252 (N_10252,N_8610,N_7258);
xnor U10253 (N_10253,N_7109,N_7480);
xnor U10254 (N_10254,N_8513,N_6670);
xnor U10255 (N_10255,N_6417,N_6532);
nor U10256 (N_10256,N_6252,N_6482);
xnor U10257 (N_10257,N_9104,N_6771);
and U10258 (N_10258,N_7063,N_8758);
nor U10259 (N_10259,N_8757,N_7711);
and U10260 (N_10260,N_7484,N_8988);
nor U10261 (N_10261,N_6971,N_7307);
nor U10262 (N_10262,N_7245,N_7143);
nor U10263 (N_10263,N_8901,N_7079);
nor U10264 (N_10264,N_8974,N_8602);
nor U10265 (N_10265,N_8034,N_6854);
xor U10266 (N_10266,N_8334,N_7145);
xor U10267 (N_10267,N_8934,N_7865);
nor U10268 (N_10268,N_6667,N_8536);
and U10269 (N_10269,N_7042,N_7878);
nand U10270 (N_10270,N_8970,N_6718);
nand U10271 (N_10271,N_9018,N_7742);
nand U10272 (N_10272,N_6851,N_8022);
nor U10273 (N_10273,N_8489,N_7364);
xor U10274 (N_10274,N_9108,N_8844);
and U10275 (N_10275,N_8777,N_6772);
nor U10276 (N_10276,N_8795,N_7724);
nand U10277 (N_10277,N_9361,N_8030);
and U10278 (N_10278,N_8116,N_7916);
nor U10279 (N_10279,N_6894,N_6768);
nor U10280 (N_10280,N_6560,N_9081);
nand U10281 (N_10281,N_6785,N_7542);
or U10282 (N_10282,N_7420,N_6502);
xnor U10283 (N_10283,N_7291,N_7686);
nand U10284 (N_10284,N_7004,N_7938);
or U10285 (N_10285,N_7850,N_9354);
nor U10286 (N_10286,N_7289,N_8292);
and U10287 (N_10287,N_6627,N_7735);
and U10288 (N_10288,N_9155,N_8725);
xnor U10289 (N_10289,N_7242,N_8318);
and U10290 (N_10290,N_8346,N_8002);
or U10291 (N_10291,N_8384,N_8448);
or U10292 (N_10292,N_9049,N_9157);
or U10293 (N_10293,N_8287,N_7718);
or U10294 (N_10294,N_8831,N_7357);
nor U10295 (N_10295,N_8512,N_7545);
and U10296 (N_10296,N_8873,N_8940);
nor U10297 (N_10297,N_6688,N_7524);
xor U10298 (N_10298,N_8947,N_7288);
nand U10299 (N_10299,N_8367,N_6738);
nor U10300 (N_10300,N_6825,N_6847);
xor U10301 (N_10301,N_8054,N_8460);
and U10302 (N_10302,N_6585,N_8487);
or U10303 (N_10303,N_7741,N_6584);
or U10304 (N_10304,N_6954,N_8521);
nor U10305 (N_10305,N_8975,N_6306);
and U10306 (N_10306,N_7934,N_7616);
nor U10307 (N_10307,N_6769,N_7286);
nor U10308 (N_10308,N_6342,N_7570);
xor U10309 (N_10309,N_7562,N_7395);
or U10310 (N_10310,N_8817,N_8923);
nand U10311 (N_10311,N_8897,N_7788);
xor U10312 (N_10312,N_8015,N_7777);
nor U10313 (N_10313,N_7712,N_8516);
nand U10314 (N_10314,N_7985,N_7996);
xnor U10315 (N_10315,N_7500,N_6643);
or U10316 (N_10316,N_8859,N_7466);
nor U10317 (N_10317,N_7050,N_7507);
and U10318 (N_10318,N_6365,N_7166);
xor U10319 (N_10319,N_7864,N_6840);
nand U10320 (N_10320,N_8323,N_6340);
and U10321 (N_10321,N_9241,N_8065);
nor U10322 (N_10322,N_7233,N_9070);
xor U10323 (N_10323,N_8863,N_6995);
and U10324 (N_10324,N_8519,N_6747);
or U10325 (N_10325,N_6384,N_6917);
nand U10326 (N_10326,N_7689,N_8471);
and U10327 (N_10327,N_7238,N_9193);
or U10328 (N_10328,N_7334,N_7117);
nor U10329 (N_10329,N_8333,N_8655);
or U10330 (N_10330,N_8364,N_7627);
and U10331 (N_10331,N_6497,N_7284);
or U10332 (N_10332,N_6765,N_7766);
or U10333 (N_10333,N_8247,N_7680);
nand U10334 (N_10334,N_7222,N_9016);
and U10335 (N_10335,N_8612,N_9111);
or U10336 (N_10336,N_9080,N_6903);
or U10337 (N_10337,N_9146,N_8680);
or U10338 (N_10338,N_7720,N_8891);
nand U10339 (N_10339,N_6777,N_8683);
nand U10340 (N_10340,N_7498,N_8202);
nor U10341 (N_10341,N_7371,N_7636);
nand U10342 (N_10342,N_8210,N_8853);
nand U10343 (N_10343,N_7544,N_7344);
nand U10344 (N_10344,N_6907,N_8386);
xor U10345 (N_10345,N_6648,N_6598);
or U10346 (N_10346,N_7485,N_6470);
or U10347 (N_10347,N_8368,N_8687);
or U10348 (N_10348,N_7965,N_6945);
nand U10349 (N_10349,N_8224,N_8965);
and U10350 (N_10350,N_6673,N_8486);
or U10351 (N_10351,N_8056,N_6344);
nor U10352 (N_10352,N_6981,N_9243);
xnor U10353 (N_10353,N_7912,N_6562);
xor U10354 (N_10354,N_7037,N_6574);
nand U10355 (N_10355,N_8964,N_7287);
or U10356 (N_10356,N_6953,N_8525);
nor U10357 (N_10357,N_8021,N_8799);
and U10358 (N_10358,N_8370,N_6315);
xnor U10359 (N_10359,N_9368,N_8783);
or U10360 (N_10360,N_8402,N_7555);
nor U10361 (N_10361,N_6606,N_8678);
or U10362 (N_10362,N_8454,N_9346);
nor U10363 (N_10363,N_9351,N_7324);
or U10364 (N_10364,N_8407,N_7396);
nor U10365 (N_10365,N_7111,N_7678);
or U10366 (N_10366,N_8909,N_6520);
xor U10367 (N_10367,N_7702,N_6305);
and U10368 (N_10368,N_8300,N_8154);
xnor U10369 (N_10369,N_8115,N_7782);
or U10370 (N_10370,N_8495,N_7265);
xor U10371 (N_10371,N_7010,N_7398);
nand U10372 (N_10372,N_6431,N_7807);
xnor U10373 (N_10373,N_6789,N_8549);
xnor U10374 (N_10374,N_6615,N_7048);
and U10375 (N_10375,N_7352,N_7538);
nor U10376 (N_10376,N_6542,N_7967);
nor U10377 (N_10377,N_7027,N_6364);
and U10378 (N_10378,N_6925,N_8717);
and U10379 (N_10379,N_6287,N_9054);
or U10380 (N_10380,N_8630,N_7981);
and U10381 (N_10381,N_7536,N_7360);
or U10382 (N_10382,N_6810,N_9297);
or U10383 (N_10383,N_7675,N_7247);
nand U10384 (N_10384,N_8192,N_8870);
or U10385 (N_10385,N_6616,N_7629);
or U10386 (N_10386,N_8443,N_9105);
or U10387 (N_10387,N_8553,N_7509);
nand U10388 (N_10388,N_8507,N_8268);
nand U10389 (N_10389,N_7331,N_9256);
nand U10390 (N_10390,N_7752,N_6745);
and U10391 (N_10391,N_8613,N_7923);
or U10392 (N_10392,N_6577,N_6815);
nand U10393 (N_10393,N_6960,N_7192);
nand U10394 (N_10394,N_7781,N_9039);
and U10395 (N_10395,N_8972,N_7887);
or U10396 (N_10396,N_8537,N_7572);
xor U10397 (N_10397,N_6547,N_8445);
and U10398 (N_10398,N_7812,N_7338);
and U10399 (N_10399,N_7226,N_6890);
nor U10400 (N_10400,N_6348,N_9195);
and U10401 (N_10401,N_9310,N_7548);
xor U10402 (N_10402,N_8576,N_8102);
or U10403 (N_10403,N_7200,N_9161);
and U10404 (N_10404,N_6456,N_6478);
nand U10405 (N_10405,N_8040,N_8003);
or U10406 (N_10406,N_7298,N_7976);
or U10407 (N_10407,N_7504,N_7644);
or U10408 (N_10408,N_6374,N_9267);
xnor U10409 (N_10409,N_7071,N_7439);
nand U10410 (N_10410,N_8966,N_8872);
or U10411 (N_10411,N_7149,N_7890);
nand U10412 (N_10412,N_6654,N_8149);
nand U10413 (N_10413,N_6519,N_8406);
xnor U10414 (N_10414,N_8332,N_8867);
nand U10415 (N_10415,N_7992,N_7706);
xnor U10416 (N_10416,N_9061,N_7126);
nor U10417 (N_10417,N_8984,N_6435);
nand U10418 (N_10418,N_6427,N_6853);
xor U10419 (N_10419,N_8914,N_8796);
xnor U10420 (N_10420,N_8779,N_7139);
nor U10421 (N_10421,N_8608,N_7786);
or U10422 (N_10422,N_9178,N_8943);
xnor U10423 (N_10423,N_7921,N_9217);
nor U10424 (N_10424,N_6338,N_8433);
xor U10425 (N_10425,N_8746,N_7089);
nand U10426 (N_10426,N_8494,N_7505);
or U10427 (N_10427,N_8677,N_7477);
or U10428 (N_10428,N_7248,N_7653);
xor U10429 (N_10429,N_7793,N_9006);
nor U10430 (N_10430,N_6984,N_8765);
and U10431 (N_10431,N_8463,N_7563);
nand U10432 (N_10432,N_6621,N_7021);
or U10433 (N_10433,N_8743,N_6674);
nand U10434 (N_10434,N_7093,N_6807);
or U10435 (N_10435,N_7745,N_6844);
or U10436 (N_10436,N_8466,N_8604);
xnor U10437 (N_10437,N_8884,N_6836);
or U10438 (N_10438,N_7405,N_7772);
or U10439 (N_10439,N_8646,N_6573);
and U10440 (N_10440,N_6605,N_7413);
or U10441 (N_10441,N_7776,N_7859);
nor U10442 (N_10442,N_6820,N_6291);
or U10443 (N_10443,N_6650,N_8459);
xor U10444 (N_10444,N_6492,N_8089);
nand U10445 (N_10445,N_7160,N_7368);
and U10446 (N_10446,N_6371,N_7227);
and U10447 (N_10447,N_7104,N_7792);
xnor U10448 (N_10448,N_6647,N_9279);
and U10449 (N_10449,N_9101,N_8531);
nand U10450 (N_10450,N_8488,N_9044);
nand U10451 (N_10451,N_7889,N_7469);
and U10452 (N_10452,N_8838,N_9023);
nand U10453 (N_10453,N_8756,N_7140);
or U10454 (N_10454,N_7771,N_9099);
and U10455 (N_10455,N_6481,N_6376);
xor U10456 (N_10456,N_8962,N_8227);
nor U10457 (N_10457,N_8726,N_9017);
nand U10458 (N_10458,N_6472,N_7326);
xor U10459 (N_10459,N_6881,N_8277);
and U10460 (N_10460,N_8651,N_7733);
xnor U10461 (N_10461,N_6719,N_7006);
or U10462 (N_10462,N_7305,N_6914);
or U10463 (N_10463,N_9107,N_6349);
nand U10464 (N_10464,N_7593,N_8276);
nor U10465 (N_10465,N_6866,N_7024);
or U10466 (N_10466,N_9207,N_8810);
nand U10467 (N_10467,N_8237,N_8852);
and U10468 (N_10468,N_9103,N_8442);
or U10469 (N_10469,N_9015,N_7057);
xor U10470 (N_10470,N_8868,N_7393);
or U10471 (N_10471,N_8871,N_8629);
nand U10472 (N_10472,N_8575,N_7124);
and U10473 (N_10473,N_6332,N_8324);
nand U10474 (N_10474,N_6420,N_7765);
and U10475 (N_10475,N_7808,N_7879);
or U10476 (N_10476,N_7151,N_7449);
and U10477 (N_10477,N_8270,N_7127);
and U10478 (N_10478,N_6474,N_7613);
and U10479 (N_10479,N_8514,N_7400);
or U10480 (N_10480,N_8431,N_6422);
nor U10481 (N_10481,N_7450,N_9165);
nand U10482 (N_10482,N_7346,N_8624);
and U10483 (N_10483,N_6770,N_8916);
or U10484 (N_10484,N_8647,N_7246);
xnor U10485 (N_10485,N_6600,N_8860);
nand U10486 (N_10486,N_7679,N_6877);
or U10487 (N_10487,N_8836,N_7699);
nand U10488 (N_10488,N_7935,N_6935);
nand U10489 (N_10489,N_7924,N_8388);
nand U10490 (N_10490,N_8605,N_8957);
xor U10491 (N_10491,N_6878,N_7003);
nand U10492 (N_10492,N_7348,N_8607);
and U10493 (N_10493,N_7353,N_7692);
and U10494 (N_10494,N_7317,N_7892);
and U10495 (N_10495,N_8467,N_8470);
xnor U10496 (N_10496,N_8664,N_7239);
xor U10497 (N_10497,N_8473,N_9223);
nor U10498 (N_10498,N_7827,N_6974);
nor U10499 (N_10499,N_9037,N_6294);
and U10500 (N_10500,N_7835,N_8419);
xnor U10501 (N_10501,N_6316,N_7155);
and U10502 (N_10502,N_7928,N_6405);
nand U10503 (N_10503,N_9264,N_9237);
and U10504 (N_10504,N_8263,N_8670);
or U10505 (N_10505,N_9097,N_8310);
nand U10506 (N_10506,N_6341,N_8979);
xor U10507 (N_10507,N_7666,N_7451);
or U10508 (N_10508,N_7571,N_6552);
and U10509 (N_10509,N_8060,N_9350);
and U10510 (N_10510,N_6932,N_7820);
nor U10511 (N_10511,N_7770,N_6919);
xnor U10512 (N_10512,N_8690,N_7225);
nand U10513 (N_10513,N_8621,N_9252);
and U10514 (N_10514,N_9009,N_8306);
nor U10515 (N_10515,N_6607,N_9011);
xor U10516 (N_10516,N_7837,N_7626);
nor U10517 (N_10517,N_6684,N_6628);
and U10518 (N_10518,N_6430,N_8372);
and U10519 (N_10519,N_7943,N_8729);
nand U10520 (N_10520,N_9320,N_7002);
and U10521 (N_10521,N_6677,N_8280);
and U10522 (N_10522,N_6779,N_6536);
nor U10523 (N_10523,N_7076,N_7565);
nand U10524 (N_10524,N_8976,N_7347);
nand U10525 (N_10525,N_6947,N_8001);
nor U10526 (N_10526,N_7028,N_6499);
nand U10527 (N_10527,N_6457,N_8350);
nand U10528 (N_10528,N_6264,N_9140);
or U10529 (N_10529,N_7234,N_8447);
xnor U10530 (N_10530,N_6846,N_6583);
xor U10531 (N_10531,N_7612,N_8759);
xor U10532 (N_10532,N_8414,N_7463);
xnor U10533 (N_10533,N_7213,N_9068);
and U10534 (N_10534,N_8360,N_7917);
and U10535 (N_10535,N_6461,N_6504);
or U10536 (N_10536,N_9198,N_7170);
and U10537 (N_10537,N_7573,N_8633);
nand U10538 (N_10538,N_9202,N_8163);
and U10539 (N_10539,N_6381,N_6313);
xnor U10540 (N_10540,N_8365,N_8997);
nor U10541 (N_10541,N_6905,N_9078);
and U10542 (N_10542,N_7775,N_8104);
xor U10543 (N_10543,N_6444,N_8781);
xor U10544 (N_10544,N_8527,N_8341);
and U10545 (N_10545,N_8371,N_7336);
or U10546 (N_10546,N_8695,N_9333);
and U10547 (N_10547,N_6827,N_6288);
or U10548 (N_10548,N_7634,N_7051);
nor U10549 (N_10549,N_8806,N_9204);
nand U10550 (N_10550,N_8809,N_7658);
or U10551 (N_10551,N_7830,N_6406);
and U10552 (N_10552,N_6476,N_6832);
and U10553 (N_10553,N_8574,N_6522);
and U10554 (N_10554,N_8805,N_6528);
or U10555 (N_10555,N_7550,N_7207);
nor U10556 (N_10556,N_8155,N_7883);
or U10557 (N_10557,N_8682,N_8504);
nand U10558 (N_10558,N_7541,N_8219);
xnor U10559 (N_10559,N_7264,N_7705);
nor U10560 (N_10560,N_7886,N_7375);
xnor U10561 (N_10561,N_8126,N_7013);
xnor U10562 (N_10562,N_8204,N_6845);
or U10563 (N_10563,N_8733,N_8176);
nand U10564 (N_10564,N_8458,N_6468);
nor U10565 (N_10565,N_8093,N_8526);
nand U10566 (N_10566,N_7088,N_9067);
nand U10567 (N_10567,N_8755,N_7085);
nor U10568 (N_10568,N_8722,N_8175);
nand U10569 (N_10569,N_7564,N_8910);
nor U10570 (N_10570,N_6311,N_6996);
nand U10571 (N_10571,N_7691,N_6530);
nand U10572 (N_10572,N_8190,N_8113);
xor U10573 (N_10573,N_8675,N_6687);
nand U10574 (N_10574,N_8416,N_9040);
xor U10575 (N_10575,N_7621,N_7096);
or U10576 (N_10576,N_6603,N_8693);
and U10577 (N_10577,N_7370,N_8179);
nand U10578 (N_10578,N_7012,N_8557);
or U10579 (N_10579,N_8705,N_8374);
and U10580 (N_10580,N_8068,N_7910);
and U10581 (N_10581,N_7325,N_6493);
nor U10582 (N_10582,N_6345,N_6533);
or U10583 (N_10583,N_6509,N_8689);
nor U10584 (N_10584,N_9074,N_6425);
nand U10585 (N_10585,N_8395,N_9087);
nor U10586 (N_10586,N_9214,N_9065);
nand U10587 (N_10587,N_6993,N_8861);
or U10588 (N_10588,N_8273,N_7637);
nor U10589 (N_10589,N_6378,N_6804);
nor U10590 (N_10590,N_6441,N_6388);
and U10591 (N_10591,N_8620,N_6940);
or U10592 (N_10592,N_8330,N_7586);
xnor U10593 (N_10593,N_7595,N_7019);
or U10594 (N_10594,N_7953,N_7877);
or U10595 (N_10595,N_7868,N_6631);
xnor U10596 (N_10596,N_7569,N_8639);
nor U10597 (N_10597,N_7561,N_8706);
nor U10598 (N_10598,N_7110,N_7435);
and U10599 (N_10599,N_7116,N_7120);
or U10600 (N_10600,N_7281,N_6568);
nand U10601 (N_10601,N_8230,N_7443);
nor U10602 (N_10602,N_8782,N_8627);
and U10603 (N_10603,N_9090,N_6495);
nor U10604 (N_10604,N_8199,N_7390);
and U10605 (N_10605,N_8231,N_8698);
or U10606 (N_10606,N_7044,N_9255);
nor U10607 (N_10607,N_8841,N_7150);
xor U10608 (N_10608,N_6875,N_7252);
nor U10609 (N_10609,N_7293,N_8285);
and U10610 (N_10610,N_7748,N_7502);
xor U10611 (N_10611,N_8595,N_7822);
xor U10612 (N_10612,N_7442,N_8044);
or U10613 (N_10613,N_6439,N_6537);
and U10614 (N_10614,N_7169,N_8641);
nor U10615 (N_10615,N_8540,N_7696);
or U10616 (N_10616,N_9022,N_8006);
or U10617 (N_10617,N_7695,N_8452);
nor U10618 (N_10618,N_8069,N_8036);
and U10619 (N_10619,N_7622,N_8835);
and U10620 (N_10620,N_6545,N_8902);
nand U10621 (N_10621,N_9257,N_6523);
nor U10622 (N_10622,N_7419,N_8720);
or U10623 (N_10623,N_8774,N_7529);
nor U10624 (N_10624,N_7520,N_6795);
or U10625 (N_10625,N_9112,N_8590);
nor U10626 (N_10626,N_8253,N_7062);
and U10627 (N_10627,N_6834,N_7880);
or U10628 (N_10628,N_8785,N_8644);
or U10629 (N_10629,N_9277,N_6740);
nand U10630 (N_10630,N_8699,N_9309);
xnor U10631 (N_10631,N_7843,N_6391);
and U10632 (N_10632,N_8735,N_6571);
and U10633 (N_10633,N_8559,N_9266);
nor U10634 (N_10634,N_9033,N_8361);
or U10635 (N_10635,N_6961,N_7332);
and U10636 (N_10636,N_7361,N_7292);
xor U10637 (N_10637,N_9075,N_6442);
nand U10638 (N_10638,N_9131,N_7645);
and U10639 (N_10639,N_7301,N_9013);
nor U10640 (N_10640,N_7579,N_8565);
nor U10641 (N_10641,N_6466,N_8244);
and U10642 (N_10642,N_7755,N_7379);
nor U10643 (N_10643,N_9280,N_9181);
or U10644 (N_10644,N_6434,N_9137);
nor U10645 (N_10645,N_7651,N_6352);
nor U10646 (N_10646,N_7790,N_9073);
or U10647 (N_10647,N_8709,N_9188);
or U10648 (N_10648,N_9171,N_6707);
or U10649 (N_10649,N_8711,N_8740);
and U10650 (N_10650,N_7373,N_7980);
nor U10651 (N_10651,N_8955,N_9359);
or U10652 (N_10652,N_8298,N_6873);
xnor U10653 (N_10653,N_8978,N_8385);
and U10654 (N_10654,N_9340,N_9177);
nand U10655 (N_10655,N_6359,N_6353);
or U10656 (N_10656,N_8456,N_6258);
xnor U10657 (N_10657,N_6826,N_7551);
nor U10658 (N_10658,N_6829,N_7251);
and U10659 (N_10659,N_7482,N_7098);
nor U10660 (N_10660,N_9300,N_8157);
and U10661 (N_10661,N_8301,N_7926);
or U10662 (N_10662,N_8208,N_6798);
xor U10663 (N_10663,N_9329,N_9308);
or U10664 (N_10664,N_6454,N_6524);
nand U10665 (N_10665,N_7077,N_7763);
or U10666 (N_10666,N_7655,N_8961);
or U10667 (N_10667,N_8379,N_6591);
and U10668 (N_10668,N_8658,N_6861);
and U10669 (N_10669,N_8238,N_8896);
xor U10670 (N_10670,N_8437,N_6299);
nor U10671 (N_10671,N_8450,N_8556);
and U10672 (N_10672,N_8971,N_6865);
nand U10673 (N_10673,N_7040,N_8245);
or U10674 (N_10674,N_8710,N_7797);
nand U10675 (N_10675,N_6334,N_8622);
nor U10676 (N_10676,N_9220,N_8200);
nor U10677 (N_10677,N_7359,N_7834);
nor U10678 (N_10678,N_8547,N_7115);
or U10679 (N_10679,N_7506,N_8520);
or U10680 (N_10680,N_8503,N_7823);
xor U10681 (N_10681,N_7391,N_7197);
or U10682 (N_10682,N_8028,N_9143);
and U10683 (N_10683,N_9224,N_9093);
nand U10684 (N_10684,N_8554,N_8517);
or U10685 (N_10685,N_9123,N_9369);
or U10686 (N_10686,N_6290,N_8530);
nand U10687 (N_10687,N_9038,N_8941);
or U10688 (N_10688,N_6567,N_7156);
or U10689 (N_10689,N_7799,N_7697);
and U10690 (N_10690,N_7540,N_8688);
nor U10691 (N_10691,N_6754,N_9298);
nand U10692 (N_10692,N_6505,N_8894);
and U10693 (N_10693,N_8712,N_8566);
and U10694 (N_10694,N_7316,N_7816);
or U10695 (N_10695,N_7798,N_6910);
xor U10696 (N_10696,N_8008,N_8787);
and U10697 (N_10697,N_7113,N_7749);
and U10698 (N_10698,N_7870,N_9139);
and U10699 (N_10699,N_8599,N_6691);
or U10700 (N_10700,N_7683,N_8833);
xnor U10701 (N_10701,N_9262,N_6541);
nand U10702 (N_10702,N_8409,N_8648);
and U10703 (N_10703,N_8326,N_9084);
xor U10704 (N_10704,N_8825,N_7811);
and U10705 (N_10705,N_8701,N_9332);
xnor U10706 (N_10706,N_7746,N_7898);
nor U10707 (N_10707,N_7374,N_7059);
and U10708 (N_10708,N_7159,N_7270);
or U10709 (N_10709,N_8029,N_7476);
and U10710 (N_10710,N_9144,N_7183);
nand U10711 (N_10711,N_6415,N_8110);
nor U10712 (N_10712,N_6986,N_7275);
nand U10713 (N_10713,N_8193,N_6726);
and U10714 (N_10714,N_8241,N_8048);
or U10715 (N_10715,N_6274,N_7927);
and U10716 (N_10716,N_6402,N_7102);
nand U10717 (N_10717,N_8653,N_6892);
xor U10718 (N_10718,N_7665,N_7750);
and U10719 (N_10719,N_6620,N_8801);
nand U10720 (N_10720,N_8123,N_7303);
or U10721 (N_10721,N_8100,N_7483);
and U10722 (N_10722,N_9042,N_7582);
or U10723 (N_10723,N_8842,N_6634);
and U10724 (N_10724,N_6377,N_8732);
xnor U10725 (N_10725,N_8344,N_9347);
nand U10726 (N_10726,N_7978,N_7851);
xor U10727 (N_10727,N_6741,N_7614);
nand U10728 (N_10728,N_6464,N_8296);
and U10729 (N_10729,N_6712,N_6823);
and U10730 (N_10730,N_6716,N_7492);
nor U10731 (N_10731,N_7053,N_9110);
or U10732 (N_10732,N_8707,N_8075);
xnor U10733 (N_10733,N_8418,N_6445);
xor U10734 (N_10734,N_8059,N_9215);
nor U10735 (N_10735,N_8462,N_8770);
nand U10736 (N_10736,N_8734,N_7977);
nand U10737 (N_10737,N_6811,N_9076);
nor U10738 (N_10738,N_7885,N_7273);
and U10739 (N_10739,N_7171,N_7464);
or U10740 (N_10740,N_6539,N_7153);
xor U10741 (N_10741,N_7377,N_9159);
or U10742 (N_10742,N_8257,N_9283);
xor U10743 (N_10743,N_6443,N_8523);
and U10744 (N_10744,N_7840,N_6644);
and U10745 (N_10745,N_8143,N_6934);
and U10746 (N_10746,N_8558,N_9169);
or U10747 (N_10747,N_6786,N_6317);
nor U10748 (N_10748,N_7635,N_8745);
xor U10749 (N_10749,N_6263,N_7738);
and U10750 (N_10750,N_7704,N_6462);
and U10751 (N_10751,N_9253,N_9187);
nor U10752 (N_10752,N_8636,N_8320);
nor U10753 (N_10753,N_8139,N_8791);
nand U10754 (N_10754,N_7942,N_8650);
or U10755 (N_10755,N_7422,N_6386);
xnor U10756 (N_10756,N_9058,N_8439);
and U10757 (N_10757,N_9210,N_6927);
or U10758 (N_10758,N_8749,N_7973);
and U10759 (N_10759,N_9203,N_7625);
xnor U10760 (N_10760,N_7082,N_7411);
nor U10761 (N_10761,N_7119,N_6617);
xor U10762 (N_10762,N_8092,N_8506);
nor U10763 (N_10763,N_7272,N_8908);
nor U10764 (N_10764,N_8843,N_7828);
and U10765 (N_10765,N_9357,N_6920);
nor U10766 (N_10766,N_6852,N_8428);
xor U10767 (N_10767,N_9162,N_9109);
or U10768 (N_10768,N_8606,N_8165);
and U10769 (N_10769,N_7638,N_9206);
and U10770 (N_10770,N_9138,N_8218);
nor U10771 (N_10771,N_8023,N_8829);
xor U10772 (N_10772,N_9083,N_7203);
xor U10773 (N_10773,N_8480,N_6916);
nand U10774 (N_10774,N_8391,N_9344);
xor U10775 (N_10775,N_9007,N_8469);
or U10776 (N_10776,N_6891,N_7425);
and U10777 (N_10777,N_6253,N_9158);
nand U10778 (N_10778,N_8887,N_8584);
nor U10779 (N_10779,N_8369,N_8500);
xor U10780 (N_10780,N_7428,N_6714);
nor U10781 (N_10781,N_7826,N_6734);
nand U10782 (N_10782,N_9234,N_8206);
or U10783 (N_10783,N_6952,N_9226);
nand U10784 (N_10784,N_8539,N_8617);
xor U10785 (N_10785,N_7188,N_6682);
or U10786 (N_10786,N_8172,N_6685);
and U10787 (N_10787,N_7407,N_6566);
xnor U10788 (N_10788,N_6904,N_8635);
nor U10789 (N_10789,N_8601,N_8603);
nor U10790 (N_10790,N_8327,N_9319);
or U10791 (N_10791,N_7946,N_6908);
or U10792 (N_10792,N_6589,N_8982);
or U10793 (N_10793,N_8713,N_7386);
or U10794 (N_10794,N_7438,N_6624);
and U10795 (N_10795,N_8169,N_8811);
or U10796 (N_10796,N_8551,N_8583);
xor U10797 (N_10797,N_8893,N_7033);
and U10798 (N_10798,N_7092,N_8403);
and U10799 (N_10799,N_8465,N_9258);
xor U10800 (N_10800,N_6806,N_6280);
or U10801 (N_10801,N_7604,N_7296);
nand U10802 (N_10802,N_7918,N_7762);
nand U10803 (N_10803,N_7433,N_7836);
or U10804 (N_10804,N_7737,N_8019);
and U10805 (N_10805,N_8820,N_8383);
and U10806 (N_10806,N_8865,N_8217);
and U10807 (N_10807,N_8944,N_7716);
nor U10808 (N_10808,N_8714,N_7744);
nand U10809 (N_10809,N_6838,N_6898);
xnor U10810 (N_10810,N_7605,N_6302);
nor U10811 (N_10811,N_7940,N_7184);
nor U10812 (N_10812,N_8187,N_7255);
and U10813 (N_10813,N_6490,N_7446);
nand U10814 (N_10814,N_7707,N_7945);
or U10815 (N_10815,N_6657,N_7600);
nor U10816 (N_10816,N_7190,N_6708);
and U10817 (N_10817,N_8490,N_6989);
xor U10818 (N_10818,N_6668,N_6250);
nor U10819 (N_10819,N_9117,N_7097);
and U10820 (N_10820,N_6801,N_8265);
and U10821 (N_10821,N_6689,N_8073);
xor U10822 (N_10822,N_6753,N_7585);
or U10823 (N_10823,N_7929,N_7372);
xor U10824 (N_10824,N_6639,N_8337);
and U10825 (N_10825,N_9311,N_8189);
nand U10826 (N_10826,N_8203,N_9004);
and U10827 (N_10827,N_6931,N_6370);
and U10828 (N_10828,N_6976,N_8753);
or U10829 (N_10829,N_7957,N_6614);
nand U10830 (N_10830,N_7017,N_6428);
or U10831 (N_10831,N_6762,N_7488);
or U10832 (N_10832,N_7095,N_7988);
nand U10833 (N_10833,N_7677,N_9229);
nor U10834 (N_10834,N_8229,N_7431);
and U10835 (N_10835,N_6912,N_9121);
nor U10836 (N_10836,N_6656,N_6783);
nor U10837 (N_10837,N_7041,N_6900);
nor U10838 (N_10838,N_7966,N_6946);
xnor U10839 (N_10839,N_6678,N_6715);
or U10840 (N_10840,N_6578,N_8446);
or U10841 (N_10841,N_6706,N_6475);
or U10842 (N_10842,N_6484,N_7221);
nand U10843 (N_10843,N_8464,N_6581);
or U10844 (N_10844,N_6488,N_9045);
nand U10845 (N_10845,N_7856,N_9114);
or U10846 (N_10846,N_8125,N_7800);
nor U10847 (N_10847,N_9293,N_6489);
nand U10848 (N_10848,N_8945,N_7349);
nand U10849 (N_10849,N_6595,N_7409);
and U10850 (N_10850,N_6862,N_6418);
nand U10851 (N_10851,N_7568,N_7815);
and U10852 (N_10852,N_7989,N_8427);
or U10853 (N_10853,N_6918,N_9136);
xor U10854 (N_10854,N_6279,N_9113);
or U10855 (N_10855,N_8440,N_8905);
xor U10856 (N_10856,N_8196,N_6666);
nor U10857 (N_10857,N_6979,N_8771);
nand U10858 (N_10858,N_6534,N_6452);
nor U10859 (N_10859,N_8499,N_6929);
xnor U10860 (N_10860,N_6817,N_7933);
nand U10861 (N_10861,N_6857,N_7952);
xor U10862 (N_10862,N_6744,N_8186);
nand U10863 (N_10863,N_8234,N_9238);
or U10864 (N_10864,N_7508,N_8161);
and U10865 (N_10865,N_8248,N_8412);
xor U10866 (N_10866,N_7983,N_7594);
and U10867 (N_10867,N_8813,N_9209);
xor U10868 (N_10868,N_6736,N_9014);
nand U10869 (N_10869,N_8983,N_6824);
nor U10870 (N_10870,N_9057,N_6982);
and U10871 (N_10871,N_6270,N_6749);
nor U10872 (N_10872,N_7700,N_8242);
or U10873 (N_10873,N_8376,N_9059);
xor U10874 (N_10874,N_7703,N_7873);
nand U10875 (N_10875,N_7761,N_6969);
or U10876 (N_10876,N_9358,N_6559);
nor U10877 (N_10877,N_6773,N_8085);
and U10878 (N_10878,N_8024,N_9285);
nand U10879 (N_10879,N_7253,N_7649);
nand U10880 (N_10880,N_7376,N_8136);
and U10881 (N_10881,N_8913,N_8138);
nand U10882 (N_10882,N_6613,N_7673);
and U10883 (N_10883,N_7285,N_7962);
and U10884 (N_10884,N_8184,N_8925);
xnor U10885 (N_10885,N_6458,N_7215);
xnor U10886 (N_10886,N_9240,N_7794);
or U10887 (N_10887,N_6593,N_8127);
xor U10888 (N_10888,N_6697,N_9275);
or U10889 (N_10889,N_7394,N_8411);
or U10890 (N_10890,N_8312,N_8614);
and U10891 (N_10891,N_6572,N_8950);
nor U10892 (N_10892,N_7897,N_8167);
nand U10893 (N_10893,N_7900,N_9173);
xor U10894 (N_10894,N_8518,N_7861);
nor U10895 (N_10895,N_7154,N_8063);
xnor U10896 (N_10896,N_6973,N_7728);
or U10897 (N_10897,N_8888,N_6467);
or U10898 (N_10898,N_8544,N_9218);
and U10899 (N_10899,N_7532,N_7432);
nand U10900 (N_10900,N_6637,N_8303);
xnor U10901 (N_10901,N_6432,N_8145);
xor U10902 (N_10902,N_9092,N_8201);
xor U10903 (N_10903,N_7065,N_9251);
nand U10904 (N_10904,N_9205,N_6962);
nand U10905 (N_10905,N_8739,N_8989);
nand U10906 (N_10906,N_7654,N_8322);
nand U10907 (N_10907,N_7214,N_7591);
or U10908 (N_10908,N_9330,N_8039);
nor U10909 (N_10909,N_8985,N_7603);
xnor U10910 (N_10910,N_6292,N_7486);
nand U10911 (N_10911,N_7907,N_8895);
xnor U10912 (N_10912,N_7664,N_8038);
and U10913 (N_10913,N_6336,N_7631);
xnor U10914 (N_10914,N_8216,N_8618);
nor U10915 (N_10915,N_7860,N_8336);
or U10916 (N_10916,N_7009,N_8994);
nor U10917 (N_10917,N_8593,N_8258);
and U10918 (N_10918,N_6339,N_7817);
or U10919 (N_10919,N_6412,N_9077);
nor U10920 (N_10920,N_8681,N_7964);
xor U10921 (N_10921,N_6814,N_8657);
nor U10922 (N_10922,N_6498,N_7574);
nand U10923 (N_10923,N_8768,N_7853);
nor U10924 (N_10924,N_6842,N_6266);
or U10925 (N_10925,N_8990,N_8594);
nor U10926 (N_10926,N_7846,N_7577);
and U10927 (N_10927,N_7813,N_8047);
or U10928 (N_10928,N_8086,N_8704);
nand U10929 (N_10929,N_7516,N_8225);
and U10930 (N_10930,N_7217,N_6351);
xor U10931 (N_10931,N_6429,N_8064);
or U10932 (N_10932,N_7261,N_6387);
and U10933 (N_10933,N_6366,N_6450);
nand U10934 (N_10934,N_8578,N_6437);
xor U10935 (N_10935,N_8183,N_7714);
or U10936 (N_10936,N_8642,N_7299);
and U10937 (N_10937,N_7674,N_9003);
and U10938 (N_10938,N_7465,N_8111);
xnor U10939 (N_10939,N_7192,N_8736);
xnor U10940 (N_10940,N_6414,N_6548);
or U10941 (N_10941,N_8936,N_9074);
nor U10942 (N_10942,N_7931,N_8986);
nor U10943 (N_10943,N_6615,N_7925);
or U10944 (N_10944,N_6364,N_6840);
nand U10945 (N_10945,N_7736,N_8273);
nor U10946 (N_10946,N_6765,N_7982);
nand U10947 (N_10947,N_8218,N_6640);
nand U10948 (N_10948,N_8019,N_9155);
nor U10949 (N_10949,N_7650,N_6804);
and U10950 (N_10950,N_7102,N_7199);
nand U10951 (N_10951,N_7814,N_7576);
nor U10952 (N_10952,N_8835,N_8245);
and U10953 (N_10953,N_8147,N_6637);
nand U10954 (N_10954,N_8131,N_7569);
and U10955 (N_10955,N_9021,N_8155);
or U10956 (N_10956,N_8705,N_6616);
nand U10957 (N_10957,N_7517,N_7967);
xnor U10958 (N_10958,N_6311,N_6493);
and U10959 (N_10959,N_8764,N_6481);
xor U10960 (N_10960,N_8363,N_8975);
xor U10961 (N_10961,N_9367,N_7528);
nor U10962 (N_10962,N_8263,N_9106);
nand U10963 (N_10963,N_6863,N_7286);
nor U10964 (N_10964,N_8231,N_8949);
and U10965 (N_10965,N_7241,N_7027);
nand U10966 (N_10966,N_7516,N_6822);
nand U10967 (N_10967,N_8956,N_9321);
xnor U10968 (N_10968,N_6799,N_6746);
or U10969 (N_10969,N_7692,N_9236);
nand U10970 (N_10970,N_6313,N_6871);
nand U10971 (N_10971,N_8590,N_9276);
nand U10972 (N_10972,N_7698,N_6459);
nand U10973 (N_10973,N_6622,N_9326);
or U10974 (N_10974,N_6814,N_6910);
or U10975 (N_10975,N_9159,N_7884);
xor U10976 (N_10976,N_7884,N_7767);
or U10977 (N_10977,N_9210,N_9061);
nand U10978 (N_10978,N_7628,N_8043);
or U10979 (N_10979,N_7148,N_9266);
nor U10980 (N_10980,N_9126,N_6804);
nor U10981 (N_10981,N_7621,N_7585);
xor U10982 (N_10982,N_9284,N_7768);
and U10983 (N_10983,N_7797,N_6844);
nand U10984 (N_10984,N_8846,N_7085);
xnor U10985 (N_10985,N_8368,N_8607);
xnor U10986 (N_10986,N_7160,N_7150);
or U10987 (N_10987,N_6580,N_9280);
or U10988 (N_10988,N_6939,N_8333);
xor U10989 (N_10989,N_7796,N_6737);
xor U10990 (N_10990,N_8810,N_6579);
or U10991 (N_10991,N_7454,N_7962);
nor U10992 (N_10992,N_7544,N_8184);
and U10993 (N_10993,N_9262,N_9170);
nor U10994 (N_10994,N_7421,N_7637);
and U10995 (N_10995,N_9212,N_6955);
and U10996 (N_10996,N_6602,N_7176);
nor U10997 (N_10997,N_9147,N_7180);
nor U10998 (N_10998,N_8688,N_7608);
nor U10999 (N_10999,N_7120,N_6319);
nand U11000 (N_11000,N_9184,N_8251);
nor U11001 (N_11001,N_6580,N_9351);
or U11002 (N_11002,N_7888,N_6719);
xor U11003 (N_11003,N_6689,N_8728);
nor U11004 (N_11004,N_7213,N_7543);
and U11005 (N_11005,N_6949,N_7222);
or U11006 (N_11006,N_6926,N_8771);
or U11007 (N_11007,N_8553,N_9290);
and U11008 (N_11008,N_8626,N_8629);
and U11009 (N_11009,N_9308,N_7263);
and U11010 (N_11010,N_7666,N_8059);
or U11011 (N_11011,N_8621,N_8964);
nand U11012 (N_11012,N_9210,N_6437);
nand U11013 (N_11013,N_7174,N_6524);
or U11014 (N_11014,N_6436,N_9173);
xor U11015 (N_11015,N_6964,N_7364);
and U11016 (N_11016,N_6517,N_7903);
nand U11017 (N_11017,N_7976,N_7558);
nor U11018 (N_11018,N_8555,N_9299);
and U11019 (N_11019,N_9296,N_8957);
and U11020 (N_11020,N_8735,N_6300);
nand U11021 (N_11021,N_9200,N_6722);
and U11022 (N_11022,N_7887,N_7500);
nor U11023 (N_11023,N_6490,N_8812);
and U11024 (N_11024,N_9286,N_7329);
and U11025 (N_11025,N_7154,N_7493);
nor U11026 (N_11026,N_6975,N_9332);
and U11027 (N_11027,N_6296,N_7469);
nand U11028 (N_11028,N_8692,N_6718);
nand U11029 (N_11029,N_7570,N_6473);
nand U11030 (N_11030,N_8466,N_8955);
nand U11031 (N_11031,N_8695,N_7333);
xnor U11032 (N_11032,N_8598,N_7773);
nor U11033 (N_11033,N_6254,N_7652);
nor U11034 (N_11034,N_6427,N_8261);
nor U11035 (N_11035,N_8623,N_6496);
or U11036 (N_11036,N_9179,N_8369);
or U11037 (N_11037,N_7498,N_6425);
and U11038 (N_11038,N_7615,N_7029);
nor U11039 (N_11039,N_7110,N_9223);
and U11040 (N_11040,N_6761,N_7445);
xnor U11041 (N_11041,N_7831,N_6809);
nand U11042 (N_11042,N_8906,N_6689);
xnor U11043 (N_11043,N_6601,N_7403);
or U11044 (N_11044,N_8168,N_7113);
or U11045 (N_11045,N_6475,N_7970);
or U11046 (N_11046,N_8612,N_6988);
nor U11047 (N_11047,N_6714,N_8952);
nand U11048 (N_11048,N_7749,N_8713);
and U11049 (N_11049,N_6990,N_6365);
xor U11050 (N_11050,N_8739,N_7081);
nor U11051 (N_11051,N_7002,N_7227);
or U11052 (N_11052,N_9124,N_8715);
nor U11053 (N_11053,N_8157,N_7485);
xor U11054 (N_11054,N_7893,N_6675);
and U11055 (N_11055,N_7144,N_6263);
nor U11056 (N_11056,N_7756,N_7184);
nor U11057 (N_11057,N_7212,N_8331);
nor U11058 (N_11058,N_7401,N_7851);
xor U11059 (N_11059,N_8309,N_8809);
or U11060 (N_11060,N_6935,N_8740);
nand U11061 (N_11061,N_9171,N_8293);
nor U11062 (N_11062,N_8732,N_8610);
nor U11063 (N_11063,N_8894,N_8859);
and U11064 (N_11064,N_7194,N_6511);
and U11065 (N_11065,N_8633,N_9347);
xor U11066 (N_11066,N_8512,N_8088);
xor U11067 (N_11067,N_6959,N_7459);
or U11068 (N_11068,N_7671,N_6674);
nor U11069 (N_11069,N_7893,N_9100);
nor U11070 (N_11070,N_7372,N_9193);
xor U11071 (N_11071,N_7532,N_7625);
or U11072 (N_11072,N_7995,N_7119);
and U11073 (N_11073,N_8977,N_7655);
nand U11074 (N_11074,N_8318,N_6892);
xor U11075 (N_11075,N_8900,N_7685);
or U11076 (N_11076,N_6820,N_8636);
xnor U11077 (N_11077,N_6932,N_9034);
xnor U11078 (N_11078,N_9354,N_8292);
nor U11079 (N_11079,N_6473,N_7536);
nand U11080 (N_11080,N_6801,N_6851);
or U11081 (N_11081,N_8020,N_7725);
or U11082 (N_11082,N_7676,N_8212);
nor U11083 (N_11083,N_8426,N_8760);
nor U11084 (N_11084,N_8850,N_8828);
xnor U11085 (N_11085,N_8020,N_8315);
xnor U11086 (N_11086,N_9350,N_7657);
or U11087 (N_11087,N_9315,N_6539);
or U11088 (N_11088,N_7669,N_9088);
nand U11089 (N_11089,N_7677,N_8026);
xnor U11090 (N_11090,N_8274,N_7946);
or U11091 (N_11091,N_9148,N_9292);
or U11092 (N_11092,N_6522,N_7610);
and U11093 (N_11093,N_6840,N_9056);
nand U11094 (N_11094,N_8158,N_7018);
xnor U11095 (N_11095,N_6846,N_8415);
nor U11096 (N_11096,N_9304,N_8527);
nor U11097 (N_11097,N_6545,N_9079);
nor U11098 (N_11098,N_8978,N_8185);
or U11099 (N_11099,N_8174,N_6524);
and U11100 (N_11100,N_7648,N_7571);
xor U11101 (N_11101,N_8165,N_7086);
xnor U11102 (N_11102,N_6431,N_6812);
or U11103 (N_11103,N_7812,N_7933);
or U11104 (N_11104,N_8489,N_8962);
or U11105 (N_11105,N_9040,N_8262);
nand U11106 (N_11106,N_8773,N_7954);
nand U11107 (N_11107,N_9290,N_6343);
and U11108 (N_11108,N_8451,N_8774);
xor U11109 (N_11109,N_6871,N_8320);
xnor U11110 (N_11110,N_7408,N_9162);
xnor U11111 (N_11111,N_7336,N_6708);
nand U11112 (N_11112,N_7764,N_6380);
nand U11113 (N_11113,N_9029,N_8791);
nor U11114 (N_11114,N_7453,N_6969);
or U11115 (N_11115,N_8448,N_9029);
nor U11116 (N_11116,N_7667,N_6853);
xor U11117 (N_11117,N_7341,N_8248);
xnor U11118 (N_11118,N_6789,N_6375);
nand U11119 (N_11119,N_7631,N_6279);
nand U11120 (N_11120,N_7231,N_6335);
nand U11121 (N_11121,N_8012,N_8127);
xnor U11122 (N_11122,N_9002,N_8402);
xnor U11123 (N_11123,N_6924,N_6548);
or U11124 (N_11124,N_7356,N_7904);
xor U11125 (N_11125,N_8359,N_7108);
and U11126 (N_11126,N_8270,N_8405);
and U11127 (N_11127,N_7448,N_8652);
and U11128 (N_11128,N_7985,N_6483);
or U11129 (N_11129,N_8855,N_8490);
xor U11130 (N_11130,N_8793,N_8872);
and U11131 (N_11131,N_7469,N_9181);
and U11132 (N_11132,N_9249,N_6576);
nor U11133 (N_11133,N_8114,N_7681);
xor U11134 (N_11134,N_6820,N_8430);
xnor U11135 (N_11135,N_7212,N_8796);
nor U11136 (N_11136,N_6363,N_7687);
and U11137 (N_11137,N_8730,N_9050);
and U11138 (N_11138,N_6578,N_9255);
nor U11139 (N_11139,N_8686,N_8094);
nor U11140 (N_11140,N_7295,N_7896);
or U11141 (N_11141,N_7697,N_8161);
and U11142 (N_11142,N_7569,N_6473);
and U11143 (N_11143,N_7495,N_8047);
or U11144 (N_11144,N_7841,N_6810);
and U11145 (N_11145,N_8799,N_7269);
xnor U11146 (N_11146,N_9007,N_8250);
and U11147 (N_11147,N_8063,N_7745);
and U11148 (N_11148,N_6761,N_8363);
and U11149 (N_11149,N_9102,N_8532);
and U11150 (N_11150,N_8848,N_7595);
or U11151 (N_11151,N_7959,N_8206);
and U11152 (N_11152,N_6323,N_7363);
and U11153 (N_11153,N_8706,N_7415);
or U11154 (N_11154,N_8084,N_8046);
and U11155 (N_11155,N_8193,N_7220);
xnor U11156 (N_11156,N_7143,N_7792);
nor U11157 (N_11157,N_8168,N_6657);
and U11158 (N_11158,N_8127,N_8016);
or U11159 (N_11159,N_8045,N_8038);
nand U11160 (N_11160,N_7195,N_6531);
nor U11161 (N_11161,N_9154,N_9151);
or U11162 (N_11162,N_7133,N_7886);
or U11163 (N_11163,N_8985,N_8477);
nand U11164 (N_11164,N_7905,N_8523);
xnor U11165 (N_11165,N_6933,N_6795);
nand U11166 (N_11166,N_8897,N_7223);
nor U11167 (N_11167,N_8418,N_7597);
nor U11168 (N_11168,N_8805,N_8357);
nor U11169 (N_11169,N_8896,N_8194);
nand U11170 (N_11170,N_8241,N_7129);
nand U11171 (N_11171,N_6704,N_6829);
nand U11172 (N_11172,N_8414,N_8286);
and U11173 (N_11173,N_7312,N_8893);
nor U11174 (N_11174,N_7054,N_9273);
or U11175 (N_11175,N_7214,N_9356);
nand U11176 (N_11176,N_6765,N_8154);
xnor U11177 (N_11177,N_6697,N_7459);
or U11178 (N_11178,N_7388,N_8837);
and U11179 (N_11179,N_6613,N_8580);
and U11180 (N_11180,N_9201,N_6987);
and U11181 (N_11181,N_8838,N_6655);
and U11182 (N_11182,N_8165,N_7883);
xnor U11183 (N_11183,N_8136,N_8901);
nand U11184 (N_11184,N_8774,N_6511);
nor U11185 (N_11185,N_8829,N_7598);
xnor U11186 (N_11186,N_6678,N_7340);
nand U11187 (N_11187,N_6715,N_9096);
nand U11188 (N_11188,N_6739,N_8040);
nand U11189 (N_11189,N_6505,N_9264);
or U11190 (N_11190,N_6364,N_8751);
or U11191 (N_11191,N_6553,N_8366);
nand U11192 (N_11192,N_8386,N_9071);
or U11193 (N_11193,N_9030,N_8543);
nor U11194 (N_11194,N_7826,N_8904);
xnor U11195 (N_11195,N_7949,N_8131);
xor U11196 (N_11196,N_6370,N_7695);
xor U11197 (N_11197,N_8339,N_7010);
or U11198 (N_11198,N_6527,N_6717);
nand U11199 (N_11199,N_7008,N_7051);
or U11200 (N_11200,N_8708,N_6922);
nor U11201 (N_11201,N_8829,N_8523);
or U11202 (N_11202,N_6849,N_7299);
or U11203 (N_11203,N_8985,N_7478);
nand U11204 (N_11204,N_8520,N_7968);
and U11205 (N_11205,N_9215,N_6324);
xor U11206 (N_11206,N_7804,N_7377);
nand U11207 (N_11207,N_8766,N_7647);
and U11208 (N_11208,N_8628,N_6704);
or U11209 (N_11209,N_6705,N_8711);
xor U11210 (N_11210,N_7380,N_8604);
nor U11211 (N_11211,N_6962,N_6941);
xor U11212 (N_11212,N_9159,N_6641);
nor U11213 (N_11213,N_6805,N_8750);
or U11214 (N_11214,N_8340,N_8426);
and U11215 (N_11215,N_8972,N_8320);
nor U11216 (N_11216,N_8330,N_8845);
and U11217 (N_11217,N_7306,N_8782);
nand U11218 (N_11218,N_7765,N_8896);
xor U11219 (N_11219,N_6754,N_8709);
xnor U11220 (N_11220,N_8858,N_7946);
xnor U11221 (N_11221,N_8261,N_7848);
and U11222 (N_11222,N_6914,N_8725);
and U11223 (N_11223,N_9172,N_6929);
nor U11224 (N_11224,N_9042,N_8590);
nand U11225 (N_11225,N_7321,N_8160);
xor U11226 (N_11226,N_9321,N_7111);
or U11227 (N_11227,N_9350,N_6981);
or U11228 (N_11228,N_8130,N_9337);
nor U11229 (N_11229,N_8102,N_8325);
and U11230 (N_11230,N_7116,N_8658);
nor U11231 (N_11231,N_9305,N_8990);
xor U11232 (N_11232,N_8830,N_8978);
nand U11233 (N_11233,N_6407,N_8856);
and U11234 (N_11234,N_8111,N_6669);
or U11235 (N_11235,N_6748,N_6275);
nor U11236 (N_11236,N_7772,N_9050);
or U11237 (N_11237,N_8496,N_8276);
and U11238 (N_11238,N_8650,N_8366);
and U11239 (N_11239,N_6666,N_7748);
nor U11240 (N_11240,N_8316,N_7911);
nor U11241 (N_11241,N_8591,N_9089);
nor U11242 (N_11242,N_9371,N_8975);
or U11243 (N_11243,N_9176,N_7781);
and U11244 (N_11244,N_6364,N_6698);
nand U11245 (N_11245,N_7307,N_8864);
xor U11246 (N_11246,N_9140,N_7220);
nand U11247 (N_11247,N_6886,N_8206);
xnor U11248 (N_11248,N_8135,N_8710);
xnor U11249 (N_11249,N_8382,N_8307);
nand U11250 (N_11250,N_7543,N_6823);
and U11251 (N_11251,N_6977,N_6646);
nand U11252 (N_11252,N_6687,N_6916);
nand U11253 (N_11253,N_7933,N_8719);
and U11254 (N_11254,N_7560,N_7227);
nor U11255 (N_11255,N_7486,N_6488);
and U11256 (N_11256,N_6755,N_9066);
and U11257 (N_11257,N_6345,N_6645);
xnor U11258 (N_11258,N_6637,N_7248);
and U11259 (N_11259,N_8725,N_6457);
and U11260 (N_11260,N_7131,N_6322);
nand U11261 (N_11261,N_7314,N_9048);
nor U11262 (N_11262,N_8215,N_8873);
and U11263 (N_11263,N_8323,N_8694);
nor U11264 (N_11264,N_7305,N_7099);
nand U11265 (N_11265,N_7182,N_8750);
nor U11266 (N_11266,N_8849,N_9037);
nor U11267 (N_11267,N_7374,N_6417);
and U11268 (N_11268,N_8204,N_7938);
or U11269 (N_11269,N_6767,N_7165);
xor U11270 (N_11270,N_8676,N_6753);
nand U11271 (N_11271,N_7005,N_8760);
and U11272 (N_11272,N_8661,N_6925);
and U11273 (N_11273,N_9268,N_8471);
xor U11274 (N_11274,N_8130,N_6861);
and U11275 (N_11275,N_6396,N_8375);
xor U11276 (N_11276,N_7358,N_6756);
or U11277 (N_11277,N_8860,N_6542);
nand U11278 (N_11278,N_8196,N_8016);
xnor U11279 (N_11279,N_9205,N_6950);
and U11280 (N_11280,N_6328,N_6850);
xor U11281 (N_11281,N_8398,N_7044);
nor U11282 (N_11282,N_8002,N_6975);
nand U11283 (N_11283,N_7376,N_7879);
nand U11284 (N_11284,N_7155,N_6292);
nand U11285 (N_11285,N_7328,N_8310);
nor U11286 (N_11286,N_8141,N_8492);
nand U11287 (N_11287,N_9070,N_9116);
or U11288 (N_11288,N_7141,N_6754);
nand U11289 (N_11289,N_6864,N_9258);
nand U11290 (N_11290,N_7894,N_7436);
or U11291 (N_11291,N_7337,N_7663);
xor U11292 (N_11292,N_6861,N_7795);
nand U11293 (N_11293,N_9133,N_6859);
and U11294 (N_11294,N_8865,N_6909);
xnor U11295 (N_11295,N_6970,N_7208);
xnor U11296 (N_11296,N_7438,N_9192);
and U11297 (N_11297,N_6719,N_8280);
or U11298 (N_11298,N_8939,N_8487);
nor U11299 (N_11299,N_9097,N_9249);
and U11300 (N_11300,N_7783,N_7421);
or U11301 (N_11301,N_7071,N_9278);
and U11302 (N_11302,N_9242,N_6440);
nand U11303 (N_11303,N_8263,N_9062);
nor U11304 (N_11304,N_7714,N_7366);
nor U11305 (N_11305,N_7133,N_9115);
or U11306 (N_11306,N_8636,N_6298);
xor U11307 (N_11307,N_8793,N_6934);
or U11308 (N_11308,N_9074,N_7823);
nor U11309 (N_11309,N_9366,N_7753);
xnor U11310 (N_11310,N_8503,N_9127);
nor U11311 (N_11311,N_8706,N_6697);
or U11312 (N_11312,N_8233,N_7355);
and U11313 (N_11313,N_6943,N_7023);
or U11314 (N_11314,N_8693,N_6970);
and U11315 (N_11315,N_8193,N_6692);
nor U11316 (N_11316,N_7878,N_7591);
nor U11317 (N_11317,N_7709,N_6889);
xnor U11318 (N_11318,N_7738,N_8049);
nand U11319 (N_11319,N_6880,N_7142);
xnor U11320 (N_11320,N_8398,N_9266);
xor U11321 (N_11321,N_6766,N_6666);
xor U11322 (N_11322,N_7557,N_8838);
or U11323 (N_11323,N_8840,N_7835);
and U11324 (N_11324,N_9090,N_9183);
or U11325 (N_11325,N_8136,N_8835);
nor U11326 (N_11326,N_9307,N_8869);
or U11327 (N_11327,N_6707,N_9258);
nand U11328 (N_11328,N_6471,N_9036);
and U11329 (N_11329,N_9331,N_8509);
or U11330 (N_11330,N_7050,N_7655);
or U11331 (N_11331,N_9336,N_8411);
nand U11332 (N_11332,N_6876,N_7901);
nor U11333 (N_11333,N_7199,N_7129);
or U11334 (N_11334,N_8755,N_8992);
nor U11335 (N_11335,N_8464,N_6393);
xor U11336 (N_11336,N_8853,N_7996);
and U11337 (N_11337,N_8468,N_6799);
xnor U11338 (N_11338,N_8582,N_6977);
nand U11339 (N_11339,N_8841,N_7964);
or U11340 (N_11340,N_9334,N_6863);
nor U11341 (N_11341,N_6461,N_6365);
nand U11342 (N_11342,N_8658,N_7259);
xnor U11343 (N_11343,N_9340,N_9327);
and U11344 (N_11344,N_7531,N_6547);
xor U11345 (N_11345,N_6404,N_7474);
or U11346 (N_11346,N_8111,N_8973);
nor U11347 (N_11347,N_8676,N_8710);
and U11348 (N_11348,N_8585,N_6874);
nor U11349 (N_11349,N_8338,N_8431);
or U11350 (N_11350,N_7129,N_6703);
nor U11351 (N_11351,N_7253,N_8772);
or U11352 (N_11352,N_6951,N_8568);
nand U11353 (N_11353,N_8879,N_9129);
xnor U11354 (N_11354,N_8471,N_7883);
nor U11355 (N_11355,N_7409,N_6755);
nor U11356 (N_11356,N_8361,N_7791);
nor U11357 (N_11357,N_8689,N_7489);
xnor U11358 (N_11358,N_7000,N_8699);
nor U11359 (N_11359,N_9115,N_7954);
or U11360 (N_11360,N_7041,N_9323);
nor U11361 (N_11361,N_7394,N_8738);
and U11362 (N_11362,N_9221,N_9344);
nand U11363 (N_11363,N_7961,N_6948);
xor U11364 (N_11364,N_9196,N_6515);
or U11365 (N_11365,N_8491,N_8145);
and U11366 (N_11366,N_7014,N_9371);
and U11367 (N_11367,N_9025,N_7505);
or U11368 (N_11368,N_6517,N_7923);
nor U11369 (N_11369,N_9023,N_6473);
and U11370 (N_11370,N_7868,N_9325);
or U11371 (N_11371,N_6510,N_6552);
or U11372 (N_11372,N_6776,N_7297);
nand U11373 (N_11373,N_8235,N_7083);
and U11374 (N_11374,N_8278,N_9127);
or U11375 (N_11375,N_7475,N_9047);
or U11376 (N_11376,N_7313,N_8200);
or U11377 (N_11377,N_8285,N_7364);
or U11378 (N_11378,N_8867,N_8962);
and U11379 (N_11379,N_8277,N_6359);
nand U11380 (N_11380,N_7896,N_7181);
nand U11381 (N_11381,N_6575,N_6727);
xor U11382 (N_11382,N_6739,N_8941);
or U11383 (N_11383,N_7964,N_8644);
nand U11384 (N_11384,N_8825,N_6257);
or U11385 (N_11385,N_6961,N_8662);
nand U11386 (N_11386,N_6772,N_7618);
nand U11387 (N_11387,N_9270,N_8101);
or U11388 (N_11388,N_6412,N_8659);
xor U11389 (N_11389,N_8319,N_9317);
and U11390 (N_11390,N_7237,N_8946);
or U11391 (N_11391,N_7146,N_8111);
nand U11392 (N_11392,N_7823,N_7773);
or U11393 (N_11393,N_7565,N_6336);
or U11394 (N_11394,N_8487,N_7753);
or U11395 (N_11395,N_9096,N_8618);
xnor U11396 (N_11396,N_8597,N_6517);
and U11397 (N_11397,N_8253,N_8375);
and U11398 (N_11398,N_7461,N_8249);
xor U11399 (N_11399,N_7354,N_6310);
nand U11400 (N_11400,N_7193,N_8083);
nor U11401 (N_11401,N_6666,N_9300);
or U11402 (N_11402,N_7289,N_6585);
or U11403 (N_11403,N_7824,N_8260);
or U11404 (N_11404,N_6511,N_8362);
and U11405 (N_11405,N_6759,N_8807);
nand U11406 (N_11406,N_8674,N_9201);
xnor U11407 (N_11407,N_8513,N_7937);
and U11408 (N_11408,N_7997,N_6656);
nand U11409 (N_11409,N_8029,N_7076);
nor U11410 (N_11410,N_6885,N_6513);
or U11411 (N_11411,N_8669,N_9126);
nor U11412 (N_11412,N_6413,N_8077);
nand U11413 (N_11413,N_8882,N_8386);
or U11414 (N_11414,N_6687,N_8602);
nand U11415 (N_11415,N_9039,N_7436);
and U11416 (N_11416,N_8815,N_7475);
and U11417 (N_11417,N_8843,N_9300);
nor U11418 (N_11418,N_6896,N_8974);
or U11419 (N_11419,N_8425,N_6297);
and U11420 (N_11420,N_9013,N_8654);
or U11421 (N_11421,N_8156,N_7954);
nand U11422 (N_11422,N_9022,N_7326);
or U11423 (N_11423,N_9368,N_8484);
nand U11424 (N_11424,N_6761,N_9321);
xor U11425 (N_11425,N_7562,N_8721);
nand U11426 (N_11426,N_6320,N_6685);
xnor U11427 (N_11427,N_7000,N_7945);
nand U11428 (N_11428,N_7689,N_8777);
and U11429 (N_11429,N_6601,N_6385);
or U11430 (N_11430,N_8649,N_7786);
and U11431 (N_11431,N_9169,N_8465);
nand U11432 (N_11432,N_6511,N_7502);
xnor U11433 (N_11433,N_8036,N_7662);
xnor U11434 (N_11434,N_6651,N_6605);
xnor U11435 (N_11435,N_8735,N_8512);
xnor U11436 (N_11436,N_7522,N_9193);
xnor U11437 (N_11437,N_7077,N_6819);
xor U11438 (N_11438,N_7788,N_7875);
and U11439 (N_11439,N_8797,N_7646);
nand U11440 (N_11440,N_7233,N_9149);
xnor U11441 (N_11441,N_9282,N_8221);
and U11442 (N_11442,N_7341,N_8928);
xor U11443 (N_11443,N_7314,N_7882);
and U11444 (N_11444,N_8736,N_9078);
nand U11445 (N_11445,N_6361,N_6340);
or U11446 (N_11446,N_9334,N_8725);
and U11447 (N_11447,N_7897,N_7262);
xor U11448 (N_11448,N_7278,N_7380);
nand U11449 (N_11449,N_7572,N_8673);
nor U11450 (N_11450,N_7781,N_7785);
nand U11451 (N_11451,N_8296,N_7141);
nor U11452 (N_11452,N_7574,N_7673);
and U11453 (N_11453,N_6307,N_8445);
or U11454 (N_11454,N_7655,N_9085);
xnor U11455 (N_11455,N_7057,N_8187);
and U11456 (N_11456,N_7863,N_7053);
and U11457 (N_11457,N_6338,N_6741);
nor U11458 (N_11458,N_8073,N_7941);
nand U11459 (N_11459,N_8546,N_7589);
or U11460 (N_11460,N_7348,N_6724);
nand U11461 (N_11461,N_8193,N_7791);
nand U11462 (N_11462,N_8466,N_7842);
xor U11463 (N_11463,N_8701,N_6586);
or U11464 (N_11464,N_6565,N_6601);
xor U11465 (N_11465,N_6960,N_8707);
xnor U11466 (N_11466,N_9095,N_6827);
nor U11467 (N_11467,N_9249,N_6522);
nand U11468 (N_11468,N_8590,N_7157);
and U11469 (N_11469,N_7452,N_8015);
nand U11470 (N_11470,N_9090,N_8375);
nand U11471 (N_11471,N_6663,N_7413);
nand U11472 (N_11472,N_6492,N_7168);
xor U11473 (N_11473,N_6292,N_7049);
nor U11474 (N_11474,N_7739,N_7874);
and U11475 (N_11475,N_6552,N_6795);
nand U11476 (N_11476,N_8048,N_8219);
and U11477 (N_11477,N_9133,N_8728);
and U11478 (N_11478,N_7569,N_8583);
nand U11479 (N_11479,N_7160,N_6896);
or U11480 (N_11480,N_8622,N_8978);
nor U11481 (N_11481,N_8619,N_9278);
nor U11482 (N_11482,N_7346,N_7004);
xnor U11483 (N_11483,N_7741,N_6782);
or U11484 (N_11484,N_8710,N_6534);
and U11485 (N_11485,N_8246,N_7872);
xor U11486 (N_11486,N_6655,N_6402);
and U11487 (N_11487,N_7218,N_7010);
xnor U11488 (N_11488,N_8927,N_7075);
or U11489 (N_11489,N_9253,N_7289);
xor U11490 (N_11490,N_8559,N_7737);
or U11491 (N_11491,N_9238,N_8382);
and U11492 (N_11492,N_8165,N_7673);
nor U11493 (N_11493,N_9262,N_7394);
nor U11494 (N_11494,N_7208,N_6562);
nor U11495 (N_11495,N_8399,N_8269);
xor U11496 (N_11496,N_7931,N_9084);
nor U11497 (N_11497,N_7700,N_6251);
nor U11498 (N_11498,N_7381,N_7362);
nor U11499 (N_11499,N_7772,N_6916);
or U11500 (N_11500,N_8376,N_9232);
xor U11501 (N_11501,N_7162,N_8616);
nor U11502 (N_11502,N_9311,N_8494);
or U11503 (N_11503,N_7744,N_7116);
or U11504 (N_11504,N_7045,N_9222);
nor U11505 (N_11505,N_7204,N_7783);
nand U11506 (N_11506,N_8367,N_9125);
and U11507 (N_11507,N_8419,N_8507);
and U11508 (N_11508,N_7812,N_6560);
nor U11509 (N_11509,N_9209,N_7232);
xor U11510 (N_11510,N_9160,N_9037);
and U11511 (N_11511,N_8538,N_7416);
nand U11512 (N_11512,N_7201,N_8499);
xnor U11513 (N_11513,N_6389,N_8813);
and U11514 (N_11514,N_6869,N_9220);
nand U11515 (N_11515,N_8781,N_7648);
or U11516 (N_11516,N_7226,N_8658);
nor U11517 (N_11517,N_7927,N_7479);
or U11518 (N_11518,N_6628,N_6789);
xnor U11519 (N_11519,N_8093,N_6276);
nor U11520 (N_11520,N_6600,N_7156);
nand U11521 (N_11521,N_7467,N_8198);
xnor U11522 (N_11522,N_6806,N_6933);
nand U11523 (N_11523,N_7212,N_8307);
nand U11524 (N_11524,N_8839,N_8910);
nand U11525 (N_11525,N_7102,N_9210);
and U11526 (N_11526,N_8954,N_6604);
nor U11527 (N_11527,N_8087,N_7418);
xor U11528 (N_11528,N_6446,N_7657);
and U11529 (N_11529,N_6487,N_8989);
or U11530 (N_11530,N_6450,N_6468);
and U11531 (N_11531,N_8221,N_8401);
and U11532 (N_11532,N_8016,N_6820);
nand U11533 (N_11533,N_7027,N_6720);
nor U11534 (N_11534,N_9082,N_8640);
and U11535 (N_11535,N_8804,N_8094);
xor U11536 (N_11536,N_6989,N_9281);
nand U11537 (N_11537,N_8766,N_9005);
and U11538 (N_11538,N_7402,N_7978);
and U11539 (N_11539,N_6510,N_7575);
or U11540 (N_11540,N_9332,N_7866);
nand U11541 (N_11541,N_9372,N_6853);
nand U11542 (N_11542,N_8733,N_7918);
nor U11543 (N_11543,N_6522,N_6356);
nor U11544 (N_11544,N_7555,N_6422);
nor U11545 (N_11545,N_8978,N_7572);
xor U11546 (N_11546,N_8158,N_7624);
xor U11547 (N_11547,N_8274,N_8940);
nor U11548 (N_11548,N_8291,N_8125);
or U11549 (N_11549,N_7532,N_8565);
xnor U11550 (N_11550,N_8122,N_9374);
nor U11551 (N_11551,N_8994,N_7984);
nor U11552 (N_11552,N_7174,N_7716);
and U11553 (N_11553,N_7356,N_8876);
nand U11554 (N_11554,N_7361,N_8936);
nand U11555 (N_11555,N_6782,N_7794);
and U11556 (N_11556,N_9039,N_6264);
xnor U11557 (N_11557,N_7635,N_9362);
and U11558 (N_11558,N_8547,N_7836);
nor U11559 (N_11559,N_8354,N_8480);
nor U11560 (N_11560,N_7642,N_9248);
nand U11561 (N_11561,N_6683,N_9336);
nor U11562 (N_11562,N_8983,N_8845);
nand U11563 (N_11563,N_7396,N_6657);
xnor U11564 (N_11564,N_7861,N_6755);
or U11565 (N_11565,N_6761,N_7283);
or U11566 (N_11566,N_9299,N_9191);
or U11567 (N_11567,N_6496,N_7223);
and U11568 (N_11568,N_9034,N_6892);
nand U11569 (N_11569,N_9121,N_7499);
nand U11570 (N_11570,N_6814,N_7717);
or U11571 (N_11571,N_7904,N_6880);
and U11572 (N_11572,N_8899,N_7164);
nor U11573 (N_11573,N_6623,N_6652);
nand U11574 (N_11574,N_9294,N_8409);
and U11575 (N_11575,N_8641,N_9093);
and U11576 (N_11576,N_8449,N_8711);
or U11577 (N_11577,N_9329,N_6981);
xor U11578 (N_11578,N_7543,N_7542);
nand U11579 (N_11579,N_9292,N_8989);
nor U11580 (N_11580,N_7399,N_7240);
xor U11581 (N_11581,N_9094,N_6534);
xor U11582 (N_11582,N_9148,N_7494);
nand U11583 (N_11583,N_8529,N_7776);
nand U11584 (N_11584,N_8071,N_8630);
and U11585 (N_11585,N_7430,N_8923);
and U11586 (N_11586,N_7776,N_9321);
nor U11587 (N_11587,N_9282,N_7630);
or U11588 (N_11588,N_8057,N_9005);
or U11589 (N_11589,N_9026,N_7100);
nand U11590 (N_11590,N_8507,N_8353);
nand U11591 (N_11591,N_9052,N_6461);
nand U11592 (N_11592,N_6422,N_7932);
or U11593 (N_11593,N_7723,N_6490);
or U11594 (N_11594,N_7115,N_7285);
or U11595 (N_11595,N_7192,N_6965);
and U11596 (N_11596,N_8018,N_6969);
and U11597 (N_11597,N_6983,N_8213);
and U11598 (N_11598,N_8987,N_8661);
and U11599 (N_11599,N_7450,N_7548);
nand U11600 (N_11600,N_9052,N_6607);
xor U11601 (N_11601,N_7461,N_9367);
nor U11602 (N_11602,N_7268,N_7878);
nor U11603 (N_11603,N_7893,N_8348);
nor U11604 (N_11604,N_8405,N_8553);
and U11605 (N_11605,N_7460,N_6530);
nor U11606 (N_11606,N_8407,N_8066);
nor U11607 (N_11607,N_8515,N_6595);
xnor U11608 (N_11608,N_8963,N_8407);
xnor U11609 (N_11609,N_8485,N_7409);
or U11610 (N_11610,N_7555,N_6732);
xor U11611 (N_11611,N_7994,N_6552);
nor U11612 (N_11612,N_9337,N_7442);
nand U11613 (N_11613,N_7263,N_7050);
xnor U11614 (N_11614,N_6274,N_7141);
nand U11615 (N_11615,N_7399,N_8266);
nor U11616 (N_11616,N_6270,N_6502);
nor U11617 (N_11617,N_7430,N_6842);
nand U11618 (N_11618,N_8162,N_6369);
nand U11619 (N_11619,N_7307,N_9009);
or U11620 (N_11620,N_8986,N_9064);
and U11621 (N_11621,N_8199,N_6916);
nor U11622 (N_11622,N_9103,N_8675);
and U11623 (N_11623,N_8293,N_8337);
nand U11624 (N_11624,N_6967,N_7389);
nand U11625 (N_11625,N_9311,N_8502);
xor U11626 (N_11626,N_8166,N_8030);
nor U11627 (N_11627,N_6527,N_6579);
or U11628 (N_11628,N_6801,N_8374);
and U11629 (N_11629,N_6517,N_9088);
or U11630 (N_11630,N_9318,N_6402);
xor U11631 (N_11631,N_8884,N_7863);
or U11632 (N_11632,N_6348,N_8124);
nor U11633 (N_11633,N_9242,N_8769);
nor U11634 (N_11634,N_8106,N_8718);
or U11635 (N_11635,N_6328,N_8084);
xor U11636 (N_11636,N_9345,N_8846);
nor U11637 (N_11637,N_8808,N_8890);
xor U11638 (N_11638,N_7409,N_6815);
and U11639 (N_11639,N_8018,N_8162);
or U11640 (N_11640,N_6773,N_8707);
nand U11641 (N_11641,N_9288,N_8708);
nand U11642 (N_11642,N_8688,N_6374);
nor U11643 (N_11643,N_8140,N_9097);
nand U11644 (N_11644,N_7520,N_6787);
or U11645 (N_11645,N_8482,N_7403);
or U11646 (N_11646,N_7765,N_8540);
nand U11647 (N_11647,N_6939,N_9289);
nor U11648 (N_11648,N_8207,N_7855);
nand U11649 (N_11649,N_8146,N_8259);
nand U11650 (N_11650,N_8586,N_6636);
and U11651 (N_11651,N_9242,N_8036);
xor U11652 (N_11652,N_7468,N_8877);
xor U11653 (N_11653,N_7232,N_9114);
nor U11654 (N_11654,N_7643,N_8693);
nor U11655 (N_11655,N_7184,N_9209);
nand U11656 (N_11656,N_7031,N_7723);
and U11657 (N_11657,N_9020,N_8054);
and U11658 (N_11658,N_7858,N_7980);
xor U11659 (N_11659,N_7464,N_7165);
nand U11660 (N_11660,N_8567,N_9356);
or U11661 (N_11661,N_7287,N_7705);
xnor U11662 (N_11662,N_9204,N_9154);
or U11663 (N_11663,N_8964,N_6903);
and U11664 (N_11664,N_7527,N_7951);
and U11665 (N_11665,N_7550,N_8266);
nand U11666 (N_11666,N_6552,N_8440);
nor U11667 (N_11667,N_9374,N_6762);
or U11668 (N_11668,N_6933,N_7631);
nor U11669 (N_11669,N_8704,N_7927);
nand U11670 (N_11670,N_8517,N_7606);
and U11671 (N_11671,N_6875,N_6440);
and U11672 (N_11672,N_9044,N_9072);
nor U11673 (N_11673,N_8755,N_8785);
and U11674 (N_11674,N_6802,N_6824);
and U11675 (N_11675,N_7650,N_8478);
xor U11676 (N_11676,N_6863,N_8289);
xor U11677 (N_11677,N_6704,N_7378);
xnor U11678 (N_11678,N_7967,N_7078);
or U11679 (N_11679,N_8402,N_6316);
xor U11680 (N_11680,N_8253,N_6384);
or U11681 (N_11681,N_8203,N_7129);
or U11682 (N_11682,N_8383,N_7258);
nor U11683 (N_11683,N_8839,N_6921);
nand U11684 (N_11684,N_8053,N_6642);
nand U11685 (N_11685,N_7928,N_8732);
and U11686 (N_11686,N_8864,N_7300);
nor U11687 (N_11687,N_8862,N_7485);
nor U11688 (N_11688,N_8580,N_7851);
and U11689 (N_11689,N_8237,N_8066);
or U11690 (N_11690,N_7795,N_6615);
xor U11691 (N_11691,N_9361,N_8234);
or U11692 (N_11692,N_8147,N_8924);
or U11693 (N_11693,N_6610,N_7457);
or U11694 (N_11694,N_7282,N_8886);
nor U11695 (N_11695,N_7321,N_8295);
or U11696 (N_11696,N_7068,N_6699);
nor U11697 (N_11697,N_7068,N_6497);
nand U11698 (N_11698,N_9346,N_8876);
nand U11699 (N_11699,N_8124,N_6427);
xor U11700 (N_11700,N_7815,N_7617);
xnor U11701 (N_11701,N_6832,N_8533);
xnor U11702 (N_11702,N_8486,N_8191);
nor U11703 (N_11703,N_8656,N_7610);
nor U11704 (N_11704,N_6713,N_9155);
nor U11705 (N_11705,N_6750,N_8581);
xor U11706 (N_11706,N_7189,N_7342);
nand U11707 (N_11707,N_8445,N_6991);
nor U11708 (N_11708,N_6344,N_7172);
and U11709 (N_11709,N_6406,N_7764);
and U11710 (N_11710,N_9278,N_6650);
nand U11711 (N_11711,N_8670,N_6874);
nor U11712 (N_11712,N_9127,N_7663);
xnor U11713 (N_11713,N_6289,N_8388);
and U11714 (N_11714,N_8329,N_6486);
and U11715 (N_11715,N_6334,N_8297);
nor U11716 (N_11716,N_8863,N_8579);
or U11717 (N_11717,N_6775,N_7124);
and U11718 (N_11718,N_9173,N_7657);
nor U11719 (N_11719,N_7881,N_8311);
nor U11720 (N_11720,N_7208,N_8439);
xnor U11721 (N_11721,N_8124,N_8433);
and U11722 (N_11722,N_8484,N_6556);
or U11723 (N_11723,N_7105,N_8056);
or U11724 (N_11724,N_7681,N_6730);
and U11725 (N_11725,N_7577,N_7445);
nor U11726 (N_11726,N_8911,N_7765);
nor U11727 (N_11727,N_7357,N_6940);
xnor U11728 (N_11728,N_8819,N_6627);
xnor U11729 (N_11729,N_8954,N_8694);
nand U11730 (N_11730,N_7216,N_6871);
and U11731 (N_11731,N_8600,N_6888);
or U11732 (N_11732,N_8438,N_6625);
xnor U11733 (N_11733,N_6299,N_8263);
nor U11734 (N_11734,N_7143,N_9012);
nor U11735 (N_11735,N_7448,N_8464);
and U11736 (N_11736,N_7121,N_6347);
nand U11737 (N_11737,N_6955,N_9105);
and U11738 (N_11738,N_8783,N_9303);
nor U11739 (N_11739,N_9343,N_8435);
nor U11740 (N_11740,N_9059,N_8217);
nor U11741 (N_11741,N_9367,N_7119);
nor U11742 (N_11742,N_9276,N_9312);
xnor U11743 (N_11743,N_7410,N_6287);
and U11744 (N_11744,N_9188,N_9285);
and U11745 (N_11745,N_8443,N_8773);
or U11746 (N_11746,N_6533,N_8675);
and U11747 (N_11747,N_6632,N_8724);
and U11748 (N_11748,N_7344,N_6786);
or U11749 (N_11749,N_8626,N_7714);
or U11750 (N_11750,N_6423,N_6555);
nand U11751 (N_11751,N_6873,N_7398);
or U11752 (N_11752,N_7176,N_8035);
or U11753 (N_11753,N_6287,N_8952);
or U11754 (N_11754,N_8645,N_7438);
nand U11755 (N_11755,N_8033,N_7070);
and U11756 (N_11756,N_8494,N_7488);
nor U11757 (N_11757,N_6828,N_8222);
xor U11758 (N_11758,N_8992,N_6280);
nand U11759 (N_11759,N_6994,N_8608);
nand U11760 (N_11760,N_8129,N_6787);
or U11761 (N_11761,N_6828,N_9160);
and U11762 (N_11762,N_6605,N_8234);
xnor U11763 (N_11763,N_7768,N_8776);
nor U11764 (N_11764,N_6635,N_6485);
nor U11765 (N_11765,N_6361,N_8492);
nor U11766 (N_11766,N_8136,N_9036);
xor U11767 (N_11767,N_6808,N_7978);
nor U11768 (N_11768,N_7133,N_7883);
or U11769 (N_11769,N_7057,N_8340);
nand U11770 (N_11770,N_7904,N_8863);
xor U11771 (N_11771,N_6817,N_6901);
nor U11772 (N_11772,N_6962,N_7599);
nand U11773 (N_11773,N_8059,N_7921);
xor U11774 (N_11774,N_9176,N_7919);
xnor U11775 (N_11775,N_8324,N_6983);
or U11776 (N_11776,N_6447,N_6984);
or U11777 (N_11777,N_9230,N_7764);
nand U11778 (N_11778,N_7233,N_8329);
nor U11779 (N_11779,N_8103,N_9139);
xor U11780 (N_11780,N_8931,N_8107);
and U11781 (N_11781,N_7284,N_6368);
and U11782 (N_11782,N_8002,N_7567);
or U11783 (N_11783,N_7436,N_7405);
or U11784 (N_11784,N_8263,N_8268);
and U11785 (N_11785,N_7547,N_6671);
and U11786 (N_11786,N_9026,N_6954);
xor U11787 (N_11787,N_7921,N_8957);
and U11788 (N_11788,N_9215,N_7849);
nand U11789 (N_11789,N_8311,N_7309);
or U11790 (N_11790,N_7825,N_6386);
or U11791 (N_11791,N_8630,N_8258);
nor U11792 (N_11792,N_6372,N_8394);
nor U11793 (N_11793,N_8043,N_6592);
nor U11794 (N_11794,N_7149,N_8339);
or U11795 (N_11795,N_6782,N_8055);
nand U11796 (N_11796,N_7719,N_8669);
or U11797 (N_11797,N_6447,N_6893);
xnor U11798 (N_11798,N_8274,N_8390);
xnor U11799 (N_11799,N_7819,N_6822);
or U11800 (N_11800,N_6407,N_9210);
xor U11801 (N_11801,N_9060,N_6860);
xor U11802 (N_11802,N_6273,N_8567);
nand U11803 (N_11803,N_8604,N_8953);
and U11804 (N_11804,N_8474,N_8727);
and U11805 (N_11805,N_7120,N_8228);
xnor U11806 (N_11806,N_9181,N_8892);
xor U11807 (N_11807,N_7288,N_8312);
and U11808 (N_11808,N_7000,N_8653);
nand U11809 (N_11809,N_6779,N_8519);
nor U11810 (N_11810,N_7232,N_8536);
or U11811 (N_11811,N_8894,N_8574);
and U11812 (N_11812,N_9352,N_7242);
nor U11813 (N_11813,N_9277,N_7569);
nand U11814 (N_11814,N_6990,N_7671);
xnor U11815 (N_11815,N_8553,N_8784);
nor U11816 (N_11816,N_7766,N_8563);
nand U11817 (N_11817,N_9021,N_9263);
or U11818 (N_11818,N_8349,N_8536);
nor U11819 (N_11819,N_8976,N_7792);
and U11820 (N_11820,N_8193,N_8562);
and U11821 (N_11821,N_7751,N_9139);
or U11822 (N_11822,N_7175,N_9256);
and U11823 (N_11823,N_8362,N_6842);
xnor U11824 (N_11824,N_7318,N_6480);
or U11825 (N_11825,N_7906,N_7942);
and U11826 (N_11826,N_9273,N_7271);
nor U11827 (N_11827,N_7112,N_7673);
or U11828 (N_11828,N_7889,N_8898);
and U11829 (N_11829,N_9215,N_6816);
or U11830 (N_11830,N_7655,N_7145);
nor U11831 (N_11831,N_6665,N_7038);
or U11832 (N_11832,N_9008,N_7161);
and U11833 (N_11833,N_6980,N_6370);
xnor U11834 (N_11834,N_6383,N_7098);
nand U11835 (N_11835,N_8074,N_6490);
or U11836 (N_11836,N_8044,N_7064);
and U11837 (N_11837,N_8468,N_8294);
and U11838 (N_11838,N_8428,N_6700);
or U11839 (N_11839,N_8363,N_8307);
nand U11840 (N_11840,N_6903,N_8038);
and U11841 (N_11841,N_6997,N_8772);
nor U11842 (N_11842,N_8638,N_7433);
and U11843 (N_11843,N_8516,N_8295);
nand U11844 (N_11844,N_8393,N_8837);
and U11845 (N_11845,N_6672,N_6947);
nand U11846 (N_11846,N_9170,N_7726);
and U11847 (N_11847,N_8712,N_8526);
or U11848 (N_11848,N_7413,N_8389);
xnor U11849 (N_11849,N_8068,N_8466);
and U11850 (N_11850,N_8666,N_8145);
nor U11851 (N_11851,N_7911,N_9134);
nor U11852 (N_11852,N_9139,N_6577);
nand U11853 (N_11853,N_6874,N_7988);
nor U11854 (N_11854,N_6276,N_7133);
or U11855 (N_11855,N_6998,N_7060);
or U11856 (N_11856,N_9091,N_6451);
nor U11857 (N_11857,N_6717,N_8994);
nor U11858 (N_11858,N_7890,N_9266);
or U11859 (N_11859,N_8538,N_7691);
or U11860 (N_11860,N_8629,N_9046);
nor U11861 (N_11861,N_9350,N_8188);
or U11862 (N_11862,N_7612,N_8991);
nand U11863 (N_11863,N_6551,N_7148);
or U11864 (N_11864,N_6368,N_9167);
or U11865 (N_11865,N_8040,N_8457);
or U11866 (N_11866,N_6401,N_6926);
nand U11867 (N_11867,N_8220,N_7741);
or U11868 (N_11868,N_7487,N_8044);
or U11869 (N_11869,N_9015,N_6582);
nand U11870 (N_11870,N_8815,N_8379);
nand U11871 (N_11871,N_7100,N_8636);
nor U11872 (N_11872,N_9223,N_9132);
nor U11873 (N_11873,N_6572,N_7027);
xnor U11874 (N_11874,N_6978,N_6478);
and U11875 (N_11875,N_6496,N_7750);
or U11876 (N_11876,N_7362,N_6522);
nor U11877 (N_11877,N_6294,N_7912);
and U11878 (N_11878,N_7180,N_6651);
or U11879 (N_11879,N_6634,N_9250);
or U11880 (N_11880,N_9095,N_6711);
nand U11881 (N_11881,N_6527,N_8152);
or U11882 (N_11882,N_8667,N_6842);
xnor U11883 (N_11883,N_6759,N_8600);
nor U11884 (N_11884,N_6857,N_7225);
nand U11885 (N_11885,N_7680,N_7854);
or U11886 (N_11886,N_7995,N_8115);
and U11887 (N_11887,N_6301,N_8577);
nor U11888 (N_11888,N_7137,N_8884);
and U11889 (N_11889,N_6474,N_9077);
or U11890 (N_11890,N_7756,N_7915);
nor U11891 (N_11891,N_8539,N_8512);
nor U11892 (N_11892,N_8782,N_8346);
nand U11893 (N_11893,N_9116,N_6995);
or U11894 (N_11894,N_6614,N_6850);
and U11895 (N_11895,N_9335,N_8287);
xor U11896 (N_11896,N_6698,N_8290);
nand U11897 (N_11897,N_8628,N_6313);
nor U11898 (N_11898,N_7589,N_7450);
and U11899 (N_11899,N_6473,N_8151);
and U11900 (N_11900,N_8791,N_7615);
or U11901 (N_11901,N_6992,N_6273);
or U11902 (N_11902,N_7973,N_8429);
xnor U11903 (N_11903,N_7811,N_8935);
nor U11904 (N_11904,N_8585,N_8080);
nand U11905 (N_11905,N_8514,N_7259);
xor U11906 (N_11906,N_7181,N_7689);
nor U11907 (N_11907,N_9174,N_8847);
xnor U11908 (N_11908,N_8204,N_9119);
or U11909 (N_11909,N_7782,N_8420);
nor U11910 (N_11910,N_7388,N_7867);
nor U11911 (N_11911,N_7477,N_6763);
xor U11912 (N_11912,N_9209,N_7360);
nor U11913 (N_11913,N_6299,N_7849);
and U11914 (N_11914,N_8784,N_9350);
or U11915 (N_11915,N_9114,N_7396);
nor U11916 (N_11916,N_8808,N_9091);
nor U11917 (N_11917,N_6594,N_8393);
nor U11918 (N_11918,N_6905,N_6424);
and U11919 (N_11919,N_6396,N_8515);
nor U11920 (N_11920,N_7856,N_9065);
xor U11921 (N_11921,N_9151,N_8345);
nand U11922 (N_11922,N_6929,N_8045);
nor U11923 (N_11923,N_6478,N_7752);
or U11924 (N_11924,N_7206,N_6657);
xnor U11925 (N_11925,N_7338,N_6692);
xnor U11926 (N_11926,N_8954,N_9241);
xor U11927 (N_11927,N_8718,N_6727);
or U11928 (N_11928,N_7668,N_7514);
nor U11929 (N_11929,N_9334,N_6876);
xnor U11930 (N_11930,N_7022,N_9321);
nand U11931 (N_11931,N_8155,N_9092);
nand U11932 (N_11932,N_7253,N_7880);
or U11933 (N_11933,N_6294,N_8943);
and U11934 (N_11934,N_6832,N_9200);
xor U11935 (N_11935,N_8893,N_8370);
or U11936 (N_11936,N_8571,N_8240);
xor U11937 (N_11937,N_6711,N_7660);
or U11938 (N_11938,N_6274,N_8239);
and U11939 (N_11939,N_7777,N_8261);
nor U11940 (N_11940,N_7658,N_8993);
nand U11941 (N_11941,N_8174,N_7092);
or U11942 (N_11942,N_7109,N_6273);
xnor U11943 (N_11943,N_6499,N_9135);
nor U11944 (N_11944,N_6485,N_8576);
nand U11945 (N_11945,N_7615,N_8116);
xnor U11946 (N_11946,N_8723,N_6939);
xnor U11947 (N_11947,N_8056,N_7612);
nor U11948 (N_11948,N_6637,N_7109);
and U11949 (N_11949,N_6704,N_8201);
xor U11950 (N_11950,N_6343,N_9108);
nor U11951 (N_11951,N_7015,N_8776);
or U11952 (N_11952,N_9323,N_7498);
or U11953 (N_11953,N_8496,N_8750);
xnor U11954 (N_11954,N_7606,N_8970);
or U11955 (N_11955,N_7940,N_9172);
xnor U11956 (N_11956,N_6445,N_7984);
nor U11957 (N_11957,N_9322,N_8108);
or U11958 (N_11958,N_7554,N_7482);
or U11959 (N_11959,N_7653,N_6780);
nand U11960 (N_11960,N_6922,N_7473);
or U11961 (N_11961,N_8641,N_7168);
and U11962 (N_11962,N_6599,N_6826);
or U11963 (N_11963,N_7269,N_7259);
and U11964 (N_11964,N_9065,N_8356);
nand U11965 (N_11965,N_7271,N_7214);
and U11966 (N_11966,N_8368,N_6468);
or U11967 (N_11967,N_7359,N_8019);
xor U11968 (N_11968,N_6340,N_8317);
nor U11969 (N_11969,N_6631,N_7931);
nor U11970 (N_11970,N_9092,N_6369);
xnor U11971 (N_11971,N_7708,N_7638);
nand U11972 (N_11972,N_6358,N_7976);
nand U11973 (N_11973,N_6476,N_9326);
xnor U11974 (N_11974,N_6578,N_9230);
and U11975 (N_11975,N_6604,N_7730);
xor U11976 (N_11976,N_7926,N_8131);
or U11977 (N_11977,N_8802,N_7289);
nor U11978 (N_11978,N_9041,N_8445);
or U11979 (N_11979,N_7343,N_6537);
xnor U11980 (N_11980,N_9188,N_8458);
nor U11981 (N_11981,N_7617,N_8830);
xnor U11982 (N_11982,N_7834,N_8583);
nand U11983 (N_11983,N_6844,N_7159);
or U11984 (N_11984,N_6466,N_6423);
or U11985 (N_11985,N_7388,N_7065);
xor U11986 (N_11986,N_8357,N_7423);
and U11987 (N_11987,N_8271,N_6620);
nor U11988 (N_11988,N_7180,N_9145);
nand U11989 (N_11989,N_7124,N_7760);
and U11990 (N_11990,N_6697,N_6710);
nand U11991 (N_11991,N_9241,N_7592);
nand U11992 (N_11992,N_7094,N_7347);
nor U11993 (N_11993,N_9190,N_8062);
nor U11994 (N_11994,N_7040,N_7552);
and U11995 (N_11995,N_7658,N_6809);
xnor U11996 (N_11996,N_7512,N_6801);
nor U11997 (N_11997,N_8266,N_6688);
xor U11998 (N_11998,N_8936,N_6490);
nor U11999 (N_11999,N_8135,N_7435);
xnor U12000 (N_12000,N_7369,N_8737);
and U12001 (N_12001,N_8134,N_6911);
nand U12002 (N_12002,N_7803,N_7686);
xnor U12003 (N_12003,N_7513,N_7511);
or U12004 (N_12004,N_6823,N_8616);
or U12005 (N_12005,N_9054,N_8532);
nor U12006 (N_12006,N_6294,N_6606);
nor U12007 (N_12007,N_7379,N_8604);
nand U12008 (N_12008,N_6984,N_7727);
nand U12009 (N_12009,N_6572,N_7583);
and U12010 (N_12010,N_8852,N_7273);
nor U12011 (N_12011,N_7954,N_6924);
nand U12012 (N_12012,N_7576,N_6738);
and U12013 (N_12013,N_8118,N_6911);
and U12014 (N_12014,N_8450,N_7239);
nand U12015 (N_12015,N_6613,N_9095);
nand U12016 (N_12016,N_7923,N_7345);
nand U12017 (N_12017,N_6913,N_7617);
nor U12018 (N_12018,N_8182,N_6989);
nor U12019 (N_12019,N_8382,N_6630);
nand U12020 (N_12020,N_7080,N_8070);
and U12021 (N_12021,N_7262,N_7233);
and U12022 (N_12022,N_6703,N_8926);
nand U12023 (N_12023,N_9211,N_7467);
nand U12024 (N_12024,N_7760,N_8623);
nor U12025 (N_12025,N_8740,N_8357);
nand U12026 (N_12026,N_6501,N_9007);
or U12027 (N_12027,N_7026,N_8213);
xnor U12028 (N_12028,N_9129,N_6645);
nor U12029 (N_12029,N_7990,N_6789);
or U12030 (N_12030,N_8052,N_8001);
nor U12031 (N_12031,N_8994,N_6857);
xnor U12032 (N_12032,N_8659,N_7437);
or U12033 (N_12033,N_9292,N_8025);
nor U12034 (N_12034,N_6795,N_8458);
nand U12035 (N_12035,N_7494,N_9314);
nand U12036 (N_12036,N_7677,N_9225);
nor U12037 (N_12037,N_9269,N_6418);
nand U12038 (N_12038,N_7299,N_9323);
or U12039 (N_12039,N_6983,N_6888);
xor U12040 (N_12040,N_7064,N_7575);
nand U12041 (N_12041,N_7392,N_6716);
nor U12042 (N_12042,N_7543,N_8196);
xnor U12043 (N_12043,N_7232,N_8203);
nand U12044 (N_12044,N_8113,N_7349);
or U12045 (N_12045,N_7496,N_7536);
nand U12046 (N_12046,N_9012,N_8011);
nor U12047 (N_12047,N_7051,N_8182);
nand U12048 (N_12048,N_8040,N_7630);
xnor U12049 (N_12049,N_8378,N_6954);
nor U12050 (N_12050,N_9331,N_6957);
and U12051 (N_12051,N_8568,N_9134);
xor U12052 (N_12052,N_9136,N_6588);
nand U12053 (N_12053,N_6318,N_9222);
and U12054 (N_12054,N_8602,N_8786);
nor U12055 (N_12055,N_6758,N_9212);
and U12056 (N_12056,N_8341,N_6423);
and U12057 (N_12057,N_9291,N_8067);
nor U12058 (N_12058,N_7731,N_8215);
and U12059 (N_12059,N_6513,N_6663);
nand U12060 (N_12060,N_6633,N_7504);
xor U12061 (N_12061,N_8531,N_8434);
and U12062 (N_12062,N_7106,N_9290);
nand U12063 (N_12063,N_7150,N_8092);
or U12064 (N_12064,N_6521,N_7539);
nand U12065 (N_12065,N_7989,N_8778);
xnor U12066 (N_12066,N_8376,N_7644);
or U12067 (N_12067,N_8758,N_9213);
nor U12068 (N_12068,N_7627,N_8589);
nor U12069 (N_12069,N_8694,N_8623);
and U12070 (N_12070,N_9110,N_7238);
xnor U12071 (N_12071,N_8790,N_9333);
and U12072 (N_12072,N_9205,N_7737);
xor U12073 (N_12073,N_9003,N_7535);
nand U12074 (N_12074,N_6587,N_6381);
or U12075 (N_12075,N_6635,N_8779);
nand U12076 (N_12076,N_8099,N_8512);
nand U12077 (N_12077,N_7897,N_8036);
and U12078 (N_12078,N_7038,N_8545);
or U12079 (N_12079,N_9267,N_9016);
and U12080 (N_12080,N_7609,N_7990);
or U12081 (N_12081,N_9103,N_7875);
xor U12082 (N_12082,N_9080,N_7815);
nor U12083 (N_12083,N_6962,N_6361);
or U12084 (N_12084,N_6683,N_9249);
nand U12085 (N_12085,N_8948,N_7566);
nor U12086 (N_12086,N_9174,N_7520);
xor U12087 (N_12087,N_8115,N_8498);
or U12088 (N_12088,N_7798,N_7946);
nor U12089 (N_12089,N_6785,N_8972);
nor U12090 (N_12090,N_7521,N_7944);
nand U12091 (N_12091,N_7950,N_8124);
xor U12092 (N_12092,N_8217,N_6580);
and U12093 (N_12093,N_7536,N_8981);
xnor U12094 (N_12094,N_7314,N_8257);
nand U12095 (N_12095,N_6445,N_7033);
nand U12096 (N_12096,N_8529,N_7153);
and U12097 (N_12097,N_7415,N_7656);
xnor U12098 (N_12098,N_7394,N_7197);
and U12099 (N_12099,N_8594,N_7796);
or U12100 (N_12100,N_6643,N_7863);
xor U12101 (N_12101,N_9075,N_8995);
xnor U12102 (N_12102,N_7334,N_8967);
nor U12103 (N_12103,N_6767,N_9130);
and U12104 (N_12104,N_7745,N_7565);
nor U12105 (N_12105,N_7979,N_9308);
xnor U12106 (N_12106,N_7648,N_7437);
xnor U12107 (N_12107,N_7631,N_6362);
nand U12108 (N_12108,N_6802,N_7165);
or U12109 (N_12109,N_6260,N_8361);
nand U12110 (N_12110,N_6426,N_7918);
and U12111 (N_12111,N_8559,N_8590);
nor U12112 (N_12112,N_7652,N_8472);
and U12113 (N_12113,N_6392,N_8787);
nor U12114 (N_12114,N_8685,N_7865);
and U12115 (N_12115,N_6425,N_7558);
xnor U12116 (N_12116,N_6892,N_8039);
and U12117 (N_12117,N_6551,N_7452);
or U12118 (N_12118,N_7673,N_7589);
or U12119 (N_12119,N_8295,N_6755);
xor U12120 (N_12120,N_7829,N_6860);
and U12121 (N_12121,N_7305,N_6874);
and U12122 (N_12122,N_6346,N_7877);
and U12123 (N_12123,N_6801,N_9349);
xor U12124 (N_12124,N_6478,N_8759);
nand U12125 (N_12125,N_9327,N_8096);
nand U12126 (N_12126,N_9044,N_7111);
or U12127 (N_12127,N_7768,N_7440);
and U12128 (N_12128,N_7009,N_7058);
and U12129 (N_12129,N_8317,N_6639);
and U12130 (N_12130,N_9047,N_8689);
nand U12131 (N_12131,N_6917,N_7418);
or U12132 (N_12132,N_8218,N_8887);
xnor U12133 (N_12133,N_9252,N_8379);
nand U12134 (N_12134,N_8539,N_7074);
nand U12135 (N_12135,N_8449,N_8535);
xnor U12136 (N_12136,N_6325,N_7256);
xnor U12137 (N_12137,N_8444,N_6761);
nand U12138 (N_12138,N_8261,N_9126);
and U12139 (N_12139,N_7160,N_8034);
and U12140 (N_12140,N_8439,N_9184);
and U12141 (N_12141,N_7904,N_9350);
or U12142 (N_12142,N_8009,N_8560);
or U12143 (N_12143,N_8861,N_6756);
and U12144 (N_12144,N_7735,N_7892);
or U12145 (N_12145,N_8441,N_7921);
and U12146 (N_12146,N_7785,N_7530);
or U12147 (N_12147,N_7321,N_9254);
nor U12148 (N_12148,N_8296,N_7380);
xor U12149 (N_12149,N_9257,N_8840);
nor U12150 (N_12150,N_6366,N_7289);
or U12151 (N_12151,N_9254,N_8847);
and U12152 (N_12152,N_7989,N_7976);
or U12153 (N_12153,N_7025,N_7936);
xnor U12154 (N_12154,N_7146,N_7755);
xor U12155 (N_12155,N_7422,N_8520);
and U12156 (N_12156,N_9151,N_8011);
xor U12157 (N_12157,N_6978,N_8147);
nand U12158 (N_12158,N_8894,N_7278);
and U12159 (N_12159,N_7355,N_7624);
and U12160 (N_12160,N_7669,N_6905);
nor U12161 (N_12161,N_8419,N_8305);
xor U12162 (N_12162,N_7930,N_6659);
nand U12163 (N_12163,N_8660,N_8449);
and U12164 (N_12164,N_8121,N_8762);
nor U12165 (N_12165,N_8256,N_8066);
xor U12166 (N_12166,N_7374,N_8310);
or U12167 (N_12167,N_8017,N_9301);
and U12168 (N_12168,N_8074,N_7385);
nand U12169 (N_12169,N_9303,N_6404);
and U12170 (N_12170,N_8098,N_9192);
nand U12171 (N_12171,N_7602,N_8491);
or U12172 (N_12172,N_6951,N_8258);
and U12173 (N_12173,N_7511,N_9293);
or U12174 (N_12174,N_7387,N_6778);
nor U12175 (N_12175,N_8063,N_7589);
and U12176 (N_12176,N_6991,N_8498);
xor U12177 (N_12177,N_6324,N_6387);
and U12178 (N_12178,N_6651,N_7680);
xor U12179 (N_12179,N_7828,N_6312);
nand U12180 (N_12180,N_8561,N_8669);
nor U12181 (N_12181,N_6675,N_7860);
nor U12182 (N_12182,N_8373,N_8991);
nor U12183 (N_12183,N_8554,N_8734);
and U12184 (N_12184,N_8164,N_6278);
and U12185 (N_12185,N_8714,N_7413);
or U12186 (N_12186,N_7131,N_7281);
nor U12187 (N_12187,N_9065,N_8426);
and U12188 (N_12188,N_8638,N_8056);
or U12189 (N_12189,N_7486,N_7399);
and U12190 (N_12190,N_6982,N_6833);
nand U12191 (N_12191,N_6954,N_7398);
nor U12192 (N_12192,N_6485,N_7476);
and U12193 (N_12193,N_9165,N_8841);
or U12194 (N_12194,N_9016,N_8810);
xnor U12195 (N_12195,N_7808,N_7095);
or U12196 (N_12196,N_8515,N_8353);
nand U12197 (N_12197,N_6942,N_8063);
and U12198 (N_12198,N_6824,N_6612);
nand U12199 (N_12199,N_6271,N_6412);
and U12200 (N_12200,N_6491,N_9224);
nand U12201 (N_12201,N_7042,N_8744);
xor U12202 (N_12202,N_9301,N_7694);
and U12203 (N_12203,N_6551,N_8569);
nor U12204 (N_12204,N_8024,N_7661);
xnor U12205 (N_12205,N_8910,N_7075);
nor U12206 (N_12206,N_6870,N_8939);
or U12207 (N_12207,N_8942,N_8974);
or U12208 (N_12208,N_7485,N_7984);
nor U12209 (N_12209,N_7731,N_7927);
or U12210 (N_12210,N_7422,N_7967);
nand U12211 (N_12211,N_8018,N_6799);
nor U12212 (N_12212,N_7950,N_6557);
nand U12213 (N_12213,N_8321,N_9038);
and U12214 (N_12214,N_8248,N_8669);
nor U12215 (N_12215,N_8694,N_6720);
and U12216 (N_12216,N_8587,N_6695);
and U12217 (N_12217,N_8044,N_6429);
or U12218 (N_12218,N_7980,N_6395);
and U12219 (N_12219,N_8703,N_8537);
nor U12220 (N_12220,N_6750,N_7553);
nor U12221 (N_12221,N_8711,N_8087);
nor U12222 (N_12222,N_7369,N_6480);
xor U12223 (N_12223,N_9186,N_9294);
nand U12224 (N_12224,N_8947,N_9244);
or U12225 (N_12225,N_7067,N_7694);
and U12226 (N_12226,N_7380,N_8744);
nand U12227 (N_12227,N_8907,N_7895);
xor U12228 (N_12228,N_7987,N_6896);
or U12229 (N_12229,N_6910,N_7196);
nor U12230 (N_12230,N_8176,N_8965);
and U12231 (N_12231,N_8072,N_6943);
xnor U12232 (N_12232,N_7624,N_7033);
xor U12233 (N_12233,N_7646,N_8736);
or U12234 (N_12234,N_8492,N_8078);
nand U12235 (N_12235,N_8680,N_6308);
or U12236 (N_12236,N_8392,N_6443);
nand U12237 (N_12237,N_8652,N_7496);
nor U12238 (N_12238,N_6984,N_8475);
xnor U12239 (N_12239,N_7986,N_9230);
or U12240 (N_12240,N_8756,N_9232);
nand U12241 (N_12241,N_7290,N_6635);
nor U12242 (N_12242,N_8708,N_7435);
and U12243 (N_12243,N_7046,N_7660);
or U12244 (N_12244,N_7357,N_7754);
nor U12245 (N_12245,N_6444,N_7532);
and U12246 (N_12246,N_7686,N_8426);
xnor U12247 (N_12247,N_7767,N_8361);
or U12248 (N_12248,N_8160,N_8007);
and U12249 (N_12249,N_7605,N_8972);
nand U12250 (N_12250,N_8318,N_8248);
or U12251 (N_12251,N_6885,N_8887);
or U12252 (N_12252,N_9218,N_8719);
or U12253 (N_12253,N_6506,N_8411);
xor U12254 (N_12254,N_7909,N_7567);
or U12255 (N_12255,N_7853,N_9038);
nor U12256 (N_12256,N_8379,N_8764);
nand U12257 (N_12257,N_7090,N_8551);
nor U12258 (N_12258,N_7162,N_6629);
and U12259 (N_12259,N_6319,N_8594);
nor U12260 (N_12260,N_7146,N_9358);
or U12261 (N_12261,N_7512,N_7700);
nand U12262 (N_12262,N_6628,N_9137);
nand U12263 (N_12263,N_6331,N_7046);
or U12264 (N_12264,N_9312,N_6921);
xor U12265 (N_12265,N_8500,N_7907);
nor U12266 (N_12266,N_6910,N_6966);
nor U12267 (N_12267,N_9374,N_7221);
nor U12268 (N_12268,N_9260,N_9209);
nor U12269 (N_12269,N_6689,N_8225);
xor U12270 (N_12270,N_8745,N_7214);
nand U12271 (N_12271,N_9265,N_9162);
nand U12272 (N_12272,N_7146,N_6532);
or U12273 (N_12273,N_8332,N_8024);
xor U12274 (N_12274,N_9066,N_7482);
or U12275 (N_12275,N_7839,N_6654);
and U12276 (N_12276,N_6898,N_6469);
or U12277 (N_12277,N_7617,N_8982);
and U12278 (N_12278,N_9148,N_9137);
and U12279 (N_12279,N_6703,N_6902);
nand U12280 (N_12280,N_9195,N_7250);
nor U12281 (N_12281,N_6341,N_8973);
nor U12282 (N_12282,N_7398,N_9258);
or U12283 (N_12283,N_8539,N_8276);
or U12284 (N_12284,N_8573,N_8902);
xor U12285 (N_12285,N_8961,N_6694);
or U12286 (N_12286,N_8572,N_9194);
nand U12287 (N_12287,N_7483,N_7346);
nand U12288 (N_12288,N_6713,N_8899);
nor U12289 (N_12289,N_8326,N_7235);
nor U12290 (N_12290,N_8048,N_7110);
nor U12291 (N_12291,N_7353,N_8580);
nor U12292 (N_12292,N_6322,N_9237);
xor U12293 (N_12293,N_8147,N_7427);
and U12294 (N_12294,N_7157,N_7248);
or U12295 (N_12295,N_8071,N_7628);
or U12296 (N_12296,N_8704,N_8263);
or U12297 (N_12297,N_9300,N_6995);
nor U12298 (N_12298,N_8575,N_7289);
nor U12299 (N_12299,N_7764,N_7609);
nor U12300 (N_12300,N_6477,N_8727);
or U12301 (N_12301,N_8295,N_8995);
xor U12302 (N_12302,N_6470,N_7854);
or U12303 (N_12303,N_6994,N_7470);
or U12304 (N_12304,N_9048,N_8405);
and U12305 (N_12305,N_7435,N_7462);
or U12306 (N_12306,N_8415,N_8265);
nor U12307 (N_12307,N_7450,N_6524);
xor U12308 (N_12308,N_7506,N_7091);
or U12309 (N_12309,N_7894,N_8075);
xor U12310 (N_12310,N_8430,N_6388);
or U12311 (N_12311,N_7790,N_9317);
or U12312 (N_12312,N_8769,N_6347);
xnor U12313 (N_12313,N_8456,N_7970);
xor U12314 (N_12314,N_9164,N_8607);
xor U12315 (N_12315,N_9120,N_6431);
or U12316 (N_12316,N_7787,N_8506);
nor U12317 (N_12317,N_8705,N_7872);
or U12318 (N_12318,N_8882,N_9196);
and U12319 (N_12319,N_9242,N_6745);
or U12320 (N_12320,N_9108,N_8358);
nor U12321 (N_12321,N_6500,N_7448);
nand U12322 (N_12322,N_6354,N_9219);
xor U12323 (N_12323,N_8394,N_7630);
and U12324 (N_12324,N_8584,N_8690);
or U12325 (N_12325,N_6262,N_7124);
or U12326 (N_12326,N_7661,N_8101);
and U12327 (N_12327,N_6361,N_8153);
xnor U12328 (N_12328,N_7596,N_7743);
xor U12329 (N_12329,N_8801,N_8551);
nand U12330 (N_12330,N_6710,N_7813);
nor U12331 (N_12331,N_8698,N_7369);
xnor U12332 (N_12332,N_7290,N_6561);
nor U12333 (N_12333,N_8172,N_9271);
and U12334 (N_12334,N_7567,N_9194);
and U12335 (N_12335,N_9316,N_9336);
nor U12336 (N_12336,N_7127,N_9253);
or U12337 (N_12337,N_7134,N_8085);
xor U12338 (N_12338,N_9233,N_8916);
or U12339 (N_12339,N_6764,N_6396);
nor U12340 (N_12340,N_9297,N_7231);
and U12341 (N_12341,N_8037,N_7472);
or U12342 (N_12342,N_8309,N_7542);
and U12343 (N_12343,N_7393,N_7164);
xor U12344 (N_12344,N_6834,N_9066);
or U12345 (N_12345,N_7267,N_7347);
xor U12346 (N_12346,N_8478,N_7697);
xor U12347 (N_12347,N_6779,N_6940);
and U12348 (N_12348,N_8153,N_9289);
or U12349 (N_12349,N_8510,N_6557);
xor U12350 (N_12350,N_7944,N_7644);
nand U12351 (N_12351,N_6777,N_7561);
and U12352 (N_12352,N_8474,N_6499);
xnor U12353 (N_12353,N_9284,N_7490);
or U12354 (N_12354,N_6580,N_7869);
nor U12355 (N_12355,N_7284,N_8558);
and U12356 (N_12356,N_8978,N_7957);
nor U12357 (N_12357,N_7901,N_9276);
or U12358 (N_12358,N_8261,N_7580);
nand U12359 (N_12359,N_6903,N_8067);
or U12360 (N_12360,N_6886,N_6936);
or U12361 (N_12361,N_7218,N_7947);
nand U12362 (N_12362,N_6425,N_6648);
xor U12363 (N_12363,N_9078,N_8616);
and U12364 (N_12364,N_7506,N_7565);
or U12365 (N_12365,N_9104,N_8063);
and U12366 (N_12366,N_7980,N_7977);
nand U12367 (N_12367,N_8815,N_8023);
xnor U12368 (N_12368,N_9321,N_8968);
xor U12369 (N_12369,N_8934,N_7523);
xor U12370 (N_12370,N_7367,N_7129);
and U12371 (N_12371,N_9157,N_8957);
nor U12372 (N_12372,N_7173,N_8795);
and U12373 (N_12373,N_8681,N_8142);
or U12374 (N_12374,N_9365,N_7623);
nor U12375 (N_12375,N_7675,N_7967);
xor U12376 (N_12376,N_8234,N_6609);
or U12377 (N_12377,N_8731,N_8410);
nor U12378 (N_12378,N_7363,N_7872);
nand U12379 (N_12379,N_9328,N_7420);
xor U12380 (N_12380,N_7671,N_7884);
xor U12381 (N_12381,N_7401,N_7299);
and U12382 (N_12382,N_7029,N_7145);
nand U12383 (N_12383,N_6475,N_7901);
or U12384 (N_12384,N_6438,N_7790);
xor U12385 (N_12385,N_8286,N_7699);
or U12386 (N_12386,N_6678,N_7163);
xnor U12387 (N_12387,N_6810,N_9279);
or U12388 (N_12388,N_8321,N_6392);
or U12389 (N_12389,N_7004,N_8176);
or U12390 (N_12390,N_8238,N_9086);
nor U12391 (N_12391,N_7538,N_8416);
xnor U12392 (N_12392,N_6679,N_8790);
or U12393 (N_12393,N_7609,N_6936);
or U12394 (N_12394,N_7133,N_9137);
and U12395 (N_12395,N_6403,N_7579);
xor U12396 (N_12396,N_7499,N_7071);
or U12397 (N_12397,N_6425,N_6832);
or U12398 (N_12398,N_8156,N_6733);
nor U12399 (N_12399,N_8242,N_7979);
or U12400 (N_12400,N_8271,N_6979);
and U12401 (N_12401,N_7573,N_8014);
or U12402 (N_12402,N_6383,N_8904);
and U12403 (N_12403,N_8896,N_8634);
nand U12404 (N_12404,N_8472,N_9310);
or U12405 (N_12405,N_9299,N_7267);
and U12406 (N_12406,N_9122,N_8963);
or U12407 (N_12407,N_7924,N_8214);
and U12408 (N_12408,N_6315,N_9329);
nor U12409 (N_12409,N_8431,N_7277);
xor U12410 (N_12410,N_8854,N_8981);
nand U12411 (N_12411,N_7521,N_7225);
nand U12412 (N_12412,N_7911,N_8425);
nor U12413 (N_12413,N_7839,N_7192);
xnor U12414 (N_12414,N_9280,N_6800);
or U12415 (N_12415,N_7517,N_9037);
xor U12416 (N_12416,N_9048,N_7901);
nor U12417 (N_12417,N_8698,N_7686);
xor U12418 (N_12418,N_8400,N_9040);
nor U12419 (N_12419,N_8288,N_7951);
and U12420 (N_12420,N_8686,N_8489);
nand U12421 (N_12421,N_6832,N_6690);
nor U12422 (N_12422,N_9330,N_6590);
and U12423 (N_12423,N_8966,N_6951);
nor U12424 (N_12424,N_8837,N_6504);
and U12425 (N_12425,N_6659,N_6521);
and U12426 (N_12426,N_9288,N_8867);
nand U12427 (N_12427,N_8967,N_7764);
nor U12428 (N_12428,N_7137,N_9367);
nor U12429 (N_12429,N_7399,N_7018);
xnor U12430 (N_12430,N_8339,N_7702);
nor U12431 (N_12431,N_8900,N_8971);
and U12432 (N_12432,N_7815,N_8168);
nor U12433 (N_12433,N_9102,N_7692);
and U12434 (N_12434,N_8535,N_8907);
xor U12435 (N_12435,N_7260,N_8549);
nor U12436 (N_12436,N_6309,N_7134);
xnor U12437 (N_12437,N_6692,N_7546);
or U12438 (N_12438,N_6704,N_7863);
and U12439 (N_12439,N_6339,N_6906);
xnor U12440 (N_12440,N_7118,N_7714);
nand U12441 (N_12441,N_9264,N_8582);
xnor U12442 (N_12442,N_7752,N_6494);
nor U12443 (N_12443,N_8373,N_7955);
or U12444 (N_12444,N_7361,N_9011);
and U12445 (N_12445,N_9195,N_6353);
nor U12446 (N_12446,N_6697,N_8382);
and U12447 (N_12447,N_7755,N_9036);
nand U12448 (N_12448,N_6381,N_8884);
nand U12449 (N_12449,N_9074,N_7467);
nand U12450 (N_12450,N_9058,N_7348);
nand U12451 (N_12451,N_7578,N_7385);
xor U12452 (N_12452,N_7306,N_8944);
and U12453 (N_12453,N_7253,N_7742);
nand U12454 (N_12454,N_9084,N_6401);
xnor U12455 (N_12455,N_7151,N_6790);
and U12456 (N_12456,N_7837,N_6850);
and U12457 (N_12457,N_8309,N_9250);
xor U12458 (N_12458,N_8910,N_6725);
nand U12459 (N_12459,N_8786,N_8770);
or U12460 (N_12460,N_6863,N_8340);
nor U12461 (N_12461,N_6778,N_9114);
nand U12462 (N_12462,N_6731,N_7824);
nor U12463 (N_12463,N_7179,N_7134);
nor U12464 (N_12464,N_7753,N_8940);
nor U12465 (N_12465,N_7311,N_7051);
xnor U12466 (N_12466,N_7432,N_7385);
nor U12467 (N_12467,N_7543,N_8113);
nor U12468 (N_12468,N_7823,N_7831);
or U12469 (N_12469,N_9343,N_7658);
xnor U12470 (N_12470,N_8016,N_6442);
xnor U12471 (N_12471,N_6965,N_7778);
nand U12472 (N_12472,N_8206,N_7027);
or U12473 (N_12473,N_6519,N_6551);
nand U12474 (N_12474,N_8333,N_6890);
xnor U12475 (N_12475,N_6949,N_6766);
nand U12476 (N_12476,N_7034,N_8095);
nor U12477 (N_12477,N_7521,N_8496);
nor U12478 (N_12478,N_8577,N_8069);
nand U12479 (N_12479,N_6515,N_7641);
nor U12480 (N_12480,N_7788,N_8379);
or U12481 (N_12481,N_6812,N_7474);
and U12482 (N_12482,N_7069,N_7147);
or U12483 (N_12483,N_8374,N_7983);
and U12484 (N_12484,N_8968,N_7798);
nor U12485 (N_12485,N_8965,N_6428);
nor U12486 (N_12486,N_7258,N_8722);
xnor U12487 (N_12487,N_7092,N_8814);
xnor U12488 (N_12488,N_7381,N_7700);
and U12489 (N_12489,N_7629,N_6753);
nor U12490 (N_12490,N_9053,N_8498);
nor U12491 (N_12491,N_6929,N_6478);
xor U12492 (N_12492,N_7123,N_6309);
nor U12493 (N_12493,N_7937,N_7580);
or U12494 (N_12494,N_7805,N_7572);
and U12495 (N_12495,N_6746,N_7407);
and U12496 (N_12496,N_6308,N_6763);
or U12497 (N_12497,N_6823,N_9281);
xnor U12498 (N_12498,N_8766,N_7991);
xor U12499 (N_12499,N_6378,N_9019);
nand U12500 (N_12500,N_10136,N_11171);
xnor U12501 (N_12501,N_10143,N_12163);
and U12502 (N_12502,N_10132,N_11798);
xor U12503 (N_12503,N_10823,N_12279);
nand U12504 (N_12504,N_10507,N_10374);
and U12505 (N_12505,N_10127,N_10742);
nor U12506 (N_12506,N_9696,N_11285);
nand U12507 (N_12507,N_10299,N_10863);
xor U12508 (N_12508,N_11206,N_10666);
and U12509 (N_12509,N_10326,N_11048);
and U12510 (N_12510,N_12066,N_11409);
nand U12511 (N_12511,N_10748,N_10777);
and U12512 (N_12512,N_9978,N_9384);
xnor U12513 (N_12513,N_9428,N_9891);
nor U12514 (N_12514,N_12491,N_11541);
nand U12515 (N_12515,N_10663,N_10112);
and U12516 (N_12516,N_10256,N_9602);
nand U12517 (N_12517,N_11888,N_10486);
and U12518 (N_12518,N_11913,N_10675);
nor U12519 (N_12519,N_10449,N_11464);
and U12520 (N_12520,N_10971,N_10684);
or U12521 (N_12521,N_11901,N_9753);
or U12522 (N_12522,N_10338,N_11963);
xnor U12523 (N_12523,N_11507,N_11069);
or U12524 (N_12524,N_9451,N_10314);
nand U12525 (N_12525,N_10910,N_12299);
and U12526 (N_12526,N_10153,N_11329);
nor U12527 (N_12527,N_11619,N_10414);
and U12528 (N_12528,N_11166,N_10465);
nand U12529 (N_12529,N_11735,N_11718);
and U12530 (N_12530,N_11013,N_10159);
nor U12531 (N_12531,N_9932,N_11761);
or U12532 (N_12532,N_9824,N_11969);
nor U12533 (N_12533,N_10196,N_10805);
and U12534 (N_12534,N_10827,N_10852);
or U12535 (N_12535,N_10339,N_11425);
or U12536 (N_12536,N_9426,N_10081);
or U12537 (N_12537,N_12119,N_11402);
or U12538 (N_12538,N_11840,N_10040);
and U12539 (N_12539,N_12339,N_12274);
or U12540 (N_12540,N_9547,N_11485);
xnor U12541 (N_12541,N_12382,N_9414);
and U12542 (N_12542,N_12071,N_11964);
or U12543 (N_12543,N_11449,N_12004);
nand U12544 (N_12544,N_11799,N_9745);
and U12545 (N_12545,N_9702,N_10526);
and U12546 (N_12546,N_10301,N_10025);
xor U12547 (N_12547,N_11232,N_12286);
nand U12548 (N_12548,N_12414,N_10458);
or U12549 (N_12549,N_9560,N_12175);
and U12550 (N_12550,N_11648,N_9876);
xor U12551 (N_12551,N_9858,N_10698);
and U12552 (N_12552,N_9959,N_9375);
nor U12553 (N_12553,N_10382,N_10445);
and U12554 (N_12554,N_12022,N_12122);
nand U12555 (N_12555,N_10415,N_10924);
nor U12556 (N_12556,N_11219,N_9862);
or U12557 (N_12557,N_10430,N_11986);
and U12558 (N_12558,N_11336,N_11008);
nand U12559 (N_12559,N_9416,N_10419);
or U12560 (N_12560,N_9864,N_11486);
xor U12561 (N_12561,N_12160,N_9831);
nor U12562 (N_12562,N_11245,N_10751);
nor U12563 (N_12563,N_11583,N_11481);
and U12564 (N_12564,N_11623,N_10831);
or U12565 (N_12565,N_10718,N_11500);
or U12566 (N_12566,N_10918,N_11601);
or U12567 (N_12567,N_9851,N_9387);
xor U12568 (N_12568,N_9513,N_12306);
nor U12569 (N_12569,N_11439,N_10131);
and U12570 (N_12570,N_9798,N_11461);
xor U12571 (N_12571,N_11027,N_9405);
or U12572 (N_12572,N_11706,N_9472);
xnor U12573 (N_12573,N_9915,N_11243);
xnor U12574 (N_12574,N_11612,N_9939);
and U12575 (N_12575,N_12124,N_10200);
nor U12576 (N_12576,N_10251,N_9742);
xnor U12577 (N_12577,N_11792,N_9713);
nand U12578 (N_12578,N_11607,N_9811);
or U12579 (N_12579,N_11104,N_12179);
xor U12580 (N_12580,N_9682,N_12287);
nor U12581 (N_12581,N_10769,N_11933);
xor U12582 (N_12582,N_10287,N_11427);
nand U12583 (N_12583,N_10460,N_10692);
xor U12584 (N_12584,N_11094,N_11899);
and U12585 (N_12585,N_10000,N_11652);
or U12586 (N_12586,N_11590,N_11633);
nor U12587 (N_12587,N_9872,N_11517);
nand U12588 (N_12588,N_11711,N_10013);
nor U12589 (N_12589,N_10803,N_12009);
nor U12590 (N_12590,N_11223,N_11044);
and U12591 (N_12591,N_11119,N_11925);
xnor U12592 (N_12592,N_11004,N_9927);
nor U12593 (N_12593,N_10295,N_11558);
xnor U12594 (N_12594,N_11781,N_10404);
nand U12595 (N_12595,N_11830,N_9608);
or U12596 (N_12596,N_10423,N_11836);
or U12597 (N_12597,N_10068,N_11542);
or U12598 (N_12598,N_10793,N_10425);
nand U12599 (N_12599,N_11802,N_9512);
xnor U12600 (N_12600,N_9531,N_11688);
nor U12601 (N_12601,N_11091,N_11155);
and U12602 (N_12602,N_11351,N_11671);
nor U12603 (N_12603,N_10631,N_10342);
xnor U12604 (N_12604,N_11992,N_12005);
nand U12605 (N_12605,N_9800,N_9543);
and U12606 (N_12606,N_9817,N_12407);
nor U12607 (N_12607,N_11084,N_12152);
xor U12608 (N_12608,N_9625,N_10491);
nand U12609 (N_12609,N_10058,N_10291);
nand U12610 (N_12610,N_11824,N_9635);
nor U12611 (N_12611,N_11366,N_11545);
nand U12612 (N_12612,N_12358,N_11376);
xnor U12613 (N_12613,N_11229,N_11076);
or U12614 (N_12614,N_11935,N_12224);
xnor U12615 (N_12615,N_10420,N_9486);
nand U12616 (N_12616,N_10847,N_11357);
xnor U12617 (N_12617,N_10222,N_9407);
nand U12618 (N_12618,N_12200,N_10026);
or U12619 (N_12619,N_12108,N_10481);
nor U12620 (N_12620,N_11551,N_10714);
and U12621 (N_12621,N_10786,N_11502);
nand U12622 (N_12622,N_10529,N_10286);
or U12623 (N_12623,N_11710,N_11478);
or U12624 (N_12624,N_10266,N_11239);
nand U12625 (N_12625,N_10494,N_10257);
and U12626 (N_12626,N_10498,N_11121);
or U12627 (N_12627,N_11509,N_12261);
xnor U12628 (N_12628,N_11360,N_11947);
and U12629 (N_12629,N_12297,N_10588);
or U12630 (N_12630,N_12390,N_10681);
nand U12631 (N_12631,N_11544,N_9985);
nor U12632 (N_12632,N_10701,N_10145);
and U12633 (N_12633,N_11730,N_11505);
or U12634 (N_12634,N_9620,N_10783);
xor U12635 (N_12635,N_10995,N_11184);
or U12636 (N_12636,N_11283,N_11864);
xnor U12637 (N_12637,N_10580,N_10792);
nand U12638 (N_12638,N_11897,N_10208);
or U12639 (N_12639,N_9609,N_11661);
xor U12640 (N_12640,N_11204,N_10613);
nand U12641 (N_12641,N_9920,N_9669);
nor U12642 (N_12642,N_10424,N_11929);
and U12643 (N_12643,N_10281,N_10697);
and U12644 (N_12644,N_9503,N_10987);
or U12645 (N_12645,N_10632,N_9413);
and U12646 (N_12646,N_10587,N_9878);
and U12647 (N_12647,N_11705,N_12000);
nor U12648 (N_12648,N_11158,N_9564);
and U12649 (N_12649,N_12276,N_9589);
nor U12650 (N_12650,N_10292,N_11668);
or U12651 (N_12651,N_11317,N_10214);
xnor U12652 (N_12652,N_11407,N_11555);
xnor U12653 (N_12653,N_10871,N_9728);
xnor U12654 (N_12654,N_10252,N_11403);
xnor U12655 (N_12655,N_10870,N_9619);
or U12656 (N_12656,N_12443,N_11404);
or U12657 (N_12657,N_9970,N_9890);
xor U12658 (N_12658,N_11755,N_10340);
nand U12659 (N_12659,N_11809,N_12336);
and U12660 (N_12660,N_11919,N_10774);
and U12661 (N_12661,N_12155,N_9983);
nor U12662 (N_12662,N_9710,N_10398);
or U12663 (N_12663,N_10213,N_12125);
nor U12664 (N_12664,N_10259,N_10215);
and U12665 (N_12665,N_11090,N_11041);
or U12666 (N_12666,N_12035,N_11884);
xor U12667 (N_12667,N_10485,N_10006);
nor U12668 (N_12668,N_11102,N_12054);
nor U12669 (N_12669,N_11458,N_12393);
xor U12670 (N_12670,N_12247,N_10380);
nor U12671 (N_12671,N_11335,N_11006);
and U12672 (N_12672,N_11079,N_9390);
xor U12673 (N_12673,N_11754,N_10097);
nor U12674 (N_12674,N_9965,N_11578);
or U12675 (N_12675,N_12476,N_12027);
and U12676 (N_12676,N_9847,N_10316);
nand U12677 (N_12677,N_9442,N_9929);
nor U12678 (N_12678,N_10216,N_12295);
xor U12679 (N_12679,N_9552,N_9925);
xnor U12680 (N_12680,N_12191,N_12199);
nand U12681 (N_12681,N_9490,N_11430);
or U12682 (N_12682,N_12241,N_11020);
nand U12683 (N_12683,N_11334,N_12383);
or U12684 (N_12684,N_9875,N_10297);
nor U12685 (N_12685,N_11131,N_12314);
and U12686 (N_12686,N_9509,N_10789);
nand U12687 (N_12687,N_11882,N_12138);
nand U12688 (N_12688,N_11617,N_11181);
nand U12689 (N_12689,N_11138,N_9991);
nor U12690 (N_12690,N_11442,N_10393);
xnor U12691 (N_12691,N_12112,N_10436);
nor U12692 (N_12692,N_9377,N_9928);
nand U12693 (N_12693,N_10590,N_9764);
and U12694 (N_12694,N_11423,N_11891);
or U12695 (N_12695,N_11391,N_12292);
nand U12696 (N_12696,N_10996,N_12073);
xor U12697 (N_12697,N_10061,N_10035);
and U12698 (N_12698,N_10344,N_10978);
nor U12699 (N_12699,N_12088,N_9952);
xor U12700 (N_12700,N_9990,N_9896);
and U12701 (N_12701,N_11364,N_9954);
or U12702 (N_12702,N_9703,N_11087);
xor U12703 (N_12703,N_9685,N_9456);
and U12704 (N_12704,N_11962,N_9586);
or U12705 (N_12705,N_10915,N_9395);
xor U12706 (N_12706,N_11807,N_12114);
nor U12707 (N_12707,N_9699,N_10411);
nand U12708 (N_12708,N_9461,N_10676);
nand U12709 (N_12709,N_12006,N_12354);
nand U12710 (N_12710,N_11172,N_10662);
xnor U12711 (N_12711,N_10290,N_9856);
xor U12712 (N_12712,N_10403,N_12485);
xor U12713 (N_12713,N_9722,N_12281);
nor U12714 (N_12714,N_10717,N_10988);
nor U12715 (N_12715,N_9849,N_11534);
or U12716 (N_12716,N_10857,N_10902);
or U12717 (N_12717,N_9680,N_11942);
nand U12718 (N_12718,N_11866,N_10079);
xor U12719 (N_12719,N_10148,N_11527);
nor U12720 (N_12720,N_11995,N_10302);
or U12721 (N_12721,N_11007,N_12334);
nand U12722 (N_12722,N_10934,N_10602);
nand U12723 (N_12723,N_10352,N_12260);
and U12724 (N_12724,N_11985,N_10320);
nand U12725 (N_12725,N_9828,N_9599);
and U12726 (N_12726,N_12194,N_11117);
and U12727 (N_12727,N_11021,N_10582);
or U12728 (N_12728,N_11740,N_12310);
nor U12729 (N_12729,N_9907,N_11565);
nor U12730 (N_12730,N_9711,N_11530);
xnor U12731 (N_12731,N_10219,N_11737);
or U12732 (N_12732,N_10188,N_11700);
or U12733 (N_12733,N_12030,N_11050);
or U12734 (N_12734,N_10730,N_9692);
nand U12735 (N_12735,N_12141,N_11703);
and U12736 (N_12736,N_9664,N_11715);
nand U12737 (N_12737,N_12494,N_11354);
and U12738 (N_12738,N_12068,N_10607);
and U12739 (N_12739,N_11297,N_11723);
or U12740 (N_12740,N_10885,N_11215);
nand U12741 (N_12741,N_11422,N_10550);
and U12742 (N_12742,N_10401,N_10307);
nor U12743 (N_12743,N_11915,N_10770);
nand U12744 (N_12744,N_10203,N_9600);
and U12745 (N_12745,N_10348,N_10811);
or U12746 (N_12746,N_11902,N_12202);
xor U12747 (N_12747,N_11605,N_9986);
nand U12748 (N_12748,N_10802,N_9726);
and U12749 (N_12749,N_11046,N_11454);
nor U12750 (N_12750,N_12015,N_10379);
xor U12751 (N_12751,N_10113,N_11061);
or U12752 (N_12752,N_11878,N_12062);
and U12753 (N_12753,N_11450,N_11295);
nand U12754 (N_12754,N_11787,N_12469);
nand U12755 (N_12755,N_9758,N_12461);
or U12756 (N_12756,N_9638,N_9510);
nand U12757 (N_12757,N_9755,N_11663);
or U12758 (N_12758,N_9701,N_10821);
xnor U12759 (N_12759,N_11865,N_10914);
xnor U12760 (N_12760,N_11849,N_11697);
xor U12761 (N_12761,N_10819,N_11637);
or U12762 (N_12762,N_9623,N_11345);
xnor U12763 (N_12763,N_11326,N_9947);
xor U12764 (N_12764,N_10033,N_9737);
xnor U12765 (N_12765,N_11525,N_11072);
and U12766 (N_12766,N_11524,N_12498);
or U12767 (N_12767,N_12198,N_9740);
nor U12768 (N_12768,N_12057,N_11523);
nor U12769 (N_12769,N_9652,N_10270);
and U12770 (N_12770,N_11681,N_11032);
nand U12771 (N_12771,N_11018,N_11940);
xor U12772 (N_12772,N_10750,N_10381);
nand U12773 (N_12773,N_9893,N_10179);
nor U12774 (N_12774,N_11214,N_10755);
and U12775 (N_12775,N_11490,N_9457);
nand U12776 (N_12776,N_10480,N_10387);
or U12777 (N_12777,N_11033,N_10965);
nor U12778 (N_12778,N_9819,N_9805);
and U12779 (N_12779,N_9671,N_10199);
and U12780 (N_12780,N_9649,N_9629);
nor U12781 (N_12781,N_12103,N_10759);
nor U12782 (N_12782,N_10711,N_10435);
nor U12783 (N_12783,N_11029,N_12365);
nor U12784 (N_12784,N_9541,N_10186);
nor U12785 (N_12785,N_10482,N_9628);
nor U12786 (N_12786,N_10739,N_10416);
nor U12787 (N_12787,N_10408,N_9980);
nor U12788 (N_12788,N_10609,N_10853);
or U12789 (N_12789,N_11968,N_9443);
nand U12790 (N_12790,N_11352,N_10462);
and U12791 (N_12791,N_10654,N_11741);
or U12792 (N_12792,N_9977,N_12203);
nor U12793 (N_12793,N_10010,N_12169);
and U12794 (N_12794,N_10469,N_9409);
or U12795 (N_12795,N_10327,N_11961);
xnor U12796 (N_12796,N_11991,N_11596);
or U12797 (N_12797,N_11197,N_11320);
nor U12798 (N_12798,N_10126,N_9850);
nor U12799 (N_12799,N_11954,N_11479);
xnor U12800 (N_12800,N_11977,N_11476);
and U12801 (N_12801,N_10323,N_11379);
nand U12802 (N_12802,N_11332,N_11395);
xnor U12803 (N_12803,N_10710,N_11952);
xnor U12804 (N_12804,N_9691,N_9873);
and U12805 (N_12805,N_9597,N_9658);
nor U12806 (N_12806,N_9749,N_12416);
and U12807 (N_12807,N_10936,N_11687);
xnor U12808 (N_12808,N_10604,N_12167);
or U12809 (N_12809,N_10734,N_12465);
nand U12810 (N_12810,N_11508,N_10896);
or U12811 (N_12811,N_10984,N_10390);
or U12812 (N_12812,N_9505,N_10052);
or U12813 (N_12813,N_11562,N_9787);
or U12814 (N_12814,N_10736,N_9842);
nand U12815 (N_12815,N_11222,N_10558);
and U12816 (N_12816,N_12413,N_9859);
nand U12817 (N_12817,N_9690,N_10262);
xor U12818 (N_12818,N_10667,N_11938);
or U12819 (N_12819,N_12178,N_11746);
or U12820 (N_12820,N_10646,N_12322);
xnor U12821 (N_12821,N_10837,N_12077);
xnor U12822 (N_12822,N_11945,N_10439);
and U12823 (N_12823,N_11709,N_12033);
nor U12824 (N_12824,N_9942,N_12262);
xnor U12825 (N_12825,N_11532,N_9822);
xor U12826 (N_12826,N_10118,N_11003);
nand U12827 (N_12827,N_11850,N_10042);
nand U12828 (N_12828,N_10804,N_11627);
and U12829 (N_12829,N_9791,N_9386);
nor U12830 (N_12830,N_12176,N_12359);
nor U12831 (N_12831,N_12143,N_9795);
or U12832 (N_12832,N_11751,N_9526);
xor U12833 (N_12833,N_11719,N_10376);
and U12834 (N_12834,N_10372,N_11895);
or U12835 (N_12835,N_11910,N_9921);
xor U12836 (N_12836,N_10832,N_9941);
xnor U12837 (N_12837,N_12184,N_12238);
nand U12838 (N_12838,N_10011,N_10970);
nand U12839 (N_12839,N_10559,N_9829);
nand U12840 (N_12840,N_11135,N_9561);
nand U12841 (N_12841,N_11990,N_10660);
nand U12842 (N_12842,N_10331,N_12438);
and U12843 (N_12843,N_11831,N_12089);
nor U12844 (N_12844,N_11296,N_12425);
and U12845 (N_12845,N_11881,N_9466);
and U12846 (N_12846,N_12135,N_11274);
and U12847 (N_12847,N_11062,N_12266);
and U12848 (N_12848,N_12316,N_9951);
xor U12849 (N_12849,N_11024,N_12228);
xor U12850 (N_12850,N_11670,N_11624);
xor U12851 (N_12851,N_12237,N_9523);
nor U12852 (N_12852,N_10767,N_12126);
or U12853 (N_12853,N_11150,N_10472);
nor U12854 (N_12854,N_11970,N_12258);
and U12855 (N_12855,N_10434,N_9821);
or U12856 (N_12856,N_11616,N_10221);
nor U12857 (N_12857,N_10232,N_11047);
or U12858 (N_12858,N_11002,N_9746);
nand U12859 (N_12859,N_10045,N_11444);
nor U12860 (N_12860,N_10239,N_10116);
nor U12861 (N_12861,N_11516,N_12154);
and U12862 (N_12862,N_11389,N_11659);
and U12863 (N_12863,N_9981,N_11160);
and U12864 (N_12864,N_11293,N_10838);
xnor U12865 (N_12865,N_10004,N_10694);
xor U12866 (N_12866,N_11622,N_11557);
nand U12867 (N_12867,N_10926,N_11328);
nor U12868 (N_12868,N_9885,N_10014);
nand U12869 (N_12869,N_11063,N_9415);
or U12870 (N_12870,N_11381,N_11739);
and U12871 (N_12871,N_10022,N_9818);
or U12872 (N_12872,N_11981,N_10083);
nor U12873 (N_12873,N_9793,N_10540);
or U12874 (N_12874,N_11122,N_10160);
or U12875 (N_12875,N_9580,N_10377);
xnor U12876 (N_12876,N_11385,N_12337);
xor U12877 (N_12877,N_10303,N_9471);
xor U12878 (N_12878,N_9975,N_9611);
and U12879 (N_12879,N_9883,N_11136);
or U12880 (N_12880,N_11598,N_10095);
nand U12881 (N_12881,N_10848,N_10842);
or U12882 (N_12882,N_11113,N_11585);
or U12883 (N_12883,N_11521,N_12134);
nand U12884 (N_12884,N_12378,N_11763);
or U12885 (N_12885,N_9478,N_12284);
or U12886 (N_12886,N_11716,N_12075);
nand U12887 (N_12887,N_10596,N_9430);
or U12888 (N_12888,N_11009,N_12102);
xor U12889 (N_12889,N_12092,N_11307);
or U12890 (N_12890,N_10993,N_9796);
or U12891 (N_12891,N_11399,N_11561);
nand U12892 (N_12892,N_9794,N_10181);
nor U12893 (N_12893,N_10016,N_12177);
and U12894 (N_12894,N_10989,N_12457);
nand U12895 (N_12895,N_9650,N_10241);
and U12896 (N_12896,N_11839,N_10183);
and U12897 (N_12897,N_11340,N_12217);
and U12898 (N_12898,N_9957,N_10610);
xor U12899 (N_12899,N_10413,N_11370);
nor U12900 (N_12900,N_9606,N_12423);
nor U12901 (N_12901,N_12479,N_10198);
nor U12902 (N_12902,N_12251,N_9744);
or U12903 (N_12903,N_12166,N_11811);
xnor U12904 (N_12904,N_11410,N_9630);
xnor U12905 (N_12905,N_12142,N_11804);
xnor U12906 (N_12906,N_11777,N_12308);
xnor U12907 (N_12907,N_10364,N_10619);
nand U12908 (N_12908,N_12150,N_11513);
or U12909 (N_12909,N_12347,N_10353);
xor U12910 (N_12910,N_9714,N_12484);
nor U12911 (N_12911,N_11808,N_9730);
nor U12912 (N_12912,N_10828,N_11996);
or U12913 (N_12913,N_10901,N_11209);
nor U12914 (N_12914,N_11914,N_11789);
or U12915 (N_12915,N_12473,N_11635);
and U12916 (N_12916,N_12415,N_9889);
and U12917 (N_12917,N_12078,N_12424);
nor U12918 (N_12918,N_11756,N_11109);
nor U12919 (N_12919,N_11058,N_9960);
xor U12920 (N_12920,N_11658,N_11495);
or U12921 (N_12921,N_12355,N_12478);
or U12922 (N_12922,N_9752,N_9935);
nor U12923 (N_12923,N_10650,N_9768);
nor U12924 (N_12924,N_10467,N_11800);
and U12925 (N_12925,N_12495,N_12361);
xor U12926 (N_12926,N_9429,N_11520);
or U12927 (N_12927,N_10606,N_11934);
xor U12928 (N_12928,N_11618,N_10069);
nor U12929 (N_12929,N_11080,N_12385);
nor U12930 (N_12930,N_12488,N_9901);
nand U12931 (N_12931,N_12253,N_11828);
xor U12932 (N_12932,N_9487,N_11489);
nor U12933 (N_12933,N_11569,N_10373);
nand U12934 (N_12934,N_10253,N_10383);
nand U12935 (N_12935,N_10564,N_10905);
or U12936 (N_12936,N_10615,N_9496);
and U12937 (N_12937,N_10608,N_10101);
or U12938 (N_12938,N_11957,N_9581);
and U12939 (N_12939,N_11776,N_10939);
xor U12940 (N_12940,N_9514,N_11116);
xor U12941 (N_12941,N_12149,N_10844);
nor U12942 (N_12942,N_11241,N_10579);
nand U12943 (N_12943,N_10788,N_11497);
nor U12944 (N_12944,N_10378,N_11178);
nand U12945 (N_12945,N_10685,N_9666);
nor U12946 (N_12946,N_11564,N_10626);
and U12947 (N_12947,N_11504,N_9607);
nand U12948 (N_12948,N_12146,N_12375);
or U12949 (N_12949,N_11156,N_10573);
xnor U12950 (N_12950,N_9868,N_9874);
xnor U12951 (N_12951,N_9610,N_10433);
xnor U12952 (N_12952,N_10651,N_11124);
and U12953 (N_12953,N_10167,N_10688);
nor U12954 (N_12954,N_10953,N_11640);
xnor U12955 (N_12955,N_12411,N_11343);
nand U12956 (N_12956,N_10900,N_10785);
nand U12957 (N_12957,N_11436,N_10636);
nor U12958 (N_12958,N_9784,N_12209);
or U12959 (N_12959,N_10845,N_11134);
nor U12960 (N_12960,N_11330,N_10992);
nor U12961 (N_12961,N_10727,N_9731);
xor U12962 (N_12962,N_12113,N_12220);
xor U12963 (N_12963,N_9439,N_9860);
nand U12964 (N_12964,N_9447,N_11108);
nand U12965 (N_12965,N_12213,N_9905);
nor U12966 (N_12966,N_9887,N_10909);
and U12967 (N_12967,N_11456,N_11695);
or U12968 (N_12968,N_9903,N_10128);
nor U12969 (N_12969,N_12181,N_11783);
and U12970 (N_12970,N_9984,N_11429);
and U12971 (N_12971,N_11547,N_9553);
and U12972 (N_12972,N_11488,N_10665);
or U12973 (N_12973,N_10043,N_11528);
nand U12974 (N_12974,N_9397,N_9879);
nor U12975 (N_12975,N_10191,N_10109);
xnor U12976 (N_12976,N_9425,N_10977);
or U12977 (N_12977,N_10410,N_11795);
and U12978 (N_12978,N_10599,N_10152);
or U12979 (N_12979,N_12395,N_11055);
and U12980 (N_12980,N_11342,N_10806);
or U12981 (N_12981,N_10696,N_9605);
or U12982 (N_12982,N_11279,N_10051);
nand U12983 (N_12983,N_11543,N_10237);
nand U12984 (N_12984,N_12435,N_10672);
or U12985 (N_12985,N_11593,N_9441);
or U12986 (N_12986,N_10272,N_9732);
and U12987 (N_12987,N_12061,N_10343);
nor U12988 (N_12988,N_10094,N_12214);
and U12989 (N_12989,N_9914,N_10567);
xor U12990 (N_12990,N_9555,N_10204);
or U12991 (N_12991,N_11437,N_10029);
nor U12992 (N_12992,N_9463,N_9644);
nor U12993 (N_12993,N_12448,N_11227);
nand U12994 (N_12994,N_12335,N_10557);
nand U12995 (N_12995,N_11603,N_10210);
nand U12996 (N_12996,N_9618,N_12246);
nand U12997 (N_12997,N_10431,N_12028);
and U12998 (N_12998,N_9974,N_10864);
or U12999 (N_12999,N_11714,N_10859);
xor U13000 (N_13000,N_10085,N_10880);
nand U13001 (N_13001,N_11315,N_9540);
nor U13002 (N_13002,N_10723,N_11841);
xnor U13003 (N_13003,N_9404,N_10501);
or U13004 (N_13004,N_11236,N_10225);
nand U13005 (N_13005,N_11322,N_11473);
or U13006 (N_13006,N_10243,N_11958);
or U13007 (N_13007,N_11704,N_10547);
and U13008 (N_13008,N_12187,N_11531);
nand U13009 (N_13009,N_11088,N_9511);
or U13010 (N_13010,N_12327,N_11732);
and U13011 (N_13011,N_9743,N_11501);
and U13012 (N_13012,N_10598,N_10284);
nand U13013 (N_13013,N_11920,N_10648);
or U13014 (N_13014,N_9958,N_10600);
or U13015 (N_13015,N_10120,N_9396);
nand U13016 (N_13016,N_11941,N_12242);
or U13017 (N_13017,N_9759,N_11696);
and U13018 (N_13018,N_11482,N_10178);
nor U13019 (N_13019,N_10594,N_11825);
nor U13020 (N_13020,N_9961,N_9533);
xnor U13021 (N_13021,N_11282,N_11321);
and U13022 (N_13022,N_10780,N_9467);
and U13023 (N_13023,N_9801,N_10964);
nand U13024 (N_13024,N_11689,N_12085);
and U13025 (N_13025,N_9551,N_11903);
xnor U13026 (N_13026,N_12055,N_9908);
or U13027 (N_13027,N_9762,N_10495);
nor U13028 (N_13028,N_12456,N_11589);
or U13029 (N_13029,N_11075,N_10499);
xor U13030 (N_13030,N_9723,N_12330);
xnor U13031 (N_13031,N_12192,N_11867);
nor U13032 (N_13032,N_11522,N_10056);
or U13033 (N_13033,N_11349,N_11550);
and U13034 (N_13034,N_11278,N_10207);
nand U13035 (N_13035,N_11951,N_10855);
xor U13036 (N_13036,N_12263,N_11054);
xor U13037 (N_13037,N_10768,N_10240);
xnor U13038 (N_13038,N_12388,N_11650);
nand U13039 (N_13039,N_12309,N_12344);
or U13040 (N_13040,N_9633,N_11014);
and U13041 (N_13041,N_9763,N_11175);
and U13042 (N_13042,N_11397,N_11731);
and U13043 (N_13043,N_10277,N_10757);
or U13044 (N_13044,N_10879,N_10913);
nor U13045 (N_13045,N_10076,N_12373);
or U13046 (N_13046,N_10409,N_10071);
nor U13047 (N_13047,N_9481,N_10358);
xor U13048 (N_13048,N_9861,N_10997);
or U13049 (N_13049,N_10223,N_9453);
xor U13050 (N_13050,N_9988,N_10994);
and U13051 (N_13051,N_9612,N_10474);
nand U13052 (N_13052,N_10511,N_10089);
and U13053 (N_13053,N_10715,N_10930);
and U13054 (N_13054,N_12399,N_10775);
and U13055 (N_13055,N_11179,N_11844);
nand U13056 (N_13056,N_12049,N_9734);
xnor U13057 (N_13057,N_10018,N_9820);
or U13058 (N_13058,N_10799,N_9909);
nor U13059 (N_13059,N_10315,N_12256);
nor U13060 (N_13060,N_11560,N_10903);
nor U13061 (N_13061,N_11827,N_12319);
nand U13062 (N_13062,N_11842,N_10937);
and U13063 (N_13063,N_9799,N_9483);
nor U13064 (N_13064,N_11979,N_9529);
nand U13065 (N_13065,N_10639,N_9641);
nor U13066 (N_13066,N_10119,N_12046);
or U13067 (N_13067,N_11380,N_9530);
nor U13068 (N_13068,N_11647,N_10361);
or U13069 (N_13069,N_10235,N_9845);
and U13070 (N_13070,N_9698,N_12267);
or U13071 (N_13071,N_10513,N_11738);
nand U13072 (N_13072,N_10180,N_10577);
xnor U13073 (N_13073,N_10657,N_10744);
nor U13074 (N_13074,N_12227,N_12379);
nor U13075 (N_13075,N_11133,N_10421);
xnor U13076 (N_13076,N_10418,N_12031);
or U13077 (N_13077,N_12007,N_10005);
xor U13078 (N_13078,N_10976,N_9528);
nand U13079 (N_13079,N_12362,N_12168);
xnor U13080 (N_13080,N_11465,N_11806);
nor U13081 (N_13081,N_12161,N_12120);
xor U13082 (N_13082,N_10493,N_10060);
xor U13083 (N_13083,N_10166,N_12447);
or U13084 (N_13084,N_10135,N_11115);
nand U13085 (N_13085,N_12278,N_10945);
or U13086 (N_13086,N_9972,N_12436);
and U13087 (N_13087,N_11118,N_9432);
or U13088 (N_13088,N_12182,N_10479);
and U13089 (N_13089,N_10535,N_10999);
nor U13090 (N_13090,N_9852,N_10618);
or U13091 (N_13091,N_11540,N_10951);
or U13092 (N_13092,N_10981,N_10090);
nand U13093 (N_13093,N_11769,N_12480);
and U13094 (N_13094,N_10904,N_10749);
xnor U13095 (N_13095,N_10980,N_9537);
nor U13096 (N_13096,N_9400,N_12272);
or U13097 (N_13097,N_12173,N_10527);
nand U13098 (N_13098,N_9807,N_12127);
nor U13099 (N_13099,N_10274,N_9445);
nand U13100 (N_13100,N_9709,N_11031);
and U13101 (N_13101,N_11858,N_10630);
nand U13102 (N_13102,N_10882,N_10790);
and U13103 (N_13103,N_11499,N_10002);
xor U13104 (N_13104,N_10952,N_11471);
or U13105 (N_13105,N_9962,N_11448);
and U13106 (N_13106,N_9645,N_10772);
nand U13107 (N_13107,N_10898,N_11099);
nor U13108 (N_13108,N_11801,N_11161);
nand U13109 (N_13109,N_12298,N_11683);
nand U13110 (N_13110,N_11142,N_10745);
or U13111 (N_13111,N_10625,N_9489);
nor U13112 (N_13112,N_10894,N_11931);
nor U13113 (N_13113,N_10078,N_11860);
and U13114 (N_13114,N_12240,N_9631);
xnor U13115 (N_13115,N_9527,N_10658);
xnor U13116 (N_13116,N_10949,N_10400);
or U13117 (N_13117,N_11821,N_10062);
nor U13118 (N_13118,N_10812,N_10743);
or U13119 (N_13119,N_9672,N_9614);
nand U13120 (N_13120,N_10721,N_10268);
nor U13121 (N_13121,N_9693,N_11774);
nor U13122 (N_13122,N_11724,N_11625);
and U13123 (N_13123,N_11924,N_10687);
nand U13124 (N_13124,N_10979,N_10623);
and U13125 (N_13125,N_12107,N_11272);
xor U13126 (N_13126,N_10887,N_10333);
and U13127 (N_13127,N_10304,N_10548);
nand U13128 (N_13128,N_9747,N_9916);
nand U13129 (N_13129,N_10968,N_11868);
and U13130 (N_13130,N_10155,N_10928);
and U13131 (N_13131,N_11611,N_9697);
xor U13132 (N_13132,N_11000,N_10556);
nand U13133 (N_13133,N_10708,N_10265);
or U13134 (N_13134,N_9781,N_12025);
nor U13135 (N_13135,N_11674,N_10086);
nor U13136 (N_13136,N_11812,N_10982);
xnor U13137 (N_13137,N_12421,N_10412);
and U13138 (N_13138,N_11675,N_12233);
or U13139 (N_13139,N_12056,N_11292);
nand U13140 (N_13140,N_9622,N_12003);
xnor U13141 (N_13141,N_9782,N_10671);
nor U13142 (N_13142,N_10144,N_10202);
nand U13143 (N_13143,N_9886,N_10758);
nor U13144 (N_13144,N_11128,N_9689);
xor U13145 (N_13145,N_11426,N_11235);
xor U13146 (N_13146,N_9834,N_10712);
nand U13147 (N_13147,N_9468,N_10897);
or U13148 (N_13148,N_9495,N_11265);
nand U13149 (N_13149,N_9906,N_12384);
nor U13150 (N_13150,N_11813,N_9474);
nor U13151 (N_13151,N_10990,N_9388);
nand U13152 (N_13152,N_11462,N_10146);
nand U13153 (N_13153,N_12304,N_12463);
nor U13154 (N_13154,N_9516,N_11226);
nand U13155 (N_13155,N_9704,N_10746);
and U13156 (N_13156,N_11244,N_11453);
or U13157 (N_13157,N_12275,N_12196);
nand U13158 (N_13158,N_12303,N_12257);
and U13159 (N_13159,N_10311,N_12058);
and U13160 (N_13160,N_11207,N_10448);
and U13161 (N_13161,N_11022,N_9601);
and U13162 (N_13162,N_12406,N_11096);
nor U13163 (N_13163,N_12036,N_9525);
nor U13164 (N_13164,N_9593,N_12429);
or U13165 (N_13165,N_10565,N_10121);
xnor U13166 (N_13166,N_11906,N_9953);
xnor U13167 (N_13167,N_10735,N_10595);
nor U13168 (N_13168,N_10450,N_11401);
nor U13169 (N_13169,N_11367,N_11908);
xor U13170 (N_13170,N_10457,N_11365);
nand U13171 (N_13171,N_11316,N_10998);
and U13172 (N_13172,N_11141,N_10634);
or U13173 (N_13173,N_12070,N_11782);
nand U13174 (N_13174,N_11566,N_10477);
and U13175 (N_13175,N_10084,N_10502);
nand U13176 (N_13176,N_11428,N_10891);
nand U13177 (N_13177,N_9389,N_10668);
nor U13178 (N_13178,N_10534,N_10836);
or U13179 (N_13179,N_9376,N_10098);
nor U13180 (N_13180,N_11869,N_9892);
and U13181 (N_13181,N_12115,N_11829);
nand U13182 (N_13182,N_11369,N_10212);
nand U13183 (N_13183,N_12368,N_12376);
nand U13184 (N_13184,N_9897,N_10028);
nand U13185 (N_13185,N_11626,N_10003);
or U13186 (N_13186,N_10176,N_10637);
xnor U13187 (N_13187,N_11539,N_9964);
xor U13188 (N_13188,N_10187,N_10907);
nor U13189 (N_13189,N_10867,N_11114);
xor U13190 (N_13190,N_11896,N_10833);
nand U13191 (N_13191,N_10034,N_11819);
nand U13192 (N_13192,N_10966,N_10839);
nand U13193 (N_13193,N_9657,N_10921);
or U13194 (N_13194,N_12426,N_10129);
xor U13195 (N_13195,N_10798,N_10260);
nand U13196 (N_13196,N_12151,N_12190);
nor U13197 (N_13197,N_10370,N_10432);
nand U13198 (N_13198,N_11348,N_12014);
and U13199 (N_13199,N_10699,N_12422);
nor U13200 (N_13200,N_9573,N_10023);
xnor U13201 (N_13201,N_9654,N_10509);
and U13202 (N_13202,N_9469,N_11288);
or U13203 (N_13203,N_12433,N_9911);
nand U13204 (N_13204,N_10689,N_10889);
nor U13205 (N_13205,N_10541,N_12441);
or U13206 (N_13206,N_11463,N_11230);
xnor U13207 (N_13207,N_11734,N_10357);
xor U13208 (N_13208,N_11989,N_12020);
or U13209 (N_13209,N_11262,N_10561);
nor U13210 (N_13210,N_10209,N_10389);
and U13211 (N_13211,N_12069,N_9992);
xnor U13212 (N_13212,N_12019,N_10391);
and U13213 (N_13213,N_11725,N_11535);
xnor U13214 (N_13214,N_11068,N_12353);
nor U13215 (N_13215,N_12016,N_10544);
and U13216 (N_13216,N_11312,N_11097);
nor U13217 (N_13217,N_10950,N_9538);
nand U13218 (N_13218,N_12264,N_10963);
and U13219 (N_13219,N_10572,N_11176);
nor U13220 (N_13220,N_11359,N_10957);
nand U13221 (N_13221,N_11553,N_9853);
nand U13222 (N_13222,N_11744,N_12044);
nor U13223 (N_13223,N_9895,N_12410);
nor U13224 (N_13224,N_10593,N_12193);
nand U13225 (N_13225,N_11341,N_11127);
xnor U13226 (N_13226,N_11413,N_10520);
nand U13227 (N_13227,N_12211,N_9655);
xor U13228 (N_13228,N_11536,N_9501);
nand U13229 (N_13229,N_10840,N_11098);
xnor U13230 (N_13230,N_12311,N_12273);
nor U13231 (N_13231,N_10102,N_12300);
nor U13232 (N_13232,N_11101,N_10603);
nor U13233 (N_13233,N_9444,N_11082);
or U13234 (N_13234,N_11538,N_11975);
xnor U13235 (N_13235,N_10962,N_11660);
xor U13236 (N_13236,N_11870,N_11786);
and U13237 (N_13237,N_11377,N_10764);
xnor U13238 (N_13238,N_10586,N_9767);
or U13239 (N_13239,N_12104,N_12249);
xor U13240 (N_13240,N_11120,N_11600);
nor U13241 (N_13241,N_12323,N_11749);
xor U13242 (N_13242,N_9995,N_10818);
nor U13243 (N_13243,N_9661,N_11567);
or U13244 (N_13244,N_12139,N_10941);
or U13245 (N_13245,N_11213,N_9716);
or U13246 (N_13246,N_9524,N_9683);
or U13247 (N_13247,N_9810,N_10490);
nor U13248 (N_13248,N_11123,N_12023);
and U13249 (N_13249,N_9708,N_10140);
xnor U13250 (N_13250,N_11011,N_11201);
nand U13251 (N_13251,N_9576,N_10088);
xnor U13252 (N_13252,N_12147,N_10168);
or U13253 (N_13253,N_11164,N_11059);
xnor U13254 (N_13254,N_11838,N_9979);
nand U13255 (N_13255,N_10228,N_9809);
or U13256 (N_13256,N_11483,N_12302);
or U13257 (N_13257,N_10446,N_11559);
and U13258 (N_13258,N_10597,N_10674);
or U13259 (N_13259,N_9498,N_12215);
nand U13260 (N_13260,N_10285,N_9695);
or U13261 (N_13261,N_10115,N_11930);
xnor U13262 (N_13262,N_9900,N_12270);
and U13263 (N_13263,N_12265,N_10756);
and U13264 (N_13264,N_10522,N_10776);
or U13265 (N_13265,N_11331,N_9494);
xnor U13266 (N_13266,N_9973,N_11826);
nand U13267 (N_13267,N_11745,N_12350);
and U13268 (N_13268,N_11736,N_12123);
nand U13269 (N_13269,N_9431,N_9592);
xnor U13270 (N_13270,N_10275,N_11609);
xnor U13271 (N_13271,N_10765,N_11653);
and U13272 (N_13272,N_11152,N_12052);
or U13273 (N_13273,N_12271,N_11846);
nor U13274 (N_13274,N_10247,N_11434);
xor U13275 (N_13275,N_11673,N_11034);
nor U13276 (N_13276,N_11639,N_11415);
and U13277 (N_13277,N_11074,N_11196);
xnor U13278 (N_13278,N_9492,N_9857);
and U13279 (N_13279,N_11748,N_10731);
nand U13280 (N_13280,N_10517,N_12008);
and U13281 (N_13281,N_11708,N_9569);
and U13282 (N_13282,N_10706,N_12408);
and U13283 (N_13283,N_9382,N_10386);
and U13284 (N_13284,N_12076,N_11887);
or U13285 (N_13285,N_11148,N_12312);
nor U13286 (N_13286,N_12106,N_9870);
nand U13287 (N_13287,N_10917,N_10834);
nor U13288 (N_13288,N_11309,N_11445);
nor U13289 (N_13289,N_10732,N_12040);
nor U13290 (N_13290,N_12232,N_10652);
nand U13291 (N_13291,N_11665,N_11574);
nand U13292 (N_13292,N_11216,N_9651);
and U13293 (N_13293,N_11948,N_10643);
xor U13294 (N_13294,N_9827,N_11217);
nor U13295 (N_13295,N_12401,N_9802);
nand U13296 (N_13296,N_10429,N_11959);
xor U13297 (N_13297,N_12280,N_10571);
and U13298 (N_13298,N_11311,N_9741);
xnor U13299 (N_13299,N_9582,N_10289);
nand U13300 (N_13300,N_12029,N_10021);
xnor U13301 (N_13301,N_12269,N_9667);
nand U13302 (N_13302,N_10392,N_10283);
nor U13303 (N_13303,N_10111,N_12013);
nor U13304 (N_13304,N_11260,N_11375);
nand U13305 (N_13305,N_11095,N_11772);
and U13306 (N_13306,N_12229,N_9421);
and U13307 (N_13307,N_10030,N_9999);
xor U13308 (N_13308,N_10705,N_11170);
or U13309 (N_13309,N_12212,N_9776);
xnor U13310 (N_13310,N_9846,N_9518);
nor U13311 (N_13311,N_10583,N_11664);
nor U13312 (N_13312,N_10053,N_10313);
and U13313 (N_13313,N_9881,N_11431);
xor U13314 (N_13314,N_10578,N_10584);
nor U13315 (N_13315,N_11484,N_9968);
xor U13316 (N_13316,N_12072,N_11684);
nor U13317 (N_13317,N_9520,N_11228);
nand U13318 (N_13318,N_11879,N_9410);
nor U13319 (N_13319,N_10633,N_9877);
or U13320 (N_13320,N_10282,N_12329);
xnor U13321 (N_13321,N_10912,N_11602);
xnor U13322 (N_13322,N_11455,N_9595);
xor U13323 (N_13323,N_10679,N_11654);
nand U13324 (N_13324,N_11266,N_10508);
and U13325 (N_13325,N_10100,N_10093);
and U13326 (N_13326,N_10298,N_11145);
or U13327 (N_13327,N_12340,N_10007);
and U13328 (N_13328,N_10700,N_11110);
and U13329 (N_13329,N_11387,N_12082);
or U13330 (N_13330,N_9440,N_11218);
or U13331 (N_13331,N_11728,N_11339);
nand U13332 (N_13332,N_10551,N_11917);
nand U13333 (N_13333,N_9790,N_11682);
nor U13334 (N_13334,N_11173,N_11514);
nor U13335 (N_13335,N_12439,N_12277);
and U13336 (N_13336,N_12389,N_10242);
nor U13337 (N_13337,N_12064,N_10310);
and U13338 (N_13338,N_9910,N_11396);
nand U13339 (N_13339,N_11303,N_10238);
nor U13340 (N_13340,N_11017,N_9700);
nand U13341 (N_13341,N_10835,N_10528);
nor U13342 (N_13342,N_11677,N_11927);
and U13343 (N_13343,N_9615,N_10720);
nand U13344 (N_13344,N_9955,N_11416);
nand U13345 (N_13345,N_10184,N_10738);
xor U13346 (N_13346,N_11515,N_10795);
nand U13347 (N_13347,N_10164,N_10273);
nand U13348 (N_13348,N_10428,N_9532);
nand U13349 (N_13349,N_11406,N_9648);
and U13350 (N_13350,N_11467,N_10886);
and U13351 (N_13351,N_12289,N_9393);
nand U13352 (N_13352,N_9926,N_10893);
xor U13353 (N_13353,N_10514,N_12364);
nor U13354 (N_13354,N_10341,N_10217);
or U13355 (N_13355,N_10141,N_10171);
and U13356 (N_13356,N_9721,N_11510);
or U13357 (N_13357,N_10677,N_11519);
nor U13358 (N_13358,N_10347,N_11506);
or U13359 (N_13359,N_10703,N_12039);
and U13360 (N_13360,N_11067,N_10354);
xnor U13361 (N_13361,N_10612,N_10077);
and U13362 (N_13362,N_12288,N_12372);
xnor U13363 (N_13363,N_12091,N_9585);
nor U13364 (N_13364,N_10224,N_11472);
or U13365 (N_13365,N_11797,N_9938);
or U13366 (N_13366,N_9422,N_9923);
nand U13367 (N_13367,N_11474,N_10591);
or U13368 (N_13368,N_9508,N_10397);
and U13369 (N_13369,N_11394,N_10233);
or U13370 (N_13370,N_9662,N_9604);
nor U13371 (N_13371,N_10539,N_12186);
and U13372 (N_13372,N_11162,N_11764);
or U13373 (N_13373,N_9643,N_11939);
or U13374 (N_13374,N_11015,N_11874);
or U13375 (N_13375,N_10130,N_10294);
nor U13376 (N_13376,N_12053,N_12140);
nand U13377 (N_13377,N_10255,N_11443);
nor U13378 (N_13378,N_11180,N_11832);
nand U13379 (N_13379,N_10447,N_10883);
xor U13380 (N_13380,N_9497,N_10575);
or U13381 (N_13381,N_10841,N_11584);
or U13382 (N_13382,N_11157,N_9544);
or U13383 (N_13383,N_9473,N_10395);
xor U13384 (N_13384,N_10614,N_11987);
xnor U13385 (N_13385,N_11875,N_11276);
and U13386 (N_13386,N_12048,N_10991);
nand U13387 (N_13387,N_12320,N_11310);
xnor U13388 (N_13388,N_9554,N_10605);
or U13389 (N_13389,N_11980,N_12451);
xor U13390 (N_13390,N_10332,N_11743);
xnor U13391 (N_13391,N_9943,N_9411);
and U13392 (N_13392,N_11634,N_11299);
nand U13393 (N_13393,N_9812,N_9836);
nor U13394 (N_13394,N_10300,N_11707);
nor U13395 (N_13395,N_9686,N_11111);
xnor U13396 (N_13396,N_11253,N_9401);
or U13397 (N_13397,N_10137,N_10122);
or U13398 (N_13398,N_10103,N_9578);
nor U13399 (N_13399,N_10760,N_10868);
or U13400 (N_13400,N_11432,N_9729);
xnor U13401 (N_13401,N_10888,N_12094);
xor U13402 (N_13402,N_9815,N_10492);
nand U13403 (N_13403,N_11144,N_9484);
and U13404 (N_13404,N_11680,N_10856);
nor U13405 (N_13405,N_10367,N_11988);
nor U13406 (N_13406,N_10475,N_10958);
or U13407 (N_13407,N_10942,N_10443);
xnor U13408 (N_13408,N_9542,N_9663);
and U13409 (N_13409,N_11905,N_12157);
or U13410 (N_13410,N_11573,N_9556);
xnor U13411 (N_13411,N_11582,N_9379);
xnor U13412 (N_13412,N_9826,N_11770);
xnor U13413 (N_13413,N_11412,N_11398);
nand U13414 (N_13414,N_10669,N_12283);
nand U13415 (N_13415,N_12394,N_11325);
nor U13416 (N_13416,N_12392,N_12051);
nor U13417 (N_13417,N_11187,N_11972);
or U13418 (N_13418,N_10440,N_11594);
and U13419 (N_13419,N_12121,N_10866);
nor U13420 (N_13420,N_11894,N_12471);
nor U13421 (N_13421,N_12218,N_10728);
and U13422 (N_13422,N_11302,N_12063);
and U13423 (N_13423,N_10363,N_10617);
and U13424 (N_13424,N_11106,N_12351);
xor U13425 (N_13425,N_11281,N_12349);
or U13426 (N_13426,N_11040,N_9760);
nor U13427 (N_13427,N_9656,N_10640);
nand U13428 (N_13428,N_11193,N_10562);
nand U13429 (N_13429,N_11889,N_9418);
and U13430 (N_13430,N_9771,N_10890);
nor U13431 (N_13431,N_9452,N_11713);
nand U13432 (N_13432,N_11393,N_12377);
or U13433 (N_13433,N_12452,N_10611);
xnor U13434 (N_13434,N_10628,N_10932);
nor U13435 (N_13435,N_12326,N_10229);
xnor U13436 (N_13436,N_10194,N_10645);
and U13437 (N_13437,N_10236,N_10895);
nor U13438 (N_13438,N_10815,N_11727);
and U13439 (N_13439,N_11036,N_11324);
nor U13440 (N_13440,N_11911,N_10762);
nor U13441 (N_13441,N_12445,N_9712);
nand U13442 (N_13442,N_10948,N_11112);
xor U13443 (N_13443,N_10532,N_9565);
nand U13444 (N_13444,N_11277,N_10065);
nor U13445 (N_13445,N_9613,N_12404);
or U13446 (N_13446,N_10417,N_11010);
xor U13447 (N_13447,N_9933,N_10059);
nor U13448 (N_13448,N_11147,N_11211);
or U13449 (N_13449,N_9994,N_10843);
nand U13450 (N_13450,N_10470,N_9660);
or U13451 (N_13451,N_11606,N_10263);
xnor U13452 (N_13452,N_10781,N_10024);
or U13453 (N_13453,N_11834,N_12206);
or U13454 (N_13454,N_9825,N_11758);
xnor U13455 (N_13455,N_10849,N_11644);
xnor U13456 (N_13456,N_11105,N_10726);
nor U13457 (N_13457,N_10046,N_9779);
nand U13458 (N_13458,N_10055,N_12369);
or U13459 (N_13459,N_11374,N_9574);
nor U13460 (N_13460,N_11372,N_9402);
or U13461 (N_13461,N_9814,N_11955);
nand U13462 (N_13462,N_10959,N_11636);
xnor U13463 (N_13463,N_10505,N_11918);
and U13464 (N_13464,N_12409,N_10601);
or U13465 (N_13465,N_11722,N_9681);
xnor U13466 (N_13466,N_9674,N_10510);
xor U13467 (N_13467,N_12205,N_9590);
or U13468 (N_13468,N_11571,N_11400);
or U13469 (N_13469,N_9617,N_11833);
nand U13470 (N_13470,N_12095,N_10319);
and U13471 (N_13471,N_12001,N_11512);
nand U13472 (N_13472,N_10149,N_10500);
and U13473 (N_13473,N_10082,N_11140);
and U13474 (N_13474,N_10955,N_11269);
and U13475 (N_13475,N_11168,N_11994);
nor U13476 (N_13476,N_11998,N_12117);
nor U13477 (N_13477,N_10350,N_11107);
nand U13478 (N_13478,N_10195,N_10906);
nand U13479 (N_13479,N_11286,N_11263);
nor U13480 (N_13480,N_10916,N_11950);
nand U13481 (N_13481,N_9940,N_11837);
nor U13482 (N_13482,N_10453,N_11248);
xnor U13483 (N_13483,N_11130,N_11580);
and U13484 (N_13484,N_9398,N_9539);
or U13485 (N_13485,N_11921,N_12204);
nor U13486 (N_13486,N_9519,N_9570);
nor U13487 (N_13487,N_9867,N_10048);
xor U13488 (N_13488,N_11563,N_9840);
xnor U13489 (N_13489,N_11820,N_9594);
nand U13490 (N_13490,N_10826,N_9394);
and U13491 (N_13491,N_9725,N_11025);
nand U13492 (N_13492,N_9458,N_10691);
and U13493 (N_13493,N_10801,N_11855);
xor U13494 (N_13494,N_10162,N_10185);
or U13495 (N_13495,N_10545,N_11420);
xor U13496 (N_13496,N_10044,N_11720);
and U13497 (N_13497,N_11900,N_9837);
xnor U13498 (N_13498,N_9460,N_12024);
or U13499 (N_13499,N_11638,N_10246);
nor U13500 (N_13500,N_10862,N_10922);
or U13501 (N_13501,N_10622,N_10779);
and U13502 (N_13502,N_12081,N_11757);
xnor U13503 (N_13503,N_10293,N_9971);
and U13504 (N_13504,N_12098,N_11753);
and U13505 (N_13505,N_11760,N_10861);
nor U13506 (N_13506,N_9403,N_11575);
nand U13507 (N_13507,N_9462,N_10813);
or U13508 (N_13508,N_12460,N_11861);
or U13509 (N_13509,N_11597,N_10039);
nand U13510 (N_13510,N_9848,N_10707);
or U13511 (N_13511,N_11803,N_9855);
nand U13512 (N_13512,N_12282,N_11189);
nand U13513 (N_13513,N_10151,N_10394);
nand U13514 (N_13514,N_10809,N_12437);
and U13515 (N_13515,N_11923,N_9464);
xnor U13516 (N_13516,N_10892,N_11685);
or U13517 (N_13517,N_12440,N_11655);
nor U13518 (N_13518,N_10778,N_10276);
and U13519 (N_13519,N_11529,N_11418);
or U13520 (N_13520,N_11742,N_12490);
and U13521 (N_13521,N_11440,N_11052);
nor U13522 (N_13522,N_9488,N_11421);
xnor U13523 (N_13523,N_10226,N_12105);
xnor U13524 (N_13524,N_11271,N_9993);
and U13525 (N_13525,N_10114,N_12021);
and U13526 (N_13526,N_9946,N_12074);
or U13527 (N_13527,N_12430,N_10324);
or U13528 (N_13528,N_11256,N_9427);
nor U13529 (N_13529,N_10288,N_11086);
nor U13530 (N_13530,N_9455,N_11721);
nand U13531 (N_13531,N_9665,N_11167);
or U13532 (N_13532,N_10729,N_10345);
nor U13533 (N_13533,N_11912,N_10554);
and U13534 (N_13534,N_9948,N_12446);
xnor U13535 (N_13535,N_12118,N_10506);
nand U13536 (N_13536,N_10452,N_9838);
nor U13537 (N_13537,N_9739,N_9449);
or U13538 (N_13538,N_11280,N_11078);
nand U13539 (N_13539,N_9433,N_12497);
nor U13540 (N_13540,N_9945,N_9634);
xor U13541 (N_13541,N_11576,N_10543);
and U13542 (N_13542,N_11154,N_10747);
nor U13543 (N_13543,N_10124,N_9391);
nor U13544 (N_13544,N_10570,N_9438);
xnor U13545 (N_13545,N_11851,N_11643);
and U13546 (N_13546,N_10519,N_10110);
and U13547 (N_13547,N_12468,N_11221);
nor U13548 (N_13548,N_11815,N_12333);
or U13549 (N_13549,N_10616,N_10267);
nand U13550 (N_13550,N_10099,N_9491);
nand U13551 (N_13551,N_11126,N_9475);
and U13552 (N_13552,N_11361,N_12221);
xnor U13553 (N_13553,N_11308,N_10170);
and U13554 (N_13554,N_10471,N_12207);
nor U13555 (N_13555,N_9884,N_10067);
or U13556 (N_13556,N_10261,N_11060);
nand U13557 (N_13557,N_10305,N_11238);
nor U13558 (N_13558,N_12444,N_11323);
xor U13559 (N_13559,N_11043,N_11268);
nor U13560 (N_13560,N_11766,N_11856);
nor U13561 (N_13561,N_11314,N_11511);
nand U13562 (N_13562,N_10754,N_12096);
nor U13563 (N_13563,N_11103,N_10264);
xnor U13564 (N_13564,N_12442,N_12458);
nand U13565 (N_13565,N_11953,N_10037);
or U13566 (N_13566,N_9866,N_9419);
or U13567 (N_13567,N_11151,N_10063);
and U13568 (N_13568,N_11965,N_11371);
and U13569 (N_13569,N_10542,N_11890);
and U13570 (N_13570,N_11001,N_11200);
xor U13571 (N_13571,N_11452,N_9733);
nand U13572 (N_13572,N_10563,N_11666);
or U13573 (N_13573,N_9772,N_11224);
and U13574 (N_13574,N_10763,N_10355);
and U13575 (N_13575,N_11202,N_9706);
and U13576 (N_13576,N_10106,N_10371);
xor U13577 (N_13577,N_9967,N_9735);
and U13578 (N_13578,N_11081,N_12482);
xnor U13579 (N_13579,N_9678,N_10163);
or U13580 (N_13580,N_9888,N_12489);
nor U13581 (N_13581,N_10322,N_11579);
or U13582 (N_13582,N_9412,N_10484);
and U13583 (N_13583,N_9724,N_11073);
nand U13584 (N_13584,N_10105,N_10944);
or U13585 (N_13585,N_10230,N_10139);
or U13586 (N_13586,N_10349,N_9579);
or U13587 (N_13587,N_10165,N_9841);
or U13588 (N_13588,N_9448,N_11712);
and U13589 (N_13589,N_10761,N_10512);
xnor U13590 (N_13590,N_12101,N_10515);
nand U13591 (N_13591,N_9385,N_11338);
and U13592 (N_13592,N_11210,N_10822);
nor U13593 (N_13593,N_10686,N_11943);
nor U13594 (N_13594,N_9987,N_10620);
or U13595 (N_13595,N_9522,N_11273);
and U13596 (N_13596,N_10642,N_10956);
and U13597 (N_13597,N_11353,N_11898);
xnor U13598 (N_13598,N_9676,N_12041);
or U13599 (N_13599,N_9406,N_11810);
nand U13600 (N_13600,N_10250,N_10986);
nand U13601 (N_13601,N_12045,N_10533);
nand U13602 (N_13602,N_10218,N_10362);
nand U13603 (N_13603,N_12294,N_9572);
nor U13604 (N_13604,N_11468,N_11649);
and U13605 (N_13605,N_11199,N_9627);
or U13606 (N_13606,N_10427,N_10549);
nand U13607 (N_13607,N_10741,N_9536);
xnor U13608 (N_13608,N_9913,N_10908);
or U13609 (N_13609,N_9434,N_9736);
nand U13610 (N_13610,N_11492,N_12470);
nand U13611 (N_13611,N_10690,N_10306);
or U13612 (N_13612,N_12268,N_11064);
xor U13613 (N_13613,N_10001,N_10925);
or U13614 (N_13614,N_12109,N_9894);
and U13615 (N_13615,N_12017,N_12483);
nor U13616 (N_13616,N_11656,N_10478);
xor U13617 (N_13617,N_11822,N_9912);
nor U13618 (N_13618,N_11814,N_10227);
nor U13619 (N_13619,N_12496,N_11793);
nor U13620 (N_13620,N_9476,N_11586);
nand U13621 (N_13621,N_9778,N_12197);
xnor U13622 (N_13622,N_12079,N_11503);
nand U13623 (N_13623,N_11388,N_10850);
nand U13624 (N_13624,N_10406,N_9687);
xnor U13625 (N_13625,N_12254,N_9587);
or U13626 (N_13626,N_9399,N_10816);
nand U13627 (N_13627,N_11188,N_9949);
xor U13628 (N_13628,N_10649,N_11548);
and U13629 (N_13629,N_9756,N_10627);
xnor U13630 (N_13630,N_9969,N_10923);
nor U13631 (N_13631,N_11747,N_10375);
or U13632 (N_13632,N_12313,N_11628);
nand U13633 (N_13633,N_9770,N_10983);
nand U13634 (N_13634,N_9996,N_11944);
xor U13635 (N_13635,N_9930,N_11212);
or U13636 (N_13636,N_10518,N_10967);
xnor U13637 (N_13637,N_11791,N_11886);
or U13638 (N_13638,N_10107,N_10954);
and U13639 (N_13639,N_10487,N_9567);
xor U13640 (N_13640,N_9477,N_9966);
or U13641 (N_13641,N_11146,N_12239);
xor U13642 (N_13642,N_10713,N_12428);
xnor U13643 (N_13643,N_11143,N_10629);
nand U13644 (N_13644,N_10337,N_11885);
nand U13645 (N_13645,N_11767,N_10366);
and U13646 (N_13646,N_10192,N_12243);
nand U13647 (N_13647,N_9786,N_11615);
nor U13648 (N_13648,N_9922,N_10161);
and U13649 (N_13649,N_12398,N_11773);
or U13650 (N_13650,N_10032,N_11877);
nand U13651 (N_13651,N_10585,N_12132);
nor U13652 (N_13652,N_12475,N_11267);
xnor U13653 (N_13653,N_11999,N_10009);
xnor U13654 (N_13654,N_11174,N_11019);
and U13655 (N_13655,N_12222,N_11498);
nor U13656 (N_13656,N_12464,N_10422);
nand U13657 (N_13657,N_9869,N_9642);
nor U13658 (N_13658,N_10455,N_12453);
xor U13659 (N_13659,N_10321,N_11928);
xnor U13660 (N_13660,N_9751,N_10536);
and U13661 (N_13661,N_10201,N_10773);
nor U13662 (N_13662,N_12225,N_9679);
nor U13663 (N_13663,N_10656,N_12188);
nand U13664 (N_13664,N_11702,N_10451);
xnor U13665 (N_13665,N_12050,N_12250);
or U13666 (N_13666,N_9854,N_9446);
nand U13667 (N_13667,N_10497,N_11568);
and U13668 (N_13668,N_9632,N_10716);
and U13669 (N_13669,N_10463,N_11480);
nor U13670 (N_13670,N_10365,N_10581);
nor U13671 (N_13671,N_10279,N_12325);
xor U13672 (N_13672,N_11362,N_11405);
nand U13673 (N_13673,N_9750,N_10489);
and U13674 (N_13674,N_10020,N_12420);
nor U13675 (N_13675,N_12293,N_11169);
nand U13676 (N_13676,N_9568,N_9549);
or U13677 (N_13677,N_9765,N_12499);
xor U13678 (N_13678,N_9546,N_11100);
nand U13679 (N_13679,N_10807,N_10530);
and U13680 (N_13680,N_12165,N_11491);
or U13681 (N_13681,N_12210,N_11632);
and U13682 (N_13682,N_11153,N_10975);
nand U13683 (N_13683,N_11645,N_11030);
nand U13684 (N_13684,N_9603,N_9823);
nand U13685 (N_13685,N_9616,N_12131);
or U13686 (N_13686,N_11185,N_10814);
and U13687 (N_13687,N_12026,N_11023);
or U13688 (N_13688,N_10473,N_9956);
nand U13689 (N_13689,N_9621,N_9566);
and U13690 (N_13690,N_9558,N_10940);
or U13691 (N_13691,N_11646,N_10459);
nor U13692 (N_13692,N_9944,N_10521);
xor U13693 (N_13693,N_12248,N_11974);
or U13694 (N_13694,N_10985,N_11466);
or U13695 (N_13695,N_10808,N_10503);
or U13696 (N_13696,N_11768,N_10680);
or U13697 (N_13697,N_10249,N_10496);
nand U13698 (N_13698,N_11289,N_12371);
nand U13699 (N_13699,N_10709,N_10012);
and U13700 (N_13700,N_11642,N_11621);
and U13701 (N_13701,N_9775,N_11251);
and U13702 (N_13702,N_9806,N_11305);
and U13703 (N_13703,N_10621,N_12328);
nand U13704 (N_13704,N_9653,N_12116);
and U13705 (N_13705,N_10278,N_12387);
xor U13706 (N_13706,N_11275,N_11587);
nor U13707 (N_13707,N_11350,N_11771);
or U13708 (N_13708,N_10368,N_10211);
or U13709 (N_13709,N_10931,N_12201);
and U13710 (N_13710,N_10576,N_9950);
nor U13711 (N_13711,N_11852,N_10523);
nand U13712 (N_13712,N_12060,N_11093);
and U13713 (N_13713,N_11186,N_10846);
nor U13714 (N_13714,N_10860,N_10825);
nand U13715 (N_13715,N_12405,N_11071);
or U13716 (N_13716,N_11414,N_10884);
nand U13717 (N_13717,N_9715,N_9797);
and U13718 (N_13718,N_9803,N_10935);
nor U13719 (N_13719,N_10108,N_11435);
or U13720 (N_13720,N_11630,N_12487);
xor U13721 (N_13721,N_10488,N_10961);
xor U13722 (N_13722,N_12018,N_10874);
xor U13723 (N_13723,N_10546,N_10644);
nand U13724 (N_13724,N_12454,N_10538);
and U13725 (N_13725,N_10464,N_11641);
nor U13726 (N_13726,N_9583,N_12467);
xor U13727 (N_13727,N_10796,N_11581);
nand U13728 (N_13728,N_11496,N_10049);
xnor U13729 (N_13729,N_9500,N_10919);
nor U13730 (N_13730,N_9420,N_11662);
nand U13731 (N_13731,N_9688,N_12230);
nand U13732 (N_13732,N_11966,N_10280);
nor U13733 (N_13733,N_11247,N_12219);
nor U13734 (N_13734,N_9865,N_11344);
xor U13735 (N_13735,N_12380,N_11233);
or U13736 (N_13736,N_12128,N_9668);
xor U13737 (N_13737,N_11459,N_9998);
or U13738 (N_13738,N_10589,N_12315);
nand U13739 (N_13739,N_12170,N_10064);
nor U13740 (N_13740,N_9465,N_11198);
nor U13741 (N_13741,N_10150,N_11460);
nor U13742 (N_13742,N_9470,N_11790);
and U13743 (N_13743,N_10092,N_12305);
or U13744 (N_13744,N_10356,N_11729);
and U13745 (N_13745,N_12223,N_10175);
or U13746 (N_13746,N_11845,N_10972);
xor U13747 (N_13747,N_11092,N_12162);
and U13748 (N_13748,N_11392,N_11620);
or U13749 (N_13749,N_11859,N_11843);
nand U13750 (N_13750,N_11373,N_10206);
or U13751 (N_13751,N_12331,N_10873);
and U13752 (N_13752,N_11976,N_10782);
or U13753 (N_13753,N_12059,N_11249);
nand U13754 (N_13754,N_10784,N_11993);
xnor U13755 (N_13755,N_11907,N_12462);
nor U13756 (N_13756,N_10177,N_11779);
xnor U13757 (N_13757,N_10312,N_10317);
and U13758 (N_13758,N_10752,N_12412);
nor U13759 (N_13759,N_11270,N_10189);
or U13760 (N_13760,N_10693,N_11159);
xnor U13761 (N_13761,N_11038,N_10702);
nor U13762 (N_13762,N_11667,N_10678);
nor U13763 (N_13763,N_10066,N_10525);
and U13764 (N_13764,N_10080,N_11252);
or U13765 (N_13765,N_10794,N_11089);
xor U13766 (N_13766,N_9934,N_10072);
or U13767 (N_13767,N_12042,N_10329);
nand U13768 (N_13768,N_9392,N_9931);
or U13769 (N_13769,N_10568,N_11242);
or U13770 (N_13770,N_12208,N_10254);
nand U13771 (N_13771,N_11264,N_10569);
and U13772 (N_13772,N_9571,N_9808);
nor U13773 (N_13773,N_9557,N_11284);
nand U13774 (N_13774,N_11672,N_12317);
xnor U13775 (N_13775,N_10531,N_10123);
and U13776 (N_13776,N_12450,N_12419);
nand U13777 (N_13777,N_11298,N_10384);
nor U13778 (N_13778,N_10969,N_11922);
and U13779 (N_13779,N_12080,N_11892);
nand U13780 (N_13780,N_9844,N_10933);
nand U13781 (N_13781,N_10664,N_10858);
and U13782 (N_13782,N_11355,N_11137);
and U13783 (N_13783,N_10876,N_11451);
nand U13784 (N_13784,N_12216,N_11192);
or U13785 (N_13785,N_11973,N_12002);
nand U13786 (N_13786,N_11679,N_11165);
or U13787 (N_13787,N_10359,N_9563);
or U13788 (N_13788,N_12348,N_10133);
nor U13789 (N_13789,N_10800,N_10574);
or U13790 (N_13790,N_11327,N_10820);
nor U13791 (N_13791,N_10172,N_12381);
or U13792 (N_13792,N_12357,N_11191);
xnor U13793 (N_13793,N_10661,N_12156);
or U13794 (N_13794,N_11570,N_12067);
xor U13795 (N_13795,N_10407,N_10193);
nand U13796 (N_13796,N_11629,N_12296);
nand U13797 (N_13797,N_9482,N_9450);
xor U13798 (N_13798,N_9937,N_12252);
and U13799 (N_13799,N_9584,N_11862);
nand U13800 (N_13800,N_10036,N_10117);
and U13801 (N_13801,N_11604,N_12486);
nand U13802 (N_13802,N_9435,N_12087);
xor U13803 (N_13803,N_10555,N_9863);
or U13804 (N_13804,N_9596,N_11438);
or U13805 (N_13805,N_9816,N_11778);
or U13806 (N_13806,N_11572,N_10125);
nor U13807 (N_13807,N_10190,N_10442);
nand U13808 (N_13808,N_11588,N_12403);
xnor U13809 (N_13809,N_12032,N_10553);
and U13810 (N_13810,N_11614,N_10031);
and U13811 (N_13811,N_10725,N_11424);
and U13812 (N_13812,N_12285,N_12180);
nand U13813 (N_13813,N_9535,N_11546);
xor U13814 (N_13814,N_9917,N_11701);
or U13815 (N_13815,N_11726,N_11893);
or U13816 (N_13816,N_10920,N_11447);
nor U13817 (N_13817,N_11045,N_11129);
xor U13818 (N_13818,N_10057,N_11258);
xor U13819 (N_13819,N_11610,N_11125);
and U13820 (N_13820,N_12367,N_10854);
xnor U13821 (N_13821,N_11785,N_12255);
nand U13822 (N_13822,N_10504,N_12236);
nand U13823 (N_13823,N_12477,N_11363);
and U13824 (N_13824,N_9880,N_11873);
and U13825 (N_13825,N_11794,N_11997);
or U13826 (N_13826,N_9918,N_10552);
nor U13827 (N_13827,N_11780,N_11053);
nand U13828 (N_13828,N_11599,N_10308);
xnor U13829 (N_13829,N_10865,N_11250);
and U13830 (N_13830,N_11883,N_10704);
and U13831 (N_13831,N_9636,N_10461);
nand U13832 (N_13832,N_9694,N_11926);
and U13833 (N_13833,N_12043,N_11225);
xnor U13834 (N_13834,N_9924,N_10635);
nand U13835 (N_13835,N_11872,N_10369);
and U13836 (N_13836,N_9423,N_9459);
or U13837 (N_13837,N_9521,N_11083);
or U13838 (N_13838,N_11026,N_11477);
xor U13839 (N_13839,N_9637,N_11077);
and U13840 (N_13840,N_10560,N_11932);
or U13841 (N_13841,N_9417,N_10881);
or U13842 (N_13842,N_12366,N_11788);
nor U13843 (N_13843,N_10335,N_11240);
and U13844 (N_13844,N_10134,N_12145);
nor U13845 (N_13845,N_11304,N_11694);
or U13846 (N_13846,N_9639,N_12342);
and U13847 (N_13847,N_11613,N_12159);
and U13848 (N_13848,N_9963,N_9670);
nor U13849 (N_13849,N_9646,N_11518);
xor U13850 (N_13850,N_9408,N_9506);
and U13851 (N_13851,N_10516,N_11691);
nand U13852 (N_13852,N_9659,N_12434);
xnor U13853 (N_13853,N_11871,N_10766);
nand U13854 (N_13854,N_12290,N_12133);
xor U13855 (N_13855,N_10075,N_12318);
nor U13856 (N_13856,N_9761,N_11411);
nand U13857 (N_13857,N_9479,N_12174);
and U13858 (N_13858,N_12449,N_10683);
nor U13859 (N_13859,N_10038,N_9727);
nor U13860 (N_13860,N_10334,N_10182);
and U13861 (N_13861,N_11805,N_9997);
xnor U13862 (N_13862,N_9545,N_12472);
nor U13863 (N_13863,N_10641,N_9766);
or U13864 (N_13864,N_12343,N_10096);
nand U13865 (N_13865,N_10929,N_9904);
nand U13866 (N_13866,N_10624,N_11446);
or U13867 (N_13867,N_12065,N_11358);
and U13868 (N_13868,N_10791,N_10197);
nor U13869 (N_13869,N_10810,N_10138);
nand U13870 (N_13870,N_11378,N_10960);
and U13871 (N_13871,N_12086,N_10328);
and U13872 (N_13872,N_10438,N_10245);
xor U13873 (N_13873,N_9548,N_12136);
xnor U13874 (N_13874,N_10877,N_11775);
and U13875 (N_13875,N_9789,N_10524);
or U13876 (N_13876,N_9720,N_12099);
xnor U13877 (N_13877,N_9833,N_10722);
or U13878 (N_13878,N_11848,N_12291);
and U13879 (N_13879,N_11291,N_11205);
xor U13880 (N_13880,N_11190,N_10205);
xnor U13881 (N_13881,N_11937,N_12427);
xnor U13882 (N_13882,N_12097,N_12402);
or U13883 (N_13883,N_11065,N_9424);
and U13884 (N_13884,N_10346,N_11984);
xor U13885 (N_13885,N_9792,N_11149);
nor U13886 (N_13886,N_10911,N_11417);
nor U13887 (N_13887,N_10231,N_10682);
or U13888 (N_13888,N_10737,N_11978);
nand U13889 (N_13889,N_12137,N_11037);
or U13890 (N_13890,N_11470,N_11386);
xor U13891 (N_13891,N_9485,N_12386);
or U13892 (N_13892,N_11847,N_12093);
or U13893 (N_13893,N_10719,N_9493);
nor U13894 (N_13894,N_9502,N_9832);
nand U13895 (N_13895,N_9437,N_9454);
or U13896 (N_13896,N_10444,N_11203);
and U13897 (N_13897,N_11177,N_10296);
nor U13898 (N_13898,N_10174,N_9718);
xor U13899 (N_13899,N_10173,N_11631);
and U13900 (N_13900,N_11457,N_9378);
xnor U13901 (N_13901,N_11595,N_10070);
or U13902 (N_13902,N_12011,N_11556);
nand U13903 (N_13903,N_12144,N_9813);
xnor U13904 (N_13904,N_11234,N_11699);
and U13905 (N_13905,N_10946,N_9640);
or U13906 (N_13906,N_10091,N_11946);
and U13907 (N_13907,N_10050,N_11949);
or U13908 (N_13908,N_10074,N_10027);
nand U13909 (N_13909,N_11085,N_11493);
nand U13910 (N_13910,N_11692,N_11012);
nand U13911 (N_13911,N_11384,N_11982);
or U13912 (N_13912,N_9754,N_9748);
nor U13913 (N_13913,N_11733,N_9936);
nand U13914 (N_13914,N_10015,N_12231);
xor U13915 (N_13915,N_10899,N_10938);
nand U13916 (N_13916,N_10830,N_11255);
and U13917 (N_13917,N_12481,N_12455);
nand U13918 (N_13918,N_9898,N_10673);
xor U13919 (N_13919,N_9598,N_11475);
nor U13920 (N_13920,N_9591,N_12492);
nand U13921 (N_13921,N_11301,N_9515);
nor U13922 (N_13922,N_10147,N_11356);
or U13923 (N_13923,N_9871,N_12226);
or U13924 (N_13924,N_11057,N_10947);
or U13925 (N_13925,N_10875,N_9774);
xor U13926 (N_13926,N_11313,N_10008);
xnor U13927 (N_13927,N_12493,N_10824);
or U13928 (N_13928,N_12332,N_10087);
nand U13929 (N_13929,N_11533,N_11383);
or U13930 (N_13930,N_11592,N_11880);
xor U13931 (N_13931,N_11347,N_9381);
nand U13932 (N_13932,N_11051,N_10157);
xor U13933 (N_13933,N_11698,N_10943);
and U13934 (N_13934,N_9626,N_12185);
or U13935 (N_13935,N_10787,N_9559);
or U13936 (N_13936,N_10647,N_12130);
and U13937 (N_13937,N_10325,N_11823);
or U13938 (N_13938,N_9499,N_11693);
or U13939 (N_13939,N_10142,N_11419);
xnor U13940 (N_13940,N_12037,N_10851);
nand U13941 (N_13941,N_10655,N_9719);
nor U13942 (N_13942,N_11433,N_12324);
or U13943 (N_13943,N_9575,N_11382);
xor U13944 (N_13944,N_12301,N_12034);
xor U13945 (N_13945,N_12345,N_12432);
nor U13946 (N_13946,N_10454,N_12084);
xor U13947 (N_13947,N_12259,N_10566);
nand U13948 (N_13948,N_10974,N_11796);
nor U13949 (N_13949,N_9830,N_10017);
and U13950 (N_13950,N_10483,N_10336);
nor U13951 (N_13951,N_9707,N_11231);
xnor U13952 (N_13952,N_12234,N_10872);
or U13953 (N_13953,N_12397,N_10244);
and U13954 (N_13954,N_9677,N_10869);
nor U13955 (N_13955,N_12189,N_11967);
or U13956 (N_13956,N_11857,N_12346);
and U13957 (N_13957,N_10878,N_11319);
and U13958 (N_13958,N_12244,N_9673);
and U13959 (N_13959,N_11028,N_10468);
or U13960 (N_13960,N_10653,N_10234);
nor U13961 (N_13961,N_10073,N_11070);
xor U13962 (N_13962,N_9843,N_12417);
nor U13963 (N_13963,N_12474,N_9588);
and U13964 (N_13964,N_10154,N_11762);
xnor U13965 (N_13965,N_10156,N_11049);
xnor U13966 (N_13966,N_11494,N_12164);
and U13967 (N_13967,N_10330,N_11818);
nor U13968 (N_13968,N_12012,N_12100);
or U13969 (N_13969,N_12431,N_11182);
and U13970 (N_13970,N_10054,N_10248);
nor U13971 (N_13971,N_9383,N_11132);
nand U13972 (N_13972,N_12391,N_10019);
nand U13973 (N_13973,N_9705,N_11487);
or U13974 (N_13974,N_12360,N_11854);
xnor U13975 (N_13975,N_11657,N_11287);
or U13976 (N_13976,N_10351,N_11139);
and U13977 (N_13977,N_12153,N_9534);
nand U13978 (N_13978,N_12418,N_10399);
nand U13979 (N_13979,N_9517,N_12341);
nand U13980 (N_13980,N_11346,N_11254);
nand U13981 (N_13981,N_12129,N_11577);
nand U13982 (N_13982,N_11676,N_9919);
and U13983 (N_13983,N_9738,N_9976);
nand U13984 (N_13984,N_11195,N_11983);
xnor U13985 (N_13985,N_9757,N_10158);
nand U13986 (N_13986,N_11876,N_10817);
or U13987 (N_13987,N_11035,N_11608);
nor U13988 (N_13988,N_10927,N_9899);
or U13989 (N_13989,N_10753,N_11554);
xnor U13990 (N_13990,N_10456,N_11306);
xnor U13991 (N_13991,N_9717,N_11853);
xor U13992 (N_13992,N_12396,N_10271);
and U13993 (N_13993,N_12352,N_12010);
xor U13994 (N_13994,N_11916,N_11717);
xor U13995 (N_13995,N_10388,N_10592);
nand U13996 (N_13996,N_11318,N_10476);
nor U13997 (N_13997,N_12370,N_11863);
and U13998 (N_13998,N_9562,N_12038);
nand U13999 (N_13999,N_11259,N_9780);
and U14000 (N_14000,N_9882,N_11549);
nor U14001 (N_14001,N_11469,N_9982);
nand U14002 (N_14002,N_11759,N_10670);
nand U14003 (N_14003,N_12363,N_9577);
and U14004 (N_14004,N_11817,N_12090);
or U14005 (N_14005,N_12245,N_11750);
xor U14006 (N_14006,N_11300,N_11220);
and U14007 (N_14007,N_9550,N_9380);
and U14008 (N_14008,N_12047,N_9839);
and U14009 (N_14009,N_9647,N_10771);
nand U14010 (N_14010,N_12195,N_12083);
nand U14011 (N_14011,N_11678,N_10318);
xnor U14012 (N_14012,N_11208,N_10041);
nor U14013 (N_14013,N_10829,N_11956);
nor U14014 (N_14014,N_11552,N_10396);
xor U14015 (N_14015,N_11765,N_11066);
nor U14016 (N_14016,N_11368,N_12110);
nand U14017 (N_14017,N_11904,N_9624);
nand U14018 (N_14018,N_9804,N_10258);
xnor U14019 (N_14019,N_11390,N_10405);
or U14020 (N_14020,N_9675,N_10466);
or U14021 (N_14021,N_9788,N_11257);
or U14022 (N_14022,N_12158,N_10659);
nand U14023 (N_14023,N_12466,N_10733);
nand U14024 (N_14024,N_11163,N_9835);
or U14025 (N_14025,N_11290,N_10169);
xor U14026 (N_14026,N_11537,N_10402);
and U14027 (N_14027,N_12235,N_11651);
nor U14028 (N_14028,N_11835,N_9785);
xor U14029 (N_14029,N_12171,N_9480);
or U14030 (N_14030,N_11669,N_11042);
xor U14031 (N_14031,N_9436,N_12111);
nor U14032 (N_14032,N_11261,N_11039);
xnor U14033 (N_14033,N_12307,N_10047);
xnor U14034 (N_14034,N_11690,N_10385);
xor U14035 (N_14035,N_11246,N_12321);
nand U14036 (N_14036,N_12459,N_11591);
and U14037 (N_14037,N_11016,N_10309);
and U14038 (N_14038,N_9504,N_9773);
nor U14039 (N_14039,N_10360,N_12148);
nor U14040 (N_14040,N_10437,N_9989);
nor U14041 (N_14041,N_11408,N_9777);
or U14042 (N_14042,N_11294,N_11194);
nor U14043 (N_14043,N_10441,N_10537);
or U14044 (N_14044,N_11005,N_11971);
or U14045 (N_14045,N_11333,N_11686);
and U14046 (N_14046,N_12338,N_12172);
nand U14047 (N_14047,N_11183,N_9507);
and U14048 (N_14048,N_10220,N_11526);
or U14049 (N_14049,N_12356,N_11784);
nand U14050 (N_14050,N_10426,N_12400);
nor U14051 (N_14051,N_10104,N_10740);
nand U14052 (N_14052,N_11816,N_10973);
or U14053 (N_14053,N_11752,N_11909);
or U14054 (N_14054,N_11936,N_10269);
and U14055 (N_14055,N_10797,N_10695);
nor U14056 (N_14056,N_12183,N_11960);
xor U14057 (N_14057,N_9684,N_11337);
and U14058 (N_14058,N_9783,N_10638);
or U14059 (N_14059,N_9902,N_11237);
and U14060 (N_14060,N_9769,N_10724);
xnor U14061 (N_14061,N_12374,N_11056);
and U14062 (N_14062,N_11441,N_11057);
xnor U14063 (N_14063,N_10939,N_10485);
or U14064 (N_14064,N_11375,N_11022);
nand U14065 (N_14065,N_10230,N_11889);
nor U14066 (N_14066,N_10297,N_11864);
nand U14067 (N_14067,N_11549,N_10718);
or U14068 (N_14068,N_10061,N_10340);
nor U14069 (N_14069,N_9445,N_10251);
nand U14070 (N_14070,N_11551,N_11579);
xnor U14071 (N_14071,N_9973,N_10509);
nor U14072 (N_14072,N_10529,N_10786);
nand U14073 (N_14073,N_12055,N_11852);
and U14074 (N_14074,N_9710,N_10736);
or U14075 (N_14075,N_12047,N_11773);
xor U14076 (N_14076,N_10705,N_9480);
and U14077 (N_14077,N_12429,N_10922);
nand U14078 (N_14078,N_9382,N_9548);
or U14079 (N_14079,N_11258,N_12195);
or U14080 (N_14080,N_11254,N_10129);
or U14081 (N_14081,N_10454,N_9842);
nand U14082 (N_14082,N_9388,N_11750);
nand U14083 (N_14083,N_9661,N_10295);
nand U14084 (N_14084,N_11417,N_10099);
nand U14085 (N_14085,N_10452,N_11592);
xor U14086 (N_14086,N_9470,N_11805);
or U14087 (N_14087,N_9762,N_12248);
nand U14088 (N_14088,N_10408,N_9885);
nor U14089 (N_14089,N_12224,N_11838);
or U14090 (N_14090,N_11132,N_10996);
nand U14091 (N_14091,N_10066,N_11682);
xnor U14092 (N_14092,N_11207,N_11087);
xnor U14093 (N_14093,N_11825,N_11326);
and U14094 (N_14094,N_10068,N_10485);
nor U14095 (N_14095,N_9408,N_9934);
nand U14096 (N_14096,N_10763,N_10154);
or U14097 (N_14097,N_10647,N_12397);
or U14098 (N_14098,N_12159,N_10579);
nand U14099 (N_14099,N_11389,N_9463);
nor U14100 (N_14100,N_10858,N_11938);
and U14101 (N_14101,N_12140,N_11173);
nor U14102 (N_14102,N_11384,N_12424);
xor U14103 (N_14103,N_12187,N_10975);
or U14104 (N_14104,N_10728,N_10942);
nand U14105 (N_14105,N_10748,N_11775);
nor U14106 (N_14106,N_10437,N_11354);
nand U14107 (N_14107,N_9659,N_11363);
and U14108 (N_14108,N_9805,N_10580);
xnor U14109 (N_14109,N_10097,N_10750);
or U14110 (N_14110,N_11280,N_9645);
and U14111 (N_14111,N_10330,N_12022);
or U14112 (N_14112,N_9720,N_11252);
nor U14113 (N_14113,N_12037,N_11790);
xor U14114 (N_14114,N_10973,N_10418);
nor U14115 (N_14115,N_12133,N_12471);
nand U14116 (N_14116,N_10027,N_9972);
and U14117 (N_14117,N_11187,N_9858);
nor U14118 (N_14118,N_11460,N_10780);
nor U14119 (N_14119,N_10167,N_11998);
nand U14120 (N_14120,N_11759,N_11189);
or U14121 (N_14121,N_10413,N_11513);
and U14122 (N_14122,N_10149,N_10435);
and U14123 (N_14123,N_10110,N_11593);
or U14124 (N_14124,N_11367,N_10529);
and U14125 (N_14125,N_10588,N_10061);
or U14126 (N_14126,N_12350,N_11995);
xnor U14127 (N_14127,N_11430,N_12360);
nand U14128 (N_14128,N_10352,N_9619);
and U14129 (N_14129,N_9810,N_11526);
or U14130 (N_14130,N_9643,N_9742);
nand U14131 (N_14131,N_9906,N_10125);
and U14132 (N_14132,N_9971,N_11414);
or U14133 (N_14133,N_9763,N_11230);
nand U14134 (N_14134,N_12003,N_11273);
nor U14135 (N_14135,N_12317,N_12327);
nand U14136 (N_14136,N_10863,N_9559);
nor U14137 (N_14137,N_9505,N_10571);
xor U14138 (N_14138,N_10400,N_10865);
xor U14139 (N_14139,N_11865,N_12233);
xor U14140 (N_14140,N_11390,N_12270);
or U14141 (N_14141,N_9982,N_10534);
nand U14142 (N_14142,N_11169,N_9547);
xor U14143 (N_14143,N_10881,N_11680);
xor U14144 (N_14144,N_12313,N_10366);
or U14145 (N_14145,N_12382,N_12217);
nand U14146 (N_14146,N_9388,N_11432);
and U14147 (N_14147,N_9497,N_12465);
or U14148 (N_14148,N_11323,N_11382);
nor U14149 (N_14149,N_11653,N_9858);
or U14150 (N_14150,N_9526,N_12168);
nand U14151 (N_14151,N_10516,N_9431);
xor U14152 (N_14152,N_9597,N_10875);
and U14153 (N_14153,N_11858,N_9965);
and U14154 (N_14154,N_12050,N_10201);
and U14155 (N_14155,N_9404,N_10852);
nand U14156 (N_14156,N_11272,N_9782);
xor U14157 (N_14157,N_9749,N_10731);
nand U14158 (N_14158,N_10227,N_10150);
and U14159 (N_14159,N_10530,N_11693);
or U14160 (N_14160,N_11895,N_12008);
nand U14161 (N_14161,N_10711,N_12408);
and U14162 (N_14162,N_11784,N_9641);
or U14163 (N_14163,N_9758,N_10839);
nand U14164 (N_14164,N_10942,N_10920);
nand U14165 (N_14165,N_12447,N_10577);
or U14166 (N_14166,N_11397,N_10296);
or U14167 (N_14167,N_10061,N_11549);
nand U14168 (N_14168,N_10903,N_11496);
nor U14169 (N_14169,N_12182,N_9846);
nor U14170 (N_14170,N_11256,N_11223);
nand U14171 (N_14171,N_11411,N_9860);
or U14172 (N_14172,N_12168,N_10676);
nor U14173 (N_14173,N_9840,N_12105);
or U14174 (N_14174,N_10879,N_12041);
nor U14175 (N_14175,N_11091,N_9439);
or U14176 (N_14176,N_9536,N_11405);
xor U14177 (N_14177,N_11284,N_11113);
xnor U14178 (N_14178,N_10837,N_10997);
xor U14179 (N_14179,N_12200,N_11667);
and U14180 (N_14180,N_10397,N_9944);
or U14181 (N_14181,N_9583,N_12470);
nor U14182 (N_14182,N_10044,N_12023);
nor U14183 (N_14183,N_11976,N_11910);
xor U14184 (N_14184,N_11176,N_10793);
or U14185 (N_14185,N_9401,N_11519);
and U14186 (N_14186,N_11756,N_9857);
nand U14187 (N_14187,N_10402,N_10226);
and U14188 (N_14188,N_10933,N_10845);
or U14189 (N_14189,N_10222,N_11514);
or U14190 (N_14190,N_11591,N_11246);
xor U14191 (N_14191,N_11075,N_11691);
and U14192 (N_14192,N_11775,N_9411);
xor U14193 (N_14193,N_10779,N_9933);
or U14194 (N_14194,N_9800,N_11787);
nand U14195 (N_14195,N_12268,N_10104);
and U14196 (N_14196,N_9728,N_11095);
nor U14197 (N_14197,N_11372,N_11804);
nand U14198 (N_14198,N_9814,N_11193);
or U14199 (N_14199,N_11627,N_9724);
xnor U14200 (N_14200,N_10129,N_10370);
xnor U14201 (N_14201,N_11585,N_11485);
or U14202 (N_14202,N_12269,N_10767);
nor U14203 (N_14203,N_10986,N_10655);
nor U14204 (N_14204,N_11630,N_9436);
and U14205 (N_14205,N_12429,N_12367);
xnor U14206 (N_14206,N_11220,N_10838);
xor U14207 (N_14207,N_11258,N_10273);
or U14208 (N_14208,N_10252,N_9814);
nand U14209 (N_14209,N_11829,N_9750);
nand U14210 (N_14210,N_11624,N_11222);
nand U14211 (N_14211,N_10858,N_10136);
xor U14212 (N_14212,N_11550,N_10334);
xnor U14213 (N_14213,N_10421,N_9767);
nor U14214 (N_14214,N_10844,N_10246);
or U14215 (N_14215,N_12266,N_10709);
xnor U14216 (N_14216,N_10397,N_12164);
nor U14217 (N_14217,N_10586,N_11421);
nand U14218 (N_14218,N_10445,N_12286);
or U14219 (N_14219,N_10058,N_11124);
and U14220 (N_14220,N_10886,N_9403);
xnor U14221 (N_14221,N_10282,N_10495);
nor U14222 (N_14222,N_11942,N_11593);
xor U14223 (N_14223,N_11505,N_9584);
xor U14224 (N_14224,N_9470,N_10214);
nand U14225 (N_14225,N_11547,N_10523);
xor U14226 (N_14226,N_10684,N_9920);
nand U14227 (N_14227,N_10516,N_11589);
or U14228 (N_14228,N_9494,N_10170);
or U14229 (N_14229,N_10405,N_11741);
or U14230 (N_14230,N_12050,N_12481);
nor U14231 (N_14231,N_10445,N_9438);
nor U14232 (N_14232,N_12170,N_11955);
nand U14233 (N_14233,N_10269,N_12123);
or U14234 (N_14234,N_9580,N_9383);
or U14235 (N_14235,N_11787,N_10760);
and U14236 (N_14236,N_12173,N_10746);
nand U14237 (N_14237,N_10185,N_9501);
and U14238 (N_14238,N_11248,N_12438);
nand U14239 (N_14239,N_11534,N_10217);
and U14240 (N_14240,N_11330,N_12053);
xnor U14241 (N_14241,N_12104,N_10110);
nor U14242 (N_14242,N_9434,N_9961);
xnor U14243 (N_14243,N_12184,N_11271);
and U14244 (N_14244,N_9512,N_10524);
and U14245 (N_14245,N_11801,N_9765);
nor U14246 (N_14246,N_10034,N_9733);
nor U14247 (N_14247,N_12409,N_9377);
xor U14248 (N_14248,N_10040,N_11512);
and U14249 (N_14249,N_10865,N_9645);
nor U14250 (N_14250,N_12194,N_9839);
and U14251 (N_14251,N_10797,N_9935);
and U14252 (N_14252,N_11680,N_12313);
and U14253 (N_14253,N_11737,N_10306);
and U14254 (N_14254,N_11542,N_11877);
or U14255 (N_14255,N_9523,N_10209);
and U14256 (N_14256,N_10005,N_10736);
nor U14257 (N_14257,N_12424,N_9745);
nor U14258 (N_14258,N_11128,N_12458);
nand U14259 (N_14259,N_12379,N_11705);
nand U14260 (N_14260,N_10330,N_9965);
and U14261 (N_14261,N_11025,N_11606);
xnor U14262 (N_14262,N_11828,N_11939);
xnor U14263 (N_14263,N_10570,N_10294);
xor U14264 (N_14264,N_10947,N_9511);
xor U14265 (N_14265,N_10537,N_10925);
and U14266 (N_14266,N_10977,N_10171);
nand U14267 (N_14267,N_10193,N_11564);
nor U14268 (N_14268,N_12318,N_9987);
xnor U14269 (N_14269,N_9658,N_10989);
nor U14270 (N_14270,N_9882,N_11000);
and U14271 (N_14271,N_11539,N_10772);
and U14272 (N_14272,N_11709,N_12455);
and U14273 (N_14273,N_11220,N_9951);
and U14274 (N_14274,N_10722,N_11741);
and U14275 (N_14275,N_9891,N_10791);
and U14276 (N_14276,N_12479,N_12035);
nand U14277 (N_14277,N_9427,N_10113);
nor U14278 (N_14278,N_10287,N_9465);
or U14279 (N_14279,N_11668,N_10490);
and U14280 (N_14280,N_9816,N_9742);
or U14281 (N_14281,N_11174,N_9572);
or U14282 (N_14282,N_9775,N_11660);
xnor U14283 (N_14283,N_9777,N_10115);
nand U14284 (N_14284,N_9609,N_12390);
or U14285 (N_14285,N_11685,N_11479);
and U14286 (N_14286,N_10800,N_10666);
and U14287 (N_14287,N_12476,N_11954);
nand U14288 (N_14288,N_11442,N_10763);
and U14289 (N_14289,N_9461,N_10471);
nand U14290 (N_14290,N_10315,N_10804);
xor U14291 (N_14291,N_9953,N_10954);
nor U14292 (N_14292,N_9495,N_10834);
or U14293 (N_14293,N_10880,N_9517);
and U14294 (N_14294,N_9440,N_9826);
or U14295 (N_14295,N_11573,N_10267);
nor U14296 (N_14296,N_11985,N_12269);
nand U14297 (N_14297,N_9640,N_11252);
nor U14298 (N_14298,N_12241,N_12351);
xor U14299 (N_14299,N_10440,N_11727);
or U14300 (N_14300,N_12360,N_10022);
xnor U14301 (N_14301,N_10017,N_9829);
xor U14302 (N_14302,N_10761,N_9626);
or U14303 (N_14303,N_10767,N_11297);
nand U14304 (N_14304,N_12438,N_10546);
nand U14305 (N_14305,N_10557,N_11425);
and U14306 (N_14306,N_12450,N_10582);
nor U14307 (N_14307,N_10507,N_10614);
or U14308 (N_14308,N_11359,N_9584);
xnor U14309 (N_14309,N_10517,N_11941);
xor U14310 (N_14310,N_12359,N_11785);
and U14311 (N_14311,N_10069,N_10034);
xnor U14312 (N_14312,N_12253,N_10643);
and U14313 (N_14313,N_12183,N_12141);
nand U14314 (N_14314,N_9650,N_11391);
xor U14315 (N_14315,N_11158,N_12222);
and U14316 (N_14316,N_11575,N_11288);
nand U14317 (N_14317,N_10315,N_10371);
nor U14318 (N_14318,N_10048,N_11472);
or U14319 (N_14319,N_9980,N_11671);
and U14320 (N_14320,N_11023,N_10240);
xnor U14321 (N_14321,N_11967,N_11771);
xnor U14322 (N_14322,N_12275,N_12268);
nand U14323 (N_14323,N_9580,N_11792);
and U14324 (N_14324,N_11406,N_12186);
nand U14325 (N_14325,N_12276,N_11027);
nand U14326 (N_14326,N_11263,N_12478);
nand U14327 (N_14327,N_9388,N_10939);
nor U14328 (N_14328,N_11280,N_11153);
or U14329 (N_14329,N_12368,N_10804);
nor U14330 (N_14330,N_11339,N_11190);
and U14331 (N_14331,N_10098,N_10764);
nor U14332 (N_14332,N_11314,N_11229);
nor U14333 (N_14333,N_10704,N_11252);
nor U14334 (N_14334,N_12316,N_12034);
or U14335 (N_14335,N_10035,N_9474);
nor U14336 (N_14336,N_11944,N_11975);
or U14337 (N_14337,N_10708,N_11971);
xnor U14338 (N_14338,N_9974,N_11384);
nand U14339 (N_14339,N_10092,N_10617);
or U14340 (N_14340,N_12353,N_10058);
nor U14341 (N_14341,N_10733,N_12471);
or U14342 (N_14342,N_10191,N_12237);
and U14343 (N_14343,N_10580,N_11401);
nand U14344 (N_14344,N_12090,N_11262);
and U14345 (N_14345,N_11625,N_12480);
and U14346 (N_14346,N_9540,N_12182);
or U14347 (N_14347,N_11995,N_10117);
and U14348 (N_14348,N_9690,N_11374);
xor U14349 (N_14349,N_9731,N_10067);
and U14350 (N_14350,N_10050,N_11147);
or U14351 (N_14351,N_10870,N_11480);
nand U14352 (N_14352,N_11000,N_12003);
nand U14353 (N_14353,N_11954,N_11776);
xor U14354 (N_14354,N_12178,N_11681);
nor U14355 (N_14355,N_10564,N_10970);
and U14356 (N_14356,N_12027,N_10950);
or U14357 (N_14357,N_10097,N_12181);
nor U14358 (N_14358,N_9965,N_11154);
or U14359 (N_14359,N_10183,N_12348);
and U14360 (N_14360,N_11725,N_10010);
and U14361 (N_14361,N_10587,N_10830);
nand U14362 (N_14362,N_11761,N_10549);
xnor U14363 (N_14363,N_10986,N_10575);
and U14364 (N_14364,N_10410,N_12178);
nor U14365 (N_14365,N_11162,N_10720);
xnor U14366 (N_14366,N_11222,N_10144);
nor U14367 (N_14367,N_11903,N_12121);
and U14368 (N_14368,N_11790,N_12018);
nor U14369 (N_14369,N_9704,N_12470);
or U14370 (N_14370,N_10879,N_10052);
or U14371 (N_14371,N_10757,N_10279);
nand U14372 (N_14372,N_9908,N_11120);
nand U14373 (N_14373,N_12457,N_9981);
or U14374 (N_14374,N_9524,N_12375);
and U14375 (N_14375,N_10969,N_10768);
nor U14376 (N_14376,N_9444,N_11253);
nand U14377 (N_14377,N_11145,N_11471);
nand U14378 (N_14378,N_9432,N_9399);
and U14379 (N_14379,N_12010,N_10487);
nor U14380 (N_14380,N_11981,N_10589);
or U14381 (N_14381,N_11606,N_9478);
xnor U14382 (N_14382,N_12365,N_12120);
or U14383 (N_14383,N_12177,N_11670);
nand U14384 (N_14384,N_10363,N_9576);
nand U14385 (N_14385,N_11125,N_12337);
or U14386 (N_14386,N_10684,N_11773);
xor U14387 (N_14387,N_10576,N_9991);
xnor U14388 (N_14388,N_9557,N_10035);
xor U14389 (N_14389,N_12191,N_11477);
nor U14390 (N_14390,N_10665,N_9451);
and U14391 (N_14391,N_10859,N_10907);
or U14392 (N_14392,N_10342,N_10624);
nand U14393 (N_14393,N_12092,N_10284);
xnor U14394 (N_14394,N_12014,N_10731);
nor U14395 (N_14395,N_9907,N_12099);
or U14396 (N_14396,N_12434,N_12442);
xnor U14397 (N_14397,N_11575,N_10798);
or U14398 (N_14398,N_12336,N_11899);
nor U14399 (N_14399,N_11078,N_10083);
or U14400 (N_14400,N_9488,N_10627);
or U14401 (N_14401,N_11108,N_11566);
nand U14402 (N_14402,N_11302,N_11011);
and U14403 (N_14403,N_9956,N_12112);
xor U14404 (N_14404,N_11462,N_11410);
and U14405 (N_14405,N_12153,N_11068);
nand U14406 (N_14406,N_9483,N_11299);
xnor U14407 (N_14407,N_11958,N_10452);
and U14408 (N_14408,N_9817,N_10686);
nand U14409 (N_14409,N_12320,N_11946);
xnor U14410 (N_14410,N_10443,N_11639);
and U14411 (N_14411,N_9524,N_9819);
nand U14412 (N_14412,N_11876,N_11931);
or U14413 (N_14413,N_9425,N_12241);
nor U14414 (N_14414,N_10677,N_10074);
and U14415 (N_14415,N_12157,N_11415);
xor U14416 (N_14416,N_10451,N_10551);
nand U14417 (N_14417,N_11211,N_11675);
or U14418 (N_14418,N_10197,N_12328);
nand U14419 (N_14419,N_10982,N_11342);
or U14420 (N_14420,N_11184,N_9750);
nand U14421 (N_14421,N_9657,N_9628);
or U14422 (N_14422,N_10341,N_9999);
nor U14423 (N_14423,N_11865,N_12289);
xnor U14424 (N_14424,N_10285,N_10247);
and U14425 (N_14425,N_9540,N_11376);
and U14426 (N_14426,N_12241,N_11534);
nand U14427 (N_14427,N_10919,N_12288);
or U14428 (N_14428,N_10374,N_11435);
or U14429 (N_14429,N_11570,N_12200);
xnor U14430 (N_14430,N_11056,N_10272);
xor U14431 (N_14431,N_9553,N_9810);
nand U14432 (N_14432,N_11701,N_11947);
xnor U14433 (N_14433,N_11442,N_10113);
xor U14434 (N_14434,N_11980,N_11379);
nand U14435 (N_14435,N_10677,N_11950);
nand U14436 (N_14436,N_9642,N_9647);
or U14437 (N_14437,N_10089,N_12331);
nor U14438 (N_14438,N_11293,N_11495);
nand U14439 (N_14439,N_11042,N_11658);
nor U14440 (N_14440,N_12255,N_10754);
and U14441 (N_14441,N_10974,N_12331);
nor U14442 (N_14442,N_12240,N_10422);
and U14443 (N_14443,N_10479,N_10618);
nand U14444 (N_14444,N_10938,N_10623);
xnor U14445 (N_14445,N_10230,N_11424);
nand U14446 (N_14446,N_12340,N_10565);
nor U14447 (N_14447,N_9737,N_11315);
nand U14448 (N_14448,N_9968,N_10893);
nand U14449 (N_14449,N_11061,N_10886);
nand U14450 (N_14450,N_10825,N_10377);
nor U14451 (N_14451,N_11557,N_10028);
xnor U14452 (N_14452,N_10881,N_11545);
xnor U14453 (N_14453,N_10357,N_12275);
xor U14454 (N_14454,N_9670,N_9742);
and U14455 (N_14455,N_10585,N_10783);
nor U14456 (N_14456,N_11906,N_11307);
nand U14457 (N_14457,N_10935,N_9548);
and U14458 (N_14458,N_10208,N_10785);
and U14459 (N_14459,N_10297,N_10079);
xnor U14460 (N_14460,N_11853,N_11681);
and U14461 (N_14461,N_12182,N_11944);
nor U14462 (N_14462,N_12171,N_11526);
and U14463 (N_14463,N_11361,N_11516);
or U14464 (N_14464,N_10075,N_10185);
xnor U14465 (N_14465,N_11650,N_11118);
nand U14466 (N_14466,N_9466,N_10900);
nand U14467 (N_14467,N_10230,N_10968);
and U14468 (N_14468,N_11483,N_10895);
nand U14469 (N_14469,N_9879,N_11737);
or U14470 (N_14470,N_11890,N_11414);
xnor U14471 (N_14471,N_11582,N_10851);
nand U14472 (N_14472,N_10230,N_10602);
or U14473 (N_14473,N_10293,N_9513);
and U14474 (N_14474,N_10760,N_12256);
or U14475 (N_14475,N_11917,N_9977);
and U14476 (N_14476,N_9719,N_11549);
nand U14477 (N_14477,N_9679,N_10557);
xnor U14478 (N_14478,N_10053,N_10491);
and U14479 (N_14479,N_11000,N_11181);
or U14480 (N_14480,N_11937,N_12473);
nand U14481 (N_14481,N_11382,N_9858);
nand U14482 (N_14482,N_10984,N_12394);
or U14483 (N_14483,N_9784,N_11056);
nand U14484 (N_14484,N_9530,N_12207);
nand U14485 (N_14485,N_10520,N_9690);
xnor U14486 (N_14486,N_11908,N_9743);
xnor U14487 (N_14487,N_11102,N_12163);
and U14488 (N_14488,N_9937,N_11449);
or U14489 (N_14489,N_9393,N_9668);
and U14490 (N_14490,N_10092,N_12115);
nand U14491 (N_14491,N_10508,N_10374);
or U14492 (N_14492,N_10068,N_11259);
and U14493 (N_14493,N_9568,N_11245);
nor U14494 (N_14494,N_9784,N_11394);
nand U14495 (N_14495,N_12263,N_10105);
and U14496 (N_14496,N_12108,N_11516);
xnor U14497 (N_14497,N_10645,N_11254);
nor U14498 (N_14498,N_10381,N_12085);
or U14499 (N_14499,N_9575,N_10402);
nor U14500 (N_14500,N_10789,N_11439);
and U14501 (N_14501,N_9545,N_9463);
and U14502 (N_14502,N_12319,N_11430);
or U14503 (N_14503,N_9686,N_12054);
nor U14504 (N_14504,N_9563,N_11780);
nor U14505 (N_14505,N_10964,N_11456);
xor U14506 (N_14506,N_11783,N_10592);
nand U14507 (N_14507,N_10577,N_10448);
nor U14508 (N_14508,N_10406,N_11051);
nand U14509 (N_14509,N_10799,N_10419);
or U14510 (N_14510,N_9738,N_10288);
and U14511 (N_14511,N_11961,N_11101);
nor U14512 (N_14512,N_11449,N_11194);
xnor U14513 (N_14513,N_12006,N_11121);
nor U14514 (N_14514,N_9427,N_11002);
and U14515 (N_14515,N_9938,N_10263);
xnor U14516 (N_14516,N_9879,N_11186);
xnor U14517 (N_14517,N_11329,N_9470);
or U14518 (N_14518,N_11436,N_12063);
and U14519 (N_14519,N_9442,N_11610);
xor U14520 (N_14520,N_11132,N_10992);
or U14521 (N_14521,N_11205,N_10753);
nand U14522 (N_14522,N_12102,N_10785);
nand U14523 (N_14523,N_9919,N_11965);
nand U14524 (N_14524,N_11632,N_12165);
xor U14525 (N_14525,N_11064,N_9878);
and U14526 (N_14526,N_11238,N_12326);
xnor U14527 (N_14527,N_11968,N_12383);
and U14528 (N_14528,N_11210,N_9429);
nor U14529 (N_14529,N_12111,N_9897);
nand U14530 (N_14530,N_11466,N_11181);
nor U14531 (N_14531,N_11254,N_11168);
or U14532 (N_14532,N_10656,N_10112);
nor U14533 (N_14533,N_10478,N_12318);
nand U14534 (N_14534,N_10064,N_10690);
or U14535 (N_14535,N_12192,N_9923);
and U14536 (N_14536,N_12167,N_11910);
xnor U14537 (N_14537,N_11954,N_11759);
nor U14538 (N_14538,N_9610,N_11849);
nand U14539 (N_14539,N_10336,N_11058);
or U14540 (N_14540,N_9764,N_12358);
nand U14541 (N_14541,N_9769,N_10420);
or U14542 (N_14542,N_12330,N_10446);
nor U14543 (N_14543,N_11548,N_9822);
nor U14544 (N_14544,N_12270,N_11157);
or U14545 (N_14545,N_10803,N_10061);
nand U14546 (N_14546,N_11397,N_11826);
nor U14547 (N_14547,N_10945,N_11397);
nor U14548 (N_14548,N_11053,N_11698);
and U14549 (N_14549,N_10410,N_9828);
nor U14550 (N_14550,N_11863,N_11846);
or U14551 (N_14551,N_12403,N_11296);
and U14552 (N_14552,N_11345,N_10688);
nor U14553 (N_14553,N_10809,N_12106);
and U14554 (N_14554,N_10862,N_11958);
xor U14555 (N_14555,N_12006,N_10777);
nor U14556 (N_14556,N_10316,N_11935);
nand U14557 (N_14557,N_10571,N_11669);
nand U14558 (N_14558,N_11539,N_11088);
and U14559 (N_14559,N_10270,N_11547);
xnor U14560 (N_14560,N_9526,N_12272);
nand U14561 (N_14561,N_9695,N_12055);
or U14562 (N_14562,N_10111,N_11270);
nor U14563 (N_14563,N_12353,N_11539);
or U14564 (N_14564,N_11010,N_10530);
xnor U14565 (N_14565,N_9934,N_11218);
nand U14566 (N_14566,N_11868,N_12341);
or U14567 (N_14567,N_10020,N_12386);
xnor U14568 (N_14568,N_10394,N_11150);
and U14569 (N_14569,N_9727,N_11705);
nor U14570 (N_14570,N_10893,N_10287);
or U14571 (N_14571,N_11548,N_10467);
nand U14572 (N_14572,N_11340,N_10653);
or U14573 (N_14573,N_12338,N_11799);
and U14574 (N_14574,N_9952,N_12047);
nor U14575 (N_14575,N_12074,N_10374);
xor U14576 (N_14576,N_11819,N_10603);
or U14577 (N_14577,N_9889,N_10824);
or U14578 (N_14578,N_12403,N_10135);
xnor U14579 (N_14579,N_11600,N_10277);
nand U14580 (N_14580,N_9692,N_12210);
and U14581 (N_14581,N_12290,N_9603);
nand U14582 (N_14582,N_9508,N_10285);
nand U14583 (N_14583,N_11254,N_11796);
and U14584 (N_14584,N_9905,N_12024);
or U14585 (N_14585,N_10779,N_11838);
nand U14586 (N_14586,N_12186,N_12229);
and U14587 (N_14587,N_12345,N_9652);
nor U14588 (N_14588,N_10376,N_11851);
nand U14589 (N_14589,N_10068,N_10275);
nand U14590 (N_14590,N_10266,N_12137);
nand U14591 (N_14591,N_9973,N_10784);
or U14592 (N_14592,N_10609,N_9463);
xnor U14593 (N_14593,N_10776,N_11986);
xor U14594 (N_14594,N_11816,N_10729);
or U14595 (N_14595,N_10344,N_12199);
nor U14596 (N_14596,N_10149,N_10175);
xor U14597 (N_14597,N_9625,N_11520);
or U14598 (N_14598,N_11169,N_9392);
or U14599 (N_14599,N_9801,N_10782);
and U14600 (N_14600,N_9920,N_9424);
or U14601 (N_14601,N_9469,N_9876);
nor U14602 (N_14602,N_11839,N_10905);
and U14603 (N_14603,N_11564,N_11132);
nor U14604 (N_14604,N_9899,N_10175);
nor U14605 (N_14605,N_11313,N_12330);
or U14606 (N_14606,N_9782,N_9692);
and U14607 (N_14607,N_12216,N_10039);
xnor U14608 (N_14608,N_9780,N_9929);
nand U14609 (N_14609,N_11936,N_10918);
or U14610 (N_14610,N_9587,N_12236);
nor U14611 (N_14611,N_11703,N_12184);
or U14612 (N_14612,N_11477,N_11520);
xor U14613 (N_14613,N_10519,N_10525);
or U14614 (N_14614,N_10531,N_11804);
nor U14615 (N_14615,N_10687,N_10320);
nand U14616 (N_14616,N_11436,N_9673);
xor U14617 (N_14617,N_9537,N_11624);
xor U14618 (N_14618,N_11670,N_10020);
and U14619 (N_14619,N_12221,N_10098);
nor U14620 (N_14620,N_11305,N_11824);
xor U14621 (N_14621,N_11473,N_11200);
nor U14622 (N_14622,N_11082,N_12023);
nand U14623 (N_14623,N_9726,N_10868);
or U14624 (N_14624,N_11946,N_11523);
nor U14625 (N_14625,N_9852,N_12417);
nor U14626 (N_14626,N_10969,N_11805);
nand U14627 (N_14627,N_12385,N_10925);
nand U14628 (N_14628,N_10852,N_9447);
and U14629 (N_14629,N_11757,N_9899);
nor U14630 (N_14630,N_10410,N_9593);
xnor U14631 (N_14631,N_11069,N_10144);
nor U14632 (N_14632,N_10652,N_12184);
nor U14633 (N_14633,N_11466,N_12276);
and U14634 (N_14634,N_10951,N_11074);
nor U14635 (N_14635,N_12217,N_11560);
or U14636 (N_14636,N_11471,N_11899);
or U14637 (N_14637,N_11927,N_10315);
and U14638 (N_14638,N_11881,N_12228);
xnor U14639 (N_14639,N_11719,N_9932);
nor U14640 (N_14640,N_11268,N_10440);
nor U14641 (N_14641,N_10744,N_11444);
and U14642 (N_14642,N_11199,N_10051);
xor U14643 (N_14643,N_11457,N_10065);
nand U14644 (N_14644,N_11863,N_10082);
xor U14645 (N_14645,N_9509,N_12373);
nand U14646 (N_14646,N_11863,N_11103);
nor U14647 (N_14647,N_11873,N_11694);
nor U14648 (N_14648,N_9904,N_12150);
nand U14649 (N_14649,N_9444,N_9979);
xnor U14650 (N_14650,N_12114,N_10285);
nand U14651 (N_14651,N_11058,N_10301);
nand U14652 (N_14652,N_11704,N_11956);
or U14653 (N_14653,N_11383,N_12437);
xnor U14654 (N_14654,N_9381,N_10247);
and U14655 (N_14655,N_12220,N_10194);
or U14656 (N_14656,N_11159,N_11657);
xnor U14657 (N_14657,N_11278,N_10162);
nor U14658 (N_14658,N_11384,N_10163);
and U14659 (N_14659,N_9615,N_12215);
nor U14660 (N_14660,N_11237,N_11785);
or U14661 (N_14661,N_10273,N_10810);
nor U14662 (N_14662,N_12181,N_12159);
or U14663 (N_14663,N_9699,N_12283);
xor U14664 (N_14664,N_9876,N_9460);
nand U14665 (N_14665,N_10012,N_10767);
xor U14666 (N_14666,N_11327,N_11182);
and U14667 (N_14667,N_11796,N_11733);
or U14668 (N_14668,N_9478,N_12164);
and U14669 (N_14669,N_11573,N_12358);
nor U14670 (N_14670,N_11893,N_10919);
nor U14671 (N_14671,N_11082,N_12146);
xnor U14672 (N_14672,N_10157,N_9781);
or U14673 (N_14673,N_12053,N_11112);
xnor U14674 (N_14674,N_12376,N_9717);
nor U14675 (N_14675,N_12079,N_11353);
nor U14676 (N_14676,N_11218,N_9701);
xnor U14677 (N_14677,N_11046,N_10570);
xor U14678 (N_14678,N_11980,N_10794);
and U14679 (N_14679,N_10277,N_10958);
xnor U14680 (N_14680,N_11906,N_10739);
xnor U14681 (N_14681,N_12373,N_9805);
nand U14682 (N_14682,N_11798,N_10744);
nand U14683 (N_14683,N_9657,N_10392);
nor U14684 (N_14684,N_9688,N_10046);
xnor U14685 (N_14685,N_11514,N_11386);
xor U14686 (N_14686,N_11013,N_12183);
nor U14687 (N_14687,N_10039,N_10408);
and U14688 (N_14688,N_10297,N_10838);
and U14689 (N_14689,N_11891,N_11157);
xnor U14690 (N_14690,N_10749,N_10556);
nand U14691 (N_14691,N_11673,N_11106);
xnor U14692 (N_14692,N_10545,N_12412);
or U14693 (N_14693,N_12434,N_10938);
xor U14694 (N_14694,N_10523,N_11865);
xnor U14695 (N_14695,N_10055,N_11740);
nor U14696 (N_14696,N_11475,N_10887);
and U14697 (N_14697,N_10318,N_9941);
xnor U14698 (N_14698,N_12351,N_10373);
nor U14699 (N_14699,N_10586,N_11132);
or U14700 (N_14700,N_11778,N_11575);
nand U14701 (N_14701,N_12144,N_11929);
xnor U14702 (N_14702,N_10084,N_11344);
xnor U14703 (N_14703,N_10540,N_10605);
xor U14704 (N_14704,N_10691,N_11192);
xnor U14705 (N_14705,N_10029,N_11182);
xor U14706 (N_14706,N_11414,N_10519);
nor U14707 (N_14707,N_12268,N_12190);
xnor U14708 (N_14708,N_9967,N_10664);
and U14709 (N_14709,N_10685,N_12497);
or U14710 (N_14710,N_9987,N_9563);
and U14711 (N_14711,N_10521,N_10923);
nor U14712 (N_14712,N_9908,N_11466);
xnor U14713 (N_14713,N_12289,N_12478);
and U14714 (N_14714,N_10474,N_10415);
or U14715 (N_14715,N_11848,N_12346);
and U14716 (N_14716,N_11839,N_10397);
nand U14717 (N_14717,N_11755,N_12289);
nand U14718 (N_14718,N_9845,N_12207);
nor U14719 (N_14719,N_11370,N_10054);
nor U14720 (N_14720,N_9618,N_9767);
and U14721 (N_14721,N_9528,N_12216);
nand U14722 (N_14722,N_10129,N_11175);
xnor U14723 (N_14723,N_10541,N_10211);
xor U14724 (N_14724,N_11356,N_9792);
and U14725 (N_14725,N_11851,N_10892);
or U14726 (N_14726,N_10883,N_11320);
nor U14727 (N_14727,N_12193,N_9960);
nand U14728 (N_14728,N_12317,N_10104);
and U14729 (N_14729,N_12140,N_10401);
nand U14730 (N_14730,N_11589,N_9967);
nor U14731 (N_14731,N_11622,N_11000);
nor U14732 (N_14732,N_12417,N_11370);
and U14733 (N_14733,N_10921,N_10001);
xor U14734 (N_14734,N_10551,N_11824);
or U14735 (N_14735,N_11914,N_12240);
xor U14736 (N_14736,N_10584,N_12459);
and U14737 (N_14737,N_10635,N_12375);
xnor U14738 (N_14738,N_10586,N_11004);
nor U14739 (N_14739,N_11577,N_11322);
nor U14740 (N_14740,N_11553,N_11146);
nor U14741 (N_14741,N_9687,N_9864);
xnor U14742 (N_14742,N_11967,N_9734);
and U14743 (N_14743,N_10091,N_11978);
nor U14744 (N_14744,N_9611,N_10530);
nor U14745 (N_14745,N_9730,N_10204);
or U14746 (N_14746,N_9921,N_11886);
or U14747 (N_14747,N_11041,N_9783);
nand U14748 (N_14748,N_10594,N_12406);
xnor U14749 (N_14749,N_9610,N_11836);
nand U14750 (N_14750,N_11276,N_10496);
xnor U14751 (N_14751,N_9430,N_10386);
and U14752 (N_14752,N_9916,N_12266);
nor U14753 (N_14753,N_12347,N_11999);
nor U14754 (N_14754,N_11855,N_12135);
xnor U14755 (N_14755,N_9928,N_9709);
nor U14756 (N_14756,N_11840,N_11403);
nand U14757 (N_14757,N_12364,N_11629);
xor U14758 (N_14758,N_11079,N_10542);
xnor U14759 (N_14759,N_11311,N_11452);
and U14760 (N_14760,N_12124,N_10696);
or U14761 (N_14761,N_9488,N_12176);
and U14762 (N_14762,N_11084,N_9612);
nand U14763 (N_14763,N_11186,N_9876);
or U14764 (N_14764,N_9907,N_11917);
and U14765 (N_14765,N_10497,N_10024);
and U14766 (N_14766,N_11441,N_11830);
nand U14767 (N_14767,N_12269,N_11993);
xor U14768 (N_14768,N_9404,N_11948);
or U14769 (N_14769,N_11827,N_9814);
xor U14770 (N_14770,N_11060,N_9819);
nor U14771 (N_14771,N_11758,N_11226);
xor U14772 (N_14772,N_10642,N_9660);
and U14773 (N_14773,N_11502,N_12193);
xor U14774 (N_14774,N_9932,N_11407);
and U14775 (N_14775,N_11358,N_12436);
nor U14776 (N_14776,N_11531,N_11850);
and U14777 (N_14777,N_11688,N_12485);
xnor U14778 (N_14778,N_10761,N_9929);
nor U14779 (N_14779,N_11464,N_12347);
xor U14780 (N_14780,N_9525,N_10405);
nand U14781 (N_14781,N_10161,N_11679);
and U14782 (N_14782,N_10719,N_12455);
nand U14783 (N_14783,N_11465,N_11301);
and U14784 (N_14784,N_10478,N_9479);
nor U14785 (N_14785,N_9445,N_11151);
or U14786 (N_14786,N_10717,N_11061);
xnor U14787 (N_14787,N_11855,N_9541);
or U14788 (N_14788,N_10608,N_11723);
xor U14789 (N_14789,N_12049,N_9591);
xor U14790 (N_14790,N_9445,N_10478);
or U14791 (N_14791,N_11427,N_11221);
nor U14792 (N_14792,N_9897,N_10023);
nand U14793 (N_14793,N_11434,N_11778);
or U14794 (N_14794,N_12338,N_10923);
xnor U14795 (N_14795,N_11914,N_12153);
nand U14796 (N_14796,N_11459,N_10686);
nand U14797 (N_14797,N_9404,N_9854);
or U14798 (N_14798,N_11012,N_11035);
nand U14799 (N_14799,N_10832,N_9494);
xor U14800 (N_14800,N_10029,N_11701);
and U14801 (N_14801,N_11543,N_11876);
nor U14802 (N_14802,N_11127,N_11318);
and U14803 (N_14803,N_10351,N_10753);
and U14804 (N_14804,N_10456,N_12415);
and U14805 (N_14805,N_9410,N_11908);
nand U14806 (N_14806,N_10880,N_12439);
and U14807 (N_14807,N_11075,N_10564);
xor U14808 (N_14808,N_11446,N_12108);
or U14809 (N_14809,N_12001,N_11533);
or U14810 (N_14810,N_9581,N_10409);
nor U14811 (N_14811,N_11828,N_11008);
nand U14812 (N_14812,N_10617,N_9455);
nor U14813 (N_14813,N_11225,N_9611);
xor U14814 (N_14814,N_10050,N_10473);
or U14815 (N_14815,N_10651,N_11271);
or U14816 (N_14816,N_9807,N_10281);
nor U14817 (N_14817,N_11454,N_11480);
xor U14818 (N_14818,N_10341,N_11343);
or U14819 (N_14819,N_10405,N_9798);
nand U14820 (N_14820,N_9894,N_12450);
xnor U14821 (N_14821,N_10954,N_10097);
xnor U14822 (N_14822,N_10324,N_12221);
nor U14823 (N_14823,N_10066,N_11565);
nand U14824 (N_14824,N_10007,N_11724);
or U14825 (N_14825,N_10593,N_10023);
or U14826 (N_14826,N_11440,N_11240);
and U14827 (N_14827,N_12277,N_11384);
nor U14828 (N_14828,N_12287,N_10388);
nand U14829 (N_14829,N_10085,N_9774);
nor U14830 (N_14830,N_10771,N_11932);
and U14831 (N_14831,N_10570,N_9781);
or U14832 (N_14832,N_10784,N_9531);
nand U14833 (N_14833,N_12110,N_11775);
nand U14834 (N_14834,N_11010,N_10021);
nand U14835 (N_14835,N_11447,N_12205);
and U14836 (N_14836,N_11471,N_11529);
or U14837 (N_14837,N_10589,N_9555);
or U14838 (N_14838,N_10364,N_10421);
and U14839 (N_14839,N_10338,N_10516);
nor U14840 (N_14840,N_10714,N_11722);
and U14841 (N_14841,N_10558,N_11936);
xor U14842 (N_14842,N_9886,N_10327);
and U14843 (N_14843,N_12346,N_12212);
nor U14844 (N_14844,N_12027,N_12037);
and U14845 (N_14845,N_11278,N_10541);
and U14846 (N_14846,N_10678,N_11318);
and U14847 (N_14847,N_11342,N_10403);
nor U14848 (N_14848,N_12426,N_10403);
and U14849 (N_14849,N_12175,N_11744);
nand U14850 (N_14850,N_10062,N_9950);
and U14851 (N_14851,N_10082,N_9629);
nand U14852 (N_14852,N_11278,N_10438);
nand U14853 (N_14853,N_11302,N_11312);
or U14854 (N_14854,N_10963,N_9789);
and U14855 (N_14855,N_12307,N_11919);
nor U14856 (N_14856,N_12437,N_12220);
and U14857 (N_14857,N_9959,N_10190);
nor U14858 (N_14858,N_10718,N_11084);
and U14859 (N_14859,N_10945,N_11590);
xor U14860 (N_14860,N_9571,N_10254);
nor U14861 (N_14861,N_11629,N_12491);
or U14862 (N_14862,N_12298,N_11959);
nand U14863 (N_14863,N_11529,N_10719);
or U14864 (N_14864,N_11053,N_10885);
nand U14865 (N_14865,N_12103,N_11010);
nor U14866 (N_14866,N_11138,N_10654);
nor U14867 (N_14867,N_12293,N_11552);
nand U14868 (N_14868,N_10784,N_9600);
and U14869 (N_14869,N_9530,N_9791);
and U14870 (N_14870,N_9610,N_11204);
nand U14871 (N_14871,N_10377,N_10771);
xnor U14872 (N_14872,N_12323,N_10392);
and U14873 (N_14873,N_9968,N_11526);
and U14874 (N_14874,N_10825,N_10985);
nor U14875 (N_14875,N_11835,N_10075);
nand U14876 (N_14876,N_10882,N_10920);
nand U14877 (N_14877,N_11755,N_11456);
and U14878 (N_14878,N_12308,N_12256);
nand U14879 (N_14879,N_11059,N_9626);
and U14880 (N_14880,N_12066,N_12458);
or U14881 (N_14881,N_11184,N_11135);
or U14882 (N_14882,N_10324,N_12137);
or U14883 (N_14883,N_9903,N_11613);
nor U14884 (N_14884,N_10651,N_11061);
nand U14885 (N_14885,N_10212,N_9886);
xnor U14886 (N_14886,N_12000,N_10063);
and U14887 (N_14887,N_10327,N_11319);
and U14888 (N_14888,N_11144,N_10769);
nand U14889 (N_14889,N_10616,N_10161);
and U14890 (N_14890,N_11837,N_11703);
nor U14891 (N_14891,N_11487,N_9852);
and U14892 (N_14892,N_12409,N_11265);
or U14893 (N_14893,N_11929,N_10749);
or U14894 (N_14894,N_11315,N_9423);
xor U14895 (N_14895,N_9867,N_11665);
nand U14896 (N_14896,N_11606,N_9765);
nand U14897 (N_14897,N_9475,N_9427);
xnor U14898 (N_14898,N_10856,N_10918);
and U14899 (N_14899,N_11537,N_10947);
and U14900 (N_14900,N_10408,N_9491);
nor U14901 (N_14901,N_11765,N_11742);
and U14902 (N_14902,N_9764,N_11773);
or U14903 (N_14903,N_9584,N_10028);
nand U14904 (N_14904,N_9630,N_10382);
and U14905 (N_14905,N_12478,N_12369);
nor U14906 (N_14906,N_10088,N_10876);
and U14907 (N_14907,N_10182,N_10654);
nor U14908 (N_14908,N_12132,N_10800);
or U14909 (N_14909,N_10592,N_10922);
nand U14910 (N_14910,N_11258,N_11464);
nand U14911 (N_14911,N_11264,N_11065);
or U14912 (N_14912,N_10734,N_12490);
xnor U14913 (N_14913,N_11802,N_9704);
nor U14914 (N_14914,N_11267,N_11114);
and U14915 (N_14915,N_9984,N_11522);
nor U14916 (N_14916,N_12367,N_12242);
xnor U14917 (N_14917,N_10773,N_11500);
and U14918 (N_14918,N_12019,N_10959);
or U14919 (N_14919,N_11710,N_11598);
nand U14920 (N_14920,N_9443,N_11169);
nand U14921 (N_14921,N_10661,N_9805);
or U14922 (N_14922,N_10121,N_12292);
or U14923 (N_14923,N_12015,N_12451);
nand U14924 (N_14924,N_10464,N_12038);
nor U14925 (N_14925,N_11892,N_11535);
nor U14926 (N_14926,N_10960,N_9711);
nand U14927 (N_14927,N_11111,N_9642);
or U14928 (N_14928,N_12498,N_11611);
nand U14929 (N_14929,N_10438,N_10529);
and U14930 (N_14930,N_10050,N_11809);
nand U14931 (N_14931,N_12497,N_10410);
nand U14932 (N_14932,N_9640,N_11063);
and U14933 (N_14933,N_9541,N_11441);
nand U14934 (N_14934,N_12184,N_11548);
nor U14935 (N_14935,N_10719,N_10318);
nand U14936 (N_14936,N_12248,N_9804);
nand U14937 (N_14937,N_11011,N_11518);
or U14938 (N_14938,N_10516,N_9658);
or U14939 (N_14939,N_11937,N_12263);
nor U14940 (N_14940,N_12236,N_11851);
xor U14941 (N_14941,N_11574,N_11473);
xor U14942 (N_14942,N_11919,N_10217);
or U14943 (N_14943,N_10220,N_11952);
nor U14944 (N_14944,N_9877,N_11144);
xnor U14945 (N_14945,N_11032,N_9664);
nor U14946 (N_14946,N_11247,N_10805);
xnor U14947 (N_14947,N_12342,N_10586);
and U14948 (N_14948,N_12417,N_11383);
or U14949 (N_14949,N_11835,N_9406);
and U14950 (N_14950,N_9887,N_10913);
or U14951 (N_14951,N_9621,N_10338);
nor U14952 (N_14952,N_10852,N_11270);
and U14953 (N_14953,N_12182,N_9692);
and U14954 (N_14954,N_11662,N_11740);
xnor U14955 (N_14955,N_11694,N_11708);
nor U14956 (N_14956,N_9722,N_11873);
nand U14957 (N_14957,N_11900,N_10132);
nand U14958 (N_14958,N_9582,N_10062);
or U14959 (N_14959,N_11431,N_12362);
nor U14960 (N_14960,N_10209,N_12045);
xnor U14961 (N_14961,N_9901,N_11103);
xnor U14962 (N_14962,N_11443,N_10668);
nor U14963 (N_14963,N_9661,N_10703);
xnor U14964 (N_14964,N_9400,N_11304);
xor U14965 (N_14965,N_11364,N_11404);
nor U14966 (N_14966,N_12049,N_10845);
nand U14967 (N_14967,N_12352,N_9436);
xor U14968 (N_14968,N_9759,N_11603);
or U14969 (N_14969,N_11860,N_9644);
or U14970 (N_14970,N_12019,N_11955);
or U14971 (N_14971,N_11722,N_10944);
nor U14972 (N_14972,N_9992,N_10599);
nor U14973 (N_14973,N_11366,N_11811);
nand U14974 (N_14974,N_9616,N_10591);
nor U14975 (N_14975,N_9794,N_9661);
nand U14976 (N_14976,N_10672,N_11955);
nor U14977 (N_14977,N_12224,N_11566);
and U14978 (N_14978,N_11382,N_11818);
nor U14979 (N_14979,N_10611,N_11331);
nand U14980 (N_14980,N_10039,N_9674);
nor U14981 (N_14981,N_9588,N_12364);
nand U14982 (N_14982,N_12029,N_12052);
xor U14983 (N_14983,N_9655,N_12381);
nand U14984 (N_14984,N_9426,N_9492);
nor U14985 (N_14985,N_11506,N_11214);
xor U14986 (N_14986,N_11367,N_11776);
and U14987 (N_14987,N_12495,N_11924);
xor U14988 (N_14988,N_10474,N_11499);
and U14989 (N_14989,N_10258,N_9962);
or U14990 (N_14990,N_9754,N_10938);
xnor U14991 (N_14991,N_11389,N_10388);
xnor U14992 (N_14992,N_9832,N_12106);
xnor U14993 (N_14993,N_11490,N_9482);
and U14994 (N_14994,N_12466,N_9489);
or U14995 (N_14995,N_11841,N_10947);
or U14996 (N_14996,N_12266,N_12326);
nor U14997 (N_14997,N_9591,N_11549);
xnor U14998 (N_14998,N_9573,N_12352);
nand U14999 (N_14999,N_12369,N_12378);
xor U15000 (N_15000,N_9608,N_9839);
xnor U15001 (N_15001,N_10409,N_10915);
nand U15002 (N_15002,N_11867,N_10946);
nand U15003 (N_15003,N_11843,N_10488);
xnor U15004 (N_15004,N_12216,N_11964);
nor U15005 (N_15005,N_11023,N_10043);
nor U15006 (N_15006,N_11359,N_11739);
or U15007 (N_15007,N_11491,N_11238);
nor U15008 (N_15008,N_10082,N_12055);
xnor U15009 (N_15009,N_11521,N_11505);
xor U15010 (N_15010,N_12112,N_9758);
or U15011 (N_15011,N_12441,N_12336);
xor U15012 (N_15012,N_11339,N_10584);
or U15013 (N_15013,N_10829,N_11004);
or U15014 (N_15014,N_11815,N_12045);
or U15015 (N_15015,N_9775,N_9588);
or U15016 (N_15016,N_9830,N_12058);
xor U15017 (N_15017,N_11746,N_9690);
nand U15018 (N_15018,N_12347,N_11534);
nor U15019 (N_15019,N_10574,N_10742);
nand U15020 (N_15020,N_12151,N_10623);
nand U15021 (N_15021,N_11439,N_11068);
nor U15022 (N_15022,N_10653,N_11387);
xnor U15023 (N_15023,N_11621,N_9489);
nor U15024 (N_15024,N_12222,N_10935);
nor U15025 (N_15025,N_9870,N_11914);
or U15026 (N_15026,N_10735,N_9574);
and U15027 (N_15027,N_11081,N_9961);
nor U15028 (N_15028,N_12305,N_10067);
nand U15029 (N_15029,N_11897,N_12342);
and U15030 (N_15030,N_10961,N_10197);
xor U15031 (N_15031,N_11013,N_12068);
nor U15032 (N_15032,N_10550,N_10380);
or U15033 (N_15033,N_11302,N_11637);
xor U15034 (N_15034,N_11614,N_10191);
xor U15035 (N_15035,N_11570,N_10742);
and U15036 (N_15036,N_11678,N_10454);
nor U15037 (N_15037,N_10028,N_10373);
or U15038 (N_15038,N_11429,N_9480);
xnor U15039 (N_15039,N_11416,N_11621);
or U15040 (N_15040,N_9405,N_12153);
xor U15041 (N_15041,N_11513,N_9577);
nand U15042 (N_15042,N_11735,N_10523);
or U15043 (N_15043,N_11916,N_10694);
or U15044 (N_15044,N_9393,N_9656);
or U15045 (N_15045,N_10770,N_11697);
nor U15046 (N_15046,N_9551,N_11875);
and U15047 (N_15047,N_12198,N_12497);
xnor U15048 (N_15048,N_11202,N_12448);
xnor U15049 (N_15049,N_11267,N_10277);
nand U15050 (N_15050,N_10635,N_12395);
nor U15051 (N_15051,N_10520,N_12092);
nand U15052 (N_15052,N_10888,N_11388);
or U15053 (N_15053,N_11366,N_11901);
nor U15054 (N_15054,N_11446,N_9548);
xor U15055 (N_15055,N_10163,N_11410);
xnor U15056 (N_15056,N_11546,N_9529);
nor U15057 (N_15057,N_10324,N_9505);
and U15058 (N_15058,N_10400,N_12089);
xor U15059 (N_15059,N_11718,N_9914);
nand U15060 (N_15060,N_10160,N_12103);
and U15061 (N_15061,N_9390,N_11255);
and U15062 (N_15062,N_11588,N_11601);
or U15063 (N_15063,N_12101,N_11595);
nand U15064 (N_15064,N_11927,N_12062);
and U15065 (N_15065,N_10678,N_11947);
or U15066 (N_15066,N_11045,N_11718);
xnor U15067 (N_15067,N_11867,N_11025);
nor U15068 (N_15068,N_10895,N_11208);
or U15069 (N_15069,N_10003,N_9460);
nand U15070 (N_15070,N_11006,N_9980);
and U15071 (N_15071,N_11120,N_12254);
nor U15072 (N_15072,N_10067,N_11746);
and U15073 (N_15073,N_11824,N_11478);
or U15074 (N_15074,N_9536,N_10466);
or U15075 (N_15075,N_10436,N_10141);
nand U15076 (N_15076,N_10657,N_10662);
and U15077 (N_15077,N_10098,N_10349);
xor U15078 (N_15078,N_9486,N_10634);
xnor U15079 (N_15079,N_10175,N_11868);
or U15080 (N_15080,N_10006,N_10686);
nor U15081 (N_15081,N_11718,N_12208);
nor U15082 (N_15082,N_10000,N_10249);
nand U15083 (N_15083,N_9451,N_12395);
nand U15084 (N_15084,N_10364,N_11038);
nand U15085 (N_15085,N_12247,N_12195);
nand U15086 (N_15086,N_12178,N_10089);
nor U15087 (N_15087,N_9598,N_10054);
nor U15088 (N_15088,N_10414,N_9715);
xnor U15089 (N_15089,N_11526,N_9533);
and U15090 (N_15090,N_10545,N_9921);
nor U15091 (N_15091,N_12336,N_10268);
nand U15092 (N_15092,N_10964,N_10713);
or U15093 (N_15093,N_11241,N_10865);
nor U15094 (N_15094,N_9450,N_12043);
and U15095 (N_15095,N_11387,N_12184);
nor U15096 (N_15096,N_12393,N_11873);
and U15097 (N_15097,N_10353,N_10224);
or U15098 (N_15098,N_10966,N_11514);
or U15099 (N_15099,N_10333,N_9461);
nor U15100 (N_15100,N_11741,N_12118);
xor U15101 (N_15101,N_11821,N_11942);
nand U15102 (N_15102,N_10077,N_9406);
and U15103 (N_15103,N_10382,N_10818);
nor U15104 (N_15104,N_11245,N_11920);
and U15105 (N_15105,N_10662,N_9871);
and U15106 (N_15106,N_10051,N_10212);
or U15107 (N_15107,N_10286,N_10909);
nor U15108 (N_15108,N_10883,N_11073);
xor U15109 (N_15109,N_10102,N_10117);
xnor U15110 (N_15110,N_9391,N_9882);
or U15111 (N_15111,N_11830,N_12191);
or U15112 (N_15112,N_11559,N_11039);
and U15113 (N_15113,N_9505,N_10503);
and U15114 (N_15114,N_9754,N_10952);
or U15115 (N_15115,N_12202,N_12143);
and U15116 (N_15116,N_12381,N_9430);
xnor U15117 (N_15117,N_12487,N_11701);
nor U15118 (N_15118,N_9473,N_10125);
or U15119 (N_15119,N_11674,N_11425);
or U15120 (N_15120,N_11047,N_9436);
nor U15121 (N_15121,N_12031,N_11838);
nand U15122 (N_15122,N_11892,N_10591);
or U15123 (N_15123,N_10218,N_10584);
nand U15124 (N_15124,N_11988,N_10125);
nor U15125 (N_15125,N_9820,N_10597);
nand U15126 (N_15126,N_11422,N_12054);
nor U15127 (N_15127,N_12077,N_11355);
nand U15128 (N_15128,N_9391,N_11611);
nand U15129 (N_15129,N_9855,N_10077);
or U15130 (N_15130,N_11940,N_12180);
nand U15131 (N_15131,N_9573,N_11361);
nand U15132 (N_15132,N_9385,N_12219);
nor U15133 (N_15133,N_11861,N_10701);
or U15134 (N_15134,N_12002,N_10845);
nand U15135 (N_15135,N_11094,N_11485);
nor U15136 (N_15136,N_11286,N_12040);
xnor U15137 (N_15137,N_10887,N_12233);
nor U15138 (N_15138,N_9767,N_11051);
xor U15139 (N_15139,N_9597,N_9377);
and U15140 (N_15140,N_9400,N_10008);
nor U15141 (N_15141,N_11359,N_12350);
xor U15142 (N_15142,N_11907,N_10259);
nand U15143 (N_15143,N_9608,N_10701);
xor U15144 (N_15144,N_10951,N_11058);
and U15145 (N_15145,N_9651,N_11260);
nor U15146 (N_15146,N_11489,N_10645);
nand U15147 (N_15147,N_11612,N_10710);
or U15148 (N_15148,N_11263,N_11142);
or U15149 (N_15149,N_9616,N_12269);
and U15150 (N_15150,N_12071,N_9919);
xor U15151 (N_15151,N_10796,N_10497);
nor U15152 (N_15152,N_10055,N_11083);
or U15153 (N_15153,N_11199,N_12225);
xor U15154 (N_15154,N_11931,N_11930);
nor U15155 (N_15155,N_11672,N_12191);
nand U15156 (N_15156,N_12310,N_12386);
or U15157 (N_15157,N_10532,N_12401);
nand U15158 (N_15158,N_11664,N_11908);
nand U15159 (N_15159,N_9515,N_9736);
xor U15160 (N_15160,N_12057,N_9566);
nor U15161 (N_15161,N_11988,N_11135);
xnor U15162 (N_15162,N_10832,N_11806);
xnor U15163 (N_15163,N_11614,N_9381);
or U15164 (N_15164,N_9672,N_11886);
and U15165 (N_15165,N_9459,N_9718);
xnor U15166 (N_15166,N_9416,N_12019);
and U15167 (N_15167,N_11496,N_10516);
xor U15168 (N_15168,N_9516,N_11165);
nand U15169 (N_15169,N_10838,N_10028);
or U15170 (N_15170,N_11846,N_11106);
or U15171 (N_15171,N_10757,N_11627);
or U15172 (N_15172,N_12069,N_12404);
or U15173 (N_15173,N_10014,N_12187);
nor U15174 (N_15174,N_10184,N_9903);
nand U15175 (N_15175,N_10720,N_11448);
and U15176 (N_15176,N_9503,N_12293);
or U15177 (N_15177,N_10449,N_11460);
and U15178 (N_15178,N_9639,N_10617);
nor U15179 (N_15179,N_10063,N_10403);
xor U15180 (N_15180,N_9828,N_12072);
nand U15181 (N_15181,N_11753,N_10929);
and U15182 (N_15182,N_11347,N_9627);
xor U15183 (N_15183,N_10432,N_12476);
nand U15184 (N_15184,N_10485,N_9391);
nor U15185 (N_15185,N_10932,N_10692);
xnor U15186 (N_15186,N_11387,N_9557);
nor U15187 (N_15187,N_12432,N_12358);
nand U15188 (N_15188,N_10544,N_10778);
and U15189 (N_15189,N_10419,N_9830);
and U15190 (N_15190,N_10026,N_9679);
or U15191 (N_15191,N_10302,N_9553);
xor U15192 (N_15192,N_11053,N_10500);
or U15193 (N_15193,N_12143,N_11025);
and U15194 (N_15194,N_9718,N_9876);
nor U15195 (N_15195,N_12108,N_10719);
or U15196 (N_15196,N_11820,N_10335);
nand U15197 (N_15197,N_9695,N_11751);
and U15198 (N_15198,N_12493,N_10559);
nand U15199 (N_15199,N_11201,N_10124);
xnor U15200 (N_15200,N_10951,N_9454);
or U15201 (N_15201,N_11327,N_10556);
xor U15202 (N_15202,N_12066,N_10570);
and U15203 (N_15203,N_11050,N_11753);
or U15204 (N_15204,N_10138,N_10164);
or U15205 (N_15205,N_9961,N_10213);
xnor U15206 (N_15206,N_12348,N_11077);
nor U15207 (N_15207,N_10614,N_10433);
nand U15208 (N_15208,N_9552,N_9842);
xor U15209 (N_15209,N_10566,N_9687);
nand U15210 (N_15210,N_10135,N_9471);
nor U15211 (N_15211,N_10572,N_10996);
nand U15212 (N_15212,N_9590,N_10706);
or U15213 (N_15213,N_11106,N_9455);
xnor U15214 (N_15214,N_12363,N_11935);
nand U15215 (N_15215,N_10199,N_12333);
and U15216 (N_15216,N_9832,N_12220);
nor U15217 (N_15217,N_12001,N_9928);
or U15218 (N_15218,N_11459,N_9576);
or U15219 (N_15219,N_10709,N_9546);
nand U15220 (N_15220,N_11004,N_9528);
nand U15221 (N_15221,N_9418,N_10111);
nor U15222 (N_15222,N_9890,N_10883);
nor U15223 (N_15223,N_10005,N_11572);
or U15224 (N_15224,N_12451,N_11764);
nor U15225 (N_15225,N_12351,N_9449);
xnor U15226 (N_15226,N_12253,N_9778);
nor U15227 (N_15227,N_9733,N_10213);
nand U15228 (N_15228,N_9572,N_10004);
nor U15229 (N_15229,N_9868,N_11368);
or U15230 (N_15230,N_9703,N_12056);
and U15231 (N_15231,N_10984,N_11756);
nand U15232 (N_15232,N_9830,N_9928);
xor U15233 (N_15233,N_9768,N_12178);
nand U15234 (N_15234,N_10231,N_9695);
and U15235 (N_15235,N_11898,N_12476);
xnor U15236 (N_15236,N_11590,N_11437);
xor U15237 (N_15237,N_10468,N_11405);
xor U15238 (N_15238,N_10815,N_11720);
xor U15239 (N_15239,N_9787,N_11085);
or U15240 (N_15240,N_11601,N_11924);
and U15241 (N_15241,N_9514,N_12115);
xnor U15242 (N_15242,N_10776,N_10938);
and U15243 (N_15243,N_9414,N_10158);
nand U15244 (N_15244,N_11414,N_10009);
nor U15245 (N_15245,N_11366,N_10889);
xor U15246 (N_15246,N_11385,N_11188);
and U15247 (N_15247,N_10818,N_11484);
and U15248 (N_15248,N_9844,N_9473);
nor U15249 (N_15249,N_12249,N_10144);
and U15250 (N_15250,N_12107,N_9851);
or U15251 (N_15251,N_11191,N_10438);
nor U15252 (N_15252,N_11598,N_9574);
nor U15253 (N_15253,N_12415,N_10275);
nand U15254 (N_15254,N_12051,N_10880);
and U15255 (N_15255,N_11552,N_11870);
and U15256 (N_15256,N_12296,N_11455);
and U15257 (N_15257,N_11528,N_11460);
nor U15258 (N_15258,N_11036,N_12433);
or U15259 (N_15259,N_11621,N_10360);
or U15260 (N_15260,N_11470,N_11494);
xor U15261 (N_15261,N_11393,N_11827);
nor U15262 (N_15262,N_11504,N_10520);
and U15263 (N_15263,N_11386,N_10041);
or U15264 (N_15264,N_11663,N_10811);
xnor U15265 (N_15265,N_10443,N_10134);
nor U15266 (N_15266,N_12296,N_10841);
and U15267 (N_15267,N_11043,N_10511);
nand U15268 (N_15268,N_11595,N_12367);
xor U15269 (N_15269,N_12198,N_11008);
xor U15270 (N_15270,N_9440,N_12061);
and U15271 (N_15271,N_10047,N_9693);
nand U15272 (N_15272,N_11093,N_11148);
and U15273 (N_15273,N_10272,N_12115);
xor U15274 (N_15274,N_12372,N_9810);
xor U15275 (N_15275,N_11462,N_11319);
nor U15276 (N_15276,N_11590,N_11921);
xnor U15277 (N_15277,N_9388,N_9841);
nand U15278 (N_15278,N_10846,N_11225);
xnor U15279 (N_15279,N_12081,N_10708);
or U15280 (N_15280,N_10332,N_10277);
xor U15281 (N_15281,N_11719,N_10089);
or U15282 (N_15282,N_11917,N_9539);
nand U15283 (N_15283,N_11897,N_11007);
nand U15284 (N_15284,N_11884,N_11797);
nand U15285 (N_15285,N_9991,N_9703);
nor U15286 (N_15286,N_12346,N_10276);
and U15287 (N_15287,N_10768,N_12069);
nor U15288 (N_15288,N_10939,N_9907);
nor U15289 (N_15289,N_12356,N_11463);
or U15290 (N_15290,N_12379,N_12156);
xnor U15291 (N_15291,N_11358,N_10398);
or U15292 (N_15292,N_9873,N_11480);
and U15293 (N_15293,N_10469,N_12055);
xor U15294 (N_15294,N_10979,N_10126);
and U15295 (N_15295,N_12401,N_11753);
nor U15296 (N_15296,N_11143,N_9601);
nand U15297 (N_15297,N_10068,N_9430);
nand U15298 (N_15298,N_11613,N_12092);
nor U15299 (N_15299,N_9429,N_12061);
nor U15300 (N_15300,N_11858,N_11423);
and U15301 (N_15301,N_12438,N_10125);
xnor U15302 (N_15302,N_11903,N_11464);
nand U15303 (N_15303,N_9637,N_9436);
or U15304 (N_15304,N_11194,N_11273);
and U15305 (N_15305,N_9516,N_11413);
or U15306 (N_15306,N_12098,N_9469);
nand U15307 (N_15307,N_12396,N_9619);
or U15308 (N_15308,N_10942,N_11394);
xor U15309 (N_15309,N_10483,N_12090);
nor U15310 (N_15310,N_9507,N_11907);
xnor U15311 (N_15311,N_12279,N_11446);
xnor U15312 (N_15312,N_10614,N_10855);
nand U15313 (N_15313,N_11205,N_12481);
and U15314 (N_15314,N_11607,N_10846);
or U15315 (N_15315,N_9545,N_10257);
nand U15316 (N_15316,N_11239,N_9895);
nand U15317 (N_15317,N_9903,N_12064);
and U15318 (N_15318,N_11929,N_11556);
and U15319 (N_15319,N_10830,N_9718);
or U15320 (N_15320,N_12455,N_10346);
nand U15321 (N_15321,N_10220,N_10804);
nand U15322 (N_15322,N_12370,N_11730);
and U15323 (N_15323,N_11952,N_9455);
xnor U15324 (N_15324,N_11171,N_10632);
and U15325 (N_15325,N_10076,N_9950);
xor U15326 (N_15326,N_10174,N_12051);
xor U15327 (N_15327,N_9492,N_10870);
nand U15328 (N_15328,N_9388,N_9803);
nand U15329 (N_15329,N_11359,N_10064);
nand U15330 (N_15330,N_9418,N_11808);
nor U15331 (N_15331,N_11568,N_10952);
nor U15332 (N_15332,N_11105,N_12222);
nor U15333 (N_15333,N_11828,N_11065);
or U15334 (N_15334,N_11661,N_11027);
nand U15335 (N_15335,N_10176,N_9582);
and U15336 (N_15336,N_9827,N_12485);
xnor U15337 (N_15337,N_9755,N_9384);
nand U15338 (N_15338,N_10596,N_11539);
xnor U15339 (N_15339,N_12198,N_10479);
nor U15340 (N_15340,N_9433,N_10863);
xor U15341 (N_15341,N_11532,N_9945);
nor U15342 (N_15342,N_12035,N_10655);
nand U15343 (N_15343,N_10024,N_10229);
xor U15344 (N_15344,N_11815,N_10021);
and U15345 (N_15345,N_10007,N_11277);
nor U15346 (N_15346,N_10431,N_10006);
or U15347 (N_15347,N_11367,N_11134);
nor U15348 (N_15348,N_12468,N_11266);
nand U15349 (N_15349,N_11090,N_11080);
nand U15350 (N_15350,N_10174,N_9674);
xor U15351 (N_15351,N_10429,N_9442);
or U15352 (N_15352,N_10654,N_9742);
and U15353 (N_15353,N_10017,N_10118);
nor U15354 (N_15354,N_11006,N_11841);
and U15355 (N_15355,N_11925,N_11492);
xor U15356 (N_15356,N_10364,N_12195);
or U15357 (N_15357,N_12046,N_12048);
and U15358 (N_15358,N_11844,N_11827);
nor U15359 (N_15359,N_10478,N_10699);
nor U15360 (N_15360,N_9400,N_11906);
nor U15361 (N_15361,N_11520,N_10541);
and U15362 (N_15362,N_9526,N_12226);
and U15363 (N_15363,N_11007,N_9898);
nand U15364 (N_15364,N_9484,N_11131);
or U15365 (N_15365,N_12162,N_10039);
and U15366 (N_15366,N_11162,N_9734);
xor U15367 (N_15367,N_9926,N_10496);
and U15368 (N_15368,N_10659,N_9768);
xnor U15369 (N_15369,N_9966,N_10036);
nand U15370 (N_15370,N_9501,N_10988);
nor U15371 (N_15371,N_12442,N_9772);
nand U15372 (N_15372,N_11165,N_10699);
nand U15373 (N_15373,N_11431,N_10191);
xor U15374 (N_15374,N_11130,N_10874);
nor U15375 (N_15375,N_10524,N_10660);
nand U15376 (N_15376,N_12200,N_10679);
xor U15377 (N_15377,N_12196,N_10550);
or U15378 (N_15378,N_11941,N_11800);
or U15379 (N_15379,N_11645,N_11384);
xor U15380 (N_15380,N_9601,N_11300);
and U15381 (N_15381,N_9918,N_10598);
and U15382 (N_15382,N_11111,N_11363);
xor U15383 (N_15383,N_9743,N_11476);
or U15384 (N_15384,N_10151,N_10221);
or U15385 (N_15385,N_10722,N_10587);
nand U15386 (N_15386,N_11899,N_11585);
nand U15387 (N_15387,N_12000,N_10602);
nor U15388 (N_15388,N_9740,N_11469);
nor U15389 (N_15389,N_12181,N_10010);
or U15390 (N_15390,N_10541,N_9490);
nand U15391 (N_15391,N_12345,N_11366);
or U15392 (N_15392,N_10146,N_11645);
xor U15393 (N_15393,N_11028,N_9522);
or U15394 (N_15394,N_10695,N_11130);
or U15395 (N_15395,N_11641,N_12152);
xnor U15396 (N_15396,N_10548,N_9864);
nor U15397 (N_15397,N_10673,N_11630);
nand U15398 (N_15398,N_9877,N_10857);
nor U15399 (N_15399,N_11649,N_11534);
xor U15400 (N_15400,N_10515,N_9677);
xnor U15401 (N_15401,N_10968,N_10696);
nand U15402 (N_15402,N_10190,N_10766);
nand U15403 (N_15403,N_12007,N_10780);
nor U15404 (N_15404,N_11141,N_10292);
and U15405 (N_15405,N_11847,N_11968);
or U15406 (N_15406,N_11438,N_11837);
nand U15407 (N_15407,N_11991,N_9974);
xor U15408 (N_15408,N_11419,N_11145);
or U15409 (N_15409,N_11058,N_9908);
and U15410 (N_15410,N_10229,N_10779);
or U15411 (N_15411,N_12308,N_10283);
nor U15412 (N_15412,N_11611,N_11553);
or U15413 (N_15413,N_11698,N_10886);
and U15414 (N_15414,N_10401,N_11840);
or U15415 (N_15415,N_10657,N_11803);
nor U15416 (N_15416,N_10406,N_9779);
xor U15417 (N_15417,N_10781,N_9628);
xor U15418 (N_15418,N_12197,N_11984);
nand U15419 (N_15419,N_12385,N_9538);
and U15420 (N_15420,N_12122,N_9961);
and U15421 (N_15421,N_12363,N_10330);
and U15422 (N_15422,N_12023,N_10185);
or U15423 (N_15423,N_11214,N_11751);
nor U15424 (N_15424,N_10233,N_11518);
nand U15425 (N_15425,N_11039,N_10949);
or U15426 (N_15426,N_9413,N_12417);
and U15427 (N_15427,N_12011,N_11512);
and U15428 (N_15428,N_9387,N_9446);
xnor U15429 (N_15429,N_10660,N_10492);
nand U15430 (N_15430,N_10173,N_12264);
and U15431 (N_15431,N_11353,N_11289);
nor U15432 (N_15432,N_10827,N_9428);
and U15433 (N_15433,N_10524,N_11652);
or U15434 (N_15434,N_9563,N_9376);
and U15435 (N_15435,N_10746,N_12029);
nand U15436 (N_15436,N_10057,N_10980);
or U15437 (N_15437,N_9401,N_11997);
and U15438 (N_15438,N_12169,N_11369);
nand U15439 (N_15439,N_11994,N_9997);
or U15440 (N_15440,N_9388,N_10052);
nand U15441 (N_15441,N_10420,N_10417);
and U15442 (N_15442,N_10842,N_11231);
or U15443 (N_15443,N_12428,N_9830);
nand U15444 (N_15444,N_9796,N_10180);
xor U15445 (N_15445,N_9957,N_10952);
nand U15446 (N_15446,N_11054,N_10207);
nor U15447 (N_15447,N_12225,N_10147);
nand U15448 (N_15448,N_10519,N_10598);
nor U15449 (N_15449,N_9442,N_12235);
nand U15450 (N_15450,N_9403,N_10168);
nand U15451 (N_15451,N_11074,N_10609);
nand U15452 (N_15452,N_10240,N_12000);
xnor U15453 (N_15453,N_11677,N_10748);
or U15454 (N_15454,N_10309,N_11421);
or U15455 (N_15455,N_10024,N_12389);
xor U15456 (N_15456,N_12125,N_10061);
nand U15457 (N_15457,N_11267,N_11747);
or U15458 (N_15458,N_10666,N_10158);
and U15459 (N_15459,N_11868,N_10389);
and U15460 (N_15460,N_11839,N_10749);
and U15461 (N_15461,N_11518,N_12241);
nand U15462 (N_15462,N_11453,N_9637);
nor U15463 (N_15463,N_10717,N_10226);
nand U15464 (N_15464,N_12155,N_11901);
and U15465 (N_15465,N_11305,N_12005);
nor U15466 (N_15466,N_10440,N_10938);
nand U15467 (N_15467,N_11896,N_11343);
nor U15468 (N_15468,N_10934,N_11170);
nor U15469 (N_15469,N_10248,N_10545);
and U15470 (N_15470,N_10550,N_10221);
nand U15471 (N_15471,N_12377,N_10849);
xnor U15472 (N_15472,N_9409,N_11727);
and U15473 (N_15473,N_11995,N_11652);
nand U15474 (N_15474,N_10230,N_9712);
nand U15475 (N_15475,N_9497,N_11590);
xor U15476 (N_15476,N_10114,N_10628);
nand U15477 (N_15477,N_10714,N_11017);
and U15478 (N_15478,N_11089,N_12253);
nor U15479 (N_15479,N_9910,N_12050);
and U15480 (N_15480,N_10639,N_12494);
or U15481 (N_15481,N_11156,N_10809);
and U15482 (N_15482,N_11357,N_10635);
or U15483 (N_15483,N_10507,N_11081);
nor U15484 (N_15484,N_10467,N_12190);
or U15485 (N_15485,N_10347,N_10699);
or U15486 (N_15486,N_10083,N_12004);
xor U15487 (N_15487,N_10238,N_12329);
nor U15488 (N_15488,N_11267,N_11752);
and U15489 (N_15489,N_11529,N_10959);
or U15490 (N_15490,N_10737,N_12114);
xor U15491 (N_15491,N_12484,N_9976);
nor U15492 (N_15492,N_10784,N_9496);
nand U15493 (N_15493,N_12417,N_11460);
or U15494 (N_15494,N_11771,N_11953);
nand U15495 (N_15495,N_10450,N_11503);
or U15496 (N_15496,N_11521,N_10491);
and U15497 (N_15497,N_10582,N_12169);
xor U15498 (N_15498,N_10867,N_10076);
nor U15499 (N_15499,N_9873,N_10496);
nor U15500 (N_15500,N_11030,N_11821);
nor U15501 (N_15501,N_12444,N_9708);
or U15502 (N_15502,N_11545,N_10056);
xor U15503 (N_15503,N_9761,N_9816);
nor U15504 (N_15504,N_9712,N_10220);
nor U15505 (N_15505,N_10980,N_11796);
nand U15506 (N_15506,N_11858,N_9886);
nand U15507 (N_15507,N_11598,N_10941);
and U15508 (N_15508,N_10372,N_10767);
and U15509 (N_15509,N_12134,N_10558);
or U15510 (N_15510,N_10046,N_9936);
nand U15511 (N_15511,N_10052,N_11679);
nor U15512 (N_15512,N_10001,N_12231);
nand U15513 (N_15513,N_10342,N_10270);
xnor U15514 (N_15514,N_11760,N_9633);
or U15515 (N_15515,N_10901,N_10657);
nand U15516 (N_15516,N_10393,N_11681);
xnor U15517 (N_15517,N_12036,N_11170);
or U15518 (N_15518,N_12283,N_10107);
nand U15519 (N_15519,N_12431,N_10083);
or U15520 (N_15520,N_9773,N_9787);
or U15521 (N_15521,N_10790,N_9827);
and U15522 (N_15522,N_10812,N_9659);
and U15523 (N_15523,N_12372,N_12094);
nor U15524 (N_15524,N_11991,N_9795);
nand U15525 (N_15525,N_9463,N_12498);
and U15526 (N_15526,N_10026,N_10364);
and U15527 (N_15527,N_10287,N_10370);
xor U15528 (N_15528,N_9844,N_9448);
or U15529 (N_15529,N_11720,N_9566);
or U15530 (N_15530,N_9951,N_10071);
xnor U15531 (N_15531,N_12344,N_9926);
and U15532 (N_15532,N_10795,N_10642);
xnor U15533 (N_15533,N_9796,N_11584);
nand U15534 (N_15534,N_12102,N_11326);
or U15535 (N_15535,N_11633,N_10695);
or U15536 (N_15536,N_11227,N_11998);
nor U15537 (N_15537,N_11970,N_11809);
or U15538 (N_15538,N_11230,N_11576);
nand U15539 (N_15539,N_11883,N_11495);
xor U15540 (N_15540,N_10379,N_10382);
and U15541 (N_15541,N_12312,N_10312);
nor U15542 (N_15542,N_10201,N_11253);
xnor U15543 (N_15543,N_10341,N_11010);
nor U15544 (N_15544,N_10533,N_12037);
and U15545 (N_15545,N_10192,N_10664);
nand U15546 (N_15546,N_12223,N_12244);
nand U15547 (N_15547,N_11362,N_10691);
nor U15548 (N_15548,N_9537,N_9986);
and U15549 (N_15549,N_10672,N_12425);
or U15550 (N_15550,N_11467,N_11621);
and U15551 (N_15551,N_11430,N_9521);
xnor U15552 (N_15552,N_11740,N_12040);
xnor U15553 (N_15553,N_11107,N_11228);
nor U15554 (N_15554,N_9981,N_9629);
nand U15555 (N_15555,N_10356,N_11697);
xnor U15556 (N_15556,N_10308,N_10154);
xnor U15557 (N_15557,N_10667,N_9549);
xor U15558 (N_15558,N_11230,N_10036);
or U15559 (N_15559,N_11381,N_10472);
or U15560 (N_15560,N_12122,N_10937);
and U15561 (N_15561,N_10413,N_11543);
or U15562 (N_15562,N_11674,N_12064);
and U15563 (N_15563,N_9454,N_10162);
nor U15564 (N_15564,N_11186,N_9555);
xor U15565 (N_15565,N_10080,N_11336);
nand U15566 (N_15566,N_10013,N_9844);
and U15567 (N_15567,N_9682,N_12299);
nor U15568 (N_15568,N_11624,N_9610);
and U15569 (N_15569,N_10073,N_10238);
nor U15570 (N_15570,N_12152,N_10555);
nor U15571 (N_15571,N_10057,N_11662);
nor U15572 (N_15572,N_12293,N_11606);
nand U15573 (N_15573,N_9820,N_10191);
nor U15574 (N_15574,N_11321,N_11045);
nand U15575 (N_15575,N_10010,N_9643);
or U15576 (N_15576,N_10070,N_10771);
and U15577 (N_15577,N_11346,N_10231);
nand U15578 (N_15578,N_12220,N_11751);
nand U15579 (N_15579,N_10157,N_10340);
or U15580 (N_15580,N_10650,N_11402);
xnor U15581 (N_15581,N_11760,N_11781);
xnor U15582 (N_15582,N_10391,N_11386);
and U15583 (N_15583,N_9965,N_12399);
nor U15584 (N_15584,N_9650,N_11962);
nor U15585 (N_15585,N_9797,N_10989);
nor U15586 (N_15586,N_11027,N_10729);
nor U15587 (N_15587,N_10663,N_9473);
nor U15588 (N_15588,N_12360,N_10044);
xor U15589 (N_15589,N_12395,N_11425);
xor U15590 (N_15590,N_11091,N_9477);
nand U15591 (N_15591,N_12065,N_12045);
nor U15592 (N_15592,N_12254,N_10435);
or U15593 (N_15593,N_10106,N_11800);
xor U15594 (N_15594,N_11588,N_9721);
xor U15595 (N_15595,N_10374,N_12312);
xnor U15596 (N_15596,N_10122,N_11983);
xnor U15597 (N_15597,N_9869,N_10007);
nor U15598 (N_15598,N_10256,N_9711);
and U15599 (N_15599,N_11294,N_10040);
nor U15600 (N_15600,N_11431,N_12010);
and U15601 (N_15601,N_11891,N_10725);
nand U15602 (N_15602,N_10120,N_9719);
xor U15603 (N_15603,N_10360,N_11930);
xor U15604 (N_15604,N_11338,N_11266);
nor U15605 (N_15605,N_9914,N_10960);
nor U15606 (N_15606,N_11773,N_9893);
nand U15607 (N_15607,N_12327,N_10736);
and U15608 (N_15608,N_10038,N_10472);
nand U15609 (N_15609,N_12410,N_9674);
or U15610 (N_15610,N_12249,N_11752);
nor U15611 (N_15611,N_12167,N_10025);
xnor U15612 (N_15612,N_11318,N_11850);
or U15613 (N_15613,N_12471,N_9746);
nor U15614 (N_15614,N_10807,N_12172);
or U15615 (N_15615,N_9817,N_9997);
xnor U15616 (N_15616,N_12354,N_12298);
and U15617 (N_15617,N_9462,N_10689);
or U15618 (N_15618,N_12152,N_11692);
or U15619 (N_15619,N_10899,N_11808);
nand U15620 (N_15620,N_11518,N_10889);
or U15621 (N_15621,N_10357,N_9878);
or U15622 (N_15622,N_11671,N_12044);
or U15623 (N_15623,N_10363,N_10708);
or U15624 (N_15624,N_12417,N_10154);
xnor U15625 (N_15625,N_13148,N_13745);
nor U15626 (N_15626,N_13957,N_15370);
nand U15627 (N_15627,N_14420,N_12640);
xor U15628 (N_15628,N_13811,N_14626);
or U15629 (N_15629,N_13255,N_15249);
or U15630 (N_15630,N_13119,N_14832);
nor U15631 (N_15631,N_12802,N_12558);
nor U15632 (N_15632,N_14559,N_14442);
xnor U15633 (N_15633,N_15598,N_12781);
xor U15634 (N_15634,N_12819,N_12913);
or U15635 (N_15635,N_13988,N_14050);
xnor U15636 (N_15636,N_13220,N_12957);
xnor U15637 (N_15637,N_14244,N_14145);
nor U15638 (N_15638,N_14208,N_14641);
nor U15639 (N_15639,N_12674,N_12772);
xor U15640 (N_15640,N_13584,N_15241);
xnor U15641 (N_15641,N_12841,N_14399);
nor U15642 (N_15642,N_13980,N_13172);
nor U15643 (N_15643,N_13117,N_14092);
or U15644 (N_15644,N_12746,N_14382);
xnor U15645 (N_15645,N_13302,N_12889);
or U15646 (N_15646,N_15574,N_15193);
nand U15647 (N_15647,N_15151,N_13150);
and U15648 (N_15648,N_15364,N_13203);
xor U15649 (N_15649,N_14448,N_14316);
or U15650 (N_15650,N_13457,N_14275);
or U15651 (N_15651,N_14983,N_14934);
nand U15652 (N_15652,N_14957,N_13273);
xor U15653 (N_15653,N_15592,N_14489);
nor U15654 (N_15654,N_14917,N_13127);
and U15655 (N_15655,N_14384,N_13412);
xor U15656 (N_15656,N_15404,N_14789);
xor U15657 (N_15657,N_14090,N_12939);
or U15658 (N_15658,N_15290,N_14870);
nand U15659 (N_15659,N_15557,N_15552);
nor U15660 (N_15660,N_14053,N_15559);
nand U15661 (N_15661,N_14783,N_13914);
nand U15662 (N_15662,N_13888,N_12550);
or U15663 (N_15663,N_14644,N_13789);
nor U15664 (N_15664,N_15329,N_15608);
or U15665 (N_15665,N_15184,N_14374);
and U15666 (N_15666,N_14181,N_13240);
and U15667 (N_15667,N_13824,N_13766);
or U15668 (N_15668,N_14681,N_12582);
xor U15669 (N_15669,N_15345,N_13553);
and U15670 (N_15670,N_15380,N_15340);
xor U15671 (N_15671,N_15415,N_12816);
xnor U15672 (N_15672,N_12820,N_14598);
and U15673 (N_15673,N_14351,N_15162);
nor U15674 (N_15674,N_12593,N_13627);
nor U15675 (N_15675,N_13405,N_13122);
nand U15676 (N_15676,N_14682,N_13937);
nand U15677 (N_15677,N_13379,N_13053);
nor U15678 (N_15678,N_12766,N_12884);
xnor U15679 (N_15679,N_13617,N_13139);
xor U15680 (N_15680,N_13008,N_13913);
nor U15681 (N_15681,N_15000,N_15225);
nor U15682 (N_15682,N_13471,N_12580);
and U15683 (N_15683,N_15150,N_13803);
or U15684 (N_15684,N_14835,N_12543);
nor U15685 (N_15685,N_12743,N_15408);
xor U15686 (N_15686,N_12633,N_13875);
nor U15687 (N_15687,N_15560,N_14920);
or U15688 (N_15688,N_14167,N_13161);
or U15689 (N_15689,N_13934,N_13852);
or U15690 (N_15690,N_13029,N_14788);
xor U15691 (N_15691,N_14478,N_14293);
xor U15692 (N_15692,N_15202,N_13443);
and U15693 (N_15693,N_13063,N_12909);
nor U15694 (N_15694,N_12976,N_14534);
nand U15695 (N_15695,N_14172,N_14565);
nor U15696 (N_15696,N_13536,N_15412);
xnor U15697 (N_15697,N_13434,N_12783);
and U15698 (N_15698,N_13187,N_13071);
nor U15699 (N_15699,N_12669,N_13258);
or U15700 (N_15700,N_15188,N_14025);
nand U15701 (N_15701,N_15034,N_13164);
xor U15702 (N_15702,N_13941,N_12584);
nand U15703 (N_15703,N_13271,N_13398);
nor U15704 (N_15704,N_15305,N_14232);
nand U15705 (N_15705,N_15291,N_14891);
or U15706 (N_15706,N_14257,N_13812);
nand U15707 (N_15707,N_12645,N_14561);
nand U15708 (N_15708,N_13085,N_13087);
nor U15709 (N_15709,N_13566,N_13606);
and U15710 (N_15710,N_13202,N_12638);
and U15711 (N_15711,N_14299,N_12993);
nor U15712 (N_15712,N_13928,N_14386);
or U15713 (N_15713,N_13147,N_13310);
nor U15714 (N_15714,N_14120,N_12951);
and U15715 (N_15715,N_14436,N_15013);
xor U15716 (N_15716,N_14919,N_14308);
or U15717 (N_15717,N_14717,N_13520);
nand U15718 (N_15718,N_15471,N_15508);
nand U15719 (N_15719,N_13808,N_14798);
nor U15720 (N_15720,N_13064,N_14005);
nand U15721 (N_15721,N_13685,N_14150);
nor U15722 (N_15722,N_13043,N_12575);
xor U15723 (N_15723,N_12549,N_14266);
or U15724 (N_15724,N_13670,N_12849);
and U15725 (N_15725,N_13309,N_13293);
xor U15726 (N_15726,N_14210,N_14871);
nor U15727 (N_15727,N_13113,N_13815);
xor U15728 (N_15728,N_13603,N_13269);
xnor U15729 (N_15729,N_13681,N_15478);
nor U15730 (N_15730,N_15264,N_14799);
nor U15731 (N_15731,N_14876,N_14056);
xor U15732 (N_15732,N_14014,N_13586);
nor U15733 (N_15733,N_15144,N_15536);
nor U15734 (N_15734,N_13032,N_12874);
nand U15735 (N_15735,N_12637,N_14036);
xnor U15736 (N_15736,N_15256,N_15604);
nor U15737 (N_15737,N_14935,N_14254);
nand U15738 (N_15738,N_13990,N_13585);
nand U15739 (N_15739,N_12878,N_12966);
or U15740 (N_15740,N_15161,N_13495);
or U15741 (N_15741,N_15158,N_12756);
nor U15742 (N_15742,N_14296,N_14412);
or U15743 (N_15743,N_12852,N_13719);
and U15744 (N_15744,N_12552,N_14973);
nor U15745 (N_15745,N_14826,N_13805);
xnor U15746 (N_15746,N_15141,N_13124);
nand U15747 (N_15747,N_13243,N_13059);
or U15748 (N_15748,N_15572,N_12591);
or U15749 (N_15749,N_14462,N_14730);
nor U15750 (N_15750,N_13082,N_14605);
xor U15751 (N_15751,N_15085,N_13193);
xor U15752 (N_15752,N_15336,N_12862);
nand U15753 (N_15753,N_15388,N_12955);
and U15754 (N_15754,N_13645,N_12696);
nor U15755 (N_15755,N_13549,N_12886);
and U15756 (N_15756,N_15439,N_12713);
nand U15757 (N_15757,N_14358,N_15414);
xor U15758 (N_15758,N_14507,N_15545);
or U15759 (N_15759,N_13706,N_14202);
and U15760 (N_15760,N_14365,N_14283);
nor U15761 (N_15761,N_15619,N_15038);
nor U15762 (N_15762,N_13908,N_14062);
xnor U15763 (N_15763,N_14415,N_13890);
nor U15764 (N_15764,N_12982,N_13447);
or U15765 (N_15765,N_13024,N_12985);
nor U15766 (N_15766,N_13788,N_15059);
nand U15767 (N_15767,N_13807,N_15548);
or U15768 (N_15768,N_14907,N_14574);
xor U15769 (N_15769,N_13488,N_13966);
and U15770 (N_15770,N_14485,N_12601);
and U15771 (N_15771,N_15219,N_14575);
and U15772 (N_15772,N_15613,N_14032);
xnor U15773 (N_15773,N_14557,N_13581);
or U15774 (N_15774,N_13497,N_13969);
xnor U15775 (N_15775,N_14470,N_14912);
or U15776 (N_15776,N_13332,N_14200);
nand U15777 (N_15777,N_15288,N_14129);
nor U15778 (N_15778,N_15010,N_14010);
and U15779 (N_15779,N_12901,N_14338);
or U15780 (N_15780,N_13880,N_14770);
nand U15781 (N_15781,N_14228,N_13287);
xnor U15782 (N_15782,N_13748,N_13967);
nand U15783 (N_15783,N_13115,N_13236);
nand U15784 (N_15784,N_13505,N_14968);
or U15785 (N_15785,N_13298,N_13297);
xnor U15786 (N_15786,N_13678,N_13440);
xnor U15787 (N_15787,N_14956,N_13643);
xnor U15788 (N_15788,N_13939,N_13104);
nor U15789 (N_15789,N_15359,N_14527);
and U15790 (N_15790,N_14864,N_15166);
and U15791 (N_15791,N_13348,N_14488);
nand U15792 (N_15792,N_13223,N_14570);
xor U15793 (N_15793,N_13311,N_12734);
nor U15794 (N_15794,N_13061,N_14974);
xor U15795 (N_15795,N_12726,N_13227);
nand U15796 (N_15796,N_13564,N_12665);
nand U15797 (N_15797,N_15179,N_15461);
nand U15798 (N_15798,N_13316,N_14411);
xor U15799 (N_15799,N_15226,N_12969);
or U15800 (N_15800,N_14528,N_13136);
nand U15801 (N_15801,N_15121,N_14556);
nor U15802 (N_15802,N_14940,N_13733);
nor U15803 (N_15803,N_15096,N_14213);
or U15804 (N_15804,N_12546,N_13918);
xnor U15805 (N_15805,N_12578,N_14022);
nor U15806 (N_15806,N_12825,N_15550);
and U15807 (N_15807,N_14427,N_15270);
or U15808 (N_15808,N_13531,N_13351);
and U15809 (N_15809,N_15523,N_14633);
nand U15810 (N_15810,N_14820,N_12809);
and U15811 (N_15811,N_15323,N_14270);
or U15812 (N_15812,N_12754,N_13355);
or U15813 (N_15813,N_15268,N_12972);
and U15814 (N_15814,N_14359,N_13668);
xnor U15815 (N_15815,N_13720,N_15172);
or U15816 (N_15816,N_14674,N_12691);
nor U15817 (N_15817,N_15204,N_14397);
or U15818 (N_15818,N_14139,N_12505);
nand U15819 (N_15819,N_12844,N_15272);
and U15820 (N_15820,N_15133,N_15434);
or U15821 (N_15821,N_13475,N_12716);
or U15822 (N_15822,N_15110,N_13660);
nand U15823 (N_15823,N_15377,N_14334);
nand U15824 (N_15824,N_12917,N_15198);
and U15825 (N_15825,N_12965,N_12532);
xor U15826 (N_15826,N_13039,N_14006);
nand U15827 (N_15827,N_13837,N_13217);
xnor U15828 (N_15828,N_13589,N_13396);
or U15829 (N_15829,N_13225,N_15147);
nand U15830 (N_15830,N_13674,N_14638);
nand U15831 (N_15831,N_15403,N_14268);
or U15832 (N_15832,N_14389,N_13828);
xnor U15833 (N_15833,N_14900,N_14651);
and U15834 (N_15834,N_13272,N_12646);
and U15835 (N_15835,N_15366,N_14125);
and U15836 (N_15836,N_14965,N_12515);
or U15837 (N_15837,N_14098,N_13796);
nand U15838 (N_15838,N_15200,N_15575);
nor U15839 (N_15839,N_15053,N_14740);
and U15840 (N_15840,N_12717,N_13793);
nand U15841 (N_15841,N_14080,N_15489);
or U15842 (N_15842,N_14807,N_15314);
or U15843 (N_15843,N_15107,N_13199);
and U15844 (N_15844,N_12830,N_14696);
and U15845 (N_15845,N_14615,N_13794);
and U15846 (N_15846,N_14848,N_13952);
and U15847 (N_15847,N_13492,N_14828);
or U15848 (N_15848,N_15534,N_14064);
and U15849 (N_15849,N_14801,N_13327);
and U15850 (N_15850,N_12540,N_12837);
nor U15851 (N_15851,N_13708,N_14055);
xnor U15852 (N_15852,N_13333,N_12512);
or U15853 (N_15853,N_15452,N_15588);
xor U15854 (N_15854,N_13346,N_13829);
nor U15855 (N_15855,N_12833,N_12980);
or U15856 (N_15856,N_13732,N_13106);
or U15857 (N_15857,N_13261,N_12857);
nand U15858 (N_15858,N_15087,N_14253);
xor U15859 (N_15859,N_14596,N_14174);
or U15860 (N_15860,N_13703,N_15116);
xnor U15861 (N_15861,N_14714,N_13864);
nand U15862 (N_15862,N_13757,N_12782);
nand U15863 (N_15863,N_14853,N_15001);
or U15864 (N_15864,N_15082,N_14960);
xnor U15865 (N_15865,N_12875,N_14039);
xor U15866 (N_15866,N_15379,N_14041);
nor U15867 (N_15867,N_13700,N_13178);
and U15868 (N_15868,N_15396,N_15501);
nand U15869 (N_15869,N_15111,N_12992);
nand U15870 (N_15870,N_13179,N_14033);
xnor U15871 (N_15871,N_14972,N_13120);
and U15872 (N_15872,N_12608,N_14921);
nor U15873 (N_15873,N_13361,N_14654);
nand U15874 (N_15874,N_13347,N_14518);
and U15875 (N_15875,N_12732,N_15218);
or U15876 (N_15876,N_15227,N_14392);
nor U15877 (N_15877,N_14444,N_15386);
and U15878 (N_15878,N_15436,N_13037);
and U15879 (N_15879,N_14993,N_13883);
nand U15880 (N_15880,N_14969,N_13233);
and U15881 (N_15881,N_13519,N_13743);
nand U15882 (N_15882,N_14417,N_13411);
xor U15883 (N_15883,N_14931,N_15612);
or U15884 (N_15884,N_15330,N_14990);
or U15885 (N_15885,N_13483,N_15553);
nand U15886 (N_15886,N_15401,N_14474);
nor U15887 (N_15887,N_14052,N_14221);
and U15888 (N_15888,N_14406,N_13782);
or U15889 (N_15889,N_14198,N_13647);
or U15890 (N_15890,N_15282,N_14065);
xnor U15891 (N_15891,N_12740,N_14685);
xnor U15892 (N_15892,N_14906,N_13409);
or U15893 (N_15893,N_13098,N_14604);
nand U15894 (N_15894,N_14043,N_14298);
or U15895 (N_15895,N_14736,N_15235);
and U15896 (N_15896,N_14842,N_12818);
or U15897 (N_15897,N_15357,N_12664);
and U15898 (N_15898,N_15618,N_13975);
xnor U15899 (N_15899,N_14400,N_13209);
nor U15900 (N_15900,N_13978,N_13641);
or U15901 (N_15901,N_15104,N_12850);
or U15902 (N_15902,N_15230,N_12708);
nand U15903 (N_15903,N_15544,N_13527);
nand U15904 (N_15904,N_15091,N_14277);
and U15905 (N_15905,N_13354,N_13274);
xnor U15906 (N_15906,N_15022,N_14622);
nand U15907 (N_15907,N_13983,N_13188);
nor U15908 (N_15908,N_14958,N_13876);
xor U15909 (N_15909,N_12660,N_14949);
or U15910 (N_15910,N_14677,N_14819);
nand U15911 (N_15911,N_13126,N_13016);
nor U15912 (N_15912,N_14816,N_12882);
and U15913 (N_15913,N_14635,N_14230);
nand U15914 (N_15914,N_12654,N_15189);
and U15915 (N_15915,N_14152,N_13431);
nand U15916 (N_15916,N_13872,N_15466);
xor U15917 (N_15917,N_14385,N_14754);
or U15918 (N_15918,N_14755,N_13715);
and U15919 (N_15919,N_13238,N_13762);
or U15920 (N_15920,N_13445,N_15344);
and U15921 (N_15921,N_14047,N_14021);
or U15922 (N_15922,N_13366,N_14926);
or U15923 (N_15923,N_15020,N_13021);
and U15924 (N_15924,N_14121,N_13932);
nand U15925 (N_15925,N_13149,N_15190);
and U15926 (N_15926,N_12667,N_13624);
or U15927 (N_15927,N_15595,N_13561);
nand U15928 (N_15928,N_15318,N_12784);
xnor U15929 (N_15929,N_14349,N_14376);
nand U15930 (N_15930,N_13056,N_13415);
xor U15931 (N_15931,N_13449,N_15546);
xor U15932 (N_15932,N_14555,N_14961);
xor U15933 (N_15933,N_12534,N_14187);
nand U15934 (N_15934,N_13823,N_15395);
nor U15935 (N_15935,N_13349,N_13341);
nor U15936 (N_15936,N_15528,N_14581);
and U15937 (N_15937,N_12791,N_14476);
and U15938 (N_15938,N_14953,N_14054);
or U15939 (N_15939,N_12661,N_14519);
nand U15940 (N_15940,N_13173,N_14107);
nor U15941 (N_15941,N_14550,N_12996);
or U15942 (N_15942,N_13785,N_13245);
xor U15943 (N_15943,N_14642,N_13128);
nand U15944 (N_15944,N_14414,N_12885);
or U15945 (N_15945,N_15012,N_15551);
xor U15946 (N_15946,N_15129,N_14149);
xnor U15947 (N_15947,N_14106,N_13752);
or U15948 (N_15948,N_13114,N_14220);
nor U15949 (N_15949,N_15497,N_13335);
nor U15950 (N_15950,N_15126,N_14171);
and U15951 (N_15951,N_15043,N_12883);
nor U15952 (N_15952,N_12806,N_13222);
and U15953 (N_15953,N_14765,N_12958);
xor U15954 (N_15954,N_14498,N_12503);
or U15955 (N_15955,N_14166,N_12610);
and U15956 (N_15956,N_14216,N_15083);
and U15957 (N_15957,N_12651,N_13548);
or U15958 (N_15958,N_15515,N_15361);
nor U15959 (N_15959,N_14303,N_15297);
and U15960 (N_15960,N_12617,N_12721);
nor U15961 (N_15961,N_14834,N_15222);
or U15962 (N_15962,N_12614,N_13138);
nor U15963 (N_15963,N_14304,N_15600);
nor U15964 (N_15964,N_14599,N_14772);
nor U15965 (N_15965,N_14795,N_15265);
xor U15966 (N_15966,N_12652,N_13731);
and U15967 (N_15967,N_13848,N_13781);
xnor U15968 (N_15968,N_12828,N_15153);
nand U15969 (N_15969,N_13590,N_12856);
or U15970 (N_15970,N_12827,N_14089);
and U15971 (N_15971,N_12625,N_15071);
xor U15972 (N_15972,N_13598,N_14209);
xor U15973 (N_15973,N_14509,N_14159);
and U15974 (N_15974,N_15581,N_14840);
nand U15975 (N_15975,N_13102,N_13911);
nand U15976 (N_15976,N_15496,N_14048);
nor U15977 (N_15977,N_15458,N_13419);
nand U15978 (N_15978,N_12673,N_15527);
nor U15979 (N_15979,N_14472,N_14839);
or U15980 (N_15980,N_15483,N_15286);
and U15981 (N_15981,N_12763,N_12587);
or U15982 (N_15982,N_12574,N_12879);
nor U15983 (N_15983,N_13458,N_13288);
xor U15984 (N_15984,N_14204,N_13529);
or U15985 (N_15985,N_13462,N_15518);
xnor U15986 (N_15986,N_12897,N_13565);
and U15987 (N_15987,N_15125,N_13231);
or U15988 (N_15988,N_15036,N_14463);
xnor U15989 (N_15989,N_14544,N_14971);
and U15990 (N_15990,N_13498,N_13323);
nand U15991 (N_15991,N_14231,N_14746);
nand U15992 (N_15992,N_12869,N_14002);
xnor U15993 (N_15993,N_15376,N_13365);
and U15994 (N_15994,N_15351,N_12688);
nand U15995 (N_15995,N_13726,N_14154);
nor U15996 (N_15996,N_13105,N_14767);
xor U15997 (N_15997,N_12589,N_13551);
nor U15998 (N_15998,N_13739,N_15040);
or U15999 (N_15999,N_14591,N_12694);
xnor U16000 (N_16000,N_15054,N_14889);
and U16001 (N_16001,N_14643,N_13058);
and U16002 (N_16002,N_14939,N_13357);
or U16003 (N_16003,N_14542,N_13997);
and U16004 (N_16004,N_13779,N_12923);
nor U16005 (N_16005,N_13418,N_12924);
xnor U16006 (N_16006,N_14784,N_15558);
nor U16007 (N_16007,N_13858,N_12592);
xor U16008 (N_16008,N_13866,N_15444);
xnor U16009 (N_16009,N_14260,N_14409);
or U16010 (N_16010,N_12769,N_12835);
nand U16011 (N_16011,N_15387,N_13067);
nand U16012 (N_16012,N_13454,N_14571);
nor U16013 (N_16013,N_15577,N_13235);
nor U16014 (N_16014,N_14922,N_15185);
nor U16015 (N_16015,N_13577,N_14726);
nand U16016 (N_16016,N_13218,N_13508);
and U16017 (N_16017,N_14758,N_12785);
xor U16018 (N_16018,N_13898,N_12518);
nor U16019 (N_16019,N_14070,N_13212);
nand U16020 (N_16020,N_13407,N_13249);
or U16021 (N_16021,N_14930,N_12704);
nand U16022 (N_16022,N_14199,N_15615);
xnor U16023 (N_16023,N_15405,N_13512);
and U16024 (N_16024,N_14739,N_13765);
and U16025 (N_16025,N_12615,N_12804);
and U16026 (N_16026,N_14806,N_12586);
xor U16027 (N_16027,N_14699,N_15167);
or U16028 (N_16028,N_13522,N_13854);
or U16029 (N_16029,N_13514,N_13007);
nand U16030 (N_16030,N_12762,N_13070);
or U16031 (N_16031,N_15494,N_13004);
nand U16032 (N_16032,N_13219,N_14743);
or U16033 (N_16033,N_13230,N_13044);
xnor U16034 (N_16034,N_12706,N_13110);
nor U16035 (N_16035,N_13046,N_13118);
or U16036 (N_16036,N_13987,N_15187);
nor U16037 (N_16037,N_13065,N_13950);
nor U16038 (N_16038,N_13033,N_12686);
nand U16039 (N_16039,N_13460,N_13501);
nor U16040 (N_16040,N_13697,N_14501);
and U16041 (N_16041,N_14863,N_15035);
or U16042 (N_16042,N_14994,N_13568);
xnor U16043 (N_16043,N_14196,N_12771);
nor U16044 (N_16044,N_14814,N_14461);
nand U16045 (N_16045,N_14028,N_12697);
and U16046 (N_16046,N_15004,N_14256);
or U16047 (N_16047,N_14989,N_14318);
or U16048 (N_16048,N_14311,N_13496);
xor U16049 (N_16049,N_15263,N_14071);
or U16050 (N_16050,N_13060,N_14796);
or U16051 (N_16051,N_13600,N_12832);
or U16052 (N_16052,N_12650,N_13638);
or U16053 (N_16053,N_14324,N_12753);
or U16054 (N_16054,N_14426,N_14103);
xnor U16055 (N_16055,N_13239,N_14526);
and U16056 (N_16056,N_14272,N_14193);
nor U16057 (N_16057,N_13844,N_14331);
and U16058 (N_16058,N_14782,N_12722);
nand U16059 (N_16059,N_14988,N_14011);
nor U16060 (N_16060,N_15052,N_14105);
or U16061 (N_16061,N_14388,N_13439);
nand U16062 (N_16062,N_14441,N_14431);
xnor U16063 (N_16063,N_14804,N_14587);
xnor U16064 (N_16064,N_14815,N_13337);
nand U16065 (N_16065,N_14785,N_12662);
nand U16066 (N_16066,N_15302,N_12947);
xor U16067 (N_16067,N_13751,N_13784);
nor U16068 (N_16068,N_14217,N_12876);
xnor U16069 (N_16069,N_12903,N_12779);
nand U16070 (N_16070,N_12551,N_15074);
nand U16071 (N_16071,N_13096,N_14639);
nor U16072 (N_16072,N_12817,N_14741);
xnor U16073 (N_16073,N_13763,N_14369);
and U16074 (N_16074,N_14661,N_15491);
and U16075 (N_16075,N_12572,N_15139);
nor U16076 (N_16076,N_13250,N_13840);
xor U16077 (N_16077,N_15365,N_13092);
xnor U16078 (N_16078,N_14950,N_14363);
and U16079 (N_16079,N_14793,N_13491);
nand U16080 (N_16080,N_12866,N_15164);
nand U16081 (N_16081,N_13414,N_14811);
or U16082 (N_16082,N_15122,N_15622);
and U16083 (N_16083,N_12870,N_13943);
or U16084 (N_16084,N_13560,N_12789);
and U16085 (N_16085,N_12964,N_13929);
and U16086 (N_16086,N_14590,N_14745);
nor U16087 (N_16087,N_14069,N_12873);
xnor U16088 (N_16088,N_15578,N_15488);
and U16089 (N_16089,N_13904,N_15367);
and U16090 (N_16090,N_12954,N_12807);
or U16091 (N_16091,N_13022,N_14947);
and U16092 (N_16092,N_15547,N_15243);
or U16093 (N_16093,N_13672,N_13874);
or U16094 (N_16094,N_15056,N_15430);
and U16095 (N_16095,N_13015,N_15018);
and U16096 (N_16096,N_15465,N_15350);
nor U16097 (N_16097,N_13390,N_14264);
and U16098 (N_16098,N_14332,N_13655);
nand U16099 (N_16099,N_14175,N_15254);
nor U16100 (N_16100,N_15078,N_14951);
nand U16101 (N_16101,N_13175,N_14295);
nand U16102 (N_16102,N_12907,N_13477);
and U16103 (N_16103,N_15542,N_13839);
or U16104 (N_16104,N_15363,N_14704);
and U16105 (N_16105,N_12542,N_14394);
and U16106 (N_16106,N_14097,N_12727);
or U16107 (N_16107,N_13755,N_13702);
xnor U16108 (N_16108,N_12703,N_14093);
xor U16109 (N_16109,N_13576,N_14733);
and U16110 (N_16110,N_12800,N_14883);
nor U16111 (N_16111,N_13049,N_13228);
or U16112 (N_16112,N_12757,N_14073);
and U16113 (N_16113,N_13413,N_14827);
nor U16114 (N_16114,N_15163,N_14396);
xor U16115 (N_16115,N_14419,N_13027);
or U16116 (N_16116,N_12863,N_14822);
nor U16117 (N_16117,N_14243,N_13772);
and U16118 (N_16118,N_15220,N_13040);
xnor U16119 (N_16119,N_13017,N_13306);
nand U16120 (N_16120,N_13718,N_13406);
xnor U16121 (N_16121,N_14724,N_13183);
or U16122 (N_16122,N_14905,N_13399);
nand U16123 (N_16123,N_14373,N_15063);
xnor U16124 (N_16124,N_13077,N_14780);
and U16125 (N_16125,N_12933,N_14475);
or U16126 (N_16126,N_13867,N_14286);
and U16127 (N_16127,N_12995,N_15457);
nand U16128 (N_16128,N_14282,N_15611);
and U16129 (N_16129,N_15234,N_13207);
xnor U16130 (N_16130,N_14333,N_14235);
and U16131 (N_16131,N_15602,N_14705);
nand U16132 (N_16132,N_13761,N_13712);
or U16133 (N_16133,N_15090,N_14143);
xor U16134 (N_16134,N_14323,N_15373);
xnor U16135 (N_16135,N_14670,N_13283);
or U16136 (N_16136,N_13651,N_14218);
nor U16137 (N_16137,N_13195,N_13370);
nor U16138 (N_16138,N_14517,N_13869);
nand U16139 (N_16139,N_15585,N_13628);
xnor U16140 (N_16140,N_14424,N_14594);
xnor U16141 (N_16141,N_14178,N_15191);
xor U16142 (N_16142,N_14138,N_13701);
xnor U16143 (N_16143,N_13896,N_13307);
xor U16144 (N_16144,N_13927,N_15448);
nor U16145 (N_16145,N_12690,N_14503);
and U16146 (N_16146,N_13038,N_13842);
nand U16147 (N_16147,N_12724,N_15248);
and U16148 (N_16148,N_15428,N_14500);
nand U16149 (N_16149,N_12655,N_13466);
or U16150 (N_16150,N_12595,N_13444);
and U16151 (N_16151,N_14013,N_14868);
xnor U16152 (N_16152,N_13953,N_14948);
xor U16153 (N_16153,N_14636,N_15420);
nor U16154 (N_16154,N_15512,N_13076);
nor U16155 (N_16155,N_15482,N_12764);
or U16156 (N_16156,N_13006,N_13003);
or U16157 (N_16157,N_13856,N_14802);
nand U16158 (N_16158,N_13125,N_15058);
nor U16159 (N_16159,N_13464,N_13539);
nor U16160 (N_16160,N_15348,N_15309);
or U16161 (N_16161,N_13516,N_13107);
or U16162 (N_16162,N_13902,N_13292);
xor U16163 (N_16163,N_14727,N_14928);
and U16164 (N_16164,N_13338,N_12758);
nand U16165 (N_16165,N_15473,N_14072);
nor U16166 (N_16166,N_15524,N_15442);
and U16167 (N_16167,N_14214,N_12702);
nor U16168 (N_16168,N_13642,N_14663);
nor U16169 (N_16169,N_13131,N_14975);
xnor U16170 (N_16170,N_14104,N_13919);
and U16171 (N_16171,N_13968,N_14482);
nand U16172 (N_16172,N_15207,N_14297);
and U16173 (N_16173,N_15047,N_13916);
nor U16174 (N_16174,N_14625,N_15539);
nor U16175 (N_16175,N_13817,N_14998);
or U16176 (N_16176,N_14878,N_13393);
xor U16177 (N_16177,N_13695,N_13894);
nor U16178 (N_16178,N_13242,N_15382);
nand U16179 (N_16179,N_14759,N_15561);
xor U16180 (N_16180,N_15565,N_15335);
nor U16181 (N_16181,N_14469,N_13737);
nand U16182 (N_16182,N_14446,N_12877);
xnor U16183 (N_16183,N_15413,N_15487);
nor U16184 (N_16184,N_14177,N_14671);
xor U16185 (N_16185,N_14247,N_13374);
or U16186 (N_16186,N_14569,N_14936);
xor U16187 (N_16187,N_15540,N_13688);
nor U16188 (N_16188,N_13859,N_14514);
nand U16189 (N_16189,N_14601,N_12500);
or U16190 (N_16190,N_13025,N_13132);
and U16191 (N_16191,N_14567,N_13797);
nor U16192 (N_16192,N_15231,N_12935);
or U16193 (N_16193,N_15095,N_13388);
nor U16194 (N_16194,N_13009,N_13582);
xnor U16195 (N_16195,N_13353,N_12525);
nand U16196 (N_16196,N_14716,N_14466);
nor U16197 (N_16197,N_13760,N_15411);
nor U16198 (N_16198,N_13621,N_15432);
or U16199 (N_16199,N_12731,N_14020);
nand U16200 (N_16200,N_14455,N_14309);
nand U16201 (N_16201,N_13378,N_14416);
nor U16202 (N_16202,N_15008,N_12916);
nor U16203 (N_16203,N_12906,N_12730);
and U16204 (N_16204,N_12684,N_14504);
nor U16205 (N_16205,N_13314,N_14668);
nand U16206 (N_16206,N_13591,N_12530);
nor U16207 (N_16207,N_13698,N_13819);
xnor U16208 (N_16208,N_13141,N_12968);
xnor U16209 (N_16209,N_13055,N_14538);
nor U16210 (N_16210,N_14449,N_13494);
or U16211 (N_16211,N_14867,N_15407);
xnor U16212 (N_16212,N_13528,N_15113);
xor U16213 (N_16213,N_13442,N_13570);
nor U16214 (N_16214,N_13486,N_15568);
and U16215 (N_16215,N_13480,N_14096);
nor U16216 (N_16216,N_13515,N_13171);
xnor U16217 (N_16217,N_15319,N_14572);
and U16218 (N_16218,N_12774,N_13773);
and U16219 (N_16219,N_15276,N_13632);
and U16220 (N_16220,N_13253,N_14234);
nor U16221 (N_16221,N_14875,N_12607);
or U16222 (N_16222,N_13707,N_13870);
nand U16223 (N_16223,N_14471,N_14088);
nand U16224 (N_16224,N_15349,N_14817);
and U16225 (N_16225,N_15050,N_13689);
nand U16226 (N_16226,N_14265,N_15045);
nand U16227 (N_16227,N_13144,N_15315);
nor U16228 (N_16228,N_13506,N_14288);
nand U16229 (N_16229,N_14831,N_15358);
and U16230 (N_16230,N_13671,N_13942);
xnor U16231 (N_16231,N_15569,N_13892);
nand U16232 (N_16232,N_14543,N_13567);
xor U16233 (N_16233,N_15168,N_15601);
nand U16234 (N_16234,N_15513,N_14608);
or U16235 (N_16235,N_13380,N_14460);
and U16236 (N_16236,N_14458,N_15521);
nor U16237 (N_16237,N_13665,N_14843);
xnor U16238 (N_16238,N_13336,N_14148);
xor U16239 (N_16239,N_12643,N_15617);
xnor U16240 (N_16240,N_13500,N_14856);
nand U16241 (N_16241,N_14037,N_13899);
xor U16242 (N_16242,N_14980,N_13383);
or U16243 (N_16243,N_13103,N_14678);
nor U16244 (N_16244,N_12921,N_13917);
nor U16245 (N_16245,N_14327,N_15587);
nand U16246 (N_16246,N_14340,N_15031);
and U16247 (N_16247,N_15427,N_14656);
nor U16248 (N_16248,N_15398,N_14742);
xnor U16249 (N_16249,N_14545,N_13244);
nor U16250 (N_16250,N_14764,N_13675);
xnor U16251 (N_16251,N_13683,N_15332);
nand U16252 (N_16252,N_12956,N_13206);
xnor U16253 (N_16253,N_14335,N_13791);
or U16254 (N_16254,N_12705,N_13639);
nor U16255 (N_16255,N_13543,N_15175);
nand U16256 (N_16256,N_13066,N_14486);
and U16257 (N_16257,N_15148,N_14580);
nor U16258 (N_16258,N_14464,N_12760);
or U16259 (N_16259,N_13503,N_13583);
or U16260 (N_16260,N_14068,N_15252);
and U16261 (N_16261,N_15099,N_14533);
xor U16262 (N_16262,N_14042,N_15307);
or U16263 (N_16263,N_13165,N_15292);
or U16264 (N_16264,N_13981,N_14946);
xor U16265 (N_16265,N_14621,N_13910);
nor U16266 (N_16266,N_13573,N_14403);
or U16267 (N_16267,N_14276,N_13650);
xnor U16268 (N_16268,N_15537,N_14893);
nor U16269 (N_16269,N_14468,N_13112);
and U16270 (N_16270,N_12629,N_12538);
nor U16271 (N_16271,N_13540,N_13404);
xnor U16272 (N_16272,N_13931,N_12915);
nand U16273 (N_16273,N_13221,N_14954);
or U16274 (N_16274,N_13831,N_14045);
and U16275 (N_16275,N_15062,N_14380);
and U16276 (N_16276,N_13857,N_13481);
or U16277 (N_16277,N_12516,N_13502);
and U16278 (N_16278,N_15069,N_14865);
nor U16279 (N_16279,N_15257,N_14360);
nor U16280 (N_16280,N_12620,N_14620);
or U16281 (N_16281,N_14046,N_13163);
nor U16282 (N_16282,N_13210,N_13108);
nor U16283 (N_16283,N_13140,N_15603);
or U16284 (N_16284,N_14857,N_13391);
xnor U16285 (N_16285,N_14982,N_15203);
and U16286 (N_16286,N_13991,N_15287);
nand U16287 (N_16287,N_12677,N_12573);
xnor U16288 (N_16288,N_13266,N_14718);
or U16289 (N_16289,N_15325,N_13091);
nand U16290 (N_16290,N_14630,N_14916);
and U16291 (N_16291,N_13759,N_15507);
nor U16292 (N_16292,N_14964,N_14886);
and U16293 (N_16293,N_13710,N_14432);
or U16294 (N_16294,N_14035,N_13270);
nor U16295 (N_16295,N_13705,N_14892);
nor U16296 (N_16296,N_13634,N_15209);
and U16297 (N_16297,N_13455,N_13186);
or U16298 (N_16298,N_12997,N_13473);
and U16299 (N_16299,N_14997,N_14186);
nand U16300 (N_16300,N_13693,N_13135);
nor U16301 (N_16301,N_13397,N_14086);
or U16302 (N_16302,N_13277,N_15154);
xor U16303 (N_16303,N_15130,N_14094);
xor U16304 (N_16304,N_13385,N_14112);
nand U16305 (N_16305,N_14371,N_12952);
and U16306 (N_16306,N_13426,N_13525);
xnor U16307 (N_16307,N_14079,N_14945);
nand U16308 (N_16308,N_14430,N_13542);
xor U16309 (N_16309,N_14616,N_15423);
nor U16310 (N_16310,N_13746,N_14236);
and U16311 (N_16311,N_12914,N_14081);
or U16312 (N_16312,N_15493,N_15048);
or U16313 (N_16313,N_13736,N_14923);
or U16314 (N_16314,N_12949,N_13605);
nand U16315 (N_16315,N_15266,N_15317);
nor U16316 (N_16316,N_12678,N_15033);
nand U16317 (N_16317,N_15081,N_13019);
nor U16318 (N_16318,N_13538,N_12910);
nor U16319 (N_16319,N_15098,N_14858);
nor U16320 (N_16320,N_13086,N_15137);
xor U16321 (N_16321,N_12642,N_12749);
and U16322 (N_16322,N_12896,N_12846);
nor U16323 (N_16323,N_15495,N_14422);
nand U16324 (N_16324,N_13813,N_12569);
nand U16325 (N_16325,N_15385,N_14879);
nand U16326 (N_16326,N_13400,N_14566);
and U16327 (N_16327,N_12600,N_15418);
or U16328 (N_16328,N_13686,N_14184);
or U16329 (N_16329,N_13547,N_14645);
xor U16330 (N_16330,N_12568,N_12928);
or U16331 (N_16331,N_14012,N_12682);
or U16332 (N_16332,N_14813,N_14810);
nor U16333 (N_16333,N_13579,N_13073);
nand U16334 (N_16334,N_12855,N_13838);
and U16335 (N_16335,N_13521,N_15057);
and U16336 (N_16336,N_14573,N_14933);
nand U16337 (N_16337,N_14752,N_14191);
nand U16338 (N_16338,N_13893,N_14881);
nand U16339 (N_16339,N_13571,N_13229);
xor U16340 (N_16340,N_13123,N_15599);
xnor U16341 (N_16341,N_14161,N_13878);
and U16342 (N_16342,N_13801,N_15118);
nor U16343 (N_16343,N_15419,N_13429);
nand U16344 (N_16344,N_12974,N_14326);
nand U16345 (N_16345,N_13232,N_13441);
nor U16346 (N_16346,N_13602,N_13159);
or U16347 (N_16347,N_14134,N_15455);
xor U16348 (N_16348,N_12892,N_12506);
or U16349 (N_16349,N_15579,N_14562);
and U16350 (N_16350,N_14866,N_13814);
nand U16351 (N_16351,N_13930,N_13679);
and U16352 (N_16352,N_13699,N_12987);
and U16353 (N_16353,N_12728,N_14761);
nor U16354 (N_16354,N_13510,N_14589);
nor U16355 (N_16355,N_15289,N_15273);
nor U16356 (N_16356,N_13532,N_13289);
and U16357 (N_16357,N_14451,N_14083);
nor U16358 (N_16358,N_14738,N_14233);
nand U16359 (N_16359,N_15221,N_14611);
or U16360 (N_16360,N_13588,N_15308);
nor U16361 (N_16361,N_13608,N_14890);
xor U16362 (N_16362,N_14675,N_15333);
nand U16363 (N_16363,N_14262,N_14578);
xnor U16364 (N_16364,N_15354,N_15088);
xnor U16365 (N_16365,N_13636,N_14437);
nor U16366 (N_16366,N_13369,N_13559);
xor U16367 (N_16367,N_12831,N_14657);
and U16368 (N_16368,N_14666,N_14381);
nor U16369 (N_16369,N_15470,N_15326);
nor U16370 (N_16370,N_14680,N_12959);
nand U16371 (N_16371,N_14132,N_13321);
nor U16372 (N_16372,N_13903,N_13537);
nand U16373 (N_16373,N_12978,N_13224);
nor U16374 (N_16374,N_15169,N_14165);
xnor U16375 (N_16375,N_13775,N_14952);
xor U16376 (N_16376,N_12566,N_12900);
nand U16377 (N_16377,N_15609,N_15417);
or U16378 (N_16378,N_13769,N_15073);
and U16379 (N_16379,N_14882,N_14885);
xor U16380 (N_16380,N_13050,N_15334);
and U16381 (N_16381,N_12765,N_14769);
xor U16382 (N_16382,N_14439,N_13900);
nor U16383 (N_16383,N_14407,N_12687);
and U16384 (N_16384,N_15502,N_14812);
xnor U16385 (N_16385,N_15119,N_15589);
or U16386 (N_16386,N_15065,N_14558);
xnor U16387 (N_16387,N_14368,N_13035);
or U16388 (N_16388,N_13234,N_15094);
nor U16389 (N_16389,N_12858,N_13633);
and U16390 (N_16390,N_14263,N_15114);
xor U16391 (N_16391,N_13986,N_14391);
nor U16392 (N_16392,N_13133,N_14689);
xnor U16393 (N_16393,N_14300,N_14941);
nand U16394 (N_16394,N_15206,N_15459);
or U16395 (N_16395,N_15352,N_13897);
and U16396 (N_16396,N_14330,N_14887);
or U16397 (N_16397,N_15402,N_15543);
nand U16398 (N_16398,N_14483,N_14756);
nand U16399 (N_16399,N_14000,N_12563);
or U16400 (N_16400,N_13871,N_12770);
or U16401 (N_16401,N_15328,N_15406);
nor U16402 (N_16402,N_12926,N_15409);
or U16403 (N_16403,N_12773,N_14141);
nor U16404 (N_16404,N_12511,N_14911);
nand U16405 (N_16405,N_13214,N_15503);
xnor U16406 (N_16406,N_15597,N_15246);
xnor U16407 (N_16407,N_14693,N_14119);
nor U16408 (N_16408,N_13356,N_12737);
nand U16409 (N_16409,N_13364,N_14118);
xnor U16410 (N_16410,N_13281,N_15519);
xor U16411 (N_16411,N_12994,N_13921);
nor U16412 (N_16412,N_15321,N_15425);
or U16413 (N_16413,N_12936,N_14434);
xnor U16414 (N_16414,N_14009,N_13821);
xnor U16415 (N_16415,N_14249,N_13256);
nor U16416 (N_16416,N_14137,N_13964);
or U16417 (N_16417,N_14751,N_14825);
nand U16418 (N_16418,N_15441,N_14018);
nand U16419 (N_16419,N_13609,N_12979);
and U16420 (N_16420,N_15030,N_13992);
xnor U16421 (N_16421,N_13030,N_12898);
nor U16422 (N_16422,N_12942,N_14102);
or U16423 (N_16423,N_15610,N_15583);
and U16424 (N_16424,N_14341,N_14720);
xnor U16425 (N_16425,N_14653,N_13296);
nor U16426 (N_16426,N_13558,N_12657);
nor U16427 (N_16427,N_15383,N_12509);
nand U16428 (N_16428,N_13569,N_13160);
nand U16429 (N_16429,N_15106,N_14610);
nand U16430 (N_16430,N_14227,N_14168);
nor U16431 (N_16431,N_12887,N_13476);
or U16432 (N_16432,N_13834,N_14708);
or U16433 (N_16433,N_14248,N_13174);
and U16434 (N_16434,N_14786,N_12679);
nand U16435 (N_16435,N_15212,N_15143);
and U16436 (N_16436,N_14583,N_12795);
or U16437 (N_16437,N_15573,N_14366);
xnor U16438 (N_16438,N_13129,N_14190);
or U16439 (N_16439,N_13607,N_14896);
nand U16440 (N_16440,N_13922,N_13728);
and U16441 (N_16441,N_14979,N_13923);
and U16442 (N_16442,N_14305,N_14357);
nand U16443 (N_16443,N_13947,N_13446);
xnor U16444 (N_16444,N_13524,N_14932);
and U16445 (N_16445,N_14729,N_14026);
xor U16446 (N_16446,N_14215,N_15170);
nor U16447 (N_16447,N_14506,N_12829);
xnor U16448 (N_16448,N_14481,N_14748);
xor U16449 (N_16449,N_13469,N_12801);
nor U16450 (N_16450,N_12521,N_15313);
nand U16451 (N_16451,N_13152,N_13973);
and U16452 (N_16452,N_14629,N_13213);
xor U16453 (N_16453,N_14548,N_12931);
or U16454 (N_16454,N_14147,N_13646);
nor U16455 (N_16455,N_12880,N_14924);
nand U16456 (N_16456,N_15177,N_15499);
nand U16457 (N_16457,N_14477,N_15017);
nand U16458 (N_16458,N_14440,N_12745);
nor U16459 (N_16459,N_13436,N_13403);
nor U16460 (N_16460,N_15181,N_14787);
nand U16461 (N_16461,N_13372,N_13552);
nor U16462 (N_16462,N_13767,N_13714);
nand U16463 (N_16463,N_15533,N_14343);
nand U16464 (N_16464,N_12675,N_15027);
nor U16465 (N_16465,N_13940,N_14003);
and U16466 (N_16466,N_14034,N_14410);
or U16467 (N_16467,N_12630,N_12680);
nor U16468 (N_16468,N_14837,N_15269);
nand U16469 (N_16469,N_13935,N_13334);
nor U16470 (N_16470,N_15504,N_12561);
and U16471 (N_16471,N_13504,N_14854);
nand U16472 (N_16472,N_13254,N_15251);
xor U16473 (N_16473,N_13820,N_13677);
nand U16474 (N_16474,N_13861,N_12894);
xnor U16475 (N_16475,N_15467,N_15049);
xnor U16476 (N_16476,N_14404,N_14467);
xor U16477 (N_16477,N_12788,N_13386);
or U16478 (N_16478,N_13345,N_14781);
and U16479 (N_16479,N_14176,N_12624);
xor U16480 (N_16480,N_14836,N_14255);
and U16481 (N_16481,N_13530,N_14797);
xnor U16482 (N_16482,N_12937,N_13395);
or U16483 (N_16483,N_12908,N_13425);
nor U16484 (N_16484,N_15124,N_13158);
nor U16485 (N_16485,N_15347,N_14287);
nand U16486 (N_16486,N_14370,N_13920);
nand U16487 (N_16487,N_13080,N_13295);
nand U16488 (N_16488,N_14450,N_12631);
nor U16489 (N_16489,N_12932,N_14194);
nor U16490 (N_16490,N_14880,N_13786);
or U16491 (N_16491,N_15192,N_14679);
nor U16492 (N_16492,N_14901,N_13612);
xnor U16493 (N_16493,N_15080,N_12938);
or U16494 (N_16494,N_14728,N_13155);
nor U16495 (N_16495,N_15520,N_14719);
xnor U16496 (N_16496,N_15039,N_14133);
xnor U16497 (N_16497,N_13626,N_14279);
nor U16498 (N_16498,N_14809,N_15481);
and U16499 (N_16499,N_15285,N_13578);
or U16500 (N_16500,N_13704,N_12567);
and U16501 (N_16501,N_13319,N_14457);
or U16502 (N_16502,N_12768,N_14694);
nor U16503 (N_16503,N_13358,N_12961);
xnor U16504 (N_16504,N_15372,N_15616);
nand U16505 (N_16505,N_14520,N_14075);
and U16506 (N_16506,N_13955,N_14593);
nand U16507 (N_16507,N_13246,N_15322);
and U16508 (N_16508,N_12984,N_13845);
nor U16509 (N_16509,N_13036,N_14531);
nand U16510 (N_16510,N_14027,N_13204);
nand U16511 (N_16511,N_13996,N_15183);
xnor U16512 (N_16512,N_14015,N_12810);
or U16513 (N_16513,N_12666,N_14938);
xor U16514 (N_16514,N_12948,N_13002);
xor U16515 (N_16515,N_13684,N_12919);
nor U16516 (N_16516,N_13926,N_12871);
nor U16517 (N_16517,N_13084,N_13069);
nor U16518 (N_16518,N_14185,N_14762);
xnor U16519 (N_16519,N_13499,N_14899);
nor U16520 (N_16520,N_13168,N_12776);
and U16521 (N_16521,N_14314,N_13325);
and U16522 (N_16522,N_12805,N_13089);
nor U16523 (N_16523,N_15570,N_15026);
nor U16524 (N_16524,N_14246,N_14805);
xor U16525 (N_16525,N_15055,N_13170);
nand U16526 (N_16526,N_12786,N_12562);
or U16527 (N_16527,N_12531,N_12934);
nor U16528 (N_16528,N_12599,N_13868);
and U16529 (N_16529,N_13339,N_15460);
xnor U16530 (N_16530,N_13318,N_12559);
nand U16531 (N_16531,N_13863,N_12689);
or U16532 (N_16532,N_15009,N_13260);
nor U16533 (N_16533,N_14320,N_14648);
nand U16534 (N_16534,N_12943,N_13180);
xor U16535 (N_16535,N_12735,N_12868);
or U16536 (N_16536,N_13974,N_14091);
and U16537 (N_16537,N_13616,N_15445);
or U16538 (N_16538,N_12510,N_15006);
nand U16539 (N_16539,N_12636,N_14631);
nand U16540 (N_16540,N_14222,N_13263);
nor U16541 (N_16541,N_13556,N_14624);
and U16542 (N_16542,N_13352,N_14051);
and U16543 (N_16543,N_13028,N_14523);
xor U16544 (N_16544,N_15165,N_14030);
xnor U16545 (N_16545,N_15245,N_15279);
and U16546 (N_16546,N_15475,N_13074);
and U16547 (N_16547,N_14219,N_14985);
nor U16548 (N_16548,N_13276,N_14977);
and U16549 (N_16549,N_15197,N_13754);
nor U16550 (N_16550,N_14546,N_14087);
xor U16551 (N_16551,N_14480,N_14659);
or U16552 (N_16552,N_15477,N_13961);
xnor U16553 (N_16553,N_13722,N_12520);
and U16554 (N_16554,N_14592,N_13574);
nand U16555 (N_16555,N_13648,N_13618);
nor U16556 (N_16556,N_12626,N_15232);
nor U16557 (N_16557,N_15075,N_15338);
nand U16558 (N_16558,N_13862,N_14057);
or U16559 (N_16559,N_14984,N_15563);
or U16560 (N_16560,N_15620,N_15029);
nor U16561 (N_16561,N_14339,N_13667);
or U16562 (N_16562,N_12590,N_14113);
and U16563 (N_16563,N_12741,N_14713);
and U16564 (N_16564,N_15281,N_13915);
xor U16565 (N_16565,N_13933,N_14877);
and U16566 (N_16566,N_13177,N_14902);
xor U16567 (N_16567,N_13157,N_14017);
and U16568 (N_16568,N_14847,N_12767);
or U16569 (N_16569,N_14530,N_13938);
nand U16570 (N_16570,N_14838,N_13047);
xnor U16571 (N_16571,N_12672,N_15454);
or U16572 (N_16572,N_14004,N_14226);
xor U16573 (N_16573,N_14554,N_14160);
nor U16574 (N_16574,N_15378,N_14564);
nand U16575 (N_16575,N_14169,N_14888);
and U16576 (N_16576,N_14372,N_13730);
or U16577 (N_16577,N_13134,N_12983);
and U16578 (N_16578,N_13886,N_15021);
xnor U16579 (N_16579,N_15194,N_15356);
xor U16580 (N_16580,N_15182,N_13982);
or U16581 (N_16581,N_14281,N_14860);
and U16582 (N_16582,N_13448,N_12797);
nor U16583 (N_16583,N_13563,N_13610);
nor U16584 (N_16584,N_15624,N_15135);
xnor U16585 (N_16585,N_13830,N_14060);
xnor U16586 (N_16586,N_14937,N_13925);
nor U16587 (N_16587,N_13375,N_12950);
xnor U16588 (N_16588,N_13012,N_13313);
or U16589 (N_16589,N_12891,N_13507);
nor U16590 (N_16590,N_15002,N_15623);
or U16591 (N_16591,N_14179,N_13735);
or U16592 (N_16592,N_13472,N_12523);
xor U16593 (N_16593,N_14603,N_12991);
nor U16594 (N_16594,N_14859,N_15571);
nor U16595 (N_16595,N_14551,N_12588);
xor U16596 (N_16596,N_13535,N_13742);
nor U16597 (N_16597,N_13420,N_14284);
or U16598 (N_16598,N_14085,N_13328);
nor U16599 (N_16599,N_12681,N_15132);
and U16600 (N_16600,N_14925,N_12986);
and U16601 (N_16601,N_12798,N_13484);
xnor U16602 (N_16602,N_13806,N_14547);
nand U16603 (N_16603,N_13185,N_14753);
and U16604 (N_16604,N_14986,N_14101);
nand U16605 (N_16605,N_12613,N_14999);
or U16606 (N_16606,N_15155,N_14433);
nand U16607 (N_16607,N_13985,N_13881);
xnor U16608 (N_16608,N_15261,N_13691);
or U16609 (N_16609,N_14001,N_13865);
nand U16610 (N_16610,N_12583,N_14640);
or U16611 (N_16611,N_13026,N_13640);
nand U16612 (N_16612,N_13604,N_15399);
nand U16613 (N_16613,N_14522,N_12990);
nor U16614 (N_16614,N_13368,N_14348);
nand U16615 (N_16615,N_13020,N_14766);
nand U16616 (N_16616,N_12925,N_12911);
and U16617 (N_16617,N_12612,N_12755);
xnor U16618 (N_16618,N_14768,N_15051);
and U16619 (N_16619,N_15213,N_14662);
and U16620 (N_16620,N_14823,N_13877);
or U16621 (N_16621,N_15301,N_13305);
or U16622 (N_16622,N_13401,N_12902);
nor U16623 (N_16623,N_12714,N_13294);
nand U16624 (N_16624,N_15011,N_15531);
nand U16625 (N_16625,N_15437,N_13509);
xor U16626 (N_16626,N_13557,N_14698);
nor U16627 (N_16627,N_14383,N_12699);
xnor U16628 (N_16628,N_14862,N_12761);
or U16629 (N_16629,N_14894,N_13887);
xnor U16630 (N_16630,N_13976,N_13014);
or U16631 (N_16631,N_12663,N_12859);
nand U16632 (N_16632,N_13944,N_15003);
and U16633 (N_16633,N_12865,N_14818);
or U16634 (N_16634,N_15079,N_15514);
nand U16635 (N_16635,N_13818,N_13197);
nor U16636 (N_16636,N_15267,N_14873);
nand U16637 (N_16637,N_14703,N_14207);
xor U16638 (N_16638,N_12571,N_13465);
xor U16639 (N_16639,N_13018,N_14319);
and U16640 (N_16640,N_15554,N_13855);
or U16641 (N_16641,N_14212,N_13013);
nor U16642 (N_16642,N_15258,N_12659);
nor U16643 (N_16643,N_14127,N_14344);
or U16644 (N_16644,N_12899,N_14016);
and U16645 (N_16645,N_14869,N_13959);
nor U16646 (N_16646,N_15476,N_12683);
nor U16647 (N_16647,N_12658,N_12544);
xor U16648 (N_16648,N_12671,N_12861);
or U16649 (N_16649,N_13279,N_12602);
xor U16650 (N_16650,N_13924,N_13461);
nor U16651 (N_16651,N_13268,N_14395);
nor U16652 (N_16652,N_15025,N_14061);
and U16653 (N_16653,N_14136,N_15157);
nor U16654 (N_16654,N_13611,N_12720);
nor U16655 (N_16655,N_13145,N_15242);
or U16656 (N_16656,N_14211,N_15535);
or U16657 (N_16657,N_14914,N_13526);
nor U16658 (N_16658,N_14535,N_14904);
nand U16659 (N_16659,N_12653,N_15490);
and U16660 (N_16660,N_14800,N_13635);
or U16661 (N_16661,N_12977,N_15456);
and U16662 (N_16662,N_13960,N_13090);
nand U16663 (N_16663,N_12963,N_15300);
and U16664 (N_16664,N_15509,N_13054);
xnor U16665 (N_16665,N_13816,N_15061);
and U16666 (N_16666,N_14627,N_15089);
and U16667 (N_16667,N_13889,N_14280);
or U16668 (N_16668,N_14390,N_12693);
nand U16669 (N_16669,N_12851,N_14872);
xnor U16670 (N_16670,N_13620,N_13387);
xnor U16671 (N_16671,N_15299,N_12790);
or U16672 (N_16672,N_13097,N_14721);
and U16673 (N_16673,N_14473,N_12513);
xnor U16674 (N_16674,N_14240,N_15346);
nor U16675 (N_16675,N_13376,N_12812);
nand U16676 (N_16676,N_13146,N_13005);
and U16677 (N_16677,N_15101,N_15451);
nor U16678 (N_16678,N_13493,N_13042);
nand U16679 (N_16679,N_15066,N_12904);
nand U16680 (N_16680,N_14529,N_14224);
nor U16681 (N_16681,N_13072,N_14379);
xnor U16682 (N_16682,N_13251,N_14524);
xnor U16683 (N_16683,N_13075,N_13694);
nand U16684 (N_16684,N_12777,N_12526);
xor U16685 (N_16685,N_13727,N_13194);
and U16686 (N_16686,N_14494,N_15046);
nand U16687 (N_16687,N_14667,N_13416);
nand U16688 (N_16688,N_14428,N_14245);
and U16689 (N_16689,N_15541,N_13664);
or U16690 (N_16690,N_15271,N_15160);
nor U16691 (N_16691,N_15304,N_15275);
and U16692 (N_16692,N_15117,N_14117);
or U16693 (N_16693,N_13666,N_14123);
nand U16694 (N_16694,N_14122,N_13723);
nand U16695 (N_16695,N_15472,N_14536);
xnor U16696 (N_16696,N_15479,N_15510);
xnor U16697 (N_16697,N_12796,N_12539);
nand U16698 (N_16698,N_14367,N_15327);
or U16699 (N_16699,N_14824,N_13709);
or U16700 (N_16700,N_13211,N_12656);
xor U16701 (N_16701,N_13320,N_14361);
and U16702 (N_16702,N_13895,N_14292);
xnor U16703 (N_16703,N_13312,N_13809);
xor U16704 (N_16704,N_14443,N_14337);
and U16705 (N_16705,N_13734,N_12793);
nor U16706 (N_16706,N_15500,N_14612);
and U16707 (N_16707,N_13827,N_13513);
xnor U16708 (N_16708,N_14315,N_12729);
nand U16709 (N_16709,N_12707,N_13795);
nor U16710 (N_16710,N_13998,N_12585);
nand U16711 (N_16711,N_14602,N_14151);
and U16712 (N_16712,N_14336,N_12619);
xor U16713 (N_16713,N_12971,N_13100);
or U16714 (N_16714,N_12751,N_13392);
nand U16715 (N_16715,N_14511,N_13891);
nor U16716 (N_16716,N_14737,N_12821);
nor U16717 (N_16717,N_13326,N_14074);
xnor U16718 (N_16718,N_14962,N_12895);
xnor U16719 (N_16719,N_14664,N_12527);
xnor U16720 (N_16720,N_15463,N_15068);
or U16721 (N_16721,N_14732,N_13653);
xor U16722 (N_16722,N_13317,N_13304);
xor U16723 (N_16723,N_15606,N_14613);
nand U16724 (N_16724,N_14252,N_14423);
nand U16725 (N_16725,N_12748,N_14058);
nor U16726 (N_16726,N_13545,N_14617);
nand U16727 (N_16727,N_14943,N_14294);
xor U16728 (N_16728,N_15596,N_12725);
xnor U16729 (N_16729,N_13182,N_13993);
and U16730 (N_16730,N_14650,N_13690);
xnor U16731 (N_16731,N_15015,N_14846);
nand U16732 (N_16732,N_12647,N_14707);
or U16733 (N_16733,N_12596,N_15274);
xor U16734 (N_16734,N_12778,N_14646);
xnor U16735 (N_16735,N_15591,N_14778);
nand U16736 (N_16736,N_15316,N_15324);
nand U16737 (N_16737,N_13882,N_14955);
and U16738 (N_16738,N_15250,N_14757);
nand U16739 (N_16739,N_13424,N_13663);
or U16740 (N_16740,N_12576,N_15355);
and U16741 (N_16741,N_15233,N_15556);
or U16742 (N_16742,N_12529,N_12577);
nor U16743 (N_16743,N_12944,N_13771);
nand U16744 (N_16744,N_12514,N_12905);
and U16745 (N_16745,N_12603,N_12946);
xnor U16746 (N_16746,N_12541,N_12579);
nand U16747 (N_16747,N_15236,N_13303);
nor U16748 (N_16748,N_14250,N_15505);
or U16749 (N_16749,N_13777,N_14493);
nand U16750 (N_16750,N_14329,N_13176);
nor U16751 (N_16751,N_13518,N_14496);
nor U16752 (N_16752,N_13810,N_12838);
and U16753 (N_16753,N_15077,N_14560);
nor U16754 (N_16754,N_13783,N_15343);
and U16755 (N_16755,N_13592,N_15131);
or U16756 (N_16756,N_14563,N_15283);
or U16757 (N_16757,N_13456,N_15576);
and U16758 (N_16758,N_13301,N_14903);
nor U16759 (N_16759,N_14744,N_13790);
xor U16760 (N_16760,N_13423,N_13965);
xor U16761 (N_16761,N_13322,N_14258);
and U16762 (N_16762,N_13792,N_15450);
or U16763 (N_16763,N_14402,N_14991);
xnor U16764 (N_16764,N_13945,N_15024);
nor U16765 (N_16765,N_14164,N_13673);
xor U16766 (N_16766,N_13631,N_13971);
or U16767 (N_16767,N_14066,N_13847);
xor U16768 (N_16768,N_14792,N_12605);
xor U16769 (N_16769,N_14111,N_15375);
nor U16770 (N_16770,N_13901,N_13850);
or U16771 (N_16771,N_13711,N_14310);
nor U16772 (N_16772,N_15443,N_13467);
and U16773 (N_16773,N_13381,N_14774);
and U16774 (N_16774,N_15525,N_13331);
or U16775 (N_16775,N_12676,N_12826);
and U16776 (N_16776,N_15105,N_14861);
nand U16777 (N_16777,N_12853,N_13849);
nand U16778 (N_16778,N_13841,N_13517);
xor U16779 (N_16779,N_13615,N_14995);
xor U16780 (N_16780,N_14607,N_12780);
and U16781 (N_16781,N_14508,N_15102);
xnor U16782 (N_16782,N_14731,N_14582);
and U16783 (N_16783,N_13422,N_13511);
or U16784 (N_16784,N_15060,N_14927);
xnor U16785 (N_16785,N_12628,N_13459);
nor U16786 (N_16786,N_15138,N_14976);
nor U16787 (N_16787,N_14850,N_13078);
nor U16788 (N_16788,N_13907,N_13166);
or U16789 (N_16789,N_12839,N_14067);
and U16790 (N_16790,N_14874,N_15422);
nand U16791 (N_16791,N_12738,N_13972);
nand U16792 (N_16792,N_14505,N_12973);
nand U16793 (N_16793,N_13825,N_12739);
nand U16794 (N_16794,N_15614,N_15229);
nand U16795 (N_16795,N_14763,N_14285);
nand U16796 (N_16796,N_14747,N_13389);
and U16797 (N_16797,N_13226,N_13162);
or U16798 (N_16798,N_14695,N_14180);
nor U16799 (N_16799,N_12864,N_13453);
and U16800 (N_16800,N_14978,N_14289);
xnor U16801 (N_16801,N_15210,N_12975);
and U16802 (N_16802,N_14709,N_13802);
xnor U16803 (N_16803,N_14660,N_12922);
nor U16804 (N_16804,N_15390,N_15394);
xor U16805 (N_16805,N_12632,N_14203);
and U16806 (N_16806,N_14552,N_12847);
or U16807 (N_16807,N_12736,N_13474);
xnor U16808 (N_16808,N_13994,N_15092);
and U16809 (N_16809,N_14251,N_13787);
or U16810 (N_16810,N_14497,N_13741);
nand U16811 (N_16811,N_13597,N_12945);
nor U16812 (N_16812,N_15368,N_12597);
and U16813 (N_16813,N_14131,N_14459);
and U16814 (N_16814,N_13593,N_15517);
or U16815 (N_16815,N_14044,N_13587);
nor U16816 (N_16816,N_14183,N_13324);
or U16817 (N_16817,N_14895,N_12836);
nand U16818 (N_16818,N_14267,N_13652);
nand U16819 (N_16819,N_12822,N_15480);
or U16820 (N_16820,N_13951,N_13377);
nor U16821 (N_16821,N_14652,N_14387);
nand U16822 (N_16822,N_13637,N_13696);
or U16823 (N_16823,N_14398,N_14710);
xnor U16824 (N_16824,N_14313,N_15109);
or U16825 (N_16825,N_13099,N_13450);
nand U16826 (N_16826,N_15019,N_14452);
nand U16827 (N_16827,N_15136,N_14967);
and U16828 (N_16828,N_13057,N_12808);
or U16829 (N_16829,N_14775,N_12787);
nor U16830 (N_16830,N_15146,N_14163);
and U16831 (N_16831,N_13758,N_15440);
xor U16832 (N_16832,N_15156,N_14634);
nor U16833 (N_16833,N_12962,N_14126);
xnor U16834 (N_16834,N_12609,N_15468);
xnor U16835 (N_16835,N_14192,N_12616);
and U16836 (N_16836,N_13095,N_14487);
xor U16837 (N_16837,N_14447,N_15337);
nand U16838 (N_16838,N_14942,N_15310);
nor U16839 (N_16839,N_14401,N_15416);
nand U16840 (N_16840,N_12524,N_14690);
xor U16841 (N_16841,N_12611,N_13121);
nor U16842 (N_16842,N_13208,N_15084);
and U16843 (N_16843,N_12988,N_12635);
nor U16844 (N_16844,N_13137,N_14614);
nand U16845 (N_16845,N_14438,N_12517);
xor U16846 (N_16846,N_15580,N_15120);
xnor U16847 (N_16847,N_15016,N_13433);
xnor U16848 (N_16848,N_14691,N_12548);
or U16849 (N_16849,N_13756,N_14242);
nand U16850 (N_16850,N_13613,N_13482);
xnor U16851 (N_16851,N_13623,N_15244);
nand U16852 (N_16852,N_14897,N_15433);
nand U16853 (N_16853,N_15498,N_15103);
and U16854 (N_16854,N_14701,N_15037);
or U16855 (N_16855,N_12930,N_13800);
xor U16856 (N_16856,N_13835,N_12622);
and U16857 (N_16857,N_12648,N_15410);
nor U16858 (N_16858,N_15566,N_13010);
or U16859 (N_16859,N_13740,N_14130);
or U16860 (N_16860,N_15171,N_14541);
nor U16861 (N_16861,N_13437,N_12715);
nor U16862 (N_16862,N_14188,N_15128);
or U16863 (N_16863,N_14317,N_13264);
nand U16864 (N_16864,N_14135,N_13724);
and U16865 (N_16865,N_13156,N_14110);
nor U16866 (N_16866,N_13470,N_13130);
and U16867 (N_16867,N_15511,N_13753);
xnor U16868 (N_16868,N_13946,N_13936);
or U16869 (N_16869,N_13523,N_14378);
xnor U16870 (N_16870,N_13649,N_14491);
xor U16871 (N_16871,N_15360,N_13776);
nor U16872 (N_16872,N_14142,N_15205);
or U16873 (N_16873,N_15532,N_14735);
and U16874 (N_16874,N_13088,N_13750);
nor U16875 (N_16875,N_14173,N_12867);
or U16876 (N_16876,N_13656,N_13280);
xnor U16877 (N_16877,N_12649,N_13201);
or U16878 (N_16878,N_15453,N_15342);
or U16879 (N_16879,N_14502,N_12744);
or U16880 (N_16880,N_15294,N_13958);
xnor U16881 (N_16881,N_13909,N_12845);
or U16882 (N_16882,N_12594,N_13184);
nand U16883 (N_16883,N_12811,N_12918);
xnor U16884 (N_16884,N_12565,N_14706);
or U16885 (N_16885,N_14830,N_14008);
or U16886 (N_16886,N_14577,N_13562);
and U16887 (N_16887,N_15260,N_14182);
or U16888 (N_16888,N_13478,N_14306);
or U16889 (N_16889,N_12941,N_15339);
nand U16890 (N_16890,N_12940,N_13949);
nand U16891 (N_16891,N_14687,N_14076);
nor U16892 (N_16892,N_13048,N_13979);
xor U16893 (N_16893,N_15032,N_12719);
nor U16894 (N_16894,N_15152,N_14929);
nand U16895 (N_16895,N_12929,N_12723);
or U16896 (N_16896,N_14350,N_15217);
xnor U16897 (N_16897,N_14271,N_13360);
and U16898 (N_16898,N_14918,N_15237);
or U16899 (N_16899,N_15127,N_14421);
or U16900 (N_16900,N_12920,N_15464);
nor U16901 (N_16901,N_13729,N_12598);
nor U16902 (N_16902,N_13200,N_13330);
nor U16903 (N_16903,N_14771,N_12522);
xor U16904 (N_16904,N_14851,N_13659);
or U16905 (N_16905,N_13658,N_14684);
or U16906 (N_16906,N_14274,N_12556);
nor U16907 (N_16907,N_15590,N_14144);
or U16908 (N_16908,N_13216,N_14206);
nand U16909 (N_16909,N_12685,N_14393);
xor U16910 (N_16910,N_15526,N_13142);
nor U16911 (N_16911,N_14734,N_14312);
or U16912 (N_16912,N_14225,N_12815);
nand U16913 (N_16913,N_13885,N_12695);
and U16914 (N_16914,N_14040,N_14418);
nor U16915 (N_16915,N_14600,N_14205);
or U16916 (N_16916,N_12618,N_12554);
and U16917 (N_16917,N_15530,N_14201);
nor U16918 (N_16918,N_12843,N_14479);
and U16919 (N_16919,N_14114,N_12709);
nand U16920 (N_16920,N_15549,N_15186);
xor U16921 (N_16921,N_12507,N_12742);
nand U16922 (N_16922,N_13594,N_14803);
or U16923 (N_16923,N_13151,N_14490);
xor U16924 (N_16924,N_13285,N_12621);
or U16925 (N_16925,N_15397,N_15180);
xnor U16926 (N_16926,N_15070,N_14259);
nand U16927 (N_16927,N_13257,N_13550);
nand U16928 (N_16928,N_13101,N_14981);
nor U16929 (N_16929,N_13373,N_15582);
xnor U16930 (N_16930,N_15112,N_13308);
nand U16931 (N_16931,N_13905,N_14992);
and U16932 (N_16932,N_14241,N_13408);
xnor U16933 (N_16933,N_15142,N_12718);
nor U16934 (N_16934,N_14453,N_13438);
and U16935 (N_16935,N_12501,N_13954);
and U16936 (N_16936,N_13041,N_14170);
xnor U16937 (N_16937,N_15369,N_14307);
nor U16938 (N_16938,N_14884,N_15041);
nand U16939 (N_16939,N_15214,N_14346);
nand U16940 (N_16940,N_13051,N_13970);
xor U16941 (N_16941,N_14549,N_14019);
and U16942 (N_16942,N_15115,N_15134);
nand U16943 (N_16943,N_15605,N_13692);
or U16944 (N_16944,N_14356,N_14750);
xor U16945 (N_16945,N_13846,N_13630);
nand U16946 (N_16946,N_12533,N_13601);
nand U16947 (N_16947,N_15215,N_13430);
and U16948 (N_16948,N_14908,N_13747);
xor U16949 (N_16949,N_15485,N_14322);
and U16950 (N_16950,N_14239,N_15438);
xor U16951 (N_16951,N_13713,N_14325);
nor U16952 (N_16952,N_12893,N_13410);
xnor U16953 (N_16953,N_14700,N_13153);
nand U16954 (N_16954,N_15529,N_13371);
and U16955 (N_16955,N_13196,N_15224);
or U16956 (N_16956,N_13062,N_15293);
or U16957 (N_16957,N_12535,N_14537);
nand U16958 (N_16958,N_14413,N_13575);
xnor U16959 (N_16959,N_15173,N_13421);
nand U16960 (N_16960,N_14794,N_12537);
and U16961 (N_16961,N_15429,N_13798);
nor U16962 (N_16962,N_13669,N_14669);
and U16963 (N_16963,N_13822,N_14576);
nand U16964 (N_16964,N_13995,N_13778);
or U16965 (N_16965,N_13428,N_13363);
nand U16966 (N_16966,N_13614,N_15277);
and U16967 (N_16967,N_13167,N_13282);
nor U16968 (N_16968,N_15093,N_13252);
or U16969 (N_16969,N_14915,N_14996);
nand U16970 (N_16970,N_13000,N_14345);
nand U16971 (N_16971,N_15567,N_14237);
xor U16972 (N_16972,N_12557,N_12670);
or U16973 (N_16973,N_12547,N_12953);
and U16974 (N_16974,N_14987,N_15076);
nand U16975 (N_16975,N_14364,N_13860);
xor U16976 (N_16976,N_12712,N_13625);
or U16977 (N_16977,N_13265,N_13344);
and U16978 (N_16978,N_15311,N_15449);
xor U16979 (N_16979,N_14153,N_13417);
nand U16980 (N_16980,N_14197,N_13286);
nand U16981 (N_16981,N_13284,N_15042);
xor U16982 (N_16982,N_15007,N_13169);
or U16983 (N_16983,N_15064,N_14510);
nand U16984 (N_16984,N_13350,N_13963);
xnor U16985 (N_16985,N_15284,N_14049);
or U16986 (N_16986,N_13832,N_13629);
and U16987 (N_16987,N_14100,N_13999);
nor U16988 (N_16988,N_15108,N_14116);
xor U16989 (N_16989,N_15159,N_15240);
xnor U16990 (N_16990,N_13948,N_14579);
nor U16991 (N_16991,N_13906,N_15607);
and U16992 (N_16992,N_14115,N_12967);
or U16993 (N_16993,N_12792,N_15239);
xnor U16994 (N_16994,N_12634,N_13081);
nand U16995 (N_16995,N_15374,N_14140);
nand U16996 (N_16996,N_12604,N_14944);
or U16997 (N_16997,N_14584,N_15391);
or U16998 (N_16998,N_13190,N_15140);
nor U16999 (N_16999,N_13977,N_15484);
or U17000 (N_17000,N_14109,N_12711);
and U17001 (N_17001,N_14585,N_14261);
nand U17002 (N_17002,N_14833,N_14606);
nor U17003 (N_17003,N_13764,N_14095);
xnor U17004 (N_17004,N_14647,N_14156);
nor U17005 (N_17005,N_14649,N_14852);
nand U17006 (N_17006,N_15262,N_14124);
nor U17007 (N_17007,N_15426,N_14229);
xor U17008 (N_17008,N_14688,N_14377);
or U17009 (N_17009,N_12528,N_13468);
nand U17010 (N_17010,N_15255,N_15320);
or U17011 (N_17011,N_15023,N_13912);
nand U17012 (N_17012,N_15195,N_15522);
nor U17013 (N_17013,N_14328,N_14655);
nand U17014 (N_17014,N_12581,N_15381);
nor U17015 (N_17015,N_13247,N_14435);
nand U17016 (N_17016,N_13045,N_14676);
xor U17017 (N_17017,N_14539,N_12623);
xnor U17018 (N_17018,N_15238,N_15474);
or U17019 (N_17019,N_14723,N_13662);
nor U17020 (N_17020,N_14146,N_15223);
or U17021 (N_17021,N_14692,N_13300);
nor U17022 (N_17022,N_14521,N_12927);
or U17023 (N_17023,N_13774,N_13962);
xnor U17024 (N_17024,N_14913,N_12752);
xnor U17025 (N_17025,N_14532,N_12823);
xnor U17026 (N_17026,N_13427,N_14586);
xnor U17027 (N_17027,N_13241,N_13749);
or U17028 (N_17028,N_14760,N_14773);
and U17029 (N_17029,N_14637,N_12960);
or U17030 (N_17030,N_14128,N_12701);
and U17031 (N_17031,N_13031,N_13384);
nor U17032 (N_17032,N_13738,N_12504);
nor U17033 (N_17033,N_14516,N_13851);
xnor U17034 (N_17034,N_12999,N_13725);
nand U17035 (N_17035,N_12553,N_13367);
nand U17036 (N_17036,N_14970,N_15199);
nor U17037 (N_17037,N_12794,N_14623);
nor U17038 (N_17038,N_13555,N_13052);
or U17039 (N_17039,N_13079,N_15562);
nand U17040 (N_17040,N_14715,N_12668);
or U17041 (N_17041,N_13657,N_12733);
or U17042 (N_17042,N_14078,N_13154);
or U17043 (N_17043,N_13534,N_15312);
or U17044 (N_17044,N_13083,N_14038);
or U17045 (N_17045,N_15564,N_15201);
xnor U17046 (N_17046,N_14301,N_15593);
or U17047 (N_17047,N_13093,N_14155);
nand U17048 (N_17048,N_13676,N_14429);
and U17049 (N_17049,N_13299,N_15421);
nand U17050 (N_17050,N_14963,N_14445);
nand U17051 (N_17051,N_13826,N_14408);
xnor U17052 (N_17052,N_13432,N_12641);
and U17053 (N_17053,N_12872,N_14484);
nor U17054 (N_17054,N_13342,N_13181);
xnor U17055 (N_17055,N_13599,N_14195);
nor U17056 (N_17056,N_13402,N_13680);
xnor U17057 (N_17057,N_14898,N_14597);
nor U17058 (N_17058,N_13329,N_12813);
or U17059 (N_17059,N_14291,N_14711);
xor U17060 (N_17060,N_15253,N_13275);
or U17061 (N_17061,N_15176,N_14223);
or U17062 (N_17062,N_12912,N_13622);
or U17063 (N_17063,N_12747,N_15446);
or U17064 (N_17064,N_13619,N_15278);
or U17065 (N_17065,N_15174,N_13546);
or U17066 (N_17066,N_12848,N_13487);
nand U17067 (N_17067,N_14375,N_12536);
or U17068 (N_17068,N_15431,N_14673);
and U17069 (N_17069,N_13259,N_14595);
xnor U17070 (N_17070,N_14966,N_12970);
nand U17071 (N_17071,N_15196,N_12842);
nor U17072 (N_17072,N_12710,N_14031);
and U17073 (N_17073,N_14495,N_15097);
nand U17074 (N_17074,N_14618,N_12989);
nor U17075 (N_17075,N_13267,N_15123);
nand U17076 (N_17076,N_15247,N_13853);
and U17077 (N_17077,N_12803,N_13804);
nor U17078 (N_17078,N_14619,N_13799);
nand U17079 (N_17079,N_14821,N_13984);
nor U17080 (N_17080,N_12555,N_13479);
nand U17081 (N_17081,N_13644,N_14845);
nand U17082 (N_17082,N_15392,N_14405);
nor U17083 (N_17083,N_13580,N_14697);
xor U17084 (N_17084,N_14658,N_14189);
nand U17085 (N_17085,N_14725,N_13770);
xor U17086 (N_17086,N_14342,N_12860);
nand U17087 (N_17087,N_13191,N_14779);
or U17088 (N_17088,N_12799,N_15005);
nor U17089 (N_17089,N_15389,N_13595);
nor U17090 (N_17090,N_15555,N_14099);
nand U17091 (N_17091,N_12639,N_13315);
nand U17092 (N_17092,N_15303,N_13485);
nor U17093 (N_17093,N_14515,N_15400);
or U17094 (N_17094,N_14157,N_12519);
and U17095 (N_17095,N_14513,N_15516);
xor U17096 (N_17096,N_14059,N_15178);
or U17097 (N_17097,N_14084,N_14672);
nand U17098 (N_17098,N_14353,N_15393);
nor U17099 (N_17099,N_14238,N_14082);
nand U17100 (N_17100,N_13452,N_13278);
nor U17101 (N_17101,N_14568,N_15044);
nand U17102 (N_17102,N_15072,N_15028);
and U17103 (N_17103,N_14588,N_14162);
nand U17104 (N_17104,N_14023,N_13291);
nand U17105 (N_17105,N_12854,N_15384);
or U17106 (N_17106,N_13023,N_13340);
nand U17107 (N_17107,N_13989,N_13290);
xnor U17108 (N_17108,N_13687,N_13435);
xnor U17109 (N_17109,N_13262,N_13463);
nor U17110 (N_17110,N_14844,N_13001);
nor U17111 (N_17111,N_15506,N_14777);
nor U17112 (N_17112,N_12698,N_13572);
or U17113 (N_17113,N_13205,N_13109);
and U17114 (N_17114,N_15228,N_14321);
and U17115 (N_17115,N_12888,N_14354);
and U17116 (N_17116,N_13780,N_14808);
or U17117 (N_17117,N_12644,N_12564);
nand U17118 (N_17118,N_14609,N_14029);
xor U17119 (N_17119,N_15424,N_12890);
or U17120 (N_17120,N_13716,N_12627);
nand U17121 (N_17121,N_13744,N_12840);
nor U17122 (N_17122,N_14712,N_15014);
nor U17123 (N_17123,N_13189,N_13094);
nand U17124 (N_17124,N_15149,N_14512);
and U17125 (N_17125,N_14007,N_14683);
nor U17126 (N_17126,N_12750,N_13554);
or U17127 (N_17127,N_12881,N_14278);
and U17128 (N_17128,N_14540,N_14665);
or U17129 (N_17129,N_15341,N_14465);
xor U17130 (N_17130,N_15145,N_15586);
nand U17131 (N_17131,N_15331,N_15447);
or U17132 (N_17132,N_14425,N_14024);
xor U17133 (N_17133,N_13394,N_13833);
xor U17134 (N_17134,N_15492,N_14492);
nand U17135 (N_17135,N_14829,N_12606);
nand U17136 (N_17136,N_12570,N_12814);
or U17137 (N_17137,N_15208,N_14959);
nand U17138 (N_17138,N_13661,N_12824);
nand U17139 (N_17139,N_13068,N_13248);
or U17140 (N_17140,N_15435,N_12692);
or U17141 (N_17141,N_13884,N_12834);
and U17142 (N_17142,N_13382,N_13843);
and U17143 (N_17143,N_14158,N_14632);
nand U17144 (N_17144,N_14273,N_13768);
and U17145 (N_17145,N_14686,N_13682);
or U17146 (N_17146,N_14077,N_14776);
nand U17147 (N_17147,N_15306,N_13198);
nand U17148 (N_17148,N_13489,N_15362);
and U17149 (N_17149,N_15469,N_14456);
and U17150 (N_17150,N_14849,N_13541);
and U17151 (N_17151,N_13343,N_13143);
xnor U17152 (N_17152,N_15371,N_14355);
nor U17153 (N_17153,N_13533,N_15216);
nand U17154 (N_17154,N_15086,N_15296);
and U17155 (N_17155,N_13654,N_13836);
nand U17156 (N_17156,N_15594,N_13873);
nor U17157 (N_17157,N_12775,N_13034);
nor U17158 (N_17158,N_15462,N_15538);
or U17159 (N_17159,N_13717,N_14302);
and U17160 (N_17160,N_14362,N_12700);
nand U17161 (N_17161,N_14269,N_14108);
xor U17162 (N_17162,N_15259,N_15621);
nor U17163 (N_17163,N_14841,N_14749);
xor U17164 (N_17164,N_15353,N_15584);
nor U17165 (N_17165,N_13111,N_14553);
nand U17166 (N_17166,N_15067,N_14702);
nand U17167 (N_17167,N_15298,N_12545);
xnor U17168 (N_17168,N_15280,N_13011);
and U17169 (N_17169,N_14347,N_13116);
nor U17170 (N_17170,N_14855,N_12508);
or U17171 (N_17171,N_12759,N_12981);
xnor U17172 (N_17172,N_14454,N_13879);
nor U17173 (N_17173,N_13192,N_15486);
and U17174 (N_17174,N_13237,N_13215);
and U17175 (N_17175,N_14525,N_14063);
nand U17176 (N_17176,N_13362,N_12502);
xor U17177 (N_17177,N_14791,N_14790);
nand U17178 (N_17178,N_13596,N_15100);
and U17179 (N_17179,N_14352,N_14628);
and U17180 (N_17180,N_14910,N_14909);
and U17181 (N_17181,N_14499,N_12560);
xor U17182 (N_17182,N_13359,N_12998);
xor U17183 (N_17183,N_15295,N_13721);
nor U17184 (N_17184,N_13544,N_14290);
nor U17185 (N_17185,N_13490,N_13956);
nand U17186 (N_17186,N_15211,N_14722);
and U17187 (N_17187,N_13451,N_12904);
xor U17188 (N_17188,N_13513,N_15029);
or U17189 (N_17189,N_13158,N_15069);
nor U17190 (N_17190,N_15605,N_13695);
nand U17191 (N_17191,N_13482,N_14828);
nor U17192 (N_17192,N_14213,N_15008);
or U17193 (N_17193,N_13733,N_14930);
nor U17194 (N_17194,N_15290,N_12569);
nand U17195 (N_17195,N_13744,N_13311);
or U17196 (N_17196,N_15492,N_13590);
nand U17197 (N_17197,N_13380,N_12587);
nor U17198 (N_17198,N_14270,N_15185);
or U17199 (N_17199,N_13539,N_12558);
and U17200 (N_17200,N_14223,N_14148);
nor U17201 (N_17201,N_14249,N_13060);
nor U17202 (N_17202,N_13527,N_13957);
or U17203 (N_17203,N_13052,N_13021);
nor U17204 (N_17204,N_15209,N_14187);
nor U17205 (N_17205,N_13918,N_15435);
or U17206 (N_17206,N_13584,N_15407);
nor U17207 (N_17207,N_14165,N_13224);
and U17208 (N_17208,N_13955,N_15125);
xor U17209 (N_17209,N_13808,N_13255);
or U17210 (N_17210,N_13530,N_12546);
nand U17211 (N_17211,N_13617,N_13778);
and U17212 (N_17212,N_12718,N_13735);
and U17213 (N_17213,N_12578,N_13821);
and U17214 (N_17214,N_12505,N_14756);
xnor U17215 (N_17215,N_15390,N_14498);
nand U17216 (N_17216,N_15393,N_12513);
or U17217 (N_17217,N_12992,N_14299);
nand U17218 (N_17218,N_14647,N_14455);
nand U17219 (N_17219,N_15121,N_14830);
xor U17220 (N_17220,N_12671,N_13774);
and U17221 (N_17221,N_12768,N_13787);
or U17222 (N_17222,N_13412,N_15317);
nor U17223 (N_17223,N_12536,N_14623);
nor U17224 (N_17224,N_12645,N_14829);
nand U17225 (N_17225,N_14165,N_14947);
xor U17226 (N_17226,N_13883,N_14739);
nand U17227 (N_17227,N_14914,N_12656);
or U17228 (N_17228,N_12660,N_15272);
or U17229 (N_17229,N_14809,N_13211);
and U17230 (N_17230,N_14008,N_14691);
or U17231 (N_17231,N_13509,N_12846);
and U17232 (N_17232,N_15397,N_13973);
or U17233 (N_17233,N_15277,N_14081);
xnor U17234 (N_17234,N_14318,N_15116);
nand U17235 (N_17235,N_13834,N_12919);
or U17236 (N_17236,N_12655,N_15283);
nand U17237 (N_17237,N_14783,N_14574);
nor U17238 (N_17238,N_15471,N_13861);
nor U17239 (N_17239,N_12603,N_13531);
nor U17240 (N_17240,N_13452,N_13918);
and U17241 (N_17241,N_13694,N_13341);
nor U17242 (N_17242,N_14649,N_13334);
nor U17243 (N_17243,N_13475,N_12800);
nand U17244 (N_17244,N_13826,N_12600);
nor U17245 (N_17245,N_14505,N_15533);
nor U17246 (N_17246,N_13381,N_12973);
xor U17247 (N_17247,N_13312,N_12758);
nor U17248 (N_17248,N_13914,N_12651);
nand U17249 (N_17249,N_13418,N_13505);
nor U17250 (N_17250,N_13150,N_12721);
and U17251 (N_17251,N_14796,N_15542);
and U17252 (N_17252,N_14022,N_13239);
xnor U17253 (N_17253,N_12718,N_14579);
nand U17254 (N_17254,N_12543,N_15445);
xor U17255 (N_17255,N_12768,N_14203);
and U17256 (N_17256,N_14845,N_14823);
nor U17257 (N_17257,N_15067,N_12811);
nand U17258 (N_17258,N_14721,N_14899);
xnor U17259 (N_17259,N_13993,N_15619);
or U17260 (N_17260,N_12563,N_13518);
or U17261 (N_17261,N_14245,N_14024);
nand U17262 (N_17262,N_13267,N_13898);
or U17263 (N_17263,N_13258,N_14112);
nor U17264 (N_17264,N_12737,N_13229);
and U17265 (N_17265,N_14636,N_13181);
nor U17266 (N_17266,N_12636,N_13108);
nor U17267 (N_17267,N_14477,N_13422);
and U17268 (N_17268,N_13915,N_14109);
xor U17269 (N_17269,N_14774,N_13794);
nor U17270 (N_17270,N_13348,N_13394);
xor U17271 (N_17271,N_14468,N_14106);
xnor U17272 (N_17272,N_14866,N_14121);
and U17273 (N_17273,N_13407,N_14411);
nor U17274 (N_17274,N_15183,N_13211);
xor U17275 (N_17275,N_12656,N_13155);
nand U17276 (N_17276,N_15240,N_14051);
and U17277 (N_17277,N_14336,N_12872);
or U17278 (N_17278,N_13671,N_14910);
or U17279 (N_17279,N_14882,N_15448);
nor U17280 (N_17280,N_12890,N_15298);
or U17281 (N_17281,N_13867,N_14902);
nor U17282 (N_17282,N_12638,N_14540);
xor U17283 (N_17283,N_13195,N_12587);
nor U17284 (N_17284,N_14997,N_13897);
xor U17285 (N_17285,N_13472,N_13579);
or U17286 (N_17286,N_15492,N_12774);
or U17287 (N_17287,N_15196,N_14044);
or U17288 (N_17288,N_13321,N_13600);
or U17289 (N_17289,N_13601,N_15452);
nand U17290 (N_17290,N_12887,N_14205);
or U17291 (N_17291,N_12938,N_13931);
nor U17292 (N_17292,N_15223,N_12952);
nand U17293 (N_17293,N_13127,N_13536);
or U17294 (N_17294,N_15013,N_15528);
nand U17295 (N_17295,N_13363,N_15615);
nor U17296 (N_17296,N_12829,N_12807);
nand U17297 (N_17297,N_14793,N_13944);
nand U17298 (N_17298,N_14996,N_14444);
nand U17299 (N_17299,N_14575,N_13256);
nor U17300 (N_17300,N_14143,N_12899);
nor U17301 (N_17301,N_15044,N_15404);
xor U17302 (N_17302,N_14761,N_12564);
xnor U17303 (N_17303,N_15623,N_15452);
and U17304 (N_17304,N_13509,N_14017);
or U17305 (N_17305,N_13301,N_12781);
nor U17306 (N_17306,N_15177,N_13828);
nor U17307 (N_17307,N_13430,N_13688);
or U17308 (N_17308,N_13574,N_15082);
and U17309 (N_17309,N_13966,N_13377);
or U17310 (N_17310,N_13045,N_15352);
nand U17311 (N_17311,N_13981,N_14265);
and U17312 (N_17312,N_14143,N_13758);
and U17313 (N_17313,N_14338,N_14330);
xor U17314 (N_17314,N_13245,N_13796);
nand U17315 (N_17315,N_12746,N_13540);
or U17316 (N_17316,N_13588,N_13137);
xnor U17317 (N_17317,N_15560,N_12543);
and U17318 (N_17318,N_13999,N_14862);
or U17319 (N_17319,N_15153,N_13104);
nand U17320 (N_17320,N_13203,N_14381);
nand U17321 (N_17321,N_15003,N_12782);
or U17322 (N_17322,N_14894,N_13699);
nor U17323 (N_17323,N_13127,N_14765);
nor U17324 (N_17324,N_15286,N_15018);
nand U17325 (N_17325,N_14390,N_13736);
xnor U17326 (N_17326,N_13218,N_12912);
xnor U17327 (N_17327,N_14687,N_15142);
xnor U17328 (N_17328,N_13302,N_14273);
or U17329 (N_17329,N_14989,N_12954);
nor U17330 (N_17330,N_15260,N_14934);
xor U17331 (N_17331,N_13979,N_15318);
or U17332 (N_17332,N_12989,N_13979);
nor U17333 (N_17333,N_13196,N_14431);
xor U17334 (N_17334,N_14797,N_13933);
and U17335 (N_17335,N_12518,N_13679);
and U17336 (N_17336,N_13918,N_14282);
xnor U17337 (N_17337,N_13613,N_14457);
nand U17338 (N_17338,N_14642,N_14122);
nor U17339 (N_17339,N_14004,N_13646);
or U17340 (N_17340,N_14599,N_14005);
xnor U17341 (N_17341,N_13403,N_13755);
nand U17342 (N_17342,N_15332,N_15271);
nand U17343 (N_17343,N_14426,N_13784);
xnor U17344 (N_17344,N_14276,N_14867);
or U17345 (N_17345,N_14913,N_12800);
nand U17346 (N_17346,N_13734,N_13083);
or U17347 (N_17347,N_15513,N_14444);
and U17348 (N_17348,N_15011,N_13435);
xnor U17349 (N_17349,N_13434,N_13166);
xnor U17350 (N_17350,N_12619,N_13760);
and U17351 (N_17351,N_15096,N_14432);
xor U17352 (N_17352,N_12946,N_12543);
or U17353 (N_17353,N_14801,N_15498);
or U17354 (N_17354,N_14828,N_14004);
or U17355 (N_17355,N_13589,N_13093);
or U17356 (N_17356,N_14247,N_13145);
xor U17357 (N_17357,N_14667,N_14738);
and U17358 (N_17358,N_15595,N_13546);
xnor U17359 (N_17359,N_12705,N_13679);
or U17360 (N_17360,N_13372,N_15074);
xnor U17361 (N_17361,N_12751,N_12594);
xnor U17362 (N_17362,N_13274,N_14122);
nand U17363 (N_17363,N_14118,N_13935);
and U17364 (N_17364,N_13106,N_13521);
and U17365 (N_17365,N_13944,N_15460);
nand U17366 (N_17366,N_15348,N_14677);
or U17367 (N_17367,N_12986,N_14260);
nor U17368 (N_17368,N_15475,N_13820);
xor U17369 (N_17369,N_14395,N_15348);
xor U17370 (N_17370,N_12639,N_14981);
or U17371 (N_17371,N_12788,N_15224);
nand U17372 (N_17372,N_12922,N_13780);
xor U17373 (N_17373,N_12699,N_14789);
or U17374 (N_17374,N_12732,N_14699);
xnor U17375 (N_17375,N_15113,N_15552);
or U17376 (N_17376,N_15058,N_14896);
or U17377 (N_17377,N_15416,N_13314);
and U17378 (N_17378,N_15622,N_13282);
or U17379 (N_17379,N_14443,N_15357);
and U17380 (N_17380,N_13264,N_12757);
nand U17381 (N_17381,N_14025,N_14887);
nand U17382 (N_17382,N_15614,N_15236);
nor U17383 (N_17383,N_14091,N_14895);
or U17384 (N_17384,N_14600,N_15363);
nand U17385 (N_17385,N_14017,N_12909);
and U17386 (N_17386,N_13298,N_12567);
or U17387 (N_17387,N_15175,N_12976);
xnor U17388 (N_17388,N_14184,N_13756);
xnor U17389 (N_17389,N_15305,N_15135);
nor U17390 (N_17390,N_15489,N_14247);
nor U17391 (N_17391,N_14659,N_13620);
or U17392 (N_17392,N_13492,N_14521);
nand U17393 (N_17393,N_14797,N_14260);
nor U17394 (N_17394,N_13282,N_13543);
nand U17395 (N_17395,N_13830,N_14354);
nand U17396 (N_17396,N_14341,N_13835);
nor U17397 (N_17397,N_13566,N_13115);
nor U17398 (N_17398,N_15550,N_13445);
and U17399 (N_17399,N_13296,N_14987);
or U17400 (N_17400,N_15315,N_15398);
nor U17401 (N_17401,N_12600,N_15421);
nor U17402 (N_17402,N_15091,N_13875);
nand U17403 (N_17403,N_14109,N_12504);
nor U17404 (N_17404,N_12547,N_13560);
and U17405 (N_17405,N_12972,N_14613);
xor U17406 (N_17406,N_13372,N_13389);
and U17407 (N_17407,N_12677,N_14080);
or U17408 (N_17408,N_15086,N_13951);
or U17409 (N_17409,N_13112,N_13917);
xnor U17410 (N_17410,N_14819,N_13944);
or U17411 (N_17411,N_15506,N_14932);
or U17412 (N_17412,N_15564,N_12787);
or U17413 (N_17413,N_12611,N_15221);
and U17414 (N_17414,N_13534,N_13824);
nor U17415 (N_17415,N_13288,N_15037);
nand U17416 (N_17416,N_14654,N_15283);
or U17417 (N_17417,N_14007,N_14880);
xor U17418 (N_17418,N_14081,N_15401);
or U17419 (N_17419,N_14343,N_15240);
or U17420 (N_17420,N_13332,N_14238);
or U17421 (N_17421,N_13679,N_15111);
or U17422 (N_17422,N_15163,N_15350);
or U17423 (N_17423,N_15379,N_12991);
nand U17424 (N_17424,N_15468,N_14174);
nor U17425 (N_17425,N_13951,N_14027);
xnor U17426 (N_17426,N_13635,N_14186);
xor U17427 (N_17427,N_13250,N_12996);
nand U17428 (N_17428,N_14857,N_12514);
or U17429 (N_17429,N_15606,N_14305);
nor U17430 (N_17430,N_12671,N_15090);
or U17431 (N_17431,N_12501,N_12625);
xnor U17432 (N_17432,N_14598,N_13299);
or U17433 (N_17433,N_14333,N_13841);
xnor U17434 (N_17434,N_12757,N_14197);
xor U17435 (N_17435,N_15150,N_14529);
xnor U17436 (N_17436,N_13051,N_15030);
xnor U17437 (N_17437,N_13112,N_13342);
or U17438 (N_17438,N_12950,N_15226);
nor U17439 (N_17439,N_14248,N_13971);
and U17440 (N_17440,N_14576,N_13708);
xnor U17441 (N_17441,N_15615,N_15572);
and U17442 (N_17442,N_13599,N_13072);
xor U17443 (N_17443,N_15103,N_13681);
nand U17444 (N_17444,N_14939,N_14776);
xnor U17445 (N_17445,N_13645,N_14758);
nand U17446 (N_17446,N_14819,N_14296);
or U17447 (N_17447,N_12747,N_14149);
xnor U17448 (N_17448,N_13710,N_14502);
or U17449 (N_17449,N_15094,N_14383);
nand U17450 (N_17450,N_13953,N_14391);
nor U17451 (N_17451,N_12554,N_14943);
nor U17452 (N_17452,N_12715,N_15271);
nor U17453 (N_17453,N_13954,N_15576);
xor U17454 (N_17454,N_14104,N_15277);
nand U17455 (N_17455,N_13010,N_13239);
or U17456 (N_17456,N_14175,N_13950);
nor U17457 (N_17457,N_13077,N_14148);
and U17458 (N_17458,N_12873,N_12811);
nor U17459 (N_17459,N_14004,N_12969);
nand U17460 (N_17460,N_12707,N_14327);
xor U17461 (N_17461,N_15166,N_14700);
or U17462 (N_17462,N_14116,N_13141);
and U17463 (N_17463,N_14717,N_14822);
or U17464 (N_17464,N_13375,N_15548);
nor U17465 (N_17465,N_15408,N_14727);
and U17466 (N_17466,N_12541,N_14952);
nor U17467 (N_17467,N_14142,N_15085);
or U17468 (N_17468,N_12761,N_15462);
nor U17469 (N_17469,N_13158,N_15247);
or U17470 (N_17470,N_13411,N_14852);
and U17471 (N_17471,N_13403,N_14192);
and U17472 (N_17472,N_13790,N_13040);
and U17473 (N_17473,N_13726,N_13111);
xnor U17474 (N_17474,N_13847,N_13947);
and U17475 (N_17475,N_14854,N_13796);
xnor U17476 (N_17476,N_13623,N_12685);
and U17477 (N_17477,N_13950,N_13350);
nand U17478 (N_17478,N_13194,N_13259);
xor U17479 (N_17479,N_15467,N_13987);
nor U17480 (N_17480,N_15102,N_12664);
nand U17481 (N_17481,N_15117,N_13286);
nand U17482 (N_17482,N_13061,N_14710);
xnor U17483 (N_17483,N_15562,N_14199);
or U17484 (N_17484,N_14606,N_14138);
or U17485 (N_17485,N_13422,N_15017);
nand U17486 (N_17486,N_13459,N_15279);
nor U17487 (N_17487,N_15221,N_13776);
nand U17488 (N_17488,N_14182,N_12517);
xnor U17489 (N_17489,N_15047,N_15594);
or U17490 (N_17490,N_14302,N_12568);
nor U17491 (N_17491,N_13059,N_13648);
or U17492 (N_17492,N_14123,N_14101);
and U17493 (N_17493,N_13653,N_15481);
xor U17494 (N_17494,N_15428,N_14050);
xnor U17495 (N_17495,N_15119,N_13310);
and U17496 (N_17496,N_13229,N_15193);
or U17497 (N_17497,N_13672,N_12855);
and U17498 (N_17498,N_14032,N_15464);
and U17499 (N_17499,N_15207,N_13213);
nor U17500 (N_17500,N_13881,N_12758);
and U17501 (N_17501,N_13749,N_12828);
xor U17502 (N_17502,N_15394,N_15572);
and U17503 (N_17503,N_13329,N_13222);
or U17504 (N_17504,N_13627,N_14611);
xnor U17505 (N_17505,N_15161,N_13229);
xnor U17506 (N_17506,N_13891,N_14657);
and U17507 (N_17507,N_13625,N_15286);
or U17508 (N_17508,N_13156,N_14265);
and U17509 (N_17509,N_13419,N_14918);
nand U17510 (N_17510,N_12679,N_12818);
xnor U17511 (N_17511,N_15303,N_14252);
nor U17512 (N_17512,N_13552,N_12505);
or U17513 (N_17513,N_13143,N_14351);
or U17514 (N_17514,N_14802,N_12676);
nor U17515 (N_17515,N_15369,N_13822);
or U17516 (N_17516,N_13027,N_15607);
nand U17517 (N_17517,N_14824,N_13678);
xnor U17518 (N_17518,N_13583,N_14602);
nand U17519 (N_17519,N_12565,N_14440);
nor U17520 (N_17520,N_14108,N_12913);
xor U17521 (N_17521,N_15259,N_13182);
nor U17522 (N_17522,N_13387,N_14587);
nor U17523 (N_17523,N_14068,N_14334);
nor U17524 (N_17524,N_15374,N_13708);
nand U17525 (N_17525,N_13344,N_12817);
nand U17526 (N_17526,N_12682,N_14847);
nand U17527 (N_17527,N_15433,N_13492);
or U17528 (N_17528,N_14842,N_13418);
xnor U17529 (N_17529,N_14831,N_14084);
nand U17530 (N_17530,N_13711,N_14332);
xnor U17531 (N_17531,N_15527,N_15093);
and U17532 (N_17532,N_12949,N_12796);
nand U17533 (N_17533,N_14157,N_13775);
nor U17534 (N_17534,N_13044,N_15253);
nand U17535 (N_17535,N_14635,N_14851);
nand U17536 (N_17536,N_14753,N_13528);
nand U17537 (N_17537,N_13688,N_13817);
or U17538 (N_17538,N_14377,N_14363);
nor U17539 (N_17539,N_14347,N_12583);
and U17540 (N_17540,N_12572,N_14256);
nor U17541 (N_17541,N_12970,N_12535);
nor U17542 (N_17542,N_12669,N_13865);
and U17543 (N_17543,N_15519,N_14540);
or U17544 (N_17544,N_13457,N_13524);
and U17545 (N_17545,N_14382,N_15470);
nor U17546 (N_17546,N_14045,N_13750);
nor U17547 (N_17547,N_14506,N_13814);
nor U17548 (N_17548,N_14361,N_14576);
and U17549 (N_17549,N_14599,N_13793);
or U17550 (N_17550,N_15410,N_13789);
nor U17551 (N_17551,N_13994,N_15457);
xor U17552 (N_17552,N_14486,N_14208);
and U17553 (N_17553,N_12958,N_13068);
nand U17554 (N_17554,N_13130,N_14382);
or U17555 (N_17555,N_13533,N_14143);
and U17556 (N_17556,N_13911,N_13830);
nor U17557 (N_17557,N_15266,N_13921);
xor U17558 (N_17558,N_12668,N_13028);
nand U17559 (N_17559,N_12784,N_13214);
nor U17560 (N_17560,N_15574,N_13368);
or U17561 (N_17561,N_14904,N_13389);
and U17562 (N_17562,N_14968,N_12971);
nor U17563 (N_17563,N_13115,N_14270);
nor U17564 (N_17564,N_13903,N_14686);
nor U17565 (N_17565,N_14317,N_13616);
or U17566 (N_17566,N_12683,N_15051);
nor U17567 (N_17567,N_15032,N_13118);
xnor U17568 (N_17568,N_13679,N_12864);
or U17569 (N_17569,N_14298,N_13560);
xnor U17570 (N_17570,N_14540,N_13038);
or U17571 (N_17571,N_13236,N_14394);
xnor U17572 (N_17572,N_13309,N_12564);
nor U17573 (N_17573,N_13259,N_14338);
xor U17574 (N_17574,N_15353,N_13239);
or U17575 (N_17575,N_13403,N_13125);
nand U17576 (N_17576,N_15278,N_13862);
nand U17577 (N_17577,N_13931,N_15601);
and U17578 (N_17578,N_12646,N_14880);
and U17579 (N_17579,N_14708,N_13823);
xnor U17580 (N_17580,N_15302,N_14555);
nand U17581 (N_17581,N_13475,N_12540);
nand U17582 (N_17582,N_14588,N_13703);
xor U17583 (N_17583,N_15226,N_14027);
nand U17584 (N_17584,N_13741,N_12827);
nor U17585 (N_17585,N_12537,N_13483);
nand U17586 (N_17586,N_12765,N_14337);
nor U17587 (N_17587,N_12848,N_12986);
xor U17588 (N_17588,N_13980,N_14351);
nand U17589 (N_17589,N_14378,N_14985);
nor U17590 (N_17590,N_12677,N_15109);
nand U17591 (N_17591,N_13472,N_15230);
or U17592 (N_17592,N_15208,N_14346);
and U17593 (N_17593,N_15597,N_14294);
nor U17594 (N_17594,N_13426,N_12790);
or U17595 (N_17595,N_15370,N_14327);
xnor U17596 (N_17596,N_14841,N_14123);
xor U17597 (N_17597,N_14622,N_14377);
xnor U17598 (N_17598,N_14329,N_13402);
and U17599 (N_17599,N_12645,N_13654);
nand U17600 (N_17600,N_14867,N_13319);
nor U17601 (N_17601,N_14028,N_12751);
xnor U17602 (N_17602,N_12730,N_12905);
and U17603 (N_17603,N_12736,N_15473);
or U17604 (N_17604,N_14547,N_15001);
nor U17605 (N_17605,N_15285,N_14809);
nor U17606 (N_17606,N_12768,N_14417);
nand U17607 (N_17607,N_14542,N_15607);
or U17608 (N_17608,N_13200,N_14381);
or U17609 (N_17609,N_13972,N_14876);
or U17610 (N_17610,N_15246,N_13468);
nor U17611 (N_17611,N_13587,N_13756);
and U17612 (N_17612,N_13780,N_12768);
nand U17613 (N_17613,N_15336,N_13305);
nand U17614 (N_17614,N_14227,N_14782);
xnor U17615 (N_17615,N_14715,N_12765);
and U17616 (N_17616,N_13069,N_13426);
xor U17617 (N_17617,N_14202,N_12766);
xnor U17618 (N_17618,N_13153,N_15119);
xnor U17619 (N_17619,N_13448,N_12511);
or U17620 (N_17620,N_15610,N_12518);
xor U17621 (N_17621,N_12873,N_15531);
and U17622 (N_17622,N_13420,N_13592);
or U17623 (N_17623,N_14367,N_12560);
xor U17624 (N_17624,N_13643,N_12795);
xnor U17625 (N_17625,N_13974,N_12838);
xor U17626 (N_17626,N_15095,N_14466);
xor U17627 (N_17627,N_14517,N_14671);
or U17628 (N_17628,N_14642,N_13021);
nor U17629 (N_17629,N_13748,N_14850);
xor U17630 (N_17630,N_14558,N_14710);
or U17631 (N_17631,N_13309,N_15596);
and U17632 (N_17632,N_13304,N_13569);
and U17633 (N_17633,N_15604,N_13031);
nand U17634 (N_17634,N_15163,N_13902);
nand U17635 (N_17635,N_15174,N_12507);
nand U17636 (N_17636,N_14784,N_13943);
and U17637 (N_17637,N_14856,N_14232);
nor U17638 (N_17638,N_14890,N_13315);
nor U17639 (N_17639,N_13527,N_14215);
and U17640 (N_17640,N_14215,N_14632);
and U17641 (N_17641,N_12731,N_12804);
xor U17642 (N_17642,N_14287,N_14352);
or U17643 (N_17643,N_14545,N_15229);
and U17644 (N_17644,N_12951,N_12515);
nand U17645 (N_17645,N_14004,N_14622);
nand U17646 (N_17646,N_14697,N_14746);
xnor U17647 (N_17647,N_14489,N_15459);
nand U17648 (N_17648,N_15349,N_13951);
nor U17649 (N_17649,N_13135,N_13287);
nor U17650 (N_17650,N_15447,N_14987);
or U17651 (N_17651,N_13791,N_14639);
nor U17652 (N_17652,N_14040,N_13395);
nand U17653 (N_17653,N_12693,N_15488);
and U17654 (N_17654,N_13551,N_13227);
nand U17655 (N_17655,N_15101,N_15084);
and U17656 (N_17656,N_13021,N_12614);
nand U17657 (N_17657,N_14494,N_12774);
nand U17658 (N_17658,N_14620,N_13299);
nor U17659 (N_17659,N_14216,N_15006);
and U17660 (N_17660,N_14082,N_14656);
nand U17661 (N_17661,N_13263,N_13266);
xnor U17662 (N_17662,N_15085,N_14600);
xnor U17663 (N_17663,N_14785,N_13637);
and U17664 (N_17664,N_13205,N_14287);
or U17665 (N_17665,N_13858,N_15332);
and U17666 (N_17666,N_14021,N_14302);
xor U17667 (N_17667,N_15553,N_13116);
xor U17668 (N_17668,N_13205,N_14243);
and U17669 (N_17669,N_13767,N_15531);
xor U17670 (N_17670,N_14638,N_13973);
or U17671 (N_17671,N_12912,N_14618);
nand U17672 (N_17672,N_13686,N_13608);
or U17673 (N_17673,N_15069,N_12524);
nand U17674 (N_17674,N_14646,N_14910);
nor U17675 (N_17675,N_13951,N_15150);
or U17676 (N_17676,N_12513,N_15123);
xnor U17677 (N_17677,N_14956,N_12956);
nor U17678 (N_17678,N_14432,N_15147);
nand U17679 (N_17679,N_14538,N_14523);
or U17680 (N_17680,N_13159,N_14787);
nand U17681 (N_17681,N_12945,N_14584);
nand U17682 (N_17682,N_13299,N_13975);
nand U17683 (N_17683,N_13422,N_12870);
xnor U17684 (N_17684,N_13387,N_13244);
xnor U17685 (N_17685,N_14439,N_12945);
nand U17686 (N_17686,N_13247,N_14228);
or U17687 (N_17687,N_15560,N_14315);
xnor U17688 (N_17688,N_12544,N_14803);
nor U17689 (N_17689,N_15514,N_13903);
nand U17690 (N_17690,N_14538,N_14148);
xor U17691 (N_17691,N_14100,N_14555);
xnor U17692 (N_17692,N_13443,N_12730);
xor U17693 (N_17693,N_13608,N_15441);
nor U17694 (N_17694,N_14916,N_15406);
nand U17695 (N_17695,N_13957,N_14060);
xnor U17696 (N_17696,N_13159,N_14945);
nor U17697 (N_17697,N_13828,N_14764);
and U17698 (N_17698,N_14342,N_15406);
xnor U17699 (N_17699,N_14458,N_12916);
xor U17700 (N_17700,N_13696,N_14999);
xnor U17701 (N_17701,N_14085,N_14226);
nand U17702 (N_17702,N_13890,N_14776);
or U17703 (N_17703,N_12981,N_14476);
or U17704 (N_17704,N_13838,N_12964);
or U17705 (N_17705,N_14747,N_13709);
xor U17706 (N_17706,N_14804,N_12755);
xnor U17707 (N_17707,N_14829,N_14853);
and U17708 (N_17708,N_15209,N_14458);
and U17709 (N_17709,N_15286,N_13019);
or U17710 (N_17710,N_12556,N_12975);
xnor U17711 (N_17711,N_14665,N_13083);
or U17712 (N_17712,N_13296,N_13351);
nand U17713 (N_17713,N_15108,N_14595);
nor U17714 (N_17714,N_15466,N_12833);
and U17715 (N_17715,N_15566,N_13542);
xor U17716 (N_17716,N_14587,N_13866);
or U17717 (N_17717,N_13697,N_14519);
xor U17718 (N_17718,N_15178,N_13531);
or U17719 (N_17719,N_13663,N_12812);
nand U17720 (N_17720,N_14539,N_15492);
xnor U17721 (N_17721,N_13056,N_15409);
xnor U17722 (N_17722,N_14712,N_14343);
and U17723 (N_17723,N_12889,N_13459);
and U17724 (N_17724,N_12991,N_13673);
or U17725 (N_17725,N_14931,N_14810);
nor U17726 (N_17726,N_12696,N_13953);
nor U17727 (N_17727,N_15367,N_14675);
nand U17728 (N_17728,N_15013,N_13285);
xnor U17729 (N_17729,N_14202,N_14366);
xnor U17730 (N_17730,N_13502,N_14924);
or U17731 (N_17731,N_14656,N_14500);
xnor U17732 (N_17732,N_13563,N_15143);
nand U17733 (N_17733,N_14055,N_13975);
and U17734 (N_17734,N_13452,N_13399);
or U17735 (N_17735,N_15492,N_14743);
xor U17736 (N_17736,N_12714,N_12585);
nand U17737 (N_17737,N_13716,N_14812);
or U17738 (N_17738,N_13442,N_12795);
or U17739 (N_17739,N_14731,N_14607);
or U17740 (N_17740,N_13960,N_13964);
or U17741 (N_17741,N_14519,N_14508);
xnor U17742 (N_17742,N_14479,N_12772);
nand U17743 (N_17743,N_14994,N_13839);
and U17744 (N_17744,N_15416,N_15527);
nor U17745 (N_17745,N_15209,N_15555);
or U17746 (N_17746,N_13911,N_13218);
or U17747 (N_17747,N_14472,N_13537);
or U17748 (N_17748,N_14092,N_13857);
or U17749 (N_17749,N_12628,N_13325);
nand U17750 (N_17750,N_15231,N_14191);
nor U17751 (N_17751,N_15129,N_15188);
nor U17752 (N_17752,N_13372,N_13691);
nand U17753 (N_17753,N_15497,N_15095);
nor U17754 (N_17754,N_12562,N_15226);
xor U17755 (N_17755,N_15247,N_14636);
nor U17756 (N_17756,N_15120,N_14471);
nor U17757 (N_17757,N_13597,N_13750);
nor U17758 (N_17758,N_14169,N_15349);
or U17759 (N_17759,N_13366,N_13642);
xnor U17760 (N_17760,N_13691,N_15048);
nor U17761 (N_17761,N_12947,N_14328);
nand U17762 (N_17762,N_15028,N_14139);
and U17763 (N_17763,N_14510,N_12837);
and U17764 (N_17764,N_13936,N_12909);
or U17765 (N_17765,N_12968,N_12771);
xor U17766 (N_17766,N_14544,N_15242);
or U17767 (N_17767,N_12873,N_13590);
xnor U17768 (N_17768,N_12864,N_13909);
and U17769 (N_17769,N_13828,N_14501);
nor U17770 (N_17770,N_13324,N_14159);
nor U17771 (N_17771,N_15215,N_14082);
xnor U17772 (N_17772,N_14490,N_15330);
and U17773 (N_17773,N_14539,N_14074);
xor U17774 (N_17774,N_14266,N_13957);
nand U17775 (N_17775,N_15288,N_12747);
and U17776 (N_17776,N_14255,N_12932);
or U17777 (N_17777,N_15323,N_13572);
or U17778 (N_17778,N_13263,N_14778);
xnor U17779 (N_17779,N_13704,N_12673);
or U17780 (N_17780,N_13401,N_15150);
nor U17781 (N_17781,N_14770,N_12681);
xor U17782 (N_17782,N_15388,N_15465);
and U17783 (N_17783,N_15489,N_15183);
or U17784 (N_17784,N_12667,N_13273);
and U17785 (N_17785,N_15395,N_14071);
or U17786 (N_17786,N_14004,N_15387);
and U17787 (N_17787,N_15219,N_13162);
nor U17788 (N_17788,N_15092,N_14649);
or U17789 (N_17789,N_13032,N_13546);
nor U17790 (N_17790,N_14547,N_15224);
nand U17791 (N_17791,N_12751,N_14564);
xnor U17792 (N_17792,N_15365,N_15167);
xor U17793 (N_17793,N_12784,N_15091);
or U17794 (N_17794,N_15535,N_14203);
and U17795 (N_17795,N_13552,N_13376);
nand U17796 (N_17796,N_14770,N_12537);
or U17797 (N_17797,N_14298,N_13566);
nand U17798 (N_17798,N_14898,N_14236);
xnor U17799 (N_17799,N_13221,N_14704);
and U17800 (N_17800,N_12572,N_12576);
xor U17801 (N_17801,N_15520,N_15604);
xor U17802 (N_17802,N_14758,N_14382);
and U17803 (N_17803,N_12679,N_15519);
or U17804 (N_17804,N_15139,N_13689);
and U17805 (N_17805,N_13430,N_13510);
or U17806 (N_17806,N_13397,N_12788);
and U17807 (N_17807,N_15487,N_13744);
xor U17808 (N_17808,N_12569,N_14421);
nor U17809 (N_17809,N_12756,N_12674);
and U17810 (N_17810,N_13300,N_13669);
nor U17811 (N_17811,N_13033,N_12691);
xor U17812 (N_17812,N_15249,N_13244);
nor U17813 (N_17813,N_14548,N_13040);
nand U17814 (N_17814,N_15172,N_15337);
and U17815 (N_17815,N_15207,N_14988);
nor U17816 (N_17816,N_12511,N_12708);
xnor U17817 (N_17817,N_15156,N_14145);
and U17818 (N_17818,N_14881,N_13095);
nor U17819 (N_17819,N_14111,N_14704);
and U17820 (N_17820,N_15058,N_13088);
or U17821 (N_17821,N_13832,N_13357);
nand U17822 (N_17822,N_14016,N_15276);
or U17823 (N_17823,N_12776,N_15280);
and U17824 (N_17824,N_13843,N_14587);
and U17825 (N_17825,N_13332,N_15378);
nand U17826 (N_17826,N_13713,N_15527);
or U17827 (N_17827,N_13087,N_13201);
nor U17828 (N_17828,N_14250,N_14908);
nand U17829 (N_17829,N_13177,N_13305);
and U17830 (N_17830,N_12933,N_13054);
nor U17831 (N_17831,N_14607,N_12829);
or U17832 (N_17832,N_14963,N_15559);
nand U17833 (N_17833,N_12807,N_15203);
and U17834 (N_17834,N_13666,N_14614);
xnor U17835 (N_17835,N_14102,N_14722);
or U17836 (N_17836,N_14102,N_14925);
xnor U17837 (N_17837,N_14745,N_13804);
nor U17838 (N_17838,N_13709,N_14407);
nand U17839 (N_17839,N_13407,N_12644);
and U17840 (N_17840,N_12567,N_14755);
or U17841 (N_17841,N_15524,N_14318);
nor U17842 (N_17842,N_15114,N_12765);
nand U17843 (N_17843,N_15539,N_14976);
nand U17844 (N_17844,N_14883,N_15433);
xor U17845 (N_17845,N_14851,N_15145);
nor U17846 (N_17846,N_13978,N_14228);
nand U17847 (N_17847,N_13235,N_15252);
nor U17848 (N_17848,N_15264,N_14953);
nor U17849 (N_17849,N_14434,N_13284);
or U17850 (N_17850,N_13105,N_13252);
xor U17851 (N_17851,N_13836,N_15356);
nand U17852 (N_17852,N_13613,N_14165);
or U17853 (N_17853,N_14729,N_14142);
xnor U17854 (N_17854,N_14915,N_13867);
nand U17855 (N_17855,N_13501,N_13869);
nor U17856 (N_17856,N_13929,N_15463);
xor U17857 (N_17857,N_14188,N_14056);
xnor U17858 (N_17858,N_15215,N_13368);
and U17859 (N_17859,N_14206,N_12713);
and U17860 (N_17860,N_14553,N_15483);
xnor U17861 (N_17861,N_13485,N_14260);
nand U17862 (N_17862,N_13331,N_14770);
and U17863 (N_17863,N_15301,N_15104);
xnor U17864 (N_17864,N_15581,N_14031);
nor U17865 (N_17865,N_15282,N_14380);
nor U17866 (N_17866,N_14814,N_12542);
nand U17867 (N_17867,N_15527,N_15565);
and U17868 (N_17868,N_14499,N_13724);
or U17869 (N_17869,N_12752,N_15301);
xor U17870 (N_17870,N_15351,N_14497);
xnor U17871 (N_17871,N_14277,N_13516);
nand U17872 (N_17872,N_14762,N_14912);
nor U17873 (N_17873,N_14673,N_12500);
or U17874 (N_17874,N_14259,N_15082);
xnor U17875 (N_17875,N_13982,N_14996);
and U17876 (N_17876,N_14263,N_14365);
nor U17877 (N_17877,N_12779,N_13074);
nand U17878 (N_17878,N_14666,N_13643);
nand U17879 (N_17879,N_15101,N_15474);
xor U17880 (N_17880,N_12642,N_14446);
xor U17881 (N_17881,N_14539,N_13522);
nand U17882 (N_17882,N_13616,N_15145);
and U17883 (N_17883,N_13473,N_12643);
nand U17884 (N_17884,N_14776,N_13184);
or U17885 (N_17885,N_13673,N_13668);
nand U17886 (N_17886,N_13873,N_13500);
xnor U17887 (N_17887,N_14650,N_15227);
nor U17888 (N_17888,N_15617,N_15620);
xor U17889 (N_17889,N_12622,N_15149);
nor U17890 (N_17890,N_13909,N_13724);
nor U17891 (N_17891,N_13357,N_15044);
nor U17892 (N_17892,N_15031,N_15002);
and U17893 (N_17893,N_14795,N_15044);
or U17894 (N_17894,N_14170,N_15071);
and U17895 (N_17895,N_13319,N_12666);
or U17896 (N_17896,N_13092,N_14417);
or U17897 (N_17897,N_14587,N_13736);
nor U17898 (N_17898,N_12684,N_13083);
nor U17899 (N_17899,N_12522,N_15179);
and U17900 (N_17900,N_14134,N_15261);
nor U17901 (N_17901,N_12761,N_15325);
or U17902 (N_17902,N_15268,N_13019);
xor U17903 (N_17903,N_13053,N_14359);
and U17904 (N_17904,N_13136,N_12784);
xnor U17905 (N_17905,N_15585,N_14396);
nor U17906 (N_17906,N_13039,N_13974);
xor U17907 (N_17907,N_15034,N_14975);
xor U17908 (N_17908,N_12637,N_13711);
or U17909 (N_17909,N_14330,N_15310);
or U17910 (N_17910,N_15387,N_15221);
and U17911 (N_17911,N_12993,N_13508);
and U17912 (N_17912,N_13417,N_15448);
and U17913 (N_17913,N_14972,N_12771);
and U17914 (N_17914,N_14156,N_13447);
and U17915 (N_17915,N_14499,N_15576);
nor U17916 (N_17916,N_13751,N_14570);
and U17917 (N_17917,N_14860,N_15265);
xor U17918 (N_17918,N_12649,N_14591);
or U17919 (N_17919,N_14667,N_15230);
nand U17920 (N_17920,N_14259,N_12880);
nand U17921 (N_17921,N_14631,N_13057);
and U17922 (N_17922,N_13964,N_13987);
and U17923 (N_17923,N_14373,N_13744);
nor U17924 (N_17924,N_13102,N_15264);
nor U17925 (N_17925,N_14621,N_13014);
xnor U17926 (N_17926,N_12922,N_15309);
xnor U17927 (N_17927,N_15086,N_12912);
xor U17928 (N_17928,N_15155,N_15460);
and U17929 (N_17929,N_15130,N_15237);
or U17930 (N_17930,N_14171,N_13658);
nand U17931 (N_17931,N_15555,N_13839);
or U17932 (N_17932,N_15365,N_15605);
xnor U17933 (N_17933,N_13369,N_12571);
nor U17934 (N_17934,N_12770,N_12542);
xnor U17935 (N_17935,N_12997,N_14927);
xnor U17936 (N_17936,N_14714,N_15414);
and U17937 (N_17937,N_13977,N_15438);
nand U17938 (N_17938,N_15413,N_13062);
nor U17939 (N_17939,N_13017,N_14788);
nand U17940 (N_17940,N_14106,N_15309);
nand U17941 (N_17941,N_13682,N_14543);
nor U17942 (N_17942,N_13139,N_15128);
and U17943 (N_17943,N_15384,N_13684);
and U17944 (N_17944,N_13940,N_14484);
or U17945 (N_17945,N_14892,N_15499);
and U17946 (N_17946,N_14044,N_14425);
nor U17947 (N_17947,N_13523,N_13111);
or U17948 (N_17948,N_14473,N_12878);
and U17949 (N_17949,N_14410,N_13179);
nand U17950 (N_17950,N_15615,N_14861);
or U17951 (N_17951,N_12917,N_14273);
and U17952 (N_17952,N_14864,N_14309);
and U17953 (N_17953,N_14473,N_15340);
or U17954 (N_17954,N_14173,N_13942);
xnor U17955 (N_17955,N_15079,N_14894);
nand U17956 (N_17956,N_13631,N_13402);
xor U17957 (N_17957,N_14177,N_14179);
nand U17958 (N_17958,N_15043,N_12502);
xnor U17959 (N_17959,N_12576,N_13494);
or U17960 (N_17960,N_14062,N_15455);
and U17961 (N_17961,N_14469,N_14345);
xnor U17962 (N_17962,N_12626,N_15373);
nor U17963 (N_17963,N_14070,N_13434);
or U17964 (N_17964,N_14273,N_15417);
xor U17965 (N_17965,N_13718,N_14214);
or U17966 (N_17966,N_12576,N_14220);
and U17967 (N_17967,N_14985,N_13176);
and U17968 (N_17968,N_12545,N_15149);
and U17969 (N_17969,N_14819,N_15041);
and U17970 (N_17970,N_15440,N_14919);
and U17971 (N_17971,N_13853,N_14226);
xnor U17972 (N_17972,N_12845,N_15112);
nor U17973 (N_17973,N_14406,N_12852);
xnor U17974 (N_17974,N_15565,N_14378);
nand U17975 (N_17975,N_13406,N_14448);
and U17976 (N_17976,N_12653,N_14126);
nor U17977 (N_17977,N_15199,N_12693);
nand U17978 (N_17978,N_14568,N_14445);
nand U17979 (N_17979,N_14368,N_14092);
xnor U17980 (N_17980,N_14458,N_15043);
nor U17981 (N_17981,N_13209,N_14396);
or U17982 (N_17982,N_14072,N_13619);
xnor U17983 (N_17983,N_15349,N_13194);
and U17984 (N_17984,N_15095,N_12792);
and U17985 (N_17985,N_14479,N_12899);
xor U17986 (N_17986,N_14081,N_12984);
nand U17987 (N_17987,N_12901,N_13518);
or U17988 (N_17988,N_15221,N_13045);
xor U17989 (N_17989,N_15276,N_13408);
or U17990 (N_17990,N_13282,N_13082);
nand U17991 (N_17991,N_13299,N_14525);
xor U17992 (N_17992,N_14666,N_14725);
or U17993 (N_17993,N_13495,N_13042);
and U17994 (N_17994,N_12659,N_13615);
nand U17995 (N_17995,N_15310,N_14856);
xor U17996 (N_17996,N_15219,N_14001);
or U17997 (N_17997,N_15316,N_14488);
nand U17998 (N_17998,N_12538,N_14371);
nand U17999 (N_17999,N_12508,N_15337);
or U18000 (N_18000,N_12845,N_13230);
nand U18001 (N_18001,N_13011,N_14246);
and U18002 (N_18002,N_12951,N_13778);
nor U18003 (N_18003,N_14044,N_13950);
nand U18004 (N_18004,N_13188,N_13155);
and U18005 (N_18005,N_13718,N_12586);
or U18006 (N_18006,N_14431,N_14585);
nand U18007 (N_18007,N_14848,N_13052);
nor U18008 (N_18008,N_12879,N_13935);
or U18009 (N_18009,N_15218,N_14449);
nor U18010 (N_18010,N_12955,N_13325);
and U18011 (N_18011,N_14000,N_14525);
and U18012 (N_18012,N_14106,N_15561);
xnor U18013 (N_18013,N_13845,N_12793);
xnor U18014 (N_18014,N_15306,N_15138);
xor U18015 (N_18015,N_14315,N_14056);
nor U18016 (N_18016,N_12961,N_13912);
nand U18017 (N_18017,N_15343,N_15415);
xor U18018 (N_18018,N_15074,N_12914);
xnor U18019 (N_18019,N_15473,N_14109);
xnor U18020 (N_18020,N_12512,N_15512);
or U18021 (N_18021,N_15452,N_14160);
and U18022 (N_18022,N_13869,N_13877);
xor U18023 (N_18023,N_14988,N_13560);
or U18024 (N_18024,N_14971,N_13222);
or U18025 (N_18025,N_13645,N_12948);
nand U18026 (N_18026,N_13643,N_15344);
nand U18027 (N_18027,N_14205,N_14856);
or U18028 (N_18028,N_15358,N_13001);
nor U18029 (N_18029,N_14367,N_12995);
nor U18030 (N_18030,N_12985,N_14867);
nand U18031 (N_18031,N_15060,N_15269);
and U18032 (N_18032,N_15435,N_14570);
nor U18033 (N_18033,N_15139,N_13346);
xor U18034 (N_18034,N_13285,N_14287);
xor U18035 (N_18035,N_13656,N_14242);
nand U18036 (N_18036,N_13116,N_14447);
and U18037 (N_18037,N_14905,N_14430);
and U18038 (N_18038,N_14635,N_13066);
and U18039 (N_18039,N_12593,N_14127);
nand U18040 (N_18040,N_15250,N_14006);
and U18041 (N_18041,N_12537,N_14436);
and U18042 (N_18042,N_15339,N_12877);
xnor U18043 (N_18043,N_13379,N_15436);
nand U18044 (N_18044,N_14140,N_14366);
or U18045 (N_18045,N_14378,N_14996);
nand U18046 (N_18046,N_15435,N_14114);
and U18047 (N_18047,N_13963,N_14553);
and U18048 (N_18048,N_12533,N_15404);
xnor U18049 (N_18049,N_13684,N_14751);
and U18050 (N_18050,N_15290,N_14764);
or U18051 (N_18051,N_14990,N_15225);
nand U18052 (N_18052,N_14606,N_14068);
nor U18053 (N_18053,N_13403,N_12867);
nand U18054 (N_18054,N_12563,N_15338);
nor U18055 (N_18055,N_12601,N_14117);
xor U18056 (N_18056,N_15216,N_15404);
xnor U18057 (N_18057,N_15622,N_13263);
and U18058 (N_18058,N_14704,N_13774);
and U18059 (N_18059,N_13906,N_14857);
nand U18060 (N_18060,N_14990,N_15286);
nor U18061 (N_18061,N_15537,N_14922);
and U18062 (N_18062,N_12784,N_15343);
nand U18063 (N_18063,N_13206,N_13670);
nor U18064 (N_18064,N_12985,N_14427);
and U18065 (N_18065,N_13494,N_13985);
xnor U18066 (N_18066,N_13434,N_13757);
or U18067 (N_18067,N_13735,N_15043);
nand U18068 (N_18068,N_12555,N_14631);
or U18069 (N_18069,N_15036,N_14588);
or U18070 (N_18070,N_14471,N_14075);
and U18071 (N_18071,N_13303,N_15559);
nand U18072 (N_18072,N_14113,N_12713);
nor U18073 (N_18073,N_14573,N_13688);
xnor U18074 (N_18074,N_14693,N_13187);
and U18075 (N_18075,N_14058,N_12708);
and U18076 (N_18076,N_13124,N_14786);
nand U18077 (N_18077,N_13909,N_14414);
and U18078 (N_18078,N_13008,N_15341);
nand U18079 (N_18079,N_12562,N_14795);
xnor U18080 (N_18080,N_13531,N_14622);
xor U18081 (N_18081,N_14642,N_13563);
nor U18082 (N_18082,N_14580,N_13812);
xor U18083 (N_18083,N_14139,N_14869);
or U18084 (N_18084,N_12646,N_14868);
nand U18085 (N_18085,N_14100,N_13754);
and U18086 (N_18086,N_13861,N_14131);
and U18087 (N_18087,N_13021,N_12913);
and U18088 (N_18088,N_15298,N_15022);
and U18089 (N_18089,N_13331,N_13110);
nand U18090 (N_18090,N_13045,N_14745);
nor U18091 (N_18091,N_12973,N_13458);
or U18092 (N_18092,N_15291,N_12791);
nor U18093 (N_18093,N_14091,N_14591);
or U18094 (N_18094,N_13610,N_12796);
nand U18095 (N_18095,N_15245,N_12900);
and U18096 (N_18096,N_14787,N_14830);
xnor U18097 (N_18097,N_14528,N_15558);
nor U18098 (N_18098,N_12727,N_13964);
xor U18099 (N_18099,N_12685,N_14957);
and U18100 (N_18100,N_13130,N_14244);
or U18101 (N_18101,N_14137,N_15248);
and U18102 (N_18102,N_14768,N_14819);
xnor U18103 (N_18103,N_13302,N_14827);
and U18104 (N_18104,N_13977,N_14116);
and U18105 (N_18105,N_14852,N_14794);
nand U18106 (N_18106,N_14073,N_14706);
nor U18107 (N_18107,N_13360,N_13827);
nor U18108 (N_18108,N_13184,N_13240);
and U18109 (N_18109,N_13320,N_13096);
nand U18110 (N_18110,N_13426,N_15216);
xor U18111 (N_18111,N_14439,N_13683);
xnor U18112 (N_18112,N_12972,N_13376);
xor U18113 (N_18113,N_12852,N_14136);
xnor U18114 (N_18114,N_13058,N_13753);
and U18115 (N_18115,N_13560,N_13488);
nor U18116 (N_18116,N_14069,N_14795);
nor U18117 (N_18117,N_13278,N_13016);
xnor U18118 (N_18118,N_15025,N_12653);
xor U18119 (N_18119,N_13154,N_14515);
or U18120 (N_18120,N_15261,N_14869);
nand U18121 (N_18121,N_13949,N_12695);
or U18122 (N_18122,N_13885,N_13708);
xnor U18123 (N_18123,N_15404,N_15262);
and U18124 (N_18124,N_13719,N_13590);
or U18125 (N_18125,N_13187,N_14564);
nand U18126 (N_18126,N_13941,N_14399);
or U18127 (N_18127,N_14822,N_13610);
and U18128 (N_18128,N_13022,N_14904);
or U18129 (N_18129,N_13131,N_14426);
or U18130 (N_18130,N_14293,N_14039);
and U18131 (N_18131,N_14095,N_12753);
or U18132 (N_18132,N_13203,N_13913);
xnor U18133 (N_18133,N_12669,N_13180);
nor U18134 (N_18134,N_15428,N_13269);
xnor U18135 (N_18135,N_13556,N_13266);
or U18136 (N_18136,N_14722,N_15609);
nand U18137 (N_18137,N_14915,N_15114);
xor U18138 (N_18138,N_13938,N_15343);
and U18139 (N_18139,N_14977,N_14167);
nor U18140 (N_18140,N_13645,N_13117);
xnor U18141 (N_18141,N_13796,N_14831);
nor U18142 (N_18142,N_12697,N_15274);
nor U18143 (N_18143,N_13777,N_14677);
nor U18144 (N_18144,N_14177,N_13005);
nor U18145 (N_18145,N_14915,N_13856);
nor U18146 (N_18146,N_13710,N_14036);
nand U18147 (N_18147,N_14737,N_14116);
nand U18148 (N_18148,N_13767,N_15037);
or U18149 (N_18149,N_14452,N_15592);
and U18150 (N_18150,N_15252,N_14655);
and U18151 (N_18151,N_13203,N_14496);
nor U18152 (N_18152,N_14189,N_15266);
xor U18153 (N_18153,N_13906,N_15089);
and U18154 (N_18154,N_13569,N_15566);
or U18155 (N_18155,N_15292,N_14226);
or U18156 (N_18156,N_14647,N_15116);
xor U18157 (N_18157,N_15177,N_15372);
xor U18158 (N_18158,N_15390,N_13046);
xor U18159 (N_18159,N_15318,N_14727);
nor U18160 (N_18160,N_12952,N_15356);
nor U18161 (N_18161,N_12858,N_15205);
nor U18162 (N_18162,N_13638,N_14584);
and U18163 (N_18163,N_14364,N_12526);
and U18164 (N_18164,N_13986,N_13440);
or U18165 (N_18165,N_12817,N_12803);
xnor U18166 (N_18166,N_14882,N_13343);
and U18167 (N_18167,N_12951,N_12775);
nor U18168 (N_18168,N_14593,N_15036);
or U18169 (N_18169,N_13662,N_14812);
xnor U18170 (N_18170,N_13094,N_14304);
nor U18171 (N_18171,N_12759,N_15013);
and U18172 (N_18172,N_13290,N_12873);
and U18173 (N_18173,N_15271,N_14863);
xor U18174 (N_18174,N_12735,N_14088);
and U18175 (N_18175,N_15059,N_15017);
xnor U18176 (N_18176,N_14440,N_13913);
nor U18177 (N_18177,N_13529,N_14355);
nand U18178 (N_18178,N_14898,N_13034);
nor U18179 (N_18179,N_13526,N_15338);
and U18180 (N_18180,N_13421,N_12673);
nor U18181 (N_18181,N_14199,N_13556);
or U18182 (N_18182,N_14475,N_13510);
xor U18183 (N_18183,N_14759,N_13986);
and U18184 (N_18184,N_15277,N_14747);
nand U18185 (N_18185,N_13959,N_12845);
or U18186 (N_18186,N_12845,N_13124);
nor U18187 (N_18187,N_14112,N_12694);
nor U18188 (N_18188,N_15623,N_15087);
and U18189 (N_18189,N_15240,N_15393);
or U18190 (N_18190,N_12554,N_13639);
nand U18191 (N_18191,N_15116,N_15436);
nand U18192 (N_18192,N_15267,N_13722);
and U18193 (N_18193,N_12568,N_13221);
and U18194 (N_18194,N_12747,N_14075);
nor U18195 (N_18195,N_12797,N_14642);
nand U18196 (N_18196,N_12728,N_13093);
xor U18197 (N_18197,N_13825,N_13972);
xnor U18198 (N_18198,N_12884,N_12702);
or U18199 (N_18199,N_13285,N_13001);
nand U18200 (N_18200,N_12875,N_12619);
and U18201 (N_18201,N_15042,N_14512);
nor U18202 (N_18202,N_12880,N_12823);
xor U18203 (N_18203,N_12663,N_13665);
xor U18204 (N_18204,N_15528,N_13444);
and U18205 (N_18205,N_12759,N_13032);
xnor U18206 (N_18206,N_15432,N_14828);
or U18207 (N_18207,N_14176,N_12905);
nor U18208 (N_18208,N_13827,N_13700);
xnor U18209 (N_18209,N_13564,N_13318);
and U18210 (N_18210,N_14163,N_12524);
xnor U18211 (N_18211,N_15265,N_14045);
nor U18212 (N_18212,N_13590,N_13496);
and U18213 (N_18213,N_14299,N_14901);
and U18214 (N_18214,N_15064,N_13877);
or U18215 (N_18215,N_13996,N_12943);
nor U18216 (N_18216,N_12720,N_12981);
and U18217 (N_18217,N_15397,N_13065);
xor U18218 (N_18218,N_12752,N_14189);
or U18219 (N_18219,N_12583,N_14616);
nor U18220 (N_18220,N_12928,N_13016);
and U18221 (N_18221,N_13231,N_13017);
xnor U18222 (N_18222,N_14511,N_15163);
nor U18223 (N_18223,N_12558,N_15349);
or U18224 (N_18224,N_13666,N_15189);
xnor U18225 (N_18225,N_15149,N_15605);
nor U18226 (N_18226,N_13484,N_14223);
nor U18227 (N_18227,N_15280,N_13195);
nor U18228 (N_18228,N_13599,N_13614);
xnor U18229 (N_18229,N_14073,N_12919);
and U18230 (N_18230,N_14459,N_13917);
or U18231 (N_18231,N_13451,N_13595);
nor U18232 (N_18232,N_14142,N_14429);
nor U18233 (N_18233,N_13628,N_14022);
and U18234 (N_18234,N_15066,N_15093);
and U18235 (N_18235,N_14854,N_14095);
nand U18236 (N_18236,N_13914,N_13653);
and U18237 (N_18237,N_13274,N_13596);
and U18238 (N_18238,N_13907,N_13763);
or U18239 (N_18239,N_12799,N_15450);
xnor U18240 (N_18240,N_13883,N_15560);
nor U18241 (N_18241,N_14787,N_14098);
xor U18242 (N_18242,N_12849,N_13766);
xnor U18243 (N_18243,N_14484,N_14264);
and U18244 (N_18244,N_15391,N_12751);
and U18245 (N_18245,N_14129,N_13991);
xor U18246 (N_18246,N_12716,N_15478);
xor U18247 (N_18247,N_15064,N_15332);
and U18248 (N_18248,N_14794,N_14875);
xor U18249 (N_18249,N_13528,N_13241);
nand U18250 (N_18250,N_14514,N_14660);
and U18251 (N_18251,N_13501,N_13346);
nor U18252 (N_18252,N_14830,N_14334);
xnor U18253 (N_18253,N_14963,N_13192);
nor U18254 (N_18254,N_15377,N_13210);
and U18255 (N_18255,N_14094,N_13952);
and U18256 (N_18256,N_13773,N_15372);
nand U18257 (N_18257,N_13503,N_13043);
nor U18258 (N_18258,N_14805,N_14131);
or U18259 (N_18259,N_13033,N_15385);
nor U18260 (N_18260,N_14056,N_14115);
xor U18261 (N_18261,N_13327,N_15030);
xnor U18262 (N_18262,N_13930,N_13484);
xor U18263 (N_18263,N_12855,N_15563);
or U18264 (N_18264,N_14389,N_13144);
or U18265 (N_18265,N_14068,N_13823);
nand U18266 (N_18266,N_15371,N_13069);
or U18267 (N_18267,N_15412,N_12734);
nor U18268 (N_18268,N_14575,N_13683);
nor U18269 (N_18269,N_14954,N_13603);
and U18270 (N_18270,N_13920,N_14485);
and U18271 (N_18271,N_14476,N_15265);
or U18272 (N_18272,N_13658,N_15425);
and U18273 (N_18273,N_12859,N_13734);
and U18274 (N_18274,N_14135,N_14430);
nand U18275 (N_18275,N_15267,N_14467);
xor U18276 (N_18276,N_13765,N_15518);
and U18277 (N_18277,N_12880,N_15079);
nor U18278 (N_18278,N_13583,N_13157);
or U18279 (N_18279,N_14224,N_14131);
and U18280 (N_18280,N_13857,N_14193);
and U18281 (N_18281,N_15305,N_14723);
and U18282 (N_18282,N_15051,N_13158);
nand U18283 (N_18283,N_14729,N_14346);
nor U18284 (N_18284,N_13899,N_12849);
and U18285 (N_18285,N_13133,N_13569);
and U18286 (N_18286,N_13996,N_13422);
xor U18287 (N_18287,N_14608,N_15563);
and U18288 (N_18288,N_14627,N_14526);
or U18289 (N_18289,N_14599,N_13107);
xor U18290 (N_18290,N_15120,N_15241);
nand U18291 (N_18291,N_14890,N_14102);
xnor U18292 (N_18292,N_14232,N_13473);
xor U18293 (N_18293,N_13796,N_14478);
and U18294 (N_18294,N_15410,N_15553);
or U18295 (N_18295,N_13441,N_12502);
nand U18296 (N_18296,N_13845,N_13827);
nor U18297 (N_18297,N_15460,N_13663);
xnor U18298 (N_18298,N_15029,N_12618);
or U18299 (N_18299,N_12862,N_15371);
nor U18300 (N_18300,N_15396,N_12867);
nor U18301 (N_18301,N_15620,N_13359);
nor U18302 (N_18302,N_15030,N_13841);
xor U18303 (N_18303,N_14879,N_14364);
xor U18304 (N_18304,N_14151,N_13845);
xor U18305 (N_18305,N_13041,N_13399);
nand U18306 (N_18306,N_13622,N_13179);
nor U18307 (N_18307,N_12707,N_13084);
or U18308 (N_18308,N_13217,N_14653);
or U18309 (N_18309,N_12929,N_14182);
nor U18310 (N_18310,N_14049,N_14531);
nand U18311 (N_18311,N_15209,N_14756);
xnor U18312 (N_18312,N_14366,N_14512);
xnor U18313 (N_18313,N_15100,N_13896);
nand U18314 (N_18314,N_14074,N_13116);
nor U18315 (N_18315,N_12659,N_15435);
nand U18316 (N_18316,N_14687,N_15139);
nand U18317 (N_18317,N_14201,N_14403);
nand U18318 (N_18318,N_13350,N_12980);
xor U18319 (N_18319,N_12707,N_14386);
and U18320 (N_18320,N_12895,N_14610);
nor U18321 (N_18321,N_13780,N_13253);
nand U18322 (N_18322,N_13048,N_15103);
or U18323 (N_18323,N_12630,N_13452);
nor U18324 (N_18324,N_12932,N_14511);
and U18325 (N_18325,N_14534,N_12797);
nor U18326 (N_18326,N_12792,N_12773);
and U18327 (N_18327,N_15143,N_13875);
or U18328 (N_18328,N_15554,N_13097);
nor U18329 (N_18329,N_14225,N_15497);
and U18330 (N_18330,N_14952,N_12546);
nand U18331 (N_18331,N_13380,N_14802);
nor U18332 (N_18332,N_12787,N_12737);
xnor U18333 (N_18333,N_12827,N_14938);
nor U18334 (N_18334,N_14009,N_14996);
and U18335 (N_18335,N_13741,N_14861);
nand U18336 (N_18336,N_13749,N_12653);
nor U18337 (N_18337,N_13418,N_15178);
or U18338 (N_18338,N_13737,N_15364);
xnor U18339 (N_18339,N_13234,N_15090);
or U18340 (N_18340,N_14260,N_15512);
nor U18341 (N_18341,N_13717,N_13990);
nor U18342 (N_18342,N_14347,N_13209);
xor U18343 (N_18343,N_15413,N_13008);
xnor U18344 (N_18344,N_14137,N_14313);
nor U18345 (N_18345,N_12539,N_12990);
or U18346 (N_18346,N_15409,N_12633);
or U18347 (N_18347,N_13949,N_15329);
or U18348 (N_18348,N_12536,N_14501);
and U18349 (N_18349,N_12694,N_13673);
nor U18350 (N_18350,N_14471,N_13023);
nor U18351 (N_18351,N_15555,N_12804);
nor U18352 (N_18352,N_12802,N_14803);
and U18353 (N_18353,N_12886,N_15271);
nor U18354 (N_18354,N_13692,N_14620);
or U18355 (N_18355,N_13917,N_12720);
nand U18356 (N_18356,N_15218,N_12751);
xor U18357 (N_18357,N_14524,N_14536);
nand U18358 (N_18358,N_13164,N_14735);
and U18359 (N_18359,N_14899,N_13333);
or U18360 (N_18360,N_14411,N_14390);
or U18361 (N_18361,N_15344,N_15385);
or U18362 (N_18362,N_14488,N_13845);
xnor U18363 (N_18363,N_15616,N_15533);
nand U18364 (N_18364,N_15095,N_13714);
or U18365 (N_18365,N_13227,N_14622);
xor U18366 (N_18366,N_14929,N_12553);
xnor U18367 (N_18367,N_14518,N_15315);
nor U18368 (N_18368,N_13323,N_13241);
and U18369 (N_18369,N_12674,N_13527);
and U18370 (N_18370,N_15141,N_15098);
nor U18371 (N_18371,N_13135,N_15437);
or U18372 (N_18372,N_12690,N_13605);
or U18373 (N_18373,N_14074,N_13500);
nor U18374 (N_18374,N_15246,N_14619);
nand U18375 (N_18375,N_14209,N_15049);
or U18376 (N_18376,N_14999,N_13680);
or U18377 (N_18377,N_12650,N_15597);
nor U18378 (N_18378,N_15462,N_12511);
nor U18379 (N_18379,N_12868,N_14473);
xnor U18380 (N_18380,N_12772,N_12609);
and U18381 (N_18381,N_15467,N_12920);
xnor U18382 (N_18382,N_12815,N_14734);
or U18383 (N_18383,N_14447,N_12794);
nor U18384 (N_18384,N_15152,N_13354);
nand U18385 (N_18385,N_14799,N_15555);
xnor U18386 (N_18386,N_13271,N_12925);
nor U18387 (N_18387,N_14875,N_14940);
or U18388 (N_18388,N_13901,N_13704);
xnor U18389 (N_18389,N_13824,N_13263);
nor U18390 (N_18390,N_12856,N_13184);
or U18391 (N_18391,N_15104,N_14221);
xor U18392 (N_18392,N_15592,N_14639);
xnor U18393 (N_18393,N_13663,N_13803);
nor U18394 (N_18394,N_15555,N_15224);
nor U18395 (N_18395,N_13373,N_13678);
nor U18396 (N_18396,N_14849,N_13997);
nor U18397 (N_18397,N_14402,N_12577);
and U18398 (N_18398,N_14443,N_13772);
nor U18399 (N_18399,N_15310,N_14610);
nand U18400 (N_18400,N_15073,N_14441);
nand U18401 (N_18401,N_13022,N_14786);
and U18402 (N_18402,N_15162,N_14526);
or U18403 (N_18403,N_13984,N_15314);
and U18404 (N_18404,N_15398,N_14210);
and U18405 (N_18405,N_12871,N_13869);
or U18406 (N_18406,N_14900,N_13930);
xnor U18407 (N_18407,N_15427,N_13225);
nand U18408 (N_18408,N_15248,N_15452);
nor U18409 (N_18409,N_14150,N_14640);
nand U18410 (N_18410,N_13648,N_13439);
and U18411 (N_18411,N_15129,N_14973);
nor U18412 (N_18412,N_15208,N_15067);
nor U18413 (N_18413,N_12755,N_14393);
or U18414 (N_18414,N_13249,N_12705);
nand U18415 (N_18415,N_14301,N_13305);
nor U18416 (N_18416,N_13034,N_12533);
and U18417 (N_18417,N_13201,N_14763);
nor U18418 (N_18418,N_14529,N_12624);
nor U18419 (N_18419,N_12984,N_13756);
nor U18420 (N_18420,N_12811,N_13028);
or U18421 (N_18421,N_14833,N_15078);
nor U18422 (N_18422,N_14540,N_12844);
and U18423 (N_18423,N_13007,N_15079);
nand U18424 (N_18424,N_14680,N_13705);
or U18425 (N_18425,N_13868,N_14585);
xor U18426 (N_18426,N_14768,N_13468);
or U18427 (N_18427,N_14086,N_12517);
nand U18428 (N_18428,N_13248,N_12564);
nor U18429 (N_18429,N_12658,N_15169);
or U18430 (N_18430,N_15351,N_15188);
nand U18431 (N_18431,N_13862,N_13261);
or U18432 (N_18432,N_13202,N_15606);
nand U18433 (N_18433,N_14741,N_13719);
xnor U18434 (N_18434,N_13341,N_13393);
or U18435 (N_18435,N_14959,N_12891);
xor U18436 (N_18436,N_13510,N_13895);
xnor U18437 (N_18437,N_12541,N_15506);
nor U18438 (N_18438,N_14528,N_15522);
or U18439 (N_18439,N_12848,N_15320);
and U18440 (N_18440,N_13087,N_14526);
nor U18441 (N_18441,N_14440,N_12741);
xor U18442 (N_18442,N_14692,N_14114);
and U18443 (N_18443,N_14321,N_14085);
nand U18444 (N_18444,N_14185,N_14804);
xnor U18445 (N_18445,N_12769,N_14152);
or U18446 (N_18446,N_14052,N_13637);
or U18447 (N_18447,N_15127,N_13560);
or U18448 (N_18448,N_15358,N_14861);
and U18449 (N_18449,N_13746,N_14112);
nor U18450 (N_18450,N_13005,N_14764);
xnor U18451 (N_18451,N_14083,N_13940);
xnor U18452 (N_18452,N_14397,N_15082);
nand U18453 (N_18453,N_15531,N_14771);
nor U18454 (N_18454,N_13357,N_13001);
xor U18455 (N_18455,N_13535,N_13097);
and U18456 (N_18456,N_13886,N_13577);
and U18457 (N_18457,N_15422,N_13303);
xnor U18458 (N_18458,N_13836,N_15038);
nand U18459 (N_18459,N_13852,N_14026);
nor U18460 (N_18460,N_13879,N_15010);
nor U18461 (N_18461,N_13882,N_14069);
nand U18462 (N_18462,N_14237,N_14561);
xor U18463 (N_18463,N_12875,N_12516);
xnor U18464 (N_18464,N_13313,N_13040);
and U18465 (N_18465,N_15305,N_15284);
nand U18466 (N_18466,N_15083,N_13079);
xnor U18467 (N_18467,N_13055,N_14412);
nor U18468 (N_18468,N_13584,N_13221);
xnor U18469 (N_18469,N_14117,N_14938);
nand U18470 (N_18470,N_14428,N_14128);
or U18471 (N_18471,N_14837,N_13431);
and U18472 (N_18472,N_13964,N_15262);
xor U18473 (N_18473,N_15377,N_15469);
and U18474 (N_18474,N_14765,N_13389);
xnor U18475 (N_18475,N_12910,N_12977);
nor U18476 (N_18476,N_13650,N_12706);
or U18477 (N_18477,N_14922,N_15299);
nand U18478 (N_18478,N_14127,N_12545);
or U18479 (N_18479,N_15417,N_15576);
and U18480 (N_18480,N_12520,N_15058);
or U18481 (N_18481,N_13193,N_12704);
and U18482 (N_18482,N_13657,N_15381);
xnor U18483 (N_18483,N_13360,N_14372);
nand U18484 (N_18484,N_15330,N_15227);
nor U18485 (N_18485,N_13907,N_13808);
and U18486 (N_18486,N_12848,N_15228);
or U18487 (N_18487,N_13709,N_14648);
and U18488 (N_18488,N_13150,N_12989);
and U18489 (N_18489,N_12589,N_13569);
and U18490 (N_18490,N_13670,N_12676);
nor U18491 (N_18491,N_15186,N_13612);
xor U18492 (N_18492,N_15094,N_13507);
xnor U18493 (N_18493,N_12945,N_14386);
and U18494 (N_18494,N_14500,N_14249);
nor U18495 (N_18495,N_14573,N_13492);
nand U18496 (N_18496,N_13036,N_15328);
xor U18497 (N_18497,N_14505,N_13575);
and U18498 (N_18498,N_14828,N_13414);
or U18499 (N_18499,N_15098,N_13860);
or U18500 (N_18500,N_14344,N_13907);
or U18501 (N_18501,N_14944,N_14568);
or U18502 (N_18502,N_13638,N_14160);
nand U18503 (N_18503,N_13206,N_15592);
or U18504 (N_18504,N_13676,N_14257);
nor U18505 (N_18505,N_12890,N_13115);
nand U18506 (N_18506,N_13661,N_12967);
nand U18507 (N_18507,N_15057,N_14653);
and U18508 (N_18508,N_14419,N_14410);
nand U18509 (N_18509,N_13557,N_14220);
nor U18510 (N_18510,N_13318,N_14252);
nand U18511 (N_18511,N_13944,N_15189);
and U18512 (N_18512,N_12565,N_13898);
xor U18513 (N_18513,N_12950,N_14879);
xnor U18514 (N_18514,N_13524,N_14866);
nand U18515 (N_18515,N_15450,N_13706);
and U18516 (N_18516,N_12554,N_15068);
and U18517 (N_18517,N_13251,N_15588);
or U18518 (N_18518,N_14511,N_14759);
xnor U18519 (N_18519,N_13929,N_13137);
nor U18520 (N_18520,N_13310,N_12549);
xnor U18521 (N_18521,N_14426,N_15596);
xnor U18522 (N_18522,N_14913,N_15609);
nand U18523 (N_18523,N_13869,N_13184);
nor U18524 (N_18524,N_14848,N_14184);
and U18525 (N_18525,N_13283,N_12985);
and U18526 (N_18526,N_12971,N_15613);
or U18527 (N_18527,N_15265,N_14107);
and U18528 (N_18528,N_14774,N_15060);
or U18529 (N_18529,N_13780,N_14772);
nor U18530 (N_18530,N_12918,N_12860);
nor U18531 (N_18531,N_14440,N_12736);
or U18532 (N_18532,N_12862,N_14186);
and U18533 (N_18533,N_13471,N_14303);
nor U18534 (N_18534,N_13890,N_13655);
nor U18535 (N_18535,N_14399,N_12698);
or U18536 (N_18536,N_15196,N_12750);
or U18537 (N_18537,N_13845,N_13586);
nand U18538 (N_18538,N_12838,N_13832);
and U18539 (N_18539,N_13769,N_14653);
nor U18540 (N_18540,N_13196,N_15115);
nand U18541 (N_18541,N_14501,N_14107);
xor U18542 (N_18542,N_13162,N_12984);
nor U18543 (N_18543,N_13274,N_14837);
and U18544 (N_18544,N_13007,N_15352);
nor U18545 (N_18545,N_14794,N_13608);
or U18546 (N_18546,N_14693,N_13958);
and U18547 (N_18547,N_14206,N_12517);
and U18548 (N_18548,N_15065,N_15464);
xor U18549 (N_18549,N_13550,N_13800);
and U18550 (N_18550,N_13283,N_13678);
and U18551 (N_18551,N_14956,N_14771);
nand U18552 (N_18552,N_14960,N_15554);
nand U18553 (N_18553,N_15268,N_13853);
nor U18554 (N_18554,N_13811,N_14619);
and U18555 (N_18555,N_12851,N_14618);
or U18556 (N_18556,N_13070,N_14500);
xnor U18557 (N_18557,N_13458,N_14276);
nor U18558 (N_18558,N_13815,N_12557);
xnor U18559 (N_18559,N_14381,N_13810);
nand U18560 (N_18560,N_15171,N_13383);
nor U18561 (N_18561,N_12583,N_13309);
or U18562 (N_18562,N_15000,N_13665);
and U18563 (N_18563,N_13209,N_12641);
or U18564 (N_18564,N_14717,N_13497);
and U18565 (N_18565,N_13655,N_14463);
and U18566 (N_18566,N_14813,N_15348);
xor U18567 (N_18567,N_13709,N_14515);
xor U18568 (N_18568,N_14483,N_12774);
xnor U18569 (N_18569,N_13178,N_14151);
xnor U18570 (N_18570,N_12554,N_12568);
nor U18571 (N_18571,N_15443,N_14387);
nor U18572 (N_18572,N_13640,N_12559);
xnor U18573 (N_18573,N_14226,N_15130);
xor U18574 (N_18574,N_14747,N_13516);
nand U18575 (N_18575,N_12870,N_13956);
nor U18576 (N_18576,N_14754,N_14739);
or U18577 (N_18577,N_14137,N_13819);
nand U18578 (N_18578,N_13810,N_15564);
nand U18579 (N_18579,N_14590,N_13762);
or U18580 (N_18580,N_13585,N_12544);
and U18581 (N_18581,N_13932,N_13909);
xnor U18582 (N_18582,N_15508,N_14825);
and U18583 (N_18583,N_15389,N_13155);
nor U18584 (N_18584,N_14991,N_13943);
nand U18585 (N_18585,N_13884,N_13629);
xnor U18586 (N_18586,N_14770,N_13538);
nor U18587 (N_18587,N_15087,N_15006);
nor U18588 (N_18588,N_13720,N_14266);
xnor U18589 (N_18589,N_15425,N_13458);
xor U18590 (N_18590,N_15546,N_15394);
nand U18591 (N_18591,N_13974,N_15385);
or U18592 (N_18592,N_14816,N_15247);
xnor U18593 (N_18593,N_13963,N_15142);
nand U18594 (N_18594,N_13810,N_15212);
and U18595 (N_18595,N_14388,N_15352);
xor U18596 (N_18596,N_14360,N_13595);
and U18597 (N_18597,N_14796,N_14813);
nor U18598 (N_18598,N_12770,N_12775);
and U18599 (N_18599,N_13931,N_13750);
nor U18600 (N_18600,N_12725,N_13402);
or U18601 (N_18601,N_15060,N_15491);
nor U18602 (N_18602,N_13649,N_13071);
or U18603 (N_18603,N_14938,N_12929);
and U18604 (N_18604,N_13531,N_13332);
nand U18605 (N_18605,N_13878,N_12615);
nor U18606 (N_18606,N_13276,N_15598);
xnor U18607 (N_18607,N_13611,N_12716);
xor U18608 (N_18608,N_13189,N_14094);
nand U18609 (N_18609,N_13593,N_14038);
and U18610 (N_18610,N_13464,N_13284);
nand U18611 (N_18611,N_15496,N_14042);
nand U18612 (N_18612,N_13566,N_13041);
nor U18613 (N_18613,N_12513,N_12875);
nand U18614 (N_18614,N_14024,N_14206);
or U18615 (N_18615,N_14932,N_14708);
and U18616 (N_18616,N_13819,N_15166);
xor U18617 (N_18617,N_14765,N_14573);
nor U18618 (N_18618,N_13303,N_14305);
xor U18619 (N_18619,N_13437,N_13266);
and U18620 (N_18620,N_14855,N_15540);
nor U18621 (N_18621,N_14409,N_13752);
and U18622 (N_18622,N_13522,N_14389);
nand U18623 (N_18623,N_12523,N_14845);
nand U18624 (N_18624,N_15370,N_12578);
xnor U18625 (N_18625,N_13504,N_13621);
and U18626 (N_18626,N_13103,N_13003);
nor U18627 (N_18627,N_13161,N_14339);
nor U18628 (N_18628,N_15138,N_12780);
or U18629 (N_18629,N_15025,N_14476);
nor U18630 (N_18630,N_14430,N_14869);
and U18631 (N_18631,N_12594,N_15379);
or U18632 (N_18632,N_15155,N_13342);
xor U18633 (N_18633,N_14205,N_15058);
nand U18634 (N_18634,N_14663,N_14105);
xor U18635 (N_18635,N_15163,N_14590);
and U18636 (N_18636,N_15389,N_13980);
xor U18637 (N_18637,N_13973,N_12627);
xor U18638 (N_18638,N_12954,N_15155);
and U18639 (N_18639,N_13788,N_14309);
xor U18640 (N_18640,N_14987,N_14712);
nor U18641 (N_18641,N_13938,N_12726);
nor U18642 (N_18642,N_13589,N_13418);
nand U18643 (N_18643,N_15094,N_15191);
or U18644 (N_18644,N_14113,N_15509);
xnor U18645 (N_18645,N_15229,N_14257);
and U18646 (N_18646,N_13814,N_14601);
nand U18647 (N_18647,N_13453,N_15134);
xor U18648 (N_18648,N_13234,N_15426);
nand U18649 (N_18649,N_14066,N_12926);
nand U18650 (N_18650,N_14201,N_13757);
nor U18651 (N_18651,N_15610,N_14791);
and U18652 (N_18652,N_15390,N_14304);
or U18653 (N_18653,N_12826,N_12771);
xor U18654 (N_18654,N_15217,N_15486);
or U18655 (N_18655,N_12533,N_15387);
xnor U18656 (N_18656,N_13724,N_13636);
and U18657 (N_18657,N_15438,N_14908);
nand U18658 (N_18658,N_14819,N_15160);
or U18659 (N_18659,N_14837,N_15104);
nand U18660 (N_18660,N_14061,N_15157);
nand U18661 (N_18661,N_15318,N_12716);
or U18662 (N_18662,N_12593,N_14690);
nand U18663 (N_18663,N_12528,N_12939);
and U18664 (N_18664,N_14018,N_13901);
and U18665 (N_18665,N_14549,N_14469);
nor U18666 (N_18666,N_13975,N_14302);
nand U18667 (N_18667,N_12824,N_13760);
nor U18668 (N_18668,N_13841,N_15255);
or U18669 (N_18669,N_14259,N_13472);
xor U18670 (N_18670,N_13336,N_15394);
nand U18671 (N_18671,N_12583,N_12541);
and U18672 (N_18672,N_13597,N_14983);
nand U18673 (N_18673,N_15196,N_14121);
nor U18674 (N_18674,N_15406,N_15425);
and U18675 (N_18675,N_15201,N_15463);
nand U18676 (N_18676,N_14860,N_12746);
or U18677 (N_18677,N_14242,N_12537);
nor U18678 (N_18678,N_14606,N_12507);
nand U18679 (N_18679,N_14844,N_15255);
xnor U18680 (N_18680,N_12599,N_14028);
nand U18681 (N_18681,N_13865,N_14700);
xor U18682 (N_18682,N_14822,N_13022);
xor U18683 (N_18683,N_12791,N_12884);
nand U18684 (N_18684,N_15590,N_15394);
or U18685 (N_18685,N_12703,N_13235);
and U18686 (N_18686,N_14393,N_13803);
or U18687 (N_18687,N_15444,N_12659);
nor U18688 (N_18688,N_13010,N_15266);
nor U18689 (N_18689,N_12578,N_14600);
nor U18690 (N_18690,N_14139,N_14626);
xor U18691 (N_18691,N_14917,N_15417);
nand U18692 (N_18692,N_14835,N_13658);
xnor U18693 (N_18693,N_13816,N_14018);
nor U18694 (N_18694,N_12823,N_13969);
or U18695 (N_18695,N_14490,N_13239);
xor U18696 (N_18696,N_12904,N_12953);
nor U18697 (N_18697,N_13261,N_14969);
xor U18698 (N_18698,N_14015,N_14515);
nand U18699 (N_18699,N_13508,N_14022);
nor U18700 (N_18700,N_13328,N_14699);
nor U18701 (N_18701,N_13645,N_14616);
and U18702 (N_18702,N_13120,N_13020);
and U18703 (N_18703,N_15347,N_12695);
xnor U18704 (N_18704,N_14998,N_14244);
or U18705 (N_18705,N_15614,N_14689);
nor U18706 (N_18706,N_14554,N_13466);
nand U18707 (N_18707,N_13794,N_15188);
or U18708 (N_18708,N_13384,N_13101);
or U18709 (N_18709,N_15052,N_14675);
nor U18710 (N_18710,N_14757,N_14716);
xor U18711 (N_18711,N_15357,N_14597);
nand U18712 (N_18712,N_12997,N_14618);
xor U18713 (N_18713,N_15075,N_13183);
or U18714 (N_18714,N_14210,N_14682);
or U18715 (N_18715,N_14129,N_14502);
or U18716 (N_18716,N_15270,N_13281);
nor U18717 (N_18717,N_13972,N_13835);
nor U18718 (N_18718,N_13129,N_14644);
nand U18719 (N_18719,N_15237,N_15475);
nor U18720 (N_18720,N_15196,N_15427);
xnor U18721 (N_18721,N_14569,N_14347);
nand U18722 (N_18722,N_13573,N_12602);
xor U18723 (N_18723,N_12929,N_14724);
nor U18724 (N_18724,N_13292,N_15082);
and U18725 (N_18725,N_13757,N_14319);
xnor U18726 (N_18726,N_13657,N_14600);
nor U18727 (N_18727,N_15184,N_13830);
nor U18728 (N_18728,N_14799,N_13877);
and U18729 (N_18729,N_14236,N_13355);
xnor U18730 (N_18730,N_13087,N_14109);
nand U18731 (N_18731,N_12784,N_14461);
xor U18732 (N_18732,N_15461,N_14099);
or U18733 (N_18733,N_12541,N_15038);
nor U18734 (N_18734,N_14492,N_13972);
or U18735 (N_18735,N_13088,N_15113);
nor U18736 (N_18736,N_14280,N_13169);
nor U18737 (N_18737,N_12631,N_14811);
nand U18738 (N_18738,N_15134,N_14092);
and U18739 (N_18739,N_13208,N_14446);
xnor U18740 (N_18740,N_13278,N_13926);
or U18741 (N_18741,N_15088,N_14024);
nand U18742 (N_18742,N_15039,N_13138);
or U18743 (N_18743,N_14184,N_13951);
xor U18744 (N_18744,N_14985,N_14544);
nand U18745 (N_18745,N_15610,N_14942);
xor U18746 (N_18746,N_13624,N_15230);
and U18747 (N_18747,N_14535,N_15286);
nand U18748 (N_18748,N_15169,N_13690);
xor U18749 (N_18749,N_15211,N_13434);
and U18750 (N_18750,N_18242,N_18401);
nand U18751 (N_18751,N_16907,N_16992);
nand U18752 (N_18752,N_17244,N_15750);
or U18753 (N_18753,N_17996,N_17889);
xnor U18754 (N_18754,N_18697,N_16960);
nor U18755 (N_18755,N_16072,N_17347);
or U18756 (N_18756,N_18325,N_17675);
nor U18757 (N_18757,N_18132,N_17789);
nor U18758 (N_18758,N_16143,N_16521);
nand U18759 (N_18759,N_16864,N_17614);
or U18760 (N_18760,N_15857,N_17512);
and U18761 (N_18761,N_15964,N_18318);
and U18762 (N_18762,N_18557,N_17034);
or U18763 (N_18763,N_16162,N_16855);
nand U18764 (N_18764,N_16311,N_17064);
xor U18765 (N_18765,N_16950,N_17989);
and U18766 (N_18766,N_18108,N_16736);
and U18767 (N_18767,N_17710,N_16623);
nor U18768 (N_18768,N_18512,N_18498);
or U18769 (N_18769,N_18040,N_16172);
or U18770 (N_18770,N_17121,N_15961);
or U18771 (N_18771,N_16880,N_15921);
or U18772 (N_18772,N_18342,N_17340);
and U18773 (N_18773,N_17550,N_16023);
nor U18774 (N_18774,N_16624,N_16375);
nor U18775 (N_18775,N_17664,N_16042);
or U18776 (N_18776,N_18319,N_16325);
xnor U18777 (N_18777,N_18485,N_17676);
nand U18778 (N_18778,N_17902,N_15922);
xnor U18779 (N_18779,N_16625,N_15655);
nand U18780 (N_18780,N_17501,N_17611);
nand U18781 (N_18781,N_17848,N_18380);
xnor U18782 (N_18782,N_18470,N_16659);
nand U18783 (N_18783,N_15901,N_16179);
or U18784 (N_18784,N_16173,N_15823);
nand U18785 (N_18785,N_17677,N_16901);
nor U18786 (N_18786,N_16323,N_16440);
nand U18787 (N_18787,N_18431,N_18373);
nor U18788 (N_18788,N_17615,N_17843);
and U18789 (N_18789,N_18117,N_18678);
nand U18790 (N_18790,N_16927,N_16879);
and U18791 (N_18791,N_18475,N_16706);
nand U18792 (N_18792,N_17195,N_15996);
or U18793 (N_18793,N_17280,N_18698);
and U18794 (N_18794,N_17791,N_18610);
or U18795 (N_18795,N_16414,N_17020);
or U18796 (N_18796,N_18227,N_15839);
nand U18797 (N_18797,N_17187,N_16175);
xnor U18798 (N_18798,N_18229,N_18454);
xnor U18799 (N_18799,N_18462,N_16987);
or U18800 (N_18800,N_16244,N_16158);
and U18801 (N_18801,N_18039,N_18712);
or U18802 (N_18802,N_16603,N_17122);
nor U18803 (N_18803,N_18527,N_16818);
nand U18804 (N_18804,N_18400,N_17780);
nand U18805 (N_18805,N_17527,N_17487);
nor U18806 (N_18806,N_17962,N_16575);
nand U18807 (N_18807,N_18734,N_17826);
nand U18808 (N_18808,N_16384,N_17531);
xor U18809 (N_18809,N_16665,N_16214);
or U18810 (N_18810,N_17157,N_16981);
nor U18811 (N_18811,N_15827,N_15738);
nand U18812 (N_18812,N_17464,N_18649);
nand U18813 (N_18813,N_17707,N_16290);
nor U18814 (N_18814,N_16117,N_15676);
nand U18815 (N_18815,N_16049,N_16641);
or U18816 (N_18816,N_18731,N_16734);
nor U18817 (N_18817,N_16144,N_17285);
xnor U18818 (N_18818,N_17085,N_16269);
or U18819 (N_18819,N_15999,N_18572);
and U18820 (N_18820,N_16620,N_16961);
nand U18821 (N_18821,N_16443,N_18410);
and U18822 (N_18822,N_15887,N_17587);
xnor U18823 (N_18823,N_16016,N_15840);
or U18824 (N_18824,N_15733,N_15792);
nand U18825 (N_18825,N_17733,N_16523);
xor U18826 (N_18826,N_15636,N_18099);
and U18827 (N_18827,N_16115,N_16590);
and U18828 (N_18828,N_15638,N_17724);
and U18829 (N_18829,N_15751,N_16487);
nand U18830 (N_18830,N_16225,N_18633);
and U18831 (N_18831,N_17875,N_17618);
xor U18832 (N_18832,N_17196,N_15930);
and U18833 (N_18833,N_17720,N_16387);
or U18834 (N_18834,N_16089,N_16608);
nand U18835 (N_18835,N_16207,N_16218);
xor U18836 (N_18836,N_17021,N_17032);
nand U18837 (N_18837,N_15943,N_16632);
xor U18838 (N_18838,N_16717,N_16490);
or U18839 (N_18839,N_17217,N_18012);
nor U18840 (N_18840,N_15966,N_18049);
and U18841 (N_18841,N_16974,N_18658);
or U18842 (N_18842,N_18134,N_16531);
and U18843 (N_18843,N_18064,N_17903);
and U18844 (N_18844,N_18044,N_17312);
xor U18845 (N_18845,N_17648,N_16810);
nor U18846 (N_18846,N_16161,N_17518);
nand U18847 (N_18847,N_18381,N_15934);
nand U18848 (N_18848,N_16655,N_16931);
and U18849 (N_18849,N_18162,N_18383);
and U18850 (N_18850,N_16837,N_15926);
nor U18851 (N_18851,N_15735,N_17380);
nand U18852 (N_18852,N_17560,N_17855);
nand U18853 (N_18853,N_16825,N_16013);
nor U18854 (N_18854,N_17907,N_16560);
nand U18855 (N_18855,N_18091,N_16555);
nor U18856 (N_18856,N_15991,N_16688);
or U18857 (N_18857,N_15853,N_17559);
or U18858 (N_18858,N_17951,N_17123);
nor U18859 (N_18859,N_17837,N_18078);
nor U18860 (N_18860,N_17808,N_18034);
and U18861 (N_18861,N_16988,N_16796);
or U18862 (N_18862,N_16871,N_17066);
nor U18863 (N_18863,N_16150,N_16829);
xor U18864 (N_18864,N_16803,N_15666);
and U18865 (N_18865,N_17114,N_16365);
and U18866 (N_18866,N_17008,N_17170);
xor U18867 (N_18867,N_16569,N_17961);
or U18868 (N_18868,N_16294,N_17221);
xnor U18869 (N_18869,N_16411,N_16128);
nor U18870 (N_18870,N_16692,N_17983);
xnor U18871 (N_18871,N_15803,N_15771);
xnor U18872 (N_18872,N_16995,N_18194);
xnor U18873 (N_18873,N_17508,N_17212);
nor U18874 (N_18874,N_15679,N_15931);
xor U18875 (N_18875,N_16121,N_18423);
nor U18876 (N_18876,N_15650,N_16631);
nor U18877 (N_18877,N_15872,N_18670);
nand U18878 (N_18878,N_16505,N_17866);
or U18879 (N_18879,N_17824,N_16522);
xor U18880 (N_18880,N_16842,N_18285);
xnor U18881 (N_18881,N_17003,N_16898);
or U18882 (N_18882,N_15911,N_15706);
xor U18883 (N_18883,N_15767,N_15932);
nor U18884 (N_18884,N_17155,N_17940);
or U18885 (N_18885,N_15625,N_16782);
nor U18886 (N_18886,N_17314,N_17214);
nand U18887 (N_18887,N_16817,N_17722);
nor U18888 (N_18888,N_17461,N_16787);
and U18889 (N_18889,N_15816,N_15742);
or U18890 (N_18890,N_16820,N_16762);
xor U18891 (N_18891,N_17143,N_15710);
and U18892 (N_18892,N_15763,N_17050);
nand U18893 (N_18893,N_16566,N_16682);
and U18894 (N_18894,N_18617,N_17140);
and U18895 (N_18895,N_18743,N_17876);
and U18896 (N_18896,N_18143,N_17953);
nor U18897 (N_18897,N_18449,N_16602);
xnor U18898 (N_18898,N_15660,N_16024);
nand U18899 (N_18899,N_18080,N_16638);
and U18900 (N_18900,N_18320,N_17905);
nand U18901 (N_18901,N_16004,N_17842);
nor U18902 (N_18902,N_16304,N_15790);
xor U18903 (N_18903,N_16199,N_16853);
nor U18904 (N_18904,N_17922,N_17575);
or U18905 (N_18905,N_15799,N_18144);
xor U18906 (N_18906,N_18556,N_16243);
nand U18907 (N_18907,N_18187,N_17916);
and U18908 (N_18908,N_16576,N_17054);
nand U18909 (N_18909,N_16288,N_17367);
or U18910 (N_18910,N_17466,N_16937);
and U18911 (N_18911,N_17556,N_15835);
nor U18912 (N_18912,N_18713,N_17514);
nor U18913 (N_18913,N_17713,N_16592);
nand U18914 (N_18914,N_16756,N_16877);
or U18915 (N_18915,N_18459,N_15651);
nor U18916 (N_18916,N_18122,N_18161);
or U18917 (N_18917,N_15800,N_17306);
nor U18918 (N_18918,N_16562,N_17330);
and U18919 (N_18919,N_17385,N_16697);
xor U18920 (N_18920,N_17685,N_17072);
nand U18921 (N_18921,N_16431,N_16125);
nor U18922 (N_18922,N_16472,N_17832);
xnor U18923 (N_18923,N_15941,N_18408);
nand U18924 (N_18924,N_17679,N_17370);
or U18925 (N_18925,N_17012,N_15987);
and U18926 (N_18926,N_17625,N_18145);
or U18927 (N_18927,N_16183,N_17831);
nand U18928 (N_18928,N_17153,N_18165);
or U18929 (N_18929,N_16619,N_18450);
nand U18930 (N_18930,N_16181,N_16684);
or U18931 (N_18931,N_18586,N_16141);
or U18932 (N_18932,N_17346,N_17304);
and U18933 (N_18933,N_18191,N_18477);
and U18934 (N_18934,N_17451,N_17599);
and U18935 (N_18935,N_18277,N_18314);
and U18936 (N_18936,N_16465,N_15741);
nand U18937 (N_18937,N_15694,N_17095);
xnor U18938 (N_18938,N_17391,N_17883);
and U18939 (N_18939,N_17551,N_16367);
nand U18940 (N_18940,N_15865,N_16654);
or U18941 (N_18941,N_16852,N_16839);
nand U18942 (N_18942,N_16498,N_18066);
nand U18943 (N_18943,N_18447,N_17488);
or U18944 (N_18944,N_18192,N_16667);
and U18945 (N_18945,N_18196,N_16231);
nand U18946 (N_18946,N_16130,N_16473);
xnor U18947 (N_18947,N_18736,N_17361);
xnor U18948 (N_18948,N_16398,N_17421);
xnor U18949 (N_18949,N_17406,N_17965);
nand U18950 (N_18950,N_16280,N_17430);
and U18951 (N_18951,N_17943,N_16957);
xor U18952 (N_18952,N_15725,N_17608);
or U18953 (N_18953,N_18024,N_18486);
nand U18954 (N_18954,N_16196,N_17019);
or U18955 (N_18955,N_16405,N_16836);
and U18956 (N_18956,N_18359,N_16788);
and U18957 (N_18957,N_17245,N_16681);
nand U18958 (N_18958,N_16362,N_18283);
nand U18959 (N_18959,N_17727,N_17117);
or U18960 (N_18960,N_17543,N_18582);
and U18961 (N_18961,N_17394,N_17165);
xor U18962 (N_18962,N_16593,N_16772);
xor U18963 (N_18963,N_16097,N_17339);
xor U18964 (N_18964,N_17337,N_18326);
nand U18965 (N_18965,N_17975,N_15808);
or U18966 (N_18966,N_17368,N_18136);
xor U18967 (N_18967,N_15635,N_16709);
nand U18968 (N_18968,N_17523,N_17649);
nand U18969 (N_18969,N_15728,N_16530);
or U18970 (N_18970,N_17735,N_18186);
and U18971 (N_18971,N_18570,N_17257);
or U18972 (N_18972,N_15830,N_16542);
and U18973 (N_18973,N_17070,N_18421);
nand U18974 (N_18974,N_16939,N_16537);
or U18975 (N_18975,N_16263,N_18732);
and U18976 (N_18976,N_16113,N_17626);
or U18977 (N_18977,N_17749,N_17432);
and U18978 (N_18978,N_18112,N_17513);
nor U18979 (N_18979,N_17183,N_16869);
or U18980 (N_18980,N_17356,N_18716);
nor U18981 (N_18981,N_17005,N_16303);
nand U18982 (N_18982,N_17783,N_17519);
and U18983 (N_18983,N_17554,N_16038);
nor U18984 (N_18984,N_17211,N_17341);
nand U18985 (N_18985,N_16336,N_17628);
and U18986 (N_18986,N_17033,N_17112);
nand U18987 (N_18987,N_17784,N_17498);
nand U18988 (N_18988,N_18173,N_18491);
or U18989 (N_18989,N_16066,N_16660);
nor U18990 (N_18990,N_17851,N_16985);
and U18991 (N_18991,N_18648,N_16731);
and U18992 (N_18992,N_15673,N_18749);
and U18993 (N_18993,N_18123,N_18175);
nand U18994 (N_18994,N_18211,N_16159);
and U18995 (N_18995,N_16201,N_16238);
or U18996 (N_18996,N_15717,N_16618);
nor U18997 (N_18997,N_18398,N_18376);
or U18998 (N_18998,N_18234,N_16563);
or U18999 (N_18999,N_17874,N_16647);
and U19000 (N_19000,N_17775,N_17793);
or U19001 (N_19001,N_16363,N_16330);
nor U19002 (N_19002,N_17145,N_17328);
nor U19003 (N_19003,N_17013,N_16503);
nand U19004 (N_19004,N_18608,N_18415);
nand U19005 (N_19005,N_16306,N_15977);
and U19006 (N_19006,N_17250,N_17094);
nor U19007 (N_19007,N_16342,N_17265);
nor U19008 (N_19008,N_16679,N_16899);
xor U19009 (N_19009,N_18038,N_16687);
nor U19010 (N_19010,N_17232,N_18439);
and U19011 (N_19011,N_18265,N_16055);
xor U19012 (N_19012,N_16636,N_17814);
nand U19013 (N_19013,N_18218,N_16751);
nand U19014 (N_19014,N_18026,N_17475);
xnor U19015 (N_19015,N_17447,N_18146);
or U19016 (N_19016,N_15925,N_15992);
xor U19017 (N_19017,N_18268,N_18082);
or U19018 (N_19018,N_18092,N_16978);
or U19019 (N_19019,N_15893,N_16467);
nor U19020 (N_19020,N_18510,N_15873);
nand U19021 (N_19021,N_16470,N_15978);
and U19022 (N_19022,N_15852,N_15713);
or U19023 (N_19023,N_18113,N_18696);
nand U19024 (N_19024,N_17087,N_17089);
or U19025 (N_19025,N_17437,N_16378);
or U19026 (N_19026,N_16257,N_17149);
and U19027 (N_19027,N_15755,N_17816);
nand U19028 (N_19028,N_16621,N_17827);
or U19029 (N_19029,N_17763,N_17416);
or U19030 (N_19030,N_17415,N_17815);
xor U19031 (N_19031,N_17926,N_16451);
nand U19032 (N_19032,N_18019,N_16613);
or U19033 (N_19033,N_18079,N_16334);
and U19034 (N_19034,N_16230,N_16020);
or U19035 (N_19035,N_16845,N_18427);
nor U19036 (N_19036,N_18666,N_16442);
or U19037 (N_19037,N_17563,N_16859);
or U19038 (N_19038,N_17798,N_17932);
nand U19039 (N_19039,N_18374,N_17018);
nor U19040 (N_19040,N_17409,N_16135);
and U19041 (N_19041,N_17662,N_16101);
and U19042 (N_19042,N_16381,N_17958);
and U19043 (N_19043,N_16552,N_18543);
nor U19044 (N_19044,N_16640,N_16471);
nand U19045 (N_19045,N_16022,N_18627);
and U19046 (N_19046,N_18336,N_17925);
and U19047 (N_19047,N_17132,N_17465);
nand U19048 (N_19048,N_18378,N_18093);
or U19049 (N_19049,N_17913,N_17452);
nor U19050 (N_19050,N_15786,N_16124);
xor U19051 (N_19051,N_18595,N_16132);
xnor U19052 (N_19052,N_16783,N_17056);
or U19053 (N_19053,N_15952,N_18180);
and U19054 (N_19054,N_16021,N_17166);
nand U19055 (N_19055,N_16675,N_18244);
nor U19056 (N_19056,N_17224,N_17116);
nand U19057 (N_19057,N_18115,N_16635);
and U19058 (N_19058,N_16938,N_17944);
nor U19059 (N_19059,N_16951,N_16652);
nor U19060 (N_19060,N_17109,N_17536);
xnor U19061 (N_19061,N_18324,N_15902);
or U19062 (N_19062,N_17717,N_18742);
nand U19063 (N_19063,N_16551,N_17841);
nand U19064 (N_19064,N_17379,N_18159);
xnor U19065 (N_19065,N_17960,N_18661);
xnor U19066 (N_19066,N_16801,N_15656);
xor U19067 (N_19067,N_18086,N_15683);
nand U19068 (N_19068,N_16104,N_16967);
nand U19069 (N_19069,N_16192,N_16668);
nand U19070 (N_19070,N_17890,N_17566);
nand U19071 (N_19071,N_15904,N_18256);
or U19072 (N_19072,N_18695,N_16459);
and U19073 (N_19073,N_15936,N_17800);
and U19074 (N_19074,N_16792,N_15971);
nand U19075 (N_19075,N_18509,N_17577);
xnor U19076 (N_19076,N_18521,N_18542);
nor U19077 (N_19077,N_18619,N_16823);
or U19078 (N_19078,N_18723,N_16401);
or U19079 (N_19079,N_18045,N_16850);
and U19080 (N_19080,N_16478,N_17100);
xor U19081 (N_19081,N_16308,N_18219);
xor U19082 (N_19082,N_16644,N_16559);
nand U19083 (N_19083,N_15628,N_16977);
xnor U19084 (N_19084,N_16744,N_18672);
nor U19085 (N_19085,N_16758,N_16476);
or U19086 (N_19086,N_15910,N_18217);
and U19087 (N_19087,N_16082,N_18601);
or U19088 (N_19088,N_16475,N_17811);
and U19089 (N_19089,N_16773,N_18693);
xor U19090 (N_19090,N_16106,N_16760);
and U19091 (N_19091,N_18530,N_16678);
nor U19092 (N_19092,N_16033,N_18225);
xnor U19093 (N_19093,N_15984,N_16002);
xor U19094 (N_19094,N_16917,N_16204);
nand U19095 (N_19095,N_18652,N_18281);
or U19096 (N_19096,N_17045,N_17027);
and U19097 (N_19097,N_18206,N_15745);
and U19098 (N_19098,N_18573,N_16955);
nor U19099 (N_19099,N_18032,N_15782);
and U19100 (N_19100,N_18356,N_16427);
nand U19101 (N_19101,N_18520,N_16509);
xnor U19102 (N_19102,N_16036,N_17291);
nor U19103 (N_19103,N_16941,N_16497);
nand U19104 (N_19104,N_16168,N_16319);
nand U19105 (N_19105,N_16942,N_17230);
or U19106 (N_19106,N_16188,N_17062);
xnor U19107 (N_19107,N_17180,N_16556);
and U19108 (N_19108,N_18630,N_16532);
nand U19109 (N_19109,N_17863,N_18369);
nand U19110 (N_19110,N_17359,N_17867);
nand U19111 (N_19111,N_18035,N_15897);
xnor U19112 (N_19112,N_18478,N_16348);
xor U19113 (N_19113,N_18167,N_18626);
or U19114 (N_19114,N_16351,N_16291);
nand U19115 (N_19115,N_16253,N_16081);
or U19116 (N_19116,N_17468,N_17968);
nor U19117 (N_19117,N_17923,N_17266);
xnor U19118 (N_19118,N_18585,N_17030);
or U19119 (N_19119,N_18558,N_18008);
nor U19120 (N_19120,N_16286,N_16360);
and U19121 (N_19121,N_18338,N_16127);
xnor U19122 (N_19122,N_18065,N_17980);
or U19123 (N_19123,N_18027,N_17194);
xor U19124 (N_19124,N_16146,N_16838);
nor U19125 (N_19125,N_16494,N_18534);
nor U19126 (N_19126,N_18523,N_17029);
nand U19127 (N_19127,N_17725,N_17795);
xnor U19128 (N_19128,N_17739,N_18298);
nand U19129 (N_19129,N_16428,N_18135);
or U19130 (N_19130,N_16458,N_17311);
nand U19131 (N_19131,N_16313,N_15898);
xnor U19132 (N_19132,N_18286,N_16627);
or U19133 (N_19133,N_16956,N_15658);
or U19134 (N_19134,N_17900,N_16163);
nor U19135 (N_19135,N_18511,N_16174);
nor U19136 (N_19136,N_17423,N_16867);
nand U19137 (N_19137,N_16843,N_15736);
nand U19138 (N_19138,N_16572,N_18334);
nor U19139 (N_19139,N_18016,N_18264);
xor U19140 (N_19140,N_18569,N_17000);
nand U19141 (N_19141,N_17290,N_16203);
and U19142 (N_19142,N_16584,N_16764);
nand U19143 (N_19143,N_15630,N_15862);
nor U19144 (N_19144,N_17759,N_15959);
or U19145 (N_19145,N_16380,N_16748);
and U19146 (N_19146,N_16982,N_17582);
or U19147 (N_19147,N_18596,N_16295);
and U19148 (N_19148,N_16239,N_18011);
and U19149 (N_19149,N_18352,N_18499);
nor U19150 (N_19150,N_16088,N_17681);
nor U19151 (N_19151,N_18289,N_16695);
and U19152 (N_19152,N_17918,N_18006);
xor U19153 (N_19153,N_15720,N_18212);
nand U19154 (N_19154,N_16601,N_15748);
nand U19155 (N_19155,N_17193,N_17317);
nor U19156 (N_19156,N_16733,N_16084);
nor U19157 (N_19157,N_16595,N_18240);
nor U19158 (N_19158,N_16702,N_18654);
and U19159 (N_19159,N_17431,N_18272);
xor U19160 (N_19160,N_18188,N_16166);
nor U19161 (N_19161,N_17134,N_16637);
nand U19162 (N_19162,N_16226,N_18055);
nor U19163 (N_19163,N_16256,N_16646);
or U19164 (N_19164,N_17239,N_16857);
nor U19165 (N_19165,N_18437,N_18405);
or U19166 (N_19166,N_15734,N_16683);
xor U19167 (N_19167,N_18166,N_16177);
nor U19168 (N_19168,N_17270,N_16714);
nor U19169 (N_19169,N_15970,N_18645);
nor U19170 (N_19170,N_17090,N_17839);
nand U19171 (N_19171,N_18153,N_15883);
xnor U19172 (N_19172,N_17641,N_18660);
nand U19173 (N_19173,N_18302,N_18124);
nor U19174 (N_19174,N_15817,N_15807);
nand U19175 (N_19175,N_18270,N_15983);
or U19176 (N_19176,N_17715,N_16276);
nand U19177 (N_19177,N_16205,N_18213);
nor U19178 (N_19178,N_16222,N_17186);
nand U19179 (N_19179,N_15701,N_17610);
nor U19180 (N_19180,N_15798,N_17490);
or U19181 (N_19181,N_17762,N_16185);
nor U19182 (N_19182,N_17711,N_16260);
or U19183 (N_19183,N_18689,N_18054);
and U19184 (N_19184,N_16495,N_16420);
and U19185 (N_19185,N_15815,N_15914);
and U19186 (N_19186,N_18399,N_18453);
xnor U19187 (N_19187,N_15882,N_16518);
and U19188 (N_19188,N_18532,N_17240);
nand U19189 (N_19189,N_16897,N_17429);
and U19190 (N_19190,N_16975,N_15659);
xnor U19191 (N_19191,N_18517,N_18390);
nor U19192 (N_19192,N_16482,N_17738);
or U19193 (N_19193,N_17173,N_16468);
xnor U19194 (N_19194,N_18476,N_15704);
and U19195 (N_19195,N_18140,N_16596);
and U19196 (N_19196,N_17017,N_18550);
nor U19197 (N_19197,N_18540,N_16212);
xnor U19198 (N_19198,N_17928,N_15796);
nor U19199 (N_19199,N_16355,N_17689);
nand U19200 (N_19200,N_16377,N_17834);
nor U19201 (N_19201,N_17769,N_17489);
and U19202 (N_19202,N_17313,N_17522);
and U19203 (N_19203,N_16670,N_16364);
xor U19204 (N_19204,N_15811,N_17573);
nand U19205 (N_19205,N_17172,N_15677);
and U19206 (N_19206,N_16945,N_16432);
or U19207 (N_19207,N_15654,N_17039);
and U19208 (N_19208,N_17603,N_16202);
xnor U19209 (N_19209,N_17102,N_15956);
nand U19210 (N_19210,N_15661,N_16298);
nor U19211 (N_19211,N_18396,N_18622);
or U19212 (N_19212,N_17504,N_16557);
or U19213 (N_19213,N_17131,N_16010);
xor U19214 (N_19214,N_18157,N_18002);
xor U19215 (N_19215,N_17700,N_16356);
or U19216 (N_19216,N_15855,N_17549);
nand U19217 (N_19217,N_17857,N_16689);
nand U19218 (N_19218,N_17301,N_18052);
nand U19219 (N_19219,N_17515,N_16711);
xnor U19220 (N_19220,N_17741,N_15876);
nand U19221 (N_19221,N_16271,N_18448);
nor U19222 (N_19222,N_17390,N_17188);
and U19223 (N_19223,N_17092,N_18358);
nor U19224 (N_19224,N_16399,N_16379);
nor U19225 (N_19225,N_18551,N_16107);
and U19226 (N_19226,N_15861,N_16481);
and U19227 (N_19227,N_16821,N_16616);
nor U19228 (N_19228,N_16197,N_18306);
nand U19229 (N_19229,N_16352,N_17009);
nor U19230 (N_19230,N_16402,N_15705);
nand U19231 (N_19231,N_16131,N_16519);
nor U19232 (N_19232,N_18360,N_17979);
nand U19233 (N_19233,N_16317,N_17539);
or U19234 (N_19234,N_18456,N_17654);
xnor U19235 (N_19235,N_17668,N_17892);
or U19236 (N_19236,N_16030,N_17927);
or U19237 (N_19237,N_17364,N_17378);
or U19238 (N_19238,N_17491,N_16320);
nand U19239 (N_19239,N_16565,N_17434);
nor U19240 (N_19240,N_17154,N_17643);
xor U19241 (N_19241,N_17872,N_16134);
xnor U19242 (N_19242,N_15986,N_16996);
and U19243 (N_19243,N_15788,N_18465);
xor U19244 (N_19244,N_16726,N_17956);
or U19245 (N_19245,N_16903,N_18015);
or U19246 (N_19246,N_16114,N_15772);
xor U19247 (N_19247,N_16582,N_17142);
nor U19248 (N_19248,N_16533,N_16567);
and U19249 (N_19249,N_15770,N_17395);
or U19250 (N_19250,N_18490,N_18254);
nand U19251 (N_19251,N_17790,N_18330);
xor U19252 (N_19252,N_15975,N_16730);
nand U19253 (N_19253,N_15685,N_16890);
nand U19254 (N_19254,N_18443,N_15859);
xnor U19255 (N_19255,N_16287,N_18579);
nand U19256 (N_19256,N_18100,N_16888);
or U19257 (N_19257,N_17865,N_16457);
or U19258 (N_19258,N_17520,N_16261);
and U19259 (N_19259,N_16064,N_17545);
or U19260 (N_19260,N_17308,N_16310);
and U19261 (N_19261,N_16909,N_17580);
and U19262 (N_19262,N_15825,N_15828);
nor U19263 (N_19263,N_17691,N_16182);
nor U19264 (N_19264,N_16354,N_17369);
nor U19265 (N_19265,N_17253,N_18593);
nor U19266 (N_19266,N_15648,N_18323);
xnor U19267 (N_19267,N_15715,N_17078);
nor U19268 (N_19268,N_17402,N_18539);
xor U19269 (N_19269,N_16191,N_16546);
and U19270 (N_19270,N_17650,N_16246);
nor U19271 (N_19271,N_15870,N_16753);
nor U19272 (N_19272,N_16242,N_17609);
and U19273 (N_19273,N_16410,N_18007);
nor U19274 (N_19274,N_16292,N_16275);
nor U19275 (N_19275,N_17829,N_18528);
and U19276 (N_19276,N_17524,N_18250);
nor U19277 (N_19277,N_17503,N_18350);
nand U19278 (N_19278,N_17321,N_18022);
nand U19279 (N_19279,N_15821,N_18245);
nor U19280 (N_19280,N_16254,N_18199);
and U19281 (N_19281,N_18018,N_15678);
nor U19282 (N_19282,N_15969,N_17098);
or U19283 (N_19283,N_16460,N_17093);
nand U19284 (N_19284,N_16190,N_17743);
or U19285 (N_19285,N_17938,N_16568);
nand U19286 (N_19286,N_16068,N_17215);
or U19287 (N_19287,N_16077,N_16433);
and U19288 (N_19288,N_18504,N_16963);
nand U19289 (N_19289,N_16933,N_18571);
and U19290 (N_19290,N_18704,N_16693);
or U19291 (N_19291,N_17723,N_18300);
and U19292 (N_19292,N_15693,N_16844);
and U19293 (N_19293,N_16847,N_18740);
nand U19294 (N_19294,N_15894,N_15851);
nor U19295 (N_19295,N_16108,N_17462);
xor U19296 (N_19296,N_17819,N_18119);
xnor U19297 (N_19297,N_16449,N_18328);
nand U19298 (N_19298,N_15831,N_17561);
nor U19299 (N_19299,N_15791,N_16591);
nor U19300 (N_19300,N_17365,N_18483);
nand U19301 (N_19301,N_15916,N_16932);
xnor U19302 (N_19302,N_16883,N_16832);
and U19303 (N_19303,N_16894,N_16430);
xor U19304 (N_19304,N_16887,N_15814);
nand U19305 (N_19305,N_18241,N_18687);
nand U19306 (N_19306,N_16949,N_18745);
or U19307 (N_19307,N_18293,N_17974);
xnor U19308 (N_19308,N_16766,N_16701);
nand U19309 (N_19309,N_16797,N_16281);
nor U19310 (N_19310,N_16170,N_18208);
xnor U19311 (N_19311,N_16496,N_17647);
or U19312 (N_19312,N_17113,N_16923);
and U19313 (N_19313,N_17624,N_18674);
or U19314 (N_19314,N_16710,N_17146);
nand U19315 (N_19315,N_16740,N_16573);
and U19316 (N_19316,N_17209,N_17480);
xnor U19317 (N_19317,N_16780,N_18118);
and U19318 (N_19318,N_17593,N_16318);
xnor U19319 (N_19319,N_18411,N_16406);
nand U19320 (N_19320,N_16483,N_18675);
nor U19321 (N_19321,N_16041,N_15626);
nor U19322 (N_19322,N_17088,N_17469);
or U19323 (N_19323,N_16598,N_17777);
or U19324 (N_19324,N_17761,N_15995);
and U19325 (N_19325,N_18299,N_15880);
nor U19326 (N_19326,N_17381,N_17198);
xnor U19327 (N_19327,N_16849,N_16129);
xnor U19328 (N_19328,N_17684,N_17315);
or U19329 (N_19329,N_17097,N_15958);
nor U19330 (N_19330,N_16926,N_18640);
or U19331 (N_19331,N_18612,N_17110);
or U19332 (N_19332,N_18163,N_16585);
nor U19333 (N_19333,N_18471,N_18105);
nor U19334 (N_19334,N_18541,N_17970);
xor U19335 (N_19335,N_16997,N_17424);
or U19336 (N_19336,N_16372,N_15634);
xor U19337 (N_19337,N_16396,N_17178);
and U19338 (N_19338,N_17758,N_17111);
nor U19339 (N_19339,N_15854,N_17274);
and U19340 (N_19340,N_16816,N_17588);
nand U19341 (N_19341,N_17383,N_16513);
nor U19342 (N_19342,N_17252,N_18735);
and U19343 (N_19343,N_18368,N_17617);
and U19344 (N_19344,N_17258,N_16370);
nor U19345 (N_19345,N_16012,N_16031);
nor U19346 (N_19346,N_18518,N_17915);
nand U19347 (N_19347,N_17342,N_17184);
or U19348 (N_19348,N_18682,N_17982);
xnor U19349 (N_19349,N_18371,N_16444);
nand U19350 (N_19350,N_16579,N_16630);
nor U19351 (N_19351,N_15919,N_16180);
and U19352 (N_19352,N_16570,N_16614);
nand U19353 (N_19353,N_18094,N_18102);
nor U19354 (N_19354,N_15973,N_16831);
nor U19355 (N_19355,N_17043,N_15924);
and U19356 (N_19356,N_18058,N_18137);
and U19357 (N_19357,N_16014,N_16969);
and U19358 (N_19358,N_17917,N_16723);
nand U19359 (N_19359,N_16112,N_15841);
and U19360 (N_19360,N_16790,N_16305);
nor U19361 (N_19361,N_18533,N_17233);
and U19362 (N_19362,N_16027,N_16011);
nand U19363 (N_19363,N_17334,N_16296);
and U19364 (N_19364,N_17655,N_16650);
nand U19365 (N_19365,N_16904,N_17332);
xor U19366 (N_19366,N_15730,N_16000);
and U19367 (N_19367,N_17190,N_18657);
nor U19368 (N_19368,N_16245,N_18574);
nor U19369 (N_19369,N_17663,N_17806);
nand U19370 (N_19370,N_17694,N_17517);
or U19371 (N_19371,N_16767,N_18525);
nand U19372 (N_19372,N_17755,N_17533);
nor U19373 (N_19373,N_17007,N_18535);
nand U19374 (N_19374,N_18284,N_17644);
and U19375 (N_19375,N_16463,N_17854);
or U19376 (N_19376,N_17442,N_17680);
xnor U19377 (N_19377,N_16333,N_17399);
and U19378 (N_19378,N_17197,N_17752);
or U19379 (N_19379,N_17828,N_16703);
or U19380 (N_19380,N_17467,N_16167);
or U19381 (N_19381,N_15822,N_17605);
and U19382 (N_19382,N_17570,N_17776);
xnor U19383 (N_19383,N_15990,N_17323);
or U19384 (N_19384,N_18364,N_18588);
nor U19385 (N_19385,N_16919,N_17191);
or U19386 (N_19386,N_16746,N_16622);
or U19387 (N_19387,N_17287,N_16283);
or U19388 (N_19388,N_18057,N_16805);
and U19389 (N_19389,N_16452,N_16340);
nor U19390 (N_19390,N_17049,N_16865);
xnor U19391 (N_19391,N_17853,N_18632);
nor U19392 (N_19392,N_17478,N_16854);
xnor U19393 (N_19393,N_15794,N_18659);
or U19394 (N_19394,N_16881,N_16139);
or U19395 (N_19395,N_18222,N_17147);
xor U19396 (N_19396,N_16065,N_15632);
xnor U19397 (N_19397,N_16833,N_17683);
and U19398 (N_19398,N_17813,N_15645);
nor U19399 (N_19399,N_15805,N_16725);
xnor U19400 (N_19400,N_17886,N_15866);
xor U19401 (N_19401,N_17978,N_16661);
or U19402 (N_19402,N_18559,N_17718);
and U19403 (N_19403,N_16133,N_16464);
or U19404 (N_19404,N_16747,N_15692);
or U19405 (N_19405,N_16233,N_16524);
or U19406 (N_19406,N_17223,N_16798);
or U19407 (N_19407,N_18395,N_15933);
nand U19408 (N_19408,N_16332,N_18098);
and U19409 (N_19409,N_18121,N_17001);
nand U19410 (N_19410,N_16578,N_17870);
and U19411 (N_19411,N_17278,N_18239);
nor U19412 (N_19412,N_16017,N_18109);
xor U19413 (N_19413,N_17282,N_17228);
xor U19414 (N_19414,N_17534,N_18583);
or U19415 (N_19415,N_16285,N_17740);
nand U19416 (N_19416,N_18650,N_17820);
and U19417 (N_19417,N_18434,N_16581);
or U19418 (N_19418,N_17120,N_15842);
nand U19419 (N_19419,N_16908,N_15641);
xor U19420 (N_19420,N_18526,N_15888);
xnor U19421 (N_19421,N_16672,N_18127);
nor U19422 (N_19422,N_16329,N_18603);
or U19423 (N_19423,N_17083,N_16111);
nor U19424 (N_19424,N_17041,N_18479);
and U19425 (N_19425,N_16093,N_16404);
or U19426 (N_19426,N_16514,N_17275);
or U19427 (N_19427,N_18513,N_18154);
or U19428 (N_19428,N_18461,N_17426);
and U19429 (N_19429,N_17389,N_18329);
xnor U19430 (N_19430,N_16300,N_15960);
or U19431 (N_19431,N_17935,N_17771);
nor U19432 (N_19432,N_15949,N_16415);
or U19433 (N_19433,N_18656,N_16074);
nor U19434 (N_19434,N_15714,N_15649);
or U19435 (N_19435,N_17712,N_17022);
nor U19436 (N_19436,N_18436,N_17807);
xor U19437 (N_19437,N_15928,N_16639);
nor U19438 (N_19438,N_17473,N_16776);
xor U19439 (N_19439,N_17479,N_15849);
nor U19440 (N_19440,N_16079,N_17036);
nor U19441 (N_19441,N_18004,N_18139);
or U19442 (N_19442,N_18294,N_17991);
xor U19443 (N_19443,N_17080,N_16103);
nand U19444 (N_19444,N_18101,N_17037);
or U19445 (N_19445,N_17445,N_17325);
or U19446 (N_19446,N_17936,N_17057);
xor U19447 (N_19447,N_17630,N_16268);
or U19448 (N_19448,N_18620,N_16946);
and U19449 (N_19449,N_16943,N_16215);
nor U19450 (N_19450,N_16599,N_16044);
and U19451 (N_19451,N_18391,N_16724);
nor U19452 (N_19452,N_15793,N_18221);
or U19453 (N_19453,N_18715,N_17859);
or U19454 (N_19454,N_16696,N_17792);
and U19455 (N_19455,N_18201,N_16213);
xnor U19456 (N_19456,N_16501,N_16438);
or U19457 (N_19457,N_15640,N_16314);
xor U19458 (N_19458,N_18385,N_18581);
nand U19459 (N_19459,N_16029,N_16015);
nor U19460 (N_19460,N_18435,N_15639);
or U19461 (N_19461,N_18273,N_17835);
and U19462 (N_19462,N_16745,N_16840);
nor U19463 (N_19463,N_17939,N_16250);
nand U19464 (N_19464,N_16344,N_15629);
and U19465 (N_19465,N_16886,N_18278);
and U19466 (N_19466,N_16187,N_18488);
or U19467 (N_19467,N_17768,N_18333);
and U19468 (N_19468,N_17028,N_17396);
xnor U19469 (N_19469,N_15689,N_15879);
or U19470 (N_19470,N_16057,N_15633);
nand U19471 (N_19471,N_17104,N_16423);
or U19472 (N_19472,N_16461,N_16965);
nor U19473 (N_19473,N_17247,N_17164);
or U19474 (N_19474,N_18553,N_15951);
or U19475 (N_19475,N_17031,N_18720);
nand U19476 (N_19476,N_15779,N_16189);
or U19477 (N_19477,N_17375,N_16076);
nand U19478 (N_19478,N_17354,N_17525);
xor U19479 (N_19479,N_16791,N_16580);
or U19480 (N_19480,N_15711,N_17272);
and U19481 (N_19481,N_17745,N_16512);
nand U19482 (N_19482,N_15627,N_18481);
or U19483 (N_19483,N_16424,N_17133);
or U19484 (N_19484,N_18248,N_18226);
or U19485 (N_19485,N_17871,N_17238);
or U19486 (N_19486,N_16110,N_16347);
or U19487 (N_19487,N_17888,N_18160);
xnor U19488 (N_19488,N_16629,N_15801);
xnor U19489 (N_19489,N_16035,N_16236);
and U19490 (N_19490,N_16535,N_17640);
nand U19491 (N_19491,N_17002,N_16437);
nor U19492 (N_19492,N_16699,N_17604);
and U19493 (N_19493,N_18416,N_16001);
nor U19494 (N_19494,N_17947,N_17405);
and U19495 (N_19495,N_16754,N_16059);
or U19496 (N_19496,N_18623,N_15864);
xnor U19497 (N_19497,N_16769,N_16369);
nand U19498 (N_19498,N_16371,N_17136);
xnor U19499 (N_19499,N_15760,N_17891);
or U19500 (N_19500,N_17404,N_17412);
xnor U19501 (N_19501,N_18203,N_15707);
xnor U19502 (N_19502,N_18663,N_17660);
nand U19503 (N_19503,N_16856,N_17812);
or U19504 (N_19504,N_17329,N_17817);
or U19505 (N_19505,N_17456,N_17063);
xor U19506 (N_19506,N_16924,N_16094);
nand U19507 (N_19507,N_18182,N_17653);
xor U19508 (N_19508,N_18501,N_16361);
or U19509 (N_19509,N_18426,N_17701);
nand U19510 (N_19510,N_17268,N_18346);
xnor U19511 (N_19511,N_17377,N_18394);
nor U19512 (N_19512,N_16418,N_18665);
nor U19513 (N_19513,N_16383,N_16058);
or U19514 (N_19514,N_18231,N_18655);
xnor U19515 (N_19515,N_18332,N_16752);
or U19516 (N_19516,N_16341,N_17557);
xnor U19517 (N_19517,N_17894,N_17035);
nand U19518 (N_19518,N_17455,N_16633);
nand U19519 (N_19519,N_17281,N_17150);
and U19520 (N_19520,N_18195,N_16910);
or U19521 (N_19521,N_17216,N_17591);
nor U19522 (N_19522,N_17645,N_16643);
nor U19523 (N_19523,N_17262,N_16067);
nor U19524 (N_19524,N_17397,N_15699);
or U19525 (N_19525,N_16925,N_16034);
xnor U19526 (N_19526,N_17457,N_17921);
or U19527 (N_19527,N_18097,N_18646);
or U19528 (N_19528,N_17623,N_16676);
nand U19529 (N_19529,N_18602,N_17408);
nand U19530 (N_19530,N_17400,N_15698);
xor U19531 (N_19531,N_16331,N_17967);
xor U19532 (N_19532,N_16025,N_18564);
xnor U19533 (N_19533,N_15946,N_15681);
nor U19534 (N_19534,N_18075,N_15820);
xor U19535 (N_19535,N_18547,N_18562);
nand U19536 (N_19536,N_16145,N_18522);
and U19537 (N_19537,N_15998,N_16768);
nor U19538 (N_19538,N_15824,N_16073);
or U19539 (N_19539,N_17460,N_18274);
and U19540 (N_19540,N_17234,N_18432);
nor U19541 (N_19541,N_17227,N_16612);
nand U19542 (N_19542,N_16793,N_17169);
nor U19543 (N_19543,N_17481,N_15948);
or U19544 (N_19544,N_17175,N_15834);
nor U19545 (N_19545,N_17673,N_17138);
or U19546 (N_19546,N_17766,N_16421);
nor U19547 (N_19547,N_15923,N_17583);
xor U19548 (N_19548,N_16835,N_16266);
and U19549 (N_19549,N_18404,N_15637);
and U19550 (N_19550,N_16998,N_17204);
nor U19551 (N_19551,N_18372,N_18220);
and U19552 (N_19552,N_17293,N_16349);
nand U19553 (N_19553,N_17407,N_16086);
and U19554 (N_19554,N_17714,N_16534);
nand U19555 (N_19555,N_17161,N_17433);
or U19556 (N_19556,N_18067,N_17439);
xnor U19557 (N_19557,N_16229,N_16400);
nor U19558 (N_19558,N_16800,N_15838);
nor U19559 (N_19559,N_17532,N_16407);
nor U19560 (N_19560,N_16169,N_17836);
and U19561 (N_19561,N_16540,N_18446);
nand U19562 (N_19562,N_16328,N_18275);
or U19563 (N_19563,N_18708,N_16651);
nor U19564 (N_19564,N_18151,N_17316);
nor U19565 (N_19565,N_18452,N_18107);
and U19566 (N_19566,N_18152,N_17185);
nand U19567 (N_19567,N_15945,N_17413);
and U19568 (N_19568,N_16737,N_17108);
xnor U19569 (N_19569,N_16217,N_16674);
and U19570 (N_19570,N_18451,N_15727);
nor U19571 (N_19571,N_18367,N_17914);
xor U19572 (N_19572,N_16738,N_18308);
xor U19573 (N_19573,N_16486,N_18133);
xor U19574 (N_19574,N_16586,N_17128);
nor U19575 (N_19575,N_17476,N_18729);
and U19576 (N_19576,N_18455,N_17450);
nand U19577 (N_19577,N_17672,N_18316);
or U19578 (N_19578,N_18337,N_15867);
nand U19579 (N_19579,N_17542,N_17772);
nand U19580 (N_19580,N_17794,N_18061);
or U19581 (N_19581,N_17417,N_16060);
or U19582 (N_19582,N_16160,N_17139);
and U19583 (N_19583,N_17500,N_15752);
and U19584 (N_19584,N_15874,N_15892);
nand U19585 (N_19585,N_16958,N_18460);
and U19586 (N_19586,N_16749,N_18168);
and U19587 (N_19587,N_17042,N_16671);
nor U19588 (N_19588,N_16658,N_16812);
xnor U19589 (N_19589,N_17411,N_15700);
or U19590 (N_19590,N_16548,N_16061);
or U19591 (N_19591,N_17284,N_15878);
nor U19592 (N_19592,N_15674,N_18741);
nor U19593 (N_19593,N_16309,N_17882);
and U19594 (N_19594,N_15988,N_16493);
xor U19595 (N_19595,N_16043,N_18184);
nand U19596 (N_19596,N_18095,N_18050);
nand U19597 (N_19597,N_17482,N_16916);
xnor U19598 (N_19598,N_17845,N_16019);
nand U19599 (N_19599,N_16928,N_18669);
or U19600 (N_19600,N_18179,N_15690);
nor U19601 (N_19601,N_18321,N_17773);
nor U19602 (N_19602,N_16232,N_16123);
xor U19603 (N_19603,N_16874,N_18215);
and U19604 (N_19604,N_17386,N_16708);
nor U19605 (N_19605,N_17981,N_17177);
nand U19606 (N_19606,N_18487,N_17163);
nand U19607 (N_19607,N_16274,N_18224);
nand U19608 (N_19608,N_16953,N_16247);
nand U19609 (N_19609,N_15912,N_17151);
xor U19610 (N_19610,N_18692,N_16392);
nor U19611 (N_19611,N_17850,N_18538);
xnor U19612 (N_19612,N_18397,N_17016);
nand U19613 (N_19613,N_18223,N_17507);
nor U19614 (N_19614,N_18315,N_16241);
or U19615 (N_19615,N_17877,N_17388);
nor U19616 (N_19616,N_16750,N_16673);
xnor U19617 (N_19617,N_18071,N_15686);
and U19618 (N_19618,N_17277,N_16171);
xor U19619 (N_19619,N_17254,N_16634);
and U19620 (N_19620,N_16249,N_17985);
xnor U19621 (N_19621,N_17627,N_16221);
and U19622 (N_19622,N_17141,N_17732);
xor U19623 (N_19623,N_17734,N_16515);
xnor U19624 (N_19624,N_18494,N_16210);
and U19625 (N_19625,N_16536,N_17067);
nand U19626 (N_19626,N_17336,N_16335);
and U19627 (N_19627,N_16456,N_15885);
nor U19628 (N_19628,N_16397,N_16050);
nand U19629 (N_19629,N_16759,N_16807);
xnor U19630 (N_19630,N_16511,N_16157);
or U19631 (N_19631,N_17937,N_16219);
or U19632 (N_19632,N_16686,N_18502);
xnor U19633 (N_19633,N_18185,N_16485);
nand U19634 (N_19634,N_18474,N_17950);
or U19635 (N_19635,N_16235,N_18083);
and U19636 (N_19636,N_16611,N_16321);
or U19637 (N_19637,N_17590,N_17419);
nand U19638 (N_19638,N_18010,N_16868);
nand U19639 (N_19639,N_16007,N_18266);
nor U19640 (N_19640,N_17382,N_17600);
nor U19641 (N_19641,N_16193,N_17189);
and U19642 (N_19642,N_17721,N_16209);
nand U19643 (N_19643,N_16474,N_16990);
nor U19644 (N_19644,N_15785,N_17844);
or U19645 (N_19645,N_18307,N_15974);
nor U19646 (N_19646,N_17091,N_16429);
and U19647 (N_19647,N_15812,N_18516);
nand U19648 (N_19648,N_17071,N_15980);
nor U19649 (N_19649,N_15899,N_18685);
nor U19650 (N_19650,N_16480,N_16248);
xnor U19651 (N_19651,N_16550,N_16739);
nor U19652 (N_19652,N_17038,N_18305);
nor U19653 (N_19653,N_18430,N_16574);
nor U19654 (N_19654,N_16359,N_17148);
nor U19655 (N_19655,N_17226,N_17255);
nor U19656 (N_19656,N_16806,N_17283);
and U19657 (N_19657,N_16900,N_16039);
and U19658 (N_19658,N_18310,N_16664);
and U19659 (N_19659,N_16571,N_16948);
or U19660 (N_19660,N_16705,N_17906);
and U19661 (N_19661,N_16720,N_16337);
nor U19662 (N_19662,N_16434,N_17472);
and U19663 (N_19663,N_16032,N_15643);
xor U19664 (N_19664,N_16911,N_18718);
xor U19665 (N_19665,N_15994,N_16062);
or U19666 (N_19666,N_17670,N_18150);
nor U19667 (N_19667,N_17860,N_18686);
nand U19668 (N_19668,N_16662,N_16417);
xor U19669 (N_19669,N_16366,N_18389);
or U19670 (N_19670,N_15756,N_16409);
xor U19671 (N_19671,N_16528,N_17300);
xor U19672 (N_19672,N_18131,N_17730);
or U19673 (N_19673,N_18178,N_18382);
or U19674 (N_19674,N_16757,N_17010);
xor U19675 (N_19675,N_17463,N_17055);
and U19676 (N_19676,N_17014,N_17620);
xnor U19677 (N_19677,N_15985,N_15784);
nor U19678 (N_19678,N_18425,N_17948);
or U19679 (N_19679,N_17074,N_16761);
nor U19680 (N_19680,N_16527,N_17271);
and U19681 (N_19681,N_17912,N_18216);
nor U19682 (N_19682,N_18392,N_16357);
nor U19683 (N_19683,N_17176,N_17754);
xor U19684 (N_19684,N_17919,N_17338);
nand U19685 (N_19685,N_16657,N_16547);
or U19686 (N_19686,N_15766,N_16137);
or U19687 (N_19687,N_16151,N_17861);
and U19688 (N_19688,N_17528,N_17371);
nor U19689 (N_19689,N_17326,N_16944);
or U19690 (N_19690,N_18331,N_16289);
nand U19691 (N_19691,N_17702,N_17595);
and U19692 (N_19692,N_17219,N_16999);
nand U19693 (N_19693,N_17895,N_18677);
xor U19694 (N_19694,N_16184,N_16155);
nor U19695 (N_19695,N_16003,N_18594);
and U19696 (N_19696,N_17898,N_17393);
nand U19697 (N_19697,N_17598,N_17260);
and U19698 (N_19698,N_16416,N_16152);
or U19699 (N_19699,N_16707,N_18261);
and U19700 (N_19700,N_16090,N_17729);
xnor U19701 (N_19701,N_16301,N_16441);
xor U19702 (N_19702,N_17474,N_16083);
xor U19703 (N_19703,N_18125,N_18174);
nor U19704 (N_19704,N_17731,N_16297);
nand U19705 (N_19705,N_15962,N_16198);
nand U19706 (N_19706,N_17908,N_15965);
xnor U19707 (N_19707,N_18128,N_15652);
xor U19708 (N_19708,N_16986,N_17809);
or U19709 (N_19709,N_17427,N_18070);
nand U19710 (N_19710,N_17537,N_16728);
nor U19711 (N_19711,N_17220,N_16326);
xnor U19712 (N_19712,N_16293,N_16053);
xor U19713 (N_19713,N_17069,N_17358);
or U19714 (N_19714,N_17757,N_15860);
nor U19715 (N_19715,N_16120,N_15722);
nand U19716 (N_19716,N_15955,N_16952);
or U19717 (N_19717,N_18249,N_17955);
and U19718 (N_19718,N_17572,N_15744);
or U19719 (N_19719,N_16122,N_17129);
nor U19720 (N_19720,N_18351,N_18303);
nand U19721 (N_19721,N_17485,N_16742);
nor U19722 (N_19722,N_16713,N_17099);
nand U19723 (N_19723,N_18296,N_16009);
xor U19724 (N_19724,N_17881,N_16373);
and U19725 (N_19725,N_17297,N_18444);
or U19726 (N_19726,N_16138,N_18207);
xnor U19727 (N_19727,N_18445,N_15981);
nor U19728 (N_19728,N_18604,N_17082);
and U19729 (N_19729,N_16453,N_18238);
nand U19730 (N_19730,N_18189,N_15775);
nand U19731 (N_19731,N_18361,N_18438);
nor U19732 (N_19732,N_18349,N_16934);
nor U19733 (N_19733,N_18484,N_17576);
nand U19734 (N_19734,N_16645,N_17538);
nand U19735 (N_19735,N_15963,N_16778);
or U19736 (N_19736,N_17682,N_17969);
and U19737 (N_19737,N_17639,N_16051);
or U19738 (N_19738,N_16588,N_17357);
xor U19739 (N_19739,N_16408,N_16102);
or U19740 (N_19740,N_17846,N_16508);
xnor U19741 (N_19741,N_18412,N_18116);
xnor U19742 (N_19742,N_16983,N_18497);
xor U19743 (N_19743,N_15929,N_16715);
nor U19744 (N_19744,N_18110,N_17318);
and U19745 (N_19745,N_15886,N_15740);
or U19746 (N_19746,N_18197,N_18714);
nand U19747 (N_19747,N_16147,N_18631);
and U19748 (N_19748,N_15702,N_17636);
nand U19749 (N_19749,N_15846,N_16153);
and U19750 (N_19750,N_18142,N_18377);
and U19751 (N_19751,N_17205,N_17856);
xnor U19752 (N_19752,N_18357,N_16070);
or U19753 (N_19753,N_15668,N_17972);
or U19754 (N_19754,N_17864,N_17295);
and U19755 (N_19755,N_17483,N_18568);
nor U19756 (N_19756,N_17348,N_15819);
nand U19757 (N_19757,N_18544,N_17688);
nor U19758 (N_19758,N_16078,N_17299);
nor U19759 (N_19759,N_16312,N_16109);
xor U19760 (N_19760,N_18515,N_16885);
xor U19761 (N_19761,N_16775,N_16455);
xnor U19762 (N_19762,N_16727,N_16466);
nor U19763 (N_19763,N_18048,N_18365);
and U19764 (N_19764,N_18344,N_15989);
and U19765 (N_19765,N_18407,N_17126);
and U19766 (N_19766,N_16265,N_17414);
nor U19767 (N_19767,N_15881,N_17687);
xor U19768 (N_19768,N_17638,N_16278);
nand U19769 (N_19769,N_17535,N_18567);
xor U19770 (N_19770,N_17622,N_18183);
xor U19771 (N_19771,N_17115,N_16529);
nor U19772 (N_19772,N_18311,N_16544);
nor U19773 (N_19773,N_15810,N_15833);
or U19774 (N_19774,N_15768,N_15688);
nor U19775 (N_19775,N_17484,N_15826);
xnor U19776 (N_19776,N_17061,N_18317);
nor U19777 (N_19777,N_15900,N_17767);
nand U19778 (N_19778,N_18282,N_17458);
nand U19779 (N_19779,N_16272,N_17690);
or U19780 (N_19780,N_15979,N_17885);
nor U19781 (N_19781,N_17241,N_18549);
or U19782 (N_19782,N_15920,N_16450);
and U19783 (N_19783,N_16940,N_16100);
and U19784 (N_19784,N_17486,N_15917);
nor U19785 (N_19785,N_18702,N_16446);
or U19786 (N_19786,N_18120,N_17044);
and U19787 (N_19787,N_17753,N_17305);
or U19788 (N_19788,N_16993,N_18158);
nand U19789 (N_19789,N_17728,N_17246);
nor U19790 (N_19790,N_16028,N_18260);
nand U19791 (N_19791,N_17053,N_17589);
or U19792 (N_19792,N_18738,N_17802);
or U19793 (N_19793,N_18717,N_18104);
nor U19794 (N_19794,N_16828,N_15670);
or U19795 (N_19795,N_17495,N_18625);
nand U19796 (N_19796,N_16860,N_17051);
nor U19797 (N_19797,N_18641,N_18560);
xnor U19798 (N_19798,N_16439,N_15868);
xor U19799 (N_19799,N_16069,N_17868);
or U19800 (N_19800,N_18616,N_16607);
xor U19801 (N_19801,N_17294,N_16435);
nand U19802 (N_19802,N_16154,N_17344);
xnor U19803 (N_19803,N_16799,N_17453);
and U19804 (N_19804,N_17678,N_16813);
and U19805 (N_19805,N_16048,N_17999);
and U19806 (N_19806,N_18388,N_18561);
nand U19807 (N_19807,N_17181,N_17179);
and U19808 (N_19808,N_16382,N_18072);
nand U19809 (N_19809,N_16698,N_15773);
xor U19810 (N_19810,N_18347,N_15993);
and U19811 (N_19811,N_15716,N_18690);
or U19812 (N_19812,N_17076,N_18613);
xor U19813 (N_19813,N_16412,N_17879);
or U19814 (N_19814,N_18524,N_15718);
nor U19815 (N_19815,N_16809,N_18279);
or U19816 (N_19816,N_16307,N_17601);
nor U19817 (N_19817,N_17995,N_16140);
nor U19818 (N_19818,N_18068,N_18667);
nor U19819 (N_19819,N_17425,N_17849);
xor U19820 (N_19820,N_15646,N_18403);
nand U19821 (N_19821,N_17756,N_17068);
and U19822 (N_19822,N_15938,N_17081);
xor U19823 (N_19823,N_15890,N_18615);
xor U19824 (N_19824,N_17709,N_17657);
or U19825 (N_19825,N_16966,N_18681);
nor U19826 (N_19826,N_17765,N_15662);
nand U19827 (N_19827,N_17026,N_17616);
nor U19828 (N_19828,N_17665,N_16510);
and U19829 (N_19829,N_16194,N_16785);
xor U19830 (N_19830,N_18639,N_17345);
xor U19831 (N_19831,N_17852,N_18263);
or U19832 (N_19832,N_17911,N_16804);
and U19833 (N_19833,N_16343,N_17540);
or U19834 (N_19834,N_17703,N_16721);
xor U19835 (N_19835,N_17366,N_15968);
nand U19836 (N_19836,N_17924,N_18472);
nor U19837 (N_19837,N_18578,N_15856);
nand U19838 (N_19838,N_16913,N_18580);
or U19839 (N_19839,N_16258,N_17060);
and U19840 (N_19840,N_18280,N_18548);
nand U19841 (N_19841,N_17901,N_17629);
or U19842 (N_19842,N_16299,N_18088);
and U19843 (N_19843,N_16385,N_17893);
and U19844 (N_19844,N_16669,N_15780);
xnor U19845 (N_19845,N_18609,N_16866);
nand U19846 (N_19846,N_15778,N_18047);
nand U19847 (N_19847,N_17949,N_18600);
nand U19848 (N_19848,N_17127,N_18546);
nor U19849 (N_19849,N_17942,N_15939);
or U19850 (N_19850,N_15759,N_17174);
and U19851 (N_19851,N_17363,N_18709);
or U19852 (N_19852,N_18335,N_18643);
nor U19853 (N_19853,N_16469,N_17564);
xnor U19854 (N_19854,N_18138,N_16099);
and U19855 (N_19855,N_16302,N_15774);
or U19856 (N_19856,N_17073,N_15813);
nor U19857 (N_19857,N_17448,N_16971);
or U19858 (N_19858,N_17248,N_18577);
nor U19859 (N_19859,N_17192,N_17303);
and U19860 (N_19860,N_15918,N_17288);
or U19861 (N_19861,N_16972,N_17403);
nand U19862 (N_19862,N_18473,N_18598);
or U19863 (N_19863,N_16691,N_17222);
xor U19864 (N_19864,N_16315,N_17310);
nor U19865 (N_19865,N_17742,N_17201);
and U19866 (N_19866,N_18073,N_17511);
nor U19867 (N_19867,N_18642,N_17309);
and U19868 (N_19868,N_18584,N_17327);
and U19869 (N_19869,N_18507,N_17931);
nor U19870 (N_19870,N_18724,N_16046);
nand U19871 (N_19871,N_17667,N_18458);
nand U19872 (N_19872,N_16649,N_16648);
or U19873 (N_19873,N_17273,N_16690);
nor U19874 (N_19874,N_17384,N_16054);
or U19875 (N_19875,N_15954,N_16884);
or U19876 (N_19876,N_16994,N_18468);
nor U19877 (N_19877,N_17493,N_17764);
or U19878 (N_19878,N_15806,N_16587);
nand U19879 (N_19879,N_17581,N_17578);
nand U19880 (N_19880,N_16984,N_16789);
nand U19881 (N_19881,N_18402,N_15747);
nand U19882 (N_19882,N_15950,N_18301);
and U19883 (N_19883,N_17118,N_17966);
nor U19884 (N_19884,N_16763,N_17669);
and U19885 (N_19885,N_16037,N_17322);
or U19886 (N_19886,N_18519,N_17079);
or U19887 (N_19887,N_18076,N_17988);
nand U19888 (N_19888,N_17441,N_16968);
or U19889 (N_19889,N_18379,N_17119);
or U19890 (N_19890,N_18707,N_18156);
and U19891 (N_19891,N_17786,N_17243);
nand U19892 (N_19892,N_15657,N_16176);
nand U19893 (N_19893,N_17443,N_16178);
and U19894 (N_19894,N_15797,N_16520);
nor U19895 (N_19895,N_15896,N_16386);
and U19896 (N_19896,N_16545,N_16895);
and U19897 (N_19897,N_17231,N_18537);
and U19898 (N_19898,N_18746,N_17084);
nand U19899 (N_19899,N_16976,N_18592);
and U19900 (N_19900,N_16492,N_15891);
or U19901 (N_19901,N_18103,N_15982);
and U19902 (N_19902,N_15708,N_16149);
or U19903 (N_19903,N_18141,N_18589);
nand U19904 (N_19904,N_17666,N_18020);
and U19905 (N_19905,N_17584,N_16227);
or U19906 (N_19906,N_16118,N_15909);
xor U19907 (N_19907,N_17324,N_15976);
nand U19908 (N_19908,N_17568,N_17499);
nor U19909 (N_19909,N_16195,N_16906);
xnor U19910 (N_19910,N_15913,N_17619);
and U19911 (N_19911,N_17263,N_16834);
and U19912 (N_19912,N_16393,N_18637);
or U19913 (N_19913,N_15903,N_16989);
nor U19914 (N_19914,N_16267,N_17213);
and U19915 (N_19915,N_15787,N_17103);
nand U19916 (N_19916,N_15723,N_17998);
or U19917 (N_19917,N_17781,N_16959);
nor U19918 (N_19918,N_16875,N_17086);
and U19919 (N_19919,N_17896,N_18177);
and U19920 (N_19920,N_16368,N_16719);
and U19921 (N_19921,N_18085,N_18291);
or U19922 (N_19922,N_17203,N_17941);
xnor U19923 (N_19923,N_17372,N_17202);
nor U19924 (N_19924,N_18701,N_16116);
nand U19925 (N_19925,N_15875,N_16594);
and U19926 (N_19926,N_15967,N_16677);
and U19927 (N_19927,N_17697,N_15642);
or U19928 (N_19928,N_16506,N_18748);
or U19929 (N_19929,N_18419,N_17805);
or U19930 (N_19930,N_16234,N_18694);
or U19931 (N_19931,N_18651,N_16722);
or U19932 (N_19932,N_15940,N_18721);
and U19933 (N_19933,N_17801,N_15776);
or U19934 (N_19934,N_18170,N_17459);
and U19935 (N_19935,N_16680,N_17632);
xnor U19936 (N_19936,N_16935,N_18628);
nand U19937 (N_19937,N_18363,N_15695);
and U19938 (N_19938,N_18699,N_15906);
nor U19939 (N_19939,N_17144,N_15858);
xor U19940 (N_19940,N_17544,N_16870);
nand U19941 (N_19941,N_18247,N_17210);
nand U19942 (N_19942,N_17920,N_17699);
xnor U19943 (N_19943,N_18739,N_17249);
nor U19944 (N_19944,N_17719,N_18339);
or U19945 (N_19945,N_18668,N_17015);
or U19946 (N_19946,N_18710,N_16583);
nand U19947 (N_19947,N_17804,N_18605);
xor U19948 (N_19948,N_17530,N_15749);
nor U19949 (N_19949,N_15972,N_17350);
xor U19950 (N_19950,N_16930,N_18493);
xor U19951 (N_19951,N_18033,N_18271);
nand U19952 (N_19952,N_17011,N_17167);
or U19953 (N_19953,N_16732,N_16889);
nand U19954 (N_19954,N_15757,N_16499);
nor U19955 (N_19955,N_18312,N_17613);
and U19956 (N_19956,N_15957,N_18726);
and U19957 (N_19957,N_15783,N_15739);
xor U19958 (N_19958,N_16040,N_15843);
xor U19959 (N_19959,N_16425,N_18209);
nand U19960 (N_19960,N_16186,N_16345);
xnor U19961 (N_19961,N_16353,N_16851);
xnor U19962 (N_19962,N_17555,N_16824);
or U19963 (N_19963,N_16422,N_17264);
xor U19964 (N_19964,N_17218,N_17633);
and U19965 (N_19965,N_17237,N_17521);
or U19966 (N_19966,N_17292,N_17964);
xor U19967 (N_19967,N_15869,N_15732);
nand U19968 (N_19968,N_18236,N_17562);
nor U19969 (N_19969,N_16223,N_15844);
and U19970 (N_19970,N_18566,N_16322);
xnor U19971 (N_19971,N_15777,N_16504);
and U19972 (N_19972,N_17075,N_17579);
xnor U19973 (N_19973,N_17822,N_18653);
or U19974 (N_19974,N_17256,N_17374);
nor U19975 (N_19975,N_17736,N_16872);
nand U19976 (N_19976,N_18442,N_17162);
or U19977 (N_19977,N_18345,N_16861);
or U19978 (N_19978,N_15664,N_18084);
or U19979 (N_19979,N_17810,N_17833);
nor U19980 (N_19980,N_16577,N_15682);
nor U19981 (N_19981,N_16729,N_17567);
nor U19982 (N_19982,N_15731,N_18413);
or U19983 (N_19983,N_18587,N_17778);
and U19984 (N_19984,N_16777,N_16394);
nand U19985 (N_19985,N_16164,N_17373);
nand U19986 (N_19986,N_18725,N_18728);
or U19987 (N_19987,N_18077,N_16609);
nor U19988 (N_19988,N_16743,N_15905);
xor U19989 (N_19989,N_15719,N_18554);
xnor U19990 (N_19990,N_17376,N_18043);
xnor U19991 (N_19991,N_16284,N_15667);
nor U19992 (N_19992,N_17235,N_17929);
and U19993 (N_19993,N_17597,N_18386);
xor U19994 (N_19994,N_18375,N_17692);
nand U19995 (N_19995,N_16771,N_18611);
nor U19996 (N_19996,N_17840,N_18384);
and U19997 (N_19997,N_16822,N_17785);
nor U19998 (N_19998,N_16454,N_18053);
and U19999 (N_19999,N_16324,N_18200);
and U20000 (N_20000,N_18730,N_16685);
and U20001 (N_20001,N_16862,N_17506);
nor U20002 (N_20002,N_15895,N_17351);
and U20003 (N_20003,N_18009,N_15665);
nor U20004 (N_20004,N_18204,N_18028);
nand U20005 (N_20005,N_16770,N_17869);
and U20006 (N_20006,N_16735,N_17651);
xnor U20007 (N_20007,N_16962,N_18327);
nor U20008 (N_20008,N_17658,N_17760);
nand U20009 (N_20009,N_18114,N_17307);
xor U20010 (N_20010,N_17992,N_16105);
or U20011 (N_20011,N_16389,N_18429);
nand U20012 (N_20012,N_17355,N_15724);
or U20013 (N_20013,N_18001,N_15631);
nor U20014 (N_20014,N_18193,N_18051);
nor U20015 (N_20015,N_18422,N_18606);
nor U20016 (N_20016,N_17934,N_18711);
and U20017 (N_20017,N_15889,N_15703);
xor U20018 (N_20018,N_18354,N_18700);
nor U20019 (N_20019,N_17242,N_17510);
or U20020 (N_20020,N_16970,N_18457);
nand U20021 (N_20021,N_18508,N_15684);
nand U20022 (N_20022,N_17990,N_18370);
nand U20023 (N_20023,N_18676,N_18287);
xnor U20024 (N_20024,N_16554,N_17418);
nand U20025 (N_20025,N_17422,N_18599);
xnor U20026 (N_20026,N_17558,N_17392);
and U20027 (N_20027,N_17586,N_17706);
nand U20028 (N_20028,N_18111,N_18252);
xnor U20029 (N_20029,N_18074,N_17505);
nand U20030 (N_20030,N_16327,N_17751);
xnor U20031 (N_20031,N_17737,N_18744);
xor U20032 (N_20032,N_17420,N_16549);
or U20033 (N_20033,N_17984,N_17207);
or U20034 (N_20034,N_18703,N_17899);
or U20035 (N_20035,N_16502,N_17635);
and U20036 (N_20036,N_17124,N_17621);
or U20037 (N_20037,N_18228,N_15764);
and U20038 (N_20038,N_16255,N_18464);
or U20039 (N_20039,N_18060,N_16920);
xnor U20040 (N_20040,N_17873,N_15765);
nand U20041 (N_20041,N_18590,N_15937);
xnor U20042 (N_20042,N_16892,N_15691);
and U20043 (N_20043,N_15847,N_16525);
or U20044 (N_20044,N_18230,N_18591);
nand U20045 (N_20045,N_17788,N_17410);
nand U20046 (N_20046,N_15997,N_16774);
or U20047 (N_20047,N_17858,N_17259);
nand U20048 (N_20048,N_18243,N_17878);
nand U20049 (N_20049,N_18634,N_18205);
nand U20050 (N_20050,N_18059,N_18705);
and U20051 (N_20051,N_17046,N_15746);
and U20052 (N_20052,N_18706,N_16516);
nand U20053 (N_20053,N_18506,N_17634);
nor U20054 (N_20054,N_16142,N_18417);
or U20055 (N_20055,N_18529,N_17782);
and U20056 (N_20056,N_17646,N_16462);
and U20057 (N_20057,N_16098,N_17435);
nor U20058 (N_20058,N_17428,N_18031);
nand U20059 (N_20059,N_15884,N_16891);
and U20060 (N_20060,N_17096,N_16484);
or U20061 (N_20061,N_15877,N_18482);
or U20062 (N_20062,N_16119,N_18719);
or U20063 (N_20063,N_17159,N_16795);
and U20064 (N_20064,N_16413,N_18251);
or U20065 (N_20065,N_16507,N_17454);
and U20066 (N_20066,N_18046,N_16391);
or U20067 (N_20067,N_18005,N_16448);
xor U20068 (N_20068,N_18147,N_17659);
or U20069 (N_20069,N_18042,N_15915);
xor U20070 (N_20070,N_18309,N_17516);
nor U20071 (N_20071,N_17708,N_17494);
xor U20072 (N_20072,N_15818,N_18171);
and U20073 (N_20073,N_18169,N_18096);
nor U20074 (N_20074,N_17594,N_18036);
and U20075 (N_20075,N_17946,N_15769);
nand U20076 (N_20076,N_16841,N_16282);
or U20077 (N_20077,N_15743,N_16553);
nor U20078 (N_20078,N_16604,N_18467);
nand U20079 (N_20079,N_16539,N_17787);
and U20080 (N_20080,N_16096,N_16741);
and U20081 (N_20081,N_15726,N_17251);
xor U20082 (N_20082,N_18353,N_16374);
nor U20083 (N_20083,N_18343,N_17492);
xor U20084 (N_20084,N_17726,N_18727);
xor U20085 (N_20085,N_16279,N_17529);
or U20086 (N_20086,N_17910,N_18341);
nand U20087 (N_20087,N_16350,N_16087);
nand U20088 (N_20088,N_17799,N_15863);
xor U20089 (N_20089,N_18056,N_17296);
nor U20090 (N_20090,N_16902,N_15907);
nor U20091 (N_20091,N_18664,N_16200);
and U20092 (N_20092,N_18149,N_17976);
and U20093 (N_20093,N_17607,N_16091);
or U20094 (N_20094,N_17065,N_18409);
nand U20095 (N_20095,N_16211,N_17656);
xnor U20096 (N_20096,N_18480,N_15669);
nor U20097 (N_20097,N_17698,N_18253);
or U20098 (N_20098,N_15644,N_18069);
or U20099 (N_20099,N_17696,N_16876);
nand U20100 (N_20100,N_17695,N_18362);
xnor U20101 (N_20101,N_18552,N_16794);
nand U20102 (N_20102,N_18424,N_18387);
nand U20103 (N_20103,N_16251,N_18463);
or U20104 (N_20104,N_17502,N_18198);
xor U20105 (N_20105,N_17352,N_18148);
or U20106 (N_20106,N_17642,N_16447);
or U20107 (N_20107,N_17362,N_16589);
and U20108 (N_20108,N_17477,N_18210);
nand U20109 (N_20109,N_16237,N_15680);
and U20110 (N_20110,N_18000,N_18255);
and U20111 (N_20111,N_17206,N_18440);
or U20112 (N_20112,N_16915,N_18607);
nor U20113 (N_20113,N_18418,N_16615);
xnor U20114 (N_20114,N_17746,N_15944);
nor U20115 (N_20115,N_15709,N_17952);
xor U20116 (N_20116,N_18262,N_16240);
and U20117 (N_20117,N_15927,N_18618);
and U20118 (N_20118,N_16403,N_17565);
or U20119 (N_20119,N_17107,N_17225);
and U20120 (N_20120,N_17661,N_17548);
nor U20121 (N_20121,N_15850,N_17954);
xor U20122 (N_20122,N_15832,N_16270);
or U20123 (N_20123,N_18514,N_15753);
nor U20124 (N_20124,N_17052,N_18673);
or U20125 (N_20125,N_16704,N_16095);
nand U20126 (N_20126,N_17024,N_18679);
nand U20127 (N_20127,N_16085,N_17959);
xor U20128 (N_20128,N_17797,N_15762);
and U20129 (N_20129,N_17569,N_18428);
and U20130 (N_20130,N_17496,N_16252);
and U20131 (N_20131,N_18355,N_15663);
nor U20132 (N_20132,N_17135,N_16419);
xnor U20133 (N_20133,N_16973,N_18269);
or U20134 (N_20134,N_16656,N_17674);
xnor U20135 (N_20135,N_17298,N_16026);
or U20136 (N_20136,N_17909,N_17546);
or U20137 (N_20137,N_18202,N_18037);
nand U20138 (N_20138,N_16390,N_17592);
and U20139 (N_20139,N_18237,N_16980);
and U20140 (N_20140,N_17897,N_16479);
and U20141 (N_20141,N_16600,N_17904);
nor U20142 (N_20142,N_17612,N_18597);
nand U20143 (N_20143,N_17199,N_17106);
xor U20144 (N_20144,N_18624,N_18638);
and U20145 (N_20145,N_18233,N_16781);
nor U20146 (N_20146,N_16047,N_17977);
nor U20147 (N_20147,N_16896,N_15653);
or U20148 (N_20148,N_16216,N_18505);
nor U20149 (N_20149,N_17261,N_17137);
or U20150 (N_20150,N_17770,N_16718);
nand U20151 (N_20151,N_18366,N_17596);
xnor U20152 (N_20152,N_16273,N_16610);
nor U20153 (N_20153,N_16395,N_16814);
or U20154 (N_20154,N_16666,N_17574);
and U20155 (N_20155,N_17438,N_18680);
nor U20156 (N_20156,N_16136,N_18017);
nor U20157 (N_20157,N_18129,N_16071);
nor U20158 (N_20158,N_18621,N_18629);
and U20159 (N_20159,N_17987,N_17993);
nor U20160 (N_20160,N_17945,N_18297);
and U20161 (N_20161,N_17994,N_17847);
and U20162 (N_20162,N_18647,N_17331);
nand U20163 (N_20163,N_17796,N_18062);
or U20164 (N_20164,N_16617,N_17957);
nor U20165 (N_20165,N_16488,N_16092);
or U20166 (N_20166,N_18340,N_16358);
xnor U20167 (N_20167,N_17444,N_16080);
and U20168 (N_20168,N_16893,N_18295);
and U20169 (N_20169,N_16979,N_15737);
nor U20170 (N_20170,N_18737,N_16063);
nand U20171 (N_20171,N_17997,N_15947);
and U20172 (N_20172,N_15935,N_17276);
nor U20173 (N_20173,N_17125,N_18348);
nor U20174 (N_20174,N_18684,N_16346);
nand U20175 (N_20175,N_16826,N_16526);
nor U20176 (N_20176,N_17349,N_17320);
nor U20177 (N_20177,N_16954,N_17158);
nor U20178 (N_20178,N_18176,N_17470);
and U20179 (N_20179,N_16517,N_18172);
or U20180 (N_20180,N_17571,N_17747);
and U20181 (N_20181,N_16827,N_16863);
xnor U20182 (N_20182,N_18087,N_16491);
and U20183 (N_20183,N_18635,N_16489);
and U20184 (N_20184,N_18164,N_16882);
and U20185 (N_20185,N_16005,N_17047);
or U20186 (N_20186,N_18081,N_18063);
and U20187 (N_20187,N_18575,N_17704);
and U20188 (N_20188,N_16936,N_17130);
nor U20189 (N_20189,N_17547,N_18235);
xor U20190 (N_20190,N_15908,N_17750);
or U20191 (N_20191,N_18683,N_17269);
xor U20192 (N_20192,N_16277,N_18466);
xnor U20193 (N_20193,N_18420,N_16426);
and U20194 (N_20194,N_16819,N_17963);
or U20195 (N_20195,N_16802,N_17229);
nor U20196 (N_20196,N_15675,N_17884);
nor U20197 (N_20197,N_17637,N_18614);
xor U20198 (N_20198,N_17289,N_15712);
or U20199 (N_20199,N_15697,N_16694);
nand U20200 (N_20200,N_16006,N_18747);
nor U20201 (N_20201,N_17509,N_17606);
nand U20202 (N_20202,N_16964,N_16541);
and U20203 (N_20203,N_16653,N_15836);
and U20204 (N_20204,N_16914,N_18290);
xor U20205 (N_20205,N_17803,N_17471);
or U20206 (N_20206,N_18531,N_16052);
xor U20207 (N_20207,N_17552,N_16388);
nor U20208 (N_20208,N_15671,N_18214);
nor U20209 (N_20209,N_16339,N_18288);
or U20210 (N_20210,N_18644,N_16905);
nand U20211 (N_20211,N_18393,N_17440);
nand U20212 (N_20212,N_16830,N_17267);
xnor U20213 (N_20213,N_16018,N_18500);
or U20214 (N_20214,N_18267,N_16224);
or U20215 (N_20215,N_16912,N_17200);
xor U20216 (N_20216,N_15789,N_15696);
and U20217 (N_20217,N_15754,N_18126);
and U20218 (N_20218,N_17631,N_17744);
nand U20219 (N_20219,N_17398,N_17236);
nor U20220 (N_20220,N_16436,N_18130);
and U20221 (N_20221,N_18636,N_17930);
nand U20222 (N_20222,N_15809,N_16056);
xor U20223 (N_20223,N_17774,N_15804);
xor U20224 (N_20224,N_16716,N_16929);
and U20225 (N_20225,N_18469,N_17821);
nand U20226 (N_20226,N_17526,N_16008);
or U20227 (N_20227,N_18565,N_18232);
or U20228 (N_20228,N_16606,N_18322);
xnor U20229 (N_20229,N_16786,N_18021);
nor U20230 (N_20230,N_17887,N_16156);
xnor U20231 (N_20231,N_17279,N_17779);
xnor U20232 (N_20232,N_17880,N_16779);
xnor U20233 (N_20233,N_15761,N_15829);
and U20234 (N_20234,N_17830,N_17171);
and U20235 (N_20235,N_16445,N_16947);
nor U20236 (N_20236,N_18576,N_16220);
and U20237 (N_20237,N_16784,N_18030);
nor U20238 (N_20238,N_18089,N_16262);
or U20239 (N_20239,N_16564,N_17353);
and U20240 (N_20240,N_16922,N_16228);
xor U20241 (N_20241,N_18257,N_15848);
xnor U20242 (N_20242,N_18013,N_17168);
nand U20243 (N_20243,N_15953,N_17006);
xor U20244 (N_20244,N_18671,N_17986);
nor U20245 (N_20245,N_17971,N_17497);
and U20246 (N_20246,N_18259,N_16873);
and U20247 (N_20247,N_15721,N_18691);
or U20248 (N_20248,N_18246,N_18304);
nor U20249 (N_20249,N_16500,N_16815);
xnor U20250 (N_20250,N_17004,N_16921);
or U20251 (N_20251,N_16338,N_18536);
and U20252 (N_20252,N_17973,N_16848);
nor U20253 (N_20253,N_18433,N_16208);
nand U20254 (N_20254,N_15845,N_16259);
nand U20255 (N_20255,N_17319,N_16477);
nor U20256 (N_20256,N_16700,N_18023);
xnor U20257 (N_20257,N_18503,N_17101);
or U20258 (N_20258,N_17059,N_17449);
or U20259 (N_20259,N_16148,N_17182);
and U20260 (N_20260,N_18563,N_17446);
xor U20261 (N_20261,N_15837,N_16126);
or U20262 (N_20262,N_16808,N_16165);
or U20263 (N_20263,N_18555,N_15687);
xnor U20264 (N_20264,N_16878,N_18190);
nand U20265 (N_20265,N_16376,N_17333);
nor U20266 (N_20266,N_17335,N_17693);
or U20267 (N_20267,N_16538,N_18733);
and U20268 (N_20268,N_16918,N_16712);
nor U20269 (N_20269,N_16561,N_17040);
and U20270 (N_20270,N_17705,N_15758);
or U20271 (N_20271,N_17152,N_17077);
xor U20272 (N_20272,N_18722,N_17286);
and U20273 (N_20273,N_18489,N_15647);
or U20274 (N_20274,N_18155,N_16264);
and U20275 (N_20275,N_17652,N_16597);
nand U20276 (N_20276,N_17671,N_16075);
or U20277 (N_20277,N_18688,N_17602);
and U20278 (N_20278,N_17401,N_18313);
nor U20279 (N_20279,N_17302,N_18292);
xor U20280 (N_20280,N_16846,N_16628);
or U20281 (N_20281,N_17862,N_17208);
and U20282 (N_20282,N_17823,N_17025);
nor U20283 (N_20283,N_17058,N_17716);
or U20284 (N_20284,N_16765,N_16811);
nor U20285 (N_20285,N_16642,N_18106);
and U20286 (N_20286,N_16045,N_17541);
xnor U20287 (N_20287,N_16626,N_16605);
nor U20288 (N_20288,N_18495,N_16858);
and U20289 (N_20289,N_18258,N_18003);
and U20290 (N_20290,N_16991,N_18276);
nand U20291 (N_20291,N_18041,N_17387);
nor U20292 (N_20292,N_16663,N_17105);
nor U20293 (N_20293,N_17686,N_17156);
and U20294 (N_20294,N_16543,N_17436);
nand U20295 (N_20295,N_17048,N_16755);
and U20296 (N_20296,N_17023,N_18441);
nor U20297 (N_20297,N_17585,N_15871);
nor U20298 (N_20298,N_18545,N_15729);
or U20299 (N_20299,N_15802,N_18414);
xor U20300 (N_20300,N_18492,N_17160);
xnor U20301 (N_20301,N_18090,N_16316);
and U20302 (N_20302,N_18496,N_18662);
nor U20303 (N_20303,N_15795,N_17838);
xnor U20304 (N_20304,N_15672,N_16558);
and U20305 (N_20305,N_17360,N_18025);
or U20306 (N_20306,N_17933,N_17343);
or U20307 (N_20307,N_17825,N_18181);
or U20308 (N_20308,N_15781,N_17748);
xor U20309 (N_20309,N_18014,N_15942);
and U20310 (N_20310,N_16206,N_18406);
or U20311 (N_20311,N_17553,N_18029);
nor U20312 (N_20312,N_17818,N_18595);
nand U20313 (N_20313,N_18024,N_17549);
nor U20314 (N_20314,N_17483,N_18355);
xnor U20315 (N_20315,N_16942,N_15931);
and U20316 (N_20316,N_17381,N_18171);
and U20317 (N_20317,N_16833,N_18243);
and U20318 (N_20318,N_16349,N_16310);
or U20319 (N_20319,N_17322,N_17618);
or U20320 (N_20320,N_16427,N_18071);
nand U20321 (N_20321,N_16371,N_17793);
and U20322 (N_20322,N_17274,N_17722);
nor U20323 (N_20323,N_17233,N_16150);
xnor U20324 (N_20324,N_16580,N_15858);
nand U20325 (N_20325,N_17252,N_15951);
nor U20326 (N_20326,N_17926,N_17367);
xnor U20327 (N_20327,N_15701,N_18064);
nor U20328 (N_20328,N_16372,N_16225);
or U20329 (N_20329,N_18602,N_18392);
and U20330 (N_20330,N_18116,N_18666);
nand U20331 (N_20331,N_18442,N_17860);
and U20332 (N_20332,N_18351,N_16008);
or U20333 (N_20333,N_16864,N_17951);
nand U20334 (N_20334,N_16960,N_16886);
or U20335 (N_20335,N_15877,N_17411);
nand U20336 (N_20336,N_18345,N_17777);
xor U20337 (N_20337,N_18550,N_17375);
xnor U20338 (N_20338,N_16454,N_18180);
xnor U20339 (N_20339,N_16711,N_16228);
nand U20340 (N_20340,N_17231,N_17016);
nor U20341 (N_20341,N_18278,N_15806);
xor U20342 (N_20342,N_15973,N_18066);
and U20343 (N_20343,N_17389,N_16068);
xor U20344 (N_20344,N_16190,N_16320);
and U20345 (N_20345,N_18149,N_18478);
nand U20346 (N_20346,N_18510,N_18440);
and U20347 (N_20347,N_18621,N_17040);
and U20348 (N_20348,N_17358,N_15841);
nor U20349 (N_20349,N_18737,N_16842);
nand U20350 (N_20350,N_15843,N_17739);
nand U20351 (N_20351,N_17174,N_18427);
nor U20352 (N_20352,N_18314,N_15775);
or U20353 (N_20353,N_18414,N_15940);
nor U20354 (N_20354,N_16981,N_18332);
xnor U20355 (N_20355,N_18605,N_16608);
and U20356 (N_20356,N_16522,N_17396);
nand U20357 (N_20357,N_17874,N_16973);
and U20358 (N_20358,N_16955,N_16390);
nand U20359 (N_20359,N_17836,N_17418);
xnor U20360 (N_20360,N_16662,N_16789);
xnor U20361 (N_20361,N_15972,N_15653);
or U20362 (N_20362,N_17375,N_15937);
or U20363 (N_20363,N_15713,N_16596);
or U20364 (N_20364,N_16940,N_16638);
nor U20365 (N_20365,N_18619,N_16503);
xor U20366 (N_20366,N_18449,N_16224);
nor U20367 (N_20367,N_18249,N_18484);
and U20368 (N_20368,N_17009,N_17030);
or U20369 (N_20369,N_18420,N_18378);
xnor U20370 (N_20370,N_15642,N_18493);
or U20371 (N_20371,N_18458,N_16686);
nand U20372 (N_20372,N_16997,N_16586);
and U20373 (N_20373,N_18277,N_18615);
nand U20374 (N_20374,N_15967,N_15674);
nor U20375 (N_20375,N_16338,N_18524);
or U20376 (N_20376,N_18437,N_18296);
xor U20377 (N_20377,N_18072,N_18415);
xor U20378 (N_20378,N_18541,N_18488);
and U20379 (N_20379,N_17415,N_17695);
nor U20380 (N_20380,N_16312,N_15637);
or U20381 (N_20381,N_17533,N_18095);
nand U20382 (N_20382,N_17850,N_16983);
xnor U20383 (N_20383,N_17019,N_16482);
nor U20384 (N_20384,N_15974,N_18159);
nand U20385 (N_20385,N_16977,N_16058);
nand U20386 (N_20386,N_16908,N_18116);
or U20387 (N_20387,N_15794,N_16175);
nand U20388 (N_20388,N_18002,N_17097);
nand U20389 (N_20389,N_18299,N_16004);
nand U20390 (N_20390,N_16286,N_15833);
or U20391 (N_20391,N_16290,N_17745);
xnor U20392 (N_20392,N_16823,N_15782);
nand U20393 (N_20393,N_18474,N_17737);
xnor U20394 (N_20394,N_16118,N_18047);
nor U20395 (N_20395,N_17715,N_17244);
nand U20396 (N_20396,N_18118,N_17717);
and U20397 (N_20397,N_17427,N_18077);
and U20398 (N_20398,N_17029,N_17152);
and U20399 (N_20399,N_16127,N_18255);
or U20400 (N_20400,N_18407,N_17292);
nand U20401 (N_20401,N_17196,N_16894);
xnor U20402 (N_20402,N_17649,N_18599);
or U20403 (N_20403,N_15987,N_17130);
or U20404 (N_20404,N_17255,N_17884);
and U20405 (N_20405,N_15865,N_18463);
xor U20406 (N_20406,N_16760,N_17141);
nand U20407 (N_20407,N_16548,N_16809);
nand U20408 (N_20408,N_17315,N_18287);
or U20409 (N_20409,N_16851,N_17243);
and U20410 (N_20410,N_16772,N_18316);
nand U20411 (N_20411,N_16718,N_16036);
nand U20412 (N_20412,N_17623,N_17632);
xor U20413 (N_20413,N_17745,N_17529);
xor U20414 (N_20414,N_18292,N_17693);
nor U20415 (N_20415,N_17432,N_16029);
nand U20416 (N_20416,N_17013,N_18560);
or U20417 (N_20417,N_18217,N_18582);
nand U20418 (N_20418,N_16769,N_18719);
or U20419 (N_20419,N_17455,N_17936);
nor U20420 (N_20420,N_18451,N_17945);
nand U20421 (N_20421,N_18619,N_17879);
or U20422 (N_20422,N_17186,N_17419);
or U20423 (N_20423,N_17654,N_16691);
nand U20424 (N_20424,N_18370,N_16232);
and U20425 (N_20425,N_16384,N_16694);
nor U20426 (N_20426,N_16643,N_18226);
nor U20427 (N_20427,N_16588,N_16883);
nand U20428 (N_20428,N_17987,N_16229);
nor U20429 (N_20429,N_16325,N_15719);
nand U20430 (N_20430,N_18126,N_18160);
or U20431 (N_20431,N_18048,N_16830);
or U20432 (N_20432,N_17851,N_17926);
nor U20433 (N_20433,N_18109,N_17728);
nor U20434 (N_20434,N_16827,N_17771);
and U20435 (N_20435,N_16981,N_18463);
nand U20436 (N_20436,N_17957,N_15951);
xor U20437 (N_20437,N_16057,N_16279);
and U20438 (N_20438,N_18457,N_16033);
nor U20439 (N_20439,N_17730,N_18243);
and U20440 (N_20440,N_17761,N_18449);
and U20441 (N_20441,N_16050,N_18746);
nor U20442 (N_20442,N_18196,N_15634);
and U20443 (N_20443,N_17617,N_17512);
and U20444 (N_20444,N_17623,N_17839);
nor U20445 (N_20445,N_16717,N_15777);
and U20446 (N_20446,N_17215,N_15862);
nor U20447 (N_20447,N_18332,N_16356);
xnor U20448 (N_20448,N_17623,N_17328);
and U20449 (N_20449,N_18737,N_17248);
xor U20450 (N_20450,N_16240,N_15899);
nand U20451 (N_20451,N_17246,N_16548);
or U20452 (N_20452,N_17527,N_17824);
or U20453 (N_20453,N_16127,N_18702);
xnor U20454 (N_20454,N_18502,N_18155);
nand U20455 (N_20455,N_16136,N_18155);
nand U20456 (N_20456,N_16328,N_16232);
nor U20457 (N_20457,N_15922,N_18543);
and U20458 (N_20458,N_18082,N_17352);
or U20459 (N_20459,N_17483,N_15806);
xor U20460 (N_20460,N_18717,N_16505);
or U20461 (N_20461,N_16818,N_15862);
xnor U20462 (N_20462,N_18463,N_17396);
and U20463 (N_20463,N_18710,N_18507);
nor U20464 (N_20464,N_17935,N_18558);
nor U20465 (N_20465,N_18004,N_16171);
and U20466 (N_20466,N_17503,N_17279);
xor U20467 (N_20467,N_16424,N_16951);
or U20468 (N_20468,N_17293,N_18729);
or U20469 (N_20469,N_17151,N_16484);
xnor U20470 (N_20470,N_18576,N_17034);
nor U20471 (N_20471,N_17271,N_18649);
xor U20472 (N_20472,N_16917,N_16705);
nand U20473 (N_20473,N_17973,N_18552);
nand U20474 (N_20474,N_17926,N_17191);
and U20475 (N_20475,N_17804,N_18205);
nor U20476 (N_20476,N_16946,N_16564);
or U20477 (N_20477,N_16556,N_16214);
and U20478 (N_20478,N_15805,N_16263);
nand U20479 (N_20479,N_16442,N_18226);
nor U20480 (N_20480,N_15690,N_17276);
and U20481 (N_20481,N_17244,N_17853);
or U20482 (N_20482,N_17599,N_15646);
or U20483 (N_20483,N_15753,N_16389);
or U20484 (N_20484,N_16403,N_16642);
or U20485 (N_20485,N_18720,N_15869);
or U20486 (N_20486,N_17148,N_16997);
nand U20487 (N_20487,N_17359,N_16477);
or U20488 (N_20488,N_16136,N_17867);
and U20489 (N_20489,N_17848,N_17499);
or U20490 (N_20490,N_16854,N_16792);
xor U20491 (N_20491,N_16837,N_16843);
and U20492 (N_20492,N_17747,N_17358);
xnor U20493 (N_20493,N_17316,N_17873);
xnor U20494 (N_20494,N_18618,N_18224);
or U20495 (N_20495,N_18622,N_17460);
nand U20496 (N_20496,N_16723,N_16370);
or U20497 (N_20497,N_15956,N_16139);
nand U20498 (N_20498,N_16019,N_17247);
nor U20499 (N_20499,N_16122,N_18534);
and U20500 (N_20500,N_18090,N_17286);
nand U20501 (N_20501,N_17295,N_17597);
xor U20502 (N_20502,N_17568,N_17550);
nor U20503 (N_20503,N_17664,N_16289);
nand U20504 (N_20504,N_18643,N_16335);
nand U20505 (N_20505,N_16392,N_16438);
nor U20506 (N_20506,N_17450,N_17456);
or U20507 (N_20507,N_17799,N_16104);
or U20508 (N_20508,N_17374,N_16784);
xor U20509 (N_20509,N_16561,N_18657);
xnor U20510 (N_20510,N_16799,N_17679);
nand U20511 (N_20511,N_15708,N_15867);
or U20512 (N_20512,N_16360,N_18450);
nand U20513 (N_20513,N_16524,N_16949);
nor U20514 (N_20514,N_18146,N_15631);
xor U20515 (N_20515,N_15811,N_17943);
or U20516 (N_20516,N_18699,N_15840);
and U20517 (N_20517,N_18401,N_17643);
nor U20518 (N_20518,N_18622,N_16240);
nor U20519 (N_20519,N_18327,N_16781);
or U20520 (N_20520,N_18415,N_17175);
xnor U20521 (N_20521,N_16881,N_15906);
nor U20522 (N_20522,N_18169,N_17962);
nand U20523 (N_20523,N_15722,N_17170);
nor U20524 (N_20524,N_17750,N_16684);
or U20525 (N_20525,N_15723,N_17111);
nor U20526 (N_20526,N_17784,N_17513);
or U20527 (N_20527,N_16355,N_16498);
nor U20528 (N_20528,N_16426,N_16351);
nand U20529 (N_20529,N_18736,N_16177);
xor U20530 (N_20530,N_15932,N_17824);
nand U20531 (N_20531,N_17578,N_16152);
nor U20532 (N_20532,N_18026,N_18394);
or U20533 (N_20533,N_17185,N_18168);
nor U20534 (N_20534,N_18729,N_17364);
nor U20535 (N_20535,N_15865,N_16328);
nand U20536 (N_20536,N_17850,N_15676);
nor U20537 (N_20537,N_15850,N_18014);
nor U20538 (N_20538,N_16901,N_17404);
xor U20539 (N_20539,N_15759,N_18693);
nand U20540 (N_20540,N_17313,N_17720);
nand U20541 (N_20541,N_18087,N_15757);
nor U20542 (N_20542,N_18647,N_18099);
nor U20543 (N_20543,N_16038,N_17208);
nand U20544 (N_20544,N_18470,N_15801);
or U20545 (N_20545,N_15897,N_16161);
and U20546 (N_20546,N_16726,N_16562);
nand U20547 (N_20547,N_15751,N_16869);
or U20548 (N_20548,N_18417,N_16769);
nor U20549 (N_20549,N_18397,N_16576);
xor U20550 (N_20550,N_17805,N_17253);
and U20551 (N_20551,N_17426,N_18295);
and U20552 (N_20552,N_16142,N_16507);
nor U20553 (N_20553,N_17567,N_16827);
or U20554 (N_20554,N_18041,N_18512);
nor U20555 (N_20555,N_15952,N_17328);
nor U20556 (N_20556,N_17783,N_16120);
and U20557 (N_20557,N_16539,N_16974);
and U20558 (N_20558,N_17986,N_18010);
and U20559 (N_20559,N_17178,N_17263);
and U20560 (N_20560,N_17217,N_17915);
xor U20561 (N_20561,N_16678,N_16747);
or U20562 (N_20562,N_18619,N_17157);
or U20563 (N_20563,N_17258,N_17698);
xnor U20564 (N_20564,N_15838,N_15743);
xor U20565 (N_20565,N_17444,N_16938);
nor U20566 (N_20566,N_17948,N_18460);
xor U20567 (N_20567,N_18098,N_18402);
nand U20568 (N_20568,N_18222,N_16073);
nor U20569 (N_20569,N_15905,N_16858);
xnor U20570 (N_20570,N_16980,N_18048);
nand U20571 (N_20571,N_16220,N_16137);
and U20572 (N_20572,N_17520,N_17176);
and U20573 (N_20573,N_17505,N_18142);
nand U20574 (N_20574,N_15768,N_18281);
and U20575 (N_20575,N_18130,N_17764);
nor U20576 (N_20576,N_17598,N_17578);
xor U20577 (N_20577,N_16187,N_16438);
xor U20578 (N_20578,N_18502,N_16054);
nor U20579 (N_20579,N_18354,N_16441);
xor U20580 (N_20580,N_17817,N_17896);
nor U20581 (N_20581,N_17142,N_17793);
and U20582 (N_20582,N_17856,N_17708);
and U20583 (N_20583,N_18098,N_15932);
nand U20584 (N_20584,N_17704,N_16877);
xnor U20585 (N_20585,N_16508,N_16269);
or U20586 (N_20586,N_17565,N_16601);
nand U20587 (N_20587,N_17044,N_17736);
nor U20588 (N_20588,N_17821,N_18670);
or U20589 (N_20589,N_16963,N_15876);
or U20590 (N_20590,N_16618,N_18188);
nor U20591 (N_20591,N_16275,N_16788);
and U20592 (N_20592,N_17732,N_17632);
xor U20593 (N_20593,N_16147,N_16329);
nor U20594 (N_20594,N_16619,N_16779);
or U20595 (N_20595,N_16132,N_17012);
xnor U20596 (N_20596,N_18415,N_17501);
xor U20597 (N_20597,N_17423,N_17403);
or U20598 (N_20598,N_16062,N_16082);
and U20599 (N_20599,N_16414,N_18237);
nand U20600 (N_20600,N_17403,N_16874);
or U20601 (N_20601,N_17498,N_18659);
and U20602 (N_20602,N_17709,N_17446);
xor U20603 (N_20603,N_16049,N_18341);
nand U20604 (N_20604,N_17770,N_17794);
or U20605 (N_20605,N_15824,N_18130);
nand U20606 (N_20606,N_17290,N_17142);
and U20607 (N_20607,N_17281,N_17543);
and U20608 (N_20608,N_17880,N_17210);
nand U20609 (N_20609,N_17510,N_16211);
nand U20610 (N_20610,N_18736,N_17184);
and U20611 (N_20611,N_18540,N_16739);
or U20612 (N_20612,N_18659,N_17229);
nor U20613 (N_20613,N_16924,N_17747);
or U20614 (N_20614,N_17369,N_18047);
xnor U20615 (N_20615,N_17663,N_17158);
nand U20616 (N_20616,N_17619,N_15699);
xnor U20617 (N_20617,N_16915,N_15673);
xnor U20618 (N_20618,N_18196,N_17290);
and U20619 (N_20619,N_16852,N_15887);
and U20620 (N_20620,N_15793,N_17630);
and U20621 (N_20621,N_16512,N_16366);
or U20622 (N_20622,N_18531,N_17689);
nor U20623 (N_20623,N_17789,N_15841);
nor U20624 (N_20624,N_16838,N_17952);
or U20625 (N_20625,N_17876,N_17614);
and U20626 (N_20626,N_18539,N_18680);
and U20627 (N_20627,N_15799,N_16788);
nor U20628 (N_20628,N_16240,N_16670);
xor U20629 (N_20629,N_18040,N_16352);
and U20630 (N_20630,N_17287,N_18635);
nand U20631 (N_20631,N_18258,N_17338);
and U20632 (N_20632,N_17867,N_17002);
xnor U20633 (N_20633,N_18115,N_17933);
and U20634 (N_20634,N_16927,N_16470);
xnor U20635 (N_20635,N_17085,N_18731);
nand U20636 (N_20636,N_17881,N_16745);
xnor U20637 (N_20637,N_17942,N_16652);
or U20638 (N_20638,N_16233,N_16119);
xnor U20639 (N_20639,N_17208,N_18638);
or U20640 (N_20640,N_15725,N_16182);
or U20641 (N_20641,N_17336,N_17785);
and U20642 (N_20642,N_16908,N_16620);
nor U20643 (N_20643,N_17530,N_17401);
nor U20644 (N_20644,N_18671,N_17379);
and U20645 (N_20645,N_18288,N_15931);
and U20646 (N_20646,N_18165,N_16792);
and U20647 (N_20647,N_18719,N_18160);
and U20648 (N_20648,N_16394,N_16959);
and U20649 (N_20649,N_17897,N_17837);
or U20650 (N_20650,N_17964,N_17028);
and U20651 (N_20651,N_18266,N_15979);
and U20652 (N_20652,N_16185,N_17867);
nand U20653 (N_20653,N_15996,N_16377);
nand U20654 (N_20654,N_16108,N_17032);
nor U20655 (N_20655,N_17368,N_16370);
xor U20656 (N_20656,N_17610,N_18636);
xor U20657 (N_20657,N_16261,N_16802);
or U20658 (N_20658,N_17922,N_18058);
xnor U20659 (N_20659,N_16494,N_16646);
and U20660 (N_20660,N_15925,N_18294);
xnor U20661 (N_20661,N_18083,N_16658);
or U20662 (N_20662,N_17655,N_18449);
nor U20663 (N_20663,N_18595,N_17572);
nor U20664 (N_20664,N_18518,N_16684);
and U20665 (N_20665,N_17385,N_16213);
xor U20666 (N_20666,N_16437,N_17055);
nor U20667 (N_20667,N_18643,N_17943);
or U20668 (N_20668,N_18563,N_16174);
and U20669 (N_20669,N_17427,N_15760);
xnor U20670 (N_20670,N_17348,N_17498);
nor U20671 (N_20671,N_17671,N_17487);
or U20672 (N_20672,N_17891,N_16112);
or U20673 (N_20673,N_18147,N_18469);
or U20674 (N_20674,N_16448,N_17726);
xnor U20675 (N_20675,N_17321,N_18381);
and U20676 (N_20676,N_18628,N_16163);
xor U20677 (N_20677,N_16687,N_15691);
xnor U20678 (N_20678,N_18007,N_17284);
and U20679 (N_20679,N_17244,N_15947);
xor U20680 (N_20680,N_15663,N_17615);
or U20681 (N_20681,N_15870,N_17027);
and U20682 (N_20682,N_17041,N_16062);
and U20683 (N_20683,N_15994,N_17312);
and U20684 (N_20684,N_17271,N_17779);
nor U20685 (N_20685,N_17594,N_16434);
and U20686 (N_20686,N_16034,N_18714);
xor U20687 (N_20687,N_18391,N_18417);
nand U20688 (N_20688,N_17485,N_18508);
xor U20689 (N_20689,N_16405,N_17200);
xnor U20690 (N_20690,N_16558,N_15893);
nor U20691 (N_20691,N_15870,N_15833);
or U20692 (N_20692,N_17947,N_17071);
and U20693 (N_20693,N_18369,N_16854);
nor U20694 (N_20694,N_15808,N_15872);
nand U20695 (N_20695,N_16290,N_18191);
and U20696 (N_20696,N_18041,N_17659);
xor U20697 (N_20697,N_17962,N_18232);
nor U20698 (N_20698,N_15647,N_17213);
nor U20699 (N_20699,N_18163,N_16309);
or U20700 (N_20700,N_16728,N_17059);
xnor U20701 (N_20701,N_16005,N_16527);
nand U20702 (N_20702,N_17253,N_15938);
nor U20703 (N_20703,N_16515,N_17748);
nor U20704 (N_20704,N_18196,N_17138);
xor U20705 (N_20705,N_18742,N_18210);
nand U20706 (N_20706,N_16845,N_16939);
xor U20707 (N_20707,N_18748,N_16016);
and U20708 (N_20708,N_17840,N_18351);
and U20709 (N_20709,N_18653,N_18714);
or U20710 (N_20710,N_18178,N_16180);
xor U20711 (N_20711,N_18178,N_16304);
nand U20712 (N_20712,N_16090,N_18150);
xor U20713 (N_20713,N_15779,N_17230);
nand U20714 (N_20714,N_16776,N_16909);
xor U20715 (N_20715,N_17883,N_16069);
nor U20716 (N_20716,N_17037,N_16378);
and U20717 (N_20717,N_17629,N_18176);
xor U20718 (N_20718,N_18382,N_18385);
nand U20719 (N_20719,N_16121,N_17794);
and U20720 (N_20720,N_16134,N_18386);
or U20721 (N_20721,N_17322,N_17414);
or U20722 (N_20722,N_17634,N_17894);
xor U20723 (N_20723,N_18541,N_18173);
xnor U20724 (N_20724,N_18490,N_18112);
xnor U20725 (N_20725,N_18697,N_16372);
nor U20726 (N_20726,N_17283,N_16003);
nand U20727 (N_20727,N_16325,N_17692);
nor U20728 (N_20728,N_18274,N_16181);
and U20729 (N_20729,N_16466,N_17214);
or U20730 (N_20730,N_18585,N_15643);
nand U20731 (N_20731,N_17109,N_16073);
nor U20732 (N_20732,N_17259,N_16249);
xnor U20733 (N_20733,N_17032,N_16647);
nor U20734 (N_20734,N_18567,N_17209);
nor U20735 (N_20735,N_17575,N_17564);
nand U20736 (N_20736,N_18084,N_18670);
and U20737 (N_20737,N_18133,N_16724);
xor U20738 (N_20738,N_16574,N_18737);
or U20739 (N_20739,N_18119,N_18611);
nand U20740 (N_20740,N_16389,N_16900);
nor U20741 (N_20741,N_17431,N_18185);
nand U20742 (N_20742,N_17771,N_16683);
nor U20743 (N_20743,N_18506,N_16843);
and U20744 (N_20744,N_18000,N_17360);
nand U20745 (N_20745,N_17378,N_17410);
or U20746 (N_20746,N_17142,N_17533);
or U20747 (N_20747,N_18250,N_18209);
xnor U20748 (N_20748,N_16932,N_16044);
xnor U20749 (N_20749,N_16616,N_18671);
and U20750 (N_20750,N_16204,N_17397);
xor U20751 (N_20751,N_18495,N_16341);
or U20752 (N_20752,N_16154,N_18602);
or U20753 (N_20753,N_17128,N_18398);
or U20754 (N_20754,N_16111,N_15871);
nand U20755 (N_20755,N_16007,N_15794);
nand U20756 (N_20756,N_18524,N_17483);
or U20757 (N_20757,N_17123,N_16111);
nand U20758 (N_20758,N_16757,N_16989);
or U20759 (N_20759,N_16537,N_17247);
nor U20760 (N_20760,N_18082,N_17861);
xor U20761 (N_20761,N_16204,N_16261);
and U20762 (N_20762,N_17160,N_16684);
nand U20763 (N_20763,N_17663,N_16265);
xor U20764 (N_20764,N_16817,N_18024);
nor U20765 (N_20765,N_18385,N_18295);
nand U20766 (N_20766,N_17486,N_15963);
or U20767 (N_20767,N_18088,N_17699);
xnor U20768 (N_20768,N_17041,N_17982);
nand U20769 (N_20769,N_16413,N_16310);
or U20770 (N_20770,N_15743,N_17513);
and U20771 (N_20771,N_17650,N_16982);
or U20772 (N_20772,N_17418,N_17522);
and U20773 (N_20773,N_16628,N_16103);
nor U20774 (N_20774,N_17330,N_16236);
or U20775 (N_20775,N_17777,N_16342);
xnor U20776 (N_20776,N_18097,N_16835);
nor U20777 (N_20777,N_17818,N_16655);
or U20778 (N_20778,N_16218,N_16708);
or U20779 (N_20779,N_17942,N_15814);
nor U20780 (N_20780,N_18553,N_16559);
nor U20781 (N_20781,N_17571,N_18104);
xnor U20782 (N_20782,N_17434,N_17766);
xor U20783 (N_20783,N_16021,N_17522);
nand U20784 (N_20784,N_18099,N_17655);
nand U20785 (N_20785,N_18118,N_16406);
nor U20786 (N_20786,N_16713,N_16223);
nand U20787 (N_20787,N_17286,N_16661);
and U20788 (N_20788,N_17747,N_16315);
xnor U20789 (N_20789,N_18041,N_15902);
or U20790 (N_20790,N_18235,N_18148);
nand U20791 (N_20791,N_16309,N_16096);
xnor U20792 (N_20792,N_18479,N_17660);
nand U20793 (N_20793,N_17018,N_17732);
xor U20794 (N_20794,N_17217,N_17913);
and U20795 (N_20795,N_17831,N_16115);
and U20796 (N_20796,N_16101,N_16651);
or U20797 (N_20797,N_15846,N_16341);
xor U20798 (N_20798,N_18453,N_17698);
and U20799 (N_20799,N_17283,N_17285);
nor U20800 (N_20800,N_16707,N_18281);
nor U20801 (N_20801,N_16143,N_16449);
nor U20802 (N_20802,N_18571,N_18063);
nor U20803 (N_20803,N_17307,N_16699);
xor U20804 (N_20804,N_16921,N_16841);
nor U20805 (N_20805,N_16515,N_17512);
nor U20806 (N_20806,N_16530,N_18388);
xor U20807 (N_20807,N_16011,N_18475);
and U20808 (N_20808,N_16165,N_17577);
xnor U20809 (N_20809,N_16923,N_15667);
nor U20810 (N_20810,N_16715,N_16436);
nor U20811 (N_20811,N_16643,N_16525);
nor U20812 (N_20812,N_15922,N_15923);
and U20813 (N_20813,N_16371,N_18277);
xnor U20814 (N_20814,N_18201,N_17920);
or U20815 (N_20815,N_17688,N_16980);
or U20816 (N_20816,N_16491,N_17057);
xor U20817 (N_20817,N_15993,N_16583);
xor U20818 (N_20818,N_16465,N_16893);
xor U20819 (N_20819,N_17275,N_18626);
nand U20820 (N_20820,N_16309,N_16492);
xor U20821 (N_20821,N_17930,N_17340);
xnor U20822 (N_20822,N_16562,N_18084);
and U20823 (N_20823,N_17305,N_18326);
and U20824 (N_20824,N_17014,N_16005);
and U20825 (N_20825,N_18466,N_17621);
nand U20826 (N_20826,N_17036,N_18012);
or U20827 (N_20827,N_16730,N_16236);
nor U20828 (N_20828,N_18343,N_17507);
xnor U20829 (N_20829,N_18624,N_16974);
nor U20830 (N_20830,N_16337,N_18647);
and U20831 (N_20831,N_15699,N_16371);
and U20832 (N_20832,N_16762,N_17304);
or U20833 (N_20833,N_17591,N_17558);
xnor U20834 (N_20834,N_16050,N_16000);
nand U20835 (N_20835,N_18133,N_17264);
and U20836 (N_20836,N_18512,N_18186);
and U20837 (N_20837,N_16222,N_18192);
or U20838 (N_20838,N_18521,N_16439);
or U20839 (N_20839,N_16923,N_17138);
and U20840 (N_20840,N_17982,N_17121);
or U20841 (N_20841,N_18736,N_17867);
xor U20842 (N_20842,N_17170,N_17697);
nor U20843 (N_20843,N_17568,N_16707);
xor U20844 (N_20844,N_18003,N_17798);
nor U20845 (N_20845,N_16516,N_17098);
or U20846 (N_20846,N_18600,N_16652);
nor U20847 (N_20847,N_18028,N_17718);
and U20848 (N_20848,N_15925,N_17367);
and U20849 (N_20849,N_18011,N_16854);
or U20850 (N_20850,N_18072,N_17494);
and U20851 (N_20851,N_18332,N_15865);
or U20852 (N_20852,N_17239,N_18314);
nand U20853 (N_20853,N_17420,N_16116);
nor U20854 (N_20854,N_16002,N_17223);
or U20855 (N_20855,N_15786,N_17509);
nor U20856 (N_20856,N_17057,N_16675);
nor U20857 (N_20857,N_16218,N_17720);
nor U20858 (N_20858,N_18405,N_17627);
nor U20859 (N_20859,N_17655,N_18638);
and U20860 (N_20860,N_17664,N_18499);
and U20861 (N_20861,N_17761,N_18386);
xor U20862 (N_20862,N_17901,N_17861);
nand U20863 (N_20863,N_17180,N_18683);
nand U20864 (N_20864,N_17206,N_17092);
or U20865 (N_20865,N_17924,N_18198);
and U20866 (N_20866,N_17995,N_16954);
nand U20867 (N_20867,N_16026,N_18073);
or U20868 (N_20868,N_16278,N_17171);
nor U20869 (N_20869,N_16974,N_18647);
nor U20870 (N_20870,N_16864,N_17846);
or U20871 (N_20871,N_16245,N_18529);
or U20872 (N_20872,N_17350,N_16827);
xnor U20873 (N_20873,N_17732,N_17822);
or U20874 (N_20874,N_18373,N_18024);
nor U20875 (N_20875,N_17308,N_16189);
xor U20876 (N_20876,N_17299,N_15698);
nand U20877 (N_20877,N_18328,N_18143);
and U20878 (N_20878,N_16786,N_17087);
and U20879 (N_20879,N_18630,N_16985);
nor U20880 (N_20880,N_18189,N_18412);
nor U20881 (N_20881,N_16680,N_16493);
xnor U20882 (N_20882,N_16887,N_17329);
or U20883 (N_20883,N_17869,N_18394);
nand U20884 (N_20884,N_17408,N_15979);
nand U20885 (N_20885,N_16222,N_17455);
xnor U20886 (N_20886,N_18454,N_16022);
xor U20887 (N_20887,N_18534,N_16794);
or U20888 (N_20888,N_18184,N_17306);
nand U20889 (N_20889,N_16280,N_16482);
nor U20890 (N_20890,N_17593,N_16097);
nor U20891 (N_20891,N_16818,N_15741);
or U20892 (N_20892,N_17309,N_15851);
nor U20893 (N_20893,N_17504,N_17747);
or U20894 (N_20894,N_16927,N_16435);
xor U20895 (N_20895,N_17705,N_16068);
or U20896 (N_20896,N_17478,N_17320);
nand U20897 (N_20897,N_17045,N_16289);
nor U20898 (N_20898,N_18605,N_16265);
or U20899 (N_20899,N_17717,N_17246);
nor U20900 (N_20900,N_16070,N_16284);
nand U20901 (N_20901,N_18036,N_16007);
or U20902 (N_20902,N_15940,N_16339);
nor U20903 (N_20903,N_15701,N_18176);
and U20904 (N_20904,N_17464,N_17877);
nor U20905 (N_20905,N_18045,N_17299);
nor U20906 (N_20906,N_17654,N_17220);
and U20907 (N_20907,N_16729,N_17324);
nand U20908 (N_20908,N_15899,N_18338);
and U20909 (N_20909,N_17019,N_17694);
or U20910 (N_20910,N_18443,N_17518);
nor U20911 (N_20911,N_16605,N_17880);
nor U20912 (N_20912,N_18659,N_17883);
nor U20913 (N_20913,N_18296,N_17659);
xnor U20914 (N_20914,N_16423,N_17478);
or U20915 (N_20915,N_16305,N_18114);
nand U20916 (N_20916,N_16916,N_16519);
nor U20917 (N_20917,N_18389,N_15807);
xor U20918 (N_20918,N_18155,N_18128);
nand U20919 (N_20919,N_16607,N_17711);
nor U20920 (N_20920,N_17640,N_17800);
xor U20921 (N_20921,N_17768,N_18316);
nor U20922 (N_20922,N_17031,N_18002);
and U20923 (N_20923,N_18131,N_16147);
nand U20924 (N_20924,N_16755,N_17088);
and U20925 (N_20925,N_17289,N_18037);
nor U20926 (N_20926,N_18431,N_16749);
nor U20927 (N_20927,N_16862,N_18500);
nand U20928 (N_20928,N_16156,N_18670);
nor U20929 (N_20929,N_18652,N_16087);
nor U20930 (N_20930,N_18729,N_17307);
or U20931 (N_20931,N_16191,N_16865);
or U20932 (N_20932,N_17046,N_17995);
nor U20933 (N_20933,N_18511,N_15666);
xnor U20934 (N_20934,N_18435,N_15931);
nor U20935 (N_20935,N_17516,N_17953);
nand U20936 (N_20936,N_16901,N_18571);
nand U20937 (N_20937,N_16531,N_16130);
xor U20938 (N_20938,N_16311,N_17933);
nor U20939 (N_20939,N_17816,N_16356);
and U20940 (N_20940,N_16365,N_17180);
nand U20941 (N_20941,N_16206,N_17934);
xnor U20942 (N_20942,N_15688,N_18197);
or U20943 (N_20943,N_16031,N_17733);
or U20944 (N_20944,N_17773,N_16908);
or U20945 (N_20945,N_17696,N_17689);
nand U20946 (N_20946,N_18181,N_17886);
or U20947 (N_20947,N_17780,N_17026);
or U20948 (N_20948,N_18191,N_16737);
xor U20949 (N_20949,N_16810,N_18128);
nor U20950 (N_20950,N_16123,N_17519);
nand U20951 (N_20951,N_16924,N_15974);
or U20952 (N_20952,N_17556,N_16850);
nand U20953 (N_20953,N_18040,N_17419);
or U20954 (N_20954,N_18264,N_16711);
or U20955 (N_20955,N_15753,N_17469);
nor U20956 (N_20956,N_17611,N_18696);
nor U20957 (N_20957,N_15628,N_17784);
or U20958 (N_20958,N_16581,N_17112);
xor U20959 (N_20959,N_17041,N_16313);
or U20960 (N_20960,N_17770,N_15806);
nor U20961 (N_20961,N_17581,N_18523);
nor U20962 (N_20962,N_16344,N_16660);
xnor U20963 (N_20963,N_16332,N_18039);
nand U20964 (N_20964,N_16223,N_16930);
or U20965 (N_20965,N_18723,N_18227);
and U20966 (N_20966,N_18649,N_18719);
nand U20967 (N_20967,N_16257,N_16059);
or U20968 (N_20968,N_18189,N_15879);
nor U20969 (N_20969,N_16009,N_17521);
nor U20970 (N_20970,N_16940,N_16943);
and U20971 (N_20971,N_17367,N_16313);
nand U20972 (N_20972,N_16201,N_17939);
nand U20973 (N_20973,N_16347,N_16787);
xor U20974 (N_20974,N_18220,N_17195);
nand U20975 (N_20975,N_17617,N_18128);
nand U20976 (N_20976,N_16105,N_18699);
nand U20977 (N_20977,N_18489,N_17789);
or U20978 (N_20978,N_17615,N_17254);
and U20979 (N_20979,N_17850,N_17306);
nor U20980 (N_20980,N_16122,N_18120);
xor U20981 (N_20981,N_16891,N_16098);
and U20982 (N_20982,N_18300,N_17873);
nand U20983 (N_20983,N_15868,N_16537);
xor U20984 (N_20984,N_17926,N_16377);
nor U20985 (N_20985,N_15698,N_17519);
nand U20986 (N_20986,N_18582,N_16441);
nor U20987 (N_20987,N_18423,N_17644);
and U20988 (N_20988,N_17306,N_16080);
nor U20989 (N_20989,N_17606,N_17056);
and U20990 (N_20990,N_18563,N_17282);
nor U20991 (N_20991,N_16263,N_16065);
xor U20992 (N_20992,N_18378,N_18700);
nand U20993 (N_20993,N_15668,N_16523);
nand U20994 (N_20994,N_17799,N_16931);
or U20995 (N_20995,N_15852,N_17024);
xor U20996 (N_20996,N_16036,N_16511);
and U20997 (N_20997,N_16286,N_18299);
xnor U20998 (N_20998,N_15940,N_17336);
nand U20999 (N_20999,N_15741,N_15967);
and U21000 (N_21000,N_17303,N_17564);
nor U21001 (N_21001,N_17045,N_16473);
nor U21002 (N_21002,N_17608,N_15627);
or U21003 (N_21003,N_15694,N_16155);
or U21004 (N_21004,N_16594,N_17732);
or U21005 (N_21005,N_18455,N_17418);
and U21006 (N_21006,N_17181,N_18715);
nand U21007 (N_21007,N_16064,N_17362);
nand U21008 (N_21008,N_15960,N_17979);
or U21009 (N_21009,N_16469,N_18204);
nand U21010 (N_21010,N_16981,N_16134);
nand U21011 (N_21011,N_16799,N_18471);
or U21012 (N_21012,N_18197,N_18239);
and U21013 (N_21013,N_18585,N_16305);
xnor U21014 (N_21014,N_17798,N_17831);
or U21015 (N_21015,N_17950,N_15900);
nor U21016 (N_21016,N_16936,N_16198);
xor U21017 (N_21017,N_16312,N_16776);
nor U21018 (N_21018,N_16382,N_17321);
or U21019 (N_21019,N_18022,N_17703);
xor U21020 (N_21020,N_16460,N_15969);
and U21021 (N_21021,N_17184,N_17928);
nand U21022 (N_21022,N_17556,N_18469);
and U21023 (N_21023,N_15958,N_16299);
nor U21024 (N_21024,N_16405,N_17332);
and U21025 (N_21025,N_16554,N_18536);
and U21026 (N_21026,N_16881,N_16105);
xor U21027 (N_21027,N_18071,N_15709);
nor U21028 (N_21028,N_17641,N_18411);
or U21029 (N_21029,N_18255,N_17091);
xor U21030 (N_21030,N_16480,N_15929);
and U21031 (N_21031,N_15960,N_18688);
and U21032 (N_21032,N_15858,N_17442);
nand U21033 (N_21033,N_17558,N_16150);
or U21034 (N_21034,N_15757,N_16467);
nand U21035 (N_21035,N_17193,N_16718);
nand U21036 (N_21036,N_17008,N_18229);
and U21037 (N_21037,N_15972,N_17458);
xnor U21038 (N_21038,N_18088,N_17912);
nor U21039 (N_21039,N_16450,N_18171);
nor U21040 (N_21040,N_16902,N_15626);
and U21041 (N_21041,N_15968,N_17621);
xnor U21042 (N_21042,N_17959,N_16790);
or U21043 (N_21043,N_18264,N_18492);
or U21044 (N_21044,N_17656,N_18072);
nor U21045 (N_21045,N_16963,N_15850);
nor U21046 (N_21046,N_15982,N_15642);
nand U21047 (N_21047,N_16684,N_15639);
nand U21048 (N_21048,N_16097,N_18453);
and U21049 (N_21049,N_16046,N_15682);
nand U21050 (N_21050,N_18423,N_17370);
nand U21051 (N_21051,N_18735,N_17119);
and U21052 (N_21052,N_16396,N_17461);
and U21053 (N_21053,N_17270,N_18667);
nor U21054 (N_21054,N_17797,N_17218);
nand U21055 (N_21055,N_18294,N_18252);
or U21056 (N_21056,N_16098,N_18713);
xor U21057 (N_21057,N_18123,N_16664);
xnor U21058 (N_21058,N_17225,N_16299);
nor U21059 (N_21059,N_16560,N_16802);
nand U21060 (N_21060,N_18341,N_17258);
and U21061 (N_21061,N_17391,N_16907);
or U21062 (N_21062,N_18721,N_15988);
nor U21063 (N_21063,N_17308,N_16635);
xor U21064 (N_21064,N_17624,N_18306);
and U21065 (N_21065,N_17227,N_16656);
nor U21066 (N_21066,N_17992,N_17695);
nor U21067 (N_21067,N_17396,N_17234);
xnor U21068 (N_21068,N_16513,N_16409);
and U21069 (N_21069,N_15723,N_18080);
and U21070 (N_21070,N_16178,N_16967);
nor U21071 (N_21071,N_18609,N_16468);
xnor U21072 (N_21072,N_16159,N_18244);
and U21073 (N_21073,N_16194,N_17719);
xor U21074 (N_21074,N_16326,N_15850);
nor U21075 (N_21075,N_17450,N_17069);
nand U21076 (N_21076,N_17351,N_16906);
xor U21077 (N_21077,N_17134,N_18008);
nand U21078 (N_21078,N_15953,N_17464);
or U21079 (N_21079,N_17072,N_18288);
and U21080 (N_21080,N_16672,N_16688);
xnor U21081 (N_21081,N_17883,N_18541);
or U21082 (N_21082,N_18448,N_16279);
and U21083 (N_21083,N_17894,N_16066);
xnor U21084 (N_21084,N_16494,N_17058);
nand U21085 (N_21085,N_16559,N_16563);
or U21086 (N_21086,N_17981,N_17107);
or U21087 (N_21087,N_18597,N_15918);
nand U21088 (N_21088,N_18698,N_15698);
and U21089 (N_21089,N_17641,N_15814);
and U21090 (N_21090,N_16147,N_16536);
xor U21091 (N_21091,N_15813,N_18498);
and U21092 (N_21092,N_18613,N_18412);
nor U21093 (N_21093,N_16207,N_17598);
nand U21094 (N_21094,N_16950,N_16345);
nor U21095 (N_21095,N_18092,N_15822);
xnor U21096 (N_21096,N_17407,N_16925);
or U21097 (N_21097,N_18533,N_16896);
xor U21098 (N_21098,N_18096,N_17982);
or U21099 (N_21099,N_17153,N_17203);
nand U21100 (N_21100,N_18734,N_18113);
and U21101 (N_21101,N_17054,N_18501);
xnor U21102 (N_21102,N_17019,N_17741);
nand U21103 (N_21103,N_18236,N_15742);
or U21104 (N_21104,N_15988,N_18166);
nor U21105 (N_21105,N_18197,N_16231);
xnor U21106 (N_21106,N_16286,N_17992);
and U21107 (N_21107,N_17939,N_16131);
xor U21108 (N_21108,N_18094,N_17590);
xnor U21109 (N_21109,N_17432,N_18567);
and U21110 (N_21110,N_16770,N_17064);
nand U21111 (N_21111,N_18104,N_16120);
and U21112 (N_21112,N_18461,N_16269);
xnor U21113 (N_21113,N_16671,N_17438);
nand U21114 (N_21114,N_15864,N_16634);
nor U21115 (N_21115,N_17362,N_16119);
and U21116 (N_21116,N_17470,N_18115);
nand U21117 (N_21117,N_18648,N_18206);
nand U21118 (N_21118,N_15813,N_18337);
xor U21119 (N_21119,N_16704,N_16945);
and U21120 (N_21120,N_16063,N_17317);
nor U21121 (N_21121,N_18475,N_17929);
nand U21122 (N_21122,N_17376,N_17558);
nor U21123 (N_21123,N_18039,N_17470);
nor U21124 (N_21124,N_17726,N_17905);
and U21125 (N_21125,N_18745,N_16991);
and U21126 (N_21126,N_17656,N_16723);
nand U21127 (N_21127,N_17290,N_15906);
and U21128 (N_21128,N_18480,N_17154);
and U21129 (N_21129,N_17007,N_17987);
nand U21130 (N_21130,N_17806,N_16386);
or U21131 (N_21131,N_16014,N_16820);
and U21132 (N_21132,N_16863,N_17163);
and U21133 (N_21133,N_16276,N_16683);
and U21134 (N_21134,N_17630,N_17528);
nor U21135 (N_21135,N_17347,N_16834);
xnor U21136 (N_21136,N_17965,N_18458);
xor U21137 (N_21137,N_16486,N_17183);
and U21138 (N_21138,N_15685,N_15828);
or U21139 (N_21139,N_17775,N_17884);
nand U21140 (N_21140,N_16775,N_18469);
nand U21141 (N_21141,N_15885,N_17202);
or U21142 (N_21142,N_16383,N_16792);
and U21143 (N_21143,N_16541,N_16995);
nand U21144 (N_21144,N_17604,N_15743);
and U21145 (N_21145,N_18210,N_18311);
nand U21146 (N_21146,N_15785,N_16448);
and U21147 (N_21147,N_17014,N_16766);
or U21148 (N_21148,N_17213,N_15706);
xnor U21149 (N_21149,N_16529,N_17456);
or U21150 (N_21150,N_17550,N_18405);
or U21151 (N_21151,N_16967,N_18256);
or U21152 (N_21152,N_17746,N_18531);
nor U21153 (N_21153,N_16869,N_16645);
and U21154 (N_21154,N_16951,N_17373);
xnor U21155 (N_21155,N_17520,N_16924);
nand U21156 (N_21156,N_15761,N_18212);
and U21157 (N_21157,N_17885,N_17555);
nor U21158 (N_21158,N_16224,N_16945);
nand U21159 (N_21159,N_18574,N_16298);
or U21160 (N_21160,N_15955,N_16911);
nand U21161 (N_21161,N_17042,N_17603);
and U21162 (N_21162,N_16205,N_17439);
nand U21163 (N_21163,N_18278,N_16291);
and U21164 (N_21164,N_16165,N_16774);
and U21165 (N_21165,N_17214,N_18550);
nor U21166 (N_21166,N_16574,N_16804);
and U21167 (N_21167,N_18701,N_18524);
nor U21168 (N_21168,N_17229,N_18705);
nand U21169 (N_21169,N_17009,N_17540);
and U21170 (N_21170,N_15995,N_18452);
xnor U21171 (N_21171,N_17089,N_17620);
nor U21172 (N_21172,N_16262,N_16001);
or U21173 (N_21173,N_16470,N_17548);
nand U21174 (N_21174,N_16419,N_17865);
or U21175 (N_21175,N_15668,N_17548);
nand U21176 (N_21176,N_17531,N_17104);
nand U21177 (N_21177,N_15786,N_17305);
or U21178 (N_21178,N_17028,N_15915);
or U21179 (N_21179,N_16776,N_18563);
nor U21180 (N_21180,N_17129,N_16862);
and U21181 (N_21181,N_17248,N_15938);
and U21182 (N_21182,N_16873,N_17270);
nor U21183 (N_21183,N_17408,N_18319);
and U21184 (N_21184,N_17391,N_18258);
xnor U21185 (N_21185,N_17423,N_16247);
nor U21186 (N_21186,N_18628,N_16798);
nand U21187 (N_21187,N_17530,N_17387);
xor U21188 (N_21188,N_17343,N_16407);
nor U21189 (N_21189,N_18187,N_18052);
or U21190 (N_21190,N_16694,N_17047);
xor U21191 (N_21191,N_18421,N_16901);
or U21192 (N_21192,N_18065,N_17277);
xor U21193 (N_21193,N_17194,N_17660);
and U21194 (N_21194,N_15939,N_18608);
xnor U21195 (N_21195,N_15741,N_15768);
nor U21196 (N_21196,N_17134,N_17098);
or U21197 (N_21197,N_18432,N_18659);
xor U21198 (N_21198,N_15895,N_16640);
and U21199 (N_21199,N_17134,N_17303);
and U21200 (N_21200,N_17631,N_17615);
and U21201 (N_21201,N_18729,N_16823);
and U21202 (N_21202,N_17978,N_16375);
nor U21203 (N_21203,N_15662,N_18433);
nor U21204 (N_21204,N_17700,N_16322);
xor U21205 (N_21205,N_16312,N_16496);
or U21206 (N_21206,N_16353,N_16216);
nand U21207 (N_21207,N_16345,N_15826);
nand U21208 (N_21208,N_17022,N_16752);
xor U21209 (N_21209,N_18443,N_17804);
and U21210 (N_21210,N_17800,N_16103);
or U21211 (N_21211,N_17325,N_17988);
or U21212 (N_21212,N_16125,N_18152);
and U21213 (N_21213,N_18705,N_18386);
xor U21214 (N_21214,N_18117,N_17995);
xnor U21215 (N_21215,N_17487,N_17659);
nor U21216 (N_21216,N_15877,N_17009);
nor U21217 (N_21217,N_16014,N_16811);
xor U21218 (N_21218,N_15854,N_17133);
nor U21219 (N_21219,N_16088,N_18517);
nor U21220 (N_21220,N_17370,N_17610);
nor U21221 (N_21221,N_17571,N_16625);
or U21222 (N_21222,N_18632,N_18474);
nor U21223 (N_21223,N_18667,N_18106);
or U21224 (N_21224,N_16174,N_16353);
and U21225 (N_21225,N_15642,N_17488);
or U21226 (N_21226,N_16837,N_17605);
xnor U21227 (N_21227,N_15928,N_16766);
and U21228 (N_21228,N_16927,N_16479);
xor U21229 (N_21229,N_16973,N_17535);
nor U21230 (N_21230,N_18630,N_17591);
nor U21231 (N_21231,N_17971,N_16529);
nor U21232 (N_21232,N_16993,N_17392);
nand U21233 (N_21233,N_18492,N_16775);
or U21234 (N_21234,N_17258,N_16233);
or U21235 (N_21235,N_18052,N_17052);
nor U21236 (N_21236,N_18136,N_18054);
nand U21237 (N_21237,N_18024,N_17229);
nor U21238 (N_21238,N_16553,N_17672);
nand U21239 (N_21239,N_16910,N_17122);
and U21240 (N_21240,N_17317,N_16525);
or U21241 (N_21241,N_17847,N_16146);
nand U21242 (N_21242,N_17572,N_18102);
nor U21243 (N_21243,N_18081,N_16913);
xnor U21244 (N_21244,N_16264,N_18216);
xnor U21245 (N_21245,N_15648,N_18240);
nor U21246 (N_21246,N_17200,N_16430);
nor U21247 (N_21247,N_18443,N_17622);
or U21248 (N_21248,N_16438,N_15629);
nand U21249 (N_21249,N_18517,N_16677);
xor U21250 (N_21250,N_18613,N_15646);
nand U21251 (N_21251,N_18232,N_18387);
nor U21252 (N_21252,N_15877,N_17090);
xnor U21253 (N_21253,N_18715,N_18603);
or U21254 (N_21254,N_15777,N_16542);
or U21255 (N_21255,N_16273,N_16125);
or U21256 (N_21256,N_17808,N_17616);
nand U21257 (N_21257,N_16474,N_17429);
nor U21258 (N_21258,N_15741,N_15855);
nand U21259 (N_21259,N_17596,N_17315);
nand U21260 (N_21260,N_18389,N_18154);
nand U21261 (N_21261,N_17550,N_16229);
nand U21262 (N_21262,N_16863,N_18189);
nor U21263 (N_21263,N_18632,N_18487);
nand U21264 (N_21264,N_17912,N_17918);
xor U21265 (N_21265,N_15957,N_18502);
nor U21266 (N_21266,N_17618,N_17820);
nor U21267 (N_21267,N_18521,N_16897);
xnor U21268 (N_21268,N_17360,N_18351);
or U21269 (N_21269,N_17078,N_15813);
xor U21270 (N_21270,N_16985,N_15699);
or U21271 (N_21271,N_17355,N_17023);
nor U21272 (N_21272,N_15662,N_16967);
nor U21273 (N_21273,N_16921,N_16764);
xnor U21274 (N_21274,N_17674,N_18023);
nor U21275 (N_21275,N_18423,N_16903);
nand U21276 (N_21276,N_17641,N_16752);
and U21277 (N_21277,N_15844,N_18671);
xnor U21278 (N_21278,N_18021,N_15782);
nor U21279 (N_21279,N_18028,N_16956);
nor U21280 (N_21280,N_18054,N_18185);
and U21281 (N_21281,N_16963,N_16986);
and U21282 (N_21282,N_18294,N_15703);
nand U21283 (N_21283,N_17288,N_16413);
nand U21284 (N_21284,N_18257,N_15872);
or U21285 (N_21285,N_17654,N_18277);
or U21286 (N_21286,N_18582,N_15674);
nand U21287 (N_21287,N_18746,N_16487);
and U21288 (N_21288,N_18370,N_16825);
and U21289 (N_21289,N_17399,N_17044);
nor U21290 (N_21290,N_17154,N_16122);
xnor U21291 (N_21291,N_18282,N_17322);
and U21292 (N_21292,N_15952,N_16236);
and U21293 (N_21293,N_16055,N_16734);
nand U21294 (N_21294,N_17135,N_18686);
xor U21295 (N_21295,N_18345,N_16372);
or U21296 (N_21296,N_17282,N_15927);
xnor U21297 (N_21297,N_16110,N_17397);
xor U21298 (N_21298,N_16415,N_16293);
xor U21299 (N_21299,N_15853,N_18164);
nor U21300 (N_21300,N_18397,N_16150);
nor U21301 (N_21301,N_16638,N_18033);
nand U21302 (N_21302,N_16535,N_17088);
nor U21303 (N_21303,N_17824,N_18000);
or U21304 (N_21304,N_17377,N_18602);
nor U21305 (N_21305,N_16854,N_17568);
or U21306 (N_21306,N_17954,N_16861);
or U21307 (N_21307,N_16987,N_15999);
or U21308 (N_21308,N_17808,N_16824);
and U21309 (N_21309,N_16332,N_15971);
nor U21310 (N_21310,N_18162,N_16024);
xor U21311 (N_21311,N_15712,N_16402);
nand U21312 (N_21312,N_15716,N_15672);
nor U21313 (N_21313,N_17494,N_18388);
nand U21314 (N_21314,N_17043,N_17058);
xor U21315 (N_21315,N_18408,N_17809);
nand U21316 (N_21316,N_15706,N_17225);
and U21317 (N_21317,N_15686,N_17092);
and U21318 (N_21318,N_17327,N_18606);
xor U21319 (N_21319,N_17031,N_16196);
xnor U21320 (N_21320,N_18188,N_15971);
and U21321 (N_21321,N_17705,N_16457);
nor U21322 (N_21322,N_16344,N_17842);
or U21323 (N_21323,N_17971,N_17227);
nand U21324 (N_21324,N_17130,N_16054);
and U21325 (N_21325,N_16473,N_16697);
xor U21326 (N_21326,N_18711,N_15660);
xor U21327 (N_21327,N_16702,N_17292);
xor U21328 (N_21328,N_17709,N_17063);
and U21329 (N_21329,N_16646,N_17585);
or U21330 (N_21330,N_15924,N_16401);
or U21331 (N_21331,N_16411,N_18540);
nor U21332 (N_21332,N_18486,N_16301);
nor U21333 (N_21333,N_17906,N_16529);
or U21334 (N_21334,N_16380,N_17937);
nand U21335 (N_21335,N_16424,N_18187);
nand U21336 (N_21336,N_17793,N_17846);
or U21337 (N_21337,N_17243,N_18489);
nand U21338 (N_21338,N_17143,N_16988);
or U21339 (N_21339,N_16980,N_18015);
xor U21340 (N_21340,N_15840,N_18011);
or U21341 (N_21341,N_18731,N_17413);
nand U21342 (N_21342,N_18256,N_16676);
nor U21343 (N_21343,N_16869,N_18380);
and U21344 (N_21344,N_18393,N_16426);
or U21345 (N_21345,N_18063,N_17104);
or U21346 (N_21346,N_17050,N_18512);
and U21347 (N_21347,N_17955,N_17138);
or U21348 (N_21348,N_17231,N_16793);
nor U21349 (N_21349,N_17159,N_18261);
nor U21350 (N_21350,N_16966,N_18069);
xnor U21351 (N_21351,N_16715,N_18356);
or U21352 (N_21352,N_16127,N_18455);
xnor U21353 (N_21353,N_16577,N_18650);
xor U21354 (N_21354,N_16952,N_16526);
xnor U21355 (N_21355,N_16927,N_16654);
xor U21356 (N_21356,N_18454,N_16741);
nand U21357 (N_21357,N_18723,N_18395);
nand U21358 (N_21358,N_18428,N_18127);
and U21359 (N_21359,N_16280,N_17237);
xor U21360 (N_21360,N_18296,N_16409);
nor U21361 (N_21361,N_17139,N_17708);
xnor U21362 (N_21362,N_16239,N_17384);
nor U21363 (N_21363,N_16826,N_18489);
nand U21364 (N_21364,N_15917,N_18029);
or U21365 (N_21365,N_16165,N_16504);
nand U21366 (N_21366,N_15894,N_16614);
nand U21367 (N_21367,N_17821,N_17036);
nand U21368 (N_21368,N_16283,N_17441);
or U21369 (N_21369,N_16442,N_15672);
nand U21370 (N_21370,N_18156,N_16758);
and U21371 (N_21371,N_18208,N_15713);
xnor U21372 (N_21372,N_17406,N_15652);
or U21373 (N_21373,N_18161,N_15640);
nand U21374 (N_21374,N_18149,N_18172);
nand U21375 (N_21375,N_17457,N_17748);
nor U21376 (N_21376,N_18486,N_16765);
and U21377 (N_21377,N_18732,N_18501);
nor U21378 (N_21378,N_18440,N_16000);
xnor U21379 (N_21379,N_16358,N_16205);
and U21380 (N_21380,N_16364,N_18010);
xnor U21381 (N_21381,N_16170,N_16751);
xor U21382 (N_21382,N_16006,N_18711);
or U21383 (N_21383,N_18445,N_18068);
nor U21384 (N_21384,N_17064,N_15905);
nand U21385 (N_21385,N_15709,N_15984);
nand U21386 (N_21386,N_17166,N_16637);
nor U21387 (N_21387,N_16985,N_16733);
or U21388 (N_21388,N_18595,N_18100);
and U21389 (N_21389,N_16504,N_17603);
xnor U21390 (N_21390,N_18644,N_16265);
or U21391 (N_21391,N_15661,N_17447);
nand U21392 (N_21392,N_17345,N_17524);
or U21393 (N_21393,N_18143,N_16147);
xnor U21394 (N_21394,N_18318,N_16919);
nor U21395 (N_21395,N_17391,N_16727);
and U21396 (N_21396,N_16648,N_18522);
nor U21397 (N_21397,N_17598,N_17989);
nor U21398 (N_21398,N_17347,N_17417);
xor U21399 (N_21399,N_18393,N_18096);
nor U21400 (N_21400,N_16606,N_15781);
xnor U21401 (N_21401,N_18353,N_16692);
nand U21402 (N_21402,N_16723,N_16783);
xnor U21403 (N_21403,N_17723,N_18591);
and U21404 (N_21404,N_15889,N_18454);
nand U21405 (N_21405,N_17758,N_15871);
nand U21406 (N_21406,N_16003,N_17521);
xor U21407 (N_21407,N_16354,N_17266);
and U21408 (N_21408,N_17557,N_16514);
or U21409 (N_21409,N_17114,N_18009);
or U21410 (N_21410,N_16823,N_18036);
nor U21411 (N_21411,N_17174,N_17170);
and U21412 (N_21412,N_17342,N_17483);
and U21413 (N_21413,N_17266,N_16489);
xor U21414 (N_21414,N_16131,N_18391);
xor U21415 (N_21415,N_18095,N_16632);
xnor U21416 (N_21416,N_18738,N_18193);
or U21417 (N_21417,N_16474,N_16053);
xor U21418 (N_21418,N_17353,N_16822);
nand U21419 (N_21419,N_17223,N_17078);
xnor U21420 (N_21420,N_15634,N_17832);
or U21421 (N_21421,N_17159,N_18486);
and U21422 (N_21422,N_16160,N_18617);
or U21423 (N_21423,N_16069,N_16808);
and U21424 (N_21424,N_16663,N_18290);
xor U21425 (N_21425,N_16376,N_17959);
nand U21426 (N_21426,N_18151,N_17597);
and U21427 (N_21427,N_15999,N_16846);
or U21428 (N_21428,N_16478,N_17850);
nand U21429 (N_21429,N_18595,N_15932);
nand U21430 (N_21430,N_18343,N_18366);
or U21431 (N_21431,N_16337,N_16910);
and U21432 (N_21432,N_18026,N_15937);
and U21433 (N_21433,N_17658,N_17146);
nand U21434 (N_21434,N_16502,N_17275);
and U21435 (N_21435,N_16343,N_18268);
nand U21436 (N_21436,N_17363,N_15945);
nand U21437 (N_21437,N_16810,N_16117);
and U21438 (N_21438,N_16320,N_16428);
xor U21439 (N_21439,N_18526,N_16930);
and U21440 (N_21440,N_17003,N_16608);
nor U21441 (N_21441,N_17849,N_18437);
xnor U21442 (N_21442,N_16368,N_17239);
and U21443 (N_21443,N_18345,N_18141);
and U21444 (N_21444,N_15827,N_17571);
xnor U21445 (N_21445,N_16391,N_18176);
and U21446 (N_21446,N_18204,N_17342);
and U21447 (N_21447,N_16813,N_17889);
nand U21448 (N_21448,N_16205,N_16673);
and U21449 (N_21449,N_18684,N_16535);
xnor U21450 (N_21450,N_18184,N_17923);
nor U21451 (N_21451,N_17627,N_16161);
xor U21452 (N_21452,N_16598,N_18637);
and U21453 (N_21453,N_16061,N_16271);
nand U21454 (N_21454,N_16393,N_16505);
nand U21455 (N_21455,N_17996,N_15757);
nor U21456 (N_21456,N_17237,N_18139);
or U21457 (N_21457,N_16202,N_16381);
nand U21458 (N_21458,N_16613,N_16342);
and U21459 (N_21459,N_18672,N_17630);
nand U21460 (N_21460,N_18620,N_17587);
and U21461 (N_21461,N_17046,N_15723);
and U21462 (N_21462,N_18562,N_17817);
nor U21463 (N_21463,N_18324,N_17938);
nand U21464 (N_21464,N_17781,N_18401);
or U21465 (N_21465,N_18050,N_17283);
nand U21466 (N_21466,N_18578,N_17181);
xnor U21467 (N_21467,N_15880,N_15776);
and U21468 (N_21468,N_18375,N_18562);
or U21469 (N_21469,N_18615,N_16941);
xor U21470 (N_21470,N_17972,N_16109);
nand U21471 (N_21471,N_16186,N_18288);
nand U21472 (N_21472,N_17427,N_17570);
and U21473 (N_21473,N_17381,N_16400);
nor U21474 (N_21474,N_17069,N_18260);
xnor U21475 (N_21475,N_16203,N_16610);
nand U21476 (N_21476,N_16986,N_18480);
nor U21477 (N_21477,N_17399,N_16935);
and U21478 (N_21478,N_16350,N_17225);
xnor U21479 (N_21479,N_16598,N_18132);
nand U21480 (N_21480,N_18087,N_17754);
nor U21481 (N_21481,N_18435,N_16903);
nand U21482 (N_21482,N_18658,N_17648);
and U21483 (N_21483,N_18441,N_17056);
and U21484 (N_21484,N_16070,N_18054);
nor U21485 (N_21485,N_16913,N_16279);
or U21486 (N_21486,N_15808,N_18740);
or U21487 (N_21487,N_17600,N_15848);
and U21488 (N_21488,N_17868,N_18315);
xnor U21489 (N_21489,N_16149,N_15901);
nor U21490 (N_21490,N_18357,N_18653);
nand U21491 (N_21491,N_16724,N_17953);
xnor U21492 (N_21492,N_16889,N_18452);
nand U21493 (N_21493,N_17387,N_18169);
nand U21494 (N_21494,N_16100,N_17880);
or U21495 (N_21495,N_18413,N_15887);
and U21496 (N_21496,N_16957,N_17503);
nand U21497 (N_21497,N_16066,N_16320);
and U21498 (N_21498,N_16863,N_18388);
and U21499 (N_21499,N_18233,N_18198);
nand U21500 (N_21500,N_18501,N_17256);
or U21501 (N_21501,N_17203,N_15806);
nor U21502 (N_21502,N_17902,N_17336);
or U21503 (N_21503,N_16800,N_16374);
nor U21504 (N_21504,N_18067,N_17759);
and U21505 (N_21505,N_18022,N_18696);
nor U21506 (N_21506,N_18127,N_15676);
xnor U21507 (N_21507,N_16697,N_18342);
nor U21508 (N_21508,N_18243,N_16682);
and U21509 (N_21509,N_15945,N_16996);
nor U21510 (N_21510,N_17770,N_17506);
nand U21511 (N_21511,N_18477,N_16335);
nand U21512 (N_21512,N_15786,N_18353);
and U21513 (N_21513,N_18519,N_18462);
xnor U21514 (N_21514,N_16706,N_17015);
and U21515 (N_21515,N_17920,N_16292);
xor U21516 (N_21516,N_17344,N_17924);
nor U21517 (N_21517,N_17588,N_15825);
nand U21518 (N_21518,N_17201,N_16918);
nor U21519 (N_21519,N_17927,N_18453);
or U21520 (N_21520,N_17693,N_15786);
or U21521 (N_21521,N_17600,N_17412);
and U21522 (N_21522,N_17026,N_18369);
nor U21523 (N_21523,N_17217,N_18168);
nor U21524 (N_21524,N_15873,N_18271);
and U21525 (N_21525,N_16130,N_16017);
and U21526 (N_21526,N_16079,N_16488);
or U21527 (N_21527,N_18619,N_16692);
nor U21528 (N_21528,N_18560,N_18047);
or U21529 (N_21529,N_17971,N_17017);
and U21530 (N_21530,N_16991,N_17015);
nand U21531 (N_21531,N_17929,N_15699);
nor U21532 (N_21532,N_16135,N_17060);
and U21533 (N_21533,N_16711,N_17597);
or U21534 (N_21534,N_16208,N_16049);
or U21535 (N_21535,N_15773,N_16740);
and U21536 (N_21536,N_18745,N_18552);
nand U21537 (N_21537,N_18527,N_17667);
and U21538 (N_21538,N_17506,N_18320);
nand U21539 (N_21539,N_16936,N_16662);
and U21540 (N_21540,N_16592,N_16490);
nand U21541 (N_21541,N_16522,N_15900);
and U21542 (N_21542,N_18525,N_17275);
nand U21543 (N_21543,N_18378,N_16708);
nor U21544 (N_21544,N_18744,N_17274);
xor U21545 (N_21545,N_15985,N_16730);
nand U21546 (N_21546,N_16751,N_17306);
nor U21547 (N_21547,N_18503,N_16609);
nor U21548 (N_21548,N_17456,N_16573);
nor U21549 (N_21549,N_17751,N_16577);
xor U21550 (N_21550,N_16107,N_17804);
nor U21551 (N_21551,N_16446,N_15812);
or U21552 (N_21552,N_17399,N_17714);
or U21553 (N_21553,N_15698,N_18559);
and U21554 (N_21554,N_17033,N_17516);
or U21555 (N_21555,N_16671,N_16836);
or U21556 (N_21556,N_18431,N_17960);
and U21557 (N_21557,N_17553,N_16907);
nor U21558 (N_21558,N_16879,N_18133);
nor U21559 (N_21559,N_16994,N_16526);
nand U21560 (N_21560,N_16391,N_17698);
nor U21561 (N_21561,N_16031,N_17983);
nand U21562 (N_21562,N_15837,N_18534);
nor U21563 (N_21563,N_18071,N_16326);
xnor U21564 (N_21564,N_17752,N_17237);
nand U21565 (N_21565,N_15670,N_18384);
and U21566 (N_21566,N_18651,N_18348);
nand U21567 (N_21567,N_16417,N_18407);
nor U21568 (N_21568,N_17135,N_17382);
xor U21569 (N_21569,N_16682,N_17505);
nand U21570 (N_21570,N_18282,N_18513);
nor U21571 (N_21571,N_18485,N_18133);
nand U21572 (N_21572,N_17910,N_18162);
or U21573 (N_21573,N_18049,N_16974);
nand U21574 (N_21574,N_18596,N_15684);
or U21575 (N_21575,N_18460,N_17837);
and U21576 (N_21576,N_16737,N_16313);
nor U21577 (N_21577,N_16073,N_17886);
nand U21578 (N_21578,N_18418,N_17707);
or U21579 (N_21579,N_17736,N_18427);
or U21580 (N_21580,N_16727,N_15919);
nand U21581 (N_21581,N_18017,N_16050);
nor U21582 (N_21582,N_18361,N_16905);
or U21583 (N_21583,N_16676,N_15629);
nor U21584 (N_21584,N_15630,N_17243);
nand U21585 (N_21585,N_18452,N_16118);
and U21586 (N_21586,N_16971,N_18174);
nand U21587 (N_21587,N_18129,N_18070);
xor U21588 (N_21588,N_17587,N_16570);
nor U21589 (N_21589,N_16660,N_15882);
nand U21590 (N_21590,N_18479,N_16088);
nor U21591 (N_21591,N_17587,N_17437);
xnor U21592 (N_21592,N_18020,N_18558);
nand U21593 (N_21593,N_17799,N_16395);
xnor U21594 (N_21594,N_18440,N_18000);
or U21595 (N_21595,N_16007,N_15715);
nor U21596 (N_21596,N_17619,N_18042);
or U21597 (N_21597,N_17468,N_18065);
or U21598 (N_21598,N_18294,N_16263);
and U21599 (N_21599,N_16528,N_16320);
nand U21600 (N_21600,N_16137,N_17614);
nand U21601 (N_21601,N_16501,N_17221);
nor U21602 (N_21602,N_16852,N_17894);
and U21603 (N_21603,N_17665,N_16444);
nor U21604 (N_21604,N_18010,N_16031);
xnor U21605 (N_21605,N_15725,N_16568);
nand U21606 (N_21606,N_17692,N_16057);
nand U21607 (N_21607,N_17782,N_18472);
or U21608 (N_21608,N_16707,N_16486);
or U21609 (N_21609,N_17166,N_18004);
nor U21610 (N_21610,N_16866,N_18725);
or U21611 (N_21611,N_18055,N_17281);
nand U21612 (N_21612,N_17284,N_16666);
xor U21613 (N_21613,N_18050,N_18157);
nand U21614 (N_21614,N_16365,N_16490);
nand U21615 (N_21615,N_17127,N_17216);
xor U21616 (N_21616,N_16142,N_15778);
nand U21617 (N_21617,N_16142,N_18473);
xnor U21618 (N_21618,N_17998,N_16151);
xor U21619 (N_21619,N_16916,N_17152);
nand U21620 (N_21620,N_16509,N_17996);
nand U21621 (N_21621,N_15851,N_16846);
and U21622 (N_21622,N_16921,N_18467);
or U21623 (N_21623,N_17342,N_17878);
nand U21624 (N_21624,N_17167,N_16625);
or U21625 (N_21625,N_17484,N_16208);
or U21626 (N_21626,N_18413,N_16496);
and U21627 (N_21627,N_18394,N_16492);
nand U21628 (N_21628,N_16747,N_18177);
nor U21629 (N_21629,N_17455,N_16961);
nor U21630 (N_21630,N_16745,N_17521);
nand U21631 (N_21631,N_15883,N_17103);
nand U21632 (N_21632,N_16586,N_18496);
and U21633 (N_21633,N_17501,N_17234);
or U21634 (N_21634,N_16322,N_16641);
and U21635 (N_21635,N_17082,N_16616);
nor U21636 (N_21636,N_18112,N_17821);
or U21637 (N_21637,N_15917,N_17359);
nor U21638 (N_21638,N_17151,N_16925);
nor U21639 (N_21639,N_17999,N_17480);
or U21640 (N_21640,N_17671,N_16453);
nand U21641 (N_21641,N_18171,N_16089);
or U21642 (N_21642,N_17241,N_17785);
nand U21643 (N_21643,N_16087,N_18162);
xnor U21644 (N_21644,N_18580,N_15673);
xnor U21645 (N_21645,N_16813,N_17330);
and U21646 (N_21646,N_18676,N_18074);
xnor U21647 (N_21647,N_17202,N_18544);
or U21648 (N_21648,N_17879,N_15894);
and U21649 (N_21649,N_15725,N_17780);
nor U21650 (N_21650,N_17381,N_18591);
nor U21651 (N_21651,N_16925,N_16958);
xnor U21652 (N_21652,N_15869,N_17581);
xnor U21653 (N_21653,N_16595,N_16422);
nor U21654 (N_21654,N_16676,N_16284);
and U21655 (N_21655,N_18504,N_16230);
and U21656 (N_21656,N_16792,N_18334);
xnor U21657 (N_21657,N_18493,N_16705);
nand U21658 (N_21658,N_18557,N_16504);
or U21659 (N_21659,N_16654,N_18670);
or U21660 (N_21660,N_18264,N_18020);
xnor U21661 (N_21661,N_16045,N_16308);
and U21662 (N_21662,N_18165,N_17996);
and U21663 (N_21663,N_17710,N_17528);
nand U21664 (N_21664,N_16966,N_18347);
nand U21665 (N_21665,N_16095,N_18674);
nor U21666 (N_21666,N_15845,N_17893);
and U21667 (N_21667,N_16926,N_15780);
xnor U21668 (N_21668,N_17092,N_15964);
or U21669 (N_21669,N_18714,N_16451);
and U21670 (N_21670,N_17584,N_17585);
nor U21671 (N_21671,N_17142,N_16206);
nor U21672 (N_21672,N_18698,N_18319);
nand U21673 (N_21673,N_17311,N_18722);
and U21674 (N_21674,N_17635,N_17233);
and U21675 (N_21675,N_16135,N_17446);
xnor U21676 (N_21676,N_16185,N_15827);
nand U21677 (N_21677,N_18070,N_18133);
nand U21678 (N_21678,N_18415,N_17443);
nand U21679 (N_21679,N_16909,N_18209);
or U21680 (N_21680,N_16978,N_18295);
nand U21681 (N_21681,N_17243,N_17528);
nand U21682 (N_21682,N_17248,N_16454);
nand U21683 (N_21683,N_15995,N_15848);
or U21684 (N_21684,N_16885,N_16908);
nand U21685 (N_21685,N_17426,N_18215);
or U21686 (N_21686,N_15859,N_17716);
xor U21687 (N_21687,N_18197,N_15666);
nor U21688 (N_21688,N_17944,N_18208);
nand U21689 (N_21689,N_17290,N_18187);
or U21690 (N_21690,N_17700,N_18403);
and U21691 (N_21691,N_17353,N_17300);
or U21692 (N_21692,N_18616,N_15929);
and U21693 (N_21693,N_16482,N_18381);
nor U21694 (N_21694,N_17121,N_16660);
nand U21695 (N_21695,N_16510,N_16304);
nand U21696 (N_21696,N_17612,N_15647);
nand U21697 (N_21697,N_17743,N_16581);
xor U21698 (N_21698,N_16197,N_16747);
and U21699 (N_21699,N_16255,N_16655);
nand U21700 (N_21700,N_18004,N_15931);
nor U21701 (N_21701,N_17789,N_17393);
xnor U21702 (N_21702,N_17911,N_16792);
and U21703 (N_21703,N_17346,N_16644);
nand U21704 (N_21704,N_17272,N_18090);
xnor U21705 (N_21705,N_17156,N_18272);
nand U21706 (N_21706,N_17615,N_16118);
or U21707 (N_21707,N_15837,N_17396);
xnor U21708 (N_21708,N_17623,N_18747);
nand U21709 (N_21709,N_18613,N_15757);
nor U21710 (N_21710,N_16946,N_16525);
nor U21711 (N_21711,N_16609,N_18069);
nor U21712 (N_21712,N_16512,N_16705);
and U21713 (N_21713,N_16552,N_17946);
nand U21714 (N_21714,N_16507,N_15906);
nor U21715 (N_21715,N_17852,N_16358);
nor U21716 (N_21716,N_15716,N_18111);
and U21717 (N_21717,N_17298,N_18690);
and U21718 (N_21718,N_17254,N_16555);
and U21719 (N_21719,N_18125,N_18555);
nor U21720 (N_21720,N_18095,N_17517);
nand U21721 (N_21721,N_18151,N_16467);
nor U21722 (N_21722,N_16491,N_15974);
nor U21723 (N_21723,N_18591,N_17813);
xor U21724 (N_21724,N_16857,N_18487);
xnor U21725 (N_21725,N_17221,N_15835);
or U21726 (N_21726,N_18027,N_17341);
or U21727 (N_21727,N_17339,N_17374);
nand U21728 (N_21728,N_17128,N_18202);
nor U21729 (N_21729,N_18212,N_18554);
xnor U21730 (N_21730,N_16903,N_16969);
xor U21731 (N_21731,N_18571,N_17710);
or U21732 (N_21732,N_18124,N_16782);
nand U21733 (N_21733,N_18139,N_16624);
nand U21734 (N_21734,N_17425,N_17205);
or U21735 (N_21735,N_18209,N_18655);
nand U21736 (N_21736,N_18364,N_16519);
or U21737 (N_21737,N_15962,N_16697);
nand U21738 (N_21738,N_16444,N_16625);
or U21739 (N_21739,N_16755,N_15654);
and U21740 (N_21740,N_16933,N_16641);
or U21741 (N_21741,N_15660,N_16623);
xor U21742 (N_21742,N_17498,N_17349);
or U21743 (N_21743,N_16002,N_15908);
xor U21744 (N_21744,N_16602,N_17779);
or U21745 (N_21745,N_17824,N_17519);
and U21746 (N_21746,N_15786,N_18703);
and U21747 (N_21747,N_16602,N_16896);
xor U21748 (N_21748,N_17553,N_17405);
or U21749 (N_21749,N_18077,N_17445);
nor U21750 (N_21750,N_18737,N_17196);
and U21751 (N_21751,N_15768,N_17822);
nor U21752 (N_21752,N_15913,N_16405);
nand U21753 (N_21753,N_17899,N_18608);
and U21754 (N_21754,N_16494,N_18203);
xnor U21755 (N_21755,N_16234,N_16331);
and U21756 (N_21756,N_16592,N_17639);
and U21757 (N_21757,N_15998,N_18049);
or U21758 (N_21758,N_17087,N_18457);
nor U21759 (N_21759,N_16612,N_17347);
and U21760 (N_21760,N_16938,N_18316);
and U21761 (N_21761,N_16459,N_17756);
xor U21762 (N_21762,N_15897,N_18262);
xor U21763 (N_21763,N_17103,N_17479);
or U21764 (N_21764,N_18280,N_16711);
nand U21765 (N_21765,N_17627,N_16703);
nor U21766 (N_21766,N_17899,N_18498);
xnor U21767 (N_21767,N_18296,N_16688);
or U21768 (N_21768,N_17409,N_17261);
nor U21769 (N_21769,N_18061,N_18495);
xnor U21770 (N_21770,N_18223,N_16360);
nor U21771 (N_21771,N_18606,N_16145);
nand U21772 (N_21772,N_18601,N_15782);
or U21773 (N_21773,N_18271,N_17920);
nor U21774 (N_21774,N_16332,N_15953);
nor U21775 (N_21775,N_17118,N_15936);
or U21776 (N_21776,N_17168,N_17040);
nor U21777 (N_21777,N_15833,N_15853);
and U21778 (N_21778,N_18259,N_17821);
xnor U21779 (N_21779,N_17191,N_18586);
and U21780 (N_21780,N_18485,N_16024);
xor U21781 (N_21781,N_16834,N_17270);
xor U21782 (N_21782,N_18548,N_15813);
and U21783 (N_21783,N_16831,N_16785);
xnor U21784 (N_21784,N_17105,N_17351);
nand U21785 (N_21785,N_16864,N_16723);
and U21786 (N_21786,N_15822,N_17003);
xor U21787 (N_21787,N_17749,N_16067);
and U21788 (N_21788,N_18684,N_18134);
nor U21789 (N_21789,N_17981,N_16686);
or U21790 (N_21790,N_16411,N_16733);
nand U21791 (N_21791,N_17040,N_15900);
nor U21792 (N_21792,N_16319,N_18171);
nor U21793 (N_21793,N_16670,N_18748);
nor U21794 (N_21794,N_17755,N_15927);
xor U21795 (N_21795,N_18111,N_16740);
nor U21796 (N_21796,N_17143,N_16578);
xnor U21797 (N_21797,N_17908,N_18678);
and U21798 (N_21798,N_16194,N_16067);
nor U21799 (N_21799,N_17443,N_18127);
nand U21800 (N_21800,N_17950,N_16913);
xnor U21801 (N_21801,N_17384,N_17480);
or U21802 (N_21802,N_18155,N_17733);
xnor U21803 (N_21803,N_17702,N_17092);
and U21804 (N_21804,N_15681,N_18137);
or U21805 (N_21805,N_17096,N_18158);
nor U21806 (N_21806,N_18365,N_16050);
nor U21807 (N_21807,N_15922,N_17416);
and U21808 (N_21808,N_15862,N_15763);
and U21809 (N_21809,N_18215,N_17485);
xor U21810 (N_21810,N_15944,N_17255);
xnor U21811 (N_21811,N_15980,N_18429);
nor U21812 (N_21812,N_15668,N_18740);
xnor U21813 (N_21813,N_16049,N_18332);
xnor U21814 (N_21814,N_18205,N_17656);
xnor U21815 (N_21815,N_16279,N_16303);
nor U21816 (N_21816,N_16552,N_17131);
nand U21817 (N_21817,N_18475,N_17157);
or U21818 (N_21818,N_18693,N_18016);
xor U21819 (N_21819,N_18176,N_17107);
and U21820 (N_21820,N_17336,N_17532);
nor U21821 (N_21821,N_15998,N_15957);
xnor U21822 (N_21822,N_16298,N_17212);
and U21823 (N_21823,N_17644,N_17363);
nand U21824 (N_21824,N_17305,N_17858);
nand U21825 (N_21825,N_16520,N_15653);
nand U21826 (N_21826,N_16409,N_16972);
nor U21827 (N_21827,N_17161,N_18562);
and U21828 (N_21828,N_15654,N_18433);
or U21829 (N_21829,N_18257,N_17209);
nand U21830 (N_21830,N_15753,N_16350);
nor U21831 (N_21831,N_18012,N_18566);
nand U21832 (N_21832,N_18040,N_16596);
nor U21833 (N_21833,N_17496,N_17840);
nand U21834 (N_21834,N_16493,N_16076);
and U21835 (N_21835,N_16361,N_17412);
nand U21836 (N_21836,N_17843,N_16180);
or U21837 (N_21837,N_17935,N_18453);
or U21838 (N_21838,N_17110,N_15790);
and U21839 (N_21839,N_17522,N_17479);
and U21840 (N_21840,N_18537,N_16274);
or U21841 (N_21841,N_15993,N_18307);
xnor U21842 (N_21842,N_17018,N_16308);
nand U21843 (N_21843,N_16144,N_15760);
nor U21844 (N_21844,N_18232,N_18467);
and U21845 (N_21845,N_17824,N_17419);
or U21846 (N_21846,N_16174,N_16881);
nor U21847 (N_21847,N_18358,N_18433);
or U21848 (N_21848,N_18296,N_18565);
nand U21849 (N_21849,N_18629,N_15968);
nor U21850 (N_21850,N_17494,N_17649);
xor U21851 (N_21851,N_17646,N_17536);
xor U21852 (N_21852,N_16577,N_16920);
nor U21853 (N_21853,N_18372,N_17922);
nor U21854 (N_21854,N_16273,N_17954);
nand U21855 (N_21855,N_16660,N_16560);
or U21856 (N_21856,N_17997,N_15631);
nor U21857 (N_21857,N_17263,N_17661);
xor U21858 (N_21858,N_16912,N_16356);
or U21859 (N_21859,N_18239,N_17036);
nor U21860 (N_21860,N_16889,N_15994);
or U21861 (N_21861,N_16698,N_17212);
and U21862 (N_21862,N_15941,N_17932);
and U21863 (N_21863,N_18061,N_17896);
or U21864 (N_21864,N_18444,N_18513);
nor U21865 (N_21865,N_15649,N_17324);
xor U21866 (N_21866,N_18040,N_17006);
xor U21867 (N_21867,N_17058,N_17313);
nand U21868 (N_21868,N_17477,N_16301);
and U21869 (N_21869,N_16468,N_17466);
nand U21870 (N_21870,N_16602,N_16983);
nor U21871 (N_21871,N_16995,N_16353);
nor U21872 (N_21872,N_16799,N_18644);
and U21873 (N_21873,N_18283,N_16383);
xnor U21874 (N_21874,N_18725,N_16727);
xnor U21875 (N_21875,N_20334,N_20956);
and U21876 (N_21876,N_21433,N_21463);
nor U21877 (N_21877,N_21153,N_19757);
or U21878 (N_21878,N_19193,N_19957);
and U21879 (N_21879,N_19215,N_21760);
and U21880 (N_21880,N_21233,N_18929);
and U21881 (N_21881,N_21690,N_19488);
and U21882 (N_21882,N_20417,N_18994);
xnor U21883 (N_21883,N_20756,N_19263);
nand U21884 (N_21884,N_21624,N_19666);
and U21885 (N_21885,N_20666,N_20827);
or U21886 (N_21886,N_21071,N_19566);
or U21887 (N_21887,N_20706,N_19416);
and U21888 (N_21888,N_21864,N_20283);
nor U21889 (N_21889,N_21493,N_20718);
or U21890 (N_21890,N_19448,N_19035);
and U21891 (N_21891,N_20160,N_20661);
or U21892 (N_21892,N_21570,N_18989);
xnor U21893 (N_21893,N_20233,N_19521);
and U21894 (N_21894,N_21273,N_18816);
and U21895 (N_21895,N_20646,N_19544);
and U21896 (N_21896,N_20958,N_18909);
nand U21897 (N_21897,N_20917,N_20112);
and U21898 (N_21898,N_21098,N_19996);
or U21899 (N_21899,N_21067,N_18890);
xnor U21900 (N_21900,N_19690,N_21562);
nand U21901 (N_21901,N_21236,N_19886);
or U21902 (N_21902,N_20945,N_19238);
or U21903 (N_21903,N_20571,N_19583);
nand U21904 (N_21904,N_20149,N_20957);
or U21905 (N_21905,N_19721,N_20327);
and U21906 (N_21906,N_21210,N_19111);
nor U21907 (N_21907,N_20590,N_20556);
xor U21908 (N_21908,N_21581,N_18789);
and U21909 (N_21909,N_19955,N_21489);
nand U21910 (N_21910,N_20132,N_19242);
or U21911 (N_21911,N_19565,N_19105);
xnor U21912 (N_21912,N_20163,N_21605);
nand U21913 (N_21913,N_21050,N_19115);
xnor U21914 (N_21914,N_19545,N_21269);
and U21915 (N_21915,N_21467,N_21752);
nor U21916 (N_21916,N_19007,N_20591);
nor U21917 (N_21917,N_21850,N_20131);
xor U21918 (N_21918,N_19301,N_21123);
nor U21919 (N_21919,N_21754,N_19716);
xor U21920 (N_21920,N_20492,N_19181);
or U21921 (N_21921,N_20007,N_20157);
nor U21922 (N_21922,N_19718,N_19205);
nand U21923 (N_21923,N_20057,N_20375);
and U21924 (N_21924,N_21803,N_19761);
or U21925 (N_21925,N_20660,N_19558);
or U21926 (N_21926,N_19348,N_21836);
or U21927 (N_21927,N_18972,N_20820);
nor U21928 (N_21928,N_20812,N_20209);
xnor U21929 (N_21929,N_19155,N_21044);
xnor U21930 (N_21930,N_19606,N_19699);
nand U21931 (N_21931,N_20741,N_19353);
nand U21932 (N_21932,N_19197,N_20815);
xor U21933 (N_21933,N_19813,N_20118);
xor U21934 (N_21934,N_20243,N_18818);
and U21935 (N_21935,N_19703,N_20844);
nand U21936 (N_21936,N_19863,N_19000);
and U21937 (N_21937,N_19417,N_20122);
nor U21938 (N_21938,N_19851,N_20483);
or U21939 (N_21939,N_21514,N_19706);
xnor U21940 (N_21940,N_19285,N_21462);
nor U21941 (N_21941,N_20041,N_19698);
xor U21942 (N_21942,N_19835,N_21120);
and U21943 (N_21943,N_19393,N_21737);
nand U21944 (N_21944,N_21688,N_20705);
and U21945 (N_21945,N_19707,N_20600);
nor U21946 (N_21946,N_19900,N_19897);
or U21947 (N_21947,N_21451,N_20199);
nor U21948 (N_21948,N_18954,N_19997);
or U21949 (N_21949,N_20025,N_18987);
or U21950 (N_21950,N_21815,N_19406);
and U21951 (N_21951,N_21183,N_20155);
nand U21952 (N_21952,N_18945,N_19094);
nor U21953 (N_21953,N_20937,N_20229);
nand U21954 (N_21954,N_20931,N_20982);
nor U21955 (N_21955,N_21114,N_20467);
nor U21956 (N_21956,N_21016,N_19758);
xor U21957 (N_21957,N_21645,N_18875);
and U21958 (N_21958,N_19574,N_20630);
nor U21959 (N_21959,N_21736,N_20030);
and U21960 (N_21960,N_21286,N_21537);
xnor U21961 (N_21961,N_21318,N_18841);
nor U21962 (N_21962,N_21424,N_19170);
xor U21963 (N_21963,N_19726,N_19842);
and U21964 (N_21964,N_19673,N_19696);
or U21965 (N_21965,N_21799,N_21542);
xnor U21966 (N_21966,N_19828,N_18976);
and U21967 (N_21967,N_20622,N_21557);
nor U21968 (N_21968,N_19923,N_21628);
or U21969 (N_21969,N_21430,N_21769);
and U21970 (N_21970,N_21580,N_18870);
and U21971 (N_21971,N_18823,N_19811);
xor U21972 (N_21972,N_20026,N_20829);
and U21973 (N_21973,N_19217,N_20091);
nor U21974 (N_21974,N_21329,N_20161);
nor U21975 (N_21975,N_21038,N_20239);
or U21976 (N_21976,N_18869,N_20384);
xnor U21977 (N_21977,N_19903,N_21500);
nand U21978 (N_21978,N_19717,N_18760);
or U21979 (N_21979,N_19099,N_21059);
nor U21980 (N_21980,N_19415,N_21352);
xor U21981 (N_21981,N_21255,N_19913);
xnor U21982 (N_21982,N_20305,N_20828);
nand U21983 (N_21983,N_20224,N_20624);
and U21984 (N_21984,N_19244,N_19605);
xnor U21985 (N_21985,N_20140,N_21844);
or U21986 (N_21986,N_20900,N_19692);
and U21987 (N_21987,N_21454,N_20468);
or U21988 (N_21988,N_19798,N_19708);
and U21989 (N_21989,N_18754,N_19365);
nor U21990 (N_21990,N_19818,N_20353);
or U21991 (N_21991,N_20880,N_20264);
nor U21992 (N_21992,N_21359,N_19057);
and U21993 (N_21993,N_19762,N_21028);
xnor U21994 (N_21994,N_21007,N_21188);
nand U21995 (N_21995,N_19737,N_20446);
nand U21996 (N_21996,N_18750,N_19753);
or U21997 (N_21997,N_19444,N_19637);
nor U21998 (N_21998,N_20307,N_20304);
nor U21999 (N_21999,N_19829,N_21381);
xnor U22000 (N_22000,N_20428,N_20870);
or U22001 (N_22001,N_20901,N_19884);
nand U22002 (N_22002,N_19777,N_21229);
nand U22003 (N_22003,N_19358,N_21407);
and U22004 (N_22004,N_20196,N_20669);
xor U22005 (N_22005,N_20036,N_20406);
or U22006 (N_22006,N_19796,N_20466);
or U22007 (N_22007,N_20075,N_19040);
nor U22008 (N_22008,N_20267,N_18828);
xnor U22009 (N_22009,N_21191,N_21728);
or U22010 (N_22010,N_21021,N_21371);
xor U22011 (N_22011,N_20516,N_20280);
nor U22012 (N_22012,N_21127,N_21148);
or U22013 (N_22013,N_20245,N_20517);
xnor U22014 (N_22014,N_19617,N_20273);
xor U22015 (N_22015,N_21778,N_21323);
or U22016 (N_22016,N_20758,N_18884);
xor U22017 (N_22017,N_18887,N_21434);
xor U22018 (N_22018,N_21609,N_21574);
or U22019 (N_22019,N_20485,N_18855);
and U22020 (N_22020,N_21608,N_19087);
and U22021 (N_22021,N_20156,N_19019);
xor U22022 (N_22022,N_20083,N_19462);
nand U22023 (N_22023,N_19723,N_20249);
and U22024 (N_22024,N_19860,N_20162);
nand U22025 (N_22025,N_20502,N_19214);
nand U22026 (N_22026,N_18952,N_19350);
nand U22027 (N_22027,N_18946,N_19715);
nand U22028 (N_22028,N_19944,N_20108);
nand U22029 (N_22029,N_20990,N_21691);
xnor U22030 (N_22030,N_21171,N_20004);
and U22031 (N_22031,N_19632,N_18764);
or U22032 (N_22032,N_19312,N_20178);
nand U22033 (N_22033,N_18799,N_21648);
nand U22034 (N_22034,N_19288,N_18775);
or U22035 (N_22035,N_21435,N_19233);
nand U22036 (N_22036,N_20848,N_20141);
xor U22037 (N_22037,N_21547,N_20651);
nor U22038 (N_22038,N_19052,N_20301);
nor U22039 (N_22039,N_18973,N_20338);
nand U22040 (N_22040,N_20659,N_20859);
or U22041 (N_22041,N_21401,N_21632);
xor U22042 (N_22042,N_20578,N_21061);
or U22043 (N_22043,N_19964,N_20970);
and U22044 (N_22044,N_20687,N_18837);
or U22045 (N_22045,N_21088,N_21106);
or U22046 (N_22046,N_21686,N_19704);
nor U22047 (N_22047,N_21009,N_19148);
xnor U22048 (N_22048,N_19167,N_18997);
nand U22049 (N_22049,N_19151,N_18774);
xor U22050 (N_22050,N_20770,N_19646);
and U22051 (N_22051,N_18988,N_19567);
nor U22052 (N_22052,N_19874,N_20792);
or U22053 (N_22053,N_18886,N_20376);
nand U22054 (N_22054,N_20015,N_19724);
nor U22055 (N_22055,N_21598,N_19306);
xnor U22056 (N_22056,N_19425,N_19808);
nor U22057 (N_22057,N_21298,N_20065);
or U22058 (N_22058,N_18939,N_21136);
xor U22059 (N_22059,N_21613,N_21477);
xor U22060 (N_22060,N_19852,N_20872);
nand U22061 (N_22061,N_21243,N_20601);
nand U22062 (N_22062,N_20103,N_21824);
nand U22063 (N_22063,N_20113,N_19668);
or U22064 (N_22064,N_20664,N_20527);
nor U22065 (N_22065,N_20274,N_21631);
or U22066 (N_22066,N_21309,N_18752);
nand U22067 (N_22067,N_20237,N_21577);
nand U22068 (N_22068,N_21792,N_21040);
nor U22069 (N_22069,N_20257,N_21703);
and U22070 (N_22070,N_20667,N_21529);
nor U22071 (N_22071,N_18766,N_21042);
nand U22072 (N_22072,N_20416,N_19321);
nand U22073 (N_22073,N_21647,N_18819);
and U22074 (N_22074,N_21419,N_19128);
nor U22075 (N_22075,N_20678,N_19581);
nor U22076 (N_22076,N_19991,N_20751);
xor U22077 (N_22077,N_21786,N_21600);
or U22078 (N_22078,N_19712,N_19603);
or U22079 (N_22079,N_20780,N_19315);
nand U22080 (N_22080,N_21013,N_21566);
nand U22081 (N_22081,N_20764,N_19002);
xor U22082 (N_22082,N_20643,N_19568);
nand U22083 (N_22083,N_19854,N_18857);
nor U22084 (N_22084,N_20185,N_20031);
nand U22085 (N_22085,N_21612,N_20377);
and U22086 (N_22086,N_20435,N_19441);
xor U22087 (N_22087,N_19806,N_20518);
and U22088 (N_22088,N_21090,N_21770);
nor U22089 (N_22089,N_21046,N_21527);
xor U22090 (N_22090,N_20555,N_21093);
xor U22091 (N_22091,N_19742,N_21867);
nor U22092 (N_22092,N_19919,N_21169);
nand U22093 (N_22093,N_20006,N_21759);
nand U22094 (N_22094,N_20801,N_20183);
nand U22095 (N_22095,N_19050,N_20135);
nand U22096 (N_22096,N_20221,N_19771);
nand U22097 (N_22097,N_19141,N_20311);
nor U22098 (N_22098,N_20124,N_21671);
nand U22099 (N_22099,N_19384,N_19994);
or U22100 (N_22100,N_20754,N_20856);
or U22101 (N_22101,N_20818,N_20519);
and U22102 (N_22102,N_21083,N_18984);
nand U22103 (N_22103,N_19586,N_20723);
nand U22104 (N_22104,N_20349,N_21094);
and U22105 (N_22105,N_20782,N_20633);
nand U22106 (N_22106,N_20379,N_21336);
and U22107 (N_22107,N_19092,N_20868);
or U22108 (N_22108,N_20440,N_20865);
xor U22109 (N_22109,N_21274,N_20064);
xor U22110 (N_22110,N_20180,N_18933);
or U22111 (N_22111,N_21170,N_18831);
or U22112 (N_22112,N_21039,N_19634);
nor U22113 (N_22113,N_20034,N_19608);
xor U22114 (N_22114,N_19982,N_19392);
or U22115 (N_22115,N_21459,N_21801);
xnor U22116 (N_22116,N_21584,N_19672);
or U22117 (N_22117,N_21279,N_19686);
xnor U22118 (N_22118,N_19754,N_20488);
nand U22119 (N_22119,N_20430,N_19270);
and U22120 (N_22120,N_20679,N_20389);
nand U22121 (N_22121,N_19477,N_19453);
nor U22122 (N_22122,N_19797,N_21396);
nor U22123 (N_22123,N_19952,N_19110);
and U22124 (N_22124,N_19885,N_21374);
xnor U22125 (N_22125,N_21767,N_19474);
nor U22126 (N_22126,N_20341,N_20743);
and U22127 (N_22127,N_21242,N_19168);
nor U22128 (N_22128,N_21414,N_20978);
and U22129 (N_22129,N_20337,N_21511);
nand U22130 (N_22130,N_18825,N_19360);
or U22131 (N_22131,N_18922,N_21139);
or U22132 (N_22132,N_19157,N_18928);
or U22133 (N_22133,N_20381,N_21256);
and U22134 (N_22134,N_21426,N_19534);
and U22135 (N_22135,N_19552,N_20340);
nand U22136 (N_22136,N_20189,N_19154);
and U22137 (N_22137,N_21828,N_18759);
or U22138 (N_22138,N_19359,N_20067);
nand U22139 (N_22139,N_20904,N_19494);
or U22140 (N_22140,N_19804,N_19053);
nand U22141 (N_22141,N_19844,N_19407);
xor U22142 (N_22142,N_21291,N_20342);
xnor U22143 (N_22143,N_19800,N_19347);
nor U22144 (N_22144,N_21670,N_21642);
xnor U22145 (N_22145,N_20954,N_20085);
or U22146 (N_22146,N_19256,N_19538);
and U22147 (N_22147,N_21490,N_20184);
nor U22148 (N_22148,N_19323,N_19104);
nand U22149 (N_22149,N_19464,N_21866);
xor U22150 (N_22150,N_20498,N_20866);
nor U22151 (N_22151,N_18969,N_18948);
or U22152 (N_22152,N_21809,N_21121);
and U22153 (N_22153,N_19594,N_19984);
and U22154 (N_22154,N_19857,N_20575);
xnor U22155 (N_22155,N_21053,N_21776);
xnor U22156 (N_22156,N_21239,N_20963);
and U22157 (N_22157,N_21651,N_21720);
nand U22158 (N_22158,N_20913,N_20763);
nand U22159 (N_22159,N_18832,N_20564);
or U22160 (N_22160,N_20942,N_20612);
and U22161 (N_22161,N_20615,N_20254);
nand U22162 (N_22162,N_20129,N_20096);
nor U22163 (N_22163,N_19005,N_19905);
xnor U22164 (N_22164,N_19228,N_19056);
nand U22165 (N_22165,N_19515,N_21304);
nor U22166 (N_22166,N_20722,N_19792);
xnor U22167 (N_22167,N_19743,N_20552);
or U22168 (N_22168,N_21162,N_20589);
and U22169 (N_22169,N_21862,N_19207);
and U22170 (N_22170,N_19388,N_21391);
nand U22171 (N_22171,N_21539,N_19372);
or U22172 (N_22172,N_21292,N_20676);
xor U22173 (N_22173,N_19473,N_19640);
and U22174 (N_22174,N_19677,N_20876);
nor U22175 (N_22175,N_20814,N_21723);
and U22176 (N_22176,N_20102,N_19071);
and U22177 (N_22177,N_21159,N_21597);
or U22178 (N_22178,N_19887,N_21128);
or U22179 (N_22179,N_18770,N_19264);
nor U22180 (N_22180,N_19898,N_19524);
xor U22181 (N_22181,N_19160,N_20852);
and U22182 (N_22182,N_21771,N_19257);
nand U22183 (N_22183,N_19076,N_20602);
nand U22184 (N_22184,N_19846,N_21060);
and U22185 (N_22185,N_20774,N_21745);
nand U22186 (N_22186,N_20699,N_19775);
or U22187 (N_22187,N_21251,N_21436);
xor U22188 (N_22188,N_20546,N_21231);
and U22189 (N_22189,N_21415,N_19017);
xnor U22190 (N_22190,N_19231,N_19279);
or U22191 (N_22191,N_19557,N_20835);
nand U22192 (N_22192,N_19625,N_20407);
xor U22193 (N_22193,N_20592,N_19506);
or U22194 (N_22194,N_19314,N_20533);
xor U22195 (N_22195,N_18991,N_19992);
and U22196 (N_22196,N_19956,N_21643);
nand U22197 (N_22197,N_20152,N_21278);
nand U22198 (N_22198,N_19072,N_21665);
and U22199 (N_22199,N_19426,N_21604);
xor U22200 (N_22200,N_20457,N_19983);
or U22201 (N_22201,N_20969,N_19117);
or U22202 (N_22202,N_20736,N_19311);
and U22203 (N_22203,N_21410,N_20449);
and U22204 (N_22204,N_21113,N_19788);
nand U22205 (N_22205,N_20262,N_19711);
xnor U22206 (N_22206,N_21143,N_19402);
nand U22207 (N_22207,N_18974,N_20604);
xnor U22208 (N_22208,N_18784,N_20839);
and U22209 (N_22209,N_19185,N_19143);
xnor U22210 (N_22210,N_19926,N_19541);
and U22211 (N_22211,N_18902,N_19065);
xnor U22212 (N_22212,N_20905,N_21476);
or U22213 (N_22213,N_19691,N_19309);
or U22214 (N_22214,N_20171,N_21213);
or U22215 (N_22215,N_18785,N_21762);
nand U22216 (N_22216,N_20345,N_21372);
xnor U22217 (N_22217,N_19122,N_18983);
or U22218 (N_22218,N_21408,N_20471);
nor U22219 (N_22219,N_21368,N_21320);
nand U22220 (N_22220,N_19739,N_20857);
or U22221 (N_22221,N_20033,N_19313);
xnor U22222 (N_22222,N_19756,N_18761);
or U22223 (N_22223,N_20186,N_21443);
nor U22224 (N_22224,N_19202,N_19179);
nand U22225 (N_22225,N_20133,N_20173);
nor U22226 (N_22226,N_20107,N_19787);
xor U22227 (N_22227,N_19664,N_20717);
nand U22228 (N_22228,N_21588,N_21035);
nand U22229 (N_22229,N_19446,N_21453);
nand U22230 (N_22230,N_19633,N_20366);
xnor U22231 (N_22231,N_21357,N_21173);
nor U22232 (N_22232,N_20760,N_21147);
xor U22233 (N_22233,N_21687,N_21194);
or U22234 (N_22234,N_18756,N_20539);
and U22235 (N_22235,N_20560,N_21413);
xor U22236 (N_22236,N_19039,N_19596);
and U22237 (N_22237,N_19918,N_19366);
xor U22238 (N_22238,N_19024,N_21364);
and U22239 (N_22239,N_21112,N_18925);
nand U22240 (N_22240,N_19239,N_19630);
or U22241 (N_22241,N_19095,N_21658);
and U22242 (N_22242,N_18794,N_21072);
nor U22243 (N_22243,N_18888,N_21783);
nor U22244 (N_22244,N_21544,N_20689);
and U22245 (N_22245,N_19631,N_19456);
nor U22246 (N_22246,N_21496,N_20040);
or U22247 (N_22247,N_20926,N_19613);
nand U22248 (N_22248,N_21019,N_19316);
xor U22249 (N_22249,N_19187,N_20029);
or U22250 (N_22250,N_20210,N_21205);
nor U22251 (N_22251,N_21474,N_19908);
nor U22252 (N_22252,N_19602,N_21807);
and U22253 (N_22253,N_21740,N_19252);
nor U22254 (N_22254,N_19182,N_21047);
xor U22255 (N_22255,N_19294,N_20074);
nand U22256 (N_22256,N_20422,N_19781);
and U22257 (N_22257,N_20965,N_19493);
nor U22258 (N_22258,N_20104,N_19871);
and U22259 (N_22259,N_19255,N_19536);
and U22260 (N_22260,N_21421,N_18773);
xor U22261 (N_22261,N_19395,N_21852);
nor U22262 (N_22262,N_19727,N_18858);
or U22263 (N_22263,N_19445,N_21513);
nor U22264 (N_22264,N_19204,N_20390);
nand U22265 (N_22265,N_20525,N_21000);
nand U22266 (N_22266,N_21795,N_21750);
xnor U22267 (N_22267,N_20120,N_20775);
nand U22268 (N_22268,N_20823,N_21222);
and U22269 (N_22269,N_19333,N_21817);
nor U22270 (N_22270,N_19853,N_20777);
nor U22271 (N_22271,N_20594,N_19577);
and U22272 (N_22272,N_21446,N_19875);
nor U22273 (N_22273,N_20863,N_21781);
nor U22274 (N_22274,N_18956,N_21860);
nand U22275 (N_22275,N_19899,N_21618);
and U22276 (N_22276,N_20629,N_19505);
or U22277 (N_22277,N_20290,N_19434);
xor U22278 (N_22278,N_21283,N_19079);
or U22279 (N_22279,N_19665,N_21025);
xor U22280 (N_22280,N_20424,N_21186);
nor U22281 (N_22281,N_20830,N_19840);
xor U22282 (N_22282,N_19888,N_19935);
nor U22283 (N_22283,N_20966,N_19153);
nand U22284 (N_22284,N_19398,N_19949);
and U22285 (N_22285,N_20748,N_21012);
xor U22286 (N_22286,N_19081,N_19376);
nand U22287 (N_22287,N_20126,N_19450);
nor U22288 (N_22288,N_19877,N_19423);
xor U22289 (N_22289,N_20690,N_20694);
xnor U22290 (N_22290,N_21714,N_20412);
nor U22291 (N_22291,N_21174,N_18763);
and U22292 (N_22292,N_19689,N_19069);
nor U22293 (N_22293,N_20553,N_20642);
or U22294 (N_22294,N_19495,N_21535);
nor U22295 (N_22295,N_19004,N_21516);
or U22296 (N_22296,N_21116,N_20144);
xor U22297 (N_22297,N_20636,N_19209);
or U22298 (N_22298,N_19123,N_20464);
nor U22299 (N_22299,N_20205,N_21322);
and U22300 (N_22300,N_20348,N_21058);
or U22301 (N_22301,N_20076,N_20153);
xnor U22302 (N_22302,N_18960,N_20778);
nor U22303 (N_22303,N_20907,N_21532);
xnor U22304 (N_22304,N_20442,N_21551);
and U22305 (N_22305,N_20663,N_19098);
nor U22306 (N_22306,N_19998,N_19995);
nand U22307 (N_22307,N_20425,N_21699);
xor U22308 (N_22308,N_20266,N_20333);
xor U22309 (N_22309,N_21383,N_19870);
nand U22310 (N_22310,N_19373,N_21842);
and U22311 (N_22311,N_18768,N_19129);
nor U22312 (N_22312,N_19149,N_21333);
or U22313 (N_22313,N_21847,N_19119);
and U22314 (N_22314,N_20403,N_20087);
nand U22315 (N_22315,N_21370,N_20732);
nand U22316 (N_22316,N_18826,N_19911);
and U22317 (N_22317,N_19560,N_20910);
nor U22318 (N_22318,N_19150,N_19188);
and U22319 (N_22319,N_20271,N_20512);
nand U22320 (N_22320,N_19046,N_20761);
nor U22321 (N_22321,N_21022,N_19237);
nor U22322 (N_22322,N_18931,N_18834);
nand U22323 (N_22323,N_19368,N_19021);
xor U22324 (N_22324,N_19165,N_21105);
nand U22325 (N_22325,N_21406,N_21196);
nand U22326 (N_22326,N_18755,N_19293);
and U22327 (N_22327,N_20671,N_19156);
or U22328 (N_22328,N_21369,N_19034);
nand U22329 (N_22329,N_21558,N_21660);
or U22330 (N_22330,N_21796,N_21538);
or U22331 (N_22331,N_19304,N_19267);
or U22332 (N_22332,N_20339,N_21846);
xor U22333 (N_22333,N_19329,N_18808);
xnor U22334 (N_22334,N_21362,N_19289);
and U22335 (N_22335,N_20577,N_20951);
nand U22336 (N_22336,N_19930,N_21829);
nand U22337 (N_22337,N_21168,N_20584);
nor U22338 (N_22338,N_18938,N_19101);
nand U22339 (N_22339,N_20220,N_21525);
or U22340 (N_22340,N_19290,N_21002);
or U22341 (N_22341,N_21611,N_20363);
nor U22342 (N_22342,N_20336,N_20716);
or U22343 (N_22343,N_19990,N_19186);
nand U22344 (N_22344,N_21076,N_18800);
and U22345 (N_22345,N_19235,N_21773);
or U22346 (N_22346,N_21793,N_21775);
or U22347 (N_22347,N_18961,N_21512);
xnor U22348 (N_22348,N_19382,N_18817);
or U22349 (N_22349,N_21394,N_19855);
nor U22350 (N_22350,N_19555,N_21638);
or U22351 (N_22351,N_21582,N_19747);
xnor U22352 (N_22352,N_18880,N_20786);
and U22353 (N_22353,N_19078,N_21308);
xor U22354 (N_22354,N_21289,N_18843);
nor U22355 (N_22355,N_21669,N_19383);
or U22356 (N_22356,N_19639,N_20912);
nand U22357 (N_22357,N_21659,N_20130);
and U22358 (N_22358,N_19283,N_21018);
or U22359 (N_22359,N_20372,N_21854);
and U22360 (N_22360,N_21478,N_20206);
xnor U22361 (N_22361,N_18993,N_18998);
nor U22362 (N_22362,N_21181,N_19868);
nand U22363 (N_22363,N_19271,N_21288);
nor U22364 (N_22364,N_18913,N_20359);
xor U22365 (N_22365,N_19736,N_21636);
xor U22366 (N_22366,N_19971,N_20095);
xnor U22367 (N_22367,N_20871,N_20843);
nand U22368 (N_22368,N_21097,N_21069);
xor U22369 (N_22369,N_20703,N_18978);
and U22370 (N_22370,N_19176,N_21839);
nor U22371 (N_22371,N_19680,N_21667);
xor U22372 (N_22372,N_21252,N_20056);
or U22373 (N_22373,N_20973,N_19500);
nand U22374 (N_22374,N_21689,N_18856);
nand U22375 (N_22375,N_20976,N_18847);
nor U22376 (N_22376,N_21700,N_21356);
or U22377 (N_22377,N_19537,N_20258);
xnor U22378 (N_22378,N_20115,N_19424);
xnor U22379 (N_22379,N_20881,N_20236);
or U22380 (N_22380,N_19447,N_20922);
nand U22381 (N_22381,N_19843,N_18916);
nand U22382 (N_22382,N_19247,N_19390);
nor U22383 (N_22383,N_18781,N_19915);
and U22384 (N_22384,N_21825,N_20724);
xor U22385 (N_22385,N_20443,N_20695);
and U22386 (N_22386,N_18804,N_20788);
or U22387 (N_22387,N_19782,N_18940);
nor U22388 (N_22388,N_20169,N_19980);
nor U22389 (N_22389,N_19807,N_19896);
nand U22390 (N_22390,N_20637,N_21550);
nor U22391 (N_22391,N_19206,N_21484);
xor U22392 (N_22392,N_21727,N_21499);
and U22393 (N_22393,N_21567,N_19542);
or U22394 (N_22394,N_20354,N_20711);
xor U22395 (N_22395,N_20314,N_21092);
nor U22396 (N_22396,N_20020,N_20360);
nor U22397 (N_22397,N_21440,N_18980);
and U22398 (N_22398,N_20677,N_19330);
nand U22399 (N_22399,N_20825,N_19124);
xnor U22400 (N_22400,N_20299,N_20005);
or U22401 (N_22401,N_21813,N_20042);
xnor U22402 (N_22402,N_21705,N_20335);
and U22403 (N_22403,N_20248,N_20369);
and U22404 (N_22404,N_21541,N_20246);
or U22405 (N_22405,N_19814,N_20579);
or U22406 (N_22406,N_20060,N_20977);
or U22407 (N_22407,N_20728,N_19381);
nand U22408 (N_22408,N_19362,N_21869);
nor U22409 (N_22409,N_18867,N_19236);
nor U22410 (N_22410,N_21505,N_19483);
or U22411 (N_22411,N_19138,N_21215);
or U22412 (N_22412,N_19909,N_21091);
or U22413 (N_22413,N_19028,N_20053);
and U22414 (N_22414,N_19970,N_19467);
or U22415 (N_22415,N_18923,N_20727);
or U22416 (N_22416,N_19478,N_20432);
nand U22417 (N_22417,N_21024,N_21258);
nor U22418 (N_22418,N_19822,N_20693);
or U22419 (N_22419,N_19501,N_20235);
nand U22420 (N_22420,N_18912,N_19295);
nand U22421 (N_22421,N_19172,N_20618);
nand U22422 (N_22422,N_21615,N_21716);
nor U22423 (N_22423,N_19009,N_21554);
or U22424 (N_22424,N_19324,N_18872);
nor U22425 (N_22425,N_21164,N_19326);
nor U22426 (N_22426,N_21133,N_21077);
nand U22427 (N_22427,N_19826,N_21548);
xnor U22428 (N_22428,N_20391,N_21652);
or U22429 (N_22429,N_19232,N_20540);
nand U22430 (N_22430,N_20987,N_20558);
xor U22431 (N_22431,N_21509,N_20674);
xnor U22432 (N_22432,N_19475,N_19589);
and U22433 (N_22433,N_20531,N_20080);
and U22434 (N_22434,N_21774,N_19163);
and U22435 (N_22435,N_19171,N_20072);
and U22436 (N_22436,N_20242,N_19859);
and U22437 (N_22437,N_20522,N_20508);
or U22438 (N_22438,N_18793,N_20569);
nand U22439 (N_22439,N_20806,N_19638);
nand U22440 (N_22440,N_20750,N_21623);
xnor U22441 (N_22441,N_20568,N_19821);
or U22442 (N_22442,N_21657,N_19073);
nor U22443 (N_22443,N_21111,N_20068);
or U22444 (N_22444,N_19027,N_20228);
nor U22445 (N_22445,N_19291,N_19675);
xor U22446 (N_22446,N_20475,N_21296);
and U22447 (N_22447,N_20585,N_19413);
or U22448 (N_22448,N_19883,N_19767);
and U22449 (N_22449,N_21065,N_20946);
xor U22450 (N_22450,N_19546,N_19275);
nand U22451 (N_22451,N_21524,N_19351);
nor U22452 (N_22452,N_21495,N_21874);
or U22453 (N_22453,N_21082,N_20000);
xor U22454 (N_22454,N_20570,N_19253);
xnor U22455 (N_22455,N_20887,N_19277);
or U22456 (N_22456,N_19340,N_21576);
nor U22457 (N_22457,N_19910,N_20992);
xor U22458 (N_22458,N_21756,N_21099);
or U22459 (N_22459,N_21684,N_19174);
and U22460 (N_22460,N_21602,N_21843);
and U22461 (N_22461,N_19922,N_21250);
or U22462 (N_22462,N_20151,N_21571);
xor U22463 (N_22463,N_19421,N_19418);
xnor U22464 (N_22464,N_18751,N_18937);
nand U22465 (N_22465,N_20465,N_21765);
nor U22466 (N_22466,N_20021,N_20644);
and U22467 (N_22467,N_20731,N_21739);
nor U22468 (N_22468,N_20459,N_21679);
nand U22469 (N_22469,N_18802,N_19459);
xor U22470 (N_22470,N_20899,N_21380);
or U22471 (N_22471,N_19953,N_21800);
xnor U22472 (N_22472,N_20477,N_20302);
nand U22473 (N_22473,N_19250,N_19022);
or U22474 (N_22474,N_20873,N_20047);
nor U22475 (N_22475,N_20841,N_20037);
nor U22476 (N_22476,N_19481,N_21870);
nand U22477 (N_22477,N_19433,N_20090);
or U22478 (N_22478,N_19773,N_21523);
nand U22479 (N_22479,N_20022,N_18934);
nor U22480 (N_22480,N_21238,N_21753);
or U22481 (N_22481,N_19612,N_19223);
xnor U22482 (N_22482,N_20947,N_19457);
or U22483 (N_22483,N_18919,N_20626);
nand U22484 (N_22484,N_20093,N_19327);
xor U22485 (N_22485,N_20528,N_19273);
and U22486 (N_22486,N_19563,N_19816);
xor U22487 (N_22487,N_18805,N_20398);
nand U22488 (N_22488,N_21693,N_21340);
or U22489 (N_22489,N_20967,N_19648);
or U22490 (N_22490,N_20240,N_19954);
nor U22491 (N_22491,N_19878,N_20395);
or U22492 (N_22492,N_21293,N_20494);
and U22493 (N_22493,N_20851,N_19619);
nand U22494 (N_22494,N_20082,N_20491);
nor U22495 (N_22495,N_20906,N_20275);
and U22496 (N_22496,N_21663,N_18942);
xor U22497 (N_22497,N_20158,N_20116);
xnor U22498 (N_22498,N_19795,N_20167);
nand U22499 (N_22499,N_20071,N_19386);
and U22500 (N_22500,N_20798,N_21485);
nor U22501 (N_22501,N_19820,N_21464);
nor U22502 (N_22502,N_20077,N_21504);
xnor U22503 (N_22503,N_21355,N_21508);
nand U22504 (N_22504,N_20561,N_21129);
and U22505 (N_22505,N_18878,N_20895);
xor U22506 (N_22506,N_21717,N_19523);
nand U22507 (N_22507,N_19713,N_19760);
and U22508 (N_22508,N_21089,N_20421);
and U22509 (N_22509,N_20172,N_19221);
and U22510 (N_22510,N_20179,N_19587);
or U22511 (N_22511,N_19108,N_20805);
and U22512 (N_22512,N_20853,N_19001);
or U22513 (N_22513,N_19765,N_20066);
or U22514 (N_22514,N_19856,N_19559);
xnor U22515 (N_22515,N_21449,N_21568);
and U22516 (N_22516,N_19337,N_21428);
or U22517 (N_22517,N_20202,N_21678);
xor U22518 (N_22518,N_20487,N_20145);
nand U22519 (N_22519,N_20526,N_19378);
nor U22520 (N_22520,N_21339,N_19419);
nor U22521 (N_22521,N_19435,N_21375);
nor U22522 (N_22522,N_21543,N_20955);
and U22523 (N_22523,N_19328,N_21721);
and U22524 (N_22524,N_19940,N_21182);
and U22525 (N_22525,N_21144,N_21849);
nand U22526 (N_22526,N_21637,N_20263);
and U22527 (N_22527,N_19272,N_20953);
nor U22528 (N_22528,N_20251,N_21855);
nand U22529 (N_22529,N_21200,N_20332);
or U22530 (N_22530,N_19136,N_20834);
and U22531 (N_22531,N_19514,N_20632);
nand U22532 (N_22532,N_19744,N_19234);
or U22533 (N_22533,N_21179,N_21095);
nor U22534 (N_22534,N_19345,N_21280);
nor U22535 (N_22535,N_20099,N_19532);
nor U22536 (N_22536,N_19580,N_21555);
nor U22537 (N_22537,N_20373,N_20890);
or U22538 (N_22538,N_20190,N_20362);
or U22539 (N_22539,N_20286,N_19759);
nand U22540 (N_22540,N_19628,N_21560);
xor U22541 (N_22541,N_19391,N_20397);
xnor U22542 (N_22542,N_20810,N_21506);
nor U22543 (N_22543,N_20110,N_19904);
or U22544 (N_22544,N_21131,N_19805);
nor U22545 (N_22545,N_21332,N_21246);
and U22546 (N_22546,N_21704,N_19082);
xnor U22547 (N_22547,N_21827,N_20523);
nor U22548 (N_22548,N_21423,N_20059);
and U22549 (N_22549,N_19023,N_18803);
and U22550 (N_22550,N_19569,N_18894);
and U22551 (N_22551,N_20358,N_21533);
or U22552 (N_22552,N_21295,N_19576);
and U22553 (N_22553,N_20799,N_21465);
nor U22554 (N_22554,N_21871,N_19011);
nor U22555 (N_22555,N_21343,N_19486);
xor U22556 (N_22556,N_19479,N_20638);
and U22557 (N_22557,N_18892,N_21119);
or U22558 (N_22558,N_19531,N_20003);
nand U22559 (N_22559,N_19029,N_19659);
xnor U22560 (N_22560,N_19089,N_20497);
and U22561 (N_22561,N_19118,N_18854);
nand U22562 (N_22562,N_21003,N_21218);
and U22563 (N_22563,N_20781,N_19296);
xor U22564 (N_22564,N_19106,N_18924);
nand U22565 (N_22565,N_19411,N_19872);
or U22566 (N_22566,N_19626,N_21306);
and U22567 (N_22567,N_19487,N_19222);
nor U22568 (N_22568,N_21303,N_18792);
xnor U22569 (N_22569,N_18986,N_18944);
or U22570 (N_22570,N_20541,N_18809);
and U22571 (N_22571,N_20392,N_19442);
nand U22572 (N_22572,N_18917,N_19730);
or U22573 (N_22573,N_18949,N_21552);
or U22574 (N_22574,N_19491,N_19458);
xnor U22575 (N_22575,N_20319,N_20745);
nand U22576 (N_22576,N_21125,N_21564);
or U22577 (N_22577,N_19091,N_21590);
nand U22578 (N_22578,N_19322,N_21675);
xnor U22579 (N_22579,N_20860,N_20084);
xnor U22580 (N_22580,N_18839,N_19729);
and U22581 (N_22581,N_21130,N_19652);
and U22582 (N_22582,N_21757,N_21232);
xor U22583 (N_22583,N_18915,N_19420);
xnor U22584 (N_22584,N_19938,N_19003);
and U22585 (N_22585,N_19030,N_20608);
xor U22586 (N_22586,N_21297,N_21045);
nor U22587 (N_22587,N_21685,N_21402);
or U22588 (N_22588,N_21545,N_20961);
xor U22589 (N_22589,N_19607,N_20445);
or U22590 (N_22590,N_20698,N_19530);
or U22591 (N_22591,N_19516,N_20755);
and U22592 (N_22592,N_19740,N_21732);
or U22593 (N_22593,N_20486,N_20012);
nand U22594 (N_22594,N_20981,N_19139);
and U22595 (N_22595,N_21835,N_19985);
or U22596 (N_22596,N_19593,N_21416);
nor U22597 (N_22597,N_19636,N_19679);
nand U22598 (N_22598,N_20444,N_19772);
and U22599 (N_22599,N_21084,N_21838);
xnor U22600 (N_22600,N_18911,N_19785);
or U22601 (N_22601,N_19305,N_21051);
nor U22602 (N_22602,N_21265,N_21442);
nand U22603 (N_22603,N_21450,N_19845);
nand U22604 (N_22604,N_20924,N_20431);
nand U22605 (N_22605,N_20737,N_18953);
xnor U22606 (N_22606,N_19578,N_20453);
nor U22607 (N_22607,N_20306,N_20598);
xor U22608 (N_22608,N_20289,N_21698);
xor U22609 (N_22609,N_19939,N_20511);
nand U22610 (N_22610,N_18968,N_19993);
nand U22611 (N_22611,N_20649,N_20989);
nor U22612 (N_22612,N_20730,N_19600);
nor U22613 (N_22613,N_21521,N_18941);
nor U22614 (N_22614,N_19437,N_20326);
or U22615 (N_22615,N_21431,N_20474);
nor U22616 (N_22616,N_20393,N_18873);
and U22617 (N_22617,N_19266,N_21534);
xnor U22618 (N_22618,N_20016,N_20735);
and U22619 (N_22619,N_19850,N_20611);
or U22620 (N_22620,N_21726,N_19770);
or U22621 (N_22621,N_21037,N_20769);
nand U22622 (N_22622,N_21719,N_19942);
nor U22623 (N_22623,N_19609,N_20148);
nand U22624 (N_22624,N_19016,N_21650);
nand U22625 (N_22625,N_20208,N_21073);
or U22626 (N_22626,N_20147,N_20673);
nor U22627 (N_22627,N_20378,N_21001);
or U22628 (N_22628,N_18900,N_19113);
xor U22629 (N_22629,N_20230,N_20504);
nand U22630 (N_22630,N_18790,N_19864);
and U22631 (N_22631,N_20874,N_20380);
and U22632 (N_22632,N_19776,N_21206);
xor U22633 (N_22633,N_19208,N_21531);
nand U22634 (N_22634,N_21692,N_21744);
and U22635 (N_22635,N_20709,N_18777);
nor U22636 (N_22636,N_19107,N_20436);
nor U22637 (N_22637,N_19461,N_21439);
or U22638 (N_22638,N_21132,N_20595);
nand U22639 (N_22639,N_19298,N_20259);
or U22640 (N_22640,N_21594,N_19145);
xor U22641 (N_22641,N_20672,N_21017);
and U22642 (N_22642,N_18830,N_20712);
nand U22643 (N_22643,N_19700,N_21857);
nand U22644 (N_22644,N_21606,N_21284);
and U22645 (N_22645,N_19669,N_19709);
and U22646 (N_22646,N_20726,N_19443);
nand U22647 (N_22647,N_18877,N_20983);
or U22648 (N_22648,N_20278,N_20999);
xor U22649 (N_22649,N_20409,N_18757);
xnor U22650 (N_22650,N_21367,N_19837);
xnor U22651 (N_22651,N_20776,N_19261);
nor U22652 (N_22652,N_21486,N_19507);
and U22653 (N_22653,N_19369,N_20019);
xor U22654 (N_22654,N_19387,N_20045);
and U22655 (N_22655,N_20893,N_20610);
xor U22656 (N_22656,N_21873,N_20696);
nand U22657 (N_22657,N_20587,N_21263);
or U22658 (N_22658,N_20452,N_18906);
nand U22659 (N_22659,N_19849,N_21491);
nand U22660 (N_22660,N_20959,N_21041);
and U22661 (N_22661,N_20284,N_19750);
xnor U22662 (N_22662,N_18797,N_19979);
nand U22663 (N_22663,N_19049,N_21747);
and U22664 (N_22664,N_20535,N_19873);
and U22665 (N_22665,N_19943,N_21317);
nor U22666 (N_22666,N_20574,N_21563);
and U22667 (N_22667,N_21152,N_21494);
xnor U22668 (N_22668,N_19439,N_19511);
xnor U22669 (N_22669,N_21520,N_20625);
nand U22670 (N_22670,N_19925,N_19663);
xnor U22671 (N_22671,N_21617,N_21335);
and U22672 (N_22672,N_19894,N_19180);
xor U22673 (N_22673,N_18885,N_19083);
nand U22674 (N_22674,N_21142,N_19768);
and U22675 (N_22675,N_21502,N_20670);
and U22676 (N_22676,N_19292,N_19428);
or U22677 (N_22677,N_20387,N_19454);
and U22678 (N_22678,N_20134,N_20729);
and U22679 (N_22679,N_19058,N_20222);
or U22680 (N_22680,N_19377,N_20675);
and U22681 (N_22681,N_20836,N_19080);
or U22682 (N_22682,N_20347,N_19074);
or U22683 (N_22683,N_20960,N_21790);
and U22684 (N_22684,N_21054,N_19549);
or U22685 (N_22685,N_18840,N_20039);
xor U22686 (N_22686,N_19015,N_21734);
nor U22687 (N_22687,N_20980,N_19476);
nor U22688 (N_22688,N_19676,N_20320);
xor U22689 (N_22689,N_19929,N_21722);
and U22690 (N_22690,N_21177,N_20499);
nor U22691 (N_22691,N_19924,N_19043);
and U22692 (N_22692,N_19695,N_20794);
nor U22693 (N_22693,N_20225,N_21241);
xor U22694 (N_22694,N_20513,N_20288);
or U22695 (N_22695,N_19597,N_20203);
and U22696 (N_22696,N_21281,N_20886);
nand U22697 (N_22697,N_18807,N_21561);
xnor U22698 (N_22698,N_21458,N_20996);
nor U22699 (N_22699,N_20367,N_20864);
nand U22700 (N_22700,N_21395,N_20382);
or U22701 (N_22701,N_19103,N_21653);
and U22702 (N_22702,N_20123,N_20923);
nor U22703 (N_22703,N_19876,N_19920);
nor U22704 (N_22704,N_19968,N_19484);
or U22705 (N_22705,N_19832,N_18829);
xor U22706 (N_22706,N_21447,N_21081);
nand U22707 (N_22707,N_21259,N_20543);
or U22708 (N_22708,N_20142,N_21411);
and U22709 (N_22709,N_20701,N_20582);
xor U22710 (N_22710,N_19431,N_18776);
and U22711 (N_22711,N_19498,N_20902);
nor U22712 (N_22712,N_19281,N_19162);
nor U22713 (N_22713,N_19794,N_20616);
nor U22714 (N_22714,N_21501,N_19950);
nor U22715 (N_22715,N_21337,N_21707);
and U22716 (N_22716,N_18848,N_19823);
nand U22717 (N_22717,N_19112,N_21230);
nand U22718 (N_22718,N_20972,N_19334);
xnor U22719 (N_22719,N_20470,N_19642);
xor U22720 (N_22720,N_21559,N_21234);
xnor U22721 (N_22721,N_21614,N_18767);
xor U22722 (N_22722,N_21070,N_20455);
xor U22723 (N_22723,N_19966,N_20481);
nor U22724 (N_22724,N_21244,N_21593);
and U22725 (N_22725,N_20495,N_20232);
nor U22726 (N_22726,N_18943,N_20562);
nand U22727 (N_22727,N_21299,N_18970);
nor U22728 (N_22728,N_20292,N_20043);
nor U22729 (N_22729,N_21625,N_21225);
or U22730 (N_22730,N_21353,N_19325);
nor U22731 (N_22731,N_21272,N_20849);
xnor U22732 (N_22732,N_19614,N_21697);
xor U22733 (N_22733,N_21237,N_21661);
and U22734 (N_22734,N_20282,N_20514);
or U22735 (N_22735,N_19685,N_19364);
or U22736 (N_22736,N_20811,N_20838);
nand U22737 (N_22737,N_20049,N_19496);
nor U22738 (N_22738,N_20450,N_21313);
nand U22739 (N_22739,N_21616,N_19621);
xor U22740 (N_22740,N_19526,N_20138);
nand U22741 (N_22741,N_21160,N_21455);
or U22742 (N_22742,N_19175,N_19133);
and U22743 (N_22743,N_20418,N_20463);
or U22744 (N_22744,N_19962,N_18862);
and U22745 (N_22745,N_21151,N_21479);
nand U22746 (N_22746,N_20009,N_20008);
nor U22747 (N_22747,N_20573,N_20563);
or U22748 (N_22748,N_21379,N_20192);
or U22749 (N_22749,N_18895,N_19455);
and U22750 (N_22750,N_20714,N_19451);
and U22751 (N_22751,N_19879,N_20460);
and U22752 (N_22752,N_21275,N_20930);
and U22753 (N_22753,N_20458,N_20175);
nor U22754 (N_22754,N_19802,N_21620);
nand U22755 (N_22755,N_19973,N_21327);
xnor U22756 (N_22756,N_20837,N_19817);
nor U22757 (N_22757,N_20888,N_20985);
or U22758 (N_22758,N_21412,N_20501);
nor U22759 (N_22759,N_21480,N_19254);
nand U22760 (N_22760,N_20200,N_20545);
and U22761 (N_22761,N_20796,N_21154);
nand U22762 (N_22762,N_19749,N_19963);
and U22763 (N_22763,N_19572,N_20882);
nor U22764 (N_22764,N_19367,N_21832);
nand U22765 (N_22765,N_20683,N_20682);
nand U22766 (N_22766,N_19553,N_20658);
or U22767 (N_22767,N_21729,N_19653);
nand U22768 (N_22768,N_19722,N_20476);
and U22769 (N_22769,N_19344,N_20063);
and U22770 (N_22770,N_21683,N_19865);
and U22771 (N_22771,N_19525,N_21388);
and U22772 (N_22772,N_20532,N_20323);
nand U22773 (N_22773,N_20803,N_19224);
nand U22774 (N_22774,N_19892,N_19485);
and U22775 (N_22775,N_20842,N_20565);
xor U22776 (N_22776,N_19410,N_18852);
and U22777 (N_22777,N_20620,N_20909);
and U22778 (N_22778,N_20896,N_20537);
and U22779 (N_22779,N_20719,N_21592);
or U22780 (N_22780,N_19622,N_20217);
and U22781 (N_22781,N_20213,N_21187);
nor U22782 (N_22782,N_21639,N_20869);
xnor U22783 (N_22783,N_21655,N_19895);
xor U22784 (N_22784,N_18962,N_21758);
or U22785 (N_22785,N_19831,N_20212);
or U22786 (N_22786,N_19591,N_19268);
or U22787 (N_22787,N_18881,N_19547);
nor U22788 (N_22788,N_19746,N_21282);
xnor U22789 (N_22789,N_19218,N_20408);
or U22790 (N_22790,N_19981,N_18822);
nor U22791 (N_22791,N_20324,N_20593);
and U22792 (N_22792,N_21360,N_21816);
and U22793 (N_22793,N_20885,N_21270);
or U22794 (N_22794,N_20219,N_19960);
nor U22795 (N_22795,N_19624,N_19867);
nor U22796 (N_22796,N_20357,N_21668);
or U22797 (N_22797,N_20111,N_18758);
and U22798 (N_22798,N_18813,N_19489);
nand U22799 (N_22799,N_21294,N_21694);
nor U22800 (N_22800,N_21165,N_20645);
or U22801 (N_22801,N_19848,N_19067);
or U22802 (N_22802,N_19183,N_19684);
nand U22803 (N_22803,N_19986,N_19482);
xor U22804 (N_22804,N_20250,N_20297);
or U22805 (N_22805,N_19585,N_19893);
and U22806 (N_22806,N_21197,N_20654);
nor U22807 (N_22807,N_21621,N_19573);
or U22808 (N_22808,N_21102,N_18882);
nand U22809 (N_22809,N_20920,N_19093);
or U22810 (N_22810,N_21300,N_20544);
and U22811 (N_22811,N_19965,N_21266);
or U22812 (N_22812,N_20309,N_21378);
and U22813 (N_22813,N_21619,N_18778);
or U22814 (N_22814,N_21109,N_20530);
xor U22815 (N_22815,N_19075,N_20260);
and U22816 (N_22816,N_21819,N_20227);
and U22817 (N_22817,N_19647,N_20797);
nor U22818 (N_22818,N_21711,N_21673);
and U22819 (N_22819,N_19006,N_18765);
or U22820 (N_22820,N_20971,N_19405);
nand U22821 (N_22821,N_21166,N_21253);
nor U22822 (N_22822,N_20374,N_21629);
xor U22823 (N_22823,N_21427,N_21797);
or U22824 (N_22824,N_18905,N_18842);
and U22825 (N_22825,N_19978,N_20136);
and U22826 (N_22826,N_20510,N_21630);
nand U22827 (N_22827,N_20789,N_19657);
nor U22828 (N_22828,N_19088,N_19125);
xor U22829 (N_22829,N_18910,N_18771);
nand U22830 (N_22830,N_20139,N_19651);
xnor U22831 (N_22831,N_18853,N_21247);
nand U22832 (N_22832,N_20294,N_19504);
or U22833 (N_22833,N_20681,N_19356);
nor U22834 (N_22834,N_20939,N_20174);
or U22835 (N_22835,N_20715,N_20069);
and U22836 (N_22836,N_19588,N_20204);
nand U22837 (N_22837,N_19308,N_20506);
and U22838 (N_22838,N_21319,N_21461);
nand U22839 (N_22839,N_21681,N_20534);
and U22840 (N_22840,N_20892,N_19246);
nand U22841 (N_22841,N_20929,N_20898);
or U22842 (N_22842,N_21399,N_21156);
nor U22843 (N_22843,N_20753,N_19032);
nor U22844 (N_22844,N_21063,N_20548);
xnor U22845 (N_22845,N_21052,N_19766);
nand U22846 (N_22846,N_19211,N_21635);
nor U22847 (N_22847,N_21644,N_19520);
nor U22848 (N_22848,N_18951,N_20554);
or U22849 (N_22849,N_19196,N_18874);
and U22850 (N_22850,N_20002,N_20388);
nand U22851 (N_22851,N_19517,N_18921);
nor U22852 (N_22852,N_20035,N_20557);
or U22853 (N_22853,N_20713,N_20884);
xnor U22854 (N_22854,N_19928,N_18861);
nor U22855 (N_22855,N_19833,N_18786);
xnor U22856 (N_22856,N_19891,N_18975);
or U22857 (N_22857,N_20597,N_19014);
and U22858 (N_22858,N_18896,N_21342);
xnor U22859 (N_22859,N_21240,N_20609);
or U22860 (N_22860,N_18927,N_19374);
nor U22861 (N_22861,N_20276,N_21315);
xor U22862 (N_22862,N_18971,N_21334);
nor U22863 (N_22863,N_19725,N_19752);
nor U22864 (N_22864,N_20321,N_20606);
nand U22865 (N_22865,N_19109,N_19720);
nand U22866 (N_22866,N_20725,N_19655);
nor U22867 (N_22867,N_19932,N_21328);
nand U22868 (N_22868,N_18868,N_19131);
nor U22869 (N_22869,N_19135,N_19318);
xor U22870 (N_22870,N_20771,N_19241);
nor U22871 (N_22871,N_20772,N_19427);
xor U22872 (N_22872,N_19120,N_20365);
or U22873 (N_22873,N_21212,N_19201);
xor U22874 (N_22874,N_20231,N_19042);
and U22875 (N_22875,N_21311,N_21746);
and U22876 (N_22876,N_19307,N_21004);
or U22877 (N_22877,N_21587,N_18990);
or U22878 (N_22878,N_20097,N_19946);
and U22879 (N_22879,N_19346,N_21487);
nor U22880 (N_22880,N_19121,N_21140);
nand U22881 (N_22881,N_19556,N_21155);
nor U22882 (N_22882,N_20410,N_19916);
xor U22883 (N_22883,N_21199,N_19535);
xnor U22884 (N_22884,N_21172,N_21350);
nor U22885 (N_22885,N_20014,N_20793);
nand U22886 (N_22886,N_20879,N_21363);
and U22887 (N_22887,N_18796,N_20787);
or U22888 (N_22888,N_19601,N_19460);
and U22889 (N_22889,N_19213,N_21386);
or U22890 (N_22890,N_20315,N_21575);
and U22891 (N_22891,N_19783,N_18889);
nor U22892 (N_22892,N_21312,N_20098);
nor U22893 (N_22893,N_20710,N_21087);
or U22894 (N_22894,N_18947,N_20596);
nand U22895 (N_22895,N_21208,N_21607);
and U22896 (N_22896,N_21358,N_21818);
and U22897 (N_22897,N_21267,N_20762);
nand U22898 (N_22898,N_19791,N_19522);
xnor U22899 (N_22899,N_20469,N_20567);
nor U22900 (N_22900,N_21601,N_20046);
nand U22901 (N_22901,N_18798,N_21831);
xnor U22902 (N_22902,N_19332,N_18936);
nor U22903 (N_22903,N_20385,N_21034);
and U22904 (N_22904,N_20051,N_19116);
xor U22905 (N_22905,N_19890,N_21314);
and U22906 (N_22906,N_21137,N_21310);
and U22907 (N_22907,N_19582,N_19641);
or U22908 (N_22908,N_21701,N_20700);
nand U22909 (N_22909,N_21808,N_20986);
nor U22910 (N_22910,N_20684,N_21064);
xor U22911 (N_22911,N_21020,N_21627);
nor U22912 (N_22912,N_21365,N_21209);
xnor U22913 (N_22913,N_20261,N_21784);
or U22914 (N_22914,N_20325,N_21749);
and U22915 (N_22915,N_21301,N_19466);
and U22916 (N_22916,N_18844,N_21822);
nand U22917 (N_22917,N_20858,N_18859);
nand U22918 (N_22918,N_19097,N_20707);
or U22919 (N_22919,N_20783,N_19799);
nand U22920 (N_22920,N_20790,N_19780);
nand U22921 (N_22921,N_20619,N_20462);
and U22922 (N_22922,N_21858,N_21696);
nor U22923 (N_22923,N_20993,N_20691);
xnor U22924 (N_22924,N_19629,N_21695);
nand U22925 (N_22925,N_20807,N_20405);
xnor U22926 (N_22926,N_20877,N_19200);
nor U22927 (N_22927,N_21316,N_19901);
nor U22928 (N_22928,N_20639,N_18779);
nor U22929 (N_22929,N_21141,N_21351);
nand U22930 (N_22930,N_19282,N_20692);
nor U22931 (N_22931,N_20176,N_20011);
xor U22932 (N_22932,N_19408,N_21706);
nor U22933 (N_22933,N_20023,N_18846);
or U22934 (N_22934,N_19169,N_19839);
xor U22935 (N_22935,N_18979,N_18864);
nand U22936 (N_22936,N_19220,N_21510);
nand U22937 (N_22937,N_21307,N_21603);
or U22938 (N_22938,N_21347,N_21709);
and U22939 (N_22939,N_21565,N_20911);
and U22940 (N_22940,N_20434,N_20244);
and U22941 (N_22941,N_20164,N_19008);
nor U22942 (N_22942,N_21497,N_19465);
nand U22943 (N_22943,N_20070,N_21204);
nand U22944 (N_22944,N_20218,N_20143);
nand U22945 (N_22945,N_20925,N_19385);
or U22946 (N_22946,N_19249,N_18982);
and U22947 (N_22947,N_19902,N_19627);
or U22948 (N_22948,N_21448,N_19357);
and U22949 (N_22949,N_21782,N_19778);
nor U22950 (N_22950,N_21540,N_21214);
or U22951 (N_22951,N_21029,N_20052);
and U22952 (N_22952,N_20168,N_21837);
nor U22953 (N_22953,N_21055,N_20188);
and U22954 (N_22954,N_20768,N_20441);
nor U22955 (N_22955,N_20300,N_20048);
xor U22956 (N_22956,N_21324,N_20415);
nand U22957 (N_22957,N_20952,N_19681);
nand U22958 (N_22958,N_19025,N_19085);
nor U22959 (N_22959,N_19660,N_20295);
nand U22960 (N_22960,N_19041,N_20505);
and U22961 (N_22961,N_21138,N_20605);
nand U22962 (N_22962,N_20657,N_20908);
and U22963 (N_22963,N_21713,N_20089);
nand U22964 (N_22964,N_19881,N_21654);
nand U22965 (N_22965,N_21223,N_21345);
nor U22966 (N_22966,N_20773,N_19610);
and U22967 (N_22967,N_19438,N_19735);
or U22968 (N_22968,N_21438,N_20507);
nand U22969 (N_22969,N_21664,N_20588);
nand U22970 (N_22970,N_19363,N_19194);
or U22971 (N_22971,N_20128,N_20688);
or U22972 (N_22972,N_20226,N_19592);
or U22973 (N_22973,N_18898,N_21518);
and U22974 (N_22974,N_21517,N_20017);
nand U22975 (N_22975,N_20094,N_19132);
nand U22976 (N_22976,N_21863,N_20627);
nand U22977 (N_22977,N_19038,N_19066);
or U22978 (N_22978,N_18753,N_20293);
nor U22979 (N_22979,N_19320,N_21189);
xnor U22980 (N_22980,N_20938,N_20472);
nor U22981 (N_22981,N_20310,N_18899);
xnor U22982 (N_22982,N_20784,N_20559);
xnor U22983 (N_22983,N_18965,N_21382);
xor U22984 (N_22984,N_19276,N_21528);
or U22985 (N_22985,N_18783,N_20988);
nand U22986 (N_22986,N_21344,N_18795);
and U22987 (N_22987,N_19917,N_19658);
nand U22988 (N_22988,N_19682,N_20013);
and U22989 (N_22989,N_19936,N_20195);
nor U22990 (N_22990,N_20964,N_21672);
nor U22991 (N_22991,N_18977,N_20438);
nor U22992 (N_22992,N_19861,N_21015);
nand U22993 (N_22993,N_19570,N_19184);
or U22994 (N_22994,N_20846,N_21195);
nand U22995 (N_22995,N_19409,N_20394);
xnor U22996 (N_22996,N_19070,N_18845);
and U22997 (N_22997,N_21268,N_19140);
xnor U22998 (N_22998,N_20915,N_21583);
and U22999 (N_22999,N_18812,N_19790);
xor U23000 (N_23000,N_21599,N_19967);
or U23001 (N_23001,N_20165,N_19810);
xnor U23002 (N_23002,N_19825,N_20994);
and U23003 (N_23003,N_21472,N_19779);
nor U23004 (N_23004,N_21325,N_21764);
nor U23005 (N_23005,N_19336,N_19731);
xnor U23006 (N_23006,N_20547,N_21074);
xor U23007 (N_23007,N_20949,N_21010);
nand U23008 (N_23008,N_19251,N_21108);
nand U23009 (N_23009,N_19972,N_19299);
or U23010 (N_23010,N_19575,N_19287);
and U23011 (N_23011,N_19240,N_19550);
and U23012 (N_23012,N_21192,N_20061);
xor U23013 (N_23013,N_20255,N_19130);
or U23014 (N_23014,N_19661,N_20117);
and U23015 (N_23015,N_19044,N_21712);
and U23016 (N_23016,N_21751,N_19934);
and U23017 (N_23017,N_21861,N_18930);
xnor U23018 (N_23018,N_20628,N_21175);
nor U23019 (N_23019,N_19248,N_19769);
and U23020 (N_23020,N_21079,N_20317);
xnor U23021 (N_23021,N_21145,N_21820);
or U23022 (N_23022,N_21596,N_20404);
or U23023 (N_23023,N_19062,N_21640);
xor U23024 (N_23024,N_21245,N_19400);
nand U23025 (N_23025,N_21507,N_18908);
nand U23026 (N_23026,N_20062,N_20451);
or U23027 (N_23027,N_21724,N_19847);
nand U23028 (N_23028,N_18996,N_20933);
and U23029 (N_23029,N_20997,N_18950);
xor U23030 (N_23030,N_19933,N_21481);
nand U23031 (N_23031,N_19077,N_20916);
nand U23032 (N_23032,N_20154,N_20826);
nor U23033 (N_23033,N_21806,N_21755);
nand U23034 (N_23034,N_19048,N_19674);
xnor U23035 (N_23035,N_20948,N_20182);
nor U23036 (N_23036,N_20583,N_19375);
and U23037 (N_23037,N_21023,N_19054);
and U23038 (N_23038,N_20800,N_19060);
and U23039 (N_23039,N_20330,N_18801);
xor U23040 (N_23040,N_19809,N_21742);
or U23041 (N_23041,N_20146,N_18814);
xor U23042 (N_23042,N_18957,N_20279);
xor U23043 (N_23043,N_19528,N_20795);
nor U23044 (N_23044,N_20429,N_21302);
nor U23045 (N_23045,N_20287,N_21226);
xnor U23046 (N_23046,N_21833,N_20328);
nand U23047 (N_23047,N_19090,N_19503);
nor U23048 (N_23048,N_19159,N_18914);
xor U23049 (N_23049,N_20647,N_21865);
xor U23050 (N_23050,N_20802,N_19502);
and U23051 (N_23051,N_21432,N_20940);
xnor U23052 (N_23052,N_20027,N_19036);
nand U23053 (N_23053,N_21216,N_20767);
xor U23054 (N_23054,N_19471,N_20044);
or U23055 (N_23055,N_21473,N_19020);
nand U23056 (N_23056,N_19355,N_20668);
or U23057 (N_23057,N_20400,N_20086);
xnor U23058 (N_23058,N_18879,N_20867);
nand U23059 (N_23059,N_21420,N_21080);
xor U23060 (N_23060,N_21043,N_20855);
and U23061 (N_23061,N_20411,N_18883);
and U23062 (N_23062,N_18850,N_19710);
nor U23063 (N_23063,N_19510,N_19564);
nor U23064 (N_23064,N_20496,N_21715);
nand U23065 (N_23065,N_18992,N_20194);
or U23066 (N_23066,N_19623,N_19190);
nor U23067 (N_23067,N_20402,N_19671);
nor U23068 (N_23068,N_21276,N_19463);
or U23069 (N_23069,N_21725,N_20749);
xor U23070 (N_23070,N_20995,N_21802);
nor U23071 (N_23071,N_18893,N_21780);
nor U23072 (N_23072,N_19068,N_21349);
xor U23073 (N_23073,N_18926,N_19697);
and U23074 (N_23074,N_20420,N_20419);
nand U23075 (N_23075,N_20277,N_21841);
or U23076 (N_23076,N_21207,N_21190);
or U23077 (N_23077,N_18964,N_19192);
nand U23078 (N_23078,N_21103,N_21262);
xnor U23079 (N_23079,N_21185,N_21134);
nand U23080 (N_23080,N_20648,N_20454);
xor U23081 (N_23081,N_20897,N_21146);
nand U23082 (N_23082,N_21662,N_21460);
nor U23083 (N_23083,N_19618,N_21354);
xnor U23084 (N_23084,N_19212,N_18772);
or U23085 (N_23085,N_19599,N_21872);
nor U23086 (N_23086,N_20473,N_21068);
or U23087 (N_23087,N_21033,N_18907);
xor U23088 (N_23088,N_19037,N_21398);
and U23089 (N_23089,N_21062,N_20914);
nand U23090 (N_23090,N_19693,N_20119);
nor U23091 (N_23091,N_20850,N_21122);
nor U23092 (N_23092,N_19988,N_20746);
nand U23093 (N_23093,N_19513,N_19999);
and U23094 (N_23094,N_21656,N_20833);
nor U23095 (N_23095,N_20296,N_21008);
and U23096 (N_23096,N_18762,N_20211);
nor U23097 (N_23097,N_20566,N_20055);
nand U23098 (N_23098,N_20331,N_21785);
nand U23099 (N_23099,N_20586,N_20928);
nand U23100 (N_23100,N_21217,N_19683);
and U23101 (N_23101,N_20414,N_20817);
xor U23102 (N_23102,N_21556,N_19866);
xnor U23103 (N_23103,N_19144,N_19352);
or U23104 (N_23104,N_18827,N_19100);
xor U23105 (N_23105,N_20322,N_21227);
and U23106 (N_23106,N_20216,N_21056);
nor U23107 (N_23107,N_20832,N_21812);
and U23108 (N_23108,N_19059,N_20740);
nor U23109 (N_23109,N_20018,N_19274);
or U23110 (N_23110,N_20413,N_20312);
and U23111 (N_23111,N_19937,N_20024);
or U23112 (N_23112,N_19958,N_21468);
xnor U23113 (N_23113,N_20542,N_19499);
nor U23114 (N_23114,N_21452,N_19258);
or U23115 (N_23115,N_20191,N_19018);
nand U23116 (N_23116,N_19278,N_21702);
nor U23117 (N_23117,N_19912,N_19595);
nand U23118 (N_23118,N_20423,N_19064);
xnor U23119 (N_23119,N_21387,N_19335);
nand U23120 (N_23120,N_21810,N_21036);
xnor U23121 (N_23121,N_19649,N_21710);
nand U23122 (N_23122,N_20538,N_20234);
and U23123 (N_23123,N_19010,N_18860);
xor U23124 (N_23124,N_21471,N_19815);
nor U23125 (N_23125,N_19562,N_19732);
nand U23126 (N_23126,N_18820,N_18963);
nor U23127 (N_23127,N_21027,N_21066);
xnor U23128 (N_23128,N_19349,N_21578);
or U23129 (N_23129,N_20549,N_19230);
or U23130 (N_23130,N_20821,N_21361);
and U23131 (N_23131,N_18863,N_19862);
xor U23132 (N_23132,N_21221,N_19644);
nor U23133 (N_23133,N_19012,N_19142);
nor U23134 (N_23134,N_19051,N_20652);
xor U23135 (N_23135,N_21743,N_20927);
or U23136 (N_23136,N_21748,N_21633);
or U23137 (N_23137,N_20550,N_21646);
nor U23138 (N_23138,N_19198,N_19527);
nand U23139 (N_23139,N_21591,N_18806);
and U23140 (N_23140,N_21086,N_19063);
and U23141 (N_23141,N_19989,N_20861);
xor U23142 (N_23142,N_19341,N_20979);
nand U23143 (N_23143,N_21048,N_19317);
xnor U23144 (N_23144,N_20752,N_20944);
xnor U23145 (N_23145,N_19134,N_20215);
or U23146 (N_23146,N_21848,N_19941);
and U23147 (N_23147,N_19219,N_19414);
or U23148 (N_23148,N_21572,N_19931);
or U23149 (N_23149,N_20785,N_20816);
or U23150 (N_23150,N_21546,N_21680);
or U23151 (N_23151,N_21851,N_19243);
xor U23152 (N_23152,N_20634,N_21075);
or U23153 (N_23153,N_18836,N_18967);
xor U23154 (N_23154,N_20490,N_21823);
nand U23155 (N_23155,N_21135,N_21107);
nor U23156 (N_23156,N_21579,N_19394);
nor U23157 (N_23157,N_20704,N_19947);
nand U23158 (N_23158,N_20193,N_19705);
or U23159 (N_23159,N_21290,N_19342);
nand U23160 (N_23160,N_20529,N_20623);
xor U23161 (N_23161,N_18891,N_20461);
or U23162 (N_23162,N_19401,N_19974);
or U23163 (N_23163,N_21220,N_20401);
and U23164 (N_23164,N_19399,N_20551);
nand U23165 (N_23165,N_21385,N_19951);
and U23166 (N_23166,N_19976,N_21124);
or U23167 (N_23167,N_21202,N_21057);
and U23168 (N_23168,N_19096,N_21526);
and U23169 (N_23169,N_20100,N_20680);
nor U23170 (N_23170,N_18966,N_19793);
nor U23171 (N_23171,N_20883,N_20247);
nand U23172 (N_23172,N_20984,N_20635);
and U23173 (N_23173,N_20875,N_18865);
or U23174 (N_23174,N_19921,N_19701);
or U23175 (N_23175,N_21338,N_20779);
nor U23176 (N_23176,N_21731,N_21264);
or U23177 (N_23177,N_19803,N_20207);
and U23178 (N_23178,N_19533,N_19229);
or U23179 (N_23179,N_19801,N_18780);
nand U23180 (N_23180,N_19225,N_21682);
nor U23181 (N_23181,N_19987,N_20607);
xnor U23182 (N_23182,N_21830,N_21158);
or U23183 (N_23183,N_18876,N_19284);
nand U23184 (N_23184,N_20088,N_21730);
xnor U23185 (N_23185,N_21733,N_21826);
and U23186 (N_23186,N_21626,N_20808);
nand U23187 (N_23187,N_20509,N_20891);
and U23188 (N_23188,N_20105,N_21798);
and U23189 (N_23189,N_19620,N_20932);
xor U23190 (N_23190,N_21779,N_21260);
or U23191 (N_23191,N_21530,N_20744);
or U23192 (N_23192,N_21466,N_21100);
nor U23193 (N_23193,N_19579,N_19379);
nor U23194 (N_23194,N_19838,N_21193);
nand U23195 (N_23195,N_20962,N_18935);
and U23196 (N_23196,N_20974,N_19819);
nor U23197 (N_23197,N_19561,N_20346);
nand U23198 (N_23198,N_20847,N_21397);
and U23199 (N_23199,N_21219,N_21634);
nor U23200 (N_23200,N_19834,N_21110);
and U23201 (N_23201,N_20520,N_19539);
and U23202 (N_23202,N_19397,N_21390);
nor U23203 (N_23203,N_21763,N_19604);
or U23204 (N_23204,N_21161,N_21211);
xor U23205 (N_23205,N_19158,N_20316);
or U23206 (N_23206,N_20734,N_19319);
nand U23207 (N_23207,N_18985,N_19127);
nor U23208 (N_23208,N_21254,N_19371);
or U23209 (N_23209,N_21811,N_21085);
nand U23210 (N_23210,N_21859,N_19216);
and U23211 (N_23211,N_20733,N_19584);
or U23212 (N_23212,N_19259,N_20170);
or U23213 (N_23213,N_20268,N_20038);
and U23214 (N_23214,N_21384,N_19102);
or U23215 (N_23215,N_19177,N_20238);
or U23216 (N_23216,N_21403,N_21488);
nor U23217 (N_23217,N_21373,N_19245);
nand U23218 (N_23218,N_20127,N_19302);
and U23219 (N_23219,N_21536,N_19280);
xor U23220 (N_23220,N_19830,N_19403);
or U23221 (N_23221,N_20187,N_20272);
and U23222 (N_23222,N_21118,N_20351);
or U23223 (N_23223,N_19195,N_19598);
nor U23224 (N_23224,N_20921,N_19654);
nor U23225 (N_23225,N_21150,N_20697);
or U23226 (N_23226,N_20641,N_20159);
xor U23227 (N_23227,N_20177,N_21115);
xnor U23228 (N_23228,N_21483,N_19061);
nand U23229 (N_23229,N_20032,N_18897);
nor U23230 (N_23230,N_19126,N_21708);
nand U23231 (N_23231,N_19687,N_20739);
xnor U23232 (N_23232,N_21184,N_21287);
nand U23233 (N_23233,N_18981,N_19858);
or U23234 (N_23234,N_20572,N_21366);
xnor U23235 (N_23235,N_19975,N_19529);
or U23236 (N_23236,N_21417,N_20368);
nand U23237 (N_23237,N_21674,N_18821);
or U23238 (N_23238,N_19173,N_20757);
and U23239 (N_23239,N_19969,N_21331);
or U23240 (N_23240,N_21248,N_19055);
nand U23241 (N_23241,N_20640,N_20650);
and U23242 (N_23242,N_21475,N_21201);
nand U23243 (N_23243,N_19440,N_20613);
nor U23244 (N_23244,N_19429,N_19763);
nor U23245 (N_23245,N_21845,N_19189);
and U23246 (N_23246,N_21498,N_21456);
xor U23247 (N_23247,N_19191,N_21178);
nand U23248 (N_23248,N_21741,N_20500);
nor U23249 (N_23249,N_20493,N_20804);
or U23250 (N_23250,N_21030,N_19227);
nand U23251 (N_23251,N_19519,N_19670);
xnor U23252 (N_23252,N_20685,N_21469);
or U23253 (N_23253,N_20738,N_19084);
nor U23254 (N_23254,N_19480,N_21515);
xnor U23255 (N_23255,N_21429,N_19662);
nor U23256 (N_23256,N_20106,N_20329);
nor U23257 (N_23257,N_19738,N_20653);
xnor U23258 (N_23258,N_19719,N_20399);
nor U23259 (N_23259,N_21389,N_20831);
nand U23260 (N_23260,N_21519,N_21049);
nor U23261 (N_23261,N_20371,N_21224);
xnor U23262 (N_23262,N_20201,N_20313);
or U23263 (N_23263,N_20197,N_18810);
nand U23264 (N_23264,N_20576,N_20081);
nand U23265 (N_23265,N_21622,N_19508);
nand U23266 (N_23266,N_21666,N_19404);
or U23267 (N_23267,N_19554,N_20822);
or U23268 (N_23268,N_21157,N_20241);
nor U23269 (N_23269,N_20489,N_19300);
xor U23270 (N_23270,N_21425,N_21649);
and U23271 (N_23271,N_18932,N_21032);
and U23272 (N_23272,N_21101,N_20166);
or U23273 (N_23273,N_21805,N_19262);
and U23274 (N_23274,N_19741,N_18901);
or U23275 (N_23275,N_19748,N_19161);
xnor U23276 (N_23276,N_19361,N_19948);
xor U23277 (N_23277,N_20935,N_20720);
and U23278 (N_23278,N_19551,N_19836);
xnor U23279 (N_23279,N_20656,N_20054);
and U23280 (N_23280,N_19755,N_19472);
nor U23281 (N_23281,N_20975,N_18999);
nand U23282 (N_23282,N_21249,N_21005);
nor U23283 (N_23283,N_21026,N_20580);
and U23284 (N_23284,N_18903,N_20447);
or U23285 (N_23285,N_20521,N_21641);
nor U23286 (N_23286,N_21814,N_20344);
nor U23287 (N_23287,N_21794,N_19303);
xnor U23288 (N_23288,N_19678,N_21735);
nor U23289 (N_23289,N_20854,N_20617);
xnor U23290 (N_23290,N_20298,N_19436);
xor U23291 (N_23291,N_20484,N_20603);
nand U23292 (N_23292,N_21078,N_19751);
xor U23293 (N_23293,N_19789,N_21437);
or U23294 (N_23294,N_20437,N_21405);
nor U23295 (N_23295,N_19396,N_20903);
and U23296 (N_23296,N_19422,N_21404);
nor U23297 (N_23297,N_21569,N_19764);
and U23298 (N_23298,N_21761,N_19370);
or U23299 (N_23299,N_20747,N_20968);
nand U23300 (N_23300,N_19389,N_19343);
or U23301 (N_23301,N_19959,N_21377);
nand U23302 (N_23302,N_19880,N_20482);
and U23303 (N_23303,N_19694,N_19114);
and U23304 (N_23304,N_21104,N_21503);
and U23305 (N_23305,N_19086,N_19199);
xnor U23306 (N_23306,N_18920,N_18788);
xnor U23307 (N_23307,N_20121,N_19714);
and U23308 (N_23308,N_19164,N_20950);
and U23309 (N_23309,N_19031,N_19656);
nor U23310 (N_23310,N_19543,N_20223);
xor U23311 (N_23311,N_21117,N_20665);
or U23312 (N_23312,N_20941,N_20515);
nand U23313 (N_23313,N_19047,N_18782);
or U23314 (N_23314,N_21392,N_20599);
xor U23315 (N_23315,N_19412,N_20265);
or U23316 (N_23316,N_19927,N_21444);
nor U23317 (N_23317,N_20114,N_19945);
and U23318 (N_23318,N_20721,N_21418);
or U23319 (N_23319,N_20010,N_21321);
or U23320 (N_23320,N_21176,N_18787);
nand U23321 (N_23321,N_19688,N_19210);
and U23322 (N_23322,N_21772,N_21522);
xor U23323 (N_23323,N_19882,N_19452);
or U23324 (N_23324,N_20655,N_21167);
or U23325 (N_23325,N_19728,N_20998);
nor U23326 (N_23326,N_20125,N_20791);
nand U23327 (N_23327,N_21011,N_20269);
or U23328 (N_23328,N_20433,N_18959);
or U23329 (N_23329,N_20092,N_19166);
xnor U23330 (N_23330,N_21031,N_21376);
xnor U23331 (N_23331,N_20478,N_20878);
nor U23332 (N_23332,N_19645,N_21738);
nand U23333 (N_23333,N_19260,N_21180);
or U23334 (N_23334,N_20318,N_19509);
or U23335 (N_23335,N_19178,N_21589);
nor U23336 (N_23336,N_20662,N_21834);
and U23337 (N_23337,N_19889,N_21006);
and U23338 (N_23338,N_18833,N_20708);
or U23339 (N_23339,N_19497,N_21856);
nand U23340 (N_23340,N_21149,N_21341);
or U23341 (N_23341,N_19518,N_18851);
xor U23342 (N_23342,N_20759,N_20918);
and U23343 (N_23343,N_21586,N_20253);
nand U23344 (N_23344,N_21277,N_19033);
nor U23345 (N_23345,N_20109,N_20150);
and U23346 (N_23346,N_21400,N_20479);
nand U23347 (N_23347,N_19146,N_21235);
xnor U23348 (N_23348,N_21305,N_19702);
or U23349 (N_23349,N_21445,N_21821);
or U23350 (N_23350,N_18866,N_21163);
xnor U23351 (N_23351,N_20396,N_21441);
or U23352 (N_23352,N_19310,N_20028);
and U23353 (N_23353,N_21096,N_20480);
xnor U23354 (N_23354,N_21840,N_19380);
nor U23355 (N_23355,N_21422,N_19540);
nor U23356 (N_23356,N_21257,N_19470);
nand U23357 (N_23357,N_20943,N_20894);
and U23358 (N_23358,N_19643,N_19339);
or U23359 (N_23359,N_19733,N_19468);
and U23360 (N_23360,N_20350,N_20383);
or U23361 (N_23361,N_19786,N_20813);
and U23362 (N_23362,N_20614,N_19013);
xnor U23363 (N_23363,N_20058,N_21126);
and U23364 (N_23364,N_19667,N_21788);
or U23365 (N_23365,N_19203,N_21595);
and U23366 (N_23366,N_20889,N_20819);
or U23367 (N_23367,N_20503,N_19650);
and U23368 (N_23368,N_20919,N_20214);
nor U23369 (N_23369,N_20101,N_21868);
and U23370 (N_23370,N_18918,N_18871);
nor U23371 (N_23371,N_20702,N_19977);
xnor U23372 (N_23372,N_20270,N_19906);
or U23373 (N_23373,N_20936,N_20352);
nand U23374 (N_23374,N_20386,N_20809);
and U23375 (N_23375,N_21326,N_19469);
nand U23376 (N_23376,N_19907,N_21853);
xnor U23377 (N_23377,N_20303,N_20581);
or U23378 (N_23378,N_19297,N_18838);
xor U23379 (N_23379,N_21718,N_20001);
and U23380 (N_23380,N_20456,N_19331);
and U23381 (N_23381,N_18958,N_20427);
nor U23382 (N_23382,N_21409,N_21198);
and U23383 (N_23383,N_20073,N_20181);
or U23384 (N_23384,N_19147,N_18811);
and U23385 (N_23385,N_19616,N_19841);
xor U23386 (N_23386,N_20252,N_18849);
nor U23387 (N_23387,N_20686,N_19827);
and U23388 (N_23388,N_21228,N_20343);
nor U23389 (N_23389,N_19784,N_19635);
nand U23390 (N_23390,N_21789,N_21492);
xor U23391 (N_23391,N_20079,N_21457);
nor U23392 (N_23392,N_19490,N_19812);
nand U23393 (N_23393,N_18815,N_19548);
and U23394 (N_23394,N_19615,N_20291);
nand U23395 (N_23395,N_19449,N_19354);
or U23396 (N_23396,N_19571,N_20840);
or U23397 (N_23397,N_21573,N_20934);
nor U23398 (N_23398,N_21203,N_21482);
or U23399 (N_23399,N_19734,N_18995);
xor U23400 (N_23400,N_20281,N_20536);
nand U23401 (N_23401,N_18835,N_18791);
or U23402 (N_23402,N_20439,N_18824);
nor U23403 (N_23403,N_20361,N_19338);
nor U23404 (N_23404,N_19961,N_19432);
and U23405 (N_23405,N_20766,N_19152);
or U23406 (N_23406,N_21271,N_20137);
or U23407 (N_23407,N_21285,N_20364);
xnor U23408 (N_23408,N_19286,N_20426);
nor U23409 (N_23409,N_20356,N_21768);
nor U23410 (N_23410,N_21261,N_19430);
and U23411 (N_23411,N_20448,N_19611);
and U23412 (N_23412,N_19226,N_19045);
or U23413 (N_23413,N_21393,N_20308);
or U23414 (N_23414,N_21804,N_19869);
nor U23415 (N_23415,N_20765,N_20355);
and U23416 (N_23416,N_20285,N_21791);
nor U23417 (N_23417,N_20621,N_20862);
nand U23418 (N_23418,N_19590,N_18769);
and U23419 (N_23419,N_19745,N_19269);
or U23420 (N_23420,N_19026,N_20050);
nor U23421 (N_23421,N_21549,N_21330);
and U23422 (N_23422,N_19512,N_20256);
nor U23423 (N_23423,N_20631,N_21348);
nand U23424 (N_23424,N_18955,N_21014);
and U23425 (N_23425,N_19265,N_21766);
and U23426 (N_23426,N_20742,N_19137);
and U23427 (N_23427,N_19774,N_20845);
nand U23428 (N_23428,N_21553,N_20524);
or U23429 (N_23429,N_21676,N_18904);
nor U23430 (N_23430,N_21470,N_21610);
and U23431 (N_23431,N_21787,N_21677);
nand U23432 (N_23432,N_20078,N_20991);
nand U23433 (N_23433,N_21585,N_20198);
and U23434 (N_23434,N_20370,N_20824);
nor U23435 (N_23435,N_19824,N_19492);
or U23436 (N_23436,N_21777,N_19914);
xor U23437 (N_23437,N_21346,N_20584);
nand U23438 (N_23438,N_20372,N_20540);
nor U23439 (N_23439,N_19456,N_19876);
or U23440 (N_23440,N_19883,N_19191);
nor U23441 (N_23441,N_19644,N_19774);
and U23442 (N_23442,N_20892,N_21293);
and U23443 (N_23443,N_21834,N_20871);
and U23444 (N_23444,N_21206,N_19864);
and U23445 (N_23445,N_20857,N_20055);
nor U23446 (N_23446,N_21542,N_20922);
and U23447 (N_23447,N_20505,N_19612);
nand U23448 (N_23448,N_21545,N_19130);
or U23449 (N_23449,N_21019,N_20266);
nand U23450 (N_23450,N_20330,N_21308);
nor U23451 (N_23451,N_20429,N_20525);
nor U23452 (N_23452,N_21022,N_21118);
xor U23453 (N_23453,N_21134,N_18945);
and U23454 (N_23454,N_20346,N_21299);
nor U23455 (N_23455,N_20419,N_19745);
nor U23456 (N_23456,N_21178,N_21241);
or U23457 (N_23457,N_19896,N_19697);
nor U23458 (N_23458,N_21428,N_21565);
nor U23459 (N_23459,N_20969,N_19987);
xor U23460 (N_23460,N_19140,N_18889);
xor U23461 (N_23461,N_19597,N_20949);
nor U23462 (N_23462,N_19051,N_20718);
and U23463 (N_23463,N_21109,N_21257);
nand U23464 (N_23464,N_19636,N_20270);
xnor U23465 (N_23465,N_20784,N_21436);
nand U23466 (N_23466,N_19352,N_18892);
nand U23467 (N_23467,N_21651,N_19588);
and U23468 (N_23468,N_20812,N_19100);
and U23469 (N_23469,N_20777,N_21402);
and U23470 (N_23470,N_21705,N_21558);
xor U23471 (N_23471,N_19560,N_21744);
and U23472 (N_23472,N_19105,N_19603);
or U23473 (N_23473,N_20230,N_19546);
or U23474 (N_23474,N_19960,N_18751);
xor U23475 (N_23475,N_21676,N_21778);
and U23476 (N_23476,N_20996,N_19129);
or U23477 (N_23477,N_20384,N_20226);
xnor U23478 (N_23478,N_20114,N_21048);
and U23479 (N_23479,N_19911,N_19438);
nor U23480 (N_23480,N_19088,N_21148);
and U23481 (N_23481,N_19982,N_21391);
or U23482 (N_23482,N_18917,N_19332);
nor U23483 (N_23483,N_19454,N_21408);
or U23484 (N_23484,N_19436,N_21224);
or U23485 (N_23485,N_20585,N_20838);
nor U23486 (N_23486,N_19648,N_21849);
and U23487 (N_23487,N_21852,N_19160);
or U23488 (N_23488,N_19192,N_18937);
xnor U23489 (N_23489,N_19472,N_21849);
or U23490 (N_23490,N_19360,N_20203);
or U23491 (N_23491,N_21738,N_20568);
and U23492 (N_23492,N_19088,N_20847);
and U23493 (N_23493,N_18845,N_21051);
nand U23494 (N_23494,N_19043,N_21857);
xor U23495 (N_23495,N_21755,N_20875);
and U23496 (N_23496,N_21852,N_21151);
nand U23497 (N_23497,N_20373,N_19505);
and U23498 (N_23498,N_20829,N_19743);
nand U23499 (N_23499,N_21592,N_20938);
and U23500 (N_23500,N_20847,N_20975);
nor U23501 (N_23501,N_18915,N_20896);
or U23502 (N_23502,N_21341,N_20873);
and U23503 (N_23503,N_20832,N_19387);
and U23504 (N_23504,N_19700,N_18920);
and U23505 (N_23505,N_21106,N_18988);
and U23506 (N_23506,N_20353,N_19923);
xor U23507 (N_23507,N_21792,N_21483);
nor U23508 (N_23508,N_21537,N_21377);
xnor U23509 (N_23509,N_21384,N_19628);
nor U23510 (N_23510,N_19473,N_19383);
and U23511 (N_23511,N_20832,N_21230);
nor U23512 (N_23512,N_20825,N_21251);
or U23513 (N_23513,N_19406,N_20402);
and U23514 (N_23514,N_20768,N_19845);
or U23515 (N_23515,N_21453,N_21347);
nand U23516 (N_23516,N_19945,N_20248);
and U23517 (N_23517,N_19205,N_20044);
nand U23518 (N_23518,N_21175,N_19740);
or U23519 (N_23519,N_20615,N_20996);
xnor U23520 (N_23520,N_18868,N_19360);
nand U23521 (N_23521,N_18896,N_20845);
xor U23522 (N_23522,N_19018,N_19651);
or U23523 (N_23523,N_21592,N_20851);
nand U23524 (N_23524,N_19672,N_21396);
nor U23525 (N_23525,N_20498,N_19979);
xnor U23526 (N_23526,N_20354,N_19194);
xnor U23527 (N_23527,N_20283,N_21459);
and U23528 (N_23528,N_20271,N_20756);
nand U23529 (N_23529,N_21071,N_21534);
nor U23530 (N_23530,N_21240,N_19573);
nor U23531 (N_23531,N_18804,N_19856);
and U23532 (N_23532,N_21394,N_20324);
nand U23533 (N_23533,N_20925,N_20529);
nand U23534 (N_23534,N_21795,N_20694);
and U23535 (N_23535,N_20430,N_21171);
and U23536 (N_23536,N_19740,N_21769);
xor U23537 (N_23537,N_18836,N_21046);
or U23538 (N_23538,N_18870,N_18770);
or U23539 (N_23539,N_20339,N_20143);
nand U23540 (N_23540,N_20458,N_20573);
nand U23541 (N_23541,N_20125,N_19431);
or U23542 (N_23542,N_21759,N_19476);
nor U23543 (N_23543,N_20117,N_19300);
nor U23544 (N_23544,N_21583,N_19901);
nand U23545 (N_23545,N_21424,N_19349);
and U23546 (N_23546,N_20644,N_20817);
nand U23547 (N_23547,N_20052,N_21063);
or U23548 (N_23548,N_21804,N_20754);
xnor U23549 (N_23549,N_19714,N_20389);
nor U23550 (N_23550,N_21611,N_19409);
nor U23551 (N_23551,N_20464,N_21110);
nand U23552 (N_23552,N_18999,N_21126);
or U23553 (N_23553,N_21546,N_20573);
or U23554 (N_23554,N_20505,N_19542);
and U23555 (N_23555,N_21554,N_21351);
or U23556 (N_23556,N_19856,N_20950);
xor U23557 (N_23557,N_21799,N_18785);
xnor U23558 (N_23558,N_19241,N_19416);
nor U23559 (N_23559,N_20883,N_19656);
and U23560 (N_23560,N_19590,N_19601);
nand U23561 (N_23561,N_18751,N_21591);
and U23562 (N_23562,N_21761,N_19603);
or U23563 (N_23563,N_20307,N_21042);
or U23564 (N_23564,N_21256,N_21558);
nand U23565 (N_23565,N_19989,N_21007);
xor U23566 (N_23566,N_21716,N_21500);
and U23567 (N_23567,N_19637,N_19076);
and U23568 (N_23568,N_19773,N_20580);
nand U23569 (N_23569,N_21486,N_21767);
nor U23570 (N_23570,N_19744,N_19829);
xor U23571 (N_23571,N_20412,N_18841);
nand U23572 (N_23572,N_20699,N_18758);
or U23573 (N_23573,N_21027,N_18805);
xnor U23574 (N_23574,N_21516,N_20944);
and U23575 (N_23575,N_20750,N_21437);
nand U23576 (N_23576,N_21521,N_18892);
xnor U23577 (N_23577,N_19380,N_19455);
xor U23578 (N_23578,N_19133,N_19252);
xor U23579 (N_23579,N_19451,N_20685);
nor U23580 (N_23580,N_20981,N_21809);
nand U23581 (N_23581,N_20915,N_19953);
nor U23582 (N_23582,N_21384,N_19685);
nor U23583 (N_23583,N_19239,N_19565);
xor U23584 (N_23584,N_21167,N_21064);
and U23585 (N_23585,N_19584,N_21385);
nand U23586 (N_23586,N_19314,N_21030);
and U23587 (N_23587,N_21197,N_18931);
nand U23588 (N_23588,N_20307,N_20297);
xnor U23589 (N_23589,N_20677,N_20833);
nand U23590 (N_23590,N_19675,N_20264);
and U23591 (N_23591,N_19123,N_18945);
nor U23592 (N_23592,N_20170,N_20597);
nand U23593 (N_23593,N_19706,N_21857);
nand U23594 (N_23594,N_19577,N_21767);
or U23595 (N_23595,N_20215,N_21243);
nor U23596 (N_23596,N_21164,N_18832);
nand U23597 (N_23597,N_19527,N_20618);
nor U23598 (N_23598,N_18779,N_20855);
nand U23599 (N_23599,N_19827,N_21739);
nand U23600 (N_23600,N_18818,N_20439);
xor U23601 (N_23601,N_21373,N_19843);
or U23602 (N_23602,N_20516,N_21315);
and U23603 (N_23603,N_21450,N_20099);
nand U23604 (N_23604,N_20462,N_21678);
and U23605 (N_23605,N_20745,N_19717);
xnor U23606 (N_23606,N_20016,N_20732);
nand U23607 (N_23607,N_19398,N_21611);
and U23608 (N_23608,N_21628,N_19461);
nor U23609 (N_23609,N_21436,N_20456);
nor U23610 (N_23610,N_20558,N_19857);
nand U23611 (N_23611,N_20079,N_21680);
or U23612 (N_23612,N_21833,N_21576);
or U23613 (N_23613,N_18996,N_21026);
or U23614 (N_23614,N_19614,N_19337);
and U23615 (N_23615,N_19488,N_21721);
nor U23616 (N_23616,N_20045,N_19697);
nor U23617 (N_23617,N_20116,N_21192);
nor U23618 (N_23618,N_21249,N_20640);
nand U23619 (N_23619,N_19748,N_20896);
nand U23620 (N_23620,N_20262,N_19013);
and U23621 (N_23621,N_19602,N_20000);
nand U23622 (N_23622,N_21701,N_20226);
xnor U23623 (N_23623,N_20384,N_19875);
and U23624 (N_23624,N_19144,N_19484);
nand U23625 (N_23625,N_20787,N_20064);
or U23626 (N_23626,N_20423,N_21192);
nor U23627 (N_23627,N_21827,N_20180);
nand U23628 (N_23628,N_21536,N_19664);
or U23629 (N_23629,N_20287,N_20279);
nor U23630 (N_23630,N_18754,N_20068);
and U23631 (N_23631,N_20765,N_21579);
nor U23632 (N_23632,N_20591,N_19357);
nor U23633 (N_23633,N_19669,N_20564);
xnor U23634 (N_23634,N_20635,N_19160);
xor U23635 (N_23635,N_20220,N_20486);
xnor U23636 (N_23636,N_18899,N_21668);
nor U23637 (N_23637,N_20824,N_20831);
nand U23638 (N_23638,N_20769,N_19128);
or U23639 (N_23639,N_19654,N_21014);
nand U23640 (N_23640,N_20354,N_20792);
nor U23641 (N_23641,N_19846,N_21555);
nor U23642 (N_23642,N_20720,N_20908);
xnor U23643 (N_23643,N_19542,N_20264);
xnor U23644 (N_23644,N_19244,N_19753);
nor U23645 (N_23645,N_21291,N_19398);
nor U23646 (N_23646,N_20266,N_21133);
nor U23647 (N_23647,N_20367,N_21306);
or U23648 (N_23648,N_20902,N_19560);
or U23649 (N_23649,N_19305,N_21662);
or U23650 (N_23650,N_21572,N_20318);
and U23651 (N_23651,N_19776,N_19912);
or U23652 (N_23652,N_20514,N_21641);
xnor U23653 (N_23653,N_20679,N_19151);
nand U23654 (N_23654,N_20699,N_21278);
xor U23655 (N_23655,N_18974,N_19152);
nand U23656 (N_23656,N_21052,N_18764);
nor U23657 (N_23657,N_19391,N_20052);
and U23658 (N_23658,N_21164,N_20205);
nand U23659 (N_23659,N_20477,N_20739);
nor U23660 (N_23660,N_21821,N_20165);
and U23661 (N_23661,N_19033,N_18797);
and U23662 (N_23662,N_20991,N_19634);
and U23663 (N_23663,N_18833,N_20495);
or U23664 (N_23664,N_19468,N_20566);
nor U23665 (N_23665,N_19408,N_20501);
xnor U23666 (N_23666,N_19863,N_21037);
nor U23667 (N_23667,N_21024,N_20458);
xnor U23668 (N_23668,N_18813,N_20640);
nand U23669 (N_23669,N_19008,N_18937);
xor U23670 (N_23670,N_20133,N_21211);
or U23671 (N_23671,N_20412,N_19959);
nand U23672 (N_23672,N_20686,N_19341);
and U23673 (N_23673,N_20359,N_19470);
nand U23674 (N_23674,N_21092,N_20367);
or U23675 (N_23675,N_19547,N_21361);
nand U23676 (N_23676,N_19924,N_19377);
or U23677 (N_23677,N_21040,N_18912);
or U23678 (N_23678,N_19992,N_21608);
xnor U23679 (N_23679,N_20793,N_21874);
nor U23680 (N_23680,N_20480,N_21505);
nor U23681 (N_23681,N_20852,N_21515);
or U23682 (N_23682,N_19868,N_20963);
nor U23683 (N_23683,N_19276,N_21866);
and U23684 (N_23684,N_20236,N_20245);
xor U23685 (N_23685,N_18831,N_20145);
nand U23686 (N_23686,N_21213,N_20533);
and U23687 (N_23687,N_20806,N_19643);
or U23688 (N_23688,N_19174,N_20712);
or U23689 (N_23689,N_21816,N_20232);
xnor U23690 (N_23690,N_20800,N_20087);
nor U23691 (N_23691,N_21160,N_18939);
and U23692 (N_23692,N_19685,N_20642);
xnor U23693 (N_23693,N_18792,N_19000);
nor U23694 (N_23694,N_19473,N_18768);
and U23695 (N_23695,N_20492,N_18871);
xnor U23696 (N_23696,N_19471,N_21709);
nand U23697 (N_23697,N_19713,N_19340);
nand U23698 (N_23698,N_21508,N_20236);
nand U23699 (N_23699,N_20822,N_19945);
and U23700 (N_23700,N_20513,N_19704);
xor U23701 (N_23701,N_19392,N_19481);
and U23702 (N_23702,N_19863,N_19405);
nor U23703 (N_23703,N_19405,N_19580);
xor U23704 (N_23704,N_20709,N_20353);
and U23705 (N_23705,N_21100,N_20265);
or U23706 (N_23706,N_19182,N_20825);
and U23707 (N_23707,N_19558,N_18970);
nand U23708 (N_23708,N_21511,N_21763);
nand U23709 (N_23709,N_20344,N_18935);
nor U23710 (N_23710,N_19467,N_21458);
xnor U23711 (N_23711,N_21015,N_19587);
xor U23712 (N_23712,N_18865,N_19234);
nand U23713 (N_23713,N_20166,N_19490);
nand U23714 (N_23714,N_20494,N_19048);
nand U23715 (N_23715,N_20935,N_19911);
or U23716 (N_23716,N_19098,N_21674);
nor U23717 (N_23717,N_20036,N_19909);
nor U23718 (N_23718,N_18921,N_19863);
nor U23719 (N_23719,N_21028,N_19568);
and U23720 (N_23720,N_19305,N_21565);
xor U23721 (N_23721,N_20653,N_19578);
or U23722 (N_23722,N_19495,N_21206);
nand U23723 (N_23723,N_19643,N_19009);
and U23724 (N_23724,N_20995,N_19133);
nor U23725 (N_23725,N_19112,N_18965);
or U23726 (N_23726,N_20909,N_19003);
nand U23727 (N_23727,N_20613,N_21083);
nor U23728 (N_23728,N_19529,N_19214);
xnor U23729 (N_23729,N_18791,N_21812);
or U23730 (N_23730,N_20734,N_20744);
and U23731 (N_23731,N_18843,N_21809);
nand U23732 (N_23732,N_20500,N_20813);
nand U23733 (N_23733,N_20930,N_21081);
nor U23734 (N_23734,N_19737,N_21109);
nor U23735 (N_23735,N_19097,N_20314);
nor U23736 (N_23736,N_21489,N_19863);
nand U23737 (N_23737,N_21597,N_20177);
or U23738 (N_23738,N_21462,N_20911);
nand U23739 (N_23739,N_19621,N_21117);
xnor U23740 (N_23740,N_21176,N_20250);
or U23741 (N_23741,N_20590,N_20618);
nand U23742 (N_23742,N_19169,N_18776);
nor U23743 (N_23743,N_21698,N_20644);
nand U23744 (N_23744,N_20692,N_19600);
nand U23745 (N_23745,N_21031,N_21573);
xor U23746 (N_23746,N_21167,N_20473);
or U23747 (N_23747,N_21471,N_19496);
xnor U23748 (N_23748,N_21537,N_19578);
nor U23749 (N_23749,N_21153,N_19353);
xnor U23750 (N_23750,N_21655,N_18811);
nand U23751 (N_23751,N_18966,N_20782);
nor U23752 (N_23752,N_19929,N_20222);
xnor U23753 (N_23753,N_20379,N_20394);
nor U23754 (N_23754,N_20416,N_20479);
nor U23755 (N_23755,N_20633,N_19452);
and U23756 (N_23756,N_20535,N_20666);
nor U23757 (N_23757,N_21007,N_21463);
or U23758 (N_23758,N_19474,N_20826);
and U23759 (N_23759,N_20525,N_18795);
and U23760 (N_23760,N_21394,N_19819);
or U23761 (N_23761,N_19002,N_20673);
xor U23762 (N_23762,N_19195,N_18947);
or U23763 (N_23763,N_20378,N_20960);
xnor U23764 (N_23764,N_20466,N_21062);
and U23765 (N_23765,N_19909,N_20669);
nor U23766 (N_23766,N_20477,N_20026);
or U23767 (N_23767,N_20743,N_19767);
nand U23768 (N_23768,N_21634,N_20308);
nor U23769 (N_23769,N_21785,N_20300);
nand U23770 (N_23770,N_18946,N_21466);
nor U23771 (N_23771,N_21457,N_19084);
or U23772 (N_23772,N_18784,N_20022);
or U23773 (N_23773,N_20344,N_20914);
nor U23774 (N_23774,N_21079,N_21437);
nand U23775 (N_23775,N_19354,N_20866);
xor U23776 (N_23776,N_20880,N_21490);
nand U23777 (N_23777,N_21290,N_20469);
and U23778 (N_23778,N_19114,N_21390);
or U23779 (N_23779,N_20380,N_19226);
nor U23780 (N_23780,N_21819,N_19660);
nor U23781 (N_23781,N_19881,N_19709);
or U23782 (N_23782,N_19976,N_19336);
nand U23783 (N_23783,N_19086,N_19672);
xnor U23784 (N_23784,N_21570,N_20321);
or U23785 (N_23785,N_19550,N_19239);
and U23786 (N_23786,N_21566,N_20507);
xor U23787 (N_23787,N_21630,N_20079);
nand U23788 (N_23788,N_20055,N_20778);
or U23789 (N_23789,N_19230,N_20174);
nor U23790 (N_23790,N_19067,N_19550);
nand U23791 (N_23791,N_20684,N_21683);
or U23792 (N_23792,N_21654,N_18919);
xnor U23793 (N_23793,N_19106,N_20894);
nor U23794 (N_23794,N_20139,N_20634);
nor U23795 (N_23795,N_20234,N_19033);
nand U23796 (N_23796,N_21185,N_20578);
or U23797 (N_23797,N_21161,N_20894);
xor U23798 (N_23798,N_20940,N_18766);
or U23799 (N_23799,N_19191,N_20359);
and U23800 (N_23800,N_19308,N_20355);
xor U23801 (N_23801,N_19869,N_19232);
xor U23802 (N_23802,N_21842,N_19781);
xor U23803 (N_23803,N_20173,N_20521);
nor U23804 (N_23804,N_19345,N_21309);
xnor U23805 (N_23805,N_19357,N_20277);
or U23806 (N_23806,N_21545,N_19305);
nor U23807 (N_23807,N_19820,N_21238);
nor U23808 (N_23808,N_20729,N_20231);
xnor U23809 (N_23809,N_21456,N_21315);
nor U23810 (N_23810,N_20659,N_20283);
nand U23811 (N_23811,N_20234,N_21065);
or U23812 (N_23812,N_20890,N_19519);
xnor U23813 (N_23813,N_19813,N_19242);
or U23814 (N_23814,N_19311,N_20883);
and U23815 (N_23815,N_20591,N_20765);
xnor U23816 (N_23816,N_21582,N_18799);
nor U23817 (N_23817,N_21400,N_21051);
nand U23818 (N_23818,N_19283,N_21111);
xnor U23819 (N_23819,N_19317,N_19821);
xnor U23820 (N_23820,N_18754,N_20288);
or U23821 (N_23821,N_19217,N_19677);
or U23822 (N_23822,N_19266,N_20695);
and U23823 (N_23823,N_18807,N_21049);
and U23824 (N_23824,N_20407,N_19925);
xor U23825 (N_23825,N_21809,N_21228);
nand U23826 (N_23826,N_21057,N_20893);
nand U23827 (N_23827,N_20463,N_20146);
nor U23828 (N_23828,N_20103,N_19947);
xnor U23829 (N_23829,N_20022,N_19324);
nand U23830 (N_23830,N_19368,N_21514);
nor U23831 (N_23831,N_20892,N_19507);
xnor U23832 (N_23832,N_20527,N_20532);
nor U23833 (N_23833,N_21766,N_20901);
nor U23834 (N_23834,N_21529,N_21434);
or U23835 (N_23835,N_21565,N_21562);
nand U23836 (N_23836,N_21128,N_21401);
xor U23837 (N_23837,N_19910,N_20760);
and U23838 (N_23838,N_21367,N_21575);
nor U23839 (N_23839,N_19760,N_21512);
or U23840 (N_23840,N_21154,N_21303);
nand U23841 (N_23841,N_18784,N_21541);
xor U23842 (N_23842,N_19193,N_20112);
nand U23843 (N_23843,N_20230,N_20442);
nand U23844 (N_23844,N_20432,N_21571);
nand U23845 (N_23845,N_19811,N_20895);
or U23846 (N_23846,N_21038,N_21420);
and U23847 (N_23847,N_21215,N_18800);
xor U23848 (N_23848,N_21429,N_20857);
or U23849 (N_23849,N_18781,N_20834);
and U23850 (N_23850,N_21065,N_19617);
or U23851 (N_23851,N_20892,N_18970);
and U23852 (N_23852,N_20520,N_19809);
nor U23853 (N_23853,N_21828,N_18878);
or U23854 (N_23854,N_19025,N_18812);
nand U23855 (N_23855,N_20650,N_19284);
xor U23856 (N_23856,N_19852,N_19403);
nand U23857 (N_23857,N_19474,N_19342);
or U23858 (N_23858,N_21434,N_21661);
and U23859 (N_23859,N_21177,N_20620);
nor U23860 (N_23860,N_20910,N_19388);
or U23861 (N_23861,N_20363,N_20269);
nor U23862 (N_23862,N_20511,N_20799);
or U23863 (N_23863,N_19119,N_21212);
nor U23864 (N_23864,N_19478,N_19637);
and U23865 (N_23865,N_19670,N_20853);
and U23866 (N_23866,N_19760,N_20723);
nand U23867 (N_23867,N_21634,N_21785);
and U23868 (N_23868,N_21142,N_21477);
xnor U23869 (N_23869,N_21715,N_20746);
and U23870 (N_23870,N_21379,N_19517);
or U23871 (N_23871,N_20607,N_18830);
nor U23872 (N_23872,N_20781,N_20876);
nor U23873 (N_23873,N_19021,N_18869);
or U23874 (N_23874,N_20838,N_20700);
nor U23875 (N_23875,N_18980,N_19526);
or U23876 (N_23876,N_21302,N_21391);
nand U23877 (N_23877,N_20583,N_19873);
and U23878 (N_23878,N_19116,N_19256);
or U23879 (N_23879,N_18774,N_20266);
xor U23880 (N_23880,N_20383,N_21590);
and U23881 (N_23881,N_20138,N_20421);
or U23882 (N_23882,N_18938,N_20998);
nor U23883 (N_23883,N_21532,N_20923);
xnor U23884 (N_23884,N_21265,N_21552);
xnor U23885 (N_23885,N_20741,N_21619);
or U23886 (N_23886,N_19913,N_21201);
and U23887 (N_23887,N_20773,N_19132);
nand U23888 (N_23888,N_19781,N_21316);
and U23889 (N_23889,N_21549,N_21803);
nor U23890 (N_23890,N_20517,N_20053);
nor U23891 (N_23891,N_19316,N_19687);
and U23892 (N_23892,N_18962,N_21050);
and U23893 (N_23893,N_21595,N_20891);
or U23894 (N_23894,N_21310,N_19624);
and U23895 (N_23895,N_20676,N_21470);
and U23896 (N_23896,N_21324,N_21244);
xor U23897 (N_23897,N_21789,N_21736);
and U23898 (N_23898,N_19304,N_19981);
xor U23899 (N_23899,N_20664,N_19946);
nand U23900 (N_23900,N_19773,N_21296);
xor U23901 (N_23901,N_20806,N_20620);
nor U23902 (N_23902,N_20792,N_18884);
nand U23903 (N_23903,N_20402,N_19168);
xnor U23904 (N_23904,N_21734,N_20035);
and U23905 (N_23905,N_19812,N_21159);
nor U23906 (N_23906,N_20981,N_19125);
xnor U23907 (N_23907,N_19048,N_18951);
and U23908 (N_23908,N_19999,N_21859);
and U23909 (N_23909,N_20841,N_20440);
xor U23910 (N_23910,N_20032,N_20172);
or U23911 (N_23911,N_21329,N_18894);
xnor U23912 (N_23912,N_21753,N_19763);
xnor U23913 (N_23913,N_19004,N_19506);
and U23914 (N_23914,N_19222,N_20232);
nor U23915 (N_23915,N_19975,N_20889);
xnor U23916 (N_23916,N_19322,N_19113);
nand U23917 (N_23917,N_21365,N_20231);
and U23918 (N_23918,N_19578,N_19296);
nor U23919 (N_23919,N_19584,N_19814);
nor U23920 (N_23920,N_20965,N_20763);
and U23921 (N_23921,N_19808,N_21256);
and U23922 (N_23922,N_21272,N_21331);
xor U23923 (N_23923,N_19584,N_18759);
nand U23924 (N_23924,N_21844,N_20661);
and U23925 (N_23925,N_21806,N_20327);
and U23926 (N_23926,N_19857,N_18969);
nand U23927 (N_23927,N_19314,N_21855);
nor U23928 (N_23928,N_19756,N_20287);
or U23929 (N_23929,N_19877,N_19927);
and U23930 (N_23930,N_21666,N_20782);
and U23931 (N_23931,N_19861,N_20189);
nand U23932 (N_23932,N_20393,N_20027);
xor U23933 (N_23933,N_19068,N_19321);
or U23934 (N_23934,N_20969,N_18912);
xnor U23935 (N_23935,N_18774,N_20492);
and U23936 (N_23936,N_20245,N_18823);
and U23937 (N_23937,N_20228,N_21863);
xnor U23938 (N_23938,N_19141,N_20908);
nand U23939 (N_23939,N_19052,N_21702);
nor U23940 (N_23940,N_20568,N_19482);
nand U23941 (N_23941,N_20489,N_21268);
or U23942 (N_23942,N_21186,N_21860);
and U23943 (N_23943,N_19348,N_19532);
nor U23944 (N_23944,N_19601,N_20198);
nor U23945 (N_23945,N_18915,N_21602);
nand U23946 (N_23946,N_21329,N_20579);
or U23947 (N_23947,N_21787,N_18923);
or U23948 (N_23948,N_20863,N_20095);
nor U23949 (N_23949,N_19938,N_19917);
and U23950 (N_23950,N_19637,N_19070);
nand U23951 (N_23951,N_21331,N_19565);
and U23952 (N_23952,N_20706,N_21475);
or U23953 (N_23953,N_19132,N_21433);
or U23954 (N_23954,N_20010,N_20227);
xnor U23955 (N_23955,N_19076,N_21524);
xnor U23956 (N_23956,N_20378,N_18922);
xor U23957 (N_23957,N_18961,N_21563);
xor U23958 (N_23958,N_21780,N_20427);
nand U23959 (N_23959,N_19513,N_19694);
and U23960 (N_23960,N_19776,N_21809);
or U23961 (N_23961,N_21079,N_19496);
nand U23962 (N_23962,N_21655,N_20634);
nand U23963 (N_23963,N_20434,N_19223);
nand U23964 (N_23964,N_19356,N_21683);
or U23965 (N_23965,N_19169,N_18873);
or U23966 (N_23966,N_19562,N_18877);
and U23967 (N_23967,N_21185,N_19173);
and U23968 (N_23968,N_21400,N_20810);
nand U23969 (N_23969,N_20414,N_21677);
xnor U23970 (N_23970,N_19627,N_20960);
nand U23971 (N_23971,N_20253,N_20322);
and U23972 (N_23972,N_21636,N_21485);
nand U23973 (N_23973,N_21504,N_21778);
xnor U23974 (N_23974,N_20445,N_20356);
or U23975 (N_23975,N_21544,N_20781);
xnor U23976 (N_23976,N_19359,N_19380);
nand U23977 (N_23977,N_21753,N_21790);
xnor U23978 (N_23978,N_21225,N_19849);
and U23979 (N_23979,N_21264,N_21127);
nor U23980 (N_23980,N_19055,N_19889);
or U23981 (N_23981,N_19336,N_20987);
and U23982 (N_23982,N_21680,N_21722);
xor U23983 (N_23983,N_20942,N_18952);
and U23984 (N_23984,N_21399,N_19488);
or U23985 (N_23985,N_21485,N_20061);
or U23986 (N_23986,N_21274,N_20353);
nand U23987 (N_23987,N_21410,N_20749);
xor U23988 (N_23988,N_20831,N_19458);
nand U23989 (N_23989,N_19578,N_20831);
or U23990 (N_23990,N_20170,N_19596);
or U23991 (N_23991,N_20427,N_20801);
nand U23992 (N_23992,N_19035,N_20299);
nor U23993 (N_23993,N_19882,N_20426);
nand U23994 (N_23994,N_18753,N_20675);
or U23995 (N_23995,N_21302,N_20704);
xnor U23996 (N_23996,N_19405,N_21487);
and U23997 (N_23997,N_19365,N_19386);
nand U23998 (N_23998,N_20255,N_21632);
nand U23999 (N_23999,N_21175,N_20220);
xnor U24000 (N_24000,N_19081,N_20789);
nor U24001 (N_24001,N_18799,N_19204);
xor U24002 (N_24002,N_19569,N_19486);
nand U24003 (N_24003,N_19264,N_20386);
or U24004 (N_24004,N_20722,N_20909);
nor U24005 (N_24005,N_21837,N_18868);
or U24006 (N_24006,N_20030,N_21312);
and U24007 (N_24007,N_21023,N_21066);
or U24008 (N_24008,N_19564,N_20571);
or U24009 (N_24009,N_20117,N_19099);
nor U24010 (N_24010,N_21793,N_19162);
nor U24011 (N_24011,N_19076,N_21558);
nand U24012 (N_24012,N_21422,N_21812);
nand U24013 (N_24013,N_19357,N_21129);
xor U24014 (N_24014,N_20977,N_19665);
nand U24015 (N_24015,N_19980,N_20858);
and U24016 (N_24016,N_20305,N_19688);
nor U24017 (N_24017,N_21793,N_21424);
xnor U24018 (N_24018,N_19894,N_20524);
nand U24019 (N_24019,N_19596,N_20682);
nand U24020 (N_24020,N_21256,N_21029);
and U24021 (N_24021,N_20840,N_21550);
nor U24022 (N_24022,N_19562,N_20558);
xor U24023 (N_24023,N_21270,N_19435);
xor U24024 (N_24024,N_19787,N_21418);
xnor U24025 (N_24025,N_19177,N_19985);
and U24026 (N_24026,N_19004,N_19307);
xnor U24027 (N_24027,N_21632,N_18921);
nand U24028 (N_24028,N_20787,N_18905);
nor U24029 (N_24029,N_21509,N_18882);
nor U24030 (N_24030,N_21354,N_19547);
nor U24031 (N_24031,N_19604,N_19880);
xor U24032 (N_24032,N_20054,N_19117);
and U24033 (N_24033,N_19210,N_19448);
nand U24034 (N_24034,N_20664,N_20167);
or U24035 (N_24035,N_19098,N_21519);
xor U24036 (N_24036,N_20359,N_21213);
nand U24037 (N_24037,N_19832,N_21226);
and U24038 (N_24038,N_19217,N_21851);
xnor U24039 (N_24039,N_20676,N_21865);
nand U24040 (N_24040,N_21134,N_20699);
nand U24041 (N_24041,N_19412,N_21788);
and U24042 (N_24042,N_19651,N_20412);
nand U24043 (N_24043,N_20747,N_21344);
nor U24044 (N_24044,N_21088,N_20498);
xnor U24045 (N_24045,N_20734,N_21827);
and U24046 (N_24046,N_20126,N_19441);
or U24047 (N_24047,N_19323,N_20442);
and U24048 (N_24048,N_19734,N_21084);
or U24049 (N_24049,N_21870,N_19075);
and U24050 (N_24050,N_21686,N_20115);
nand U24051 (N_24051,N_21674,N_21321);
or U24052 (N_24052,N_20707,N_20041);
xnor U24053 (N_24053,N_20071,N_21781);
xor U24054 (N_24054,N_20641,N_21303);
nor U24055 (N_24055,N_21619,N_18930);
and U24056 (N_24056,N_19206,N_21111);
xor U24057 (N_24057,N_19434,N_20061);
and U24058 (N_24058,N_20337,N_21212);
nor U24059 (N_24059,N_19634,N_21730);
xor U24060 (N_24060,N_21618,N_19603);
nor U24061 (N_24061,N_21795,N_19810);
and U24062 (N_24062,N_19516,N_20397);
or U24063 (N_24063,N_19926,N_19139);
and U24064 (N_24064,N_20239,N_19853);
nand U24065 (N_24065,N_19796,N_19503);
xor U24066 (N_24066,N_19088,N_20140);
nor U24067 (N_24067,N_20114,N_21260);
xor U24068 (N_24068,N_21537,N_20632);
or U24069 (N_24069,N_19795,N_21447);
or U24070 (N_24070,N_19323,N_21062);
nand U24071 (N_24071,N_20184,N_20110);
and U24072 (N_24072,N_21451,N_21233);
xor U24073 (N_24073,N_19542,N_20181);
xnor U24074 (N_24074,N_18895,N_21604);
or U24075 (N_24075,N_20358,N_20570);
and U24076 (N_24076,N_18880,N_19031);
or U24077 (N_24077,N_20560,N_19230);
nand U24078 (N_24078,N_21323,N_19539);
xor U24079 (N_24079,N_19271,N_21661);
or U24080 (N_24080,N_18869,N_20174);
nor U24081 (N_24081,N_19252,N_19075);
xor U24082 (N_24082,N_21221,N_21321);
nor U24083 (N_24083,N_19918,N_20025);
and U24084 (N_24084,N_21172,N_20833);
or U24085 (N_24085,N_21231,N_20054);
xor U24086 (N_24086,N_21335,N_21621);
nand U24087 (N_24087,N_18980,N_20366);
and U24088 (N_24088,N_19879,N_21244);
and U24089 (N_24089,N_21768,N_20638);
nor U24090 (N_24090,N_19112,N_21001);
or U24091 (N_24091,N_18968,N_21241);
xnor U24092 (N_24092,N_20969,N_20075);
xnor U24093 (N_24093,N_20837,N_19217);
nor U24094 (N_24094,N_19328,N_20248);
xor U24095 (N_24095,N_19628,N_20538);
xnor U24096 (N_24096,N_19150,N_18916);
xor U24097 (N_24097,N_20013,N_20787);
or U24098 (N_24098,N_19639,N_21009);
or U24099 (N_24099,N_20412,N_19438);
or U24100 (N_24100,N_20181,N_20674);
nand U24101 (N_24101,N_21182,N_20283);
xor U24102 (N_24102,N_20603,N_19640);
or U24103 (N_24103,N_20617,N_20097);
or U24104 (N_24104,N_19830,N_21113);
nand U24105 (N_24105,N_21610,N_20157);
nand U24106 (N_24106,N_21217,N_19718);
nand U24107 (N_24107,N_19822,N_20894);
xor U24108 (N_24108,N_21691,N_19331);
and U24109 (N_24109,N_20920,N_19877);
xor U24110 (N_24110,N_21315,N_21738);
and U24111 (N_24111,N_21802,N_19714);
nand U24112 (N_24112,N_19356,N_20314);
nor U24113 (N_24113,N_20866,N_21357);
and U24114 (N_24114,N_20205,N_19840);
and U24115 (N_24115,N_21472,N_19670);
nand U24116 (N_24116,N_19977,N_21213);
xor U24117 (N_24117,N_19253,N_19394);
nor U24118 (N_24118,N_19781,N_18757);
and U24119 (N_24119,N_19946,N_20214);
nand U24120 (N_24120,N_20049,N_21344);
and U24121 (N_24121,N_21343,N_20719);
and U24122 (N_24122,N_20690,N_20853);
xnor U24123 (N_24123,N_21224,N_21042);
nand U24124 (N_24124,N_20327,N_19312);
xnor U24125 (N_24125,N_19379,N_21074);
and U24126 (N_24126,N_20382,N_18868);
or U24127 (N_24127,N_20559,N_19130);
nand U24128 (N_24128,N_20036,N_21299);
or U24129 (N_24129,N_19089,N_19629);
nor U24130 (N_24130,N_18828,N_21599);
and U24131 (N_24131,N_21709,N_18963);
nand U24132 (N_24132,N_20015,N_21455);
or U24133 (N_24133,N_19555,N_20023);
nand U24134 (N_24134,N_20134,N_20440);
and U24135 (N_24135,N_19376,N_21069);
nand U24136 (N_24136,N_20885,N_18765);
nor U24137 (N_24137,N_19599,N_19001);
or U24138 (N_24138,N_19243,N_20082);
nand U24139 (N_24139,N_21809,N_20296);
xor U24140 (N_24140,N_19196,N_20215);
xnor U24141 (N_24141,N_21246,N_20206);
or U24142 (N_24142,N_20352,N_21097);
xnor U24143 (N_24143,N_19187,N_21109);
and U24144 (N_24144,N_21219,N_19805);
and U24145 (N_24145,N_21580,N_19232);
and U24146 (N_24146,N_20406,N_19061);
or U24147 (N_24147,N_19145,N_21744);
and U24148 (N_24148,N_18876,N_20289);
and U24149 (N_24149,N_20594,N_19964);
xor U24150 (N_24150,N_21287,N_21144);
or U24151 (N_24151,N_19147,N_20967);
nand U24152 (N_24152,N_18975,N_20084);
nor U24153 (N_24153,N_20060,N_19114);
nor U24154 (N_24154,N_21694,N_21289);
and U24155 (N_24155,N_19280,N_19794);
nor U24156 (N_24156,N_21158,N_19742);
and U24157 (N_24157,N_20594,N_21091);
nand U24158 (N_24158,N_20297,N_21244);
nand U24159 (N_24159,N_18953,N_20758);
nor U24160 (N_24160,N_20760,N_20743);
or U24161 (N_24161,N_19606,N_20022);
and U24162 (N_24162,N_19372,N_19488);
nand U24163 (N_24163,N_20084,N_20013);
nor U24164 (N_24164,N_21404,N_18919);
and U24165 (N_24165,N_19057,N_21702);
nand U24166 (N_24166,N_21779,N_18958);
nand U24167 (N_24167,N_19384,N_21017);
xnor U24168 (N_24168,N_20062,N_21741);
nand U24169 (N_24169,N_20527,N_19638);
xnor U24170 (N_24170,N_20538,N_21452);
nand U24171 (N_24171,N_19921,N_20368);
nand U24172 (N_24172,N_19972,N_20658);
or U24173 (N_24173,N_20518,N_19379);
nand U24174 (N_24174,N_19855,N_21380);
and U24175 (N_24175,N_19197,N_20372);
and U24176 (N_24176,N_20282,N_18911);
or U24177 (N_24177,N_20755,N_20389);
nor U24178 (N_24178,N_19748,N_21588);
or U24179 (N_24179,N_19078,N_21337);
or U24180 (N_24180,N_19912,N_21267);
and U24181 (N_24181,N_18872,N_18815);
or U24182 (N_24182,N_20370,N_21478);
xor U24183 (N_24183,N_20333,N_19958);
xnor U24184 (N_24184,N_19263,N_20021);
nand U24185 (N_24185,N_21717,N_19776);
nand U24186 (N_24186,N_21709,N_20775);
or U24187 (N_24187,N_21001,N_21683);
or U24188 (N_24188,N_21215,N_19859);
nor U24189 (N_24189,N_20821,N_19236);
nand U24190 (N_24190,N_21783,N_21668);
and U24191 (N_24191,N_21649,N_21217);
nor U24192 (N_24192,N_20503,N_20807);
nor U24193 (N_24193,N_19205,N_20451);
or U24194 (N_24194,N_20266,N_20256);
nand U24195 (N_24195,N_21739,N_19252);
xor U24196 (N_24196,N_20191,N_20421);
and U24197 (N_24197,N_21854,N_20412);
or U24198 (N_24198,N_19370,N_19807);
and U24199 (N_24199,N_21333,N_20410);
and U24200 (N_24200,N_19652,N_19241);
and U24201 (N_24201,N_19660,N_19723);
nor U24202 (N_24202,N_20396,N_20403);
xnor U24203 (N_24203,N_18893,N_20367);
nand U24204 (N_24204,N_20568,N_19297);
nor U24205 (N_24205,N_19182,N_19285);
or U24206 (N_24206,N_20108,N_21449);
xnor U24207 (N_24207,N_18820,N_19504);
and U24208 (N_24208,N_20143,N_21487);
nand U24209 (N_24209,N_19792,N_19013);
or U24210 (N_24210,N_21343,N_21071);
nand U24211 (N_24211,N_20665,N_21796);
nor U24212 (N_24212,N_18885,N_21722);
nand U24213 (N_24213,N_21549,N_20339);
or U24214 (N_24214,N_20045,N_19535);
and U24215 (N_24215,N_19139,N_21295);
xnor U24216 (N_24216,N_19068,N_21356);
nand U24217 (N_24217,N_21611,N_19721);
and U24218 (N_24218,N_21128,N_18990);
xor U24219 (N_24219,N_18850,N_21687);
nor U24220 (N_24220,N_19047,N_20328);
nand U24221 (N_24221,N_19517,N_18862);
xor U24222 (N_24222,N_21122,N_21298);
nor U24223 (N_24223,N_21572,N_19963);
and U24224 (N_24224,N_20998,N_19141);
nand U24225 (N_24225,N_19361,N_21248);
nand U24226 (N_24226,N_19213,N_21426);
and U24227 (N_24227,N_19918,N_19159);
and U24228 (N_24228,N_21177,N_20985);
and U24229 (N_24229,N_19329,N_20148);
xor U24230 (N_24230,N_21505,N_19470);
nand U24231 (N_24231,N_20711,N_18936);
and U24232 (N_24232,N_19813,N_20102);
nor U24233 (N_24233,N_18867,N_21554);
or U24234 (N_24234,N_21868,N_18905);
nand U24235 (N_24235,N_18922,N_19590);
nand U24236 (N_24236,N_20446,N_19974);
or U24237 (N_24237,N_21443,N_21762);
or U24238 (N_24238,N_20948,N_21455);
nor U24239 (N_24239,N_19656,N_19486);
and U24240 (N_24240,N_19513,N_20857);
xnor U24241 (N_24241,N_18984,N_21041);
or U24242 (N_24242,N_19426,N_21642);
xnor U24243 (N_24243,N_20129,N_20337);
and U24244 (N_24244,N_19329,N_19618);
nor U24245 (N_24245,N_21562,N_19495);
nor U24246 (N_24246,N_21037,N_19005);
and U24247 (N_24247,N_19148,N_19186);
xor U24248 (N_24248,N_21802,N_21321);
nor U24249 (N_24249,N_19179,N_19161);
and U24250 (N_24250,N_20752,N_19307);
or U24251 (N_24251,N_19390,N_18966);
nor U24252 (N_24252,N_20774,N_19315);
xnor U24253 (N_24253,N_21500,N_18758);
nor U24254 (N_24254,N_20708,N_20785);
nand U24255 (N_24255,N_20965,N_21766);
nand U24256 (N_24256,N_20301,N_20389);
and U24257 (N_24257,N_19323,N_21712);
nand U24258 (N_24258,N_19528,N_20492);
or U24259 (N_24259,N_21026,N_19109);
xnor U24260 (N_24260,N_19744,N_18844);
nand U24261 (N_24261,N_19278,N_21669);
nor U24262 (N_24262,N_20044,N_19289);
nor U24263 (N_24263,N_21594,N_19741);
nor U24264 (N_24264,N_19031,N_21097);
nand U24265 (N_24265,N_19160,N_18883);
or U24266 (N_24266,N_19528,N_20419);
nand U24267 (N_24267,N_20923,N_21643);
nand U24268 (N_24268,N_19246,N_19157);
xor U24269 (N_24269,N_21322,N_18868);
xor U24270 (N_24270,N_21531,N_20242);
or U24271 (N_24271,N_19745,N_21124);
xnor U24272 (N_24272,N_19817,N_20371);
nand U24273 (N_24273,N_21101,N_19159);
nor U24274 (N_24274,N_20123,N_20222);
nor U24275 (N_24275,N_20219,N_18750);
and U24276 (N_24276,N_20520,N_19915);
or U24277 (N_24277,N_20577,N_21817);
xnor U24278 (N_24278,N_21232,N_20921);
nand U24279 (N_24279,N_21123,N_19998);
or U24280 (N_24280,N_19237,N_21600);
or U24281 (N_24281,N_19414,N_21405);
or U24282 (N_24282,N_19845,N_19600);
or U24283 (N_24283,N_19386,N_20533);
nor U24284 (N_24284,N_20087,N_21872);
and U24285 (N_24285,N_21411,N_20516);
or U24286 (N_24286,N_21075,N_21156);
and U24287 (N_24287,N_21061,N_20018);
and U24288 (N_24288,N_20752,N_19965);
nand U24289 (N_24289,N_21140,N_21081);
nand U24290 (N_24290,N_21281,N_19996);
nor U24291 (N_24291,N_20083,N_20642);
xor U24292 (N_24292,N_21025,N_18984);
nor U24293 (N_24293,N_20355,N_19573);
nand U24294 (N_24294,N_21524,N_19276);
nor U24295 (N_24295,N_19105,N_19684);
nor U24296 (N_24296,N_21322,N_20319);
nand U24297 (N_24297,N_21364,N_21210);
nand U24298 (N_24298,N_18912,N_20759);
and U24299 (N_24299,N_19447,N_18779);
nand U24300 (N_24300,N_20448,N_21691);
nand U24301 (N_24301,N_21733,N_21772);
and U24302 (N_24302,N_21109,N_19631);
nand U24303 (N_24303,N_20860,N_20984);
xnor U24304 (N_24304,N_19175,N_19656);
nor U24305 (N_24305,N_21375,N_20402);
nand U24306 (N_24306,N_18827,N_20830);
or U24307 (N_24307,N_19922,N_19394);
and U24308 (N_24308,N_21653,N_19131);
nor U24309 (N_24309,N_21024,N_18868);
nor U24310 (N_24310,N_19560,N_21870);
nor U24311 (N_24311,N_19868,N_21340);
xor U24312 (N_24312,N_19828,N_21693);
xor U24313 (N_24313,N_19664,N_19738);
nand U24314 (N_24314,N_21821,N_20064);
and U24315 (N_24315,N_21743,N_21152);
nor U24316 (N_24316,N_19698,N_20082);
nand U24317 (N_24317,N_19530,N_20980);
or U24318 (N_24318,N_20067,N_20884);
xor U24319 (N_24319,N_18833,N_20764);
xor U24320 (N_24320,N_19671,N_19130);
nor U24321 (N_24321,N_19041,N_19185);
nand U24322 (N_24322,N_18941,N_21324);
nand U24323 (N_24323,N_20046,N_19331);
or U24324 (N_24324,N_19528,N_20661);
nand U24325 (N_24325,N_19116,N_19386);
and U24326 (N_24326,N_19961,N_20404);
nand U24327 (N_24327,N_20941,N_21597);
nor U24328 (N_24328,N_21262,N_19526);
and U24329 (N_24329,N_21833,N_20163);
nand U24330 (N_24330,N_18878,N_19859);
or U24331 (N_24331,N_21625,N_21557);
nand U24332 (N_24332,N_21086,N_18836);
nor U24333 (N_24333,N_18769,N_21207);
xor U24334 (N_24334,N_21017,N_20224);
xor U24335 (N_24335,N_21137,N_20488);
nor U24336 (N_24336,N_19661,N_20724);
nand U24337 (N_24337,N_19574,N_21231);
nor U24338 (N_24338,N_21524,N_19829);
nand U24339 (N_24339,N_21031,N_21618);
or U24340 (N_24340,N_20380,N_18909);
nand U24341 (N_24341,N_20592,N_19047);
nand U24342 (N_24342,N_19791,N_20660);
xnor U24343 (N_24343,N_18781,N_19948);
xor U24344 (N_24344,N_19956,N_21551);
xnor U24345 (N_24345,N_18759,N_20121);
nand U24346 (N_24346,N_20241,N_21508);
or U24347 (N_24347,N_20438,N_20579);
or U24348 (N_24348,N_21199,N_20462);
nor U24349 (N_24349,N_18822,N_18790);
or U24350 (N_24350,N_21097,N_19322);
nor U24351 (N_24351,N_21435,N_20611);
xor U24352 (N_24352,N_19905,N_19262);
nand U24353 (N_24353,N_18937,N_19321);
xor U24354 (N_24354,N_20939,N_19684);
and U24355 (N_24355,N_20224,N_20406);
nand U24356 (N_24356,N_21780,N_19484);
xnor U24357 (N_24357,N_20845,N_20377);
nor U24358 (N_24358,N_19952,N_18992);
or U24359 (N_24359,N_19974,N_19104);
nor U24360 (N_24360,N_21630,N_21485);
or U24361 (N_24361,N_19930,N_21641);
or U24362 (N_24362,N_21788,N_20667);
xnor U24363 (N_24363,N_21098,N_19397);
or U24364 (N_24364,N_19409,N_20089);
nand U24365 (N_24365,N_21672,N_21410);
or U24366 (N_24366,N_18809,N_21787);
nor U24367 (N_24367,N_20705,N_19341);
nand U24368 (N_24368,N_18807,N_19733);
xor U24369 (N_24369,N_19688,N_20021);
nor U24370 (N_24370,N_20376,N_21537);
nand U24371 (N_24371,N_20685,N_19794);
or U24372 (N_24372,N_19200,N_19986);
and U24373 (N_24373,N_19678,N_20300);
xor U24374 (N_24374,N_21179,N_19307);
or U24375 (N_24375,N_20736,N_21113);
xnor U24376 (N_24376,N_19200,N_19835);
nor U24377 (N_24377,N_20787,N_19540);
and U24378 (N_24378,N_20749,N_21785);
nand U24379 (N_24379,N_20529,N_19714);
and U24380 (N_24380,N_21199,N_21525);
xnor U24381 (N_24381,N_21136,N_20624);
nand U24382 (N_24382,N_20125,N_20295);
and U24383 (N_24383,N_20780,N_21436);
or U24384 (N_24384,N_18962,N_18920);
and U24385 (N_24385,N_21411,N_21794);
xor U24386 (N_24386,N_20269,N_20073);
xor U24387 (N_24387,N_18877,N_21187);
or U24388 (N_24388,N_20661,N_20654);
nand U24389 (N_24389,N_21145,N_21014);
and U24390 (N_24390,N_19141,N_19974);
and U24391 (N_24391,N_20974,N_21153);
xnor U24392 (N_24392,N_19658,N_20099);
nor U24393 (N_24393,N_18822,N_20621);
or U24394 (N_24394,N_19042,N_21867);
and U24395 (N_24395,N_18865,N_19714);
and U24396 (N_24396,N_20001,N_19582);
and U24397 (N_24397,N_21187,N_19248);
nor U24398 (N_24398,N_21165,N_20635);
xnor U24399 (N_24399,N_20478,N_19496);
nor U24400 (N_24400,N_20847,N_19400);
and U24401 (N_24401,N_20322,N_21402);
and U24402 (N_24402,N_20901,N_21155);
xor U24403 (N_24403,N_21873,N_18795);
xnor U24404 (N_24404,N_20182,N_19459);
or U24405 (N_24405,N_21486,N_20937);
nand U24406 (N_24406,N_19573,N_21370);
nand U24407 (N_24407,N_20408,N_21177);
nor U24408 (N_24408,N_20947,N_20481);
xor U24409 (N_24409,N_19548,N_20733);
or U24410 (N_24410,N_18882,N_19477);
xnor U24411 (N_24411,N_19724,N_21362);
xnor U24412 (N_24412,N_21800,N_20451);
and U24413 (N_24413,N_19041,N_18868);
nor U24414 (N_24414,N_21667,N_21373);
nand U24415 (N_24415,N_20166,N_18797);
or U24416 (N_24416,N_20173,N_18794);
or U24417 (N_24417,N_19053,N_19854);
xor U24418 (N_24418,N_21011,N_20144);
or U24419 (N_24419,N_20763,N_20250);
xor U24420 (N_24420,N_21586,N_20859);
xor U24421 (N_24421,N_19797,N_21819);
xnor U24422 (N_24422,N_20087,N_21152);
nand U24423 (N_24423,N_19914,N_20663);
or U24424 (N_24424,N_21607,N_18975);
and U24425 (N_24425,N_20016,N_19715);
or U24426 (N_24426,N_20762,N_21797);
or U24427 (N_24427,N_19797,N_20920);
or U24428 (N_24428,N_20322,N_18894);
nor U24429 (N_24429,N_21204,N_20942);
and U24430 (N_24430,N_21746,N_21082);
nand U24431 (N_24431,N_20471,N_20129);
nand U24432 (N_24432,N_21492,N_20760);
xor U24433 (N_24433,N_19671,N_20259);
and U24434 (N_24434,N_20973,N_19744);
nor U24435 (N_24435,N_19221,N_21512);
and U24436 (N_24436,N_19173,N_21541);
or U24437 (N_24437,N_19825,N_21496);
and U24438 (N_24438,N_21162,N_20863);
and U24439 (N_24439,N_20348,N_21851);
and U24440 (N_24440,N_19895,N_18782);
or U24441 (N_24441,N_20111,N_20883);
or U24442 (N_24442,N_20436,N_19733);
nand U24443 (N_24443,N_21490,N_21155);
or U24444 (N_24444,N_21756,N_21355);
or U24445 (N_24445,N_19415,N_21347);
xor U24446 (N_24446,N_20986,N_20979);
or U24447 (N_24447,N_21611,N_20385);
nor U24448 (N_24448,N_20539,N_20677);
or U24449 (N_24449,N_19203,N_21185);
xnor U24450 (N_24450,N_20639,N_18902);
nand U24451 (N_24451,N_19619,N_20424);
xnor U24452 (N_24452,N_19525,N_20123);
or U24453 (N_24453,N_19307,N_20259);
and U24454 (N_24454,N_20633,N_21381);
and U24455 (N_24455,N_20120,N_20639);
xor U24456 (N_24456,N_21429,N_19070);
and U24457 (N_24457,N_20781,N_21025);
or U24458 (N_24458,N_19836,N_19676);
nor U24459 (N_24459,N_20201,N_20951);
or U24460 (N_24460,N_21479,N_21288);
nand U24461 (N_24461,N_19111,N_20127);
xor U24462 (N_24462,N_19600,N_21604);
xnor U24463 (N_24463,N_19752,N_21583);
nor U24464 (N_24464,N_20223,N_20185);
and U24465 (N_24465,N_20600,N_19813);
nand U24466 (N_24466,N_21725,N_20698);
and U24467 (N_24467,N_20888,N_20393);
xnor U24468 (N_24468,N_18887,N_18776);
or U24469 (N_24469,N_20454,N_20383);
xor U24470 (N_24470,N_19378,N_20694);
xor U24471 (N_24471,N_20210,N_20168);
and U24472 (N_24472,N_20591,N_21625);
and U24473 (N_24473,N_19000,N_19011);
nand U24474 (N_24474,N_21309,N_19559);
nand U24475 (N_24475,N_21718,N_18781);
xor U24476 (N_24476,N_20747,N_21102);
or U24477 (N_24477,N_19855,N_21196);
or U24478 (N_24478,N_20903,N_20977);
or U24479 (N_24479,N_21809,N_21076);
or U24480 (N_24480,N_19478,N_18868);
xor U24481 (N_24481,N_21396,N_20805);
and U24482 (N_24482,N_21813,N_20951);
xnor U24483 (N_24483,N_20210,N_21585);
or U24484 (N_24484,N_20744,N_21008);
and U24485 (N_24485,N_21154,N_21574);
xnor U24486 (N_24486,N_21174,N_19104);
or U24487 (N_24487,N_19394,N_20900);
and U24488 (N_24488,N_20355,N_20853);
xnor U24489 (N_24489,N_21264,N_21209);
nor U24490 (N_24490,N_19509,N_19242);
and U24491 (N_24491,N_18974,N_20841);
and U24492 (N_24492,N_19842,N_18880);
nand U24493 (N_24493,N_21301,N_21145);
nand U24494 (N_24494,N_20281,N_19648);
xor U24495 (N_24495,N_19184,N_21324);
nand U24496 (N_24496,N_19301,N_20773);
and U24497 (N_24497,N_19558,N_21369);
nor U24498 (N_24498,N_19663,N_21540);
xor U24499 (N_24499,N_20414,N_19068);
nand U24500 (N_24500,N_21032,N_19753);
nor U24501 (N_24501,N_20278,N_20534);
or U24502 (N_24502,N_20592,N_20644);
xnor U24503 (N_24503,N_20947,N_21632);
nor U24504 (N_24504,N_20246,N_19095);
nor U24505 (N_24505,N_19525,N_20060);
nor U24506 (N_24506,N_19965,N_20933);
or U24507 (N_24507,N_20158,N_20944);
nor U24508 (N_24508,N_21572,N_20133);
and U24509 (N_24509,N_20484,N_19230);
nand U24510 (N_24510,N_19003,N_20824);
nand U24511 (N_24511,N_21781,N_20118);
and U24512 (N_24512,N_21759,N_19835);
or U24513 (N_24513,N_20790,N_19730);
or U24514 (N_24514,N_19016,N_20187);
nor U24515 (N_24515,N_20567,N_20823);
xnor U24516 (N_24516,N_19815,N_20200);
nand U24517 (N_24517,N_20878,N_20695);
xor U24518 (N_24518,N_19536,N_19529);
xnor U24519 (N_24519,N_21257,N_20075);
nor U24520 (N_24520,N_19476,N_19446);
xnor U24521 (N_24521,N_21662,N_19178);
nor U24522 (N_24522,N_21125,N_21793);
or U24523 (N_24523,N_20500,N_20816);
xor U24524 (N_24524,N_19571,N_21843);
nand U24525 (N_24525,N_20669,N_20334);
nand U24526 (N_24526,N_19952,N_19659);
xor U24527 (N_24527,N_21240,N_20044);
xor U24528 (N_24528,N_20731,N_20668);
xor U24529 (N_24529,N_20056,N_20294);
or U24530 (N_24530,N_19819,N_21040);
nor U24531 (N_24531,N_20301,N_19499);
or U24532 (N_24532,N_19937,N_19747);
and U24533 (N_24533,N_21858,N_19718);
and U24534 (N_24534,N_21828,N_20429);
nand U24535 (N_24535,N_20839,N_18986);
nand U24536 (N_24536,N_19228,N_19179);
nand U24537 (N_24537,N_20274,N_19722);
or U24538 (N_24538,N_19055,N_20494);
nand U24539 (N_24539,N_20389,N_19283);
xnor U24540 (N_24540,N_18914,N_19955);
xor U24541 (N_24541,N_18816,N_20965);
and U24542 (N_24542,N_19018,N_19119);
or U24543 (N_24543,N_21192,N_19867);
and U24544 (N_24544,N_19331,N_20888);
or U24545 (N_24545,N_21480,N_21482);
and U24546 (N_24546,N_20574,N_21573);
and U24547 (N_24547,N_18778,N_19937);
nand U24548 (N_24548,N_20095,N_20794);
nor U24549 (N_24549,N_21768,N_19912);
nand U24550 (N_24550,N_20070,N_19220);
or U24551 (N_24551,N_21756,N_20811);
xnor U24552 (N_24552,N_18905,N_21268);
nand U24553 (N_24553,N_20767,N_18771);
and U24554 (N_24554,N_21499,N_21504);
nor U24555 (N_24555,N_19042,N_19359);
or U24556 (N_24556,N_21766,N_19881);
nand U24557 (N_24557,N_21504,N_19336);
nor U24558 (N_24558,N_21430,N_20514);
nor U24559 (N_24559,N_19175,N_19065);
nand U24560 (N_24560,N_20028,N_21617);
and U24561 (N_24561,N_19120,N_19617);
and U24562 (N_24562,N_18764,N_21199);
xnor U24563 (N_24563,N_21715,N_21838);
xor U24564 (N_24564,N_19078,N_19243);
nand U24565 (N_24565,N_21820,N_19790);
nor U24566 (N_24566,N_18974,N_19759);
or U24567 (N_24567,N_19515,N_21179);
xnor U24568 (N_24568,N_20986,N_19610);
nand U24569 (N_24569,N_20446,N_20124);
or U24570 (N_24570,N_21229,N_20601);
or U24571 (N_24571,N_19605,N_21234);
nor U24572 (N_24572,N_19131,N_20672);
nor U24573 (N_24573,N_20204,N_21517);
nor U24574 (N_24574,N_20065,N_20616);
xnor U24575 (N_24575,N_20984,N_20684);
and U24576 (N_24576,N_19514,N_19353);
nand U24577 (N_24577,N_21033,N_20714);
nand U24578 (N_24578,N_19041,N_20527);
or U24579 (N_24579,N_21523,N_19520);
and U24580 (N_24580,N_18851,N_19725);
or U24581 (N_24581,N_21450,N_19314);
nand U24582 (N_24582,N_21853,N_20548);
or U24583 (N_24583,N_18875,N_21056);
nand U24584 (N_24584,N_21033,N_19288);
or U24585 (N_24585,N_20374,N_20777);
nand U24586 (N_24586,N_19407,N_19919);
nor U24587 (N_24587,N_21145,N_18778);
xnor U24588 (N_24588,N_21854,N_20489);
nor U24589 (N_24589,N_19666,N_20647);
and U24590 (N_24590,N_19494,N_20269);
xor U24591 (N_24591,N_20906,N_20102);
nor U24592 (N_24592,N_19783,N_21135);
or U24593 (N_24593,N_19944,N_20711);
and U24594 (N_24594,N_19299,N_21637);
nor U24595 (N_24595,N_19582,N_20579);
xor U24596 (N_24596,N_21648,N_20497);
and U24597 (N_24597,N_19279,N_20750);
and U24598 (N_24598,N_21690,N_20833);
and U24599 (N_24599,N_19502,N_19505);
and U24600 (N_24600,N_21425,N_20713);
and U24601 (N_24601,N_21753,N_18942);
nor U24602 (N_24602,N_21682,N_18962);
nand U24603 (N_24603,N_21818,N_21546);
or U24604 (N_24604,N_19745,N_20078);
nand U24605 (N_24605,N_18943,N_19066);
xor U24606 (N_24606,N_19363,N_20122);
or U24607 (N_24607,N_20171,N_19338);
nor U24608 (N_24608,N_21140,N_21064);
or U24609 (N_24609,N_20921,N_18816);
nor U24610 (N_24610,N_20859,N_20872);
xnor U24611 (N_24611,N_21488,N_18919);
nor U24612 (N_24612,N_19289,N_21225);
or U24613 (N_24613,N_21752,N_21519);
xor U24614 (N_24614,N_20364,N_19531);
nor U24615 (N_24615,N_20097,N_20834);
xnor U24616 (N_24616,N_21725,N_21776);
nand U24617 (N_24617,N_21044,N_19021);
nor U24618 (N_24618,N_20322,N_21068);
and U24619 (N_24619,N_19652,N_20201);
xnor U24620 (N_24620,N_19645,N_20419);
nand U24621 (N_24621,N_19724,N_21470);
xor U24622 (N_24622,N_21219,N_19434);
xor U24623 (N_24623,N_19243,N_19383);
or U24624 (N_24624,N_19354,N_19766);
and U24625 (N_24625,N_18947,N_19315);
nor U24626 (N_24626,N_19638,N_21552);
and U24627 (N_24627,N_21752,N_19679);
nor U24628 (N_24628,N_18837,N_19535);
and U24629 (N_24629,N_18816,N_21172);
and U24630 (N_24630,N_19467,N_21321);
nor U24631 (N_24631,N_21747,N_20292);
nand U24632 (N_24632,N_19167,N_19385);
and U24633 (N_24633,N_21306,N_21564);
and U24634 (N_24634,N_20950,N_18918);
nand U24635 (N_24635,N_21073,N_18817);
and U24636 (N_24636,N_19584,N_21187);
nand U24637 (N_24637,N_20367,N_21613);
nor U24638 (N_24638,N_19139,N_19587);
xor U24639 (N_24639,N_20136,N_20365);
nor U24640 (N_24640,N_21360,N_19328);
xor U24641 (N_24641,N_20649,N_19396);
nand U24642 (N_24642,N_20482,N_19338);
nor U24643 (N_24643,N_20202,N_19909);
xor U24644 (N_24644,N_19538,N_19168);
nand U24645 (N_24645,N_19291,N_21040);
nand U24646 (N_24646,N_20344,N_21264);
nor U24647 (N_24647,N_19131,N_19938);
or U24648 (N_24648,N_20536,N_20570);
xor U24649 (N_24649,N_20256,N_19416);
nor U24650 (N_24650,N_20731,N_21838);
nand U24651 (N_24651,N_21638,N_20937);
nor U24652 (N_24652,N_19730,N_21145);
nand U24653 (N_24653,N_21874,N_19724);
and U24654 (N_24654,N_19692,N_20735);
nor U24655 (N_24655,N_21501,N_19164);
nand U24656 (N_24656,N_19203,N_20643);
and U24657 (N_24657,N_19672,N_19007);
and U24658 (N_24658,N_20596,N_19353);
nor U24659 (N_24659,N_19761,N_19260);
or U24660 (N_24660,N_20894,N_19760);
xnor U24661 (N_24661,N_21751,N_20309);
nor U24662 (N_24662,N_21652,N_18967);
or U24663 (N_24663,N_20624,N_21809);
or U24664 (N_24664,N_20689,N_21576);
or U24665 (N_24665,N_19829,N_19684);
nand U24666 (N_24666,N_19536,N_19754);
nor U24667 (N_24667,N_19667,N_21836);
nand U24668 (N_24668,N_20470,N_20956);
and U24669 (N_24669,N_19388,N_18943);
nor U24670 (N_24670,N_19930,N_20339);
and U24671 (N_24671,N_19310,N_20821);
or U24672 (N_24672,N_21382,N_20629);
and U24673 (N_24673,N_20936,N_21732);
and U24674 (N_24674,N_18905,N_20292);
or U24675 (N_24675,N_19470,N_20531);
and U24676 (N_24676,N_21358,N_20462);
nand U24677 (N_24677,N_18979,N_21522);
and U24678 (N_24678,N_21177,N_21057);
xor U24679 (N_24679,N_18925,N_18788);
or U24680 (N_24680,N_19201,N_21609);
nand U24681 (N_24681,N_20652,N_20943);
or U24682 (N_24682,N_21448,N_20368);
nand U24683 (N_24683,N_20603,N_21441);
xnor U24684 (N_24684,N_21050,N_21394);
nor U24685 (N_24685,N_20638,N_18992);
and U24686 (N_24686,N_19706,N_19965);
and U24687 (N_24687,N_20592,N_20561);
nand U24688 (N_24688,N_18814,N_21754);
nor U24689 (N_24689,N_20812,N_18924);
or U24690 (N_24690,N_21728,N_19430);
nand U24691 (N_24691,N_21605,N_20321);
nor U24692 (N_24692,N_20182,N_20710);
or U24693 (N_24693,N_21733,N_19199);
xor U24694 (N_24694,N_20787,N_19327);
and U24695 (N_24695,N_19557,N_20620);
nand U24696 (N_24696,N_20828,N_20272);
nand U24697 (N_24697,N_19447,N_19305);
xnor U24698 (N_24698,N_19014,N_21391);
or U24699 (N_24699,N_21412,N_20116);
or U24700 (N_24700,N_21033,N_19384);
xnor U24701 (N_24701,N_19417,N_19658);
xor U24702 (N_24702,N_21157,N_19735);
and U24703 (N_24703,N_21229,N_21451);
xnor U24704 (N_24704,N_20498,N_21574);
nor U24705 (N_24705,N_18779,N_19547);
and U24706 (N_24706,N_20978,N_19619);
nor U24707 (N_24707,N_20440,N_20639);
or U24708 (N_24708,N_19520,N_19000);
and U24709 (N_24709,N_21415,N_20870);
and U24710 (N_24710,N_21308,N_20311);
or U24711 (N_24711,N_21573,N_20944);
xor U24712 (N_24712,N_19164,N_19788);
and U24713 (N_24713,N_20695,N_18892);
nor U24714 (N_24714,N_21818,N_20012);
xor U24715 (N_24715,N_19859,N_19974);
xnor U24716 (N_24716,N_19360,N_21665);
xor U24717 (N_24717,N_21368,N_20414);
nor U24718 (N_24718,N_20493,N_19159);
and U24719 (N_24719,N_18769,N_20084);
or U24720 (N_24720,N_20721,N_18899);
or U24721 (N_24721,N_19923,N_21537);
and U24722 (N_24722,N_20423,N_20331);
nor U24723 (N_24723,N_21723,N_19260);
or U24724 (N_24724,N_21779,N_21569);
xor U24725 (N_24725,N_19879,N_19324);
nand U24726 (N_24726,N_21278,N_19306);
or U24727 (N_24727,N_18931,N_18909);
xnor U24728 (N_24728,N_19883,N_20929);
and U24729 (N_24729,N_20734,N_20194);
xnor U24730 (N_24730,N_21355,N_20368);
and U24731 (N_24731,N_19322,N_21099);
or U24732 (N_24732,N_19762,N_20458);
nand U24733 (N_24733,N_19055,N_20837);
xnor U24734 (N_24734,N_21184,N_20190);
or U24735 (N_24735,N_19853,N_20607);
nor U24736 (N_24736,N_21804,N_20601);
xor U24737 (N_24737,N_19309,N_20085);
nor U24738 (N_24738,N_21103,N_20421);
nor U24739 (N_24739,N_20661,N_18989);
xnor U24740 (N_24740,N_20849,N_19725);
and U24741 (N_24741,N_21089,N_19646);
nor U24742 (N_24742,N_21298,N_19559);
xnor U24743 (N_24743,N_19773,N_20740);
nand U24744 (N_24744,N_20008,N_20982);
or U24745 (N_24745,N_19555,N_20253);
or U24746 (N_24746,N_20014,N_18974);
and U24747 (N_24747,N_20307,N_21023);
or U24748 (N_24748,N_21024,N_20424);
nand U24749 (N_24749,N_20452,N_20796);
nand U24750 (N_24750,N_21206,N_18769);
and U24751 (N_24751,N_20857,N_20721);
nand U24752 (N_24752,N_21738,N_19539);
nor U24753 (N_24753,N_20867,N_20953);
nand U24754 (N_24754,N_19395,N_20974);
nor U24755 (N_24755,N_19271,N_21587);
nor U24756 (N_24756,N_20016,N_20087);
nand U24757 (N_24757,N_21510,N_21724);
or U24758 (N_24758,N_18904,N_20570);
nor U24759 (N_24759,N_20185,N_20981);
nor U24760 (N_24760,N_21603,N_20164);
and U24761 (N_24761,N_20185,N_19052);
and U24762 (N_24762,N_20687,N_21257);
or U24763 (N_24763,N_20435,N_20134);
or U24764 (N_24764,N_18992,N_20489);
nor U24765 (N_24765,N_21342,N_19137);
and U24766 (N_24766,N_21474,N_20522);
nor U24767 (N_24767,N_18849,N_21530);
nor U24768 (N_24768,N_21538,N_20416);
or U24769 (N_24769,N_19716,N_20473);
or U24770 (N_24770,N_19158,N_21213);
or U24771 (N_24771,N_19376,N_21189);
nor U24772 (N_24772,N_19963,N_20009);
and U24773 (N_24773,N_21559,N_20146);
nor U24774 (N_24774,N_19839,N_20864);
nand U24775 (N_24775,N_20920,N_20572);
xnor U24776 (N_24776,N_19213,N_20709);
and U24777 (N_24777,N_21849,N_19428);
xnor U24778 (N_24778,N_21364,N_19481);
and U24779 (N_24779,N_19936,N_21743);
and U24780 (N_24780,N_21041,N_19556);
and U24781 (N_24781,N_19235,N_21467);
or U24782 (N_24782,N_20272,N_20713);
nor U24783 (N_24783,N_19582,N_21065);
nand U24784 (N_24784,N_20599,N_19680);
and U24785 (N_24785,N_19888,N_21336);
nand U24786 (N_24786,N_21187,N_21573);
nand U24787 (N_24787,N_20810,N_19277);
xnor U24788 (N_24788,N_20917,N_21853);
or U24789 (N_24789,N_18996,N_19681);
xor U24790 (N_24790,N_21081,N_21576);
nor U24791 (N_24791,N_21072,N_19567);
xnor U24792 (N_24792,N_19211,N_20546);
xnor U24793 (N_24793,N_20155,N_21815);
and U24794 (N_24794,N_21705,N_20929);
nand U24795 (N_24795,N_20335,N_21552);
nand U24796 (N_24796,N_20021,N_20607);
nor U24797 (N_24797,N_21497,N_20091);
or U24798 (N_24798,N_20221,N_18852);
nor U24799 (N_24799,N_20863,N_21841);
nor U24800 (N_24800,N_20244,N_20868);
xnor U24801 (N_24801,N_19656,N_21688);
xnor U24802 (N_24802,N_19679,N_19818);
xnor U24803 (N_24803,N_19909,N_19213);
xnor U24804 (N_24804,N_20233,N_20185);
or U24805 (N_24805,N_20556,N_18865);
xor U24806 (N_24806,N_19267,N_21703);
or U24807 (N_24807,N_20447,N_20474);
nor U24808 (N_24808,N_20455,N_20248);
nor U24809 (N_24809,N_21834,N_20943);
and U24810 (N_24810,N_19721,N_20738);
nand U24811 (N_24811,N_20975,N_21412);
nor U24812 (N_24812,N_21681,N_19053);
and U24813 (N_24813,N_20116,N_20326);
nor U24814 (N_24814,N_20614,N_19016);
and U24815 (N_24815,N_20957,N_19194);
and U24816 (N_24816,N_20290,N_19982);
xnor U24817 (N_24817,N_21279,N_19862);
or U24818 (N_24818,N_21004,N_21736);
nand U24819 (N_24819,N_20496,N_21759);
and U24820 (N_24820,N_18919,N_21133);
nor U24821 (N_24821,N_19696,N_19332);
and U24822 (N_24822,N_19701,N_19506);
xnor U24823 (N_24823,N_20698,N_20590);
and U24824 (N_24824,N_20376,N_20745);
nand U24825 (N_24825,N_21243,N_20386);
nor U24826 (N_24826,N_20982,N_19765);
nand U24827 (N_24827,N_21748,N_19929);
nand U24828 (N_24828,N_20754,N_19446);
xnor U24829 (N_24829,N_19722,N_20199);
nor U24830 (N_24830,N_21642,N_21098);
xor U24831 (N_24831,N_19358,N_21050);
or U24832 (N_24832,N_18836,N_19055);
nor U24833 (N_24833,N_20411,N_19346);
nand U24834 (N_24834,N_21813,N_21275);
or U24835 (N_24835,N_20106,N_20170);
and U24836 (N_24836,N_19591,N_19421);
nor U24837 (N_24837,N_21383,N_21242);
nand U24838 (N_24838,N_20261,N_21652);
or U24839 (N_24839,N_21319,N_19015);
nand U24840 (N_24840,N_20978,N_20622);
nor U24841 (N_24841,N_21546,N_21709);
xor U24842 (N_24842,N_20754,N_21589);
nor U24843 (N_24843,N_19229,N_21148);
and U24844 (N_24844,N_21553,N_21198);
xor U24845 (N_24845,N_20079,N_19492);
nand U24846 (N_24846,N_21622,N_19359);
nand U24847 (N_24847,N_20413,N_21046);
and U24848 (N_24848,N_19944,N_21653);
xor U24849 (N_24849,N_19319,N_18954);
and U24850 (N_24850,N_21009,N_21819);
or U24851 (N_24851,N_19090,N_19307);
or U24852 (N_24852,N_20505,N_20012);
or U24853 (N_24853,N_19803,N_19552);
nor U24854 (N_24854,N_19811,N_20446);
nor U24855 (N_24855,N_19277,N_20997);
or U24856 (N_24856,N_19412,N_21076);
xnor U24857 (N_24857,N_21067,N_19510);
nand U24858 (N_24858,N_20872,N_20686);
nor U24859 (N_24859,N_18771,N_20292);
nand U24860 (N_24860,N_20239,N_21722);
and U24861 (N_24861,N_19621,N_20088);
nor U24862 (N_24862,N_21748,N_20240);
or U24863 (N_24863,N_21074,N_18870);
xnor U24864 (N_24864,N_21656,N_20826);
and U24865 (N_24865,N_20739,N_19064);
and U24866 (N_24866,N_21836,N_19003);
and U24867 (N_24867,N_21302,N_21827);
xnor U24868 (N_24868,N_19536,N_19336);
and U24869 (N_24869,N_21121,N_20708);
nand U24870 (N_24870,N_21089,N_21063);
nand U24871 (N_24871,N_20930,N_19225);
or U24872 (N_24872,N_19793,N_20409);
xor U24873 (N_24873,N_21341,N_20504);
nand U24874 (N_24874,N_19013,N_19903);
and U24875 (N_24875,N_21528,N_19356);
nor U24876 (N_24876,N_19948,N_20483);
nand U24877 (N_24877,N_21561,N_20173);
or U24878 (N_24878,N_20106,N_20479);
or U24879 (N_24879,N_21014,N_19450);
or U24880 (N_24880,N_21463,N_20555);
nand U24881 (N_24881,N_18907,N_19889);
nor U24882 (N_24882,N_20242,N_20564);
and U24883 (N_24883,N_19729,N_21676);
xnor U24884 (N_24884,N_18892,N_20795);
nor U24885 (N_24885,N_19868,N_21485);
or U24886 (N_24886,N_21397,N_20594);
or U24887 (N_24887,N_21727,N_19513);
or U24888 (N_24888,N_20799,N_20054);
xnor U24889 (N_24889,N_19551,N_20014);
nand U24890 (N_24890,N_18992,N_21482);
nand U24891 (N_24891,N_19647,N_21356);
and U24892 (N_24892,N_21711,N_20619);
xnor U24893 (N_24893,N_20799,N_20372);
or U24894 (N_24894,N_19088,N_21787);
xnor U24895 (N_24895,N_18980,N_19743);
nor U24896 (N_24896,N_21065,N_19522);
xor U24897 (N_24897,N_20613,N_19607);
or U24898 (N_24898,N_21845,N_19555);
and U24899 (N_24899,N_21860,N_20979);
and U24900 (N_24900,N_20576,N_21175);
xor U24901 (N_24901,N_21101,N_19855);
or U24902 (N_24902,N_19866,N_20001);
nor U24903 (N_24903,N_20247,N_20526);
and U24904 (N_24904,N_21459,N_20660);
or U24905 (N_24905,N_19152,N_19774);
and U24906 (N_24906,N_20890,N_19706);
nor U24907 (N_24907,N_19002,N_19831);
or U24908 (N_24908,N_21689,N_19052);
nand U24909 (N_24909,N_20636,N_19959);
and U24910 (N_24910,N_21101,N_19602);
or U24911 (N_24911,N_19000,N_21439);
nor U24912 (N_24912,N_19517,N_21418);
nand U24913 (N_24913,N_20219,N_20374);
xor U24914 (N_24914,N_19039,N_19889);
nand U24915 (N_24915,N_19032,N_19289);
and U24916 (N_24916,N_21805,N_18956);
and U24917 (N_24917,N_18901,N_20068);
and U24918 (N_24918,N_19678,N_20055);
or U24919 (N_24919,N_19184,N_19188);
or U24920 (N_24920,N_19497,N_21763);
or U24921 (N_24921,N_20872,N_19422);
and U24922 (N_24922,N_21032,N_19223);
and U24923 (N_24923,N_20479,N_20847);
and U24924 (N_24924,N_19011,N_19079);
and U24925 (N_24925,N_19199,N_20094);
and U24926 (N_24926,N_20364,N_21008);
or U24927 (N_24927,N_18756,N_19790);
nand U24928 (N_24928,N_20343,N_20285);
nand U24929 (N_24929,N_20253,N_20848);
xor U24930 (N_24930,N_19044,N_21839);
nand U24931 (N_24931,N_19365,N_21732);
nand U24932 (N_24932,N_20179,N_20954);
nor U24933 (N_24933,N_20125,N_19236);
nor U24934 (N_24934,N_21254,N_20056);
and U24935 (N_24935,N_20271,N_21636);
or U24936 (N_24936,N_19801,N_21117);
or U24937 (N_24937,N_21549,N_19215);
xor U24938 (N_24938,N_21865,N_21353);
xnor U24939 (N_24939,N_19643,N_19900);
nand U24940 (N_24940,N_20165,N_20225);
nor U24941 (N_24941,N_18813,N_20304);
or U24942 (N_24942,N_19224,N_20975);
or U24943 (N_24943,N_21235,N_19588);
xor U24944 (N_24944,N_18780,N_20610);
or U24945 (N_24945,N_20990,N_19648);
nand U24946 (N_24946,N_20917,N_21791);
nor U24947 (N_24947,N_19026,N_18814);
nand U24948 (N_24948,N_20484,N_21785);
and U24949 (N_24949,N_19100,N_21692);
or U24950 (N_24950,N_19265,N_21291);
nor U24951 (N_24951,N_21671,N_20708);
or U24952 (N_24952,N_20561,N_19199);
and U24953 (N_24953,N_20078,N_18750);
nand U24954 (N_24954,N_19121,N_21644);
xor U24955 (N_24955,N_20693,N_19687);
and U24956 (N_24956,N_21352,N_20536);
nand U24957 (N_24957,N_21655,N_20334);
or U24958 (N_24958,N_21224,N_20115);
and U24959 (N_24959,N_18904,N_19379);
nand U24960 (N_24960,N_20036,N_19308);
and U24961 (N_24961,N_19847,N_20322);
nand U24962 (N_24962,N_21172,N_20479);
or U24963 (N_24963,N_19478,N_20320);
xnor U24964 (N_24964,N_21458,N_19906);
and U24965 (N_24965,N_19276,N_19598);
or U24966 (N_24966,N_19488,N_20968);
nor U24967 (N_24967,N_20087,N_20713);
nand U24968 (N_24968,N_19642,N_21851);
nand U24969 (N_24969,N_18954,N_19097);
nor U24970 (N_24970,N_21220,N_21019);
nand U24971 (N_24971,N_19190,N_18959);
or U24972 (N_24972,N_20805,N_21385);
xnor U24973 (N_24973,N_19534,N_19023);
xor U24974 (N_24974,N_18838,N_21201);
or U24975 (N_24975,N_19774,N_21831);
xor U24976 (N_24976,N_21328,N_20982);
xnor U24977 (N_24977,N_19155,N_20193);
or U24978 (N_24978,N_20441,N_20278);
nand U24979 (N_24979,N_20059,N_21519);
nand U24980 (N_24980,N_19935,N_18838);
nor U24981 (N_24981,N_19831,N_20039);
or U24982 (N_24982,N_19468,N_20741);
nand U24983 (N_24983,N_20053,N_19453);
or U24984 (N_24984,N_20891,N_20919);
nor U24985 (N_24985,N_21097,N_19310);
and U24986 (N_24986,N_19705,N_21051);
xnor U24987 (N_24987,N_21759,N_20914);
nand U24988 (N_24988,N_21455,N_19786);
nor U24989 (N_24989,N_20576,N_20025);
nand U24990 (N_24990,N_21068,N_20374);
nor U24991 (N_24991,N_20071,N_19580);
nor U24992 (N_24992,N_21373,N_19755);
or U24993 (N_24993,N_20728,N_19802);
nand U24994 (N_24994,N_21085,N_21283);
nor U24995 (N_24995,N_19521,N_20755);
and U24996 (N_24996,N_20170,N_21404);
nand U24997 (N_24997,N_18988,N_19646);
nand U24998 (N_24998,N_19008,N_18951);
nor U24999 (N_24999,N_19535,N_19659);
and UO_0 (O_0,N_22278,N_22838);
nor UO_1 (O_1,N_22489,N_22486);
nand UO_2 (O_2,N_22629,N_21891);
nor UO_3 (O_3,N_21974,N_22848);
nor UO_4 (O_4,N_21882,N_22410);
nand UO_5 (O_5,N_23942,N_21939);
nor UO_6 (O_6,N_22693,N_24476);
and UO_7 (O_7,N_24088,N_23636);
xnor UO_8 (O_8,N_23356,N_23780);
or UO_9 (O_9,N_24444,N_23847);
and UO_10 (O_10,N_23988,N_22977);
and UO_11 (O_11,N_23564,N_24780);
nand UO_12 (O_12,N_23435,N_22034);
nand UO_13 (O_13,N_23080,N_23016);
nor UO_14 (O_14,N_24796,N_23285);
xor UO_15 (O_15,N_23656,N_24855);
and UO_16 (O_16,N_24682,N_24896);
nor UO_17 (O_17,N_24218,N_23253);
and UO_18 (O_18,N_23110,N_24948);
nand UO_19 (O_19,N_24635,N_24652);
nand UO_20 (O_20,N_24078,N_22895);
and UO_21 (O_21,N_24670,N_24607);
nor UO_22 (O_22,N_23925,N_22585);
and UO_23 (O_23,N_22301,N_24057);
nand UO_24 (O_24,N_24334,N_22095);
nand UO_25 (O_25,N_24025,N_22267);
xor UO_26 (O_26,N_23149,N_23087);
nor UO_27 (O_27,N_24574,N_22658);
and UO_28 (O_28,N_24632,N_24806);
xnor UO_29 (O_29,N_23146,N_23451);
xnor UO_30 (O_30,N_22208,N_22437);
or UO_31 (O_31,N_24602,N_22344);
nand UO_32 (O_32,N_23241,N_24917);
nor UO_33 (O_33,N_22409,N_23368);
nor UO_34 (O_34,N_22317,N_22780);
nor UO_35 (O_35,N_24363,N_24936);
nand UO_36 (O_36,N_24684,N_24991);
nand UO_37 (O_37,N_23294,N_22953);
xor UO_38 (O_38,N_21893,N_22180);
nor UO_39 (O_39,N_21972,N_22498);
nor UO_40 (O_40,N_22916,N_24337);
or UO_41 (O_41,N_21926,N_23585);
xnor UO_42 (O_42,N_23433,N_22287);
nand UO_43 (O_43,N_22984,N_22198);
xnor UO_44 (O_44,N_21951,N_23125);
nand UO_45 (O_45,N_23626,N_23319);
nor UO_46 (O_46,N_24825,N_22762);
and UO_47 (O_47,N_22169,N_24410);
or UO_48 (O_48,N_24767,N_22005);
xor UO_49 (O_49,N_22500,N_23429);
and UO_50 (O_50,N_24145,N_24085);
xor UO_51 (O_51,N_24086,N_23842);
and UO_52 (O_52,N_21977,N_23587);
or UO_53 (O_53,N_23015,N_22215);
or UO_54 (O_54,N_24318,N_24878);
nand UO_55 (O_55,N_24886,N_23601);
nand UO_56 (O_56,N_24719,N_23295);
nor UO_57 (O_57,N_24597,N_22909);
or UO_58 (O_58,N_22030,N_24250);
xnor UO_59 (O_59,N_22761,N_24155);
nand UO_60 (O_60,N_24469,N_23409);
and UO_61 (O_61,N_24683,N_24952);
or UO_62 (O_62,N_23474,N_24842);
or UO_63 (O_63,N_24675,N_23277);
nor UO_64 (O_64,N_23662,N_23164);
nor UO_65 (O_65,N_24508,N_22995);
or UO_66 (O_66,N_22485,N_24465);
nand UO_67 (O_67,N_24553,N_24560);
and UO_68 (O_68,N_24576,N_23224);
nand UO_69 (O_69,N_22682,N_21879);
nand UO_70 (O_70,N_22702,N_22860);
xnor UO_71 (O_71,N_24461,N_24768);
xnor UO_72 (O_72,N_23683,N_23766);
and UO_73 (O_73,N_24150,N_24380);
nor UO_74 (O_74,N_22948,N_22634);
or UO_75 (O_75,N_23620,N_22816);
or UO_76 (O_76,N_23380,N_24620);
and UO_77 (O_77,N_24133,N_22767);
xor UO_78 (O_78,N_22681,N_24152);
nand UO_79 (O_79,N_23234,N_23185);
or UO_80 (O_80,N_22022,N_23046);
or UO_81 (O_81,N_22806,N_22567);
xnor UO_82 (O_82,N_24450,N_21906);
nand UO_83 (O_83,N_24887,N_24548);
xor UO_84 (O_84,N_23562,N_22796);
or UO_85 (O_85,N_23961,N_23273);
nor UO_86 (O_86,N_24499,N_22297);
xor UO_87 (O_87,N_22366,N_23283);
or UO_88 (O_88,N_22367,N_22216);
nand UO_89 (O_89,N_23109,N_23346);
nand UO_90 (O_90,N_23931,N_22440);
and UO_91 (O_91,N_24624,N_23750);
or UO_92 (O_92,N_22908,N_22457);
xor UO_93 (O_93,N_23117,N_23054);
and UO_94 (O_94,N_24930,N_22803);
xor UO_95 (O_95,N_23619,N_23765);
xor UO_96 (O_96,N_24726,N_22122);
nor UO_97 (O_97,N_22662,N_23084);
nor UO_98 (O_98,N_21892,N_23603);
nand UO_99 (O_99,N_24464,N_24906);
or UO_100 (O_100,N_22353,N_24281);
nand UO_101 (O_101,N_24591,N_24154);
or UO_102 (O_102,N_22362,N_23193);
nand UO_103 (O_103,N_23240,N_24966);
or UO_104 (O_104,N_22322,N_21995);
nor UO_105 (O_105,N_24783,N_23332);
or UO_106 (O_106,N_22894,N_22219);
nor UO_107 (O_107,N_24378,N_24484);
nand UO_108 (O_108,N_24904,N_23903);
nand UO_109 (O_109,N_24891,N_24716);
xnor UO_110 (O_110,N_21927,N_23539);
and UO_111 (O_111,N_23375,N_24434);
or UO_112 (O_112,N_22432,N_24206);
xor UO_113 (O_113,N_24999,N_24105);
xor UO_114 (O_114,N_22959,N_24995);
and UO_115 (O_115,N_22117,N_24800);
or UO_116 (O_116,N_23630,N_24278);
xnor UO_117 (O_117,N_24126,N_22231);
nand UO_118 (O_118,N_21985,N_24113);
and UO_119 (O_119,N_22102,N_23712);
nand UO_120 (O_120,N_22017,N_23915);
xnor UO_121 (O_121,N_23764,N_22480);
xor UO_122 (O_122,N_24753,N_24093);
nor UO_123 (O_123,N_23650,N_22471);
nor UO_124 (O_124,N_24423,N_22944);
xor UO_125 (O_125,N_22191,N_23227);
nor UO_126 (O_126,N_24920,N_23422);
or UO_127 (O_127,N_24397,N_22318);
nand UO_128 (O_128,N_23821,N_22652);
xor UO_129 (O_129,N_22165,N_23716);
xnor UO_130 (O_130,N_24103,N_23657);
nor UO_131 (O_131,N_23349,N_22919);
and UO_132 (O_132,N_23640,N_24622);
and UO_133 (O_133,N_24164,N_24890);
or UO_134 (O_134,N_22637,N_22164);
or UO_135 (O_135,N_23904,N_24998);
or UO_136 (O_136,N_23641,N_23778);
and UO_137 (O_137,N_24854,N_23031);
or UO_138 (O_138,N_22354,N_24513);
xor UO_139 (O_139,N_24926,N_23525);
and UO_140 (O_140,N_22113,N_23112);
or UO_141 (O_141,N_24177,N_24095);
nor UO_142 (O_142,N_24340,N_23089);
nand UO_143 (O_143,N_22282,N_24431);
or UO_144 (O_144,N_24416,N_22782);
xnor UO_145 (O_145,N_24784,N_23906);
nand UO_146 (O_146,N_24128,N_23408);
nor UO_147 (O_147,N_22091,N_23577);
or UO_148 (O_148,N_23222,N_22669);
nand UO_149 (O_149,N_23327,N_24394);
and UO_150 (O_150,N_23049,N_23604);
nand UO_151 (O_151,N_24244,N_23479);
nor UO_152 (O_152,N_24102,N_23397);
xor UO_153 (O_153,N_24943,N_22859);
and UO_154 (O_154,N_23258,N_22512);
xor UO_155 (O_155,N_22904,N_23195);
or UO_156 (O_156,N_22651,N_23898);
or UO_157 (O_157,N_24918,N_24437);
nand UO_158 (O_158,N_24667,N_24251);
xor UO_159 (O_159,N_23901,N_22356);
nor UO_160 (O_160,N_24644,N_21901);
nand UO_161 (O_161,N_22999,N_24766);
nor UO_162 (O_162,N_24846,N_22826);
or UO_163 (O_163,N_23524,N_24373);
or UO_164 (O_164,N_22997,N_22068);
nand UO_165 (O_165,N_23043,N_22056);
xor UO_166 (O_166,N_22177,N_24472);
nand UO_167 (O_167,N_24064,N_22127);
nand UO_168 (O_168,N_24613,N_23105);
xor UO_169 (O_169,N_23774,N_23320);
nor UO_170 (O_170,N_22416,N_22808);
xor UO_171 (O_171,N_21905,N_24941);
xor UO_172 (O_172,N_22163,N_22308);
or UO_173 (O_173,N_22578,N_24122);
or UO_174 (O_174,N_22740,N_24140);
and UO_175 (O_175,N_23999,N_23364);
xnor UO_176 (O_176,N_23698,N_22115);
nor UO_177 (O_177,N_24819,N_24467);
nor UO_178 (O_178,N_24295,N_24045);
nand UO_179 (O_179,N_23651,N_22636);
xor UO_180 (O_180,N_23315,N_24353);
nand UO_181 (O_181,N_22481,N_22288);
nand UO_182 (O_182,N_23873,N_23994);
nand UO_183 (O_183,N_22212,N_23790);
nand UO_184 (O_184,N_23384,N_24880);
nand UO_185 (O_185,N_23247,N_22070);
or UO_186 (O_186,N_23310,N_24672);
or UO_187 (O_187,N_24138,N_24238);
nor UO_188 (O_188,N_23827,N_23861);
and UO_189 (O_189,N_21922,N_22910);
nor UO_190 (O_190,N_21877,N_22565);
or UO_191 (O_191,N_22229,N_22533);
nor UO_192 (O_192,N_24744,N_23184);
nor UO_193 (O_193,N_22284,N_24587);
and UO_194 (O_194,N_23893,N_22986);
xor UO_195 (O_195,N_23501,N_23884);
nand UO_196 (O_196,N_22444,N_23967);
and UO_197 (O_197,N_24175,N_21971);
and UO_198 (O_198,N_23625,N_24023);
and UO_199 (O_199,N_24374,N_24640);
nand UO_200 (O_200,N_22139,N_22739);
nor UO_201 (O_201,N_24984,N_22172);
and UO_202 (O_202,N_24961,N_22843);
xnor UO_203 (O_203,N_22188,N_22744);
nand UO_204 (O_204,N_24003,N_24993);
nor UO_205 (O_205,N_23550,N_22508);
xnor UO_206 (O_206,N_23246,N_24745);
nor UO_207 (O_207,N_21986,N_22869);
and UO_208 (O_208,N_22442,N_24965);
nor UO_209 (O_209,N_23148,N_24165);
nor UO_210 (O_210,N_21888,N_24741);
nand UO_211 (O_211,N_22086,N_22880);
nor UO_212 (O_212,N_22729,N_22793);
or UO_213 (O_213,N_23991,N_23341);
nand UO_214 (O_214,N_21887,N_24322);
xnor UO_215 (O_215,N_24723,N_23088);
nor UO_216 (O_216,N_23161,N_24132);
xor UO_217 (O_217,N_23508,N_22016);
and UO_218 (O_218,N_24047,N_21928);
xnor UO_219 (O_219,N_24990,N_24844);
and UO_220 (O_220,N_24951,N_22732);
nand UO_221 (O_221,N_23167,N_23731);
and UO_222 (O_222,N_24972,N_23589);
nor UO_223 (O_223,N_24069,N_24939);
xor UO_224 (O_224,N_22764,N_23573);
xnor UO_225 (O_225,N_21909,N_23201);
or UO_226 (O_226,N_23869,N_22296);
nand UO_227 (O_227,N_24571,N_24293);
or UO_228 (O_228,N_24687,N_22801);
nor UO_229 (O_229,N_24158,N_23093);
or UO_230 (O_230,N_24751,N_24409);
and UO_231 (O_231,N_22445,N_23358);
xnor UO_232 (O_232,N_24160,N_22590);
and UO_233 (O_233,N_22612,N_24792);
xor UO_234 (O_234,N_23183,N_24289);
nand UO_235 (O_235,N_24714,N_22323);
and UO_236 (O_236,N_22026,N_24178);
nor UO_237 (O_237,N_23993,N_23369);
xnor UO_238 (O_238,N_22772,N_24121);
xnor UO_239 (O_239,N_23092,N_23949);
xor UO_240 (O_240,N_23916,N_23137);
nand UO_241 (O_241,N_22196,N_23530);
or UO_242 (O_242,N_21996,N_22831);
nor UO_243 (O_243,N_23387,N_23472);
nor UO_244 (O_244,N_22062,N_23521);
xor UO_245 (O_245,N_22077,N_23517);
xor UO_246 (O_246,N_24830,N_24094);
xor UO_247 (O_247,N_23954,N_23527);
or UO_248 (O_248,N_24899,N_24705);
and UO_249 (O_249,N_23237,N_24949);
or UO_250 (O_250,N_23071,N_24486);
nand UO_251 (O_251,N_22725,N_24211);
or UO_252 (O_252,N_22623,N_23519);
and UO_253 (O_253,N_23749,N_23446);
or UO_254 (O_254,N_24971,N_24435);
nor UO_255 (O_255,N_22294,N_23814);
or UO_256 (O_256,N_21914,N_22265);
nand UO_257 (O_257,N_22233,N_24430);
and UO_258 (O_258,N_22561,N_22888);
or UO_259 (O_259,N_24457,N_24605);
or UO_260 (O_260,N_24722,N_24071);
nand UO_261 (O_261,N_23639,N_24843);
or UO_262 (O_262,N_24312,N_23826);
nor UO_263 (O_263,N_22506,N_22186);
xnor UO_264 (O_264,N_22600,N_24427);
nor UO_265 (O_265,N_22584,N_22811);
xor UO_266 (O_266,N_24139,N_23303);
nor UO_267 (O_267,N_22815,N_22560);
and UO_268 (O_268,N_24053,N_23432);
nor UO_269 (O_269,N_22528,N_22543);
nand UO_270 (O_270,N_23726,N_22784);
or UO_271 (O_271,N_21923,N_23823);
nand UO_272 (O_272,N_24273,N_24310);
or UO_273 (O_273,N_22333,N_23282);
xnor UO_274 (O_274,N_23718,N_23645);
or UO_275 (O_275,N_24717,N_22941);
or UO_276 (O_276,N_23238,N_24223);
nand UO_277 (O_277,N_24847,N_22329);
xnor UO_278 (O_278,N_22853,N_24029);
nand UO_279 (O_279,N_23744,N_23487);
nand UO_280 (O_280,N_23052,N_24169);
and UO_281 (O_281,N_22920,N_23617);
nor UO_282 (O_282,N_22008,N_22421);
and UO_283 (O_283,N_23175,N_23436);
nor UO_284 (O_284,N_23325,N_22663);
nand UO_285 (O_285,N_22738,N_24627);
xnor UO_286 (O_286,N_23628,N_24616);
nand UO_287 (O_287,N_24889,N_24983);
nor UO_288 (O_288,N_21981,N_23202);
or UO_289 (O_289,N_22391,N_21998);
xor UO_290 (O_290,N_22555,N_23615);
or UO_291 (O_291,N_24260,N_22829);
and UO_292 (O_292,N_22569,N_24383);
nand UO_293 (O_293,N_24543,N_23733);
or UO_294 (O_294,N_21962,N_21886);
xor UO_295 (O_295,N_23666,N_23066);
xor UO_296 (O_296,N_24505,N_23249);
nor UO_297 (O_297,N_23439,N_24236);
and UO_298 (O_298,N_23413,N_24243);
or UO_299 (O_299,N_22502,N_23857);
and UO_300 (O_300,N_23810,N_24204);
nor UO_301 (O_301,N_23464,N_24647);
or UO_302 (O_302,N_24219,N_23153);
xor UO_303 (O_303,N_23162,N_23523);
nor UO_304 (O_304,N_24452,N_22210);
and UO_305 (O_305,N_23978,N_23165);
xnor UO_306 (O_306,N_21921,N_22351);
and UO_307 (O_307,N_24987,N_22695);
nand UO_308 (O_308,N_24030,N_24041);
nor UO_309 (O_309,N_24845,N_22598);
or UO_310 (O_310,N_23189,N_24076);
and UO_311 (O_311,N_24573,N_22802);
and UO_312 (O_312,N_24657,N_23278);
xnor UO_313 (O_313,N_23710,N_23050);
xnor UO_314 (O_314,N_24341,N_22388);
nand UO_315 (O_315,N_22896,N_24737);
xnor UO_316 (O_316,N_21918,N_22657);
nand UO_317 (O_317,N_22987,N_24633);
xnor UO_318 (O_318,N_22203,N_22148);
or UO_319 (O_319,N_22339,N_24284);
nor UO_320 (O_320,N_22577,N_24167);
and UO_321 (O_321,N_24658,N_23748);
nor UO_322 (O_322,N_24557,N_22734);
and UO_323 (O_323,N_24817,N_22958);
or UO_324 (O_324,N_22721,N_22493);
or UO_325 (O_325,N_23041,N_24720);
nor UO_326 (O_326,N_22307,N_22377);
nor UO_327 (O_327,N_24733,N_23350);
nand UO_328 (O_328,N_23219,N_21938);
xor UO_329 (O_329,N_23541,N_22065);
nor UO_330 (O_330,N_21942,N_24955);
and UO_331 (O_331,N_23099,N_23402);
nor UO_332 (O_332,N_23196,N_23377);
nor UO_333 (O_333,N_21973,N_24407);
nor UO_334 (O_334,N_23854,N_22406);
nor UO_335 (O_335,N_22546,N_21884);
xnor UO_336 (O_336,N_24022,N_21944);
nor UO_337 (O_337,N_22456,N_23329);
and UO_338 (O_338,N_22060,N_24162);
nor UO_339 (O_339,N_22756,N_22821);
nand UO_340 (O_340,N_24364,N_22428);
nand UO_341 (O_341,N_24763,N_23998);
or UO_342 (O_342,N_22972,N_23878);
xnor UO_343 (O_343,N_23902,N_24021);
or UO_344 (O_344,N_22272,N_22358);
and UO_345 (O_345,N_22971,N_24600);
nor UO_346 (O_346,N_22970,N_24699);
or UO_347 (O_347,N_22677,N_22211);
or UO_348 (O_348,N_23629,N_24782);
xnor UO_349 (O_349,N_22683,N_22407);
nand UO_350 (O_350,N_22545,N_23691);
xor UO_351 (O_351,N_22217,N_24487);
xor UO_352 (O_352,N_24738,N_21982);
and UO_353 (O_353,N_22069,N_22010);
xor UO_354 (O_354,N_22884,N_24732);
or UO_355 (O_355,N_21975,N_23836);
or UO_356 (O_356,N_23646,N_23305);
nor UO_357 (O_357,N_21955,N_22025);
and UO_358 (O_358,N_22104,N_24436);
nand UO_359 (O_359,N_23082,N_24498);
nand UO_360 (O_360,N_23073,N_22690);
nor UO_361 (O_361,N_22059,N_23095);
and UO_362 (O_362,N_23142,N_23830);
nor UO_363 (O_363,N_24901,N_22643);
xnor UO_364 (O_364,N_22464,N_22704);
nand UO_365 (O_365,N_22051,N_23172);
xnor UO_366 (O_366,N_24893,N_22072);
and UO_367 (O_367,N_23879,N_24382);
xor UO_368 (O_368,N_23383,N_23828);
xor UO_369 (O_369,N_24665,N_22722);
and UO_370 (O_370,N_23627,N_24166);
and UO_371 (O_371,N_22544,N_22038);
nor UO_372 (O_372,N_22542,N_24215);
and UO_373 (O_373,N_23024,N_23753);
nand UO_374 (O_374,N_22589,N_23692);
nor UO_375 (O_375,N_23876,N_22522);
and UO_376 (O_376,N_23445,N_22580);
or UO_377 (O_377,N_23534,N_23379);
nand UO_378 (O_378,N_23460,N_22269);
nand UO_379 (O_379,N_23463,N_23211);
and UO_380 (O_380,N_24570,N_22789);
nand UO_381 (O_381,N_22047,N_22559);
nand UO_382 (O_382,N_22338,N_23160);
and UO_383 (O_383,N_24376,N_23055);
xnor UO_384 (O_384,N_23311,N_23602);
xor UO_385 (O_385,N_22201,N_23104);
and UO_386 (O_386,N_22586,N_22627);
or UO_387 (O_387,N_23980,N_24718);
xor UO_388 (O_388,N_21994,N_23069);
nor UO_389 (O_389,N_22509,N_22023);
or UO_390 (O_390,N_23326,N_24187);
xor UO_391 (O_391,N_23803,N_22531);
or UO_392 (O_392,N_23226,N_22001);
nor UO_393 (O_393,N_23702,N_22730);
xnor UO_394 (O_394,N_23840,N_23169);
and UO_395 (O_395,N_22688,N_22737);
and UO_396 (O_396,N_22587,N_24894);
and UO_397 (O_397,N_24969,N_24533);
nand UO_398 (O_398,N_22315,N_24836);
xor UO_399 (O_399,N_21902,N_22342);
and UO_400 (O_400,N_24693,N_24496);
xor UO_401 (O_401,N_23886,N_24460);
xor UO_402 (O_402,N_23735,N_24905);
nor UO_403 (O_403,N_22374,N_22571);
nand UO_404 (O_404,N_22973,N_23461);
or UO_405 (O_405,N_22446,N_23313);
xnor UO_406 (O_406,N_22520,N_24707);
or UO_407 (O_407,N_24402,N_23509);
or UO_408 (O_408,N_24606,N_21987);
or UO_409 (O_409,N_23526,N_24096);
xnor UO_410 (O_410,N_22967,N_24144);
and UO_411 (O_411,N_24892,N_24040);
nand UO_412 (O_412,N_24090,N_23133);
xor UO_413 (O_413,N_24660,N_21947);
and UO_414 (O_414,N_23754,N_22628);
and UO_415 (O_415,N_23819,N_23996);
xnor UO_416 (O_416,N_23267,N_22431);
xor UO_417 (O_417,N_24556,N_24365);
xnor UO_418 (O_418,N_23121,N_23768);
nor UO_419 (O_419,N_24522,N_22252);
xor UO_420 (O_420,N_22731,N_22805);
or UO_421 (O_421,N_23897,N_24933);
and UO_422 (O_422,N_23373,N_23357);
or UO_423 (O_423,N_23862,N_23470);
nand UO_424 (O_424,N_23200,N_24946);
nor UO_425 (O_425,N_22257,N_22451);
and UO_426 (O_426,N_24208,N_24968);
nand UO_427 (O_427,N_23887,N_23838);
or UO_428 (O_428,N_23136,N_24115);
nor UO_429 (O_429,N_21945,N_24695);
nand UO_430 (O_430,N_21959,N_23740);
or UO_431 (O_431,N_23450,N_24216);
xor UO_432 (O_432,N_24801,N_24455);
xor UO_433 (O_433,N_24769,N_23660);
xnor UO_434 (O_434,N_24676,N_24109);
nand UO_435 (O_435,N_22511,N_24601);
and UO_436 (O_436,N_24540,N_23404);
xnor UO_437 (O_437,N_23317,N_24519);
nor UO_438 (O_438,N_22146,N_22867);
and UO_439 (O_439,N_23122,N_24879);
or UO_440 (O_440,N_24253,N_24392);
xor UO_441 (O_441,N_23382,N_22616);
or UO_442 (O_442,N_24756,N_22084);
and UO_443 (O_443,N_23538,N_24161);
nor UO_444 (O_444,N_22911,N_22205);
and UO_445 (O_445,N_22675,N_22131);
nor UO_446 (O_446,N_22844,N_22689);
nand UO_447 (O_447,N_23720,N_22534);
xnor UO_448 (O_448,N_22147,N_23248);
nand UO_449 (O_449,N_24014,N_23159);
nand UO_450 (O_450,N_23107,N_23351);
xor UO_451 (O_451,N_23483,N_22243);
and UO_452 (O_452,N_23773,N_23223);
or UO_453 (O_453,N_23934,N_24781);
and UO_454 (O_454,N_24485,N_22705);
and UO_455 (O_455,N_23658,N_24012);
nor UO_456 (O_456,N_23667,N_24862);
or UO_457 (O_457,N_23336,N_22951);
or UO_458 (O_458,N_24291,N_22668);
or UO_459 (O_459,N_24181,N_22766);
xnor UO_460 (O_460,N_23536,N_23844);
and UO_461 (O_461,N_24403,N_21949);
xnor UO_462 (O_462,N_22174,N_22370);
or UO_463 (O_463,N_22699,N_24307);
and UO_464 (O_464,N_22454,N_24013);
or UO_465 (O_465,N_22273,N_22939);
nand UO_466 (O_466,N_23608,N_24956);
or UO_467 (O_467,N_24550,N_24112);
xor UO_468 (O_468,N_24863,N_24202);
nor UO_469 (O_469,N_24921,N_23434);
nand UO_470 (O_470,N_23775,N_24747);
xor UO_471 (O_471,N_22040,N_24209);
or UO_472 (O_472,N_21984,N_23010);
nor UO_473 (O_473,N_24681,N_23900);
or UO_474 (O_474,N_23290,N_22264);
nand UO_475 (O_475,N_23118,N_24580);
and UO_476 (O_476,N_24354,N_23500);
xnor UO_477 (O_477,N_22564,N_23938);
xnor UO_478 (O_478,N_23616,N_24925);
nor UO_479 (O_479,N_24074,N_24470);
or UO_480 (O_480,N_23548,N_23067);
or UO_481 (O_481,N_24123,N_22866);
and UO_482 (O_482,N_22513,N_23704);
nand UO_483 (O_483,N_23076,N_23263);
nor UO_484 (O_484,N_24339,N_24758);
and UO_485 (O_485,N_24420,N_22864);
xnor UO_486 (O_486,N_24765,N_24006);
or UO_487 (O_487,N_22014,N_24297);
nand UO_488 (O_488,N_23552,N_22039);
and UO_489 (O_489,N_22413,N_22966);
xnor UO_490 (O_490,N_24549,N_24639);
and UO_491 (O_491,N_22684,N_24860);
nand UO_492 (O_492,N_22343,N_22305);
nor UO_493 (O_493,N_22798,N_24422);
nor UO_494 (O_494,N_23695,N_24044);
or UO_495 (O_495,N_23496,N_23174);
nor UO_496 (O_496,N_22304,N_22400);
nand UO_497 (O_497,N_22820,N_22223);
or UO_498 (O_498,N_23051,N_22582);
nand UO_499 (O_499,N_23466,N_22327);
nand UO_500 (O_500,N_24612,N_22107);
xnor UO_501 (O_501,N_22303,N_24775);
xnor UO_502 (O_502,N_24835,N_24327);
xor UO_503 (O_503,N_22783,N_23399);
nor UO_504 (O_504,N_23157,N_24494);
xnor UO_505 (O_505,N_23808,N_23837);
and UO_506 (O_506,N_24367,N_22314);
or UO_507 (O_507,N_23114,N_22061);
xnor UO_508 (O_508,N_23742,N_22097);
xor UO_509 (O_509,N_23575,N_23255);
and UO_510 (O_510,N_23782,N_22020);
nor UO_511 (O_511,N_22621,N_22785);
nand UO_512 (O_512,N_24653,N_22466);
and UO_513 (O_513,N_23037,N_22779);
or UO_514 (O_514,N_22408,N_22249);
nand UO_515 (O_515,N_24406,N_21916);
or UO_516 (O_516,N_22752,N_22963);
or UO_517 (O_517,N_24696,N_22755);
nand UO_518 (O_518,N_23870,N_22340);
and UO_519 (O_519,N_24527,N_24134);
nor UO_520 (O_520,N_24170,N_22603);
or UO_521 (O_521,N_22402,N_24881);
or UO_522 (O_522,N_23727,N_22570);
or UO_523 (O_523,N_23334,N_24668);
nor UO_524 (O_524,N_22483,N_23940);
or UO_525 (O_525,N_23039,N_23476);
xnor UO_526 (O_526,N_23846,N_23685);
or UO_527 (O_527,N_24292,N_22591);
and UO_528 (O_528,N_23001,N_23992);
xor UO_529 (O_529,N_22822,N_23251);
xor UO_530 (O_530,N_22929,N_24350);
or UO_531 (O_531,N_22746,N_23062);
or UO_532 (O_532,N_24604,N_24249);
and UO_533 (O_533,N_23987,N_23406);
nand UO_534 (O_534,N_21956,N_24666);
nor UO_535 (O_535,N_23210,N_23624);
or UO_536 (O_536,N_23554,N_24362);
xor UO_537 (O_537,N_22708,N_24812);
nand UO_538 (O_538,N_23719,N_24791);
and UO_539 (O_539,N_24288,N_22736);
or UO_540 (O_540,N_23594,N_21964);
nor UO_541 (O_541,N_23511,N_22554);
nor UO_542 (O_542,N_23514,N_21915);
or UO_543 (O_543,N_23986,N_23187);
and UO_544 (O_544,N_22271,N_24481);
nand UO_545 (O_545,N_23056,N_23694);
nand UO_546 (O_546,N_24272,N_23877);
nand UO_547 (O_547,N_24685,N_22042);
nor UO_548 (O_548,N_22774,N_21885);
xor UO_549 (O_549,N_22300,N_24729);
nand UO_550 (O_550,N_24584,N_22742);
or UO_551 (O_551,N_23990,N_23739);
and UO_552 (O_552,N_23231,N_21968);
nand UO_553 (O_553,N_22548,N_24964);
nand UO_554 (O_554,N_23324,N_23289);
and UO_555 (O_555,N_24978,N_23299);
and UO_556 (O_556,N_22463,N_23111);
nor UO_557 (O_557,N_24412,N_24552);
nand UO_558 (O_558,N_23057,N_22108);
nand UO_559 (O_559,N_21935,N_22239);
xnor UO_560 (O_560,N_23535,N_22477);
and UO_561 (O_561,N_24989,N_24563);
xor UO_562 (O_562,N_23264,N_24443);
nor UO_563 (O_563,N_22202,N_22936);
or UO_564 (O_564,N_22726,N_23690);
or UO_565 (O_565,N_22962,N_22983);
and UO_566 (O_566,N_22857,N_24721);
nor UO_567 (O_567,N_23102,N_22041);
nand UO_568 (O_568,N_22897,N_22817);
nand UO_569 (O_569,N_23457,N_22192);
nor UO_570 (O_570,N_22676,N_24869);
xor UO_571 (O_571,N_22747,N_23917);
nand UO_572 (O_572,N_22281,N_24054);
or UO_573 (O_573,N_22274,N_23592);
nor UO_574 (O_574,N_24748,N_23883);
or UO_575 (O_575,N_24042,N_23342);
xor UO_576 (O_576,N_23804,N_22033);
and UO_577 (O_577,N_24355,N_23937);
nor UO_578 (O_578,N_22289,N_24063);
nand UO_579 (O_579,N_22771,N_24149);
nor UO_580 (O_580,N_23681,N_24578);
nor UO_581 (O_581,N_24306,N_23572);
nor UO_582 (O_582,N_24478,N_22873);
nor UO_583 (O_583,N_23190,N_24913);
xnor UO_584 (O_584,N_24254,N_23599);
xnor UO_585 (O_585,N_22968,N_24032);
nor UO_586 (O_586,N_22248,N_22847);
xnor UO_587 (O_587,N_24561,N_22449);
xnor UO_588 (O_588,N_24075,N_24277);
nand UO_589 (O_589,N_23437,N_23287);
or UO_590 (O_590,N_22532,N_24179);
and UO_591 (O_591,N_23722,N_24509);
nor UO_592 (O_592,N_21934,N_22240);
xnor UO_593 (O_593,N_23975,N_22640);
or UO_594 (O_594,N_24912,N_23068);
xor UO_595 (O_595,N_24997,N_22604);
nor UO_596 (O_596,N_22758,N_24865);
nor UO_597 (O_597,N_21896,N_24520);
nand UO_598 (O_598,N_24368,N_23791);
and UO_599 (O_599,N_22101,N_22638);
nand UO_600 (O_600,N_23096,N_23281);
nor UO_601 (O_601,N_24586,N_24671);
and UO_602 (O_602,N_22320,N_23308);
nand UO_603 (O_603,N_22063,N_24495);
xnor UO_604 (O_604,N_23779,N_23777);
nand UO_605 (O_605,N_22098,N_22552);
or UO_606 (O_606,N_22331,N_22635);
or UO_607 (O_607,N_23168,N_22980);
nor UO_608 (O_608,N_22791,N_24529);
xor UO_609 (O_609,N_23895,N_22714);
and UO_610 (O_610,N_24332,N_24771);
or UO_611 (O_611,N_23256,N_24649);
nor UO_612 (O_612,N_23272,N_22781);
xnor UO_613 (O_613,N_22387,N_24197);
nand UO_614 (O_614,N_24104,N_22423);
nand UO_615 (O_615,N_22516,N_22872);
xnor UO_616 (O_616,N_23420,N_22182);
nand UO_617 (O_617,N_23428,N_23239);
nand UO_618 (O_618,N_23932,N_22112);
xor UO_619 (O_619,N_22458,N_24824);
and UO_620 (O_620,N_23497,N_23858);
or UO_621 (O_621,N_22365,N_22363);
and UO_622 (O_622,N_23053,N_23458);
xor UO_623 (O_623,N_24523,N_23386);
and UO_624 (O_624,N_24559,N_24621);
or UO_625 (O_625,N_24379,N_23401);
nor UO_626 (O_626,N_22381,N_24996);
nor UO_627 (O_627,N_24531,N_23952);
xor UO_628 (O_628,N_24538,N_22144);
xor UO_629 (O_629,N_22797,N_24451);
and UO_630 (O_630,N_22484,N_24518);
nor UO_631 (O_631,N_22247,N_22081);
nor UO_632 (O_632,N_22769,N_23298);
nor UO_633 (O_633,N_23331,N_22660);
and UO_634 (O_634,N_21908,N_23250);
nand UO_635 (O_635,N_23423,N_23444);
and UO_636 (O_636,N_24081,N_22242);
nand UO_637 (O_637,N_22361,N_23378);
nand UO_638 (O_638,N_23529,N_24787);
or UO_639 (O_639,N_24942,N_23418);
and UO_640 (O_640,N_21976,N_24240);
and UO_641 (O_641,N_23686,N_23147);
nor UO_642 (O_642,N_22846,N_22106);
nand UO_643 (O_643,N_24608,N_23367);
nor UO_644 (O_644,N_24127,N_24414);
xnor UO_645 (O_645,N_23506,N_22349);
or UO_646 (O_646,N_22357,N_24141);
nor UO_647 (O_647,N_22647,N_23708);
xnor UO_648 (O_648,N_23551,N_24871);
or UO_649 (O_649,N_23044,N_24136);
and UO_650 (O_650,N_24258,N_24415);
nor UO_651 (O_651,N_21954,N_24903);
xor UO_652 (O_652,N_23522,N_23794);
xor UO_653 (O_653,N_22698,N_22645);
and UO_654 (O_654,N_23119,N_22452);
nand UO_655 (O_655,N_24828,N_24188);
and UO_656 (O_656,N_22003,N_22099);
or UO_657 (O_657,N_22109,N_22433);
xor UO_658 (O_658,N_23610,N_23578);
and UO_659 (O_659,N_22221,N_24902);
or UO_660 (O_660,N_24813,N_24809);
or UO_661 (O_661,N_23703,N_23547);
and UO_662 (O_662,N_22405,N_23701);
nand UO_663 (O_663,N_23297,N_24692);
nor UO_664 (O_664,N_24459,N_24590);
nor UO_665 (O_665,N_22415,N_24347);
nand UO_666 (O_666,N_22334,N_24287);
and UO_667 (O_667,N_22854,N_23669);
and UO_668 (O_668,N_24916,N_24342);
nor UO_669 (O_669,N_24829,N_24019);
or UO_670 (O_670,N_23270,N_22141);
xor UO_671 (O_671,N_24271,N_23922);
nor UO_672 (O_672,N_22892,N_23540);
or UO_673 (O_673,N_22159,N_21919);
or UO_674 (O_674,N_24959,N_22426);
or UO_675 (O_675,N_24852,N_24727);
nand UO_676 (O_676,N_24338,N_22906);
and UO_677 (O_677,N_24343,N_23293);
and UO_678 (O_678,N_23376,N_23957);
nand UO_679 (O_679,N_23905,N_21988);
and UO_680 (O_680,N_23385,N_24445);
nand UO_681 (O_681,N_24884,N_23154);
nand UO_682 (O_682,N_24594,N_24017);
nor UO_683 (O_683,N_23060,N_22251);
or UO_684 (O_684,N_22644,N_22476);
nand UO_685 (O_685,N_22309,N_23229);
or UO_686 (O_686,N_22491,N_24269);
nand UO_687 (O_687,N_23822,N_23353);
nor UO_688 (O_688,N_22390,N_22825);
xnor UO_689 (O_689,N_22706,N_23571);
and UO_690 (O_690,N_24703,N_24184);
xnor UO_691 (O_691,N_22132,N_22874);
nand UO_692 (O_692,N_22696,N_23505);
xor UO_693 (O_693,N_23557,N_24567);
and UO_694 (O_694,N_23323,N_23503);
xor UO_695 (O_695,N_24539,N_22596);
xor UO_696 (O_696,N_23676,N_23032);
or UO_697 (O_697,N_24706,N_23284);
nor UO_698 (O_698,N_23700,N_22957);
xnor UO_699 (O_699,N_24661,N_23787);
nor UO_700 (O_700,N_23674,N_22214);
nor UO_701 (O_701,N_23221,N_22563);
nor UO_702 (O_702,N_23124,N_22277);
and UO_703 (O_703,N_24524,N_22788);
nor UO_704 (O_704,N_22235,N_22712);
or UO_705 (O_705,N_24497,N_23033);
xnor UO_706 (O_706,N_22507,N_23953);
nor UO_707 (O_707,N_22954,N_24399);
xor UO_708 (O_708,N_21965,N_21993);
nand UO_709 (O_709,N_24542,N_22804);
and UO_710 (O_710,N_23907,N_22094);
xnor UO_711 (O_711,N_24739,N_24009);
and UO_712 (O_712,N_24491,N_24275);
xnor UO_713 (O_713,N_24092,N_24153);
nand UO_714 (O_714,N_23516,N_22665);
and UO_715 (O_715,N_22879,N_23699);
or UO_716 (O_716,N_23340,N_24979);
and UO_717 (O_717,N_23848,N_24331);
and UO_718 (O_718,N_24222,N_24233);
nor UO_719 (O_719,N_22049,N_24172);
xor UO_720 (O_720,N_22286,N_23962);
or UO_721 (O_721,N_24004,N_23772);
and UO_722 (O_722,N_24011,N_23352);
or UO_723 (O_723,N_24280,N_22443);
xnor UO_724 (O_724,N_22460,N_24173);
nor UO_725 (O_725,N_23205,N_24231);
nand UO_726 (O_726,N_22467,N_24033);
nand UO_727 (O_727,N_24116,N_22019);
nor UO_728 (O_728,N_23061,N_23348);
or UO_729 (O_729,N_23825,N_24344);
nor UO_730 (O_730,N_23482,N_23785);
nor UO_731 (O_731,N_22383,N_22523);
or UO_732 (O_732,N_22540,N_22943);
or UO_733 (O_733,N_23442,N_24036);
xnor UO_734 (O_734,N_23835,N_23918);
xnor UO_735 (O_735,N_24038,N_22671);
and UO_736 (O_736,N_23997,N_22076);
and UO_737 (O_737,N_21989,N_23491);
and UO_738 (O_738,N_23414,N_24439);
xor UO_739 (O_739,N_24345,N_24709);
xnor UO_740 (O_740,N_21970,N_23834);
or UO_741 (O_741,N_22678,N_24193);
xnor UO_742 (O_742,N_24595,N_23426);
xor UO_743 (O_743,N_24811,N_23654);
xor UO_744 (O_744,N_23622,N_24927);
xnor UO_745 (O_745,N_23370,N_24631);
and UO_746 (O_746,N_24528,N_22597);
xor UO_747 (O_747,N_22376,N_23542);
xnor UO_748 (O_748,N_22152,N_23689);
nand UO_749 (O_749,N_22004,N_22018);
nor UO_750 (O_750,N_24778,N_23811);
or UO_751 (O_751,N_24689,N_22087);
and UO_752 (O_752,N_22727,N_23781);
nand UO_753 (O_753,N_24565,N_23851);
nand UO_754 (O_754,N_24393,N_23243);
and UO_755 (O_755,N_23486,N_22302);
or UO_756 (O_756,N_23252,N_22438);
and UO_757 (O_757,N_22588,N_22818);
nor UO_758 (O_758,N_22928,N_24832);
or UO_759 (O_759,N_22079,N_24401);
or UO_760 (O_760,N_23705,N_23973);
xnor UO_761 (O_761,N_22369,N_22680);
or UO_762 (O_762,N_24448,N_22492);
nand UO_763 (O_763,N_22757,N_23815);
nor UO_764 (O_764,N_22593,N_24617);
xnor UO_765 (O_765,N_21932,N_22841);
xor UO_766 (O_766,N_24596,N_24356);
nand UO_767 (O_767,N_22568,N_23038);
nand UO_768 (O_768,N_22751,N_22855);
and UO_769 (O_769,N_23812,N_22455);
nor UO_770 (O_770,N_22524,N_23910);
xnor UO_771 (O_771,N_23965,N_22207);
and UO_772 (O_772,N_23945,N_23590);
xnor UO_773 (O_773,N_23309,N_24055);
xnor UO_774 (O_774,N_23204,N_21878);
or UO_775 (O_775,N_23492,N_23948);
and UO_776 (O_776,N_24050,N_22851);
xnor UO_777 (O_777,N_23724,N_22868);
or UO_778 (O_778,N_23199,N_23242);
or UO_779 (O_779,N_24265,N_22666);
and UO_780 (O_780,N_23919,N_23914);
xor UO_781 (O_781,N_24314,N_22990);
xor UO_782 (O_782,N_23158,N_23984);
xor UO_783 (O_783,N_22656,N_23259);
nand UO_784 (O_784,N_23374,N_24686);
and UO_785 (O_785,N_22710,N_24929);
nand UO_786 (O_786,N_23027,N_22686);
xor UO_787 (O_787,N_23471,N_22261);
xnor UO_788 (O_788,N_24861,N_21907);
and UO_789 (O_789,N_22648,N_23801);
nor UO_790 (O_790,N_23481,N_24777);
or UO_791 (O_791,N_24118,N_24919);
and UO_792 (O_792,N_22557,N_23063);
or UO_793 (O_793,N_24659,N_24820);
nor UO_794 (O_794,N_22979,N_24475);
or UO_795 (O_795,N_24625,N_22674);
or UO_796 (O_796,N_23396,N_24168);
xnor UO_797 (O_797,N_24750,N_23950);
nor UO_798 (O_798,N_22161,N_24493);
nor UO_799 (O_799,N_24877,N_24283);
nand UO_800 (O_800,N_21992,N_22504);
xor UO_801 (O_801,N_22661,N_22064);
nor UO_802 (O_802,N_22200,N_24016);
and UO_803 (O_803,N_24186,N_21933);
xnor UO_804 (O_804,N_23579,N_23447);
or UO_805 (O_805,N_22724,N_22181);
and UO_806 (O_806,N_24097,N_22162);
nand UO_807 (O_807,N_22711,N_22283);
and UO_808 (O_808,N_24575,N_24977);
nand UO_809 (O_809,N_21898,N_22630);
nand UO_810 (O_810,N_24818,N_22360);
or UO_811 (O_811,N_22700,N_23499);
or UO_812 (O_812,N_24384,N_23042);
xor UO_813 (O_813,N_22133,N_23598);
and UO_814 (O_814,N_23618,N_24980);
or UO_815 (O_815,N_24062,N_23469);
nor UO_816 (O_816,N_24710,N_23467);
or UO_817 (O_817,N_23789,N_23405);
nor UO_818 (O_818,N_24923,N_23882);
nor UO_819 (O_819,N_24458,N_23795);
or UO_820 (O_820,N_24735,N_23020);
or UO_821 (O_821,N_21913,N_22156);
nor UO_822 (O_822,N_23194,N_23236);
nor UO_823 (O_823,N_24975,N_22394);
nand UO_824 (O_824,N_23824,N_23180);
xor UO_825 (O_825,N_22149,N_22618);
nand UO_826 (O_826,N_22735,N_22754);
nand UO_827 (O_827,N_22840,N_22080);
nand UO_828 (O_828,N_24020,N_23969);
nor UO_829 (O_829,N_24315,N_24589);
and UO_830 (O_830,N_23806,N_24788);
or UO_831 (O_831,N_21931,N_24083);
nor UO_832 (O_832,N_23507,N_22931);
xnor UO_833 (O_833,N_24774,N_24388);
xnor UO_834 (O_834,N_22126,N_22404);
nor UO_835 (O_835,N_24227,N_24385);
nor UO_836 (O_836,N_22052,N_22352);
nor UO_837 (O_837,N_23711,N_23473);
xnor UO_838 (O_838,N_24425,N_23707);
nor UO_839 (O_839,N_24958,N_24654);
nor UO_840 (O_840,N_22280,N_24361);
and UO_841 (O_841,N_24981,N_22878);
and UO_842 (O_842,N_23929,N_23456);
nand UO_843 (O_843,N_22672,N_22089);
xor UO_844 (O_844,N_24874,N_23797);
and UO_845 (O_845,N_22071,N_24224);
or UO_846 (O_846,N_24110,N_22316);
or UO_847 (O_847,N_24754,N_24091);
nand UO_848 (O_848,N_22625,N_23668);
and UO_849 (O_849,N_24537,N_23563);
and UO_850 (O_850,N_24702,N_23321);
xor UO_851 (O_851,N_22298,N_22748);
nor UO_852 (O_852,N_21881,N_24708);
and UO_853 (O_853,N_23648,N_23366);
nand UO_854 (O_854,N_24858,N_22013);
or UO_855 (O_855,N_21953,N_22886);
xnor UO_856 (O_856,N_23989,N_24366);
and UO_857 (O_857,N_23745,N_24950);
xor UO_858 (O_858,N_22573,N_22291);
or UO_859 (O_859,N_23792,N_23981);
nand UO_860 (O_860,N_24526,N_24308);
xnor UO_861 (O_861,N_22697,N_22193);
xnor UO_862 (O_862,N_22707,N_21903);
nand UO_863 (O_863,N_23301,N_23763);
xnor UO_864 (O_864,N_23513,N_21924);
nor UO_865 (O_865,N_23151,N_22539);
xnor UO_866 (O_866,N_24833,N_23372);
nand UO_867 (O_867,N_23833,N_24734);
or UO_868 (O_868,N_23863,N_24566);
nor UO_869 (O_869,N_22624,N_23318);
nand UO_870 (O_870,N_23717,N_21876);
nand UO_871 (O_871,N_23478,N_24056);
or UO_872 (O_872,N_22253,N_23127);
or UO_873 (O_873,N_22043,N_22833);
xor UO_874 (O_874,N_24447,N_23520);
nand UO_875 (O_875,N_22420,N_23946);
nor UO_876 (O_876,N_23568,N_24688);
nor UO_877 (O_877,N_23874,N_22121);
nor UO_878 (O_878,N_22347,N_23913);
nand UO_879 (O_879,N_22021,N_22395);
nand UO_880 (O_880,N_22002,N_23359);
nor UO_881 (O_881,N_22228,N_23217);
xor UO_882 (O_882,N_24015,N_22007);
xnor UO_883 (O_883,N_23438,N_22024);
nand UO_884 (O_884,N_23747,N_22914);
nand UO_885 (O_885,N_24489,N_24079);
nand UO_886 (O_886,N_23074,N_22143);
or UO_887 (O_887,N_23762,N_24248);
xor UO_888 (O_888,N_23207,N_22617);
and UO_889 (O_889,N_23415,N_22994);
nand UO_890 (O_890,N_22975,N_24241);
nand UO_891 (O_891,N_23490,N_24808);
nor UO_892 (O_892,N_22392,N_24588);
or UO_893 (O_893,N_24043,N_21999);
and UO_894 (O_894,N_24530,N_22526);
and UO_895 (O_895,N_22222,N_24915);
or UO_896 (O_896,N_24610,N_24049);
nand UO_897 (O_897,N_24603,N_24073);
nor UO_898 (O_898,N_24711,N_22750);
and UO_899 (O_899,N_22382,N_24502);
nand UO_900 (O_900,N_22227,N_22856);
nor UO_901 (O_901,N_24151,N_24577);
xnor UO_902 (O_902,N_22380,N_24108);
nand UO_903 (O_903,N_22922,N_22270);
and UO_904 (O_904,N_22364,N_24471);
or UO_905 (O_905,N_23355,N_23218);
and UO_906 (O_906,N_23495,N_23025);
xor UO_907 (O_907,N_23330,N_22883);
nand UO_908 (O_908,N_22158,N_24031);
or UO_909 (O_909,N_24191,N_23454);
nor UO_910 (O_910,N_23872,N_22399);
and UO_911 (O_911,N_23019,N_22142);
nor UO_912 (O_912,N_22581,N_24311);
and UO_913 (O_913,N_21912,N_23206);
xnor UO_914 (O_914,N_24885,N_22905);
xnor UO_915 (O_915,N_22691,N_24882);
xnor UO_916 (O_916,N_23581,N_22375);
xnor UO_917 (O_917,N_23613,N_24107);
xor UO_918 (O_918,N_23982,N_24928);
or UO_919 (O_919,N_24147,N_22275);
and UO_920 (O_920,N_23653,N_24581);
nor UO_921 (O_921,N_22173,N_24137);
nor UO_922 (O_922,N_21948,N_22760);
or UO_923 (O_923,N_23484,N_22123);
xnor UO_924 (O_924,N_24562,N_24174);
xnor UO_925 (O_925,N_22134,N_22813);
nand UO_926 (O_926,N_22103,N_23028);
and UO_927 (O_927,N_23007,N_22128);
or UO_928 (O_928,N_22090,N_23881);
xor UO_929 (O_929,N_22799,N_22137);
nand UO_930 (O_930,N_24282,N_24510);
or UO_931 (O_931,N_23561,N_22178);
xor UO_932 (O_932,N_24521,N_22055);
xor UO_933 (O_933,N_24856,N_22850);
nand UO_934 (O_934,N_24387,N_22472);
or UO_935 (O_935,N_22902,N_23126);
xor UO_936 (O_936,N_23065,N_22537);
and UO_937 (O_937,N_24089,N_22610);
nor UO_938 (O_938,N_24772,N_23941);
and UO_939 (O_939,N_23855,N_24648);
nor UO_940 (O_940,N_22553,N_24514);
nand UO_941 (O_941,N_22439,N_24413);
or UO_942 (O_942,N_23736,N_22608);
or UO_943 (O_943,N_24662,N_24404);
xor UO_944 (O_944,N_24839,N_22225);
or UO_945 (O_945,N_22312,N_23113);
and UO_946 (O_946,N_23809,N_24822);
and UO_947 (O_947,N_22118,N_22965);
nand UO_948 (O_948,N_23143,N_21983);
xor UO_949 (O_949,N_23771,N_23213);
nand UO_950 (O_950,N_22501,N_22497);
nor UO_951 (O_951,N_22907,N_22631);
or UO_952 (O_952,N_23959,N_22058);
and UO_953 (O_953,N_22379,N_23680);
or UO_954 (O_954,N_22599,N_23652);
xor UO_955 (O_955,N_23784,N_24619);
or UO_956 (O_956,N_22538,N_24010);
nand UO_957 (O_957,N_24230,N_23679);
nor UO_958 (O_958,N_23276,N_23390);
and UO_959 (O_959,N_24516,N_23493);
nor UO_960 (O_960,N_22918,N_24357);
nor UO_961 (O_961,N_22324,N_24294);
nor UO_962 (O_962,N_24910,N_24477);
nand UO_963 (O_963,N_23776,N_23924);
nand UO_964 (O_964,N_24183,N_22012);
nor UO_965 (O_965,N_22720,N_23100);
and UO_966 (O_966,N_23788,N_23081);
xor UO_967 (O_967,N_22535,N_23131);
nor UO_968 (O_968,N_23203,N_24454);
nor UO_969 (O_969,N_21890,N_22925);
nand UO_970 (O_970,N_24655,N_24377);
and UO_971 (O_971,N_22138,N_23936);
nand UO_972 (O_972,N_24715,N_23209);
nand UO_973 (O_973,N_22468,N_22238);
nor UO_974 (O_974,N_24701,N_24803);
nand UO_975 (O_975,N_22998,N_22157);
nor UO_976 (O_976,N_23560,N_22937);
xnor UO_977 (O_977,N_24000,N_22389);
nor UO_978 (O_978,N_22403,N_24725);
xor UO_979 (O_979,N_22418,N_22518);
nand UO_980 (O_980,N_23083,N_24037);
or UO_981 (O_981,N_22550,N_23191);
or UO_982 (O_982,N_24554,N_24503);
and UO_983 (O_983,N_24072,N_24868);
xnor UO_984 (O_984,N_21997,N_23152);
nand UO_985 (O_985,N_22031,N_24473);
nor UO_986 (O_986,N_22028,N_23269);
nand UO_987 (O_987,N_22622,N_23725);
nand UO_988 (O_988,N_24506,N_22901);
and UO_989 (O_989,N_24569,N_24463);
xor UO_990 (O_990,N_22515,N_24176);
nor UO_991 (O_991,N_22125,N_24400);
or UO_992 (O_992,N_23135,N_23116);
or UO_993 (O_993,N_23888,N_23567);
or UO_994 (O_994,N_23150,N_23737);
nor UO_995 (O_995,N_23412,N_24068);
nand UO_996 (O_996,N_22978,N_22913);
nand UO_997 (O_997,N_24309,N_22258);
nand UO_998 (O_998,N_22336,N_22827);
nor UO_999 (O_999,N_23022,N_24268);
nor UO_1000 (O_1000,N_21895,N_22870);
nand UO_1001 (O_1001,N_24546,N_24262);
and UO_1002 (O_1002,N_22236,N_24691);
nand UO_1003 (O_1003,N_22849,N_21969);
nor UO_1004 (O_1004,N_23090,N_23468);
xnor UO_1005 (O_1005,N_23155,N_24638);
nand UO_1006 (O_1006,N_22295,N_24125);
or UO_1007 (O_1007,N_23951,N_23262);
or UO_1008 (O_1008,N_23909,N_24194);
xnor UO_1009 (O_1009,N_23271,N_22397);
nand UO_1010 (O_1010,N_24159,N_22871);
nor UO_1011 (O_1011,N_22530,N_22679);
nand UO_1012 (O_1012,N_24805,N_23850);
and UO_1013 (O_1013,N_23176,N_24866);
nand UO_1014 (O_1014,N_23338,N_22794);
nor UO_1015 (O_1015,N_22474,N_24545);
xnor UO_1016 (O_1016,N_22209,N_23477);
nor UO_1017 (O_1017,N_24199,N_23480);
nor UO_1018 (O_1018,N_23141,N_24117);
nand UO_1019 (O_1019,N_22473,N_24740);
nand UO_1020 (O_1020,N_22845,N_22259);
or UO_1021 (O_1021,N_23443,N_22254);
nor UO_1022 (O_1022,N_23108,N_24579);
nand UO_1023 (O_1023,N_23086,N_22469);
nor UO_1024 (O_1024,N_24005,N_22891);
nor UO_1025 (O_1025,N_22111,N_24797);
xnor UO_1026 (O_1026,N_22244,N_24349);
nor UO_1027 (O_1027,N_24517,N_23960);
nor UO_1028 (O_1028,N_22810,N_22184);
or UO_1029 (O_1029,N_22517,N_24200);
xor UO_1030 (O_1030,N_22921,N_22359);
xnor UO_1031 (O_1031,N_22032,N_22417);
or UO_1032 (O_1032,N_22960,N_23891);
nor UO_1033 (O_1033,N_22000,N_24761);
nor UO_1034 (O_1034,N_24831,N_21904);
and UO_1035 (O_1035,N_24390,N_22932);
nand UO_1036 (O_1036,N_22558,N_22985);
and UO_1037 (O_1037,N_22786,N_24135);
nand UO_1038 (O_1038,N_23462,N_21894);
nand UO_1039 (O_1039,N_24536,N_22290);
and UO_1040 (O_1040,N_23586,N_24888);
nand UO_1041 (O_1041,N_22741,N_22982);
or UO_1042 (O_1042,N_22807,N_22749);
xnor UO_1043 (O_1043,N_23971,N_23220);
nor UO_1044 (O_1044,N_22350,N_22974);
nor UO_1045 (O_1045,N_24947,N_22326);
nor UO_1046 (O_1046,N_24067,N_22981);
or UO_1047 (O_1047,N_22124,N_23606);
nand UO_1048 (O_1048,N_23129,N_23178);
and UO_1049 (O_1049,N_21980,N_23128);
xor UO_1050 (O_1050,N_22574,N_23600);
or UO_1051 (O_1051,N_22717,N_23306);
xor UO_1052 (O_1052,N_24994,N_22419);
and UO_1053 (O_1053,N_23335,N_23655);
nor UO_1054 (O_1054,N_22576,N_23921);
nand UO_1055 (O_1055,N_22642,N_22519);
and UO_1056 (O_1056,N_24039,N_24764);
or UO_1057 (O_1057,N_24490,N_24663);
or UO_1058 (O_1058,N_22955,N_23935);
nand UO_1059 (O_1059,N_24229,N_22330);
xor UO_1060 (O_1060,N_24438,N_22398);
or UO_1061 (O_1061,N_23233,N_23770);
or UO_1062 (O_1062,N_23322,N_23758);
and UO_1063 (O_1063,N_24541,N_23569);
xnor UO_1064 (O_1064,N_24359,N_23280);
or UO_1065 (O_1065,N_24551,N_23144);
or UO_1066 (O_1066,N_22823,N_22462);
xor UO_1067 (O_1067,N_24834,N_24205);
xor UO_1068 (O_1068,N_22942,N_23115);
or UO_1069 (O_1069,N_24228,N_24534);
nor UO_1070 (O_1070,N_23582,N_23621);
nand UO_1071 (O_1071,N_24432,N_23746);
nor UO_1072 (O_1072,N_23584,N_23926);
or UO_1073 (O_1073,N_24163,N_24305);
or UO_1074 (O_1074,N_21979,N_22667);
nand UO_1075 (O_1075,N_24585,N_23757);
nand UO_1076 (O_1076,N_23453,N_23035);
or UO_1077 (O_1077,N_24757,N_23755);
nor UO_1078 (O_1078,N_23715,N_24963);
or UO_1079 (O_1079,N_23663,N_22450);
xor UO_1080 (O_1080,N_22505,N_23673);
and UO_1081 (O_1081,N_23623,N_23609);
nor UO_1082 (O_1082,N_24564,N_23566);
nand UO_1083 (O_1083,N_22814,N_22447);
xnor UO_1084 (O_1084,N_23631,N_23908);
or UO_1085 (O_1085,N_24018,N_22422);
xnor UO_1086 (O_1086,N_23983,N_24488);
and UO_1087 (O_1087,N_23852,N_22626);
and UO_1088 (O_1088,N_22956,N_22195);
nor UO_1089 (O_1089,N_23892,N_23659);
nand UO_1090 (O_1090,N_22006,N_23866);
or UO_1091 (O_1091,N_24911,N_22594);
nand UO_1092 (O_1092,N_23832,N_22646);
nor UO_1093 (O_1093,N_22430,N_24034);
xnor UO_1094 (O_1094,N_24786,N_22601);
nor UO_1095 (O_1095,N_22085,N_22475);
nand UO_1096 (O_1096,N_24483,N_23421);
or UO_1097 (O_1097,N_24974,N_23171);
nand UO_1098 (O_1098,N_24798,N_22348);
and UO_1099 (O_1099,N_23974,N_22938);
nand UO_1100 (O_1100,N_22029,N_24087);
xor UO_1101 (O_1101,N_24462,N_22503);
or UO_1102 (O_1102,N_23245,N_23958);
or UO_1103 (O_1103,N_23894,N_21958);
nor UO_1104 (O_1104,N_24897,N_22185);
and UO_1105 (O_1105,N_23244,N_22313);
or UO_1106 (O_1106,N_24598,N_22579);
nand UO_1107 (O_1107,N_22276,N_22105);
xor UO_1108 (O_1108,N_23871,N_23186);
xnor UO_1109 (O_1109,N_24555,N_23029);
xnor UO_1110 (O_1110,N_23502,N_23026);
nand UO_1111 (O_1111,N_24992,N_22321);
nor UO_1112 (O_1112,N_23014,N_22411);
nand UO_1113 (O_1113,N_22429,N_24680);
and UO_1114 (O_1114,N_22763,N_22924);
xnor UO_1115 (O_1115,N_23488,N_22441);
xor UO_1116 (O_1116,N_22241,N_23452);
xnor UO_1117 (O_1117,N_24246,N_24171);
xor UO_1118 (O_1118,N_22541,N_22893);
or UO_1119 (O_1119,N_24848,N_24099);
xnor UO_1120 (O_1120,N_23543,N_23783);
or UO_1121 (O_1121,N_24418,N_22800);
or UO_1122 (O_1122,N_23459,N_22887);
or UO_1123 (O_1123,N_24203,N_24351);
nor UO_1124 (O_1124,N_22790,N_22311);
nand UO_1125 (O_1125,N_23696,N_22633);
or UO_1126 (O_1126,N_21920,N_23416);
nor UO_1127 (O_1127,N_24674,N_24650);
or UO_1128 (O_1128,N_24922,N_23966);
nor UO_1129 (O_1129,N_22262,N_22378);
or UO_1130 (O_1130,N_24480,N_23079);
nor UO_1131 (O_1131,N_22861,N_24815);
and UO_1132 (O_1132,N_22949,N_23004);
xnor UO_1133 (O_1133,N_24694,N_24369);
nand UO_1134 (O_1134,N_24713,N_24259);
and UO_1135 (O_1135,N_22992,N_22842);
nor UO_1136 (O_1136,N_24746,N_24730);
xor UO_1137 (O_1137,N_22778,N_23091);
and UO_1138 (O_1138,N_23841,N_23638);
xor UO_1139 (O_1139,N_22961,N_22346);
xnor UO_1140 (O_1140,N_23400,N_22337);
nand UO_1141 (O_1141,N_24759,N_23212);
nor UO_1142 (O_1142,N_24468,N_23389);
nand UO_1143 (O_1143,N_22053,N_24180);
and UO_1144 (O_1144,N_22199,N_24256);
xnor UO_1145 (O_1145,N_24419,N_22834);
xnor UO_1146 (O_1146,N_23644,N_22150);
and UO_1147 (O_1147,N_24507,N_22527);
or UO_1148 (O_1148,N_22057,N_21957);
nand UO_1149 (O_1149,N_23286,N_23448);
nand UO_1150 (O_1150,N_24558,N_23101);
nor UO_1151 (O_1151,N_23140,N_24114);
or UO_1152 (O_1152,N_24061,N_24245);
xor UO_1153 (O_1153,N_23672,N_24263);
and UO_1154 (O_1154,N_22054,N_22703);
nand UO_1155 (O_1155,N_24799,N_22592);
and UO_1156 (O_1156,N_22136,N_22187);
nor UO_1157 (O_1157,N_23976,N_24386);
xnor UO_1158 (O_1158,N_23728,N_24532);
nand UO_1159 (O_1159,N_23970,N_22510);
or UO_1160 (O_1160,N_23395,N_24325);
xor UO_1161 (O_1161,N_24914,N_23928);
and UO_1162 (O_1162,N_22067,N_23333);
or UO_1163 (O_1163,N_24982,N_24743);
and UO_1164 (O_1164,N_22809,N_24593);
nand UO_1165 (O_1165,N_22926,N_24785);
xnor UO_1166 (O_1166,N_22412,N_22204);
or UO_1167 (O_1167,N_23730,N_23995);
xor UO_1168 (O_1168,N_24106,N_21978);
xnor UO_1169 (O_1169,N_23002,N_24908);
or UO_1170 (O_1170,N_23260,N_24101);
or UO_1171 (O_1171,N_23559,N_24474);
nor UO_1172 (O_1172,N_22659,N_22619);
or UO_1173 (O_1173,N_24424,N_24736);
nand UO_1174 (O_1174,N_23767,N_23607);
and UO_1175 (O_1175,N_24192,N_23985);
or UO_1176 (O_1176,N_23688,N_22073);
xor UO_1177 (O_1177,N_24945,N_22614);
and UO_1178 (O_1178,N_23923,N_24515);
or UO_1179 (O_1179,N_23813,N_24302);
and UO_1180 (O_1180,N_24242,N_24853);
or UO_1181 (O_1181,N_22166,N_24060);
and UO_1182 (O_1182,N_22670,N_24429);
or UO_1183 (O_1183,N_24084,N_24614);
or UO_1184 (O_1184,N_22988,N_22319);
and UO_1185 (O_1185,N_24426,N_23741);
xor UO_1186 (O_1186,N_23077,N_22889);
and UO_1187 (O_1187,N_24637,N_24938);
xnor UO_1188 (O_1188,N_23714,N_22923);
nand UO_1189 (O_1189,N_23343,N_22260);
nand UO_1190 (O_1190,N_23403,N_24953);
nor UO_1191 (O_1191,N_24300,N_22819);
nor UO_1192 (O_1192,N_21950,N_23614);
xor UO_1193 (O_1193,N_22556,N_24148);
nor UO_1194 (O_1194,N_24146,N_24210);
nand UO_1195 (O_1195,N_23647,N_23134);
nand UO_1196 (O_1196,N_22876,N_23106);
xnor UO_1197 (O_1197,N_24823,N_24646);
or UO_1198 (O_1198,N_22372,N_23709);
nand UO_1199 (O_1199,N_23064,N_24677);
xor UO_1200 (O_1200,N_23528,N_24252);
nand UO_1201 (O_1201,N_22881,N_23544);
and UO_1202 (O_1202,N_22393,N_22733);
nand UO_1203 (O_1203,N_23040,N_22299);
or UO_1204 (O_1204,N_23510,N_21897);
or UO_1205 (O_1205,N_22899,N_24851);
nand UO_1206 (O_1206,N_23036,N_24900);
or UO_1207 (O_1207,N_23853,N_23475);
nor UO_1208 (O_1208,N_22583,N_24773);
xor UO_1209 (O_1209,N_22547,N_21937);
and UO_1210 (O_1210,N_22465,N_23279);
nor UO_1211 (O_1211,N_24501,N_22120);
xor UO_1212 (O_1212,N_24323,N_21911);
and UO_1213 (O_1213,N_22490,N_24630);
xor UO_1214 (O_1214,N_24225,N_24411);
and UO_1215 (O_1215,N_22773,N_22865);
nand UO_1216 (O_1216,N_22167,N_23381);
nor UO_1217 (O_1217,N_23665,N_22890);
or UO_1218 (O_1218,N_23261,N_23889);
xnor UO_1219 (O_1219,N_24371,N_22135);
and UO_1220 (O_1220,N_23920,N_23558);
nor UO_1221 (O_1221,N_23005,N_23075);
nand UO_1222 (O_1222,N_22828,N_21960);
nand UO_1223 (O_1223,N_22940,N_22770);
xnor UO_1224 (O_1224,N_24547,N_23130);
nor UO_1225 (O_1225,N_22777,N_22226);
and UO_1226 (O_1226,N_22096,N_24651);
and UO_1227 (O_1227,N_22461,N_24324);
and UO_1228 (O_1228,N_23532,N_22335);
or UO_1229 (O_1229,N_23799,N_24333);
nor UO_1230 (O_1230,N_22263,N_24001);
and UO_1231 (O_1231,N_22572,N_23394);
xor UO_1232 (O_1232,N_22434,N_23094);
and UO_1233 (O_1233,N_22649,N_22194);
xor UO_1234 (O_1234,N_22494,N_22976);
nand UO_1235 (O_1235,N_24789,N_24035);
and UO_1236 (O_1236,N_23070,N_23291);
and UO_1237 (O_1237,N_22759,N_21929);
nor UO_1238 (O_1238,N_24221,N_23633);
nand UO_1239 (O_1239,N_24742,N_22197);
and UO_1240 (O_1240,N_24841,N_23605);
and UO_1241 (O_1241,N_22655,N_22946);
or UO_1242 (O_1242,N_24582,N_23643);
nand UO_1243 (O_1243,N_23177,N_23786);
xnor UO_1244 (O_1244,N_22927,N_22011);
and UO_1245 (O_1245,N_23687,N_23818);
or UO_1246 (O_1246,N_24634,N_24120);
nor UO_1247 (O_1247,N_23899,N_22448);
nor UO_1248 (O_1248,N_23430,N_23677);
or UO_1249 (O_1249,N_23455,N_22082);
or UO_1250 (O_1250,N_22292,N_23751);
xnor UO_1251 (O_1251,N_24804,N_23296);
nor UO_1252 (O_1252,N_23664,N_23533);
nand UO_1253 (O_1253,N_23388,N_23021);
nor UO_1254 (O_1254,N_22996,N_24008);
xnor UO_1255 (O_1255,N_24408,N_23215);
and UO_1256 (O_1256,N_24449,N_24213);
nor UO_1257 (O_1257,N_23682,N_23440);
nand UO_1258 (O_1258,N_24940,N_22692);
or UO_1259 (O_1259,N_23365,N_22917);
nor UO_1260 (O_1260,N_23214,N_23964);
nand UO_1261 (O_1261,N_22190,N_23839);
and UO_1262 (O_1262,N_23732,N_23512);
xnor UO_1263 (O_1263,N_23179,N_22673);
nor UO_1264 (O_1264,N_23292,N_24795);
nand UO_1265 (O_1265,N_23302,N_23419);
and UO_1266 (O_1266,N_22189,N_22325);
xnor UO_1267 (O_1267,N_23831,N_22479);
nor UO_1268 (O_1268,N_22728,N_24909);
or UO_1269 (O_1269,N_22787,N_23588);
nand UO_1270 (O_1270,N_24932,N_22709);
or UO_1271 (O_1271,N_24279,N_22154);
nand UO_1272 (O_1272,N_23829,N_24807);
and UO_1273 (O_1273,N_22035,N_23867);
and UO_1274 (O_1274,N_23360,N_24196);
nor UO_1275 (O_1275,N_24024,N_24370);
nor UO_1276 (O_1276,N_24182,N_24441);
and UO_1277 (O_1277,N_23977,N_22950);
or UO_1278 (O_1278,N_24026,N_22224);
nor UO_1279 (O_1279,N_24535,N_24669);
nor UO_1280 (O_1280,N_23761,N_24592);
nand UO_1281 (O_1281,N_23634,N_24814);
or UO_1282 (O_1282,N_21946,N_23875);
nand UO_1283 (O_1283,N_22496,N_24446);
nand UO_1284 (O_1284,N_22183,N_22371);
nand UO_1285 (O_1285,N_22386,N_23555);
or UO_1286 (O_1286,N_23274,N_23947);
or UO_1287 (O_1287,N_24453,N_24875);
or UO_1288 (O_1288,N_22345,N_23023);
nor UO_1289 (O_1289,N_22964,N_23498);
or UO_1290 (O_1290,N_24261,N_23880);
xor UO_1291 (O_1291,N_22487,N_23849);
nand UO_1292 (O_1292,N_22745,N_22650);
xnor UO_1293 (O_1293,N_24479,N_24270);
xnor UO_1294 (O_1294,N_23103,N_24934);
nand UO_1295 (O_1295,N_23030,N_24895);
or UO_1296 (O_1296,N_24793,N_23307);
or UO_1297 (O_1297,N_24728,N_23859);
nand UO_1298 (O_1298,N_23424,N_22915);
nor UO_1299 (O_1299,N_21990,N_23596);
and UO_1300 (O_1300,N_23706,N_24876);
and UO_1301 (O_1301,N_24618,N_24960);
nand UO_1302 (O_1302,N_23684,N_23411);
nor UO_1303 (O_1303,N_24762,N_24098);
nor UO_1304 (O_1304,N_22478,N_24237);
or UO_1305 (O_1305,N_22765,N_23018);
xnor UO_1306 (O_1306,N_23612,N_23182);
or UO_1307 (O_1307,N_22046,N_22171);
nand UO_1308 (O_1308,N_22293,N_22606);
and UO_1309 (O_1309,N_22715,N_23611);
and UO_1310 (O_1310,N_24070,N_24348);
xnor UO_1311 (O_1311,N_22160,N_22551);
xor UO_1312 (O_1312,N_24214,N_22753);
nand UO_1313 (O_1313,N_24967,N_24027);
or UO_1314 (O_1314,N_23649,N_24988);
nand UO_1315 (O_1315,N_24645,N_24883);
nor UO_1316 (O_1316,N_23008,N_21991);
or UO_1317 (O_1317,N_24456,N_22234);
nor UO_1318 (O_1318,N_24381,N_24007);
nand UO_1319 (O_1319,N_22723,N_22718);
or UO_1320 (O_1320,N_24276,N_23972);
xnor UO_1321 (O_1321,N_22100,N_23362);
or UO_1322 (O_1322,N_23048,N_22903);
nand UO_1323 (O_1323,N_22495,N_22332);
nor UO_1324 (O_1324,N_23013,N_24628);
nor UO_1325 (O_1325,N_23132,N_24264);
and UO_1326 (O_1326,N_24760,N_23339);
nand UO_1327 (O_1327,N_22401,N_23798);
or UO_1328 (O_1328,N_24303,N_24330);
xor UO_1329 (O_1329,N_23266,N_23407);
nand UO_1330 (O_1330,N_23230,N_24826);
nor UO_1331 (O_1331,N_21943,N_23697);
xor UO_1332 (O_1332,N_24816,N_23047);
or UO_1333 (O_1333,N_23034,N_24321);
and UO_1334 (O_1334,N_24082,N_22836);
nor UO_1335 (O_1335,N_24749,N_23188);
xor UO_1336 (O_1336,N_24704,N_24234);
and UO_1337 (O_1337,N_21899,N_23556);
nand UO_1338 (O_1338,N_23504,N_21952);
or UO_1339 (O_1339,N_23300,N_21936);
nor UO_1340 (O_1340,N_23431,N_22246);
nor UO_1341 (O_1341,N_22009,N_23597);
xnor UO_1342 (O_1342,N_22912,N_22812);
xor UO_1343 (O_1343,N_23637,N_22470);
or UO_1344 (O_1344,N_24313,N_23817);
nor UO_1345 (O_1345,N_24157,N_24317);
or UO_1346 (O_1346,N_22632,N_24274);
nor UO_1347 (O_1347,N_24124,N_23006);
and UO_1348 (O_1348,N_24296,N_24924);
or UO_1349 (O_1349,N_24077,N_24304);
nand UO_1350 (O_1350,N_24731,N_22179);
or UO_1351 (O_1351,N_24226,N_23860);
and UO_1352 (O_1352,N_24217,N_24611);
nor UO_1353 (O_1353,N_24700,N_23139);
nor UO_1354 (O_1354,N_24048,N_23939);
or UO_1355 (O_1355,N_23721,N_24867);
nand UO_1356 (O_1356,N_23583,N_22609);
and UO_1357 (O_1357,N_24142,N_23843);
nand UO_1358 (O_1358,N_22875,N_23802);
and UO_1359 (O_1359,N_22863,N_22664);
and UO_1360 (O_1360,N_23675,N_23345);
nand UO_1361 (O_1361,N_24360,N_24346);
xnor UO_1362 (O_1362,N_22885,N_22153);
nor UO_1363 (O_1363,N_24779,N_23314);
and UO_1364 (O_1364,N_23097,N_22232);
nand UO_1365 (O_1365,N_22119,N_21889);
or UO_1366 (O_1366,N_22036,N_24673);
nand UO_1367 (O_1367,N_22130,N_24398);
nand UO_1368 (O_1368,N_24544,N_24636);
or UO_1369 (O_1369,N_22066,N_23856);
nand UO_1370 (O_1370,N_24266,N_22255);
or UO_1371 (O_1371,N_21925,N_22653);
xnor UO_1372 (O_1372,N_23192,N_22934);
nor UO_1373 (O_1373,N_24058,N_23361);
xnor UO_1374 (O_1374,N_22839,N_23800);
nand UO_1375 (O_1375,N_24850,N_22078);
nor UO_1376 (O_1376,N_23642,N_22424);
nand UO_1377 (O_1377,N_22373,N_23145);
xor UO_1378 (O_1378,N_22088,N_24970);
xnor UO_1379 (O_1379,N_23738,N_23410);
nand UO_1380 (O_1380,N_23235,N_21940);
or UO_1381 (O_1381,N_23009,N_22151);
or UO_1382 (O_1382,N_24873,N_22140);
and UO_1383 (O_1383,N_24985,N_22050);
nand UO_1384 (O_1384,N_23363,N_24664);
xor UO_1385 (O_1385,N_24724,N_23756);
nor UO_1386 (O_1386,N_24492,N_24935);
nor UO_1387 (O_1387,N_24944,N_24417);
or UO_1388 (O_1388,N_24525,N_22575);
or UO_1389 (O_1389,N_23545,N_24335);
xor UO_1390 (O_1390,N_22713,N_24810);
and UO_1391 (O_1391,N_24837,N_23734);
or UO_1392 (O_1392,N_24212,N_23820);
xor UO_1393 (O_1393,N_24395,N_24405);
and UO_1394 (O_1394,N_24111,N_23912);
or UO_1395 (O_1395,N_23546,N_23228);
xnor UO_1396 (O_1396,N_24320,N_22213);
nor UO_1397 (O_1397,N_22341,N_22250);
or UO_1398 (O_1398,N_24973,N_22027);
and UO_1399 (O_1399,N_22611,N_21966);
nand UO_1400 (O_1400,N_22488,N_23570);
or UO_1401 (O_1401,N_22048,N_23208);
and UO_1402 (O_1402,N_22256,N_24290);
xnor UO_1403 (O_1403,N_24827,N_23865);
or UO_1404 (O_1404,N_21941,N_24352);
or UO_1405 (O_1405,N_23769,N_22328);
xnor UO_1406 (O_1406,N_23427,N_24511);
xor UO_1407 (O_1407,N_24195,N_24267);
xnor UO_1408 (O_1408,N_23417,N_22641);
nand UO_1409 (O_1409,N_23955,N_23398);
or UO_1410 (O_1410,N_22482,N_22176);
nand UO_1411 (O_1411,N_23391,N_22882);
nor UO_1412 (O_1412,N_24391,N_23576);
nor UO_1413 (O_1413,N_21930,N_22306);
or UO_1414 (O_1414,N_22427,N_24679);
nor UO_1415 (O_1415,N_24752,N_22279);
or UO_1416 (O_1416,N_22685,N_22285);
xor UO_1417 (O_1417,N_23593,N_22175);
or UO_1418 (O_1418,N_24962,N_23890);
nand UO_1419 (O_1419,N_23098,N_23163);
xor UO_1420 (O_1420,N_24872,N_22170);
or UO_1421 (O_1421,N_22425,N_23072);
xor UO_1422 (O_1422,N_23268,N_23166);
xnor UO_1423 (O_1423,N_22832,N_24421);
xor UO_1424 (O_1424,N_24931,N_22858);
or UO_1425 (O_1425,N_24504,N_22989);
nor UO_1426 (O_1426,N_24207,N_22613);
nand UO_1427 (O_1427,N_24201,N_23393);
or UO_1428 (O_1428,N_24697,N_24466);
xnor UO_1429 (O_1429,N_23670,N_23956);
nor UO_1430 (O_1430,N_24298,N_22933);
and UO_1431 (O_1431,N_24299,N_23963);
xnor UO_1432 (O_1432,N_24301,N_21900);
and UO_1433 (O_1433,N_24131,N_22536);
or UO_1434 (O_1434,N_23671,N_24059);
or UO_1435 (O_1435,N_22459,N_24156);
or UO_1436 (O_1436,N_23225,N_24285);
xor UO_1437 (O_1437,N_23316,N_24143);
and UO_1438 (O_1438,N_22549,N_23449);
and UO_1439 (O_1439,N_24129,N_22525);
xor UO_1440 (O_1440,N_23078,N_24643);
or UO_1441 (O_1441,N_24119,N_22768);
and UO_1442 (O_1442,N_23759,N_24100);
xor UO_1443 (O_1443,N_22092,N_23181);
xnor UO_1444 (O_1444,N_23537,N_22220);
xnor UO_1445 (O_1445,N_23425,N_24838);
and UO_1446 (O_1446,N_23494,N_24326);
nor UO_1447 (O_1447,N_23661,N_24954);
xor UO_1448 (O_1448,N_23304,N_23173);
nand UO_1449 (O_1449,N_23232,N_24500);
nand UO_1450 (O_1450,N_23312,N_24986);
and UO_1451 (O_1451,N_24433,N_23968);
or UO_1452 (O_1452,N_22521,N_24583);
or UO_1453 (O_1453,N_24239,N_23805);
or UO_1454 (O_1454,N_24849,N_22837);
or UO_1455 (O_1455,N_24396,N_22168);
or UO_1456 (O_1456,N_21963,N_24220);
xor UO_1457 (O_1457,N_22385,N_24615);
nand UO_1458 (O_1458,N_24028,N_23058);
nor UO_1459 (O_1459,N_23017,N_22694);
and UO_1460 (O_1460,N_22206,N_23085);
nor UO_1461 (O_1461,N_24257,N_22310);
or UO_1462 (O_1462,N_24698,N_23518);
nor UO_1463 (O_1463,N_23553,N_23216);
nor UO_1464 (O_1464,N_24678,N_22268);
nor UO_1465 (O_1465,N_24755,N_23000);
nand UO_1466 (O_1466,N_24375,N_23489);
nand UO_1467 (O_1467,N_23003,N_23337);
xor UO_1468 (O_1468,N_24358,N_22562);
nand UO_1469 (O_1469,N_24623,N_22514);
nor UO_1470 (O_1470,N_24336,N_23265);
nand UO_1471 (O_1471,N_23943,N_23170);
and UO_1472 (O_1472,N_24286,N_24130);
or UO_1473 (O_1473,N_24794,N_24372);
and UO_1474 (O_1474,N_22075,N_22743);
nand UO_1475 (O_1475,N_23120,N_23011);
xnor UO_1476 (O_1476,N_22110,N_24198);
xnor UO_1477 (O_1477,N_23760,N_22775);
and UO_1478 (O_1478,N_23441,N_22607);
xnor UO_1479 (O_1479,N_23156,N_22499);
nor UO_1480 (O_1480,N_23344,N_22654);
and UO_1481 (O_1481,N_22898,N_23275);
nand UO_1482 (O_1482,N_24642,N_24002);
nor UO_1483 (O_1483,N_24821,N_24641);
nor UO_1484 (O_1484,N_22835,N_23565);
xnor UO_1485 (O_1485,N_22015,N_24898);
or UO_1486 (O_1486,N_22862,N_22414);
and UO_1487 (O_1487,N_24389,N_23595);
xor UO_1488 (O_1488,N_23896,N_24316);
xnor UO_1489 (O_1489,N_24609,N_22952);
or UO_1490 (O_1490,N_23515,N_23198);
or UO_1491 (O_1491,N_23012,N_23635);
xnor UO_1492 (O_1492,N_24235,N_21961);
xor UO_1493 (O_1493,N_22436,N_21875);
nor UO_1494 (O_1494,N_22083,N_21917);
nand UO_1495 (O_1495,N_22877,N_23885);
and UO_1496 (O_1496,N_24599,N_24328);
nor UO_1497 (O_1497,N_22947,N_22605);
or UO_1498 (O_1498,N_24512,N_22155);
or UO_1499 (O_1499,N_23933,N_23713);
and UO_1500 (O_1500,N_24442,N_24629);
or UO_1501 (O_1501,N_23485,N_23807);
or UO_1502 (O_1502,N_24859,N_22074);
nor UO_1503 (O_1503,N_21910,N_23752);
nand UO_1504 (O_1504,N_24937,N_22776);
nor UO_1505 (O_1505,N_22237,N_24255);
or UO_1506 (O_1506,N_22266,N_24626);
and UO_1507 (O_1507,N_24572,N_24864);
or UO_1508 (O_1508,N_22900,N_24046);
xor UO_1509 (O_1509,N_23816,N_22093);
and UO_1510 (O_1510,N_24052,N_23743);
and UO_1511 (O_1511,N_24185,N_22435);
nand UO_1512 (O_1512,N_22991,N_24690);
nor UO_1513 (O_1513,N_22930,N_24329);
nor UO_1514 (O_1514,N_22620,N_24066);
and UO_1515 (O_1515,N_24857,N_23845);
and UO_1516 (O_1516,N_22719,N_23549);
nand UO_1517 (O_1517,N_23197,N_23693);
nor UO_1518 (O_1518,N_22993,N_23868);
xnor UO_1519 (O_1519,N_23531,N_23465);
and UO_1520 (O_1520,N_23591,N_24051);
and UO_1521 (O_1521,N_22792,N_24065);
and UO_1522 (O_1522,N_22218,N_22969);
nor UO_1523 (O_1523,N_22453,N_23927);
nand UO_1524 (O_1524,N_23254,N_23793);
and UO_1525 (O_1525,N_22935,N_22687);
nor UO_1526 (O_1526,N_22824,N_23796);
and UO_1527 (O_1527,N_24189,N_22716);
and UO_1528 (O_1528,N_22145,N_23678);
or UO_1529 (O_1529,N_23288,N_24232);
or UO_1530 (O_1530,N_23371,N_23723);
xor UO_1531 (O_1531,N_24957,N_23979);
and UO_1532 (O_1532,N_23580,N_23045);
nand UO_1533 (O_1533,N_24907,N_24319);
nand UO_1534 (O_1534,N_22615,N_22639);
nor UO_1535 (O_1535,N_24776,N_24190);
or UO_1536 (O_1536,N_24840,N_24428);
or UO_1537 (O_1537,N_21880,N_22566);
or UO_1538 (O_1538,N_24247,N_22129);
xor UO_1539 (O_1539,N_22595,N_24656);
xnor UO_1540 (O_1540,N_24976,N_22396);
and UO_1541 (O_1541,N_24770,N_22529);
xor UO_1542 (O_1542,N_22245,N_22045);
or UO_1543 (O_1543,N_23123,N_24870);
nor UO_1544 (O_1544,N_22368,N_23059);
nand UO_1545 (O_1545,N_23138,N_22114);
nand UO_1546 (O_1546,N_22116,N_23911);
xor UO_1547 (O_1547,N_24712,N_23574);
xor UO_1548 (O_1548,N_22852,N_24080);
xor UO_1549 (O_1549,N_23944,N_23632);
or UO_1550 (O_1550,N_22945,N_22701);
and UO_1551 (O_1551,N_23392,N_23257);
nor UO_1552 (O_1552,N_23930,N_22037);
xor UO_1553 (O_1553,N_23328,N_22830);
or UO_1554 (O_1554,N_23864,N_22230);
and UO_1555 (O_1555,N_22795,N_21883);
and UO_1556 (O_1556,N_24568,N_21967);
nor UO_1557 (O_1557,N_22044,N_24482);
xor UO_1558 (O_1558,N_24802,N_22384);
nand UO_1559 (O_1559,N_23347,N_23729);
and UO_1560 (O_1560,N_24790,N_22355);
or UO_1561 (O_1561,N_24440,N_23354);
and UO_1562 (O_1562,N_22602,N_23782);
or UO_1563 (O_1563,N_23462,N_23090);
nor UO_1564 (O_1564,N_24675,N_24790);
and UO_1565 (O_1565,N_24285,N_24326);
and UO_1566 (O_1566,N_21944,N_22404);
nand UO_1567 (O_1567,N_23656,N_23969);
and UO_1568 (O_1568,N_24345,N_24056);
nor UO_1569 (O_1569,N_23897,N_24402);
xor UO_1570 (O_1570,N_21891,N_24897);
and UO_1571 (O_1571,N_22677,N_22710);
and UO_1572 (O_1572,N_24246,N_21958);
or UO_1573 (O_1573,N_22660,N_24454);
xor UO_1574 (O_1574,N_23349,N_24733);
or UO_1575 (O_1575,N_24364,N_23507);
nand UO_1576 (O_1576,N_22254,N_24736);
xor UO_1577 (O_1577,N_23950,N_23411);
nor UO_1578 (O_1578,N_22486,N_22957);
xor UO_1579 (O_1579,N_23606,N_21946);
and UO_1580 (O_1580,N_24819,N_24653);
nand UO_1581 (O_1581,N_22274,N_23462);
nor UO_1582 (O_1582,N_24398,N_21967);
nor UO_1583 (O_1583,N_22892,N_24781);
xnor UO_1584 (O_1584,N_22189,N_23774);
nor UO_1585 (O_1585,N_22108,N_23582);
or UO_1586 (O_1586,N_23048,N_24938);
nand UO_1587 (O_1587,N_22697,N_22590);
nor UO_1588 (O_1588,N_22259,N_22021);
or UO_1589 (O_1589,N_23971,N_23988);
xnor UO_1590 (O_1590,N_22808,N_22254);
xnor UO_1591 (O_1591,N_23406,N_24793);
and UO_1592 (O_1592,N_22474,N_22055);
nand UO_1593 (O_1593,N_23597,N_22206);
and UO_1594 (O_1594,N_23428,N_22082);
xor UO_1595 (O_1595,N_23741,N_24388);
nand UO_1596 (O_1596,N_21953,N_22307);
and UO_1597 (O_1597,N_22080,N_23406);
nand UO_1598 (O_1598,N_23947,N_24240);
and UO_1599 (O_1599,N_24500,N_23641);
xnor UO_1600 (O_1600,N_23379,N_22364);
and UO_1601 (O_1601,N_22133,N_23867);
nand UO_1602 (O_1602,N_24844,N_22297);
xor UO_1603 (O_1603,N_24519,N_23924);
and UO_1604 (O_1604,N_22947,N_22659);
and UO_1605 (O_1605,N_23538,N_22445);
or UO_1606 (O_1606,N_23937,N_24605);
or UO_1607 (O_1607,N_23064,N_23589);
nor UO_1608 (O_1608,N_24107,N_24122);
xor UO_1609 (O_1609,N_22000,N_24230);
nor UO_1610 (O_1610,N_24845,N_22659);
nand UO_1611 (O_1611,N_22463,N_23524);
nand UO_1612 (O_1612,N_24302,N_23980);
and UO_1613 (O_1613,N_23275,N_22429);
nor UO_1614 (O_1614,N_22234,N_22014);
or UO_1615 (O_1615,N_21973,N_23972);
nor UO_1616 (O_1616,N_22041,N_23973);
or UO_1617 (O_1617,N_23995,N_23007);
and UO_1618 (O_1618,N_24633,N_23811);
nand UO_1619 (O_1619,N_22551,N_22051);
or UO_1620 (O_1620,N_24065,N_24840);
nor UO_1621 (O_1621,N_23067,N_24306);
nand UO_1622 (O_1622,N_24429,N_24953);
nand UO_1623 (O_1623,N_23320,N_22073);
or UO_1624 (O_1624,N_23102,N_23706);
xor UO_1625 (O_1625,N_23762,N_24194);
nand UO_1626 (O_1626,N_22099,N_24949);
and UO_1627 (O_1627,N_23732,N_22437);
xor UO_1628 (O_1628,N_22607,N_22957);
and UO_1629 (O_1629,N_23417,N_24916);
nand UO_1630 (O_1630,N_24432,N_23518);
and UO_1631 (O_1631,N_23955,N_24572);
and UO_1632 (O_1632,N_23587,N_24900);
and UO_1633 (O_1633,N_22103,N_23543);
and UO_1634 (O_1634,N_24163,N_24395);
xor UO_1635 (O_1635,N_23123,N_24251);
nor UO_1636 (O_1636,N_23424,N_22019);
nand UO_1637 (O_1637,N_22644,N_22223);
or UO_1638 (O_1638,N_22828,N_22083);
or UO_1639 (O_1639,N_24942,N_24908);
xnor UO_1640 (O_1640,N_23107,N_23569);
nand UO_1641 (O_1641,N_24728,N_23285);
and UO_1642 (O_1642,N_24452,N_22736);
and UO_1643 (O_1643,N_24009,N_23063);
and UO_1644 (O_1644,N_22360,N_23298);
and UO_1645 (O_1645,N_23808,N_24031);
or UO_1646 (O_1646,N_22007,N_22539);
nand UO_1647 (O_1647,N_22170,N_24594);
or UO_1648 (O_1648,N_22840,N_23888);
nand UO_1649 (O_1649,N_23214,N_24846);
xnor UO_1650 (O_1650,N_23589,N_24097);
nor UO_1651 (O_1651,N_22951,N_23555);
and UO_1652 (O_1652,N_23561,N_22730);
nand UO_1653 (O_1653,N_24165,N_23188);
nor UO_1654 (O_1654,N_22504,N_24727);
nor UO_1655 (O_1655,N_23332,N_22610);
or UO_1656 (O_1656,N_22756,N_23117);
and UO_1657 (O_1657,N_22473,N_22396);
or UO_1658 (O_1658,N_23776,N_22641);
xor UO_1659 (O_1659,N_24076,N_24721);
and UO_1660 (O_1660,N_22058,N_23764);
xor UO_1661 (O_1661,N_24447,N_24022);
nor UO_1662 (O_1662,N_22289,N_23831);
and UO_1663 (O_1663,N_24721,N_23653);
and UO_1664 (O_1664,N_24351,N_24311);
nand UO_1665 (O_1665,N_23088,N_24024);
nor UO_1666 (O_1666,N_22252,N_22210);
nand UO_1667 (O_1667,N_24904,N_24964);
and UO_1668 (O_1668,N_23990,N_24217);
or UO_1669 (O_1669,N_22275,N_23111);
and UO_1670 (O_1670,N_22499,N_22843);
and UO_1671 (O_1671,N_22195,N_22135);
nand UO_1672 (O_1672,N_23099,N_23009);
nand UO_1673 (O_1673,N_23196,N_22597);
or UO_1674 (O_1674,N_22884,N_24977);
or UO_1675 (O_1675,N_22826,N_23916);
nand UO_1676 (O_1676,N_24590,N_24708);
xor UO_1677 (O_1677,N_24265,N_22443);
or UO_1678 (O_1678,N_24155,N_24581);
xor UO_1679 (O_1679,N_22669,N_23225);
xnor UO_1680 (O_1680,N_22713,N_23097);
and UO_1681 (O_1681,N_23959,N_22002);
and UO_1682 (O_1682,N_24914,N_24196);
or UO_1683 (O_1683,N_22480,N_22884);
or UO_1684 (O_1684,N_24646,N_24808);
or UO_1685 (O_1685,N_23554,N_24007);
and UO_1686 (O_1686,N_24954,N_24012);
xor UO_1687 (O_1687,N_23685,N_22626);
or UO_1688 (O_1688,N_22911,N_22103);
nand UO_1689 (O_1689,N_23126,N_23097);
nand UO_1690 (O_1690,N_24087,N_23449);
and UO_1691 (O_1691,N_23247,N_24600);
and UO_1692 (O_1692,N_24168,N_22286);
xnor UO_1693 (O_1693,N_21943,N_24276);
nand UO_1694 (O_1694,N_24505,N_22137);
nor UO_1695 (O_1695,N_24852,N_24693);
and UO_1696 (O_1696,N_24291,N_23322);
nand UO_1697 (O_1697,N_24186,N_23299);
and UO_1698 (O_1698,N_22724,N_23065);
nor UO_1699 (O_1699,N_22425,N_24795);
nor UO_1700 (O_1700,N_22369,N_24175);
xor UO_1701 (O_1701,N_24070,N_22645);
or UO_1702 (O_1702,N_23627,N_23618);
nand UO_1703 (O_1703,N_22479,N_22449);
and UO_1704 (O_1704,N_23855,N_22199);
xnor UO_1705 (O_1705,N_24419,N_23424);
xor UO_1706 (O_1706,N_21935,N_22529);
and UO_1707 (O_1707,N_24659,N_22237);
or UO_1708 (O_1708,N_22819,N_23888);
xnor UO_1709 (O_1709,N_23778,N_24404);
nand UO_1710 (O_1710,N_24287,N_23587);
nand UO_1711 (O_1711,N_24134,N_24106);
or UO_1712 (O_1712,N_22343,N_22427);
and UO_1713 (O_1713,N_23839,N_23730);
xnor UO_1714 (O_1714,N_24748,N_22477);
or UO_1715 (O_1715,N_24434,N_24758);
nor UO_1716 (O_1716,N_23114,N_24415);
or UO_1717 (O_1717,N_22301,N_24474);
or UO_1718 (O_1718,N_24943,N_24120);
nand UO_1719 (O_1719,N_22937,N_24507);
and UO_1720 (O_1720,N_23365,N_22409);
or UO_1721 (O_1721,N_22807,N_23231);
nand UO_1722 (O_1722,N_21975,N_21962);
and UO_1723 (O_1723,N_23227,N_24965);
or UO_1724 (O_1724,N_24854,N_24559);
or UO_1725 (O_1725,N_23062,N_23691);
xnor UO_1726 (O_1726,N_23395,N_21982);
or UO_1727 (O_1727,N_21887,N_24814);
or UO_1728 (O_1728,N_22316,N_22383);
or UO_1729 (O_1729,N_24143,N_22506);
xor UO_1730 (O_1730,N_23090,N_21966);
or UO_1731 (O_1731,N_22031,N_23377);
or UO_1732 (O_1732,N_24056,N_24352);
nand UO_1733 (O_1733,N_23683,N_24660);
xnor UO_1734 (O_1734,N_24436,N_22962);
and UO_1735 (O_1735,N_21922,N_24095);
nand UO_1736 (O_1736,N_23711,N_24215);
nor UO_1737 (O_1737,N_23110,N_22163);
nor UO_1738 (O_1738,N_22907,N_23007);
nor UO_1739 (O_1739,N_22908,N_24559);
and UO_1740 (O_1740,N_22477,N_23634);
nand UO_1741 (O_1741,N_24955,N_22555);
nand UO_1742 (O_1742,N_24771,N_22621);
nand UO_1743 (O_1743,N_24980,N_22880);
nor UO_1744 (O_1744,N_23591,N_24653);
xor UO_1745 (O_1745,N_21986,N_23400);
xor UO_1746 (O_1746,N_23924,N_23698);
nand UO_1747 (O_1747,N_22516,N_23114);
nor UO_1748 (O_1748,N_22503,N_22194);
nand UO_1749 (O_1749,N_24636,N_23354);
xnor UO_1750 (O_1750,N_23058,N_23777);
or UO_1751 (O_1751,N_23490,N_23955);
nor UO_1752 (O_1752,N_22111,N_22607);
nor UO_1753 (O_1753,N_23612,N_23771);
nor UO_1754 (O_1754,N_23494,N_23613);
or UO_1755 (O_1755,N_22420,N_24982);
nand UO_1756 (O_1756,N_24295,N_22750);
and UO_1757 (O_1757,N_22370,N_24939);
and UO_1758 (O_1758,N_21882,N_22520);
nand UO_1759 (O_1759,N_22129,N_24813);
nor UO_1760 (O_1760,N_24632,N_23809);
and UO_1761 (O_1761,N_23447,N_24072);
or UO_1762 (O_1762,N_24880,N_24521);
xnor UO_1763 (O_1763,N_22302,N_24751);
nand UO_1764 (O_1764,N_23717,N_22812);
xor UO_1765 (O_1765,N_21979,N_22147);
xor UO_1766 (O_1766,N_22299,N_24160);
nor UO_1767 (O_1767,N_24438,N_22988);
xnor UO_1768 (O_1768,N_24820,N_24384);
nor UO_1769 (O_1769,N_24695,N_22038);
nand UO_1770 (O_1770,N_22077,N_24545);
or UO_1771 (O_1771,N_22544,N_23427);
or UO_1772 (O_1772,N_24160,N_23899);
or UO_1773 (O_1773,N_23383,N_23710);
nand UO_1774 (O_1774,N_23954,N_22697);
nor UO_1775 (O_1775,N_24300,N_22578);
and UO_1776 (O_1776,N_23465,N_23175);
nor UO_1777 (O_1777,N_22546,N_22794);
or UO_1778 (O_1778,N_23695,N_24564);
nor UO_1779 (O_1779,N_23688,N_22722);
nand UO_1780 (O_1780,N_22844,N_24839);
nand UO_1781 (O_1781,N_22610,N_24648);
or UO_1782 (O_1782,N_24244,N_24047);
nor UO_1783 (O_1783,N_22947,N_22630);
nor UO_1784 (O_1784,N_22383,N_24261);
and UO_1785 (O_1785,N_23505,N_23712);
xnor UO_1786 (O_1786,N_22819,N_24061);
or UO_1787 (O_1787,N_22462,N_24101);
xnor UO_1788 (O_1788,N_24083,N_23242);
nor UO_1789 (O_1789,N_24587,N_22929);
nor UO_1790 (O_1790,N_24968,N_23046);
nand UO_1791 (O_1791,N_22965,N_24795);
nor UO_1792 (O_1792,N_23998,N_22149);
xor UO_1793 (O_1793,N_22977,N_24692);
or UO_1794 (O_1794,N_22054,N_23736);
or UO_1795 (O_1795,N_24185,N_23420);
nor UO_1796 (O_1796,N_24873,N_23843);
and UO_1797 (O_1797,N_24667,N_21885);
and UO_1798 (O_1798,N_22904,N_22743);
xnor UO_1799 (O_1799,N_22326,N_24873);
and UO_1800 (O_1800,N_24741,N_22923);
or UO_1801 (O_1801,N_22475,N_23112);
xor UO_1802 (O_1802,N_22079,N_23193);
or UO_1803 (O_1803,N_24790,N_23707);
nand UO_1804 (O_1804,N_24746,N_24442);
nand UO_1805 (O_1805,N_22170,N_22607);
and UO_1806 (O_1806,N_24483,N_22849);
and UO_1807 (O_1807,N_24028,N_24958);
nand UO_1808 (O_1808,N_23146,N_23081);
and UO_1809 (O_1809,N_24464,N_22957);
or UO_1810 (O_1810,N_22514,N_22304);
xor UO_1811 (O_1811,N_24157,N_22901);
or UO_1812 (O_1812,N_23016,N_23240);
nand UO_1813 (O_1813,N_22034,N_23967);
and UO_1814 (O_1814,N_22036,N_23486);
or UO_1815 (O_1815,N_24587,N_21994);
nand UO_1816 (O_1816,N_23120,N_24723);
nor UO_1817 (O_1817,N_22506,N_22261);
and UO_1818 (O_1818,N_23304,N_23947);
nand UO_1819 (O_1819,N_23643,N_23309);
nand UO_1820 (O_1820,N_24589,N_24912);
xor UO_1821 (O_1821,N_23151,N_24141);
nor UO_1822 (O_1822,N_23203,N_22705);
nand UO_1823 (O_1823,N_24052,N_22597);
or UO_1824 (O_1824,N_22404,N_22156);
xnor UO_1825 (O_1825,N_24251,N_22882);
and UO_1826 (O_1826,N_22615,N_24644);
xnor UO_1827 (O_1827,N_23197,N_22713);
and UO_1828 (O_1828,N_22489,N_24610);
nor UO_1829 (O_1829,N_23028,N_23177);
xnor UO_1830 (O_1830,N_22977,N_22404);
xor UO_1831 (O_1831,N_24332,N_24062);
xor UO_1832 (O_1832,N_23630,N_24226);
nor UO_1833 (O_1833,N_24274,N_22879);
nor UO_1834 (O_1834,N_22367,N_22423);
nand UO_1835 (O_1835,N_23474,N_22869);
and UO_1836 (O_1836,N_24807,N_24032);
nand UO_1837 (O_1837,N_24225,N_24397);
nand UO_1838 (O_1838,N_22895,N_23404);
or UO_1839 (O_1839,N_22248,N_22169);
or UO_1840 (O_1840,N_23401,N_24107);
xnor UO_1841 (O_1841,N_22784,N_22730);
nand UO_1842 (O_1842,N_22006,N_23160);
or UO_1843 (O_1843,N_22135,N_22892);
nand UO_1844 (O_1844,N_22360,N_23168);
or UO_1845 (O_1845,N_24690,N_22988);
or UO_1846 (O_1846,N_22161,N_23436);
nand UO_1847 (O_1847,N_21981,N_22007);
xor UO_1848 (O_1848,N_21992,N_24644);
nor UO_1849 (O_1849,N_23530,N_22773);
or UO_1850 (O_1850,N_22371,N_23043);
and UO_1851 (O_1851,N_22736,N_22652);
or UO_1852 (O_1852,N_23319,N_23027);
or UO_1853 (O_1853,N_22664,N_23172);
or UO_1854 (O_1854,N_24615,N_23573);
nor UO_1855 (O_1855,N_22281,N_22504);
xnor UO_1856 (O_1856,N_24242,N_22683);
or UO_1857 (O_1857,N_24313,N_24778);
or UO_1858 (O_1858,N_23727,N_21946);
xor UO_1859 (O_1859,N_21974,N_23610);
and UO_1860 (O_1860,N_23375,N_22002);
nor UO_1861 (O_1861,N_24143,N_21913);
and UO_1862 (O_1862,N_22482,N_22123);
nor UO_1863 (O_1863,N_23197,N_22353);
nor UO_1864 (O_1864,N_24682,N_21917);
nor UO_1865 (O_1865,N_23366,N_24991);
nor UO_1866 (O_1866,N_24086,N_23315);
nor UO_1867 (O_1867,N_24737,N_21991);
nor UO_1868 (O_1868,N_24398,N_22711);
or UO_1869 (O_1869,N_22805,N_22428);
and UO_1870 (O_1870,N_24313,N_24231);
xnor UO_1871 (O_1871,N_24546,N_24315);
and UO_1872 (O_1872,N_23063,N_22930);
nand UO_1873 (O_1873,N_22381,N_24650);
xnor UO_1874 (O_1874,N_22899,N_23581);
and UO_1875 (O_1875,N_22288,N_24068);
xor UO_1876 (O_1876,N_23062,N_22254);
or UO_1877 (O_1877,N_23560,N_22662);
xor UO_1878 (O_1878,N_22949,N_24077);
and UO_1879 (O_1879,N_24666,N_24974);
xor UO_1880 (O_1880,N_22918,N_23141);
or UO_1881 (O_1881,N_23373,N_24369);
and UO_1882 (O_1882,N_24420,N_22798);
or UO_1883 (O_1883,N_24506,N_23737);
nor UO_1884 (O_1884,N_23982,N_23455);
and UO_1885 (O_1885,N_23378,N_24634);
nor UO_1886 (O_1886,N_22252,N_24399);
xor UO_1887 (O_1887,N_22007,N_22865);
or UO_1888 (O_1888,N_22327,N_23364);
nand UO_1889 (O_1889,N_22841,N_24794);
and UO_1890 (O_1890,N_23451,N_24415);
and UO_1891 (O_1891,N_22891,N_23750);
and UO_1892 (O_1892,N_23928,N_23020);
xor UO_1893 (O_1893,N_23517,N_24837);
and UO_1894 (O_1894,N_23099,N_22698);
nand UO_1895 (O_1895,N_23133,N_23641);
xnor UO_1896 (O_1896,N_24862,N_23592);
and UO_1897 (O_1897,N_24009,N_22438);
nor UO_1898 (O_1898,N_22341,N_24923);
xnor UO_1899 (O_1899,N_24383,N_24070);
nand UO_1900 (O_1900,N_22025,N_22929);
xnor UO_1901 (O_1901,N_24608,N_23141);
xor UO_1902 (O_1902,N_24825,N_24342);
or UO_1903 (O_1903,N_24006,N_24039);
nor UO_1904 (O_1904,N_22613,N_24623);
and UO_1905 (O_1905,N_24740,N_24834);
xnor UO_1906 (O_1906,N_24164,N_23231);
and UO_1907 (O_1907,N_23339,N_22687);
xor UO_1908 (O_1908,N_24148,N_24613);
xor UO_1909 (O_1909,N_24605,N_22734);
nand UO_1910 (O_1910,N_22015,N_22882);
nand UO_1911 (O_1911,N_23594,N_24042);
nand UO_1912 (O_1912,N_23175,N_23244);
nand UO_1913 (O_1913,N_24983,N_21927);
nor UO_1914 (O_1914,N_23519,N_24224);
and UO_1915 (O_1915,N_22215,N_23350);
nor UO_1916 (O_1916,N_22676,N_22632);
nand UO_1917 (O_1917,N_24616,N_23034);
nor UO_1918 (O_1918,N_23137,N_22838);
xnor UO_1919 (O_1919,N_22740,N_24406);
and UO_1920 (O_1920,N_24442,N_22346);
and UO_1921 (O_1921,N_22729,N_24442);
nand UO_1922 (O_1922,N_22585,N_24275);
and UO_1923 (O_1923,N_21899,N_22336);
nor UO_1924 (O_1924,N_24792,N_23745);
or UO_1925 (O_1925,N_24936,N_24414);
and UO_1926 (O_1926,N_21978,N_24792);
xnor UO_1927 (O_1927,N_24078,N_23078);
and UO_1928 (O_1928,N_24944,N_22624);
nor UO_1929 (O_1929,N_24169,N_22760);
and UO_1930 (O_1930,N_24820,N_23351);
or UO_1931 (O_1931,N_23301,N_23033);
or UO_1932 (O_1932,N_22655,N_22795);
and UO_1933 (O_1933,N_21933,N_24743);
nand UO_1934 (O_1934,N_23514,N_24500);
and UO_1935 (O_1935,N_23602,N_22834);
nor UO_1936 (O_1936,N_24222,N_22475);
nand UO_1937 (O_1937,N_22081,N_22446);
nand UO_1938 (O_1938,N_24882,N_24983);
or UO_1939 (O_1939,N_23311,N_22403);
xor UO_1940 (O_1940,N_24691,N_21951);
nor UO_1941 (O_1941,N_24134,N_24434);
or UO_1942 (O_1942,N_22058,N_22322);
and UO_1943 (O_1943,N_24192,N_23099);
nor UO_1944 (O_1944,N_24472,N_23232);
nand UO_1945 (O_1945,N_23523,N_22005);
or UO_1946 (O_1946,N_22121,N_24660);
xor UO_1947 (O_1947,N_24381,N_24397);
nor UO_1948 (O_1948,N_23239,N_22213);
nand UO_1949 (O_1949,N_23544,N_23064);
or UO_1950 (O_1950,N_22377,N_24795);
nor UO_1951 (O_1951,N_21881,N_24560);
and UO_1952 (O_1952,N_24510,N_24498);
nand UO_1953 (O_1953,N_24329,N_22112);
nand UO_1954 (O_1954,N_23014,N_23886);
xnor UO_1955 (O_1955,N_21901,N_24006);
nand UO_1956 (O_1956,N_21947,N_24960);
nand UO_1957 (O_1957,N_22417,N_23419);
and UO_1958 (O_1958,N_22447,N_22922);
and UO_1959 (O_1959,N_23375,N_24280);
or UO_1960 (O_1960,N_23738,N_24909);
xor UO_1961 (O_1961,N_24672,N_23095);
or UO_1962 (O_1962,N_24966,N_24372);
xor UO_1963 (O_1963,N_23455,N_22985);
or UO_1964 (O_1964,N_24626,N_24497);
xnor UO_1965 (O_1965,N_24877,N_23935);
or UO_1966 (O_1966,N_22676,N_23749);
nor UO_1967 (O_1967,N_22704,N_24743);
nor UO_1968 (O_1968,N_23119,N_23031);
nor UO_1969 (O_1969,N_23109,N_24117);
nand UO_1970 (O_1970,N_23174,N_24836);
nand UO_1971 (O_1971,N_24290,N_23004);
or UO_1972 (O_1972,N_22822,N_22815);
or UO_1973 (O_1973,N_23028,N_23653);
and UO_1974 (O_1974,N_24656,N_22118);
nor UO_1975 (O_1975,N_23989,N_23194);
and UO_1976 (O_1976,N_23310,N_24567);
xnor UO_1977 (O_1977,N_22441,N_23363);
xor UO_1978 (O_1978,N_23171,N_22897);
or UO_1979 (O_1979,N_24021,N_23725);
nand UO_1980 (O_1980,N_24204,N_21933);
nor UO_1981 (O_1981,N_23677,N_23037);
xor UO_1982 (O_1982,N_24999,N_22133);
xor UO_1983 (O_1983,N_23987,N_23324);
nand UO_1984 (O_1984,N_22464,N_22059);
or UO_1985 (O_1985,N_22495,N_23284);
xnor UO_1986 (O_1986,N_22579,N_23642);
xor UO_1987 (O_1987,N_22492,N_23329);
and UO_1988 (O_1988,N_24090,N_23040);
or UO_1989 (O_1989,N_22093,N_24001);
nor UO_1990 (O_1990,N_22897,N_24767);
or UO_1991 (O_1991,N_24714,N_24405);
xor UO_1992 (O_1992,N_23683,N_21909);
nand UO_1993 (O_1993,N_23817,N_24335);
xor UO_1994 (O_1994,N_23705,N_24863);
xor UO_1995 (O_1995,N_24595,N_23460);
and UO_1996 (O_1996,N_23250,N_22260);
nand UO_1997 (O_1997,N_22087,N_22896);
nor UO_1998 (O_1998,N_23378,N_22207);
or UO_1999 (O_1999,N_22721,N_23328);
xor UO_2000 (O_2000,N_22084,N_23419);
and UO_2001 (O_2001,N_22015,N_24018);
nor UO_2002 (O_2002,N_21957,N_22496);
or UO_2003 (O_2003,N_23066,N_23007);
xor UO_2004 (O_2004,N_21882,N_23709);
or UO_2005 (O_2005,N_23751,N_22443);
nor UO_2006 (O_2006,N_22004,N_24601);
xnor UO_2007 (O_2007,N_22642,N_22649);
nor UO_2008 (O_2008,N_22990,N_23959);
or UO_2009 (O_2009,N_22637,N_24479);
nand UO_2010 (O_2010,N_22521,N_22409);
or UO_2011 (O_2011,N_22987,N_23064);
nand UO_2012 (O_2012,N_23439,N_24720);
and UO_2013 (O_2013,N_24527,N_24301);
nand UO_2014 (O_2014,N_23360,N_23767);
xor UO_2015 (O_2015,N_21875,N_23921);
nor UO_2016 (O_2016,N_22271,N_22645);
nor UO_2017 (O_2017,N_24097,N_22184);
and UO_2018 (O_2018,N_23911,N_22443);
or UO_2019 (O_2019,N_24083,N_23142);
nand UO_2020 (O_2020,N_24751,N_22649);
nand UO_2021 (O_2021,N_22121,N_21885);
xor UO_2022 (O_2022,N_22598,N_23910);
xor UO_2023 (O_2023,N_24000,N_23756);
and UO_2024 (O_2024,N_21881,N_24504);
or UO_2025 (O_2025,N_24142,N_23028);
nor UO_2026 (O_2026,N_22153,N_23450);
or UO_2027 (O_2027,N_22049,N_23576);
nand UO_2028 (O_2028,N_24619,N_24107);
nand UO_2029 (O_2029,N_22977,N_24056);
nor UO_2030 (O_2030,N_22503,N_23344);
and UO_2031 (O_2031,N_23473,N_22470);
xor UO_2032 (O_2032,N_23485,N_24564);
xnor UO_2033 (O_2033,N_23320,N_24172);
and UO_2034 (O_2034,N_24455,N_22652);
nand UO_2035 (O_2035,N_23486,N_24095);
and UO_2036 (O_2036,N_24398,N_22114);
nand UO_2037 (O_2037,N_23112,N_24227);
or UO_2038 (O_2038,N_22260,N_24458);
nor UO_2039 (O_2039,N_24082,N_23556);
nor UO_2040 (O_2040,N_23061,N_22403);
nand UO_2041 (O_2041,N_24596,N_22964);
xor UO_2042 (O_2042,N_23508,N_24393);
and UO_2043 (O_2043,N_23247,N_22464);
nand UO_2044 (O_2044,N_24877,N_23132);
or UO_2045 (O_2045,N_24453,N_22111);
nand UO_2046 (O_2046,N_21934,N_22083);
nand UO_2047 (O_2047,N_22837,N_22393);
nand UO_2048 (O_2048,N_21995,N_22967);
and UO_2049 (O_2049,N_24698,N_23333);
and UO_2050 (O_2050,N_23021,N_23460);
or UO_2051 (O_2051,N_24244,N_24413);
xnor UO_2052 (O_2052,N_24355,N_23998);
nor UO_2053 (O_2053,N_24320,N_24552);
and UO_2054 (O_2054,N_22879,N_22542);
nand UO_2055 (O_2055,N_22911,N_22061);
and UO_2056 (O_2056,N_24602,N_24090);
and UO_2057 (O_2057,N_22014,N_22151);
nand UO_2058 (O_2058,N_22370,N_22300);
and UO_2059 (O_2059,N_24158,N_22400);
and UO_2060 (O_2060,N_24676,N_22392);
xor UO_2061 (O_2061,N_22419,N_22179);
and UO_2062 (O_2062,N_24903,N_23548);
and UO_2063 (O_2063,N_23691,N_22577);
xor UO_2064 (O_2064,N_23290,N_21884);
xnor UO_2065 (O_2065,N_22192,N_22200);
or UO_2066 (O_2066,N_22885,N_23558);
or UO_2067 (O_2067,N_23557,N_22752);
and UO_2068 (O_2068,N_22333,N_24810);
or UO_2069 (O_2069,N_24192,N_22722);
xor UO_2070 (O_2070,N_21994,N_21883);
nor UO_2071 (O_2071,N_23751,N_23091);
and UO_2072 (O_2072,N_23227,N_23898);
and UO_2073 (O_2073,N_24835,N_23489);
xnor UO_2074 (O_2074,N_24792,N_22881);
xnor UO_2075 (O_2075,N_23909,N_22641);
nand UO_2076 (O_2076,N_24092,N_24299);
and UO_2077 (O_2077,N_23933,N_23322);
or UO_2078 (O_2078,N_24018,N_24681);
or UO_2079 (O_2079,N_23521,N_22713);
nor UO_2080 (O_2080,N_24383,N_24477);
nor UO_2081 (O_2081,N_24945,N_24410);
and UO_2082 (O_2082,N_24509,N_22389);
nand UO_2083 (O_2083,N_24399,N_23207);
xor UO_2084 (O_2084,N_22088,N_23571);
xnor UO_2085 (O_2085,N_22611,N_24804);
or UO_2086 (O_2086,N_24056,N_24162);
and UO_2087 (O_2087,N_22901,N_23486);
xnor UO_2088 (O_2088,N_24880,N_24742);
or UO_2089 (O_2089,N_24598,N_23553);
or UO_2090 (O_2090,N_24450,N_22111);
and UO_2091 (O_2091,N_22692,N_24557);
nand UO_2092 (O_2092,N_22057,N_24625);
or UO_2093 (O_2093,N_23280,N_22352);
nand UO_2094 (O_2094,N_22114,N_23543);
xor UO_2095 (O_2095,N_22005,N_24835);
and UO_2096 (O_2096,N_22114,N_22466);
or UO_2097 (O_2097,N_24665,N_22622);
and UO_2098 (O_2098,N_21948,N_24449);
xnor UO_2099 (O_2099,N_21992,N_24420);
nand UO_2100 (O_2100,N_22701,N_23603);
xnor UO_2101 (O_2101,N_24907,N_24390);
and UO_2102 (O_2102,N_23738,N_22639);
xor UO_2103 (O_2103,N_23955,N_23684);
nor UO_2104 (O_2104,N_22972,N_22038);
and UO_2105 (O_2105,N_24962,N_22689);
xor UO_2106 (O_2106,N_23593,N_22318);
and UO_2107 (O_2107,N_21926,N_24761);
or UO_2108 (O_2108,N_22653,N_22798);
xnor UO_2109 (O_2109,N_22581,N_23561);
nor UO_2110 (O_2110,N_23818,N_22943);
or UO_2111 (O_2111,N_22462,N_24927);
or UO_2112 (O_2112,N_24312,N_22589);
xnor UO_2113 (O_2113,N_22367,N_21885);
nand UO_2114 (O_2114,N_23604,N_23339);
and UO_2115 (O_2115,N_23997,N_24607);
nand UO_2116 (O_2116,N_24041,N_24171);
nand UO_2117 (O_2117,N_24328,N_23757);
nor UO_2118 (O_2118,N_24932,N_24233);
xor UO_2119 (O_2119,N_23259,N_24518);
nor UO_2120 (O_2120,N_23451,N_23962);
xor UO_2121 (O_2121,N_23593,N_24997);
or UO_2122 (O_2122,N_23184,N_23250);
and UO_2123 (O_2123,N_22031,N_22830);
nor UO_2124 (O_2124,N_22442,N_24257);
nor UO_2125 (O_2125,N_22501,N_24749);
xor UO_2126 (O_2126,N_22392,N_22774);
or UO_2127 (O_2127,N_23878,N_24201);
or UO_2128 (O_2128,N_24949,N_22314);
nand UO_2129 (O_2129,N_23344,N_24776);
nand UO_2130 (O_2130,N_24280,N_22173);
nand UO_2131 (O_2131,N_23625,N_23054);
or UO_2132 (O_2132,N_24004,N_23522);
xor UO_2133 (O_2133,N_23310,N_22050);
and UO_2134 (O_2134,N_22292,N_22524);
and UO_2135 (O_2135,N_22631,N_24092);
nor UO_2136 (O_2136,N_23531,N_22844);
nand UO_2137 (O_2137,N_24602,N_24684);
xor UO_2138 (O_2138,N_23752,N_22758);
nor UO_2139 (O_2139,N_22813,N_21989);
and UO_2140 (O_2140,N_24897,N_23496);
nand UO_2141 (O_2141,N_23849,N_23364);
xor UO_2142 (O_2142,N_23201,N_22326);
nor UO_2143 (O_2143,N_23042,N_21883);
xor UO_2144 (O_2144,N_23766,N_23817);
nand UO_2145 (O_2145,N_22512,N_24708);
xnor UO_2146 (O_2146,N_22604,N_22071);
or UO_2147 (O_2147,N_23019,N_24573);
or UO_2148 (O_2148,N_24675,N_22190);
xor UO_2149 (O_2149,N_22024,N_24255);
nand UO_2150 (O_2150,N_24080,N_23490);
nand UO_2151 (O_2151,N_24317,N_24354);
or UO_2152 (O_2152,N_22934,N_24409);
or UO_2153 (O_2153,N_22704,N_24161);
nand UO_2154 (O_2154,N_24380,N_23415);
nor UO_2155 (O_2155,N_23532,N_23088);
or UO_2156 (O_2156,N_23110,N_23355);
and UO_2157 (O_2157,N_24411,N_24264);
xor UO_2158 (O_2158,N_24884,N_23796);
xor UO_2159 (O_2159,N_23793,N_23881);
xnor UO_2160 (O_2160,N_24276,N_22700);
and UO_2161 (O_2161,N_22654,N_23294);
and UO_2162 (O_2162,N_22667,N_23869);
nor UO_2163 (O_2163,N_22233,N_23579);
nor UO_2164 (O_2164,N_23548,N_23964);
nor UO_2165 (O_2165,N_24567,N_23420);
xnor UO_2166 (O_2166,N_23510,N_23425);
nand UO_2167 (O_2167,N_24698,N_22201);
or UO_2168 (O_2168,N_21969,N_24763);
xor UO_2169 (O_2169,N_23794,N_24326);
and UO_2170 (O_2170,N_22909,N_22754);
nor UO_2171 (O_2171,N_24765,N_22405);
or UO_2172 (O_2172,N_24239,N_24016);
and UO_2173 (O_2173,N_23746,N_23502);
nand UO_2174 (O_2174,N_24694,N_23275);
and UO_2175 (O_2175,N_22715,N_23684);
nand UO_2176 (O_2176,N_21884,N_22697);
nand UO_2177 (O_2177,N_24946,N_23252);
nand UO_2178 (O_2178,N_23622,N_22640);
nand UO_2179 (O_2179,N_22228,N_24035);
nor UO_2180 (O_2180,N_23024,N_24435);
xnor UO_2181 (O_2181,N_22740,N_23458);
nor UO_2182 (O_2182,N_24902,N_22109);
nor UO_2183 (O_2183,N_22046,N_23484);
and UO_2184 (O_2184,N_24021,N_23428);
nand UO_2185 (O_2185,N_24014,N_24611);
nor UO_2186 (O_2186,N_23827,N_22873);
or UO_2187 (O_2187,N_24662,N_22262);
and UO_2188 (O_2188,N_24643,N_22604);
nand UO_2189 (O_2189,N_23277,N_22235);
nand UO_2190 (O_2190,N_22406,N_22894);
nand UO_2191 (O_2191,N_22773,N_23673);
and UO_2192 (O_2192,N_21979,N_24530);
or UO_2193 (O_2193,N_23584,N_24114);
nand UO_2194 (O_2194,N_24707,N_22347);
nand UO_2195 (O_2195,N_24470,N_22590);
nor UO_2196 (O_2196,N_24842,N_23954);
xnor UO_2197 (O_2197,N_23972,N_24310);
xor UO_2198 (O_2198,N_24951,N_22153);
and UO_2199 (O_2199,N_23328,N_23317);
nor UO_2200 (O_2200,N_24829,N_24345);
nand UO_2201 (O_2201,N_24130,N_24869);
and UO_2202 (O_2202,N_22524,N_22186);
or UO_2203 (O_2203,N_23549,N_22674);
or UO_2204 (O_2204,N_24312,N_23164);
or UO_2205 (O_2205,N_23032,N_23924);
or UO_2206 (O_2206,N_22815,N_22644);
nor UO_2207 (O_2207,N_22050,N_24210);
nor UO_2208 (O_2208,N_22846,N_21935);
and UO_2209 (O_2209,N_22116,N_22089);
and UO_2210 (O_2210,N_22876,N_22971);
and UO_2211 (O_2211,N_22093,N_22795);
nand UO_2212 (O_2212,N_22890,N_23975);
xnor UO_2213 (O_2213,N_22432,N_24087);
or UO_2214 (O_2214,N_24101,N_21900);
xor UO_2215 (O_2215,N_21938,N_22229);
xnor UO_2216 (O_2216,N_22360,N_23931);
nand UO_2217 (O_2217,N_24893,N_24322);
and UO_2218 (O_2218,N_22796,N_24856);
xnor UO_2219 (O_2219,N_23260,N_23609);
xnor UO_2220 (O_2220,N_24528,N_24605);
nor UO_2221 (O_2221,N_22463,N_24000);
and UO_2222 (O_2222,N_22535,N_23123);
nand UO_2223 (O_2223,N_22260,N_24432);
nand UO_2224 (O_2224,N_24344,N_24316);
and UO_2225 (O_2225,N_24967,N_24766);
nor UO_2226 (O_2226,N_24036,N_23386);
nand UO_2227 (O_2227,N_24436,N_23163);
xor UO_2228 (O_2228,N_24384,N_22186);
and UO_2229 (O_2229,N_22188,N_23499);
and UO_2230 (O_2230,N_24298,N_22334);
xor UO_2231 (O_2231,N_24164,N_24242);
nand UO_2232 (O_2232,N_23406,N_23106);
and UO_2233 (O_2233,N_23549,N_24579);
xor UO_2234 (O_2234,N_22420,N_21881);
nor UO_2235 (O_2235,N_21879,N_21976);
nor UO_2236 (O_2236,N_23328,N_22491);
nor UO_2237 (O_2237,N_23935,N_24510);
and UO_2238 (O_2238,N_24161,N_24431);
or UO_2239 (O_2239,N_23367,N_23606);
and UO_2240 (O_2240,N_24616,N_23569);
nand UO_2241 (O_2241,N_24652,N_24002);
nor UO_2242 (O_2242,N_23915,N_22288);
and UO_2243 (O_2243,N_24541,N_22676);
nor UO_2244 (O_2244,N_22384,N_22753);
nand UO_2245 (O_2245,N_24277,N_23581);
xor UO_2246 (O_2246,N_24922,N_22532);
nand UO_2247 (O_2247,N_23496,N_24250);
nor UO_2248 (O_2248,N_22838,N_24461);
or UO_2249 (O_2249,N_21939,N_21987);
xnor UO_2250 (O_2250,N_23165,N_21923);
or UO_2251 (O_2251,N_23640,N_22164);
nor UO_2252 (O_2252,N_22785,N_24766);
and UO_2253 (O_2253,N_24828,N_22421);
and UO_2254 (O_2254,N_23450,N_23641);
xnor UO_2255 (O_2255,N_22250,N_22488);
xor UO_2256 (O_2256,N_22136,N_24849);
or UO_2257 (O_2257,N_24992,N_23001);
nor UO_2258 (O_2258,N_22234,N_22959);
nand UO_2259 (O_2259,N_24732,N_23308);
xnor UO_2260 (O_2260,N_23124,N_22674);
nand UO_2261 (O_2261,N_21895,N_23531);
or UO_2262 (O_2262,N_24075,N_24452);
nor UO_2263 (O_2263,N_24112,N_24419);
nor UO_2264 (O_2264,N_23762,N_22418);
and UO_2265 (O_2265,N_24534,N_23789);
or UO_2266 (O_2266,N_22941,N_22569);
nor UO_2267 (O_2267,N_24889,N_22765);
nand UO_2268 (O_2268,N_24765,N_23570);
nand UO_2269 (O_2269,N_23562,N_23525);
nor UO_2270 (O_2270,N_24445,N_22242);
nor UO_2271 (O_2271,N_23168,N_23306);
and UO_2272 (O_2272,N_24691,N_23912);
nor UO_2273 (O_2273,N_23030,N_24887);
nor UO_2274 (O_2274,N_24072,N_24163);
xnor UO_2275 (O_2275,N_21906,N_24700);
nor UO_2276 (O_2276,N_24000,N_23478);
xnor UO_2277 (O_2277,N_23543,N_22672);
xor UO_2278 (O_2278,N_22604,N_23460);
nor UO_2279 (O_2279,N_23459,N_24043);
nor UO_2280 (O_2280,N_22921,N_23512);
or UO_2281 (O_2281,N_22706,N_23094);
nand UO_2282 (O_2282,N_24284,N_22154);
xor UO_2283 (O_2283,N_23352,N_22155);
nand UO_2284 (O_2284,N_23684,N_22867);
xnor UO_2285 (O_2285,N_22425,N_22232);
nand UO_2286 (O_2286,N_24841,N_22895);
xnor UO_2287 (O_2287,N_24009,N_22826);
or UO_2288 (O_2288,N_24398,N_23028);
and UO_2289 (O_2289,N_23082,N_23408);
and UO_2290 (O_2290,N_23112,N_24003);
nor UO_2291 (O_2291,N_22139,N_24311);
and UO_2292 (O_2292,N_22647,N_21964);
and UO_2293 (O_2293,N_23240,N_21984);
nand UO_2294 (O_2294,N_22151,N_23312);
nor UO_2295 (O_2295,N_24872,N_22736);
or UO_2296 (O_2296,N_24455,N_24199);
and UO_2297 (O_2297,N_24861,N_23324);
nor UO_2298 (O_2298,N_22635,N_22055);
and UO_2299 (O_2299,N_22580,N_22413);
xor UO_2300 (O_2300,N_21992,N_22268);
xor UO_2301 (O_2301,N_22344,N_23919);
and UO_2302 (O_2302,N_24394,N_22299);
nor UO_2303 (O_2303,N_24641,N_24317);
nand UO_2304 (O_2304,N_23068,N_22653);
and UO_2305 (O_2305,N_23737,N_24540);
nor UO_2306 (O_2306,N_23541,N_22589);
xnor UO_2307 (O_2307,N_24100,N_22746);
and UO_2308 (O_2308,N_22115,N_22116);
nand UO_2309 (O_2309,N_23409,N_23682);
xor UO_2310 (O_2310,N_22685,N_23702);
xnor UO_2311 (O_2311,N_23971,N_23569);
nor UO_2312 (O_2312,N_22901,N_24751);
xor UO_2313 (O_2313,N_24642,N_23523);
and UO_2314 (O_2314,N_24398,N_22062);
xor UO_2315 (O_2315,N_24139,N_24400);
or UO_2316 (O_2316,N_24145,N_22825);
nor UO_2317 (O_2317,N_24291,N_22998);
or UO_2318 (O_2318,N_24232,N_24325);
xor UO_2319 (O_2319,N_23598,N_23217);
nand UO_2320 (O_2320,N_22510,N_24975);
and UO_2321 (O_2321,N_24483,N_23343);
or UO_2322 (O_2322,N_24980,N_24847);
and UO_2323 (O_2323,N_23518,N_22786);
xor UO_2324 (O_2324,N_21951,N_24052);
or UO_2325 (O_2325,N_23662,N_22138);
or UO_2326 (O_2326,N_22428,N_23449);
xnor UO_2327 (O_2327,N_23171,N_23491);
nand UO_2328 (O_2328,N_24427,N_21978);
xnor UO_2329 (O_2329,N_22650,N_23992);
nor UO_2330 (O_2330,N_21910,N_24078);
xor UO_2331 (O_2331,N_22906,N_24591);
nand UO_2332 (O_2332,N_23437,N_22208);
xnor UO_2333 (O_2333,N_23812,N_21955);
nor UO_2334 (O_2334,N_22425,N_22380);
or UO_2335 (O_2335,N_23914,N_23382);
and UO_2336 (O_2336,N_24566,N_22935);
and UO_2337 (O_2337,N_23912,N_22202);
xor UO_2338 (O_2338,N_22123,N_22715);
nand UO_2339 (O_2339,N_22724,N_23212);
nand UO_2340 (O_2340,N_22975,N_23544);
nor UO_2341 (O_2341,N_24894,N_22899);
xor UO_2342 (O_2342,N_24804,N_23980);
xnor UO_2343 (O_2343,N_22496,N_22746);
xor UO_2344 (O_2344,N_23448,N_23017);
xor UO_2345 (O_2345,N_24980,N_22408);
nor UO_2346 (O_2346,N_23142,N_22686);
nor UO_2347 (O_2347,N_23676,N_23891);
nor UO_2348 (O_2348,N_22538,N_24227);
xor UO_2349 (O_2349,N_24015,N_24905);
xor UO_2350 (O_2350,N_22688,N_22485);
xnor UO_2351 (O_2351,N_22353,N_24355);
and UO_2352 (O_2352,N_24264,N_24684);
nor UO_2353 (O_2353,N_22336,N_24747);
xor UO_2354 (O_2354,N_23307,N_21891);
nand UO_2355 (O_2355,N_24302,N_22858);
or UO_2356 (O_2356,N_22598,N_22691);
nor UO_2357 (O_2357,N_24384,N_22453);
nor UO_2358 (O_2358,N_22937,N_24637);
xnor UO_2359 (O_2359,N_22347,N_24133);
and UO_2360 (O_2360,N_22674,N_23288);
nor UO_2361 (O_2361,N_22201,N_23156);
xor UO_2362 (O_2362,N_23613,N_22288);
nand UO_2363 (O_2363,N_24000,N_22981);
nand UO_2364 (O_2364,N_22004,N_22168);
or UO_2365 (O_2365,N_24247,N_24121);
and UO_2366 (O_2366,N_24483,N_22756);
nand UO_2367 (O_2367,N_22787,N_22719);
and UO_2368 (O_2368,N_23343,N_22832);
or UO_2369 (O_2369,N_24659,N_22688);
and UO_2370 (O_2370,N_24984,N_22133);
and UO_2371 (O_2371,N_24729,N_24212);
nand UO_2372 (O_2372,N_23279,N_24575);
nand UO_2373 (O_2373,N_23860,N_24677);
xnor UO_2374 (O_2374,N_24639,N_24264);
or UO_2375 (O_2375,N_22788,N_24747);
nor UO_2376 (O_2376,N_23800,N_24726);
xnor UO_2377 (O_2377,N_23316,N_22163);
or UO_2378 (O_2378,N_22024,N_24206);
or UO_2379 (O_2379,N_24626,N_23804);
nor UO_2380 (O_2380,N_22851,N_23756);
xnor UO_2381 (O_2381,N_24966,N_24239);
xor UO_2382 (O_2382,N_23983,N_24737);
or UO_2383 (O_2383,N_22899,N_24903);
xnor UO_2384 (O_2384,N_22361,N_22752);
and UO_2385 (O_2385,N_23694,N_23169);
or UO_2386 (O_2386,N_21959,N_23561);
and UO_2387 (O_2387,N_22416,N_24992);
or UO_2388 (O_2388,N_22187,N_22144);
xnor UO_2389 (O_2389,N_24497,N_24070);
xor UO_2390 (O_2390,N_23570,N_24190);
nor UO_2391 (O_2391,N_22840,N_22306);
nand UO_2392 (O_2392,N_24585,N_24869);
nand UO_2393 (O_2393,N_24685,N_23730);
and UO_2394 (O_2394,N_22339,N_24049);
xnor UO_2395 (O_2395,N_23344,N_24036);
xor UO_2396 (O_2396,N_22903,N_22263);
nor UO_2397 (O_2397,N_23315,N_22243);
nor UO_2398 (O_2398,N_24318,N_23594);
nor UO_2399 (O_2399,N_22809,N_22660);
nand UO_2400 (O_2400,N_22612,N_22170);
and UO_2401 (O_2401,N_22880,N_23444);
nand UO_2402 (O_2402,N_22245,N_22655);
nor UO_2403 (O_2403,N_24176,N_23916);
nand UO_2404 (O_2404,N_24918,N_24594);
nand UO_2405 (O_2405,N_23173,N_24062);
xnor UO_2406 (O_2406,N_22585,N_22694);
or UO_2407 (O_2407,N_22620,N_23208);
xnor UO_2408 (O_2408,N_23910,N_24135);
nand UO_2409 (O_2409,N_24619,N_24497);
and UO_2410 (O_2410,N_22638,N_23510);
or UO_2411 (O_2411,N_22355,N_23764);
xor UO_2412 (O_2412,N_22403,N_22139);
nor UO_2413 (O_2413,N_24808,N_24401);
or UO_2414 (O_2414,N_23165,N_22871);
or UO_2415 (O_2415,N_24624,N_22033);
or UO_2416 (O_2416,N_23046,N_24561);
and UO_2417 (O_2417,N_24615,N_22925);
nand UO_2418 (O_2418,N_24482,N_22652);
nand UO_2419 (O_2419,N_22425,N_23473);
xnor UO_2420 (O_2420,N_22540,N_23234);
xnor UO_2421 (O_2421,N_22208,N_22528);
nor UO_2422 (O_2422,N_24410,N_22922);
nor UO_2423 (O_2423,N_24577,N_23920);
and UO_2424 (O_2424,N_24176,N_24637);
and UO_2425 (O_2425,N_22620,N_23625);
or UO_2426 (O_2426,N_23670,N_23609);
and UO_2427 (O_2427,N_22679,N_22058);
nor UO_2428 (O_2428,N_24444,N_22738);
and UO_2429 (O_2429,N_24396,N_23131);
nor UO_2430 (O_2430,N_22738,N_24788);
nor UO_2431 (O_2431,N_22295,N_23990);
nor UO_2432 (O_2432,N_22179,N_22246);
xor UO_2433 (O_2433,N_24655,N_23610);
xor UO_2434 (O_2434,N_22992,N_24214);
xor UO_2435 (O_2435,N_24230,N_23147);
and UO_2436 (O_2436,N_22319,N_24273);
and UO_2437 (O_2437,N_22013,N_24668);
nand UO_2438 (O_2438,N_23305,N_23482);
nand UO_2439 (O_2439,N_22676,N_22083);
nand UO_2440 (O_2440,N_23687,N_22493);
nand UO_2441 (O_2441,N_22978,N_23066);
xnor UO_2442 (O_2442,N_24270,N_21994);
xor UO_2443 (O_2443,N_24598,N_22528);
or UO_2444 (O_2444,N_24837,N_24221);
nor UO_2445 (O_2445,N_22495,N_23089);
xnor UO_2446 (O_2446,N_22580,N_23376);
nand UO_2447 (O_2447,N_24463,N_23423);
xnor UO_2448 (O_2448,N_22249,N_22053);
nor UO_2449 (O_2449,N_24505,N_24890);
nand UO_2450 (O_2450,N_23658,N_23712);
nor UO_2451 (O_2451,N_22334,N_23414);
xor UO_2452 (O_2452,N_22512,N_22030);
xnor UO_2453 (O_2453,N_22627,N_23551);
nor UO_2454 (O_2454,N_23234,N_24095);
xnor UO_2455 (O_2455,N_24397,N_24553);
xnor UO_2456 (O_2456,N_22224,N_23755);
xnor UO_2457 (O_2457,N_21897,N_24068);
nor UO_2458 (O_2458,N_24819,N_22772);
nor UO_2459 (O_2459,N_24029,N_21978);
or UO_2460 (O_2460,N_23646,N_24806);
and UO_2461 (O_2461,N_24015,N_24819);
or UO_2462 (O_2462,N_23841,N_23466);
and UO_2463 (O_2463,N_21876,N_24806);
nor UO_2464 (O_2464,N_22628,N_23907);
nor UO_2465 (O_2465,N_24488,N_22774);
xor UO_2466 (O_2466,N_24837,N_21925);
or UO_2467 (O_2467,N_24809,N_22184);
nand UO_2468 (O_2468,N_22751,N_24896);
or UO_2469 (O_2469,N_22103,N_24135);
nor UO_2470 (O_2470,N_23937,N_22304);
xnor UO_2471 (O_2471,N_22401,N_22589);
xor UO_2472 (O_2472,N_24083,N_24589);
nor UO_2473 (O_2473,N_24908,N_22224);
xnor UO_2474 (O_2474,N_24316,N_22859);
and UO_2475 (O_2475,N_24857,N_24243);
nand UO_2476 (O_2476,N_22535,N_23242);
and UO_2477 (O_2477,N_21920,N_22684);
nand UO_2478 (O_2478,N_22401,N_24976);
xnor UO_2479 (O_2479,N_22108,N_23017);
or UO_2480 (O_2480,N_23751,N_22693);
and UO_2481 (O_2481,N_22923,N_24800);
xor UO_2482 (O_2482,N_24909,N_23037);
nor UO_2483 (O_2483,N_22243,N_24983);
xor UO_2484 (O_2484,N_22313,N_24582);
nand UO_2485 (O_2485,N_22121,N_24739);
nand UO_2486 (O_2486,N_24746,N_22797);
nand UO_2487 (O_2487,N_24772,N_22086);
nand UO_2488 (O_2488,N_23745,N_23547);
and UO_2489 (O_2489,N_24200,N_21945);
nand UO_2490 (O_2490,N_23327,N_22253);
or UO_2491 (O_2491,N_24337,N_24008);
nand UO_2492 (O_2492,N_22709,N_22817);
nor UO_2493 (O_2493,N_22321,N_23888);
and UO_2494 (O_2494,N_24147,N_22124);
or UO_2495 (O_2495,N_24883,N_22489);
and UO_2496 (O_2496,N_22299,N_24860);
nor UO_2497 (O_2497,N_23339,N_22224);
nand UO_2498 (O_2498,N_24663,N_23209);
or UO_2499 (O_2499,N_23539,N_22944);
and UO_2500 (O_2500,N_23505,N_22729);
and UO_2501 (O_2501,N_24588,N_22397);
or UO_2502 (O_2502,N_24826,N_23568);
nor UO_2503 (O_2503,N_22844,N_22646);
xor UO_2504 (O_2504,N_24405,N_22567);
xnor UO_2505 (O_2505,N_24579,N_23828);
nor UO_2506 (O_2506,N_22683,N_23424);
nand UO_2507 (O_2507,N_24893,N_22042);
xor UO_2508 (O_2508,N_23341,N_24028);
xnor UO_2509 (O_2509,N_23562,N_24474);
xor UO_2510 (O_2510,N_22990,N_23666);
xor UO_2511 (O_2511,N_24527,N_23078);
nand UO_2512 (O_2512,N_24334,N_22828);
xnor UO_2513 (O_2513,N_24475,N_22463);
and UO_2514 (O_2514,N_23509,N_24507);
nor UO_2515 (O_2515,N_24087,N_24816);
xnor UO_2516 (O_2516,N_24227,N_24151);
xnor UO_2517 (O_2517,N_23653,N_23769);
xor UO_2518 (O_2518,N_22412,N_23610);
xor UO_2519 (O_2519,N_23944,N_23170);
or UO_2520 (O_2520,N_22860,N_22589);
nand UO_2521 (O_2521,N_24215,N_24797);
and UO_2522 (O_2522,N_22228,N_24305);
nand UO_2523 (O_2523,N_23741,N_24686);
nor UO_2524 (O_2524,N_24422,N_23789);
nor UO_2525 (O_2525,N_24319,N_22172);
or UO_2526 (O_2526,N_22779,N_21909);
and UO_2527 (O_2527,N_22206,N_22403);
or UO_2528 (O_2528,N_24653,N_23800);
xnor UO_2529 (O_2529,N_24927,N_22191);
or UO_2530 (O_2530,N_22418,N_23970);
or UO_2531 (O_2531,N_22715,N_23931);
xor UO_2532 (O_2532,N_21881,N_22553);
or UO_2533 (O_2533,N_24409,N_23464);
nand UO_2534 (O_2534,N_23390,N_22225);
xnor UO_2535 (O_2535,N_22074,N_22124);
nor UO_2536 (O_2536,N_24934,N_23091);
nand UO_2537 (O_2537,N_22459,N_22756);
nand UO_2538 (O_2538,N_23863,N_24744);
nor UO_2539 (O_2539,N_23457,N_23215);
nor UO_2540 (O_2540,N_23394,N_22114);
and UO_2541 (O_2541,N_24415,N_23787);
and UO_2542 (O_2542,N_24832,N_24515);
and UO_2543 (O_2543,N_24274,N_24237);
or UO_2544 (O_2544,N_23881,N_22593);
nand UO_2545 (O_2545,N_24553,N_24484);
and UO_2546 (O_2546,N_24236,N_23071);
and UO_2547 (O_2547,N_22077,N_23440);
nor UO_2548 (O_2548,N_22089,N_23475);
and UO_2549 (O_2549,N_22632,N_22663);
nand UO_2550 (O_2550,N_24750,N_24742);
or UO_2551 (O_2551,N_22257,N_22176);
xor UO_2552 (O_2552,N_21953,N_24808);
nor UO_2553 (O_2553,N_24421,N_23248);
xnor UO_2554 (O_2554,N_21890,N_23113);
or UO_2555 (O_2555,N_23179,N_24208);
nor UO_2556 (O_2556,N_24178,N_24327);
nor UO_2557 (O_2557,N_23430,N_22280);
or UO_2558 (O_2558,N_23733,N_24685);
xnor UO_2559 (O_2559,N_22397,N_23835);
nand UO_2560 (O_2560,N_23652,N_23222);
or UO_2561 (O_2561,N_24216,N_22598);
or UO_2562 (O_2562,N_23779,N_22738);
and UO_2563 (O_2563,N_22140,N_21994);
and UO_2564 (O_2564,N_24199,N_24885);
or UO_2565 (O_2565,N_23870,N_23160);
xor UO_2566 (O_2566,N_23006,N_23886);
and UO_2567 (O_2567,N_24766,N_24431);
nand UO_2568 (O_2568,N_22501,N_24113);
or UO_2569 (O_2569,N_24234,N_22894);
and UO_2570 (O_2570,N_23039,N_22598);
or UO_2571 (O_2571,N_22099,N_22808);
nand UO_2572 (O_2572,N_23773,N_23260);
nor UO_2573 (O_2573,N_22468,N_23529);
nor UO_2574 (O_2574,N_22185,N_23200);
xnor UO_2575 (O_2575,N_22738,N_22180);
and UO_2576 (O_2576,N_22214,N_23004);
and UO_2577 (O_2577,N_22679,N_22568);
or UO_2578 (O_2578,N_22064,N_23946);
and UO_2579 (O_2579,N_22200,N_22882);
or UO_2580 (O_2580,N_22841,N_21960);
xor UO_2581 (O_2581,N_24012,N_22281);
xnor UO_2582 (O_2582,N_23517,N_23335);
and UO_2583 (O_2583,N_24464,N_24911);
nor UO_2584 (O_2584,N_24928,N_23723);
nor UO_2585 (O_2585,N_21941,N_24562);
nor UO_2586 (O_2586,N_23367,N_23826);
nor UO_2587 (O_2587,N_22121,N_24714);
or UO_2588 (O_2588,N_24664,N_24231);
nor UO_2589 (O_2589,N_22862,N_22785);
xor UO_2590 (O_2590,N_22293,N_24135);
nor UO_2591 (O_2591,N_24447,N_22211);
nand UO_2592 (O_2592,N_22539,N_24563);
xnor UO_2593 (O_2593,N_22616,N_24115);
nor UO_2594 (O_2594,N_23652,N_21888);
nand UO_2595 (O_2595,N_24537,N_24292);
xor UO_2596 (O_2596,N_23786,N_24734);
nor UO_2597 (O_2597,N_22468,N_22386);
nor UO_2598 (O_2598,N_22571,N_22679);
nand UO_2599 (O_2599,N_23464,N_23753);
nand UO_2600 (O_2600,N_24429,N_24043);
nand UO_2601 (O_2601,N_22644,N_22346);
nand UO_2602 (O_2602,N_22033,N_24953);
and UO_2603 (O_2603,N_22284,N_23202);
and UO_2604 (O_2604,N_23608,N_22948);
nand UO_2605 (O_2605,N_22747,N_22527);
or UO_2606 (O_2606,N_24179,N_23631);
nand UO_2607 (O_2607,N_23292,N_22532);
nor UO_2608 (O_2608,N_22266,N_24261);
and UO_2609 (O_2609,N_22210,N_22308);
nand UO_2610 (O_2610,N_24382,N_22973);
nand UO_2611 (O_2611,N_22788,N_21926);
nor UO_2612 (O_2612,N_22459,N_22931);
nand UO_2613 (O_2613,N_24108,N_24370);
or UO_2614 (O_2614,N_22680,N_24325);
or UO_2615 (O_2615,N_23558,N_21961);
and UO_2616 (O_2616,N_22023,N_21888);
nor UO_2617 (O_2617,N_24759,N_24114);
nor UO_2618 (O_2618,N_24480,N_22167);
nor UO_2619 (O_2619,N_22061,N_23069);
nand UO_2620 (O_2620,N_23023,N_23948);
nand UO_2621 (O_2621,N_24034,N_23196);
and UO_2622 (O_2622,N_22711,N_22986);
and UO_2623 (O_2623,N_24700,N_24709);
xor UO_2624 (O_2624,N_24437,N_23278);
or UO_2625 (O_2625,N_23159,N_23294);
nand UO_2626 (O_2626,N_24460,N_24439);
xor UO_2627 (O_2627,N_24329,N_24241);
nor UO_2628 (O_2628,N_23632,N_22753);
xor UO_2629 (O_2629,N_24435,N_23447);
and UO_2630 (O_2630,N_22329,N_24077);
or UO_2631 (O_2631,N_22810,N_23402);
nor UO_2632 (O_2632,N_22190,N_23735);
xor UO_2633 (O_2633,N_23740,N_22442);
or UO_2634 (O_2634,N_24051,N_23551);
nand UO_2635 (O_2635,N_23433,N_24855);
and UO_2636 (O_2636,N_24878,N_22477);
nand UO_2637 (O_2637,N_22848,N_22276);
or UO_2638 (O_2638,N_23085,N_22510);
xor UO_2639 (O_2639,N_24516,N_22668);
and UO_2640 (O_2640,N_23411,N_24417);
xor UO_2641 (O_2641,N_22556,N_23324);
nor UO_2642 (O_2642,N_23383,N_23670);
nor UO_2643 (O_2643,N_23875,N_22617);
and UO_2644 (O_2644,N_24736,N_22758);
nor UO_2645 (O_2645,N_23282,N_21902);
and UO_2646 (O_2646,N_23768,N_24345);
and UO_2647 (O_2647,N_23384,N_22520);
and UO_2648 (O_2648,N_22593,N_24266);
and UO_2649 (O_2649,N_23969,N_22025);
or UO_2650 (O_2650,N_23894,N_24863);
xnor UO_2651 (O_2651,N_24418,N_23042);
nand UO_2652 (O_2652,N_24483,N_23420);
or UO_2653 (O_2653,N_22676,N_24691);
and UO_2654 (O_2654,N_23735,N_22308);
or UO_2655 (O_2655,N_24668,N_24986);
nand UO_2656 (O_2656,N_22848,N_24963);
nand UO_2657 (O_2657,N_23074,N_23605);
and UO_2658 (O_2658,N_22830,N_22177);
nor UO_2659 (O_2659,N_24301,N_22455);
or UO_2660 (O_2660,N_23217,N_24432);
nand UO_2661 (O_2661,N_24222,N_23850);
or UO_2662 (O_2662,N_24819,N_22681);
xnor UO_2663 (O_2663,N_22310,N_23846);
nand UO_2664 (O_2664,N_23563,N_24801);
and UO_2665 (O_2665,N_24230,N_24317);
and UO_2666 (O_2666,N_24791,N_24826);
nor UO_2667 (O_2667,N_23476,N_24806);
nand UO_2668 (O_2668,N_24899,N_22841);
or UO_2669 (O_2669,N_21877,N_24691);
nand UO_2670 (O_2670,N_24417,N_23113);
and UO_2671 (O_2671,N_21972,N_22517);
xnor UO_2672 (O_2672,N_23164,N_22658);
nand UO_2673 (O_2673,N_23886,N_23284);
xnor UO_2674 (O_2674,N_24224,N_24029);
and UO_2675 (O_2675,N_24541,N_22617);
or UO_2676 (O_2676,N_24386,N_22650);
or UO_2677 (O_2677,N_22994,N_22197);
nand UO_2678 (O_2678,N_24316,N_24846);
and UO_2679 (O_2679,N_23710,N_24350);
or UO_2680 (O_2680,N_22455,N_24615);
xnor UO_2681 (O_2681,N_23953,N_24683);
nand UO_2682 (O_2682,N_22664,N_22097);
nand UO_2683 (O_2683,N_24933,N_23231);
nor UO_2684 (O_2684,N_24290,N_22687);
xor UO_2685 (O_2685,N_24656,N_22738);
or UO_2686 (O_2686,N_23960,N_24406);
or UO_2687 (O_2687,N_24605,N_24404);
nand UO_2688 (O_2688,N_22300,N_23746);
nand UO_2689 (O_2689,N_22861,N_24810);
nor UO_2690 (O_2690,N_23383,N_23799);
and UO_2691 (O_2691,N_22278,N_23127);
nand UO_2692 (O_2692,N_22354,N_22861);
or UO_2693 (O_2693,N_24928,N_23986);
and UO_2694 (O_2694,N_22789,N_23368);
xor UO_2695 (O_2695,N_23288,N_22603);
nor UO_2696 (O_2696,N_23438,N_23112);
nand UO_2697 (O_2697,N_24608,N_24728);
nor UO_2698 (O_2698,N_22164,N_23961);
nand UO_2699 (O_2699,N_24893,N_24765);
or UO_2700 (O_2700,N_24922,N_24620);
nand UO_2701 (O_2701,N_23801,N_22589);
and UO_2702 (O_2702,N_24689,N_23000);
xor UO_2703 (O_2703,N_23847,N_24529);
xnor UO_2704 (O_2704,N_24029,N_22508);
nor UO_2705 (O_2705,N_24189,N_23961);
and UO_2706 (O_2706,N_24951,N_22081);
or UO_2707 (O_2707,N_22492,N_22170);
xnor UO_2708 (O_2708,N_24719,N_23111);
or UO_2709 (O_2709,N_24401,N_22402);
and UO_2710 (O_2710,N_23102,N_22677);
xor UO_2711 (O_2711,N_24934,N_24479);
nand UO_2712 (O_2712,N_22214,N_24979);
and UO_2713 (O_2713,N_21932,N_24017);
or UO_2714 (O_2714,N_23074,N_22967);
or UO_2715 (O_2715,N_24146,N_23219);
or UO_2716 (O_2716,N_24904,N_22389);
nand UO_2717 (O_2717,N_24156,N_23746);
and UO_2718 (O_2718,N_23892,N_22310);
xnor UO_2719 (O_2719,N_23680,N_24126);
nand UO_2720 (O_2720,N_21932,N_22795);
xnor UO_2721 (O_2721,N_22014,N_22390);
nor UO_2722 (O_2722,N_23912,N_22361);
nor UO_2723 (O_2723,N_24780,N_24880);
nand UO_2724 (O_2724,N_23998,N_22396);
xnor UO_2725 (O_2725,N_23489,N_23049);
xor UO_2726 (O_2726,N_24851,N_24305);
and UO_2727 (O_2727,N_22733,N_21879);
or UO_2728 (O_2728,N_23831,N_23803);
or UO_2729 (O_2729,N_21964,N_23466);
nor UO_2730 (O_2730,N_22226,N_24190);
nand UO_2731 (O_2731,N_22623,N_22497);
or UO_2732 (O_2732,N_24458,N_24601);
nand UO_2733 (O_2733,N_23217,N_24790);
xor UO_2734 (O_2734,N_22498,N_22859);
nand UO_2735 (O_2735,N_22653,N_23716);
or UO_2736 (O_2736,N_23548,N_23633);
nand UO_2737 (O_2737,N_22590,N_24660);
or UO_2738 (O_2738,N_22764,N_23310);
nand UO_2739 (O_2739,N_22614,N_23830);
and UO_2740 (O_2740,N_23652,N_24064);
xor UO_2741 (O_2741,N_23040,N_21985);
nand UO_2742 (O_2742,N_22517,N_23590);
nand UO_2743 (O_2743,N_24427,N_24125);
or UO_2744 (O_2744,N_23555,N_24165);
or UO_2745 (O_2745,N_22189,N_24723);
and UO_2746 (O_2746,N_23291,N_23540);
nand UO_2747 (O_2747,N_23900,N_22397);
xnor UO_2748 (O_2748,N_24040,N_22786);
and UO_2749 (O_2749,N_24371,N_22512);
xnor UO_2750 (O_2750,N_24166,N_22569);
or UO_2751 (O_2751,N_23539,N_21931);
xnor UO_2752 (O_2752,N_22668,N_22103);
nor UO_2753 (O_2753,N_24941,N_22283);
nand UO_2754 (O_2754,N_24552,N_23188);
and UO_2755 (O_2755,N_24289,N_24138);
nor UO_2756 (O_2756,N_23464,N_24385);
nand UO_2757 (O_2757,N_22210,N_21939);
and UO_2758 (O_2758,N_21915,N_23384);
or UO_2759 (O_2759,N_24006,N_22059);
or UO_2760 (O_2760,N_24205,N_22816);
or UO_2761 (O_2761,N_23662,N_23311);
nand UO_2762 (O_2762,N_22579,N_23567);
nand UO_2763 (O_2763,N_23327,N_23991);
or UO_2764 (O_2764,N_24182,N_23815);
xnor UO_2765 (O_2765,N_23376,N_22067);
xnor UO_2766 (O_2766,N_23303,N_24953);
or UO_2767 (O_2767,N_24124,N_22394);
or UO_2768 (O_2768,N_23877,N_22825);
or UO_2769 (O_2769,N_24808,N_22276);
or UO_2770 (O_2770,N_23734,N_22955);
nand UO_2771 (O_2771,N_22277,N_22692);
or UO_2772 (O_2772,N_22996,N_21876);
nand UO_2773 (O_2773,N_24297,N_23255);
and UO_2774 (O_2774,N_23909,N_22571);
or UO_2775 (O_2775,N_22767,N_24906);
xor UO_2776 (O_2776,N_22276,N_23204);
xor UO_2777 (O_2777,N_24742,N_23131);
xor UO_2778 (O_2778,N_24139,N_23167);
nand UO_2779 (O_2779,N_23254,N_23018);
xor UO_2780 (O_2780,N_23370,N_23108);
or UO_2781 (O_2781,N_24419,N_24744);
nand UO_2782 (O_2782,N_24209,N_23395);
xor UO_2783 (O_2783,N_24782,N_23450);
nor UO_2784 (O_2784,N_24285,N_22176);
nand UO_2785 (O_2785,N_22498,N_22445);
nand UO_2786 (O_2786,N_23427,N_22132);
nand UO_2787 (O_2787,N_23286,N_24401);
nor UO_2788 (O_2788,N_24331,N_24799);
nand UO_2789 (O_2789,N_22484,N_24907);
nor UO_2790 (O_2790,N_24118,N_23109);
and UO_2791 (O_2791,N_22581,N_22920);
nor UO_2792 (O_2792,N_24803,N_24515);
and UO_2793 (O_2793,N_23731,N_24511);
nor UO_2794 (O_2794,N_21905,N_24033);
nor UO_2795 (O_2795,N_24297,N_24022);
or UO_2796 (O_2796,N_23180,N_22371);
or UO_2797 (O_2797,N_22727,N_24065);
nand UO_2798 (O_2798,N_22135,N_23849);
nand UO_2799 (O_2799,N_22770,N_22509);
or UO_2800 (O_2800,N_23609,N_23961);
nand UO_2801 (O_2801,N_23248,N_22103);
xor UO_2802 (O_2802,N_22482,N_23247);
and UO_2803 (O_2803,N_23149,N_23818);
nand UO_2804 (O_2804,N_24682,N_22802);
xor UO_2805 (O_2805,N_22890,N_23495);
or UO_2806 (O_2806,N_22839,N_23854);
nor UO_2807 (O_2807,N_22335,N_23232);
nor UO_2808 (O_2808,N_24925,N_24370);
or UO_2809 (O_2809,N_23878,N_22674);
nand UO_2810 (O_2810,N_24294,N_23686);
nand UO_2811 (O_2811,N_22278,N_23113);
and UO_2812 (O_2812,N_24710,N_22062);
nand UO_2813 (O_2813,N_22250,N_22073);
and UO_2814 (O_2814,N_23435,N_24496);
nand UO_2815 (O_2815,N_23449,N_24176);
nor UO_2816 (O_2816,N_24330,N_23135);
xnor UO_2817 (O_2817,N_21985,N_24531);
and UO_2818 (O_2818,N_24027,N_21935);
nand UO_2819 (O_2819,N_23332,N_24699);
and UO_2820 (O_2820,N_23086,N_22767);
and UO_2821 (O_2821,N_24250,N_24517);
nand UO_2822 (O_2822,N_23359,N_22248);
xor UO_2823 (O_2823,N_22772,N_24025);
and UO_2824 (O_2824,N_23041,N_22310);
or UO_2825 (O_2825,N_23380,N_23132);
nand UO_2826 (O_2826,N_24358,N_24045);
nor UO_2827 (O_2827,N_24695,N_23545);
nand UO_2828 (O_2828,N_24099,N_22252);
nor UO_2829 (O_2829,N_23643,N_23483);
xnor UO_2830 (O_2830,N_23144,N_23229);
and UO_2831 (O_2831,N_24921,N_23500);
and UO_2832 (O_2832,N_24751,N_22916);
nor UO_2833 (O_2833,N_23728,N_23881);
xor UO_2834 (O_2834,N_24265,N_24871);
and UO_2835 (O_2835,N_23598,N_24289);
xor UO_2836 (O_2836,N_24895,N_22928);
or UO_2837 (O_2837,N_24993,N_22640);
and UO_2838 (O_2838,N_22371,N_21895);
or UO_2839 (O_2839,N_24944,N_24858);
or UO_2840 (O_2840,N_22127,N_21913);
or UO_2841 (O_2841,N_22909,N_23503);
nand UO_2842 (O_2842,N_22839,N_22910);
or UO_2843 (O_2843,N_24650,N_24758);
xnor UO_2844 (O_2844,N_24301,N_24489);
nand UO_2845 (O_2845,N_24384,N_24412);
or UO_2846 (O_2846,N_24769,N_23649);
or UO_2847 (O_2847,N_24978,N_22652);
or UO_2848 (O_2848,N_24074,N_24902);
nor UO_2849 (O_2849,N_24633,N_23673);
and UO_2850 (O_2850,N_22218,N_24010);
nor UO_2851 (O_2851,N_22444,N_23761);
nand UO_2852 (O_2852,N_24897,N_23339);
nor UO_2853 (O_2853,N_22339,N_23215);
nand UO_2854 (O_2854,N_23259,N_23854);
xnor UO_2855 (O_2855,N_23170,N_21960);
and UO_2856 (O_2856,N_22639,N_22653);
or UO_2857 (O_2857,N_24156,N_23576);
xnor UO_2858 (O_2858,N_23281,N_24335);
xnor UO_2859 (O_2859,N_24374,N_24808);
nand UO_2860 (O_2860,N_22174,N_24072);
or UO_2861 (O_2861,N_24335,N_23066);
or UO_2862 (O_2862,N_23028,N_23933);
and UO_2863 (O_2863,N_24694,N_24178);
nor UO_2864 (O_2864,N_24509,N_22096);
and UO_2865 (O_2865,N_24700,N_22940);
or UO_2866 (O_2866,N_22518,N_23147);
nor UO_2867 (O_2867,N_23346,N_23327);
or UO_2868 (O_2868,N_23957,N_22738);
nand UO_2869 (O_2869,N_24894,N_22227);
nor UO_2870 (O_2870,N_23292,N_24994);
or UO_2871 (O_2871,N_23350,N_22135);
or UO_2872 (O_2872,N_22794,N_22571);
and UO_2873 (O_2873,N_22332,N_24044);
or UO_2874 (O_2874,N_23475,N_23106);
and UO_2875 (O_2875,N_23840,N_23552);
nor UO_2876 (O_2876,N_21985,N_22614);
nand UO_2877 (O_2877,N_23143,N_23976);
and UO_2878 (O_2878,N_23380,N_22979);
nand UO_2879 (O_2879,N_22583,N_24803);
or UO_2880 (O_2880,N_22519,N_23422);
xnor UO_2881 (O_2881,N_22663,N_22865);
xor UO_2882 (O_2882,N_22387,N_22391);
or UO_2883 (O_2883,N_23227,N_24688);
or UO_2884 (O_2884,N_22644,N_22729);
or UO_2885 (O_2885,N_21971,N_23892);
nor UO_2886 (O_2886,N_23219,N_23795);
or UO_2887 (O_2887,N_22340,N_23473);
nand UO_2888 (O_2888,N_24174,N_22069);
or UO_2889 (O_2889,N_23166,N_24924);
nor UO_2890 (O_2890,N_22845,N_22288);
xnor UO_2891 (O_2891,N_21984,N_24068);
and UO_2892 (O_2892,N_24216,N_22215);
xor UO_2893 (O_2893,N_22727,N_24706);
nor UO_2894 (O_2894,N_22097,N_23983);
xor UO_2895 (O_2895,N_22577,N_23543);
nand UO_2896 (O_2896,N_22052,N_23403);
and UO_2897 (O_2897,N_22183,N_22243);
and UO_2898 (O_2898,N_23201,N_24899);
nor UO_2899 (O_2899,N_22594,N_24780);
xnor UO_2900 (O_2900,N_22955,N_23098);
and UO_2901 (O_2901,N_23643,N_24692);
nand UO_2902 (O_2902,N_24020,N_22877);
or UO_2903 (O_2903,N_24122,N_23521);
and UO_2904 (O_2904,N_23015,N_24754);
nand UO_2905 (O_2905,N_24000,N_21986);
or UO_2906 (O_2906,N_22268,N_22016);
nand UO_2907 (O_2907,N_23161,N_23376);
and UO_2908 (O_2908,N_24961,N_23534);
xnor UO_2909 (O_2909,N_22886,N_23079);
nand UO_2910 (O_2910,N_22502,N_24228);
xor UO_2911 (O_2911,N_22864,N_24110);
or UO_2912 (O_2912,N_24621,N_22776);
xnor UO_2913 (O_2913,N_22203,N_24800);
nor UO_2914 (O_2914,N_24223,N_22946);
nor UO_2915 (O_2915,N_24367,N_24557);
and UO_2916 (O_2916,N_22426,N_22805);
nor UO_2917 (O_2917,N_24342,N_21932);
and UO_2918 (O_2918,N_24638,N_22819);
nand UO_2919 (O_2919,N_24293,N_24883);
nand UO_2920 (O_2920,N_22050,N_24188);
or UO_2921 (O_2921,N_21911,N_24958);
and UO_2922 (O_2922,N_23040,N_23373);
nor UO_2923 (O_2923,N_23725,N_22586);
nand UO_2924 (O_2924,N_23743,N_23830);
nor UO_2925 (O_2925,N_21971,N_23071);
nand UO_2926 (O_2926,N_24805,N_22102);
or UO_2927 (O_2927,N_23283,N_24864);
xor UO_2928 (O_2928,N_24292,N_24419);
nor UO_2929 (O_2929,N_22330,N_23175);
and UO_2930 (O_2930,N_23528,N_23162);
nor UO_2931 (O_2931,N_23829,N_24336);
nand UO_2932 (O_2932,N_22518,N_23457);
nor UO_2933 (O_2933,N_23142,N_22864);
or UO_2934 (O_2934,N_24798,N_23247);
and UO_2935 (O_2935,N_24751,N_24651);
nor UO_2936 (O_2936,N_24275,N_24806);
nand UO_2937 (O_2937,N_22040,N_22015);
and UO_2938 (O_2938,N_23715,N_24444);
and UO_2939 (O_2939,N_24875,N_23532);
xnor UO_2940 (O_2940,N_24223,N_24207);
nand UO_2941 (O_2941,N_24108,N_23521);
or UO_2942 (O_2942,N_23471,N_23555);
nand UO_2943 (O_2943,N_23065,N_24857);
or UO_2944 (O_2944,N_22550,N_23591);
nor UO_2945 (O_2945,N_22979,N_24171);
xor UO_2946 (O_2946,N_22576,N_24768);
xnor UO_2947 (O_2947,N_24751,N_24632);
nor UO_2948 (O_2948,N_24045,N_23068);
or UO_2949 (O_2949,N_24089,N_24292);
xor UO_2950 (O_2950,N_22009,N_24079);
xor UO_2951 (O_2951,N_24276,N_23995);
nand UO_2952 (O_2952,N_24743,N_22016);
and UO_2953 (O_2953,N_21957,N_24714);
nand UO_2954 (O_2954,N_23985,N_24382);
and UO_2955 (O_2955,N_24281,N_24781);
or UO_2956 (O_2956,N_22504,N_23112);
and UO_2957 (O_2957,N_23106,N_22915);
nand UO_2958 (O_2958,N_24893,N_23148);
and UO_2959 (O_2959,N_22188,N_24895);
and UO_2960 (O_2960,N_24629,N_23764);
nor UO_2961 (O_2961,N_23338,N_23462);
nor UO_2962 (O_2962,N_24024,N_23144);
and UO_2963 (O_2963,N_22661,N_23247);
nor UO_2964 (O_2964,N_22670,N_24841);
or UO_2965 (O_2965,N_22571,N_23300);
xnor UO_2966 (O_2966,N_23602,N_23388);
or UO_2967 (O_2967,N_23843,N_24454);
nor UO_2968 (O_2968,N_21904,N_24224);
nor UO_2969 (O_2969,N_23492,N_24827);
and UO_2970 (O_2970,N_23330,N_23386);
or UO_2971 (O_2971,N_22885,N_23046);
nand UO_2972 (O_2972,N_22364,N_21890);
and UO_2973 (O_2973,N_24794,N_22158);
xor UO_2974 (O_2974,N_21896,N_24165);
xor UO_2975 (O_2975,N_22977,N_24391);
nand UO_2976 (O_2976,N_23785,N_22675);
xnor UO_2977 (O_2977,N_22566,N_24513);
and UO_2978 (O_2978,N_21892,N_24796);
nand UO_2979 (O_2979,N_22519,N_24752);
or UO_2980 (O_2980,N_22832,N_22769);
xnor UO_2981 (O_2981,N_24562,N_23313);
xor UO_2982 (O_2982,N_23778,N_23104);
nor UO_2983 (O_2983,N_23686,N_22574);
nand UO_2984 (O_2984,N_24927,N_21991);
and UO_2985 (O_2985,N_24650,N_24535);
and UO_2986 (O_2986,N_22323,N_23750);
nand UO_2987 (O_2987,N_23105,N_24263);
and UO_2988 (O_2988,N_23855,N_24623);
and UO_2989 (O_2989,N_23106,N_23043);
or UO_2990 (O_2990,N_22983,N_24624);
nor UO_2991 (O_2991,N_23158,N_24096);
nand UO_2992 (O_2992,N_24200,N_23171);
nand UO_2993 (O_2993,N_24842,N_23372);
nor UO_2994 (O_2994,N_23786,N_23697);
or UO_2995 (O_2995,N_23958,N_23884);
nand UO_2996 (O_2996,N_22803,N_22067);
nor UO_2997 (O_2997,N_24730,N_24947);
nand UO_2998 (O_2998,N_22144,N_22813);
nand UO_2999 (O_2999,N_23018,N_24441);
endmodule