module basic_2000_20000_2500_10_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_1398,In_132);
and U1 (N_1,In_257,In_566);
nor U2 (N_2,In_880,In_1038);
and U3 (N_3,In_58,In_349);
nor U4 (N_4,In_1947,In_142);
or U5 (N_5,In_243,In_202);
or U6 (N_6,In_1774,In_1921);
or U7 (N_7,In_1417,In_838);
nand U8 (N_8,In_1838,In_1261);
xor U9 (N_9,In_864,In_401);
and U10 (N_10,In_876,In_522);
nor U11 (N_11,In_34,In_1968);
nand U12 (N_12,In_1394,In_48);
and U13 (N_13,In_151,In_568);
and U14 (N_14,In_1413,In_23);
nor U15 (N_15,In_1965,In_1804);
xnor U16 (N_16,In_1125,In_1870);
nor U17 (N_17,In_930,In_67);
and U18 (N_18,In_613,In_532);
nor U19 (N_19,In_817,In_915);
xor U20 (N_20,In_1752,In_1118);
and U21 (N_21,In_314,In_1879);
and U22 (N_22,In_491,In_321);
nand U23 (N_23,In_1946,In_1541);
or U24 (N_24,In_1633,In_604);
nor U25 (N_25,In_1908,In_1942);
nand U26 (N_26,In_1450,In_1717);
or U27 (N_27,In_984,In_1584);
or U28 (N_28,In_1084,In_700);
or U29 (N_29,In_160,In_1520);
nand U30 (N_30,In_1052,In_430);
nand U31 (N_31,In_499,In_1409);
nand U32 (N_32,In_1978,In_705);
nor U33 (N_33,In_1185,In_1535);
nand U34 (N_34,In_572,In_500);
and U35 (N_35,In_1618,In_1777);
nand U36 (N_36,In_626,In_1845);
or U37 (N_37,In_1191,In_1435);
nand U38 (N_38,In_1987,In_258);
or U39 (N_39,In_559,In_737);
xor U40 (N_40,In_1540,In_636);
nand U41 (N_41,In_74,In_1739);
xnor U42 (N_42,In_341,In_459);
and U43 (N_43,In_133,In_553);
nand U44 (N_44,In_480,In_1104);
nand U45 (N_45,In_198,In_666);
or U46 (N_46,In_32,In_652);
nand U47 (N_47,In_71,In_1682);
nand U48 (N_48,In_1677,In_280);
xor U49 (N_49,In_1243,In_1044);
xnor U50 (N_50,In_1267,In_503);
xor U51 (N_51,In_281,In_954);
nor U52 (N_52,In_1276,In_965);
nand U53 (N_53,In_609,In_55);
or U54 (N_54,In_1762,In_1933);
or U55 (N_55,In_1501,In_1523);
nor U56 (N_56,In_795,In_37);
xnor U57 (N_57,In_1577,In_1491);
xnor U58 (N_58,In_749,In_733);
and U59 (N_59,In_813,In_1740);
or U60 (N_60,In_1241,In_301);
nor U61 (N_61,In_1317,In_1952);
xnor U62 (N_62,In_1672,In_1602);
xor U63 (N_63,In_1625,In_247);
and U64 (N_64,In_428,In_1221);
nand U65 (N_65,In_688,In_200);
xor U66 (N_66,In_1371,In_981);
nand U67 (N_67,In_106,In_1109);
xor U68 (N_68,In_110,In_881);
and U69 (N_69,In_35,In_972);
and U70 (N_70,In_508,In_1055);
and U71 (N_71,In_858,In_1755);
nor U72 (N_72,In_1454,In_1658);
nor U73 (N_73,In_339,In_1381);
nand U74 (N_74,In_1126,In_1863);
and U75 (N_75,In_1641,In_820);
or U76 (N_76,In_1843,In_1715);
and U77 (N_77,In_1343,In_496);
xor U78 (N_78,In_282,In_318);
nor U79 (N_79,In_1709,In_454);
xnor U80 (N_80,In_674,In_1420);
or U81 (N_81,In_1472,In_939);
or U82 (N_82,In_676,In_1585);
and U83 (N_83,In_1418,In_958);
xor U84 (N_84,In_1822,In_1610);
and U85 (N_85,In_1669,In_1369);
xor U86 (N_86,In_1265,In_1462);
and U87 (N_87,In_1237,In_533);
or U88 (N_88,In_1915,In_1581);
nand U89 (N_89,In_1897,In_81);
nor U90 (N_90,In_125,In_1090);
nand U91 (N_91,In_951,In_1884);
nand U92 (N_92,In_1920,In_1252);
xnor U93 (N_93,In_1964,In_1687);
nand U94 (N_94,In_1455,In_346);
nor U95 (N_95,In_36,In_543);
nor U96 (N_96,In_738,In_1207);
nor U97 (N_97,In_268,In_1594);
and U98 (N_98,In_1598,In_1567);
and U99 (N_99,In_1823,In_1324);
xnor U100 (N_100,In_902,In_1157);
nor U101 (N_101,In_860,In_1176);
xor U102 (N_102,In_1189,In_1726);
nor U103 (N_103,In_873,In_1169);
nand U104 (N_104,In_1129,In_344);
nand U105 (N_105,In_938,In_851);
nor U106 (N_106,In_1414,In_1539);
nor U107 (N_107,In_1917,In_1528);
nand U108 (N_108,In_596,In_1384);
nand U109 (N_109,In_1145,In_1851);
nor U110 (N_110,In_1623,In_424);
and U111 (N_111,In_1922,In_647);
nor U112 (N_112,In_659,In_1323);
nand U113 (N_113,In_933,In_461);
xnor U114 (N_114,In_161,In_837);
and U115 (N_115,In_1991,In_1608);
nand U116 (N_116,In_859,In_1825);
nor U117 (N_117,In_1914,In_1620);
nor U118 (N_118,In_1927,In_1614);
xor U119 (N_119,In_1305,In_1192);
and U120 (N_120,In_623,In_1375);
and U121 (N_121,In_1654,In_1582);
nand U122 (N_122,In_1484,In_1511);
and U123 (N_123,In_43,In_869);
xnor U124 (N_124,In_1216,In_2);
xnor U125 (N_125,In_1911,In_218);
and U126 (N_126,In_1986,In_1864);
xor U127 (N_127,In_645,In_1123);
or U128 (N_128,In_1703,In_669);
or U129 (N_129,In_630,In_152);
and U130 (N_130,In_1500,In_1200);
xnor U131 (N_131,In_1337,In_358);
or U132 (N_132,In_129,In_1552);
or U133 (N_133,In_1961,In_422);
nand U134 (N_134,In_548,In_1502);
nand U135 (N_135,In_1756,In_914);
and U136 (N_136,In_1956,In_657);
nor U137 (N_137,In_1763,In_692);
xor U138 (N_138,In_810,In_455);
nand U139 (N_139,In_1219,In_1376);
or U140 (N_140,In_174,In_1302);
nor U141 (N_141,In_671,In_1701);
nor U142 (N_142,In_94,In_1199);
or U143 (N_143,In_926,In_1174);
xor U144 (N_144,In_656,In_1209);
and U145 (N_145,In_1112,In_1729);
nor U146 (N_146,In_238,In_62);
nor U147 (N_147,In_662,In_169);
or U148 (N_148,In_56,In_342);
xor U149 (N_149,In_1827,In_1030);
and U150 (N_150,In_1613,In_1561);
and U151 (N_151,In_479,In_1270);
nand U152 (N_152,In_994,In_1143);
and U153 (N_153,In_70,In_554);
and U154 (N_154,In_610,In_897);
nor U155 (N_155,In_1114,In_396);
nor U156 (N_156,In_1635,In_1378);
or U157 (N_157,In_1116,In_381);
xnor U158 (N_158,In_911,In_478);
xnor U159 (N_159,In_1210,In_262);
nand U160 (N_160,In_557,In_1634);
xnor U161 (N_161,In_112,In_1045);
and U162 (N_162,In_865,In_1285);
xor U163 (N_163,In_1494,In_1767);
nand U164 (N_164,In_1251,In_421);
xnor U165 (N_165,In_1686,In_99);
nand U166 (N_166,In_1108,In_638);
and U167 (N_167,In_822,In_416);
or U168 (N_168,In_288,In_1306);
nor U169 (N_169,In_1008,In_473);
and U170 (N_170,In_376,In_1892);
or U171 (N_171,In_1440,In_1699);
nand U172 (N_172,In_1712,In_1458);
xnor U173 (N_173,In_304,In_360);
or U174 (N_174,In_80,In_483);
nor U175 (N_175,In_1431,In_1446);
nor U176 (N_176,In_1648,In_0);
or U177 (N_177,In_707,In_1731);
or U178 (N_178,In_1070,In_368);
nor U179 (N_179,In_1967,In_265);
or U180 (N_180,In_1548,In_516);
nand U181 (N_181,In_307,In_1031);
or U182 (N_182,In_527,In_690);
and U183 (N_183,In_1645,In_111);
and U184 (N_184,In_599,In_298);
xnor U185 (N_185,In_606,In_1773);
xnor U186 (N_186,In_1029,In_1906);
or U187 (N_187,In_825,In_1573);
and U188 (N_188,In_1258,In_661);
nor U189 (N_189,In_154,In_1903);
nor U190 (N_190,In_1292,In_1142);
nor U191 (N_191,In_1382,In_1061);
or U192 (N_192,In_577,In_155);
xnor U193 (N_193,In_847,In_38);
nand U194 (N_194,In_734,In_1867);
nor U195 (N_195,In_47,In_770);
nand U196 (N_196,In_745,In_1977);
nor U197 (N_197,In_1497,In_1795);
and U198 (N_198,In_1950,In_1487);
and U199 (N_199,In_1155,In_1283);
or U200 (N_200,In_1432,In_1589);
or U201 (N_201,In_1820,In_921);
xnor U202 (N_202,In_1543,In_1374);
nor U203 (N_203,In_1093,In_852);
or U204 (N_204,In_551,In_1346);
or U205 (N_205,In_1363,In_509);
xnor U206 (N_206,In_841,In_726);
nor U207 (N_207,In_168,In_150);
xnor U208 (N_208,In_1590,In_1367);
xor U209 (N_209,In_1099,In_937);
and U210 (N_210,In_1295,In_518);
xnor U211 (N_211,In_1460,In_196);
and U212 (N_212,In_333,In_1442);
or U213 (N_213,In_242,In_394);
and U214 (N_214,In_1779,In_1271);
nand U215 (N_215,In_1524,In_1507);
or U216 (N_216,In_840,In_1106);
nand U217 (N_217,In_1807,In_137);
nand U218 (N_218,In_1833,In_1678);
nand U219 (N_219,In_493,In_898);
and U220 (N_220,In_1385,In_1647);
and U221 (N_221,In_955,In_992);
nor U222 (N_222,In_205,In_1888);
and U223 (N_223,In_1165,In_1529);
nand U224 (N_224,In_1357,In_1105);
nor U225 (N_225,In_113,In_1742);
nor U226 (N_226,In_264,In_1336);
nor U227 (N_227,In_79,In_1916);
and U228 (N_228,In_970,In_59);
xnor U229 (N_229,In_1178,In_1799);
xor U230 (N_230,In_224,In_1904);
or U231 (N_231,In_251,In_791);
nor U232 (N_232,In_1347,In_547);
nor U233 (N_233,In_555,In_208);
nand U234 (N_234,In_886,In_1056);
nor U235 (N_235,In_124,In_767);
nand U236 (N_236,In_1344,In_250);
or U237 (N_237,In_1042,In_1248);
nand U238 (N_238,In_1203,In_1941);
nand U239 (N_239,In_1018,In_668);
nand U240 (N_240,In_52,In_269);
or U241 (N_241,In_350,In_906);
and U242 (N_242,In_1865,In_1342);
nand U243 (N_243,In_338,In_316);
or U244 (N_244,In_1495,In_140);
nor U245 (N_245,In_53,In_1201);
nor U246 (N_246,In_434,In_237);
and U247 (N_247,In_1315,In_1003);
nand U248 (N_248,In_404,In_611);
nand U249 (N_249,In_506,In_221);
or U250 (N_250,In_327,In_591);
xor U251 (N_251,In_1652,In_1452);
and U252 (N_252,In_57,In_724);
nand U253 (N_253,In_1282,In_1022);
and U254 (N_254,In_1229,In_1107);
and U255 (N_255,In_815,In_855);
or U256 (N_256,In_1300,In_1653);
or U257 (N_257,In_210,In_244);
and U258 (N_258,In_17,In_1049);
nand U259 (N_259,In_1828,In_903);
and U260 (N_260,In_313,In_76);
nor U261 (N_261,In_203,In_751);
nor U262 (N_262,In_386,In_138);
xnor U263 (N_263,In_718,In_417);
nor U264 (N_264,In_1738,In_904);
nor U265 (N_265,In_1788,In_1951);
or U266 (N_266,In_236,In_383);
nand U267 (N_267,In_1890,In_1747);
or U268 (N_268,In_1776,In_1745);
xnor U269 (N_269,In_413,In_393);
or U270 (N_270,In_1883,In_816);
xnor U271 (N_271,In_1429,In_165);
nor U272 (N_272,In_754,In_1547);
nand U273 (N_273,In_336,In_684);
or U274 (N_274,In_176,In_1069);
and U275 (N_275,In_1616,In_206);
nor U276 (N_276,In_698,In_995);
nand U277 (N_277,In_436,In_1041);
nand U278 (N_278,In_1887,In_1688);
and U279 (N_279,In_863,In_1604);
and U280 (N_280,In_1526,In_1422);
nand U281 (N_281,In_1278,In_447);
xnor U282 (N_282,In_1624,In_1316);
or U283 (N_283,In_530,In_340);
and U284 (N_284,In_1134,In_1530);
nor U285 (N_285,In_525,In_714);
xnor U286 (N_286,In_529,In_363);
nand U287 (N_287,In_60,In_1026);
and U288 (N_288,In_1962,In_655);
xor U289 (N_289,In_145,In_741);
nor U290 (N_290,In_1082,In_1274);
nor U291 (N_291,In_477,In_1483);
or U292 (N_292,In_432,In_390);
xnor U293 (N_293,In_1796,In_1100);
nand U294 (N_294,In_375,In_844);
nor U295 (N_295,In_940,In_1586);
xnor U296 (N_296,In_437,In_1372);
or U297 (N_297,In_1253,In_1621);
and U298 (N_298,In_1309,In_429);
nand U299 (N_299,In_632,In_1558);
nor U300 (N_300,In_1141,In_1945);
or U301 (N_301,In_1364,In_1628);
nor U302 (N_302,In_30,In_50);
and U303 (N_303,In_1240,In_905);
xnor U304 (N_304,In_1448,In_427);
and U305 (N_305,In_1263,In_1576);
nand U306 (N_306,In_91,In_1016);
nor U307 (N_307,In_1175,In_1683);
xor U308 (N_308,In_649,In_1695);
xor U309 (N_309,In_520,In_353);
nor U310 (N_310,In_1146,In_13);
or U311 (N_311,In_1733,In_1858);
and U312 (N_312,In_1939,In_848);
or U313 (N_313,In_1707,In_1362);
xor U314 (N_314,In_1330,In_252);
and U315 (N_315,In_1102,In_1238);
or U316 (N_316,In_687,In_1938);
and U317 (N_317,In_1859,In_123);
and U318 (N_318,In_971,In_1606);
or U319 (N_319,In_231,In_1296);
or U320 (N_320,In_209,In_107);
nand U321 (N_321,In_295,In_1474);
or U322 (N_322,In_845,In_470);
nor U323 (N_323,In_1937,In_1161);
nor U324 (N_324,In_788,In_1588);
nand U325 (N_325,In_722,In_809);
xor U326 (N_326,In_267,In_562);
nand U327 (N_327,In_1765,In_226);
nand U328 (N_328,In_354,In_488);
xor U329 (N_329,In_597,In_181);
xor U330 (N_330,In_1676,In_1486);
nor U331 (N_331,In_1087,In_255);
nand U332 (N_332,In_1025,In_1400);
xor U333 (N_333,In_1513,In_273);
nor U334 (N_334,In_1925,In_153);
and U335 (N_335,In_474,In_369);
xor U336 (N_336,In_1136,In_1640);
and U337 (N_337,In_1401,In_990);
and U338 (N_338,In_853,In_290);
xor U339 (N_339,In_234,In_1275);
xor U340 (N_340,In_31,In_157);
and U341 (N_341,In_512,In_1974);
or U342 (N_342,In_1813,In_576);
or U343 (N_343,In_69,In_1743);
nand U344 (N_344,In_1060,In_389);
nor U345 (N_345,In_9,In_1578);
nand U346 (N_346,In_1894,In_729);
nor U347 (N_347,In_1924,In_1352);
or U348 (N_348,In_1510,In_1272);
and U349 (N_349,In_245,In_792);
and U350 (N_350,In_410,In_539);
or U351 (N_351,In_634,In_1128);
and U352 (N_352,In_1390,In_85);
or U353 (N_353,In_1131,In_806);
nor U354 (N_354,In_1218,In_116);
xnor U355 (N_355,In_650,In_450);
or U356 (N_356,In_179,In_1047);
nand U357 (N_357,In_419,In_1284);
xor U358 (N_358,In_1919,In_117);
nand U359 (N_359,In_908,In_315);
or U360 (N_360,In_1525,In_1303);
and U361 (N_361,In_747,In_1195);
or U362 (N_362,In_872,In_783);
xnor U363 (N_363,In_1277,In_29);
nand U364 (N_364,In_789,In_292);
nand U365 (N_365,In_1963,In_183);
and U366 (N_366,In_736,In_949);
nor U367 (N_367,In_1913,In_1656);
nor U368 (N_368,In_1948,In_1032);
xor U369 (N_369,In_1990,In_579);
nand U370 (N_370,In_1465,In_833);
nand U371 (N_371,In_1716,In_286);
and U372 (N_372,In_1681,In_1516);
nor U373 (N_373,In_507,In_1753);
and U374 (N_374,In_637,In_1664);
nand U375 (N_375,In_1875,In_912);
or U376 (N_376,In_1711,In_1830);
nand U377 (N_377,In_888,In_1170);
and U378 (N_378,In_719,In_1425);
and U379 (N_379,In_808,In_1113);
nand U380 (N_380,In_600,In_228);
and U381 (N_381,In_448,In_974);
or U382 (N_382,In_374,In_446);
xor U383 (N_383,In_449,In_222);
or U384 (N_384,In_748,In_780);
xnor U385 (N_385,In_811,In_484);
nor U386 (N_386,In_18,In_925);
and U387 (N_387,In_1886,In_411);
and U388 (N_388,In_325,In_1995);
xor U389 (N_389,In_1231,In_384);
nor U390 (N_390,In_1975,In_605);
and U391 (N_391,In_1815,In_1862);
nand U392 (N_392,In_1365,In_235);
nor U393 (N_393,In_1644,In_1698);
nand U394 (N_394,In_100,In_412);
nor U395 (N_395,In_1002,In_608);
and U396 (N_396,In_1173,In_730);
nor U397 (N_397,In_82,In_1268);
nand U398 (N_398,In_287,In_119);
nor U399 (N_399,In_8,In_26);
nor U400 (N_400,In_1607,In_495);
nor U401 (N_401,In_900,In_1934);
nand U402 (N_402,In_1158,In_993);
nand U403 (N_403,In_1480,In_973);
xnor U404 (N_404,In_220,In_1852);
and U405 (N_405,In_1900,In_728);
or U406 (N_406,In_1531,In_1728);
or U407 (N_407,In_758,In_854);
and U408 (N_408,In_1983,In_969);
nand U409 (N_409,In_1368,In_320);
or U410 (N_410,In_1971,In_1569);
nor U411 (N_411,In_83,In_1782);
nor U412 (N_412,In_960,In_945);
xor U413 (N_413,In_1310,In_1122);
or U414 (N_414,In_1015,In_170);
nand U415 (N_415,In_1086,In_1338);
nand U416 (N_416,In_364,In_1675);
or U417 (N_417,In_934,In_263);
and U418 (N_418,In_1889,In_442);
or U419 (N_419,In_1979,In_1481);
and U420 (N_420,In_1407,In_1505);
xnor U421 (N_421,In_686,In_162);
nand U422 (N_422,In_1334,In_178);
and U423 (N_423,In_607,In_1000);
nand U424 (N_424,In_1720,In_143);
nor U425 (N_425,In_768,In_1609);
nand U426 (N_426,In_1423,In_452);
nand U427 (N_427,In_614,In_86);
nand U428 (N_428,In_1930,In_1622);
nor U429 (N_429,In_1844,In_941);
xnor U430 (N_430,In_306,In_1627);
xnor U431 (N_431,In_1719,In_842);
xor U432 (N_432,In_1842,In_1943);
or U433 (N_433,In_1094,In_850);
xnor U434 (N_434,In_15,In_1957);
and U435 (N_435,In_1124,In_310);
nand U436 (N_436,In_1792,In_753);
xor U437 (N_437,In_731,In_1466);
nor U438 (N_438,In_682,In_1768);
xnor U439 (N_439,In_1181,In_317);
nand U440 (N_440,In_1970,In_431);
nor U441 (N_441,In_1144,In_409);
nand U442 (N_442,In_771,In_1488);
xnor U443 (N_443,In_293,In_1341);
and U444 (N_444,In_1205,In_1832);
nor U445 (N_445,In_896,In_1410);
or U446 (N_446,In_128,In_1004);
and U447 (N_447,In_1724,In_1345);
nand U448 (N_448,In_584,In_787);
xnor U449 (N_449,In_778,In_1553);
xnor U450 (N_450,In_642,In_1533);
or U451 (N_451,In_1193,In_1212);
xnor U452 (N_452,In_352,In_528);
xnor U453 (N_453,In_362,In_378);
xnor U454 (N_454,In_204,In_126);
or U455 (N_455,In_1899,In_1451);
and U456 (N_456,In_1089,In_457);
nor U457 (N_457,In_1521,In_78);
nand U458 (N_458,In_330,In_1517);
xor U459 (N_459,In_118,In_348);
nor U460 (N_460,In_1377,In_523);
nor U461 (N_461,In_1713,In_526);
and U462 (N_462,In_1873,In_592);
and U463 (N_463,In_492,In_439);
and U464 (N_464,In_821,In_536);
xor U465 (N_465,In_1078,In_219);
and U466 (N_466,In_7,In_1037);
nor U467 (N_467,In_324,In_946);
nand U468 (N_468,In_977,In_173);
and U469 (N_469,In_1992,In_171);
nor U470 (N_470,In_980,In_1898);
nor U471 (N_471,In_453,In_136);
or U472 (N_472,In_1115,In_1233);
and U473 (N_473,In_1288,In_355);
or U474 (N_474,In_1655,In_866);
or U475 (N_475,In_1399,In_148);
and U476 (N_476,In_878,In_426);
nand U477 (N_477,In_702,In_985);
or U478 (N_478,In_1408,In_472);
nor U479 (N_479,In_1079,In_1312);
or U480 (N_480,In_1806,In_1819);
nor U481 (N_481,In_1691,In_1814);
nor U482 (N_482,In_1651,In_1436);
nor U483 (N_483,In_764,In_357);
and U484 (N_484,In_1428,In_147);
or U485 (N_485,In_326,In_1459);
nor U486 (N_486,In_1149,In_1010);
and U487 (N_487,In_1121,In_552);
nand U488 (N_488,In_513,In_1011);
nor U489 (N_489,In_93,In_96);
or U490 (N_490,In_1198,In_1512);
or U491 (N_491,In_1236,In_505);
nor U492 (N_492,In_1318,In_1461);
nor U493 (N_493,In_305,In_590);
or U494 (N_494,In_534,In_1163);
xor U495 (N_495,In_1893,In_1932);
and U496 (N_496,In_583,In_621);
nor U497 (N_497,In_1098,In_254);
nand U498 (N_498,In_1135,In_1697);
and U499 (N_499,In_130,In_1319);
nand U500 (N_500,In_836,In_149);
and U501 (N_501,In_1468,In_1476);
and U502 (N_502,In_1358,In_1350);
xnor U503 (N_503,In_467,In_1213);
nor U504 (N_504,In_1847,In_185);
nor U505 (N_505,In_1211,In_894);
xor U506 (N_506,In_1006,In_1393);
xor U507 (N_507,In_1257,In_542);
xor U508 (N_508,In_1239,In_400);
or U509 (N_509,In_115,In_233);
and U510 (N_510,In_616,In_1159);
or U511 (N_511,In_1048,In_1264);
nand U512 (N_512,In_1575,In_103);
or U513 (N_513,In_1058,In_1835);
nor U514 (N_514,In_720,In_601);
and U515 (N_515,In_755,In_582);
and U516 (N_516,In_665,In_1940);
xnor U517 (N_517,In_1333,In_1993);
and U518 (N_518,In_625,In_1710);
or U519 (N_519,In_403,In_1255);
and U520 (N_520,In_445,In_6);
and U521 (N_521,In_1737,In_786);
nor U522 (N_522,In_1848,In_1250);
nand U523 (N_523,In_830,In_1696);
or U524 (N_524,In_1758,In_1999);
nor U525 (N_525,In_585,In_760);
and U526 (N_526,In_1412,In_1190);
xor U527 (N_527,In_1560,In_885);
and U528 (N_528,In_978,In_775);
and U529 (N_529,In_824,In_1489);
or U530 (N_530,In_1034,In_1095);
and U531 (N_531,In_1339,In_1111);
or U532 (N_532,In_1019,In_1262);
and U533 (N_533,In_3,In_1546);
nand U534 (N_534,In_460,In_395);
or U535 (N_535,In_1171,In_211);
nand U536 (N_536,In_987,In_465);
xor U537 (N_537,In_1662,In_1532);
or U538 (N_538,In_1692,In_1117);
nor U539 (N_539,In_1611,In_991);
nand U540 (N_540,In_658,In_270);
nand U541 (N_541,In_1554,In_1356);
nand U542 (N_542,In_1801,In_1242);
xor U543 (N_543,In_654,In_1787);
and U544 (N_544,In_909,In_1021);
nand U545 (N_545,In_1901,In_1615);
or U546 (N_546,In_927,In_289);
or U547 (N_547,In_1766,In_740);
xnor U548 (N_548,In_586,In_882);
xnor U549 (N_549,In_1260,In_595);
nand U550 (N_550,In_20,In_166);
and U551 (N_551,In_329,In_458);
xnor U552 (N_552,In_660,In_1156);
or U553 (N_553,In_164,In_797);
nor U554 (N_554,In_1297,In_1861);
xnor U555 (N_555,In_701,In_1663);
nor U556 (N_556,In_765,In_42);
nor U557 (N_557,In_1379,In_976);
nand U558 (N_558,In_560,In_802);
nand U559 (N_559,In_917,In_1220);
nor U560 (N_560,In_5,In_1439);
or U561 (N_561,In_628,In_1080);
and U562 (N_562,In_1314,In_1321);
and U563 (N_563,In_1182,In_1595);
and U564 (N_564,In_874,In_1503);
and U565 (N_565,In_1103,In_1406);
nand U566 (N_566,In_1496,In_870);
or U567 (N_567,In_541,In_1224);
xor U568 (N_568,In_1424,In_957);
or U569 (N_569,In_1805,In_1869);
nor U570 (N_570,In_1473,In_929);
nand U571 (N_571,In_98,In_1404);
or U572 (N_572,In_1036,In_1536);
xor U573 (N_573,In_1206,In_1690);
or U574 (N_574,In_618,In_1053);
nor U575 (N_575,In_746,In_1279);
nand U576 (N_576,In_1162,In_425);
and U577 (N_577,In_1583,In_1876);
and U578 (N_578,In_1133,In_680);
xor U579 (N_579,In_1396,In_249);
or U580 (N_580,In_867,In_1172);
and U581 (N_581,In_831,In_644);
xor U582 (N_582,In_294,In_1132);
and U583 (N_583,In_1059,In_952);
xor U584 (N_584,In_1160,In_217);
or U585 (N_585,In_884,In_1817);
and U586 (N_586,In_1445,In_1874);
or U587 (N_587,In_766,In_1693);
and U588 (N_588,In_1714,In_135);
xor U589 (N_589,In_779,In_664);
nor U590 (N_590,In_790,In_1230);
nand U591 (N_591,In_524,In_537);
nand U592 (N_592,In_373,In_1139);
and U593 (N_593,In_1269,In_51);
nand U594 (N_594,In_1065,In_1769);
and U595 (N_595,In_1028,In_923);
or U596 (N_596,In_1559,In_44);
nor U597 (N_597,In_159,In_1499);
xor U598 (N_598,In_213,In_1154);
xor U599 (N_599,In_88,In_494);
nor U600 (N_600,In_101,In_983);
and U601 (N_601,In_415,In_382);
and U602 (N_602,In_1855,In_716);
nor U603 (N_603,In_769,In_712);
and U604 (N_604,In_1639,In_188);
xnor U605 (N_605,In_256,In_191);
xor U606 (N_606,In_988,In_1478);
and U607 (N_607,In_1718,In_372);
nand U608 (N_608,In_1519,In_1101);
and U609 (N_609,In_490,In_1092);
nor U610 (N_610,In_1383,In_1985);
xor U611 (N_611,In_1434,In_1840);
nor U612 (N_612,In_641,In_891);
or U613 (N_613,In_757,In_207);
xor U614 (N_614,In_501,In_670);
xor U615 (N_615,In_679,In_1757);
and U616 (N_616,In_1809,In_1416);
xor U617 (N_617,In_1504,In_1138);
and U618 (N_618,In_261,In_581);
or U619 (N_619,In_1245,In_182);
nor U620 (N_620,In_1631,In_1557);
and U621 (N_621,In_481,In_1072);
xnor U622 (N_622,In_1403,In_274);
xor U623 (N_623,In_1325,In_1427);
or U624 (N_624,In_283,In_1075);
or U625 (N_625,In_986,In_456);
xnor U626 (N_626,In_331,In_471);
and U627 (N_627,In_414,In_612);
or U628 (N_628,In_1373,In_1327);
or U629 (N_629,In_1826,In_1035);
and U630 (N_630,In_1085,In_1402);
and U631 (N_631,In_578,In_359);
nand U632 (N_632,In_975,In_1301);
nor U633 (N_633,In_916,In_1054);
xnor U634 (N_634,In_1600,In_504);
nand U635 (N_635,In_1549,In_1127);
and U636 (N_636,In_1074,In_563);
or U637 (N_637,In_1329,In_967);
xor U638 (N_638,In_936,In_1868);
nor U639 (N_639,In_1793,In_683);
and U640 (N_640,In_1839,In_942);
xor U641 (N_641,In_1130,In_1811);
or U642 (N_642,In_1204,In_677);
xnor U643 (N_643,In_1936,In_1249);
or U644 (N_644,In_944,In_1668);
or U645 (N_645,In_1040,In_1120);
xor U646 (N_646,In_1490,In_108);
and U647 (N_647,In_312,In_648);
or U648 (N_648,In_1626,In_589);
and U649 (N_649,In_875,In_545);
xor U650 (N_650,In_144,In_685);
nand U651 (N_651,In_131,In_476);
nand U652 (N_652,In_423,In_1166);
nand U653 (N_653,In_1397,In_1910);
or U654 (N_654,In_901,In_1148);
or U655 (N_655,In_1685,In_487);
or U656 (N_656,In_565,In_1147);
or U657 (N_657,In_784,In_54);
xnor U658 (N_658,In_1361,In_90);
and U659 (N_659,In_1764,In_1039);
and U660 (N_660,In_1395,In_1467);
xor U661 (N_661,In_240,In_1902);
and U662 (N_662,In_227,In_947);
nor U663 (N_663,In_931,In_883);
or U664 (N_664,In_772,In_102);
and U665 (N_665,In_1097,In_1150);
and U666 (N_666,In_1068,In_1340);
nand U667 (N_667,In_996,In_1649);
nand U668 (N_668,In_1856,In_65);
or U669 (N_669,In_1702,In_1706);
nor U670 (N_670,In_1194,In_1960);
nor U671 (N_671,In_782,In_1349);
xnor U672 (N_672,In_1493,In_73);
xor U673 (N_673,In_643,In_49);
and U674 (N_674,In_1180,In_1670);
nor U675 (N_675,In_781,In_556);
xnor U676 (N_676,In_1387,In_1332);
nand U677 (N_677,In_1066,In_377);
or U678 (N_678,In_588,In_502);
xor U679 (N_679,In_1596,In_899);
nor U680 (N_680,In_1803,In_1671);
nand U681 (N_681,In_75,In_832);
nor U682 (N_682,In_805,In_63);
or U683 (N_683,In_1430,In_175);
nor U684 (N_684,In_167,In_713);
or U685 (N_685,In_122,In_1555);
and U686 (N_686,In_22,In_72);
nand U687 (N_687,In_1722,In_571);
nand U688 (N_688,In_172,In_14);
xnor U689 (N_689,In_1033,In_691);
nor U690 (N_690,In_61,In_1259);
nand U691 (N_691,In_134,In_935);
and U692 (N_692,In_146,In_39);
nor U693 (N_693,In_1642,In_879);
or U694 (N_694,In_1657,In_1636);
xor U695 (N_695,In_1179,In_309);
and U696 (N_696,In_950,In_1007);
and U697 (N_697,In_709,In_345);
or U698 (N_698,In_1959,In_1);
nor U699 (N_699,In_593,In_184);
and U700 (N_700,In_1479,In_1348);
and U701 (N_701,In_877,In_328);
and U702 (N_702,In_380,In_284);
nand U703 (N_703,In_998,In_1014);
or U704 (N_704,In_1780,In_1522);
nor U705 (N_705,In_706,In_999);
xor U706 (N_706,In_573,In_1772);
nor U707 (N_707,In_1545,In_594);
nor U708 (N_708,In_361,In_408);
nor U709 (N_709,In_696,In_485);
and U710 (N_710,In_1137,In_1846);
or U711 (N_711,In_540,In_1281);
or U712 (N_712,In_1771,In_1565);
and U713 (N_713,In_932,In_1477);
nand U714 (N_714,In_1580,In_1679);
nor U715 (N_715,In_1794,In_435);
and U716 (N_716,In_398,In_462);
and U717 (N_717,In_1485,In_727);
or U718 (N_718,In_405,In_1617);
or U719 (N_719,In_87,In_546);
and U720 (N_720,In_1091,In_1304);
and U721 (N_721,In_1208,In_1660);
xor U722 (N_722,In_371,In_343);
nand U723 (N_723,In_1931,In_1853);
nor U724 (N_724,In_197,In_982);
xor U725 (N_725,In_828,In_1612);
xnor U726 (N_726,In_735,In_28);
nand U727 (N_727,In_190,In_569);
or U728 (N_728,In_214,In_1298);
or U729 (N_729,In_773,In_1326);
nor U730 (N_730,In_1544,In_216);
nor U731 (N_731,In_1012,In_1187);
nor U732 (N_732,In_1183,In_1666);
nor U733 (N_733,In_1984,In_232);
xnor U734 (N_734,In_839,In_1287);
or U735 (N_735,In_438,In_1816);
and U736 (N_736,In_1944,In_1599);
nand U737 (N_737,In_1954,In_1514);
nand U738 (N_738,In_697,In_66);
xnor U739 (N_739,In_323,In_856);
xor U740 (N_740,In_311,In_819);
xor U741 (N_741,In_260,In_1438);
and U742 (N_742,In_667,In_1601);
nor U743 (N_743,In_793,In_266);
nand U744 (N_744,In_1732,In_774);
or U745 (N_745,In_1005,In_402);
or U746 (N_746,In_1023,In_1907);
nor U747 (N_747,In_1444,In_279);
xor U748 (N_748,In_1498,In_275);
and U749 (N_749,In_1151,In_407);
or U750 (N_750,In_704,In_1996);
nand U751 (N_751,In_1538,In_1227);
xnor U752 (N_752,In_1311,In_1912);
xnor U753 (N_753,In_177,In_807);
and U754 (N_754,In_1322,In_1643);
nor U755 (N_755,In_739,In_763);
and U756 (N_756,In_843,In_1419);
and U757 (N_757,In_1197,In_379);
nor U758 (N_758,In_1232,In_928);
nand U759 (N_759,In_796,In_1088);
xor U760 (N_760,In_549,In_1453);
or U761 (N_761,In_1235,In_1405);
nand U762 (N_762,In_1638,In_511);
nor U763 (N_763,In_433,In_710);
xnor U764 (N_764,In_715,In_1013);
nand U765 (N_765,In_699,In_1073);
and U766 (N_766,In_1184,In_230);
or U767 (N_767,In_114,In_1024);
nand U768 (N_768,In_1071,In_16);
nand U769 (N_769,In_1818,In_1293);
or U770 (N_770,In_948,In_1750);
xor U771 (N_771,In_1587,In_1222);
xor U772 (N_772,In_750,In_1878);
nor U773 (N_773,In_399,In_1568);
or U774 (N_774,In_334,In_498);
xnor U775 (N_775,In_356,In_693);
xnor U776 (N_776,In_1723,In_1027);
or U777 (N_777,In_139,In_1605);
xor U778 (N_778,In_229,In_895);
nand U779 (N_779,In_672,In_1759);
nor U780 (N_780,In_277,In_1593);
nor U781 (N_781,In_1689,In_1760);
nand U782 (N_782,In_818,In_1335);
nor U783 (N_783,In_1994,In_1571);
and U784 (N_784,In_598,In_1784);
nor U785 (N_785,In_1083,In_253);
nor U786 (N_786,In_1570,In_1603);
and U787 (N_787,In_25,In_1223);
nor U788 (N_788,In_1215,In_1988);
nand U789 (N_789,In_1800,In_1247);
nand U790 (N_790,In_1896,In_1808);
nand U791 (N_791,In_1572,In_40);
nor U792 (N_792,In_519,In_1217);
nand U793 (N_793,In_1328,In_849);
xnor U794 (N_794,In_370,In_1727);
and U795 (N_795,In_1388,In_308);
or U796 (N_796,In_1976,In_387);
nand U797 (N_797,In_121,In_1926);
and U798 (N_798,In_1355,In_1592);
or U799 (N_799,In_84,In_794);
nor U800 (N_800,In_1064,In_1556);
or U801 (N_801,In_1294,In_889);
nor U802 (N_802,In_12,In_887);
nand U803 (N_803,In_1632,In_919);
and U804 (N_804,In_1829,In_1234);
nor U805 (N_805,In_1836,In_215);
or U806 (N_806,In_1953,In_1067);
nand U807 (N_807,In_1527,In_1110);
nor U808 (N_808,In_1981,In_857);
nor U809 (N_809,In_1659,In_814);
or U810 (N_810,In_186,In_1177);
and U811 (N_811,In_444,In_732);
or U812 (N_812,In_1824,In_1009);
nand U813 (N_813,In_1791,In_675);
and U814 (N_814,In_1307,In_463);
nor U815 (N_815,In_922,In_742);
and U816 (N_816,In_189,In_1789);
or U817 (N_817,In_1841,In_695);
xor U818 (N_818,In_1542,In_1786);
xor U819 (N_819,In_617,In_1972);
or U820 (N_820,In_158,In_1370);
nor U821 (N_821,In_580,In_486);
or U822 (N_822,In_92,In_959);
and U823 (N_823,In_703,In_776);
nand U824 (N_824,In_1854,In_441);
nor U825 (N_825,In_1515,In_1790);
nand U826 (N_826,In_1849,In_961);
xnor U827 (N_827,In_1433,In_759);
nor U828 (N_828,In_1290,In_1918);
nand U829 (N_829,In_1891,In_1997);
or U830 (N_830,In_1508,In_246);
or U831 (N_831,In_689,In_1164);
or U832 (N_832,In_1534,In_1492);
or U833 (N_833,In_1872,In_1380);
nand U834 (N_834,In_1881,In_1246);
or U835 (N_835,In_276,In_1469);
and U836 (N_836,In_550,In_33);
nand U837 (N_837,In_1831,In_785);
nand U838 (N_838,In_1020,In_322);
nor U839 (N_839,In_777,In_1551);
nor U840 (N_840,In_1291,In_1471);
nor U841 (N_841,In_1646,In_1810);
nor U842 (N_842,In_1441,In_1391);
nand U843 (N_843,In_366,In_1389);
or U844 (N_844,In_332,In_561);
and U845 (N_845,In_1273,In_1684);
or U846 (N_846,In_804,In_1153);
nand U847 (N_847,In_156,In_1751);
nand U848 (N_848,In_1437,In_1680);
xnor U849 (N_849,In_1673,In_514);
or U850 (N_850,In_19,In_180);
and U851 (N_851,In_1050,In_1140);
xor U852 (N_852,In_564,In_1877);
nor U853 (N_853,In_1449,In_1629);
nand U854 (N_854,In_892,In_187);
nand U855 (N_855,In_1456,In_1286);
or U856 (N_856,In_1834,In_297);
or U857 (N_857,In_1630,In_640);
or U858 (N_858,In_694,In_635);
nor U859 (N_859,In_46,In_835);
nand U860 (N_860,In_721,In_1186);
and U861 (N_861,In_517,In_1725);
xor U862 (N_862,In_440,In_1447);
nand U863 (N_863,In_673,In_1885);
and U864 (N_864,In_212,In_575);
or U865 (N_865,In_989,In_1443);
nand U866 (N_866,In_1857,In_587);
or U867 (N_867,In_602,In_68);
and U868 (N_868,In_1866,In_109);
nor U869 (N_869,In_1935,In_1802);
or U870 (N_870,In_1949,In_1989);
and U871 (N_871,In_1797,In_1850);
and U872 (N_872,In_241,In_21);
nor U873 (N_873,In_868,In_1077);
nand U874 (N_874,In_1256,In_1202);
nor U875 (N_875,In_225,In_120);
or U876 (N_876,In_1509,In_27);
nor U877 (N_877,In_1761,In_1735);
nand U878 (N_878,In_1966,In_391);
nor U879 (N_879,In_475,In_631);
and U880 (N_880,In_756,In_1871);
nor U881 (N_881,In_1860,In_278);
nor U882 (N_882,In_1650,In_1392);
or U883 (N_883,In_1837,In_558);
or U884 (N_884,In_1411,In_834);
or U885 (N_885,In_531,In_388);
or U886 (N_886,In_1929,In_299);
nor U887 (N_887,In_1661,In_337);
and U888 (N_888,In_1812,In_829);
xor U889 (N_889,In_752,In_515);
or U890 (N_890,In_1280,In_1308);
or U891 (N_891,In_223,In_291);
nor U892 (N_892,In_1754,In_1228);
xnor U893 (N_893,In_1537,In_653);
nor U894 (N_894,In_574,In_846);
nor U895 (N_895,In_708,In_1057);
nand U896 (N_896,In_1360,In_1980);
or U897 (N_897,In_1667,In_1564);
nand U898 (N_898,In_248,In_538);
and U899 (N_899,In_1351,In_603);
or U900 (N_900,In_1998,In_812);
nor U901 (N_901,In_743,In_1905);
or U902 (N_902,In_1225,In_141);
xnor U903 (N_903,In_1457,In_1597);
xor U904 (N_904,In_1973,In_1563);
xnor U905 (N_905,In_259,In_633);
nor U906 (N_906,In_1254,In_1299);
or U907 (N_907,In_907,In_468);
xor U908 (N_908,In_335,In_918);
nand U909 (N_909,In_489,In_681);
and U910 (N_910,In_1721,In_1619);
and U911 (N_911,In_1266,In_1770);
and U912 (N_912,In_319,In_193);
or U913 (N_913,In_1359,In_744);
and U914 (N_914,In_1188,In_913);
xor U915 (N_915,In_464,In_1415);
nor U916 (N_916,In_1354,In_104);
and U917 (N_917,In_1167,In_64);
nor U918 (N_918,In_1470,In_1785);
xor U919 (N_919,In_862,In_296);
xor U920 (N_920,In_199,In_443);
nand U921 (N_921,In_510,In_619);
nor U922 (N_922,In_1051,In_1482);
or U923 (N_923,In_723,In_1562);
nand U924 (N_924,In_651,In_1955);
nand U925 (N_925,In_620,In_963);
or U926 (N_926,In_1665,In_77);
and U927 (N_927,In_420,In_1366);
nor U928 (N_928,In_302,In_1882);
nand U929 (N_929,In_497,In_1969);
and U930 (N_930,In_962,In_920);
nand U931 (N_931,In_956,In_1062);
and U932 (N_932,In_272,In_1289);
or U933 (N_933,In_397,In_567);
and U934 (N_934,In_1574,In_1749);
nor U935 (N_935,In_1096,In_347);
nor U936 (N_936,In_997,In_1730);
and U937 (N_937,In_406,In_1196);
nand U938 (N_938,In_1386,In_1226);
nor U939 (N_939,In_871,In_469);
xnor U940 (N_940,In_482,In_1579);
nand U941 (N_941,In_385,In_762);
and U942 (N_942,In_285,In_4);
nand U943 (N_943,In_1518,In_41);
nor U944 (N_944,In_924,In_271);
or U945 (N_945,In_1320,In_351);
nand U946 (N_946,In_966,In_300);
nand U947 (N_947,In_964,In_1463);
nor U948 (N_948,In_89,In_861);
and U949 (N_949,In_1017,In_717);
or U950 (N_950,In_1744,In_663);
xnor U951 (N_951,In_1708,In_1464);
or U952 (N_952,In_239,In_629);
or U953 (N_953,In_194,In_1591);
nand U954 (N_954,In_823,In_11);
and U955 (N_955,In_201,In_622);
nand U956 (N_956,In_1880,In_890);
nand U957 (N_957,In_1421,In_535);
and U958 (N_958,In_798,In_1982);
nand U959 (N_959,In_365,In_195);
xnor U960 (N_960,In_627,In_1700);
xnor U961 (N_961,In_1748,In_725);
xnor U962 (N_962,In_521,In_1781);
xor U963 (N_963,In_466,In_163);
and U964 (N_964,In_1637,In_799);
xnor U965 (N_965,In_1694,In_827);
nand U966 (N_966,In_1244,In_1043);
nand U967 (N_967,In_1566,In_392);
and U968 (N_968,In_1704,In_1119);
xor U969 (N_969,In_1353,In_1152);
nand U970 (N_970,In_761,In_303);
nor U971 (N_971,In_1736,In_1778);
and U972 (N_972,In_1923,In_968);
nand U973 (N_973,In_1821,In_1798);
nor U974 (N_974,In_1746,In_1775);
and U975 (N_975,In_1475,In_192);
nor U976 (N_976,In_1734,In_97);
xor U977 (N_977,In_24,In_1895);
and U978 (N_978,In_1214,In_10);
nand U979 (N_979,In_1063,In_624);
nor U980 (N_980,In_45,In_615);
or U981 (N_981,In_544,In_639);
nand U982 (N_982,In_1001,In_1046);
xor U983 (N_983,In_1909,In_1705);
or U984 (N_984,In_1168,In_826);
nand U985 (N_985,In_1674,In_646);
nand U986 (N_986,In_1506,In_801);
and U987 (N_987,In_367,In_953);
nor U988 (N_988,In_943,In_979);
or U989 (N_989,In_803,In_910);
xnor U990 (N_990,In_893,In_1550);
nand U991 (N_991,In_105,In_1081);
and U992 (N_992,In_1426,In_570);
and U993 (N_993,In_1958,In_1783);
and U994 (N_994,In_418,In_451);
nand U995 (N_995,In_1331,In_1741);
nor U996 (N_996,In_1313,In_95);
nand U997 (N_997,In_800,In_711);
and U998 (N_998,In_127,In_1928);
xnor U999 (N_999,In_1076,In_678);
and U1000 (N_1000,In_1956,In_214);
nor U1001 (N_1001,In_1607,In_993);
nand U1002 (N_1002,In_307,In_382);
xnor U1003 (N_1003,In_910,In_1293);
or U1004 (N_1004,In_1629,In_586);
xnor U1005 (N_1005,In_8,In_1993);
and U1006 (N_1006,In_494,In_1845);
and U1007 (N_1007,In_70,In_180);
and U1008 (N_1008,In_1633,In_1764);
nor U1009 (N_1009,In_1699,In_1560);
or U1010 (N_1010,In_715,In_461);
or U1011 (N_1011,In_1414,In_1901);
nand U1012 (N_1012,In_1135,In_1024);
and U1013 (N_1013,In_1399,In_1655);
or U1014 (N_1014,In_1529,In_713);
nor U1015 (N_1015,In_1358,In_1609);
nand U1016 (N_1016,In_1548,In_1812);
nor U1017 (N_1017,In_216,In_306);
xor U1018 (N_1018,In_1437,In_781);
or U1019 (N_1019,In_886,In_1723);
and U1020 (N_1020,In_878,In_95);
nand U1021 (N_1021,In_1729,In_1091);
and U1022 (N_1022,In_1052,In_239);
nor U1023 (N_1023,In_701,In_195);
or U1024 (N_1024,In_796,In_1113);
or U1025 (N_1025,In_316,In_1297);
nand U1026 (N_1026,In_892,In_448);
nor U1027 (N_1027,In_1065,In_518);
xnor U1028 (N_1028,In_1547,In_1113);
nand U1029 (N_1029,In_1664,In_1940);
nand U1030 (N_1030,In_579,In_910);
and U1031 (N_1031,In_216,In_1110);
and U1032 (N_1032,In_1761,In_524);
nor U1033 (N_1033,In_292,In_116);
and U1034 (N_1034,In_473,In_868);
nor U1035 (N_1035,In_1327,In_873);
xnor U1036 (N_1036,In_448,In_1311);
or U1037 (N_1037,In_627,In_540);
nand U1038 (N_1038,In_653,In_1229);
or U1039 (N_1039,In_1329,In_259);
or U1040 (N_1040,In_758,In_1117);
nand U1041 (N_1041,In_257,In_1445);
nand U1042 (N_1042,In_1864,In_386);
xnor U1043 (N_1043,In_74,In_78);
and U1044 (N_1044,In_1785,In_768);
xnor U1045 (N_1045,In_1045,In_1525);
or U1046 (N_1046,In_269,In_783);
or U1047 (N_1047,In_1711,In_657);
xor U1048 (N_1048,In_1503,In_716);
xnor U1049 (N_1049,In_1373,In_1358);
or U1050 (N_1050,In_1602,In_830);
xor U1051 (N_1051,In_1622,In_1059);
and U1052 (N_1052,In_1963,In_518);
nor U1053 (N_1053,In_269,In_15);
xor U1054 (N_1054,In_938,In_1182);
nand U1055 (N_1055,In_496,In_1009);
nand U1056 (N_1056,In_677,In_96);
nand U1057 (N_1057,In_1053,In_1265);
nor U1058 (N_1058,In_176,In_33);
and U1059 (N_1059,In_216,In_1633);
nor U1060 (N_1060,In_1374,In_1332);
or U1061 (N_1061,In_1092,In_1117);
nor U1062 (N_1062,In_925,In_1323);
xnor U1063 (N_1063,In_718,In_1620);
or U1064 (N_1064,In_1408,In_760);
and U1065 (N_1065,In_1608,In_592);
nor U1066 (N_1066,In_621,In_540);
xnor U1067 (N_1067,In_1773,In_1178);
or U1068 (N_1068,In_184,In_848);
xnor U1069 (N_1069,In_1159,In_1407);
and U1070 (N_1070,In_743,In_1670);
nor U1071 (N_1071,In_1355,In_451);
nor U1072 (N_1072,In_218,In_1430);
nand U1073 (N_1073,In_1685,In_1850);
xnor U1074 (N_1074,In_736,In_1080);
xor U1075 (N_1075,In_748,In_1207);
nand U1076 (N_1076,In_696,In_967);
nand U1077 (N_1077,In_1302,In_328);
nand U1078 (N_1078,In_1114,In_1456);
and U1079 (N_1079,In_807,In_190);
nor U1080 (N_1080,In_1040,In_1506);
or U1081 (N_1081,In_525,In_726);
nor U1082 (N_1082,In_40,In_590);
nand U1083 (N_1083,In_818,In_730);
nor U1084 (N_1084,In_1160,In_23);
nor U1085 (N_1085,In_540,In_860);
and U1086 (N_1086,In_601,In_434);
nor U1087 (N_1087,In_418,In_1220);
or U1088 (N_1088,In_125,In_1358);
xnor U1089 (N_1089,In_1697,In_98);
nand U1090 (N_1090,In_1891,In_1908);
xnor U1091 (N_1091,In_1696,In_980);
xor U1092 (N_1092,In_633,In_1937);
nand U1093 (N_1093,In_1807,In_1321);
or U1094 (N_1094,In_1875,In_1471);
xor U1095 (N_1095,In_1704,In_531);
nand U1096 (N_1096,In_168,In_677);
xor U1097 (N_1097,In_377,In_1582);
nor U1098 (N_1098,In_146,In_329);
or U1099 (N_1099,In_1151,In_1375);
and U1100 (N_1100,In_1347,In_116);
nand U1101 (N_1101,In_1203,In_1251);
and U1102 (N_1102,In_1920,In_801);
xor U1103 (N_1103,In_1375,In_793);
and U1104 (N_1104,In_243,In_887);
nand U1105 (N_1105,In_123,In_1237);
or U1106 (N_1106,In_1365,In_1464);
and U1107 (N_1107,In_783,In_375);
nand U1108 (N_1108,In_1766,In_1673);
xor U1109 (N_1109,In_262,In_1933);
or U1110 (N_1110,In_115,In_1139);
nand U1111 (N_1111,In_1326,In_310);
and U1112 (N_1112,In_1447,In_1643);
or U1113 (N_1113,In_778,In_1947);
xor U1114 (N_1114,In_1070,In_1333);
xnor U1115 (N_1115,In_1270,In_1490);
or U1116 (N_1116,In_446,In_236);
and U1117 (N_1117,In_388,In_1831);
xor U1118 (N_1118,In_1307,In_922);
or U1119 (N_1119,In_1380,In_1567);
nor U1120 (N_1120,In_1634,In_270);
nor U1121 (N_1121,In_1662,In_1986);
xor U1122 (N_1122,In_19,In_599);
nand U1123 (N_1123,In_1777,In_886);
nand U1124 (N_1124,In_188,In_1324);
nor U1125 (N_1125,In_1180,In_328);
xnor U1126 (N_1126,In_39,In_1234);
xnor U1127 (N_1127,In_1213,In_119);
nand U1128 (N_1128,In_312,In_412);
or U1129 (N_1129,In_1760,In_1959);
nor U1130 (N_1130,In_1822,In_298);
or U1131 (N_1131,In_1427,In_1589);
xor U1132 (N_1132,In_543,In_661);
xnor U1133 (N_1133,In_896,In_954);
xor U1134 (N_1134,In_1247,In_931);
xor U1135 (N_1135,In_653,In_912);
and U1136 (N_1136,In_1708,In_351);
and U1137 (N_1137,In_1835,In_1309);
nand U1138 (N_1138,In_1010,In_1251);
nor U1139 (N_1139,In_574,In_177);
or U1140 (N_1140,In_1464,In_1935);
nor U1141 (N_1141,In_1931,In_1859);
nand U1142 (N_1142,In_1599,In_47);
xnor U1143 (N_1143,In_1050,In_1803);
nor U1144 (N_1144,In_973,In_672);
or U1145 (N_1145,In_698,In_1868);
and U1146 (N_1146,In_586,In_1588);
nand U1147 (N_1147,In_821,In_213);
and U1148 (N_1148,In_338,In_49);
nand U1149 (N_1149,In_1542,In_925);
nor U1150 (N_1150,In_1095,In_643);
nor U1151 (N_1151,In_1118,In_1467);
xor U1152 (N_1152,In_1208,In_280);
or U1153 (N_1153,In_557,In_1982);
and U1154 (N_1154,In_1243,In_520);
xor U1155 (N_1155,In_1248,In_1474);
or U1156 (N_1156,In_864,In_559);
nand U1157 (N_1157,In_1256,In_9);
and U1158 (N_1158,In_1108,In_713);
nand U1159 (N_1159,In_66,In_814);
nand U1160 (N_1160,In_1445,In_235);
nand U1161 (N_1161,In_1915,In_47);
xnor U1162 (N_1162,In_189,In_1503);
xor U1163 (N_1163,In_1463,In_73);
nor U1164 (N_1164,In_1517,In_1278);
nand U1165 (N_1165,In_344,In_845);
or U1166 (N_1166,In_47,In_141);
xnor U1167 (N_1167,In_192,In_790);
or U1168 (N_1168,In_494,In_1018);
or U1169 (N_1169,In_409,In_167);
xor U1170 (N_1170,In_568,In_1304);
and U1171 (N_1171,In_987,In_995);
xor U1172 (N_1172,In_771,In_1405);
xor U1173 (N_1173,In_960,In_89);
or U1174 (N_1174,In_1777,In_359);
and U1175 (N_1175,In_218,In_180);
nor U1176 (N_1176,In_1214,In_919);
nor U1177 (N_1177,In_1038,In_957);
xnor U1178 (N_1178,In_1315,In_916);
nor U1179 (N_1179,In_700,In_1593);
nor U1180 (N_1180,In_1405,In_1323);
nand U1181 (N_1181,In_1084,In_720);
nand U1182 (N_1182,In_1496,In_106);
nor U1183 (N_1183,In_122,In_1663);
nor U1184 (N_1184,In_1552,In_1923);
nand U1185 (N_1185,In_1127,In_1210);
xor U1186 (N_1186,In_1635,In_1245);
nor U1187 (N_1187,In_373,In_274);
nand U1188 (N_1188,In_92,In_886);
and U1189 (N_1189,In_375,In_847);
or U1190 (N_1190,In_25,In_655);
nand U1191 (N_1191,In_1853,In_1630);
nor U1192 (N_1192,In_715,In_593);
nand U1193 (N_1193,In_974,In_1400);
nor U1194 (N_1194,In_280,In_796);
nor U1195 (N_1195,In_1602,In_84);
nor U1196 (N_1196,In_496,In_615);
and U1197 (N_1197,In_1918,In_613);
and U1198 (N_1198,In_276,In_1396);
or U1199 (N_1199,In_1517,In_729);
and U1200 (N_1200,In_1872,In_333);
nand U1201 (N_1201,In_1623,In_3);
nand U1202 (N_1202,In_870,In_1266);
and U1203 (N_1203,In_1050,In_1207);
nor U1204 (N_1204,In_87,In_154);
or U1205 (N_1205,In_783,In_416);
xor U1206 (N_1206,In_1138,In_1819);
xor U1207 (N_1207,In_244,In_1938);
xor U1208 (N_1208,In_1124,In_1396);
and U1209 (N_1209,In_438,In_299);
nor U1210 (N_1210,In_1417,In_927);
nor U1211 (N_1211,In_355,In_1685);
or U1212 (N_1212,In_1267,In_1325);
nand U1213 (N_1213,In_1519,In_67);
and U1214 (N_1214,In_586,In_1665);
or U1215 (N_1215,In_697,In_140);
xor U1216 (N_1216,In_1527,In_125);
nand U1217 (N_1217,In_647,In_996);
and U1218 (N_1218,In_174,In_1094);
xor U1219 (N_1219,In_519,In_168);
xnor U1220 (N_1220,In_227,In_1945);
and U1221 (N_1221,In_1832,In_587);
or U1222 (N_1222,In_1955,In_675);
nand U1223 (N_1223,In_1823,In_800);
xor U1224 (N_1224,In_1635,In_110);
nor U1225 (N_1225,In_1965,In_424);
nor U1226 (N_1226,In_202,In_506);
xor U1227 (N_1227,In_1847,In_431);
and U1228 (N_1228,In_1417,In_82);
nand U1229 (N_1229,In_593,In_69);
and U1230 (N_1230,In_1122,In_1604);
nor U1231 (N_1231,In_1726,In_714);
or U1232 (N_1232,In_529,In_1331);
and U1233 (N_1233,In_1872,In_1613);
or U1234 (N_1234,In_297,In_1230);
nand U1235 (N_1235,In_142,In_1990);
xor U1236 (N_1236,In_1000,In_1394);
nor U1237 (N_1237,In_1424,In_280);
and U1238 (N_1238,In_1928,In_1799);
nor U1239 (N_1239,In_1253,In_284);
nand U1240 (N_1240,In_820,In_1683);
and U1241 (N_1241,In_289,In_618);
xor U1242 (N_1242,In_1377,In_60);
or U1243 (N_1243,In_1939,In_1805);
nor U1244 (N_1244,In_1215,In_766);
nand U1245 (N_1245,In_971,In_874);
nor U1246 (N_1246,In_524,In_811);
and U1247 (N_1247,In_264,In_1147);
and U1248 (N_1248,In_1814,In_499);
xor U1249 (N_1249,In_738,In_1245);
xor U1250 (N_1250,In_137,In_836);
nor U1251 (N_1251,In_998,In_1568);
or U1252 (N_1252,In_866,In_377);
xnor U1253 (N_1253,In_343,In_1521);
nand U1254 (N_1254,In_569,In_1757);
and U1255 (N_1255,In_167,In_308);
nand U1256 (N_1256,In_805,In_583);
and U1257 (N_1257,In_1443,In_1838);
nor U1258 (N_1258,In_618,In_126);
nand U1259 (N_1259,In_1471,In_1701);
or U1260 (N_1260,In_1202,In_660);
nand U1261 (N_1261,In_876,In_811);
and U1262 (N_1262,In_1262,In_841);
nand U1263 (N_1263,In_882,In_499);
nand U1264 (N_1264,In_263,In_1029);
and U1265 (N_1265,In_237,In_114);
nor U1266 (N_1266,In_1901,In_395);
or U1267 (N_1267,In_1438,In_566);
nor U1268 (N_1268,In_397,In_237);
nand U1269 (N_1269,In_734,In_1275);
nand U1270 (N_1270,In_561,In_1077);
and U1271 (N_1271,In_994,In_1319);
or U1272 (N_1272,In_612,In_496);
or U1273 (N_1273,In_1875,In_132);
nand U1274 (N_1274,In_356,In_472);
and U1275 (N_1275,In_1717,In_1330);
nand U1276 (N_1276,In_1291,In_360);
xnor U1277 (N_1277,In_1551,In_771);
or U1278 (N_1278,In_314,In_530);
nand U1279 (N_1279,In_897,In_285);
nor U1280 (N_1280,In_450,In_1976);
xnor U1281 (N_1281,In_684,In_1230);
xor U1282 (N_1282,In_622,In_781);
nor U1283 (N_1283,In_1812,In_1540);
nand U1284 (N_1284,In_952,In_268);
nand U1285 (N_1285,In_1824,In_915);
nand U1286 (N_1286,In_424,In_1952);
nor U1287 (N_1287,In_435,In_491);
and U1288 (N_1288,In_1763,In_279);
nor U1289 (N_1289,In_534,In_896);
or U1290 (N_1290,In_1932,In_368);
nor U1291 (N_1291,In_1739,In_1419);
and U1292 (N_1292,In_1872,In_814);
and U1293 (N_1293,In_1180,In_762);
nand U1294 (N_1294,In_1172,In_789);
nand U1295 (N_1295,In_1687,In_815);
and U1296 (N_1296,In_76,In_1742);
and U1297 (N_1297,In_1550,In_534);
or U1298 (N_1298,In_1248,In_473);
or U1299 (N_1299,In_85,In_538);
and U1300 (N_1300,In_718,In_1884);
nand U1301 (N_1301,In_886,In_283);
nand U1302 (N_1302,In_1918,In_1982);
or U1303 (N_1303,In_540,In_181);
and U1304 (N_1304,In_1290,In_1880);
and U1305 (N_1305,In_950,In_985);
nor U1306 (N_1306,In_878,In_1001);
and U1307 (N_1307,In_289,In_1537);
xor U1308 (N_1308,In_791,In_1108);
nor U1309 (N_1309,In_649,In_1515);
and U1310 (N_1310,In_232,In_1546);
nor U1311 (N_1311,In_1387,In_1983);
nor U1312 (N_1312,In_84,In_1873);
nand U1313 (N_1313,In_1997,In_189);
xor U1314 (N_1314,In_1355,In_1192);
nand U1315 (N_1315,In_1306,In_1783);
xor U1316 (N_1316,In_411,In_1183);
nor U1317 (N_1317,In_1978,In_1354);
nand U1318 (N_1318,In_1360,In_689);
nand U1319 (N_1319,In_1959,In_41);
or U1320 (N_1320,In_1771,In_963);
nand U1321 (N_1321,In_537,In_517);
or U1322 (N_1322,In_1013,In_1023);
nand U1323 (N_1323,In_966,In_1619);
and U1324 (N_1324,In_582,In_48);
xnor U1325 (N_1325,In_774,In_1396);
and U1326 (N_1326,In_1963,In_401);
and U1327 (N_1327,In_342,In_1212);
xnor U1328 (N_1328,In_860,In_1770);
xnor U1329 (N_1329,In_1514,In_1145);
nand U1330 (N_1330,In_126,In_392);
nand U1331 (N_1331,In_587,In_1348);
or U1332 (N_1332,In_388,In_365);
or U1333 (N_1333,In_571,In_1146);
or U1334 (N_1334,In_1557,In_287);
nor U1335 (N_1335,In_1135,In_43);
nand U1336 (N_1336,In_1008,In_1557);
xor U1337 (N_1337,In_1380,In_775);
xor U1338 (N_1338,In_1120,In_1465);
nand U1339 (N_1339,In_410,In_1315);
or U1340 (N_1340,In_1256,In_200);
nor U1341 (N_1341,In_1936,In_1557);
nand U1342 (N_1342,In_1095,In_1297);
nor U1343 (N_1343,In_443,In_805);
and U1344 (N_1344,In_1015,In_1467);
or U1345 (N_1345,In_634,In_67);
and U1346 (N_1346,In_221,In_563);
xor U1347 (N_1347,In_1262,In_1650);
nor U1348 (N_1348,In_1594,In_662);
nor U1349 (N_1349,In_962,In_29);
nand U1350 (N_1350,In_1087,In_1084);
nand U1351 (N_1351,In_815,In_4);
xor U1352 (N_1352,In_1543,In_1838);
or U1353 (N_1353,In_918,In_327);
nor U1354 (N_1354,In_1582,In_1828);
xnor U1355 (N_1355,In_1564,In_1515);
and U1356 (N_1356,In_272,In_1113);
and U1357 (N_1357,In_639,In_1828);
or U1358 (N_1358,In_1421,In_1090);
and U1359 (N_1359,In_1533,In_1739);
or U1360 (N_1360,In_111,In_656);
xnor U1361 (N_1361,In_1535,In_1027);
xor U1362 (N_1362,In_1993,In_1293);
nor U1363 (N_1363,In_880,In_1925);
xor U1364 (N_1364,In_1679,In_1434);
or U1365 (N_1365,In_339,In_1162);
nand U1366 (N_1366,In_614,In_1637);
nor U1367 (N_1367,In_550,In_1601);
and U1368 (N_1368,In_16,In_1175);
nand U1369 (N_1369,In_1012,In_1462);
nor U1370 (N_1370,In_1827,In_340);
and U1371 (N_1371,In_411,In_500);
nand U1372 (N_1372,In_403,In_766);
and U1373 (N_1373,In_1585,In_669);
and U1374 (N_1374,In_293,In_1174);
xor U1375 (N_1375,In_515,In_339);
and U1376 (N_1376,In_685,In_922);
nor U1377 (N_1377,In_1528,In_455);
xnor U1378 (N_1378,In_371,In_1942);
and U1379 (N_1379,In_1999,In_31);
or U1380 (N_1380,In_742,In_1244);
or U1381 (N_1381,In_507,In_200);
nand U1382 (N_1382,In_1876,In_1959);
nand U1383 (N_1383,In_7,In_1070);
and U1384 (N_1384,In_1733,In_680);
and U1385 (N_1385,In_1091,In_1370);
or U1386 (N_1386,In_314,In_1666);
or U1387 (N_1387,In_497,In_1813);
xnor U1388 (N_1388,In_1467,In_1793);
and U1389 (N_1389,In_1252,In_1430);
xor U1390 (N_1390,In_721,In_1212);
nor U1391 (N_1391,In_1651,In_369);
nor U1392 (N_1392,In_1893,In_1001);
nand U1393 (N_1393,In_1528,In_1872);
or U1394 (N_1394,In_72,In_1805);
nor U1395 (N_1395,In_1567,In_912);
xor U1396 (N_1396,In_391,In_1570);
and U1397 (N_1397,In_62,In_318);
xnor U1398 (N_1398,In_1942,In_699);
or U1399 (N_1399,In_1307,In_1309);
and U1400 (N_1400,In_1253,In_371);
nor U1401 (N_1401,In_1986,In_1773);
xnor U1402 (N_1402,In_1777,In_1833);
nand U1403 (N_1403,In_1752,In_390);
or U1404 (N_1404,In_521,In_1747);
or U1405 (N_1405,In_754,In_804);
nor U1406 (N_1406,In_514,In_187);
nor U1407 (N_1407,In_1815,In_175);
xnor U1408 (N_1408,In_1281,In_596);
nand U1409 (N_1409,In_988,In_1793);
xnor U1410 (N_1410,In_1605,In_1441);
nor U1411 (N_1411,In_374,In_1652);
or U1412 (N_1412,In_495,In_103);
and U1413 (N_1413,In_489,In_1685);
nand U1414 (N_1414,In_881,In_1992);
nor U1415 (N_1415,In_1562,In_1624);
xor U1416 (N_1416,In_540,In_435);
and U1417 (N_1417,In_684,In_1532);
xor U1418 (N_1418,In_550,In_796);
nor U1419 (N_1419,In_1224,In_122);
or U1420 (N_1420,In_1525,In_1246);
xor U1421 (N_1421,In_1204,In_234);
and U1422 (N_1422,In_1033,In_1672);
nor U1423 (N_1423,In_1042,In_1612);
and U1424 (N_1424,In_1446,In_1377);
nor U1425 (N_1425,In_799,In_1072);
or U1426 (N_1426,In_160,In_1181);
nand U1427 (N_1427,In_825,In_1549);
xnor U1428 (N_1428,In_1430,In_30);
nor U1429 (N_1429,In_335,In_1918);
nor U1430 (N_1430,In_781,In_343);
nor U1431 (N_1431,In_1572,In_1635);
nor U1432 (N_1432,In_1124,In_1423);
or U1433 (N_1433,In_953,In_748);
xor U1434 (N_1434,In_603,In_253);
and U1435 (N_1435,In_605,In_944);
and U1436 (N_1436,In_827,In_125);
xnor U1437 (N_1437,In_624,In_1406);
or U1438 (N_1438,In_963,In_950);
xor U1439 (N_1439,In_1831,In_1413);
xnor U1440 (N_1440,In_1183,In_803);
nand U1441 (N_1441,In_1165,In_1314);
or U1442 (N_1442,In_644,In_249);
or U1443 (N_1443,In_861,In_1626);
or U1444 (N_1444,In_1041,In_1090);
nand U1445 (N_1445,In_1378,In_1940);
nand U1446 (N_1446,In_1691,In_1839);
xnor U1447 (N_1447,In_416,In_1482);
xnor U1448 (N_1448,In_970,In_1422);
xnor U1449 (N_1449,In_75,In_1342);
nor U1450 (N_1450,In_685,In_20);
nand U1451 (N_1451,In_1779,In_398);
or U1452 (N_1452,In_186,In_624);
or U1453 (N_1453,In_400,In_1941);
or U1454 (N_1454,In_1312,In_1684);
nor U1455 (N_1455,In_927,In_346);
xnor U1456 (N_1456,In_1039,In_620);
nor U1457 (N_1457,In_978,In_485);
nand U1458 (N_1458,In_1115,In_896);
or U1459 (N_1459,In_1453,In_403);
nor U1460 (N_1460,In_790,In_1282);
nand U1461 (N_1461,In_749,In_530);
nor U1462 (N_1462,In_528,In_1987);
nor U1463 (N_1463,In_1575,In_1592);
or U1464 (N_1464,In_1536,In_1775);
and U1465 (N_1465,In_1258,In_528);
nand U1466 (N_1466,In_1262,In_1841);
nor U1467 (N_1467,In_1268,In_344);
xnor U1468 (N_1468,In_1261,In_1085);
and U1469 (N_1469,In_37,In_1015);
or U1470 (N_1470,In_269,In_436);
and U1471 (N_1471,In_691,In_409);
xnor U1472 (N_1472,In_1006,In_1365);
and U1473 (N_1473,In_299,In_1544);
xnor U1474 (N_1474,In_1846,In_1132);
nand U1475 (N_1475,In_292,In_1429);
xor U1476 (N_1476,In_1357,In_1212);
and U1477 (N_1477,In_368,In_1795);
nor U1478 (N_1478,In_508,In_496);
xnor U1479 (N_1479,In_336,In_1540);
xnor U1480 (N_1480,In_1465,In_1843);
or U1481 (N_1481,In_444,In_658);
xor U1482 (N_1482,In_1157,In_556);
xor U1483 (N_1483,In_1250,In_1805);
nor U1484 (N_1484,In_1034,In_1116);
nand U1485 (N_1485,In_1089,In_1565);
nand U1486 (N_1486,In_504,In_1992);
and U1487 (N_1487,In_1069,In_1050);
xnor U1488 (N_1488,In_389,In_1996);
nor U1489 (N_1489,In_753,In_1800);
and U1490 (N_1490,In_282,In_1826);
xnor U1491 (N_1491,In_1118,In_1316);
or U1492 (N_1492,In_1545,In_1306);
xnor U1493 (N_1493,In_522,In_857);
xor U1494 (N_1494,In_1230,In_1173);
xor U1495 (N_1495,In_889,In_396);
xnor U1496 (N_1496,In_663,In_575);
and U1497 (N_1497,In_544,In_1474);
nand U1498 (N_1498,In_91,In_1634);
xor U1499 (N_1499,In_1914,In_1989);
nand U1500 (N_1500,In_1533,In_312);
nand U1501 (N_1501,In_808,In_389);
xor U1502 (N_1502,In_578,In_306);
xor U1503 (N_1503,In_975,In_794);
xor U1504 (N_1504,In_1517,In_304);
or U1505 (N_1505,In_1763,In_400);
and U1506 (N_1506,In_899,In_1171);
or U1507 (N_1507,In_671,In_1810);
and U1508 (N_1508,In_1911,In_915);
and U1509 (N_1509,In_202,In_1252);
and U1510 (N_1510,In_732,In_702);
nand U1511 (N_1511,In_1962,In_846);
or U1512 (N_1512,In_1966,In_638);
xnor U1513 (N_1513,In_31,In_1978);
nand U1514 (N_1514,In_325,In_1960);
nor U1515 (N_1515,In_679,In_1416);
and U1516 (N_1516,In_1230,In_442);
nand U1517 (N_1517,In_1673,In_811);
nor U1518 (N_1518,In_1199,In_98);
or U1519 (N_1519,In_724,In_408);
nor U1520 (N_1520,In_813,In_656);
or U1521 (N_1521,In_512,In_1992);
and U1522 (N_1522,In_891,In_1417);
nor U1523 (N_1523,In_180,In_1072);
and U1524 (N_1524,In_138,In_1705);
xnor U1525 (N_1525,In_658,In_945);
xor U1526 (N_1526,In_1827,In_644);
or U1527 (N_1527,In_943,In_1177);
xor U1528 (N_1528,In_1264,In_975);
nand U1529 (N_1529,In_564,In_697);
nand U1530 (N_1530,In_280,In_921);
and U1531 (N_1531,In_1485,In_664);
xor U1532 (N_1532,In_237,In_1425);
nor U1533 (N_1533,In_1385,In_1006);
nand U1534 (N_1534,In_1649,In_1849);
or U1535 (N_1535,In_1608,In_1044);
and U1536 (N_1536,In_1339,In_1463);
nor U1537 (N_1537,In_1156,In_882);
nor U1538 (N_1538,In_1998,In_129);
and U1539 (N_1539,In_1349,In_1446);
or U1540 (N_1540,In_1704,In_1795);
xnor U1541 (N_1541,In_1935,In_1361);
nor U1542 (N_1542,In_1870,In_606);
xor U1543 (N_1543,In_1449,In_1622);
nor U1544 (N_1544,In_1488,In_978);
or U1545 (N_1545,In_1542,In_668);
nor U1546 (N_1546,In_575,In_1874);
xnor U1547 (N_1547,In_499,In_566);
nand U1548 (N_1548,In_852,In_579);
xor U1549 (N_1549,In_563,In_910);
and U1550 (N_1550,In_1054,In_40);
nor U1551 (N_1551,In_642,In_1853);
nor U1552 (N_1552,In_436,In_696);
or U1553 (N_1553,In_1960,In_1475);
nor U1554 (N_1554,In_527,In_1565);
xor U1555 (N_1555,In_186,In_1720);
nand U1556 (N_1556,In_1150,In_1910);
and U1557 (N_1557,In_1224,In_679);
nor U1558 (N_1558,In_372,In_1568);
xnor U1559 (N_1559,In_1201,In_1935);
nor U1560 (N_1560,In_1112,In_196);
nor U1561 (N_1561,In_258,In_1622);
xnor U1562 (N_1562,In_517,In_1572);
or U1563 (N_1563,In_1272,In_43);
nor U1564 (N_1564,In_181,In_343);
or U1565 (N_1565,In_259,In_1583);
and U1566 (N_1566,In_248,In_125);
xor U1567 (N_1567,In_479,In_1781);
nor U1568 (N_1568,In_624,In_806);
xor U1569 (N_1569,In_1526,In_1846);
or U1570 (N_1570,In_1705,In_1910);
and U1571 (N_1571,In_368,In_662);
and U1572 (N_1572,In_536,In_1985);
or U1573 (N_1573,In_642,In_641);
and U1574 (N_1574,In_619,In_446);
or U1575 (N_1575,In_1346,In_964);
and U1576 (N_1576,In_560,In_769);
xor U1577 (N_1577,In_1470,In_1143);
nor U1578 (N_1578,In_605,In_1972);
xnor U1579 (N_1579,In_451,In_18);
xor U1580 (N_1580,In_343,In_735);
and U1581 (N_1581,In_1759,In_812);
or U1582 (N_1582,In_949,In_1667);
and U1583 (N_1583,In_870,In_458);
nor U1584 (N_1584,In_1502,In_598);
or U1585 (N_1585,In_270,In_1711);
nand U1586 (N_1586,In_1485,In_751);
nor U1587 (N_1587,In_1282,In_527);
and U1588 (N_1588,In_1876,In_613);
nor U1589 (N_1589,In_1321,In_555);
xor U1590 (N_1590,In_1219,In_1043);
xnor U1591 (N_1591,In_306,In_1671);
or U1592 (N_1592,In_259,In_1262);
xor U1593 (N_1593,In_654,In_1199);
or U1594 (N_1594,In_1204,In_1644);
and U1595 (N_1595,In_1856,In_649);
nor U1596 (N_1596,In_919,In_651);
and U1597 (N_1597,In_1596,In_1743);
nor U1598 (N_1598,In_527,In_1940);
and U1599 (N_1599,In_377,In_669);
and U1600 (N_1600,In_1897,In_1220);
and U1601 (N_1601,In_1397,In_1667);
and U1602 (N_1602,In_92,In_1507);
or U1603 (N_1603,In_587,In_1694);
and U1604 (N_1604,In_655,In_1333);
and U1605 (N_1605,In_729,In_382);
xnor U1606 (N_1606,In_558,In_593);
or U1607 (N_1607,In_356,In_1284);
and U1608 (N_1608,In_411,In_633);
xnor U1609 (N_1609,In_1245,In_1070);
xnor U1610 (N_1610,In_1189,In_130);
xnor U1611 (N_1611,In_983,In_1683);
xor U1612 (N_1612,In_504,In_230);
nand U1613 (N_1613,In_96,In_1186);
nand U1614 (N_1614,In_991,In_1897);
xor U1615 (N_1615,In_237,In_1893);
nand U1616 (N_1616,In_1713,In_956);
and U1617 (N_1617,In_795,In_201);
or U1618 (N_1618,In_1654,In_201);
nand U1619 (N_1619,In_1431,In_1349);
nand U1620 (N_1620,In_65,In_68);
nor U1621 (N_1621,In_294,In_986);
nand U1622 (N_1622,In_83,In_1046);
or U1623 (N_1623,In_360,In_198);
nor U1624 (N_1624,In_1011,In_895);
and U1625 (N_1625,In_1168,In_1214);
or U1626 (N_1626,In_1706,In_1773);
and U1627 (N_1627,In_121,In_1040);
and U1628 (N_1628,In_1993,In_220);
nand U1629 (N_1629,In_636,In_128);
nand U1630 (N_1630,In_37,In_1382);
nor U1631 (N_1631,In_919,In_452);
nand U1632 (N_1632,In_1668,In_696);
nor U1633 (N_1633,In_1217,In_1318);
or U1634 (N_1634,In_1287,In_1254);
xnor U1635 (N_1635,In_1473,In_1180);
or U1636 (N_1636,In_1787,In_1908);
nor U1637 (N_1637,In_1776,In_163);
or U1638 (N_1638,In_1654,In_1543);
nor U1639 (N_1639,In_610,In_612);
and U1640 (N_1640,In_1682,In_911);
and U1641 (N_1641,In_229,In_1220);
xor U1642 (N_1642,In_863,In_507);
and U1643 (N_1643,In_601,In_733);
or U1644 (N_1644,In_501,In_598);
and U1645 (N_1645,In_1588,In_1894);
and U1646 (N_1646,In_1137,In_432);
or U1647 (N_1647,In_362,In_1700);
xnor U1648 (N_1648,In_1840,In_271);
and U1649 (N_1649,In_158,In_358);
nor U1650 (N_1650,In_965,In_1879);
nand U1651 (N_1651,In_1644,In_914);
and U1652 (N_1652,In_1203,In_750);
xnor U1653 (N_1653,In_503,In_127);
or U1654 (N_1654,In_1658,In_1928);
and U1655 (N_1655,In_353,In_343);
nor U1656 (N_1656,In_1079,In_1711);
or U1657 (N_1657,In_337,In_1249);
nor U1658 (N_1658,In_1185,In_1854);
and U1659 (N_1659,In_545,In_1712);
and U1660 (N_1660,In_598,In_1941);
nand U1661 (N_1661,In_222,In_815);
and U1662 (N_1662,In_1765,In_239);
xor U1663 (N_1663,In_1075,In_1006);
nand U1664 (N_1664,In_1193,In_913);
or U1665 (N_1665,In_1683,In_1283);
or U1666 (N_1666,In_1255,In_1011);
xnor U1667 (N_1667,In_1106,In_71);
nand U1668 (N_1668,In_1560,In_683);
nor U1669 (N_1669,In_398,In_1481);
xor U1670 (N_1670,In_893,In_1873);
nand U1671 (N_1671,In_1168,In_516);
or U1672 (N_1672,In_632,In_1384);
or U1673 (N_1673,In_841,In_1815);
and U1674 (N_1674,In_1788,In_19);
nand U1675 (N_1675,In_146,In_413);
nand U1676 (N_1676,In_1808,In_994);
or U1677 (N_1677,In_1394,In_1146);
nand U1678 (N_1678,In_694,In_1487);
nor U1679 (N_1679,In_1817,In_944);
nor U1680 (N_1680,In_372,In_567);
or U1681 (N_1681,In_523,In_83);
and U1682 (N_1682,In_1897,In_1345);
and U1683 (N_1683,In_753,In_829);
nand U1684 (N_1684,In_56,In_579);
and U1685 (N_1685,In_963,In_429);
nand U1686 (N_1686,In_1151,In_131);
and U1687 (N_1687,In_1289,In_758);
nand U1688 (N_1688,In_1805,In_652);
xor U1689 (N_1689,In_1097,In_858);
nor U1690 (N_1690,In_1570,In_1959);
or U1691 (N_1691,In_93,In_1559);
or U1692 (N_1692,In_22,In_980);
nor U1693 (N_1693,In_1858,In_27);
nor U1694 (N_1694,In_1205,In_12);
nor U1695 (N_1695,In_801,In_1221);
or U1696 (N_1696,In_1601,In_1413);
and U1697 (N_1697,In_53,In_981);
nor U1698 (N_1698,In_800,In_313);
nor U1699 (N_1699,In_1407,In_753);
or U1700 (N_1700,In_215,In_1415);
xnor U1701 (N_1701,In_1230,In_1781);
nand U1702 (N_1702,In_880,In_1239);
or U1703 (N_1703,In_130,In_1081);
nor U1704 (N_1704,In_1952,In_555);
and U1705 (N_1705,In_1692,In_1193);
nand U1706 (N_1706,In_1618,In_1050);
nand U1707 (N_1707,In_404,In_1384);
or U1708 (N_1708,In_1901,In_112);
nand U1709 (N_1709,In_509,In_1579);
xor U1710 (N_1710,In_881,In_1706);
nor U1711 (N_1711,In_4,In_245);
nor U1712 (N_1712,In_246,In_1313);
or U1713 (N_1713,In_209,In_249);
or U1714 (N_1714,In_1750,In_884);
xor U1715 (N_1715,In_966,In_1974);
nor U1716 (N_1716,In_1491,In_39);
and U1717 (N_1717,In_924,In_1041);
nor U1718 (N_1718,In_1198,In_1157);
nor U1719 (N_1719,In_1376,In_839);
and U1720 (N_1720,In_417,In_1229);
and U1721 (N_1721,In_1112,In_1674);
and U1722 (N_1722,In_1444,In_301);
and U1723 (N_1723,In_173,In_1694);
xnor U1724 (N_1724,In_865,In_1190);
and U1725 (N_1725,In_1176,In_761);
nand U1726 (N_1726,In_1424,In_687);
nor U1727 (N_1727,In_60,In_1249);
and U1728 (N_1728,In_1089,In_1221);
nor U1729 (N_1729,In_1629,In_1114);
nor U1730 (N_1730,In_208,In_37);
and U1731 (N_1731,In_1991,In_839);
nand U1732 (N_1732,In_112,In_1487);
or U1733 (N_1733,In_1647,In_1719);
and U1734 (N_1734,In_1125,In_266);
nand U1735 (N_1735,In_722,In_1117);
nand U1736 (N_1736,In_1457,In_1512);
and U1737 (N_1737,In_442,In_351);
and U1738 (N_1738,In_1569,In_1238);
and U1739 (N_1739,In_1941,In_1356);
xnor U1740 (N_1740,In_1888,In_1832);
xnor U1741 (N_1741,In_663,In_1291);
or U1742 (N_1742,In_114,In_1497);
and U1743 (N_1743,In_1021,In_92);
nand U1744 (N_1744,In_1764,In_64);
nor U1745 (N_1745,In_1503,In_85);
or U1746 (N_1746,In_1396,In_55);
nand U1747 (N_1747,In_751,In_1649);
or U1748 (N_1748,In_823,In_706);
or U1749 (N_1749,In_334,In_14);
nor U1750 (N_1750,In_313,In_22);
xnor U1751 (N_1751,In_782,In_389);
or U1752 (N_1752,In_1671,In_1115);
and U1753 (N_1753,In_770,In_273);
xor U1754 (N_1754,In_1450,In_562);
and U1755 (N_1755,In_1428,In_107);
xor U1756 (N_1756,In_686,In_1043);
and U1757 (N_1757,In_848,In_230);
or U1758 (N_1758,In_1396,In_1954);
nand U1759 (N_1759,In_745,In_1673);
and U1760 (N_1760,In_1905,In_1814);
or U1761 (N_1761,In_254,In_416);
nand U1762 (N_1762,In_1536,In_1801);
nor U1763 (N_1763,In_1326,In_1051);
and U1764 (N_1764,In_1762,In_943);
xnor U1765 (N_1765,In_802,In_556);
nand U1766 (N_1766,In_1921,In_1009);
xnor U1767 (N_1767,In_1749,In_1469);
or U1768 (N_1768,In_664,In_1033);
xor U1769 (N_1769,In_1894,In_432);
nand U1770 (N_1770,In_1518,In_1685);
xnor U1771 (N_1771,In_662,In_1801);
or U1772 (N_1772,In_210,In_111);
or U1773 (N_1773,In_1618,In_69);
nand U1774 (N_1774,In_1148,In_618);
nor U1775 (N_1775,In_230,In_144);
or U1776 (N_1776,In_1006,In_40);
and U1777 (N_1777,In_456,In_1264);
nand U1778 (N_1778,In_157,In_858);
or U1779 (N_1779,In_1142,In_1751);
or U1780 (N_1780,In_1892,In_1731);
nor U1781 (N_1781,In_1076,In_258);
and U1782 (N_1782,In_1893,In_717);
xor U1783 (N_1783,In_810,In_1625);
nor U1784 (N_1784,In_1680,In_163);
or U1785 (N_1785,In_397,In_903);
or U1786 (N_1786,In_1561,In_178);
and U1787 (N_1787,In_777,In_1250);
xnor U1788 (N_1788,In_1628,In_1981);
nand U1789 (N_1789,In_990,In_641);
nor U1790 (N_1790,In_1558,In_535);
xor U1791 (N_1791,In_754,In_958);
xnor U1792 (N_1792,In_1917,In_1603);
xor U1793 (N_1793,In_757,In_718);
and U1794 (N_1794,In_1305,In_1422);
nand U1795 (N_1795,In_1649,In_1192);
or U1796 (N_1796,In_1474,In_415);
xnor U1797 (N_1797,In_138,In_1021);
nand U1798 (N_1798,In_1274,In_838);
xor U1799 (N_1799,In_1480,In_279);
nand U1800 (N_1800,In_1524,In_1859);
and U1801 (N_1801,In_887,In_1486);
or U1802 (N_1802,In_1386,In_298);
or U1803 (N_1803,In_937,In_1439);
and U1804 (N_1804,In_407,In_616);
and U1805 (N_1805,In_268,In_1929);
or U1806 (N_1806,In_905,In_362);
or U1807 (N_1807,In_510,In_1485);
xor U1808 (N_1808,In_1186,In_642);
or U1809 (N_1809,In_491,In_522);
nor U1810 (N_1810,In_1687,In_719);
nor U1811 (N_1811,In_1164,In_449);
nand U1812 (N_1812,In_221,In_935);
or U1813 (N_1813,In_958,In_609);
or U1814 (N_1814,In_16,In_521);
or U1815 (N_1815,In_1531,In_128);
nor U1816 (N_1816,In_474,In_931);
nand U1817 (N_1817,In_549,In_1413);
nand U1818 (N_1818,In_273,In_1316);
and U1819 (N_1819,In_408,In_1518);
or U1820 (N_1820,In_1376,In_996);
xnor U1821 (N_1821,In_751,In_1113);
or U1822 (N_1822,In_1137,In_1076);
nand U1823 (N_1823,In_178,In_647);
xnor U1824 (N_1824,In_1712,In_1374);
nand U1825 (N_1825,In_1114,In_1156);
and U1826 (N_1826,In_1035,In_1355);
nand U1827 (N_1827,In_1727,In_1633);
xor U1828 (N_1828,In_1449,In_1921);
or U1829 (N_1829,In_555,In_1865);
or U1830 (N_1830,In_102,In_1165);
xnor U1831 (N_1831,In_300,In_1198);
nand U1832 (N_1832,In_1291,In_195);
nand U1833 (N_1833,In_1896,In_1083);
or U1834 (N_1834,In_1307,In_977);
or U1835 (N_1835,In_210,In_1420);
or U1836 (N_1836,In_1512,In_1422);
nand U1837 (N_1837,In_969,In_1601);
nor U1838 (N_1838,In_1121,In_149);
nand U1839 (N_1839,In_883,In_1708);
xor U1840 (N_1840,In_79,In_545);
nand U1841 (N_1841,In_810,In_1282);
nor U1842 (N_1842,In_1090,In_599);
and U1843 (N_1843,In_928,In_26);
or U1844 (N_1844,In_1757,In_952);
nor U1845 (N_1845,In_229,In_601);
nand U1846 (N_1846,In_332,In_1008);
xnor U1847 (N_1847,In_546,In_657);
nand U1848 (N_1848,In_1022,In_24);
and U1849 (N_1849,In_529,In_129);
nand U1850 (N_1850,In_898,In_1152);
or U1851 (N_1851,In_1981,In_1960);
nor U1852 (N_1852,In_586,In_34);
and U1853 (N_1853,In_12,In_1023);
nor U1854 (N_1854,In_17,In_1823);
nand U1855 (N_1855,In_364,In_511);
or U1856 (N_1856,In_329,In_1119);
or U1857 (N_1857,In_1926,In_555);
nand U1858 (N_1858,In_592,In_804);
or U1859 (N_1859,In_1880,In_1697);
or U1860 (N_1860,In_1063,In_1944);
nand U1861 (N_1861,In_283,In_233);
or U1862 (N_1862,In_1821,In_843);
and U1863 (N_1863,In_60,In_642);
or U1864 (N_1864,In_1925,In_169);
nor U1865 (N_1865,In_980,In_8);
xor U1866 (N_1866,In_1428,In_1214);
or U1867 (N_1867,In_970,In_135);
and U1868 (N_1868,In_551,In_1462);
and U1869 (N_1869,In_1598,In_1399);
nor U1870 (N_1870,In_1800,In_828);
and U1871 (N_1871,In_64,In_1073);
and U1872 (N_1872,In_747,In_104);
nor U1873 (N_1873,In_1854,In_391);
and U1874 (N_1874,In_350,In_1620);
xor U1875 (N_1875,In_1946,In_1930);
nor U1876 (N_1876,In_815,In_1865);
xor U1877 (N_1877,In_1798,In_1118);
and U1878 (N_1878,In_1276,In_1305);
nand U1879 (N_1879,In_1820,In_1756);
or U1880 (N_1880,In_160,In_1696);
and U1881 (N_1881,In_848,In_351);
and U1882 (N_1882,In_1674,In_325);
or U1883 (N_1883,In_856,In_818);
xor U1884 (N_1884,In_324,In_1769);
or U1885 (N_1885,In_31,In_830);
nand U1886 (N_1886,In_1374,In_42);
nor U1887 (N_1887,In_1484,In_469);
nand U1888 (N_1888,In_66,In_268);
or U1889 (N_1889,In_1711,In_1119);
or U1890 (N_1890,In_1592,In_1931);
xnor U1891 (N_1891,In_964,In_946);
xor U1892 (N_1892,In_1433,In_1362);
xnor U1893 (N_1893,In_1288,In_858);
xnor U1894 (N_1894,In_1616,In_1513);
or U1895 (N_1895,In_1973,In_591);
and U1896 (N_1896,In_1638,In_1815);
and U1897 (N_1897,In_1467,In_1306);
nand U1898 (N_1898,In_1833,In_1166);
xnor U1899 (N_1899,In_1946,In_590);
and U1900 (N_1900,In_1863,In_112);
nor U1901 (N_1901,In_846,In_101);
or U1902 (N_1902,In_975,In_1864);
or U1903 (N_1903,In_1882,In_736);
nor U1904 (N_1904,In_1379,In_1008);
nor U1905 (N_1905,In_908,In_721);
xnor U1906 (N_1906,In_1787,In_434);
nand U1907 (N_1907,In_691,In_375);
xnor U1908 (N_1908,In_1929,In_740);
xnor U1909 (N_1909,In_825,In_136);
nor U1910 (N_1910,In_754,In_869);
nand U1911 (N_1911,In_642,In_1655);
xor U1912 (N_1912,In_236,In_545);
xnor U1913 (N_1913,In_296,In_962);
and U1914 (N_1914,In_1548,In_1381);
and U1915 (N_1915,In_1442,In_1689);
xor U1916 (N_1916,In_740,In_1456);
nand U1917 (N_1917,In_1584,In_1638);
xor U1918 (N_1918,In_1707,In_280);
or U1919 (N_1919,In_103,In_1728);
xnor U1920 (N_1920,In_835,In_641);
or U1921 (N_1921,In_1532,In_1350);
xnor U1922 (N_1922,In_828,In_1960);
or U1923 (N_1923,In_481,In_1365);
nor U1924 (N_1924,In_1387,In_1558);
or U1925 (N_1925,In_390,In_1204);
nor U1926 (N_1926,In_317,In_1371);
and U1927 (N_1927,In_736,In_1993);
nor U1928 (N_1928,In_1161,In_1142);
and U1929 (N_1929,In_458,In_1862);
nand U1930 (N_1930,In_1277,In_259);
or U1931 (N_1931,In_817,In_1153);
nand U1932 (N_1932,In_997,In_1477);
or U1933 (N_1933,In_1827,In_1148);
nor U1934 (N_1934,In_968,In_1958);
and U1935 (N_1935,In_63,In_878);
and U1936 (N_1936,In_151,In_1238);
nor U1937 (N_1937,In_667,In_1624);
xnor U1938 (N_1938,In_323,In_1326);
xnor U1939 (N_1939,In_804,In_1194);
xor U1940 (N_1940,In_618,In_1525);
nor U1941 (N_1941,In_619,In_1689);
and U1942 (N_1942,In_1820,In_140);
xnor U1943 (N_1943,In_1347,In_305);
and U1944 (N_1944,In_656,In_1471);
nand U1945 (N_1945,In_297,In_1330);
xor U1946 (N_1946,In_528,In_33);
and U1947 (N_1947,In_335,In_1827);
and U1948 (N_1948,In_917,In_862);
nor U1949 (N_1949,In_256,In_1844);
and U1950 (N_1950,In_628,In_1588);
and U1951 (N_1951,In_720,In_580);
nand U1952 (N_1952,In_1260,In_1483);
or U1953 (N_1953,In_1382,In_295);
nand U1954 (N_1954,In_1699,In_76);
or U1955 (N_1955,In_427,In_358);
and U1956 (N_1956,In_906,In_756);
nand U1957 (N_1957,In_108,In_962);
nand U1958 (N_1958,In_68,In_13);
nand U1959 (N_1959,In_895,In_575);
nand U1960 (N_1960,In_1185,In_881);
or U1961 (N_1961,In_945,In_52);
and U1962 (N_1962,In_1246,In_741);
or U1963 (N_1963,In_93,In_199);
nor U1964 (N_1964,In_1895,In_636);
and U1965 (N_1965,In_579,In_1630);
nor U1966 (N_1966,In_1042,In_1169);
nor U1967 (N_1967,In_1113,In_1177);
nor U1968 (N_1968,In_652,In_359);
nor U1969 (N_1969,In_487,In_6);
nand U1970 (N_1970,In_203,In_1765);
nor U1971 (N_1971,In_1719,In_91);
or U1972 (N_1972,In_1491,In_1091);
nor U1973 (N_1973,In_1423,In_381);
or U1974 (N_1974,In_459,In_1298);
nand U1975 (N_1975,In_1521,In_1703);
nand U1976 (N_1976,In_792,In_526);
nand U1977 (N_1977,In_1718,In_921);
nor U1978 (N_1978,In_1770,In_1587);
and U1979 (N_1979,In_1727,In_491);
nand U1980 (N_1980,In_181,In_254);
nor U1981 (N_1981,In_1644,In_1468);
xnor U1982 (N_1982,In_1671,In_1745);
nand U1983 (N_1983,In_1568,In_1392);
xnor U1984 (N_1984,In_1813,In_192);
nand U1985 (N_1985,In_545,In_167);
nor U1986 (N_1986,In_1611,In_941);
nand U1987 (N_1987,In_1461,In_1872);
and U1988 (N_1988,In_1947,In_1845);
xnor U1989 (N_1989,In_836,In_1734);
nand U1990 (N_1990,In_25,In_1287);
or U1991 (N_1991,In_305,In_147);
xnor U1992 (N_1992,In_597,In_1935);
nand U1993 (N_1993,In_1036,In_181);
or U1994 (N_1994,In_1458,In_1018);
xor U1995 (N_1995,In_1119,In_961);
nor U1996 (N_1996,In_1203,In_1746);
xor U1997 (N_1997,In_931,In_58);
xnor U1998 (N_1998,In_1636,In_835);
xnor U1999 (N_1999,In_185,In_1337);
and U2000 (N_2000,N_564,N_1060);
or U2001 (N_2001,N_197,N_874);
or U2002 (N_2002,N_710,N_1037);
xor U2003 (N_2003,N_1872,N_1260);
and U2004 (N_2004,N_1043,N_1828);
or U2005 (N_2005,N_179,N_512);
or U2006 (N_2006,N_831,N_1875);
or U2007 (N_2007,N_1590,N_305);
or U2008 (N_2008,N_143,N_464);
nor U2009 (N_2009,N_1323,N_1614);
and U2010 (N_2010,N_190,N_766);
xnor U2011 (N_2011,N_642,N_906);
nand U2012 (N_2012,N_291,N_838);
nand U2013 (N_2013,N_819,N_136);
xnor U2014 (N_2014,N_259,N_164);
xnor U2015 (N_2015,N_545,N_873);
and U2016 (N_2016,N_1477,N_1038);
nand U2017 (N_2017,N_165,N_1298);
nand U2018 (N_2018,N_416,N_173);
or U2019 (N_2019,N_1290,N_1336);
nor U2020 (N_2020,N_1543,N_117);
nor U2021 (N_2021,N_1777,N_1107);
nand U2022 (N_2022,N_355,N_567);
and U2023 (N_2023,N_1294,N_1801);
nor U2024 (N_2024,N_296,N_69);
nand U2025 (N_2025,N_1678,N_1272);
nand U2026 (N_2026,N_262,N_1878);
xnor U2027 (N_2027,N_46,N_1132);
xor U2028 (N_2028,N_1669,N_1075);
nand U2029 (N_2029,N_1432,N_1244);
and U2030 (N_2030,N_875,N_1685);
nor U2031 (N_2031,N_1933,N_387);
xnor U2032 (N_2032,N_1149,N_1976);
or U2033 (N_2033,N_514,N_93);
nor U2034 (N_2034,N_1092,N_1708);
xnor U2035 (N_2035,N_243,N_1210);
and U2036 (N_2036,N_188,N_348);
or U2037 (N_2037,N_756,N_771);
nor U2038 (N_2038,N_1276,N_147);
nor U2039 (N_2039,N_1209,N_1994);
and U2040 (N_2040,N_1219,N_636);
nand U2041 (N_2041,N_949,N_985);
nand U2042 (N_2042,N_1482,N_1188);
or U2043 (N_2043,N_1494,N_154);
nand U2044 (N_2044,N_212,N_1212);
and U2045 (N_2045,N_1512,N_1183);
xor U2046 (N_2046,N_1312,N_1196);
nand U2047 (N_2047,N_1844,N_1803);
nor U2048 (N_2048,N_303,N_896);
xnor U2049 (N_2049,N_1481,N_655);
and U2050 (N_2050,N_1966,N_1069);
and U2051 (N_2051,N_1090,N_1837);
nor U2052 (N_2052,N_499,N_658);
or U2053 (N_2053,N_1325,N_1772);
or U2054 (N_2054,N_36,N_1306);
and U2055 (N_2055,N_1560,N_1694);
nand U2056 (N_2056,N_91,N_437);
or U2057 (N_2057,N_1174,N_868);
and U2058 (N_2058,N_552,N_972);
nand U2059 (N_2059,N_1213,N_227);
and U2060 (N_2060,N_1400,N_1808);
nor U2061 (N_2061,N_1378,N_1430);
and U2062 (N_2062,N_556,N_174);
nand U2063 (N_2063,N_1089,N_1029);
and U2064 (N_2064,N_1124,N_1819);
nand U2065 (N_2065,N_384,N_942);
nand U2066 (N_2066,N_1653,N_1176);
nand U2067 (N_2067,N_1216,N_1756);
nor U2068 (N_2068,N_1137,N_358);
and U2069 (N_2069,N_1798,N_1940);
nor U2070 (N_2070,N_269,N_1252);
and U2071 (N_2071,N_915,N_1740);
nand U2072 (N_2072,N_391,N_1867);
nor U2073 (N_2073,N_360,N_1195);
xnor U2074 (N_2074,N_578,N_90);
and U2075 (N_2075,N_721,N_550);
and U2076 (N_2076,N_853,N_1850);
xor U2077 (N_2077,N_943,N_682);
and U2078 (N_2078,N_1690,N_1552);
or U2079 (N_2079,N_687,N_1957);
nand U2080 (N_2080,N_155,N_1319);
or U2081 (N_2081,N_412,N_1473);
or U2082 (N_2082,N_231,N_422);
nand U2083 (N_2083,N_1501,N_901);
or U2084 (N_2084,N_479,N_1185);
nor U2085 (N_2085,N_325,N_169);
nor U2086 (N_2086,N_633,N_38);
or U2087 (N_2087,N_245,N_1833);
nand U2088 (N_2088,N_632,N_373);
and U2089 (N_2089,N_607,N_531);
or U2090 (N_2090,N_1567,N_804);
and U2091 (N_2091,N_1963,N_175);
nand U2092 (N_2092,N_624,N_108);
and U2093 (N_2093,N_1502,N_859);
or U2094 (N_2094,N_1287,N_1486);
nor U2095 (N_2095,N_343,N_835);
or U2096 (N_2096,N_181,N_585);
nor U2097 (N_2097,N_229,N_1579);
nand U2098 (N_2098,N_1734,N_1846);
xor U2099 (N_2099,N_1108,N_1654);
xor U2100 (N_2100,N_442,N_813);
xnor U2101 (N_2101,N_557,N_1585);
and U2102 (N_2102,N_1592,N_614);
or U2103 (N_2103,N_1748,N_501);
xnor U2104 (N_2104,N_1427,N_788);
nor U2105 (N_2105,N_1650,N_1563);
nand U2106 (N_2106,N_581,N_237);
nand U2107 (N_2107,N_64,N_857);
nand U2108 (N_2108,N_297,N_1620);
nor U2109 (N_2109,N_1309,N_1937);
xor U2110 (N_2110,N_18,N_1380);
xnor U2111 (N_2111,N_265,N_573);
nor U2112 (N_2112,N_529,N_1768);
nor U2113 (N_2113,N_1417,N_1376);
nand U2114 (N_2114,N_8,N_1001);
xor U2115 (N_2115,N_605,N_1123);
xnor U2116 (N_2116,N_448,N_1433);
nor U2117 (N_2117,N_638,N_1688);
nor U2118 (N_2118,N_1139,N_309);
nor U2119 (N_2119,N_1628,N_1058);
xor U2120 (N_2120,N_534,N_861);
xnor U2121 (N_2121,N_474,N_1278);
nand U2122 (N_2122,N_1022,N_1337);
or U2123 (N_2123,N_398,N_802);
nor U2124 (N_2124,N_1076,N_698);
and U2125 (N_2125,N_1184,N_958);
or U2126 (N_2126,N_1693,N_1647);
nand U2127 (N_2127,N_508,N_132);
or U2128 (N_2128,N_1364,N_1015);
xnor U2129 (N_2129,N_1515,N_1610);
nand U2130 (N_2130,N_745,N_1944);
nand U2131 (N_2131,N_1436,N_1416);
nand U2132 (N_2132,N_574,N_1282);
nand U2133 (N_2133,N_818,N_648);
nand U2134 (N_2134,N_1351,N_1634);
nor U2135 (N_2135,N_1695,N_1999);
or U2136 (N_2136,N_326,N_664);
and U2137 (N_2137,N_1539,N_484);
nand U2138 (N_2138,N_71,N_1909);
and U2139 (N_2139,N_829,N_718);
nand U2140 (N_2140,N_367,N_456);
xnor U2141 (N_2141,N_1152,N_246);
or U2142 (N_2142,N_752,N_333);
nor U2143 (N_2143,N_238,N_1117);
nand U2144 (N_2144,N_1392,N_1947);
xor U2145 (N_2145,N_667,N_21);
and U2146 (N_2146,N_1659,N_1052);
or U2147 (N_2147,N_1946,N_1091);
nand U2148 (N_2148,N_1084,N_1169);
nor U2149 (N_2149,N_404,N_1266);
and U2150 (N_2150,N_59,N_527);
nand U2151 (N_2151,N_1147,N_1063);
or U2152 (N_2152,N_1381,N_1072);
xor U2153 (N_2153,N_1612,N_150);
or U2154 (N_2154,N_496,N_1607);
nor U2155 (N_2155,N_1326,N_1240);
nor U2156 (N_2156,N_1883,N_386);
or U2157 (N_2157,N_849,N_1549);
xor U2158 (N_2158,N_1071,N_20);
and U2159 (N_2159,N_1913,N_258);
xnor U2160 (N_2160,N_536,N_661);
nand U2161 (N_2161,N_1646,N_869);
xor U2162 (N_2162,N_299,N_1382);
and U2163 (N_2163,N_1227,N_1778);
nand U2164 (N_2164,N_1797,N_1273);
nand U2165 (N_2165,N_1277,N_1100);
nor U2166 (N_2166,N_396,N_1370);
and U2167 (N_2167,N_129,N_172);
or U2168 (N_2168,N_1067,N_344);
xor U2169 (N_2169,N_1877,N_1814);
xor U2170 (N_2170,N_469,N_774);
nor U2171 (N_2171,N_1904,N_1434);
or U2172 (N_2172,N_1042,N_1341);
and U2173 (N_2173,N_1897,N_1645);
or U2174 (N_2174,N_891,N_488);
nand U2175 (N_2175,N_481,N_1223);
or U2176 (N_2176,N_880,N_1489);
nand U2177 (N_2177,N_122,N_425);
xnor U2178 (N_2178,N_1484,N_366);
nor U2179 (N_2179,N_42,N_580);
and U2180 (N_2180,N_579,N_1995);
nand U2181 (N_2181,N_611,N_1225);
and U2182 (N_2182,N_780,N_921);
nand U2183 (N_2183,N_604,N_1179);
and U2184 (N_2184,N_843,N_912);
xor U2185 (N_2185,N_1793,N_860);
or U2186 (N_2186,N_1345,N_1405);
xnor U2187 (N_2187,N_1031,N_250);
and U2188 (N_2188,N_1902,N_961);
nand U2189 (N_2189,N_1702,N_881);
nand U2190 (N_2190,N_544,N_603);
and U2191 (N_2191,N_968,N_458);
nor U2192 (N_2192,N_1622,N_1105);
or U2193 (N_2193,N_220,N_795);
or U2194 (N_2194,N_33,N_428);
and U2195 (N_2195,N_58,N_1411);
xor U2196 (N_2196,N_940,N_183);
nor U2197 (N_2197,N_408,N_1035);
nor U2198 (N_2198,N_1232,N_954);
xor U2199 (N_2199,N_466,N_962);
nand U2200 (N_2200,N_1332,N_855);
nand U2201 (N_2201,N_953,N_463);
and U2202 (N_2202,N_841,N_35);
nand U2203 (N_2203,N_2,N_1507);
nand U2204 (N_2204,N_993,N_39);
and U2205 (N_2205,N_1573,N_739);
nor U2206 (N_2206,N_1488,N_539);
and U2207 (N_2207,N_1941,N_1127);
xor U2208 (N_2208,N_1581,N_960);
or U2209 (N_2209,N_1253,N_1943);
or U2210 (N_2210,N_1204,N_805);
nand U2211 (N_2211,N_1300,N_994);
and U2212 (N_2212,N_984,N_1738);
xnor U2213 (N_2213,N_1633,N_685);
xnor U2214 (N_2214,N_1885,N_992);
xnor U2215 (N_2215,N_289,N_1615);
nor U2216 (N_2216,N_644,N_1821);
nor U2217 (N_2217,N_1193,N_1192);
xnor U2218 (N_2218,N_867,N_1849);
and U2219 (N_2219,N_1865,N_1766);
xor U2220 (N_2220,N_1208,N_279);
nor U2221 (N_2221,N_1722,N_1888);
nand U2222 (N_2222,N_284,N_207);
or U2223 (N_2223,N_1460,N_890);
and U2224 (N_2224,N_1041,N_1156);
nand U2225 (N_2225,N_500,N_1816);
xnor U2226 (N_2226,N_170,N_286);
xnor U2227 (N_2227,N_267,N_918);
and U2228 (N_2228,N_1971,N_421);
xnor U2229 (N_2229,N_1073,N_1536);
nor U2230 (N_2230,N_1180,N_1687);
nand U2231 (N_2231,N_1970,N_290);
and U2232 (N_2232,N_346,N_0);
nor U2233 (N_2233,N_1161,N_145);
nand U2234 (N_2234,N_1544,N_1529);
or U2235 (N_2235,N_569,N_1949);
nor U2236 (N_2236,N_903,N_761);
xnor U2237 (N_2237,N_216,N_318);
nand U2238 (N_2238,N_1742,N_1830);
and U2239 (N_2239,N_1269,N_1407);
nor U2240 (N_2240,N_1039,N_1088);
nor U2241 (N_2241,N_1514,N_602);
and U2242 (N_2242,N_1894,N_528);
or U2243 (N_2243,N_1683,N_472);
nor U2244 (N_2244,N_465,N_25);
and U2245 (N_2245,N_971,N_493);
and U2246 (N_2246,N_72,N_1157);
and U2247 (N_2247,N_1027,N_452);
or U2248 (N_2248,N_1498,N_1613);
xor U2249 (N_2249,N_1542,N_1);
and U2250 (N_2250,N_316,N_506);
nor U2251 (N_2251,N_563,N_734);
nand U2252 (N_2252,N_1985,N_1189);
nand U2253 (N_2253,N_1438,N_1118);
nor U2254 (N_2254,N_314,N_131);
and U2255 (N_2255,N_641,N_877);
or U2256 (N_2256,N_517,N_640);
or U2257 (N_2257,N_225,N_478);
nor U2258 (N_2258,N_242,N_226);
xor U2259 (N_2259,N_1905,N_997);
or U2260 (N_2260,N_213,N_568);
or U2261 (N_2261,N_897,N_619);
and U2262 (N_2262,N_973,N_483);
nand U2263 (N_2263,N_610,N_705);
and U2264 (N_2264,N_120,N_53);
nor U2265 (N_2265,N_1666,N_974);
or U2266 (N_2266,N_356,N_457);
nand U2267 (N_2267,N_1007,N_1931);
nand U2268 (N_2268,N_1595,N_130);
or U2269 (N_2269,N_160,N_783);
or U2270 (N_2270,N_162,N_403);
and U2271 (N_2271,N_1725,N_361);
nor U2272 (N_2272,N_1327,N_178);
or U2273 (N_2273,N_16,N_659);
or U2274 (N_2274,N_983,N_288);
nor U2275 (N_2275,N_1984,N_1357);
nand U2276 (N_2276,N_487,N_228);
and U2277 (N_2277,N_1975,N_647);
nand U2278 (N_2278,N_1737,N_549);
and U2279 (N_2279,N_1239,N_79);
nand U2280 (N_2280,N_864,N_1288);
or U2281 (N_2281,N_1393,N_1608);
nand U2282 (N_2282,N_1900,N_293);
xor U2283 (N_2283,N_998,N_1810);
and U2284 (N_2284,N_47,N_1866);
and U2285 (N_2285,N_1452,N_1248);
nor U2286 (N_2286,N_1827,N_1490);
or U2287 (N_2287,N_945,N_1961);
or U2288 (N_2288,N_68,N_1788);
nand U2289 (N_2289,N_88,N_1371);
and U2290 (N_2290,N_524,N_800);
and U2291 (N_2291,N_1661,N_1085);
nand U2292 (N_2292,N_1377,N_1191);
nand U2293 (N_2293,N_1631,N_1575);
xnor U2294 (N_2294,N_1924,N_824);
nor U2295 (N_2295,N_27,N_1333);
nand U2296 (N_2296,N_833,N_609);
nor U2297 (N_2297,N_1479,N_980);
and U2298 (N_2298,N_1228,N_1714);
nand U2299 (N_2299,N_317,N_438);
nand U2300 (N_2300,N_553,N_1297);
or U2301 (N_2301,N_75,N_1068);
nand U2302 (N_2302,N_1136,N_635);
nor U2303 (N_2303,N_67,N_793);
nand U2304 (N_2304,N_106,N_1116);
nor U2305 (N_2305,N_792,N_1596);
nor U2306 (N_2306,N_1206,N_620);
or U2307 (N_2307,N_436,N_202);
or U2308 (N_2308,N_1112,N_1832);
nand U2309 (N_2309,N_1051,N_1207);
nor U2310 (N_2310,N_1361,N_1550);
nand U2311 (N_2311,N_1648,N_400);
or U2312 (N_2312,N_1780,N_551);
or U2313 (N_2313,N_230,N_822);
or U2314 (N_2314,N_1958,N_751);
and U2315 (N_2315,N_1214,N_1732);
and U2316 (N_2316,N_311,N_917);
and U2317 (N_2317,N_847,N_1135);
nor U2318 (N_2318,N_1884,N_631);
or U2319 (N_2319,N_1403,N_1283);
nor U2320 (N_2320,N_1471,N_1760);
xor U2321 (N_2321,N_617,N_1983);
or U2322 (N_2322,N_1813,N_1665);
or U2323 (N_2323,N_768,N_1491);
and U2324 (N_2324,N_754,N_1762);
or U2325 (N_2325,N_406,N_922);
and U2326 (N_2326,N_336,N_652);
and U2327 (N_2327,N_765,N_1601);
nand U2328 (N_2328,N_1247,N_342);
nand U2329 (N_2329,N_251,N_1243);
nor U2330 (N_2330,N_1449,N_1728);
xor U2331 (N_2331,N_742,N_900);
nor U2332 (N_2332,N_1422,N_345);
nor U2333 (N_2333,N_1083,N_392);
or U2334 (N_2334,N_1518,N_105);
and U2335 (N_2335,N_426,N_1483);
nor U2336 (N_2336,N_304,N_1098);
nand U2337 (N_2337,N_696,N_1321);
nor U2338 (N_2338,N_1673,N_895);
nand U2339 (N_2339,N_292,N_963);
and U2340 (N_2340,N_1824,N_97);
and U2341 (N_2341,N_1811,N_1053);
and U2342 (N_2342,N_1598,N_1868);
xor U2343 (N_2343,N_1997,N_263);
and U2344 (N_2344,N_1437,N_275);
and U2345 (N_2345,N_916,N_60);
xnor U2346 (N_2346,N_1876,N_475);
nand U2347 (N_2347,N_1362,N_975);
nand U2348 (N_2348,N_629,N_1880);
nand U2349 (N_2349,N_1641,N_820);
xnor U2350 (N_2350,N_1159,N_206);
xor U2351 (N_2351,N_882,N_287);
and U2352 (N_2352,N_1274,N_65);
nand U2353 (N_2353,N_920,N_1081);
xnor U2354 (N_2354,N_654,N_399);
xnor U2355 (N_2355,N_594,N_797);
nand U2356 (N_2356,N_144,N_1699);
nand U2357 (N_2357,N_1716,N_1697);
xnor U2358 (N_2358,N_1020,N_844);
and U2359 (N_2359,N_1129,N_1746);
nor U2360 (N_2360,N_1523,N_934);
xnor U2361 (N_2361,N_1735,N_812);
and U2362 (N_2362,N_1205,N_699);
and U2363 (N_2363,N_1701,N_700);
nand U2364 (N_2364,N_10,N_1799);
nand U2365 (N_2365,N_98,N_196);
or U2366 (N_2366,N_608,N_184);
or U2367 (N_2367,N_722,N_334);
or U2368 (N_2368,N_1374,N_414);
and U2369 (N_2369,N_727,N_1532);
and U2370 (N_2370,N_54,N_1925);
xor U2371 (N_2371,N_1354,N_307);
xor U2372 (N_2372,N_1388,N_1700);
nor U2373 (N_2373,N_374,N_1980);
and U2374 (N_2374,N_1328,N_592);
or U2375 (N_2375,N_1487,N_837);
or U2376 (N_2376,N_720,N_755);
nor U2377 (N_2377,N_353,N_424);
nand U2378 (N_2378,N_836,N_757);
or U2379 (N_2379,N_255,N_1887);
xnor U2380 (N_2380,N_743,N_1765);
nor U2381 (N_2381,N_1565,N_716);
nor U2382 (N_2382,N_1676,N_814);
nand U2383 (N_2383,N_410,N_189);
nand U2384 (N_2384,N_1235,N_61);
or U2385 (N_2385,N_401,N_785);
nand U2386 (N_2386,N_124,N_1397);
and U2387 (N_2387,N_1724,N_480);
nand U2388 (N_2388,N_1953,N_1903);
and U2389 (N_2389,N_540,N_1404);
nor U2390 (N_2390,N_429,N_241);
xor U2391 (N_2391,N_1664,N_541);
nor U2392 (N_2392,N_198,N_589);
and U2393 (N_2393,N_1752,N_1704);
xnor U2394 (N_2394,N_477,N_1070);
and U2395 (N_2395,N_236,N_503);
nor U2396 (N_2396,N_639,N_746);
nand U2397 (N_2397,N_1713,N_1093);
and U2398 (N_2398,N_1143,N_146);
and U2399 (N_2399,N_656,N_415);
and U2400 (N_2400,N_1731,N_1082);
xor U2401 (N_2401,N_925,N_977);
nor U2402 (N_2402,N_1292,N_740);
or U2403 (N_2403,N_31,N_468);
and U2404 (N_2404,N_1730,N_1018);
xor U2405 (N_2405,N_956,N_1630);
nor U2406 (N_2406,N_1790,N_1717);
nand U2407 (N_2407,N_1617,N_1591);
nor U2408 (N_2408,N_1006,N_1318);
nor U2409 (N_2409,N_1969,N_234);
nand U2410 (N_2410,N_1453,N_1822);
xor U2411 (N_2411,N_253,N_74);
or U2412 (N_2412,N_865,N_92);
xnor U2413 (N_2413,N_695,N_1265);
or U2414 (N_2414,N_1537,N_1146);
nand U2415 (N_2415,N_908,N_1733);
and U2416 (N_2416,N_913,N_665);
or U2417 (N_2417,N_1144,N_1727);
xnor U2418 (N_2418,N_84,N_959);
nand U2419 (N_2419,N_357,N_876);
nand U2420 (N_2420,N_502,N_1114);
or U2421 (N_2421,N_248,N_1128);
nor U2422 (N_2422,N_1019,N_846);
nor U2423 (N_2423,N_1317,N_1577);
nand U2424 (N_2424,N_1632,N_737);
and U2425 (N_2425,N_601,N_1763);
xor U2426 (N_2426,N_1800,N_1853);
nand U2427 (N_2427,N_615,N_273);
nor U2428 (N_2428,N_1528,N_613);
nand U2429 (N_2429,N_82,N_1588);
nand U2430 (N_2430,N_952,N_1111);
nand U2431 (N_2431,N_4,N_26);
nand U2432 (N_2432,N_856,N_858);
nand U2433 (N_2433,N_1506,N_1133);
or U2434 (N_2434,N_96,N_1719);
or U2435 (N_2435,N_1285,N_1165);
nand U2436 (N_2436,N_156,N_1852);
nand U2437 (N_2437,N_1838,N_526);
or U2438 (N_2438,N_507,N_1442);
nand U2439 (N_2439,N_1597,N_277);
and U2440 (N_2440,N_215,N_914);
xor U2441 (N_2441,N_1757,N_1526);
xnor U2442 (N_2442,N_1175,N_302);
and U2443 (N_2443,N_1505,N_554);
nor U2444 (N_2444,N_1055,N_1246);
nand U2445 (N_2445,N_419,N_1485);
or U2446 (N_2446,N_1275,N_1807);
nor U2447 (N_2447,N_1251,N_708);
nand U2448 (N_2448,N_1930,N_911);
or U2449 (N_2449,N_1825,N_1954);
nand U2450 (N_2450,N_1342,N_467);
nor U2451 (N_2451,N_1950,N_1150);
xnor U2452 (N_2452,N_257,N_219);
nor U2453 (N_2453,N_1166,N_397);
or U2454 (N_2454,N_418,N_1097);
xnor U2455 (N_2455,N_1461,N_1658);
or U2456 (N_2456,N_266,N_902);
nand U2457 (N_2457,N_180,N_1835);
nand U2458 (N_2458,N_320,N_753);
or U2459 (N_2459,N_1548,N_380);
nor U2460 (N_2460,N_577,N_1729);
nand U2461 (N_2461,N_1414,N_80);
nand U2462 (N_2462,N_1681,N_680);
or U2463 (N_2463,N_950,N_142);
xor U2464 (N_2464,N_1406,N_1258);
nand U2465 (N_2465,N_803,N_1519);
xnor U2466 (N_2466,N_1047,N_1675);
nor U2467 (N_2467,N_1064,N_1649);
nor U2468 (N_2468,N_407,N_1353);
nand U2469 (N_2469,N_1776,N_702);
nand U2470 (N_2470,N_133,N_798);
xor U2471 (N_2471,N_56,N_1454);
and U2472 (N_2472,N_1256,N_158);
and U2473 (N_2473,N_1843,N_1497);
and U2474 (N_2474,N_395,N_1257);
and U2475 (N_2475,N_301,N_907);
nor U2476 (N_2476,N_845,N_1138);
nand U2477 (N_2477,N_1308,N_94);
nor U2478 (N_2478,N_649,N_167);
xor U2479 (N_2479,N_350,N_1522);
nand U2480 (N_2480,N_1050,N_651);
nand U2481 (N_2481,N_1032,N_1939);
nand U2482 (N_2482,N_1330,N_1220);
xor U2483 (N_2483,N_1671,N_650);
or U2484 (N_2484,N_280,N_1314);
nand U2485 (N_2485,N_1197,N_55);
or U2486 (N_2486,N_24,N_681);
xnor U2487 (N_2487,N_686,N_128);
and U2488 (N_2488,N_627,N_1535);
and U2489 (N_2489,N_85,N_1839);
nand U2490 (N_2490,N_240,N_730);
nand U2491 (N_2491,N_492,N_497);
and U2492 (N_2492,N_1624,N_460);
xor U2493 (N_2493,N_81,N_417);
nand U2494 (N_2494,N_694,N_1686);
or U2495 (N_2495,N_347,N_930);
xor U2496 (N_2496,N_368,N_1583);
or U2497 (N_2497,N_717,N_208);
nand U2498 (N_2498,N_1492,N_1935);
xnor U2499 (N_2499,N_1462,N_491);
nor U2500 (N_2500,N_1259,N_1024);
nor U2501 (N_2501,N_138,N_177);
and U2502 (N_2502,N_454,N_1164);
nor U2503 (N_2503,N_1831,N_1307);
xor U2504 (N_2504,N_9,N_171);
or U2505 (N_2505,N_1359,N_1652);
xnor U2506 (N_2506,N_151,N_1786);
and U2507 (N_2507,N_741,N_570);
nand U2508 (N_2508,N_1080,N_459);
xor U2509 (N_2509,N_928,N_473);
and U2510 (N_2510,N_1104,N_1315);
and U2511 (N_2511,N_1626,N_893);
and U2512 (N_2512,N_1186,N_1236);
nor U2513 (N_2513,N_1026,N_411);
or U2514 (N_2514,N_1992,N_176);
nor U2515 (N_2515,N_1066,N_308);
nor U2516 (N_2516,N_295,N_1268);
or U2517 (N_2517,N_1245,N_1546);
xnor U2518 (N_2518,N_1304,N_712);
nor U2519 (N_2519,N_1480,N_1785);
and U2520 (N_2520,N_1440,N_1349);
nand U2521 (N_2521,N_1131,N_1516);
xor U2522 (N_2522,N_1079,N_1177);
xnor U2523 (N_2523,N_715,N_596);
and U2524 (N_2524,N_281,N_719);
and U2525 (N_2525,N_1692,N_1603);
and U2526 (N_2526,N_1101,N_1365);
and U2527 (N_2527,N_1769,N_738);
or U2528 (N_2528,N_1540,N_1789);
and U2529 (N_2529,N_1698,N_1200);
nor U2530 (N_2530,N_523,N_22);
xor U2531 (N_2531,N_1815,N_886);
nand U2532 (N_2532,N_331,N_1511);
xor U2533 (N_2533,N_340,N_1812);
nor U2534 (N_2534,N_1625,N_369);
nor U2535 (N_2535,N_828,N_1099);
xor U2536 (N_2536,N_1973,N_1201);
xor U2537 (N_2537,N_1141,N_1974);
nand U2538 (N_2538,N_28,N_1870);
or U2539 (N_2539,N_443,N_375);
nand U2540 (N_2540,N_114,N_815);
xor U2541 (N_2541,N_490,N_938);
xnor U2542 (N_2542,N_1410,N_1711);
nor U2543 (N_2543,N_1238,N_1446);
nor U2544 (N_2544,N_1680,N_510);
xor U2545 (N_2545,N_769,N_12);
nand U2546 (N_2546,N_1102,N_1736);
xnor U2547 (N_2547,N_1920,N_672);
nor U2548 (N_2548,N_990,N_1387);
nor U2549 (N_2549,N_561,N_1305);
and U2550 (N_2550,N_1566,N_809);
xnor U2551 (N_2551,N_1293,N_1412);
nor U2552 (N_2552,N_1572,N_703);
nor U2553 (N_2553,N_1606,N_187);
or U2554 (N_2554,N_970,N_1324);
or U2555 (N_2555,N_182,N_759);
and U2556 (N_2556,N_1656,N_999);
nand U2557 (N_2557,N_283,N_1222);
xor U2558 (N_2558,N_584,N_435);
nand U2559 (N_2559,N_103,N_14);
nor U2560 (N_2560,N_1747,N_1873);
nor U2561 (N_2561,N_1435,N_191);
nand U2562 (N_2562,N_1372,N_486);
and U2563 (N_2563,N_744,N_597);
xnor U2564 (N_2564,N_546,N_1521);
xnor U2565 (N_2565,N_100,N_83);
xnor U2566 (N_2566,N_1425,N_200);
or U2567 (N_2567,N_623,N_306);
or U2568 (N_2568,N_1122,N_668);
nand U2569 (N_2569,N_1034,N_1524);
nand U2570 (N_2570,N_1662,N_1932);
and U2571 (N_2571,N_365,N_1621);
nor U2572 (N_2572,N_626,N_670);
xnor U2573 (N_2573,N_445,N_1331);
nor U2574 (N_2574,N_264,N_957);
or U2575 (N_2575,N_714,N_1923);
nand U2576 (N_2576,N_1919,N_1048);
nand U2577 (N_2577,N_1979,N_89);
and U2578 (N_2578,N_704,N_1784);
or U2579 (N_2579,N_806,N_1423);
or U2580 (N_2580,N_1234,N_244);
nand U2581 (N_2581,N_315,N_919);
and U2582 (N_2582,N_195,N_1025);
and U2583 (N_2583,N_1352,N_834);
xnor U2584 (N_2584,N_1751,N_989);
and U2585 (N_2585,N_1795,N_628);
and U2586 (N_2586,N_731,N_779);
or U2587 (N_2587,N_799,N_1016);
nand U2588 (N_2588,N_379,N_451);
xnor U2589 (N_2589,N_1582,N_1310);
xor U2590 (N_2590,N_1464,N_1908);
nand U2591 (N_2591,N_1569,N_119);
nor U2592 (N_2592,N_1301,N_87);
and U2593 (N_2593,N_256,N_1028);
and U2594 (N_2594,N_1616,N_842);
nor U2595 (N_2595,N_1350,N_327);
or U2596 (N_2596,N_854,N_709);
nor U2597 (N_2597,N_153,N_898);
or U2598 (N_2598,N_1395,N_1030);
xor U2599 (N_2599,N_674,N_450);
or U2600 (N_2600,N_23,N_905);
and U2601 (N_2601,N_1379,N_1960);
and U2602 (N_2602,N_645,N_588);
nand U2603 (N_2603,N_1218,N_723);
and U2604 (N_2604,N_1805,N_1750);
and U2605 (N_2605,N_1509,N_439);
or U2606 (N_2606,N_532,N_1782);
or U2607 (N_2607,N_666,N_107);
or U2608 (N_2608,N_678,N_112);
nor U2609 (N_2609,N_1474,N_747);
or U2610 (N_2610,N_1964,N_560);
nand U2611 (N_2611,N_1928,N_1420);
and U2612 (N_2612,N_542,N_1657);
and U2613 (N_2613,N_1962,N_1000);
nand U2614 (N_2614,N_599,N_1570);
and U2615 (N_2615,N_1600,N_1926);
xnor U2616 (N_2616,N_214,N_1869);
xnor U2617 (N_2617,N_78,N_1527);
nand U2618 (N_2618,N_1428,N_1987);
and U2619 (N_2619,N_1190,N_966);
xor U2620 (N_2620,N_110,N_30);
nor U2621 (N_2621,N_1340,N_444);
nor U2622 (N_2622,N_1443,N_1906);
xor U2623 (N_2623,N_1967,N_104);
and U2624 (N_2624,N_1303,N_1221);
nand U2625 (N_2625,N_773,N_555);
or U2626 (N_2626,N_1401,N_979);
or U2627 (N_2627,N_363,N_364);
or U2628 (N_2628,N_1503,N_185);
nand U2629 (N_2629,N_711,N_113);
and U2630 (N_2630,N_892,N_967);
or U2631 (N_2631,N_1672,N_1916);
nand U2632 (N_2632,N_1231,N_1396);
or U2633 (N_2633,N_1951,N_409);
and U2634 (N_2634,N_118,N_1533);
and U2635 (N_2635,N_1945,N_1242);
xnor U2636 (N_2636,N_352,N_634);
and U2637 (N_2637,N_1755,N_879);
xnor U2638 (N_2638,N_1296,N_1609);
nor U2639 (N_2639,N_1942,N_1637);
nor U2640 (N_2640,N_1989,N_1046);
and U2641 (N_2641,N_261,N_485);
nand U2642 (N_2642,N_372,N_462);
nand U2643 (N_2643,N_1106,N_1119);
nor U2644 (N_2644,N_1074,N_870);
and U2645 (N_2645,N_1517,N_351);
or U2646 (N_2646,N_1571,N_1689);
nor U2647 (N_2647,N_1705,N_894);
nand U2648 (N_2648,N_767,N_1316);
or U2649 (N_2649,N_11,N_1623);
nor U2650 (N_2650,N_1668,N_600);
and U2651 (N_2651,N_270,N_489);
or U2652 (N_2652,N_978,N_1682);
or U2653 (N_2653,N_1530,N_390);
nor U2654 (N_2654,N_1663,N_518);
or U2655 (N_2655,N_1466,N_1578);
and U2656 (N_2656,N_378,N_276);
or U2657 (N_2657,N_1602,N_1774);
or U2658 (N_2658,N_724,N_848);
or U2659 (N_2659,N_1644,N_57);
and U2660 (N_2660,N_127,N_1773);
xnor U2661 (N_2661,N_1710,N_653);
nand U2662 (N_2662,N_1500,N_801);
nand U2663 (N_2663,N_637,N_1142);
xnor U2664 (N_2664,N_504,N_1495);
nor U2665 (N_2665,N_446,N_1450);
and U2666 (N_2666,N_1329,N_498);
or U2667 (N_2667,N_1413,N_1390);
nor U2668 (N_2668,N_1262,N_786);
nor U2669 (N_2669,N_149,N_764);
and U2670 (N_2670,N_1224,N_1547);
nand U2671 (N_2671,N_1599,N_382);
nand U2672 (N_2672,N_547,N_796);
or U2673 (N_2673,N_1399,N_1429);
or U2674 (N_2674,N_1743,N_924);
and U2675 (N_2675,N_1062,N_1130);
xnor U2676 (N_2676,N_1818,N_1295);
nor U2677 (N_2677,N_1154,N_910);
nor U2678 (N_2678,N_1927,N_1834);
nand U2679 (N_2679,N_148,N_337);
nand U2680 (N_2680,N_159,N_1978);
xor U2681 (N_2681,N_1120,N_44);
nor U2682 (N_2682,N_995,N_116);
or U2683 (N_2683,N_1322,N_612);
nand U2684 (N_2684,N_1472,N_1934);
nand U2685 (N_2685,N_1861,N_1982);
xor U2686 (N_2686,N_1467,N_1525);
xnor U2687 (N_2687,N_1968,N_123);
and U2688 (N_2688,N_851,N_1424);
nor U2689 (N_2689,N_37,N_1863);
and U2690 (N_2690,N_1721,N_817);
xnor U2691 (N_2691,N_1642,N_1469);
and U2692 (N_2692,N_324,N_66);
xor U2693 (N_2693,N_850,N_947);
or U2694 (N_2694,N_1643,N_1211);
xor U2695 (N_2695,N_683,N_1611);
xnor U2696 (N_2696,N_1448,N_1504);
xnor U2697 (N_2697,N_1917,N_736);
and U2698 (N_2698,N_449,N_268);
and U2699 (N_2699,N_1783,N_17);
and U2700 (N_2700,N_1289,N_1151);
nor U2701 (N_2701,N_1096,N_663);
and U2702 (N_2702,N_562,N_933);
nor U2703 (N_2703,N_689,N_371);
nor U2704 (N_2704,N_1110,N_199);
nor U2705 (N_2705,N_1299,N_1871);
and U2706 (N_2706,N_1929,N_1796);
xor U2707 (N_2707,N_224,N_1703);
nor U2708 (N_2708,N_1557,N_1667);
nand U2709 (N_2709,N_1054,N_40);
nor U2710 (N_2710,N_1910,N_982);
nor U2711 (N_2711,N_691,N_1094);
xor U2712 (N_2712,N_1558,N_679);
nand U2713 (N_2713,N_1457,N_99);
nand U2714 (N_2714,N_1959,N_1568);
and U2715 (N_2715,N_221,N_1886);
and U2716 (N_2716,N_811,N_1172);
nand U2717 (N_2717,N_781,N_109);
and U2718 (N_2718,N_1023,N_1233);
or U2719 (N_2719,N_1121,N_1520);
or U2720 (N_2720,N_1912,N_1358);
and U2721 (N_2721,N_1826,N_1408);
and U2722 (N_2722,N_1468,N_669);
nand U2723 (N_2723,N_1155,N_1045);
and U2724 (N_2724,N_582,N_1754);
xnor U2725 (N_2725,N_1952,N_951);
xor U2726 (N_2726,N_235,N_808);
and U2727 (N_2727,N_29,N_821);
or U2728 (N_2728,N_51,N_1021);
nand U2729 (N_2729,N_322,N_1078);
or U2730 (N_2730,N_1439,N_1313);
nand U2731 (N_2731,N_1918,N_1881);
and U2732 (N_2732,N_6,N_1168);
and U2733 (N_2733,N_1126,N_252);
nand U2734 (N_2734,N_1263,N_816);
nand U2735 (N_2735,N_420,N_453);
and U2736 (N_2736,N_152,N_1249);
and U2737 (N_2737,N_657,N_1478);
and U2738 (N_2738,N_163,N_52);
nand U2739 (N_2739,N_533,N_271);
nand U2740 (N_2740,N_621,N_1004);
nor U2741 (N_2741,N_1344,N_1840);
nor U2742 (N_2742,N_789,N_1922);
nand U2743 (N_2743,N_937,N_125);
or U2744 (N_2744,N_1555,N_878);
nor U2745 (N_2745,N_1384,N_1421);
nor U2746 (N_2746,N_201,N_247);
nand U2747 (N_2747,N_826,N_1375);
and U2748 (N_2748,N_883,N_1402);
xor U2749 (N_2749,N_976,N_15);
and U2750 (N_2750,N_1574,N_688);
and U2751 (N_2751,N_73,N_1418);
or U2752 (N_2752,N_1911,N_476);
xnor U2753 (N_2753,N_1153,N_1451);
or U2754 (N_2754,N_274,N_1551);
xor U2755 (N_2755,N_482,N_575);
and U2756 (N_2756,N_1764,N_590);
nor U2757 (N_2757,N_775,N_1366);
nor U2758 (N_2758,N_1230,N_1115);
nor U2759 (N_2759,N_209,N_1965);
nand U2760 (N_2760,N_1261,N_1334);
or U2761 (N_2761,N_1874,N_1145);
xnor U2762 (N_2762,N_591,N_986);
or U2763 (N_2763,N_1077,N_1629);
nand U2764 (N_2764,N_1348,N_434);
or U2765 (N_2765,N_1003,N_86);
xor U2766 (N_2766,N_1745,N_1158);
xnor U2767 (N_2767,N_1771,N_1651);
xnor U2768 (N_2768,N_7,N_790);
xnor U2769 (N_2769,N_1363,N_758);
nor U2770 (N_2770,N_1279,N_1707);
nand U2771 (N_2771,N_593,N_885);
or U2772 (N_2772,N_1103,N_749);
or U2773 (N_2773,N_690,N_671);
or U2774 (N_2774,N_260,N_1302);
and U2775 (N_2775,N_565,N_76);
nor U2776 (N_2776,N_1593,N_1194);
nor U2777 (N_2777,N_1709,N_1389);
nand U2778 (N_2778,N_1792,N_1017);
xor U2779 (N_2779,N_310,N_1459);
nand U2780 (N_2780,N_359,N_1531);
nor U2781 (N_2781,N_63,N_1758);
xnor U2782 (N_2782,N_662,N_725);
or U2783 (N_2783,N_140,N_1171);
xor U2784 (N_2784,N_349,N_732);
and U2785 (N_2785,N_1061,N_519);
nand U2786 (N_2786,N_760,N_300);
and U2787 (N_2787,N_1576,N_643);
nor U2788 (N_2788,N_1033,N_385);
and U2789 (N_2789,N_1556,N_249);
and U2790 (N_2790,N_193,N_1005);
nand U2791 (N_2791,N_1271,N_1759);
xor U2792 (N_2792,N_1554,N_381);
xnor U2793 (N_2793,N_946,N_1056);
and U2794 (N_2794,N_991,N_194);
nand U2795 (N_2795,N_1538,N_823);
nor U2796 (N_2796,N_41,N_1972);
nor U2797 (N_2797,N_1040,N_701);
nand U2798 (N_2798,N_1996,N_1320);
or U2799 (N_2799,N_441,N_1691);
xnor U2800 (N_2800,N_1860,N_222);
xnor U2801 (N_2801,N_1011,N_762);
or U2802 (N_2802,N_232,N_1684);
nor U2803 (N_2803,N_505,N_1890);
xnor U2804 (N_2804,N_3,N_328);
nand U2805 (N_2805,N_1936,N_839);
xor U2806 (N_2806,N_1360,N_810);
and U2807 (N_2807,N_1847,N_1604);
nor U2808 (N_2808,N_1049,N_939);
nand U2809 (N_2809,N_1541,N_676);
xor U2810 (N_2810,N_587,N_1109);
or U2811 (N_2811,N_1859,N_137);
nor U2812 (N_2812,N_1013,N_777);
nand U2813 (N_2813,N_427,N_218);
or U2814 (N_2814,N_383,N_1373);
and U2815 (N_2815,N_1002,N_1475);
nor U2816 (N_2816,N_1712,N_1476);
and U2817 (N_2817,N_827,N_1956);
and U2818 (N_2818,N_571,N_389);
and U2819 (N_2819,N_1286,N_825);
or U2820 (N_2820,N_1998,N_941);
xor U2821 (N_2821,N_1057,N_1455);
and U2822 (N_2822,N_1696,N_1586);
or U2823 (N_2823,N_338,N_832);
and U2824 (N_2824,N_576,N_126);
and U2825 (N_2825,N_513,N_1167);
nand U2826 (N_2826,N_1203,N_298);
xor U2827 (N_2827,N_1767,N_852);
and U2828 (N_2828,N_735,N_733);
and U2829 (N_2829,N_1761,N_1343);
and U2830 (N_2830,N_1618,N_1938);
xor U2831 (N_2831,N_559,N_522);
or U2832 (N_2832,N_1896,N_1977);
nor U2833 (N_2833,N_1791,N_566);
nand U2834 (N_2834,N_1841,N_1009);
or U2835 (N_2835,N_1368,N_1889);
nor U2836 (N_2836,N_330,N_1178);
or U2837 (N_2837,N_1419,N_1636);
nor U2838 (N_2838,N_239,N_1202);
nand U2839 (N_2839,N_1802,N_5);
or U2840 (N_2840,N_50,N_1545);
or U2841 (N_2841,N_1836,N_543);
nor U2842 (N_2842,N_139,N_1857);
or U2843 (N_2843,N_1895,N_1605);
or U2844 (N_2844,N_1753,N_48);
and U2845 (N_2845,N_455,N_494);
nand U2846 (N_2846,N_1065,N_630);
xor U2847 (N_2847,N_872,N_34);
nor U2848 (N_2848,N_1993,N_684);
nand U2849 (N_2849,N_728,N_1369);
nand U2850 (N_2850,N_511,N_1638);
nor U2851 (N_2851,N_1990,N_388);
and U2852 (N_2852,N_471,N_1014);
and U2853 (N_2853,N_1858,N_622);
nor U2854 (N_2854,N_1584,N_186);
nand U2855 (N_2855,N_927,N_1655);
nand U2856 (N_2856,N_776,N_440);
nand U2857 (N_2857,N_955,N_1749);
nand U2858 (N_2858,N_1781,N_899);
and U2859 (N_2859,N_996,N_433);
and U2860 (N_2860,N_393,N_413);
xnor U2861 (N_2861,N_530,N_535);
nand U2862 (N_2862,N_470,N_1640);
or U2863 (N_2863,N_19,N_770);
nor U2864 (N_2864,N_1311,N_618);
xnor U2865 (N_2865,N_62,N_1356);
or U2866 (N_2866,N_1346,N_1162);
or U2867 (N_2867,N_447,N_782);
nor U2868 (N_2868,N_1215,N_1893);
or U2869 (N_2869,N_697,N_1465);
nor U2870 (N_2870,N_157,N_1134);
nand U2871 (N_2871,N_1385,N_830);
nor U2872 (N_2872,N_377,N_1639);
and U2873 (N_2873,N_111,N_525);
and U2874 (N_2874,N_763,N_887);
or U2875 (N_2875,N_332,N_729);
or U2876 (N_2876,N_1044,N_932);
nor U2877 (N_2877,N_1988,N_964);
xor U2878 (N_2878,N_866,N_1493);
and U2879 (N_2879,N_1806,N_1415);
nor U2880 (N_2880,N_884,N_1898);
or U2881 (N_2881,N_625,N_1431);
or U2882 (N_2882,N_595,N_1237);
and U2883 (N_2883,N_1899,N_1012);
or U2884 (N_2884,N_965,N_1447);
xnor U2885 (N_2885,N_45,N_1892);
nor U2886 (N_2886,N_168,N_495);
or U2887 (N_2887,N_278,N_313);
nor U2888 (N_2888,N_354,N_1660);
nor U2889 (N_2889,N_516,N_1499);
xnor U2890 (N_2890,N_203,N_1463);
and U2891 (N_2891,N_1008,N_1113);
xnor U2892 (N_2892,N_787,N_1229);
and U2893 (N_2893,N_1087,N_660);
nor U2894 (N_2894,N_1264,N_272);
nand U2895 (N_2895,N_254,N_675);
xnor U2896 (N_2896,N_1848,N_1726);
nor U2897 (N_2897,N_1391,N_537);
xnor U2898 (N_2898,N_115,N_1280);
nand U2899 (N_2899,N_376,N_1804);
nor U2900 (N_2900,N_1744,N_1456);
xnor U2901 (N_2901,N_321,N_223);
nor U2902 (N_2902,N_931,N_1559);
xnor U2903 (N_2903,N_43,N_713);
nor U2904 (N_2904,N_423,N_217);
or U2905 (N_2905,N_1787,N_1794);
or U2906 (N_2906,N_936,N_706);
and U2907 (N_2907,N_969,N_1441);
and U2908 (N_2908,N_616,N_1561);
nand U2909 (N_2909,N_1182,N_192);
xnor U2910 (N_2910,N_294,N_1444);
nand U2911 (N_2911,N_558,N_871);
nor U2912 (N_2912,N_1891,N_1882);
or U2913 (N_2913,N_586,N_402);
xnor U2914 (N_2914,N_141,N_319);
nor U2915 (N_2915,N_926,N_1496);
or U2916 (N_2916,N_1879,N_784);
and U2917 (N_2917,N_1723,N_923);
or U2918 (N_2918,N_101,N_904);
and U2919 (N_2919,N_909,N_772);
nor U2920 (N_2920,N_1255,N_981);
nand U2921 (N_2921,N_1508,N_521);
or U2922 (N_2922,N_1059,N_285);
nor U2923 (N_2923,N_77,N_693);
nor U2924 (N_2924,N_583,N_1635);
nor U2925 (N_2925,N_520,N_987);
xor U2926 (N_2926,N_646,N_1339);
nor U2927 (N_2927,N_1914,N_1820);
nand U2928 (N_2928,N_598,N_461);
or U2929 (N_2929,N_948,N_1338);
xor U2930 (N_2930,N_1470,N_1715);
and U2931 (N_2931,N_1458,N_677);
nor U2932 (N_2932,N_432,N_1706);
nand U2933 (N_2933,N_1809,N_1817);
xor U2934 (N_2934,N_726,N_1854);
nor U2935 (N_2935,N_1986,N_1907);
nand U2936 (N_2936,N_362,N_1739);
or U2937 (N_2937,N_282,N_748);
or U2938 (N_2938,N_1619,N_1627);
and U2939 (N_2939,N_1367,N_1140);
and U2940 (N_2940,N_1187,N_1335);
and U2941 (N_2941,N_134,N_1281);
and U2942 (N_2942,N_161,N_1862);
nand U2943 (N_2943,N_863,N_1445);
or U2944 (N_2944,N_204,N_888);
or U2945 (N_2945,N_1564,N_1741);
nand U2946 (N_2946,N_1291,N_1589);
or U2947 (N_2947,N_1125,N_1855);
nor U2948 (N_2948,N_329,N_13);
xnor U2949 (N_2949,N_1594,N_935);
nor U2950 (N_2950,N_430,N_335);
and U2951 (N_2951,N_862,N_431);
or U2952 (N_2952,N_394,N_1254);
xor U2953 (N_2953,N_889,N_1347);
or U2954 (N_2954,N_1534,N_1241);
or U2955 (N_2955,N_1267,N_929);
nand U2956 (N_2956,N_1181,N_1823);
xor U2957 (N_2957,N_1086,N_1426);
nor U2958 (N_2958,N_1394,N_102);
nand U2959 (N_2959,N_1674,N_1845);
nand U2960 (N_2960,N_944,N_121);
or U2961 (N_2961,N_750,N_312);
or U2962 (N_2962,N_70,N_1553);
or U2963 (N_2963,N_538,N_205);
xor U2964 (N_2964,N_1720,N_1562);
xnor U2965 (N_2965,N_1921,N_1148);
nor U2966 (N_2966,N_1284,N_1409);
nor U2967 (N_2967,N_791,N_1580);
or U2968 (N_2968,N_1160,N_1170);
nor U2969 (N_2969,N_166,N_548);
xor U2970 (N_2970,N_1163,N_32);
nand U2971 (N_2971,N_323,N_1270);
and U2972 (N_2972,N_370,N_339);
nand U2973 (N_2973,N_988,N_211);
and U2974 (N_2974,N_135,N_1250);
nor U2975 (N_2975,N_509,N_807);
and U2976 (N_2976,N_1670,N_1587);
xnor U2977 (N_2977,N_1991,N_1718);
xnor U2978 (N_2978,N_1036,N_794);
or U2979 (N_2979,N_1842,N_233);
or U2980 (N_2980,N_1383,N_1198);
nand U2981 (N_2981,N_1915,N_95);
nand U2982 (N_2982,N_1199,N_707);
xor U2983 (N_2983,N_1829,N_778);
and U2984 (N_2984,N_1513,N_1856);
nand U2985 (N_2985,N_572,N_1679);
or U2986 (N_2986,N_49,N_1010);
and U2987 (N_2987,N_1775,N_1955);
xnor U2988 (N_2988,N_210,N_405);
nor U2989 (N_2989,N_1948,N_1217);
nor U2990 (N_2990,N_1226,N_1173);
or U2991 (N_2991,N_1398,N_1386);
xnor U2992 (N_2992,N_515,N_1864);
nor U2993 (N_2993,N_1779,N_606);
or U2994 (N_2994,N_692,N_341);
xor U2995 (N_2995,N_1981,N_1510);
nand U2996 (N_2996,N_1901,N_1095);
or U2997 (N_2997,N_673,N_1355);
nand U2998 (N_2998,N_1851,N_1770);
or U2999 (N_2999,N_1677,N_840);
and U3000 (N_3000,N_983,N_1080);
and U3001 (N_3001,N_1587,N_194);
and U3002 (N_3002,N_310,N_822);
nand U3003 (N_3003,N_1775,N_1353);
nor U3004 (N_3004,N_1290,N_1820);
nor U3005 (N_3005,N_1493,N_429);
nand U3006 (N_3006,N_1696,N_643);
or U3007 (N_3007,N_1930,N_1713);
xor U3008 (N_3008,N_1880,N_747);
or U3009 (N_3009,N_517,N_1606);
nand U3010 (N_3010,N_1435,N_587);
nor U3011 (N_3011,N_437,N_1672);
and U3012 (N_3012,N_424,N_1369);
xor U3013 (N_3013,N_501,N_1991);
nand U3014 (N_3014,N_1271,N_8);
xnor U3015 (N_3015,N_488,N_797);
xor U3016 (N_3016,N_804,N_1479);
nand U3017 (N_3017,N_100,N_1343);
xnor U3018 (N_3018,N_53,N_1017);
and U3019 (N_3019,N_681,N_1118);
nand U3020 (N_3020,N_494,N_665);
or U3021 (N_3021,N_1941,N_243);
nor U3022 (N_3022,N_106,N_810);
nor U3023 (N_3023,N_1224,N_1006);
nand U3024 (N_3024,N_617,N_1958);
and U3025 (N_3025,N_276,N_483);
nor U3026 (N_3026,N_775,N_524);
or U3027 (N_3027,N_1958,N_733);
and U3028 (N_3028,N_1938,N_209);
or U3029 (N_3029,N_957,N_28);
nor U3030 (N_3030,N_1336,N_13);
or U3031 (N_3031,N_1867,N_1477);
nor U3032 (N_3032,N_1972,N_410);
nor U3033 (N_3033,N_1047,N_1335);
xor U3034 (N_3034,N_1523,N_138);
nor U3035 (N_3035,N_1700,N_1234);
or U3036 (N_3036,N_628,N_203);
nor U3037 (N_3037,N_1046,N_1350);
nor U3038 (N_3038,N_378,N_994);
xnor U3039 (N_3039,N_781,N_1220);
nor U3040 (N_3040,N_585,N_1110);
or U3041 (N_3041,N_787,N_877);
nor U3042 (N_3042,N_1290,N_70);
nor U3043 (N_3043,N_785,N_1746);
and U3044 (N_3044,N_606,N_1912);
xnor U3045 (N_3045,N_1529,N_1480);
or U3046 (N_3046,N_3,N_1984);
xor U3047 (N_3047,N_380,N_452);
nor U3048 (N_3048,N_921,N_585);
or U3049 (N_3049,N_1687,N_1540);
and U3050 (N_3050,N_71,N_1707);
and U3051 (N_3051,N_292,N_1252);
and U3052 (N_3052,N_53,N_833);
xor U3053 (N_3053,N_1622,N_771);
xor U3054 (N_3054,N_982,N_1956);
nor U3055 (N_3055,N_1237,N_556);
nand U3056 (N_3056,N_1686,N_434);
nand U3057 (N_3057,N_1822,N_612);
nor U3058 (N_3058,N_1905,N_381);
xnor U3059 (N_3059,N_1717,N_1566);
nor U3060 (N_3060,N_1907,N_865);
nand U3061 (N_3061,N_1269,N_1129);
nor U3062 (N_3062,N_317,N_989);
or U3063 (N_3063,N_1373,N_1974);
and U3064 (N_3064,N_275,N_420);
nor U3065 (N_3065,N_1582,N_277);
xnor U3066 (N_3066,N_1372,N_1336);
nor U3067 (N_3067,N_247,N_819);
nand U3068 (N_3068,N_1344,N_939);
nor U3069 (N_3069,N_534,N_690);
nand U3070 (N_3070,N_1673,N_1495);
xnor U3071 (N_3071,N_1386,N_1580);
nand U3072 (N_3072,N_977,N_1796);
xnor U3073 (N_3073,N_909,N_678);
xor U3074 (N_3074,N_1585,N_1624);
xor U3075 (N_3075,N_90,N_552);
xnor U3076 (N_3076,N_798,N_511);
xor U3077 (N_3077,N_793,N_1398);
or U3078 (N_3078,N_273,N_1185);
or U3079 (N_3079,N_9,N_1740);
nor U3080 (N_3080,N_1935,N_1517);
xor U3081 (N_3081,N_161,N_1638);
or U3082 (N_3082,N_1355,N_484);
and U3083 (N_3083,N_1870,N_196);
nor U3084 (N_3084,N_347,N_399);
nor U3085 (N_3085,N_1182,N_459);
nor U3086 (N_3086,N_1088,N_442);
nor U3087 (N_3087,N_1437,N_551);
or U3088 (N_3088,N_1,N_947);
nand U3089 (N_3089,N_430,N_278);
or U3090 (N_3090,N_1534,N_570);
nor U3091 (N_3091,N_1480,N_1759);
nor U3092 (N_3092,N_1900,N_1463);
nor U3093 (N_3093,N_850,N_1070);
nor U3094 (N_3094,N_1193,N_75);
nor U3095 (N_3095,N_332,N_1959);
or U3096 (N_3096,N_1681,N_813);
nor U3097 (N_3097,N_858,N_1046);
or U3098 (N_3098,N_222,N_651);
and U3099 (N_3099,N_653,N_413);
xnor U3100 (N_3100,N_1918,N_1739);
xnor U3101 (N_3101,N_1615,N_653);
or U3102 (N_3102,N_936,N_1678);
or U3103 (N_3103,N_1368,N_581);
or U3104 (N_3104,N_1097,N_1782);
nor U3105 (N_3105,N_908,N_1514);
and U3106 (N_3106,N_1710,N_439);
xor U3107 (N_3107,N_358,N_1743);
or U3108 (N_3108,N_1601,N_1559);
nand U3109 (N_3109,N_856,N_1742);
and U3110 (N_3110,N_14,N_1983);
or U3111 (N_3111,N_89,N_1163);
nand U3112 (N_3112,N_1407,N_564);
or U3113 (N_3113,N_1744,N_1064);
or U3114 (N_3114,N_548,N_126);
and U3115 (N_3115,N_513,N_1543);
nor U3116 (N_3116,N_1419,N_1508);
nand U3117 (N_3117,N_1703,N_1453);
nor U3118 (N_3118,N_1681,N_1168);
xnor U3119 (N_3119,N_1068,N_281);
xnor U3120 (N_3120,N_1905,N_749);
nor U3121 (N_3121,N_534,N_47);
nor U3122 (N_3122,N_1214,N_339);
xor U3123 (N_3123,N_1594,N_1972);
nand U3124 (N_3124,N_1861,N_972);
and U3125 (N_3125,N_5,N_1103);
and U3126 (N_3126,N_347,N_693);
nor U3127 (N_3127,N_1990,N_193);
xnor U3128 (N_3128,N_1290,N_1090);
and U3129 (N_3129,N_482,N_599);
xnor U3130 (N_3130,N_657,N_1105);
xor U3131 (N_3131,N_1519,N_1955);
and U3132 (N_3132,N_1380,N_1446);
nor U3133 (N_3133,N_1876,N_1149);
and U3134 (N_3134,N_1843,N_1087);
or U3135 (N_3135,N_1160,N_228);
and U3136 (N_3136,N_1109,N_1029);
and U3137 (N_3137,N_1976,N_256);
and U3138 (N_3138,N_1325,N_600);
or U3139 (N_3139,N_1151,N_1624);
nand U3140 (N_3140,N_1594,N_648);
or U3141 (N_3141,N_344,N_967);
or U3142 (N_3142,N_1705,N_932);
xnor U3143 (N_3143,N_1588,N_881);
and U3144 (N_3144,N_1399,N_4);
xnor U3145 (N_3145,N_103,N_811);
nor U3146 (N_3146,N_750,N_833);
nand U3147 (N_3147,N_1670,N_974);
xor U3148 (N_3148,N_582,N_50);
or U3149 (N_3149,N_1608,N_1583);
nand U3150 (N_3150,N_752,N_1577);
or U3151 (N_3151,N_1384,N_1035);
or U3152 (N_3152,N_1765,N_0);
nor U3153 (N_3153,N_1697,N_1485);
nand U3154 (N_3154,N_1592,N_157);
nor U3155 (N_3155,N_355,N_1496);
nor U3156 (N_3156,N_1372,N_1770);
or U3157 (N_3157,N_1323,N_877);
xor U3158 (N_3158,N_820,N_1681);
xnor U3159 (N_3159,N_1672,N_1691);
and U3160 (N_3160,N_1494,N_1576);
xor U3161 (N_3161,N_778,N_1744);
nand U3162 (N_3162,N_15,N_1756);
nand U3163 (N_3163,N_1443,N_286);
xor U3164 (N_3164,N_235,N_977);
and U3165 (N_3165,N_1879,N_1387);
or U3166 (N_3166,N_1983,N_577);
and U3167 (N_3167,N_650,N_730);
nand U3168 (N_3168,N_72,N_1539);
nand U3169 (N_3169,N_1065,N_704);
nor U3170 (N_3170,N_1911,N_889);
and U3171 (N_3171,N_1041,N_1540);
xnor U3172 (N_3172,N_1466,N_447);
or U3173 (N_3173,N_214,N_324);
and U3174 (N_3174,N_428,N_808);
nor U3175 (N_3175,N_864,N_1668);
nor U3176 (N_3176,N_87,N_542);
nand U3177 (N_3177,N_1932,N_1513);
xnor U3178 (N_3178,N_1937,N_1663);
nand U3179 (N_3179,N_1525,N_928);
nand U3180 (N_3180,N_1812,N_350);
or U3181 (N_3181,N_1595,N_1845);
xnor U3182 (N_3182,N_589,N_108);
xor U3183 (N_3183,N_1186,N_359);
and U3184 (N_3184,N_1695,N_1233);
nand U3185 (N_3185,N_425,N_1908);
and U3186 (N_3186,N_779,N_877);
xnor U3187 (N_3187,N_934,N_722);
nand U3188 (N_3188,N_758,N_725);
or U3189 (N_3189,N_1072,N_1121);
nand U3190 (N_3190,N_14,N_256);
nand U3191 (N_3191,N_1159,N_518);
and U3192 (N_3192,N_1418,N_1331);
and U3193 (N_3193,N_1492,N_484);
and U3194 (N_3194,N_1329,N_1379);
and U3195 (N_3195,N_1236,N_654);
and U3196 (N_3196,N_752,N_1150);
or U3197 (N_3197,N_1904,N_1217);
and U3198 (N_3198,N_1796,N_935);
nand U3199 (N_3199,N_37,N_1026);
and U3200 (N_3200,N_21,N_126);
or U3201 (N_3201,N_718,N_1774);
nor U3202 (N_3202,N_39,N_1722);
nand U3203 (N_3203,N_818,N_1726);
nor U3204 (N_3204,N_393,N_1411);
nand U3205 (N_3205,N_590,N_1937);
nand U3206 (N_3206,N_1572,N_1859);
nand U3207 (N_3207,N_1002,N_9);
or U3208 (N_3208,N_1204,N_336);
xor U3209 (N_3209,N_1401,N_904);
or U3210 (N_3210,N_1845,N_1462);
xnor U3211 (N_3211,N_1967,N_1654);
and U3212 (N_3212,N_469,N_1556);
xor U3213 (N_3213,N_886,N_1686);
nor U3214 (N_3214,N_1895,N_193);
and U3215 (N_3215,N_360,N_325);
and U3216 (N_3216,N_1045,N_1156);
nand U3217 (N_3217,N_79,N_1054);
xnor U3218 (N_3218,N_1567,N_1809);
xor U3219 (N_3219,N_1902,N_535);
nor U3220 (N_3220,N_72,N_1836);
nor U3221 (N_3221,N_1872,N_757);
nand U3222 (N_3222,N_382,N_646);
nand U3223 (N_3223,N_1267,N_670);
nand U3224 (N_3224,N_45,N_642);
and U3225 (N_3225,N_869,N_456);
xor U3226 (N_3226,N_504,N_1646);
or U3227 (N_3227,N_1646,N_1748);
nor U3228 (N_3228,N_1109,N_662);
nor U3229 (N_3229,N_77,N_319);
nor U3230 (N_3230,N_770,N_1501);
xnor U3231 (N_3231,N_967,N_1785);
or U3232 (N_3232,N_1589,N_1464);
and U3233 (N_3233,N_192,N_1551);
and U3234 (N_3234,N_401,N_1096);
xor U3235 (N_3235,N_904,N_404);
or U3236 (N_3236,N_690,N_1398);
nor U3237 (N_3237,N_42,N_1192);
nand U3238 (N_3238,N_988,N_1613);
and U3239 (N_3239,N_287,N_439);
xor U3240 (N_3240,N_174,N_324);
nand U3241 (N_3241,N_1064,N_305);
nand U3242 (N_3242,N_1400,N_1168);
or U3243 (N_3243,N_11,N_267);
nand U3244 (N_3244,N_1745,N_1013);
or U3245 (N_3245,N_1831,N_277);
xnor U3246 (N_3246,N_1457,N_1199);
xnor U3247 (N_3247,N_707,N_1636);
xnor U3248 (N_3248,N_1644,N_593);
or U3249 (N_3249,N_1026,N_629);
nand U3250 (N_3250,N_1789,N_421);
nand U3251 (N_3251,N_1204,N_1351);
or U3252 (N_3252,N_877,N_1557);
and U3253 (N_3253,N_1818,N_719);
nor U3254 (N_3254,N_1329,N_724);
nor U3255 (N_3255,N_994,N_367);
nor U3256 (N_3256,N_1685,N_543);
xnor U3257 (N_3257,N_577,N_264);
and U3258 (N_3258,N_1412,N_128);
xnor U3259 (N_3259,N_145,N_167);
nand U3260 (N_3260,N_1511,N_153);
nor U3261 (N_3261,N_1446,N_700);
and U3262 (N_3262,N_1446,N_1972);
and U3263 (N_3263,N_1071,N_824);
xor U3264 (N_3264,N_8,N_1560);
nand U3265 (N_3265,N_1722,N_1742);
nor U3266 (N_3266,N_399,N_57);
xor U3267 (N_3267,N_954,N_1191);
nand U3268 (N_3268,N_546,N_1786);
and U3269 (N_3269,N_1902,N_1626);
or U3270 (N_3270,N_1956,N_333);
nand U3271 (N_3271,N_1568,N_1293);
and U3272 (N_3272,N_508,N_1901);
xor U3273 (N_3273,N_1352,N_824);
and U3274 (N_3274,N_317,N_1494);
xnor U3275 (N_3275,N_528,N_1093);
or U3276 (N_3276,N_1269,N_15);
and U3277 (N_3277,N_604,N_1281);
nand U3278 (N_3278,N_1813,N_189);
and U3279 (N_3279,N_80,N_1235);
and U3280 (N_3280,N_1929,N_842);
nand U3281 (N_3281,N_1522,N_979);
nand U3282 (N_3282,N_1957,N_1633);
or U3283 (N_3283,N_716,N_1023);
nor U3284 (N_3284,N_247,N_1939);
nand U3285 (N_3285,N_1179,N_1066);
nand U3286 (N_3286,N_867,N_957);
xnor U3287 (N_3287,N_1032,N_1451);
nor U3288 (N_3288,N_1328,N_1892);
xnor U3289 (N_3289,N_219,N_1352);
nor U3290 (N_3290,N_181,N_658);
or U3291 (N_3291,N_910,N_68);
nand U3292 (N_3292,N_1040,N_1146);
or U3293 (N_3293,N_802,N_1914);
nand U3294 (N_3294,N_1766,N_681);
and U3295 (N_3295,N_1830,N_930);
and U3296 (N_3296,N_405,N_60);
nand U3297 (N_3297,N_961,N_175);
or U3298 (N_3298,N_644,N_1658);
nor U3299 (N_3299,N_1696,N_1927);
and U3300 (N_3300,N_980,N_229);
xor U3301 (N_3301,N_463,N_650);
nor U3302 (N_3302,N_11,N_1529);
nor U3303 (N_3303,N_911,N_275);
xnor U3304 (N_3304,N_468,N_1305);
and U3305 (N_3305,N_1961,N_413);
and U3306 (N_3306,N_1612,N_968);
or U3307 (N_3307,N_1133,N_1601);
nand U3308 (N_3308,N_218,N_1291);
or U3309 (N_3309,N_271,N_1339);
or U3310 (N_3310,N_152,N_1392);
nor U3311 (N_3311,N_1468,N_1961);
nor U3312 (N_3312,N_408,N_678);
or U3313 (N_3313,N_682,N_302);
nor U3314 (N_3314,N_811,N_1315);
and U3315 (N_3315,N_995,N_944);
nand U3316 (N_3316,N_1015,N_1519);
or U3317 (N_3317,N_1633,N_1823);
nand U3318 (N_3318,N_752,N_472);
or U3319 (N_3319,N_1169,N_1584);
xor U3320 (N_3320,N_524,N_226);
or U3321 (N_3321,N_36,N_117);
nand U3322 (N_3322,N_1786,N_1644);
nor U3323 (N_3323,N_1357,N_45);
nor U3324 (N_3324,N_407,N_1273);
or U3325 (N_3325,N_1389,N_1352);
nand U3326 (N_3326,N_1054,N_260);
nor U3327 (N_3327,N_1940,N_1563);
and U3328 (N_3328,N_186,N_1358);
xnor U3329 (N_3329,N_546,N_1997);
or U3330 (N_3330,N_1452,N_470);
or U3331 (N_3331,N_837,N_955);
or U3332 (N_3332,N_293,N_1367);
and U3333 (N_3333,N_1063,N_1231);
nand U3334 (N_3334,N_279,N_1029);
and U3335 (N_3335,N_368,N_1249);
or U3336 (N_3336,N_299,N_1986);
or U3337 (N_3337,N_62,N_1776);
or U3338 (N_3338,N_1744,N_570);
nand U3339 (N_3339,N_201,N_5);
xnor U3340 (N_3340,N_352,N_652);
and U3341 (N_3341,N_940,N_840);
nor U3342 (N_3342,N_805,N_1483);
and U3343 (N_3343,N_1894,N_1422);
nor U3344 (N_3344,N_1324,N_1311);
nand U3345 (N_3345,N_1567,N_1653);
nand U3346 (N_3346,N_1916,N_891);
nor U3347 (N_3347,N_1628,N_221);
and U3348 (N_3348,N_432,N_521);
nor U3349 (N_3349,N_668,N_483);
or U3350 (N_3350,N_409,N_1618);
nand U3351 (N_3351,N_1840,N_1545);
nor U3352 (N_3352,N_1642,N_166);
xor U3353 (N_3353,N_456,N_198);
nand U3354 (N_3354,N_1802,N_955);
or U3355 (N_3355,N_1860,N_1497);
nor U3356 (N_3356,N_1285,N_739);
nand U3357 (N_3357,N_53,N_1724);
nand U3358 (N_3358,N_1077,N_112);
and U3359 (N_3359,N_658,N_1186);
nor U3360 (N_3360,N_1710,N_1487);
or U3361 (N_3361,N_1132,N_900);
xnor U3362 (N_3362,N_518,N_517);
and U3363 (N_3363,N_1716,N_508);
or U3364 (N_3364,N_91,N_1628);
nor U3365 (N_3365,N_1024,N_1218);
and U3366 (N_3366,N_601,N_942);
nand U3367 (N_3367,N_86,N_819);
and U3368 (N_3368,N_240,N_716);
xor U3369 (N_3369,N_1764,N_563);
or U3370 (N_3370,N_1388,N_1553);
nand U3371 (N_3371,N_730,N_1913);
xor U3372 (N_3372,N_1132,N_1478);
and U3373 (N_3373,N_400,N_894);
nand U3374 (N_3374,N_114,N_1350);
and U3375 (N_3375,N_1206,N_251);
xor U3376 (N_3376,N_610,N_1278);
nand U3377 (N_3377,N_1863,N_1249);
or U3378 (N_3378,N_757,N_1514);
xor U3379 (N_3379,N_365,N_154);
or U3380 (N_3380,N_1636,N_559);
xor U3381 (N_3381,N_155,N_1657);
nor U3382 (N_3382,N_174,N_428);
nand U3383 (N_3383,N_1352,N_840);
xor U3384 (N_3384,N_55,N_1494);
xnor U3385 (N_3385,N_1467,N_1718);
xnor U3386 (N_3386,N_326,N_1316);
or U3387 (N_3387,N_1427,N_307);
nor U3388 (N_3388,N_674,N_562);
nand U3389 (N_3389,N_107,N_932);
nand U3390 (N_3390,N_371,N_1284);
nand U3391 (N_3391,N_1709,N_447);
or U3392 (N_3392,N_1584,N_346);
nor U3393 (N_3393,N_108,N_349);
xnor U3394 (N_3394,N_1650,N_1966);
nor U3395 (N_3395,N_703,N_234);
nand U3396 (N_3396,N_1483,N_1929);
xor U3397 (N_3397,N_1030,N_712);
xnor U3398 (N_3398,N_409,N_647);
xnor U3399 (N_3399,N_564,N_1387);
nand U3400 (N_3400,N_1040,N_1625);
nor U3401 (N_3401,N_1652,N_211);
nor U3402 (N_3402,N_435,N_1282);
nand U3403 (N_3403,N_1284,N_1756);
xnor U3404 (N_3404,N_1509,N_1233);
nor U3405 (N_3405,N_59,N_209);
and U3406 (N_3406,N_1794,N_1237);
nand U3407 (N_3407,N_391,N_504);
or U3408 (N_3408,N_401,N_1883);
xnor U3409 (N_3409,N_195,N_648);
xnor U3410 (N_3410,N_990,N_93);
or U3411 (N_3411,N_1356,N_1351);
and U3412 (N_3412,N_228,N_1017);
nand U3413 (N_3413,N_1141,N_220);
xor U3414 (N_3414,N_317,N_1940);
or U3415 (N_3415,N_208,N_1514);
nor U3416 (N_3416,N_1504,N_1579);
and U3417 (N_3417,N_671,N_1374);
and U3418 (N_3418,N_181,N_382);
and U3419 (N_3419,N_635,N_370);
xnor U3420 (N_3420,N_406,N_1474);
nor U3421 (N_3421,N_93,N_307);
nor U3422 (N_3422,N_1087,N_1804);
xor U3423 (N_3423,N_1278,N_1034);
xnor U3424 (N_3424,N_806,N_1850);
xor U3425 (N_3425,N_1313,N_1819);
nand U3426 (N_3426,N_47,N_1610);
or U3427 (N_3427,N_149,N_1841);
xnor U3428 (N_3428,N_421,N_438);
or U3429 (N_3429,N_633,N_1137);
or U3430 (N_3430,N_1364,N_443);
nand U3431 (N_3431,N_976,N_24);
or U3432 (N_3432,N_1903,N_469);
nor U3433 (N_3433,N_1109,N_1895);
xnor U3434 (N_3434,N_708,N_78);
and U3435 (N_3435,N_31,N_534);
nand U3436 (N_3436,N_1601,N_1985);
and U3437 (N_3437,N_1768,N_314);
nor U3438 (N_3438,N_118,N_1450);
xnor U3439 (N_3439,N_519,N_366);
nand U3440 (N_3440,N_989,N_19);
and U3441 (N_3441,N_1228,N_1679);
nand U3442 (N_3442,N_1394,N_1450);
xnor U3443 (N_3443,N_1485,N_1098);
or U3444 (N_3444,N_315,N_597);
nand U3445 (N_3445,N_418,N_30);
nand U3446 (N_3446,N_353,N_714);
xnor U3447 (N_3447,N_761,N_99);
or U3448 (N_3448,N_312,N_772);
xor U3449 (N_3449,N_520,N_1965);
or U3450 (N_3450,N_1212,N_345);
xnor U3451 (N_3451,N_750,N_1134);
xnor U3452 (N_3452,N_828,N_199);
nor U3453 (N_3453,N_196,N_895);
nor U3454 (N_3454,N_1128,N_1005);
nand U3455 (N_3455,N_1780,N_1976);
or U3456 (N_3456,N_1899,N_899);
nor U3457 (N_3457,N_261,N_1414);
nor U3458 (N_3458,N_595,N_64);
xor U3459 (N_3459,N_1752,N_917);
nand U3460 (N_3460,N_490,N_1730);
xor U3461 (N_3461,N_389,N_144);
and U3462 (N_3462,N_125,N_1311);
nand U3463 (N_3463,N_319,N_1199);
nand U3464 (N_3464,N_1802,N_1436);
xnor U3465 (N_3465,N_1965,N_1004);
and U3466 (N_3466,N_1660,N_85);
xor U3467 (N_3467,N_1482,N_1153);
xnor U3468 (N_3468,N_1003,N_838);
xor U3469 (N_3469,N_1298,N_1894);
and U3470 (N_3470,N_1524,N_1669);
xor U3471 (N_3471,N_1922,N_1428);
xnor U3472 (N_3472,N_962,N_1509);
and U3473 (N_3473,N_1760,N_872);
nand U3474 (N_3474,N_1459,N_1549);
nor U3475 (N_3475,N_1196,N_1111);
or U3476 (N_3476,N_771,N_1149);
and U3477 (N_3477,N_1524,N_985);
nor U3478 (N_3478,N_947,N_1774);
nand U3479 (N_3479,N_547,N_1527);
and U3480 (N_3480,N_862,N_1767);
or U3481 (N_3481,N_1708,N_1333);
or U3482 (N_3482,N_82,N_1114);
nand U3483 (N_3483,N_1267,N_820);
nand U3484 (N_3484,N_319,N_1346);
and U3485 (N_3485,N_495,N_585);
nand U3486 (N_3486,N_1411,N_1689);
and U3487 (N_3487,N_1343,N_890);
nand U3488 (N_3488,N_1049,N_1425);
nor U3489 (N_3489,N_1430,N_28);
nor U3490 (N_3490,N_1002,N_1495);
or U3491 (N_3491,N_990,N_355);
nor U3492 (N_3492,N_142,N_1834);
nand U3493 (N_3493,N_1839,N_746);
or U3494 (N_3494,N_82,N_1634);
nor U3495 (N_3495,N_268,N_237);
and U3496 (N_3496,N_1276,N_98);
nor U3497 (N_3497,N_1346,N_543);
xnor U3498 (N_3498,N_1409,N_174);
or U3499 (N_3499,N_554,N_250);
and U3500 (N_3500,N_241,N_851);
nor U3501 (N_3501,N_1673,N_1580);
and U3502 (N_3502,N_1047,N_377);
and U3503 (N_3503,N_1057,N_792);
nor U3504 (N_3504,N_1830,N_1532);
nor U3505 (N_3505,N_97,N_1433);
or U3506 (N_3506,N_1274,N_1819);
nand U3507 (N_3507,N_604,N_1456);
and U3508 (N_3508,N_1314,N_1033);
xnor U3509 (N_3509,N_1161,N_1245);
and U3510 (N_3510,N_541,N_554);
or U3511 (N_3511,N_1079,N_1155);
nand U3512 (N_3512,N_889,N_495);
nand U3513 (N_3513,N_1916,N_1114);
or U3514 (N_3514,N_522,N_1500);
nor U3515 (N_3515,N_269,N_736);
nand U3516 (N_3516,N_1648,N_1315);
or U3517 (N_3517,N_1754,N_26);
or U3518 (N_3518,N_1526,N_482);
nand U3519 (N_3519,N_71,N_1039);
xor U3520 (N_3520,N_949,N_1762);
and U3521 (N_3521,N_1816,N_1979);
nand U3522 (N_3522,N_951,N_674);
or U3523 (N_3523,N_504,N_831);
or U3524 (N_3524,N_333,N_59);
nand U3525 (N_3525,N_862,N_1094);
and U3526 (N_3526,N_384,N_854);
xor U3527 (N_3527,N_333,N_495);
and U3528 (N_3528,N_958,N_1240);
nand U3529 (N_3529,N_933,N_1255);
nand U3530 (N_3530,N_1194,N_867);
nand U3531 (N_3531,N_1969,N_1326);
xor U3532 (N_3532,N_1020,N_57);
nor U3533 (N_3533,N_1247,N_1120);
nand U3534 (N_3534,N_1317,N_1480);
nor U3535 (N_3535,N_505,N_1953);
and U3536 (N_3536,N_363,N_998);
nand U3537 (N_3537,N_1746,N_1090);
and U3538 (N_3538,N_1078,N_1605);
nand U3539 (N_3539,N_1080,N_1717);
nand U3540 (N_3540,N_396,N_1386);
nor U3541 (N_3541,N_1350,N_629);
nand U3542 (N_3542,N_1391,N_62);
nand U3543 (N_3543,N_1131,N_1085);
or U3544 (N_3544,N_469,N_1992);
and U3545 (N_3545,N_1079,N_300);
nand U3546 (N_3546,N_1897,N_1663);
nand U3547 (N_3547,N_1824,N_942);
or U3548 (N_3548,N_45,N_811);
and U3549 (N_3549,N_1541,N_575);
nand U3550 (N_3550,N_498,N_1580);
and U3551 (N_3551,N_909,N_1796);
xnor U3552 (N_3552,N_1577,N_1109);
and U3553 (N_3553,N_1001,N_1657);
xnor U3554 (N_3554,N_1345,N_907);
xnor U3555 (N_3555,N_488,N_793);
nor U3556 (N_3556,N_1238,N_370);
nand U3557 (N_3557,N_1358,N_703);
or U3558 (N_3558,N_368,N_119);
xnor U3559 (N_3559,N_816,N_462);
or U3560 (N_3560,N_864,N_651);
nor U3561 (N_3561,N_985,N_336);
nor U3562 (N_3562,N_1589,N_1398);
and U3563 (N_3563,N_1307,N_1932);
nor U3564 (N_3564,N_1133,N_1060);
nand U3565 (N_3565,N_1408,N_1446);
nand U3566 (N_3566,N_1392,N_1226);
xor U3567 (N_3567,N_700,N_722);
nor U3568 (N_3568,N_620,N_1025);
and U3569 (N_3569,N_1290,N_1447);
xnor U3570 (N_3570,N_168,N_645);
nor U3571 (N_3571,N_603,N_1054);
and U3572 (N_3572,N_325,N_953);
xnor U3573 (N_3573,N_679,N_1217);
xor U3574 (N_3574,N_1729,N_711);
or U3575 (N_3575,N_1348,N_1479);
and U3576 (N_3576,N_212,N_1038);
nor U3577 (N_3577,N_198,N_546);
nor U3578 (N_3578,N_83,N_89);
nand U3579 (N_3579,N_280,N_124);
nor U3580 (N_3580,N_1559,N_12);
nand U3581 (N_3581,N_1713,N_349);
nand U3582 (N_3582,N_1518,N_1930);
nor U3583 (N_3583,N_1284,N_1833);
or U3584 (N_3584,N_314,N_1025);
or U3585 (N_3585,N_1069,N_104);
nand U3586 (N_3586,N_1484,N_39);
xor U3587 (N_3587,N_64,N_198);
and U3588 (N_3588,N_814,N_1195);
and U3589 (N_3589,N_1312,N_1207);
or U3590 (N_3590,N_1145,N_1959);
nor U3591 (N_3591,N_1450,N_1048);
nor U3592 (N_3592,N_995,N_882);
nand U3593 (N_3593,N_511,N_1308);
nor U3594 (N_3594,N_208,N_450);
nand U3595 (N_3595,N_1379,N_424);
or U3596 (N_3596,N_1842,N_816);
and U3597 (N_3597,N_1971,N_918);
xor U3598 (N_3598,N_1800,N_1754);
and U3599 (N_3599,N_902,N_1805);
nand U3600 (N_3600,N_309,N_882);
nor U3601 (N_3601,N_1317,N_1505);
and U3602 (N_3602,N_263,N_1724);
nor U3603 (N_3603,N_345,N_1429);
xnor U3604 (N_3604,N_67,N_80);
nand U3605 (N_3605,N_110,N_1253);
xnor U3606 (N_3606,N_1567,N_659);
and U3607 (N_3607,N_96,N_473);
and U3608 (N_3608,N_179,N_982);
xnor U3609 (N_3609,N_1561,N_604);
nor U3610 (N_3610,N_81,N_689);
nand U3611 (N_3611,N_509,N_937);
and U3612 (N_3612,N_1917,N_1921);
nor U3613 (N_3613,N_581,N_540);
and U3614 (N_3614,N_146,N_1951);
xnor U3615 (N_3615,N_159,N_1986);
nor U3616 (N_3616,N_106,N_39);
nor U3617 (N_3617,N_744,N_1718);
nand U3618 (N_3618,N_1474,N_1940);
nor U3619 (N_3619,N_1860,N_1564);
nor U3620 (N_3620,N_317,N_1762);
or U3621 (N_3621,N_905,N_732);
xnor U3622 (N_3622,N_1287,N_1990);
and U3623 (N_3623,N_1552,N_1806);
nand U3624 (N_3624,N_247,N_725);
nor U3625 (N_3625,N_57,N_1332);
xnor U3626 (N_3626,N_1991,N_1275);
xor U3627 (N_3627,N_1335,N_300);
nand U3628 (N_3628,N_1239,N_1576);
xnor U3629 (N_3629,N_1638,N_181);
nor U3630 (N_3630,N_157,N_1104);
and U3631 (N_3631,N_1915,N_1826);
xnor U3632 (N_3632,N_558,N_1813);
and U3633 (N_3633,N_1123,N_154);
and U3634 (N_3634,N_1414,N_1225);
nor U3635 (N_3635,N_998,N_616);
or U3636 (N_3636,N_672,N_1568);
and U3637 (N_3637,N_1760,N_1474);
xnor U3638 (N_3638,N_11,N_1717);
xor U3639 (N_3639,N_1662,N_1495);
and U3640 (N_3640,N_966,N_244);
nor U3641 (N_3641,N_145,N_55);
xnor U3642 (N_3642,N_1723,N_252);
nand U3643 (N_3643,N_1769,N_317);
or U3644 (N_3644,N_612,N_499);
xor U3645 (N_3645,N_1046,N_1213);
xnor U3646 (N_3646,N_1249,N_1704);
or U3647 (N_3647,N_1102,N_1806);
xnor U3648 (N_3648,N_1372,N_782);
nor U3649 (N_3649,N_1202,N_1003);
xor U3650 (N_3650,N_1866,N_559);
or U3651 (N_3651,N_840,N_648);
xnor U3652 (N_3652,N_422,N_1676);
and U3653 (N_3653,N_954,N_410);
nand U3654 (N_3654,N_1241,N_1561);
or U3655 (N_3655,N_229,N_1957);
or U3656 (N_3656,N_1412,N_1189);
or U3657 (N_3657,N_1018,N_125);
nand U3658 (N_3658,N_216,N_49);
and U3659 (N_3659,N_54,N_1777);
and U3660 (N_3660,N_118,N_870);
xnor U3661 (N_3661,N_630,N_1059);
nand U3662 (N_3662,N_1051,N_1266);
nor U3663 (N_3663,N_1899,N_1735);
nand U3664 (N_3664,N_131,N_1472);
nand U3665 (N_3665,N_792,N_435);
nand U3666 (N_3666,N_1135,N_332);
and U3667 (N_3667,N_1019,N_1201);
and U3668 (N_3668,N_185,N_1459);
nor U3669 (N_3669,N_1576,N_1697);
or U3670 (N_3670,N_337,N_1929);
xor U3671 (N_3671,N_243,N_353);
and U3672 (N_3672,N_557,N_1803);
nor U3673 (N_3673,N_1521,N_1239);
and U3674 (N_3674,N_265,N_1923);
nor U3675 (N_3675,N_1712,N_208);
xnor U3676 (N_3676,N_1894,N_1203);
and U3677 (N_3677,N_1586,N_1682);
xor U3678 (N_3678,N_1527,N_1507);
nor U3679 (N_3679,N_171,N_643);
and U3680 (N_3680,N_12,N_959);
nand U3681 (N_3681,N_417,N_890);
and U3682 (N_3682,N_1486,N_1686);
and U3683 (N_3683,N_1741,N_1780);
and U3684 (N_3684,N_1732,N_1729);
xnor U3685 (N_3685,N_1554,N_704);
nor U3686 (N_3686,N_29,N_517);
and U3687 (N_3687,N_1260,N_1291);
nor U3688 (N_3688,N_793,N_1418);
xor U3689 (N_3689,N_37,N_1462);
nor U3690 (N_3690,N_1314,N_1663);
and U3691 (N_3691,N_1699,N_321);
nand U3692 (N_3692,N_185,N_1015);
or U3693 (N_3693,N_391,N_796);
or U3694 (N_3694,N_901,N_1810);
xor U3695 (N_3695,N_620,N_1749);
nor U3696 (N_3696,N_268,N_1092);
nor U3697 (N_3697,N_1893,N_1620);
xor U3698 (N_3698,N_1063,N_1085);
and U3699 (N_3699,N_679,N_860);
nor U3700 (N_3700,N_1770,N_977);
or U3701 (N_3701,N_1798,N_985);
and U3702 (N_3702,N_491,N_1962);
and U3703 (N_3703,N_1000,N_1108);
or U3704 (N_3704,N_1830,N_1556);
nor U3705 (N_3705,N_502,N_1077);
and U3706 (N_3706,N_1787,N_1923);
xor U3707 (N_3707,N_752,N_1778);
xnor U3708 (N_3708,N_1341,N_1721);
xor U3709 (N_3709,N_1727,N_1435);
nor U3710 (N_3710,N_1997,N_1278);
xor U3711 (N_3711,N_1396,N_281);
and U3712 (N_3712,N_181,N_511);
xnor U3713 (N_3713,N_1393,N_747);
nand U3714 (N_3714,N_512,N_1321);
nand U3715 (N_3715,N_282,N_1097);
and U3716 (N_3716,N_729,N_1606);
xnor U3717 (N_3717,N_796,N_944);
xnor U3718 (N_3718,N_1573,N_990);
nor U3719 (N_3719,N_1775,N_1093);
or U3720 (N_3720,N_957,N_990);
and U3721 (N_3721,N_270,N_1108);
and U3722 (N_3722,N_1687,N_1244);
nor U3723 (N_3723,N_66,N_578);
nor U3724 (N_3724,N_723,N_1872);
xnor U3725 (N_3725,N_1598,N_532);
nand U3726 (N_3726,N_202,N_541);
and U3727 (N_3727,N_1949,N_808);
xor U3728 (N_3728,N_816,N_164);
and U3729 (N_3729,N_1940,N_1732);
nand U3730 (N_3730,N_1937,N_1714);
and U3731 (N_3731,N_1962,N_1945);
nand U3732 (N_3732,N_540,N_1739);
nand U3733 (N_3733,N_462,N_954);
and U3734 (N_3734,N_1112,N_114);
nand U3735 (N_3735,N_1798,N_142);
nor U3736 (N_3736,N_1051,N_1425);
or U3737 (N_3737,N_1773,N_259);
xor U3738 (N_3738,N_1060,N_1039);
nor U3739 (N_3739,N_758,N_28);
or U3740 (N_3740,N_1621,N_1653);
nor U3741 (N_3741,N_1766,N_1449);
nor U3742 (N_3742,N_702,N_942);
nor U3743 (N_3743,N_456,N_1478);
nor U3744 (N_3744,N_723,N_485);
or U3745 (N_3745,N_1883,N_715);
nor U3746 (N_3746,N_883,N_1026);
nor U3747 (N_3747,N_1206,N_1690);
nand U3748 (N_3748,N_1148,N_1786);
and U3749 (N_3749,N_617,N_716);
nor U3750 (N_3750,N_1873,N_1823);
nand U3751 (N_3751,N_468,N_7);
or U3752 (N_3752,N_1915,N_363);
nor U3753 (N_3753,N_1682,N_163);
or U3754 (N_3754,N_1878,N_1500);
xnor U3755 (N_3755,N_172,N_1631);
nor U3756 (N_3756,N_383,N_2);
nand U3757 (N_3757,N_1253,N_957);
or U3758 (N_3758,N_1254,N_414);
or U3759 (N_3759,N_1614,N_789);
nor U3760 (N_3760,N_1555,N_194);
and U3761 (N_3761,N_1649,N_558);
or U3762 (N_3762,N_1049,N_1062);
xor U3763 (N_3763,N_204,N_1263);
nand U3764 (N_3764,N_1873,N_1800);
and U3765 (N_3765,N_255,N_1158);
nand U3766 (N_3766,N_1348,N_1763);
and U3767 (N_3767,N_1777,N_1815);
nand U3768 (N_3768,N_1807,N_1059);
xnor U3769 (N_3769,N_929,N_1795);
nor U3770 (N_3770,N_1422,N_985);
nor U3771 (N_3771,N_841,N_971);
or U3772 (N_3772,N_1806,N_726);
nor U3773 (N_3773,N_1475,N_1258);
or U3774 (N_3774,N_341,N_1901);
nor U3775 (N_3775,N_501,N_982);
xor U3776 (N_3776,N_1544,N_487);
xnor U3777 (N_3777,N_173,N_209);
nand U3778 (N_3778,N_916,N_1852);
xor U3779 (N_3779,N_1482,N_1285);
xor U3780 (N_3780,N_1372,N_1578);
xnor U3781 (N_3781,N_215,N_400);
and U3782 (N_3782,N_1027,N_618);
nor U3783 (N_3783,N_1236,N_816);
xnor U3784 (N_3784,N_1748,N_1229);
nand U3785 (N_3785,N_1055,N_426);
or U3786 (N_3786,N_1688,N_1269);
or U3787 (N_3787,N_1061,N_1280);
and U3788 (N_3788,N_1355,N_1120);
nand U3789 (N_3789,N_1316,N_238);
or U3790 (N_3790,N_266,N_983);
nor U3791 (N_3791,N_1311,N_1859);
and U3792 (N_3792,N_918,N_1468);
and U3793 (N_3793,N_926,N_1037);
xor U3794 (N_3794,N_322,N_785);
xor U3795 (N_3795,N_22,N_393);
xor U3796 (N_3796,N_839,N_577);
nand U3797 (N_3797,N_1961,N_1795);
nor U3798 (N_3798,N_1413,N_702);
and U3799 (N_3799,N_1503,N_551);
and U3800 (N_3800,N_1260,N_1986);
and U3801 (N_3801,N_337,N_439);
or U3802 (N_3802,N_1763,N_356);
xnor U3803 (N_3803,N_1252,N_1830);
xnor U3804 (N_3804,N_1798,N_1306);
nand U3805 (N_3805,N_1563,N_1894);
xor U3806 (N_3806,N_162,N_1190);
or U3807 (N_3807,N_1172,N_403);
nor U3808 (N_3808,N_340,N_337);
and U3809 (N_3809,N_308,N_1886);
or U3810 (N_3810,N_1494,N_21);
or U3811 (N_3811,N_1495,N_1821);
or U3812 (N_3812,N_934,N_1351);
and U3813 (N_3813,N_1531,N_582);
and U3814 (N_3814,N_1494,N_1802);
and U3815 (N_3815,N_996,N_761);
nor U3816 (N_3816,N_1797,N_1817);
xnor U3817 (N_3817,N_944,N_446);
xnor U3818 (N_3818,N_585,N_1209);
nor U3819 (N_3819,N_1080,N_1509);
nor U3820 (N_3820,N_443,N_298);
xnor U3821 (N_3821,N_1283,N_1667);
nor U3822 (N_3822,N_1355,N_1394);
nor U3823 (N_3823,N_26,N_1176);
nor U3824 (N_3824,N_1959,N_1928);
nand U3825 (N_3825,N_1658,N_799);
or U3826 (N_3826,N_478,N_785);
and U3827 (N_3827,N_1154,N_1438);
or U3828 (N_3828,N_1732,N_1381);
and U3829 (N_3829,N_348,N_621);
or U3830 (N_3830,N_232,N_1637);
nand U3831 (N_3831,N_647,N_343);
and U3832 (N_3832,N_439,N_1034);
nor U3833 (N_3833,N_1689,N_1132);
nor U3834 (N_3834,N_1826,N_1109);
xor U3835 (N_3835,N_1090,N_1383);
nand U3836 (N_3836,N_1808,N_312);
nand U3837 (N_3837,N_682,N_475);
nand U3838 (N_3838,N_1573,N_826);
and U3839 (N_3839,N_1347,N_1409);
or U3840 (N_3840,N_6,N_1541);
nand U3841 (N_3841,N_1147,N_1191);
and U3842 (N_3842,N_571,N_841);
nor U3843 (N_3843,N_525,N_1023);
xor U3844 (N_3844,N_1151,N_1150);
nor U3845 (N_3845,N_572,N_618);
nand U3846 (N_3846,N_1950,N_202);
or U3847 (N_3847,N_402,N_484);
or U3848 (N_3848,N_1152,N_1912);
nor U3849 (N_3849,N_1148,N_679);
or U3850 (N_3850,N_1240,N_1265);
or U3851 (N_3851,N_1454,N_504);
nor U3852 (N_3852,N_833,N_470);
xnor U3853 (N_3853,N_959,N_1372);
xnor U3854 (N_3854,N_59,N_1998);
and U3855 (N_3855,N_1842,N_1949);
xor U3856 (N_3856,N_106,N_669);
nor U3857 (N_3857,N_593,N_787);
nor U3858 (N_3858,N_17,N_50);
and U3859 (N_3859,N_365,N_412);
or U3860 (N_3860,N_23,N_268);
or U3861 (N_3861,N_667,N_1275);
nor U3862 (N_3862,N_102,N_1731);
or U3863 (N_3863,N_808,N_1891);
and U3864 (N_3864,N_220,N_1190);
nor U3865 (N_3865,N_1593,N_830);
xor U3866 (N_3866,N_836,N_1920);
nor U3867 (N_3867,N_1139,N_764);
or U3868 (N_3868,N_1874,N_114);
and U3869 (N_3869,N_1270,N_638);
or U3870 (N_3870,N_878,N_1982);
or U3871 (N_3871,N_1660,N_1527);
xor U3872 (N_3872,N_1314,N_296);
and U3873 (N_3873,N_24,N_1241);
and U3874 (N_3874,N_683,N_1811);
nand U3875 (N_3875,N_1498,N_1211);
and U3876 (N_3876,N_1304,N_1429);
and U3877 (N_3877,N_428,N_832);
and U3878 (N_3878,N_1054,N_946);
nor U3879 (N_3879,N_880,N_368);
nor U3880 (N_3880,N_70,N_1467);
nand U3881 (N_3881,N_1161,N_1521);
nor U3882 (N_3882,N_1894,N_662);
nor U3883 (N_3883,N_1776,N_461);
or U3884 (N_3884,N_1178,N_1610);
nand U3885 (N_3885,N_185,N_1232);
and U3886 (N_3886,N_1759,N_299);
or U3887 (N_3887,N_1473,N_369);
nor U3888 (N_3888,N_170,N_1849);
or U3889 (N_3889,N_1338,N_1889);
xor U3890 (N_3890,N_499,N_618);
and U3891 (N_3891,N_1460,N_217);
nand U3892 (N_3892,N_1270,N_1238);
nor U3893 (N_3893,N_212,N_4);
and U3894 (N_3894,N_812,N_1525);
nor U3895 (N_3895,N_43,N_560);
or U3896 (N_3896,N_989,N_448);
and U3897 (N_3897,N_596,N_697);
nor U3898 (N_3898,N_319,N_1325);
nor U3899 (N_3899,N_1283,N_1810);
nor U3900 (N_3900,N_1743,N_63);
xor U3901 (N_3901,N_1502,N_132);
nor U3902 (N_3902,N_94,N_112);
nand U3903 (N_3903,N_1539,N_879);
nand U3904 (N_3904,N_1427,N_1973);
or U3905 (N_3905,N_1135,N_104);
xor U3906 (N_3906,N_1960,N_603);
nor U3907 (N_3907,N_1845,N_365);
nor U3908 (N_3908,N_1213,N_1133);
nand U3909 (N_3909,N_1959,N_1707);
xnor U3910 (N_3910,N_1541,N_1831);
or U3911 (N_3911,N_290,N_1442);
or U3912 (N_3912,N_1321,N_264);
nor U3913 (N_3913,N_1612,N_457);
nand U3914 (N_3914,N_1805,N_569);
nor U3915 (N_3915,N_539,N_187);
nand U3916 (N_3916,N_1303,N_67);
xnor U3917 (N_3917,N_1805,N_1202);
and U3918 (N_3918,N_1896,N_1342);
or U3919 (N_3919,N_1778,N_1411);
nand U3920 (N_3920,N_1797,N_1309);
or U3921 (N_3921,N_1588,N_893);
or U3922 (N_3922,N_1020,N_416);
or U3923 (N_3923,N_1882,N_1717);
or U3924 (N_3924,N_1500,N_674);
and U3925 (N_3925,N_1579,N_1616);
nor U3926 (N_3926,N_1997,N_605);
nor U3927 (N_3927,N_743,N_1788);
xnor U3928 (N_3928,N_534,N_886);
nor U3929 (N_3929,N_321,N_297);
nor U3930 (N_3930,N_1482,N_1863);
and U3931 (N_3931,N_1529,N_1784);
nor U3932 (N_3932,N_139,N_126);
or U3933 (N_3933,N_1631,N_842);
and U3934 (N_3934,N_1190,N_561);
and U3935 (N_3935,N_1640,N_1929);
and U3936 (N_3936,N_106,N_1149);
nand U3937 (N_3937,N_102,N_219);
nand U3938 (N_3938,N_444,N_392);
nand U3939 (N_3939,N_561,N_1153);
nor U3940 (N_3940,N_1318,N_1097);
nor U3941 (N_3941,N_1630,N_453);
nand U3942 (N_3942,N_693,N_858);
nand U3943 (N_3943,N_1100,N_1221);
nor U3944 (N_3944,N_1019,N_1542);
and U3945 (N_3945,N_730,N_1383);
or U3946 (N_3946,N_506,N_192);
xnor U3947 (N_3947,N_848,N_1829);
and U3948 (N_3948,N_1533,N_44);
or U3949 (N_3949,N_1992,N_324);
nand U3950 (N_3950,N_919,N_733);
and U3951 (N_3951,N_1632,N_1409);
nand U3952 (N_3952,N_1780,N_1495);
or U3953 (N_3953,N_741,N_1253);
xor U3954 (N_3954,N_1397,N_432);
nor U3955 (N_3955,N_1451,N_46);
nor U3956 (N_3956,N_1075,N_30);
and U3957 (N_3957,N_771,N_33);
nand U3958 (N_3958,N_318,N_1517);
or U3959 (N_3959,N_268,N_678);
nand U3960 (N_3960,N_954,N_952);
nand U3961 (N_3961,N_1155,N_305);
nor U3962 (N_3962,N_542,N_52);
nor U3963 (N_3963,N_1497,N_1609);
or U3964 (N_3964,N_236,N_1882);
or U3965 (N_3965,N_1764,N_1812);
and U3966 (N_3966,N_1204,N_1329);
and U3967 (N_3967,N_277,N_1755);
and U3968 (N_3968,N_25,N_1424);
and U3969 (N_3969,N_586,N_1427);
xnor U3970 (N_3970,N_1103,N_424);
nand U3971 (N_3971,N_857,N_841);
or U3972 (N_3972,N_1527,N_108);
and U3973 (N_3973,N_65,N_1555);
nor U3974 (N_3974,N_1129,N_962);
xnor U3975 (N_3975,N_1715,N_1202);
nand U3976 (N_3976,N_897,N_1497);
or U3977 (N_3977,N_443,N_923);
nor U3978 (N_3978,N_277,N_73);
or U3979 (N_3979,N_1583,N_1145);
nand U3980 (N_3980,N_1901,N_1049);
and U3981 (N_3981,N_1060,N_118);
and U3982 (N_3982,N_48,N_1629);
nand U3983 (N_3983,N_1451,N_429);
nand U3984 (N_3984,N_1660,N_978);
xnor U3985 (N_3985,N_742,N_671);
or U3986 (N_3986,N_1051,N_1465);
or U3987 (N_3987,N_1856,N_1449);
nor U3988 (N_3988,N_1376,N_366);
nand U3989 (N_3989,N_1851,N_113);
and U3990 (N_3990,N_218,N_845);
and U3991 (N_3991,N_155,N_645);
nor U3992 (N_3992,N_1503,N_298);
nand U3993 (N_3993,N_811,N_1902);
and U3994 (N_3994,N_1375,N_1173);
or U3995 (N_3995,N_1856,N_700);
nand U3996 (N_3996,N_1841,N_285);
nor U3997 (N_3997,N_869,N_1672);
nand U3998 (N_3998,N_923,N_1857);
or U3999 (N_3999,N_1960,N_426);
xnor U4000 (N_4000,N_2566,N_3838);
and U4001 (N_4001,N_3863,N_2316);
nor U4002 (N_4002,N_2754,N_2141);
or U4003 (N_4003,N_3037,N_2496);
xnor U4004 (N_4004,N_2099,N_3137);
nand U4005 (N_4005,N_3948,N_3759);
xor U4006 (N_4006,N_3974,N_3343);
and U4007 (N_4007,N_2290,N_2713);
or U4008 (N_4008,N_3513,N_2537);
xnor U4009 (N_4009,N_2365,N_2088);
xor U4010 (N_4010,N_2192,N_2643);
xor U4011 (N_4011,N_2687,N_2350);
xnor U4012 (N_4012,N_3786,N_3896);
nand U4013 (N_4013,N_2025,N_2143);
xor U4014 (N_4014,N_2959,N_2356);
nor U4015 (N_4015,N_2684,N_2852);
nand U4016 (N_4016,N_2925,N_2701);
xor U4017 (N_4017,N_2726,N_3163);
xor U4018 (N_4018,N_2013,N_3847);
and U4019 (N_4019,N_2724,N_2457);
nor U4020 (N_4020,N_2512,N_3151);
and U4021 (N_4021,N_2111,N_3980);
xnor U4022 (N_4022,N_2884,N_2881);
or U4023 (N_4023,N_3624,N_3443);
or U4024 (N_4024,N_2979,N_3779);
or U4025 (N_4025,N_2636,N_3601);
and U4026 (N_4026,N_2733,N_2879);
xnor U4027 (N_4027,N_3632,N_2763);
nand U4028 (N_4028,N_2862,N_3212);
nor U4029 (N_4029,N_3219,N_2407);
nand U4030 (N_4030,N_2026,N_3803);
nand U4031 (N_4031,N_2760,N_2390);
nor U4032 (N_4032,N_3520,N_2259);
nand U4033 (N_4033,N_2739,N_2461);
nor U4034 (N_4034,N_3679,N_2723);
xnor U4035 (N_4035,N_3501,N_3815);
and U4036 (N_4036,N_2393,N_2396);
or U4037 (N_4037,N_3606,N_2584);
nor U4038 (N_4038,N_2757,N_3511);
nand U4039 (N_4039,N_2888,N_3422);
xnor U4040 (N_4040,N_3428,N_2110);
and U4041 (N_4041,N_3008,N_2593);
nor U4042 (N_4042,N_2891,N_2284);
or U4043 (N_4043,N_3063,N_3699);
xnor U4044 (N_4044,N_3462,N_3584);
nand U4045 (N_4045,N_3197,N_3377);
and U4046 (N_4046,N_2460,N_2800);
xor U4047 (N_4047,N_3603,N_2834);
nor U4048 (N_4048,N_2789,N_2963);
nor U4049 (N_4049,N_2160,N_2294);
or U4050 (N_4050,N_3147,N_2231);
nand U4051 (N_4051,N_2326,N_3844);
or U4052 (N_4052,N_3716,N_3011);
nor U4053 (N_4053,N_2694,N_3857);
and U4054 (N_4054,N_3537,N_2454);
nand U4055 (N_4055,N_3684,N_3814);
or U4056 (N_4056,N_3991,N_2405);
nand U4057 (N_4057,N_3269,N_2742);
xor U4058 (N_4058,N_3527,N_2240);
nor U4059 (N_4059,N_3136,N_2258);
nand U4060 (N_4060,N_3719,N_2187);
or U4061 (N_4061,N_3528,N_3496);
nor U4062 (N_4062,N_3555,N_2164);
nor U4063 (N_4063,N_2422,N_2533);
or U4064 (N_4064,N_3899,N_3125);
or U4065 (N_4065,N_2277,N_3795);
xnor U4066 (N_4066,N_3502,N_2436);
nor U4067 (N_4067,N_2897,N_3696);
or U4068 (N_4068,N_3039,N_3972);
xnor U4069 (N_4069,N_3425,N_3308);
xnor U4070 (N_4070,N_2960,N_3346);
nand U4071 (N_4071,N_2886,N_3467);
xnor U4072 (N_4072,N_3956,N_2796);
or U4073 (N_4073,N_2131,N_3214);
nand U4074 (N_4074,N_2112,N_2541);
or U4075 (N_4075,N_3851,N_2139);
nor U4076 (N_4076,N_3303,N_2354);
nand U4077 (N_4077,N_3328,N_2828);
or U4078 (N_4078,N_3869,N_3506);
xnor U4079 (N_4079,N_3352,N_3598);
nand U4080 (N_4080,N_3327,N_2664);
xor U4081 (N_4081,N_3194,N_3764);
nand U4082 (N_4082,N_2753,N_2621);
nand U4083 (N_4083,N_2264,N_3454);
xnor U4084 (N_4084,N_2462,N_2179);
nand U4085 (N_4085,N_2295,N_3121);
or U4086 (N_4086,N_2971,N_2603);
and U4087 (N_4087,N_3044,N_3808);
nor U4088 (N_4088,N_2338,N_2311);
and U4089 (N_4089,N_2340,N_3668);
and U4090 (N_4090,N_3401,N_3191);
nor U4091 (N_4091,N_2469,N_3973);
or U4092 (N_4092,N_2820,N_2571);
and U4093 (N_4093,N_2178,N_2146);
and U4094 (N_4094,N_3834,N_2681);
xor U4095 (N_4095,N_2586,N_3762);
nand U4096 (N_4096,N_3867,N_3643);
nand U4097 (N_4097,N_3231,N_2648);
nor U4098 (N_4098,N_3497,N_2317);
and U4099 (N_4099,N_3638,N_2916);
or U4100 (N_4100,N_3267,N_2361);
or U4101 (N_4101,N_2434,N_2638);
nand U4102 (N_4102,N_3409,N_3066);
or U4103 (N_4103,N_3205,N_2659);
nand U4104 (N_4104,N_2425,N_3203);
nor U4105 (N_4105,N_3914,N_2423);
xor U4106 (N_4106,N_2734,N_2500);
nand U4107 (N_4107,N_2810,N_2251);
and U4108 (N_4108,N_2988,N_3288);
xnor U4109 (N_4109,N_3547,N_3718);
nand U4110 (N_4110,N_3540,N_2610);
nor U4111 (N_4111,N_3741,N_3217);
nor U4112 (N_4112,N_3423,N_3397);
and U4113 (N_4113,N_2710,N_3441);
nor U4114 (N_4114,N_2438,N_3969);
or U4115 (N_4115,N_3550,N_2181);
or U4116 (N_4116,N_2003,N_3342);
nand U4117 (N_4117,N_2174,N_3539);
nor U4118 (N_4118,N_2081,N_2993);
and U4119 (N_4119,N_3061,N_3260);
xor U4120 (N_4120,N_2282,N_2902);
xnor U4121 (N_4121,N_2556,N_2836);
xor U4122 (N_4122,N_2587,N_2996);
and U4123 (N_4123,N_2458,N_3596);
xnor U4124 (N_4124,N_3849,N_2074);
and U4125 (N_4125,N_3617,N_3033);
and U4126 (N_4126,N_2216,N_3070);
nor U4127 (N_4127,N_2649,N_2832);
or U4128 (N_4128,N_2589,N_2903);
xor U4129 (N_4129,N_3531,N_2008);
nand U4130 (N_4130,N_2673,N_3530);
xor U4131 (N_4131,N_3772,N_2823);
and U4132 (N_4132,N_2762,N_3856);
xnor U4133 (N_4133,N_3650,N_2369);
xor U4134 (N_4134,N_3180,N_3870);
nand U4135 (N_4135,N_2297,N_3154);
or U4136 (N_4136,N_3592,N_3349);
nand U4137 (N_4137,N_2005,N_2287);
nand U4138 (N_4138,N_2104,N_2947);
nor U4139 (N_4139,N_3712,N_2036);
xor U4140 (N_4140,N_3209,N_3153);
xor U4141 (N_4141,N_2332,N_2688);
xnor U4142 (N_4142,N_3266,N_3736);
and U4143 (N_4143,N_3620,N_3521);
xor U4144 (N_4144,N_3618,N_3590);
or U4145 (N_4145,N_3612,N_3608);
nor U4146 (N_4146,N_2633,N_3049);
and U4147 (N_4147,N_3631,N_3281);
xnor U4148 (N_4148,N_3913,N_3418);
and U4149 (N_4149,N_3305,N_2871);
nor U4150 (N_4150,N_3235,N_2414);
xor U4151 (N_4151,N_3414,N_3324);
and U4152 (N_4152,N_2235,N_3571);
and U4153 (N_4153,N_3236,N_2601);
and U4154 (N_4154,N_2484,N_2676);
nand U4155 (N_4155,N_2339,N_2301);
and U4156 (N_4156,N_3561,N_3080);
or U4157 (N_4157,N_3742,N_3187);
xor U4158 (N_4158,N_2464,N_3623);
nor U4159 (N_4159,N_3196,N_3130);
or U4160 (N_4160,N_3720,N_2585);
xnor U4161 (N_4161,N_3495,N_2012);
xor U4162 (N_4162,N_2825,N_3797);
or U4163 (N_4163,N_2218,N_2315);
nor U4164 (N_4164,N_3802,N_3126);
or U4165 (N_4165,N_2391,N_2530);
nand U4166 (N_4166,N_3490,N_2854);
and U4167 (N_4167,N_2037,N_2715);
and U4168 (N_4168,N_3320,N_3569);
xor U4169 (N_4169,N_3998,N_2529);
nor U4170 (N_4170,N_3532,N_2728);
and U4171 (N_4171,N_3007,N_2552);
xor U4172 (N_4172,N_2653,N_3192);
nand U4173 (N_4173,N_2278,N_3947);
nor U4174 (N_4174,N_2043,N_2949);
and U4175 (N_4175,N_3483,N_2722);
nor U4176 (N_4176,N_3118,N_3405);
or U4177 (N_4177,N_3613,N_2213);
xnor U4178 (N_4178,N_2750,N_2867);
nand U4179 (N_4179,N_2892,N_2280);
xnor U4180 (N_4180,N_3564,N_3104);
xor U4181 (N_4181,N_2120,N_3651);
nor U4182 (N_4182,N_3081,N_3408);
and U4183 (N_4183,N_2882,N_2686);
or U4184 (N_4184,N_3204,N_2794);
nor U4185 (N_4185,N_2766,N_2122);
and U4186 (N_4186,N_3745,N_3293);
or U4187 (N_4187,N_2581,N_3404);
xnor U4188 (N_4188,N_2743,N_2241);
and U4189 (N_4189,N_3107,N_2144);
nand U4190 (N_4190,N_2072,N_3050);
and U4191 (N_4191,N_2207,N_2569);
or U4192 (N_4192,N_3032,N_3333);
nor U4193 (N_4193,N_3680,N_2906);
nor U4194 (N_4194,N_3744,N_2576);
xnor U4195 (N_4195,N_3472,N_3394);
xor U4196 (N_4196,N_3378,N_2738);
and U4197 (N_4197,N_3416,N_2166);
and U4198 (N_4198,N_2558,N_3583);
xnor U4199 (N_4199,N_2439,N_2616);
nor U4200 (N_4200,N_2864,N_3774);
and U4201 (N_4201,N_3591,N_3085);
xnor U4202 (N_4202,N_3934,N_2783);
nor U4203 (N_4203,N_3445,N_2437);
or U4204 (N_4204,N_2957,N_2334);
or U4205 (N_4205,N_2094,N_2087);
nor U4206 (N_4206,N_2101,N_2986);
nand U4207 (N_4207,N_2381,N_3082);
and U4208 (N_4208,N_3227,N_3239);
nor U4209 (N_4209,N_2215,N_3156);
xor U4210 (N_4210,N_2124,N_3688);
nor U4211 (N_4211,N_2914,N_2736);
nor U4212 (N_4212,N_3941,N_3709);
or U4213 (N_4213,N_2815,N_3117);
and U4214 (N_4214,N_3315,N_3283);
xnor U4215 (N_4215,N_3514,N_2430);
nand U4216 (N_4216,N_3412,N_3999);
xnor U4217 (N_4217,N_3048,N_3337);
nand U4218 (N_4218,N_3548,N_3076);
and U4219 (N_4219,N_3348,N_3339);
or U4220 (N_4220,N_2698,N_3903);
or U4221 (N_4221,N_3477,N_3186);
nand U4222 (N_4222,N_2497,N_3955);
nor U4223 (N_4223,N_3637,N_2296);
xnor U4224 (N_4224,N_2032,N_3034);
nor U4225 (N_4225,N_2699,N_3731);
nand U4226 (N_4226,N_2225,N_2307);
or U4227 (N_4227,N_3993,N_2837);
xnor U4228 (N_4228,N_2261,N_3458);
nor U4229 (N_4229,N_3480,N_3439);
xor U4230 (N_4230,N_3202,N_2358);
or U4231 (N_4231,N_2378,N_3110);
xnor U4232 (N_4232,N_2983,N_2406);
or U4233 (N_4233,N_3355,N_3058);
nor U4234 (N_4234,N_2158,N_2588);
and U4235 (N_4235,N_2525,N_2106);
nand U4236 (N_4236,N_3662,N_2780);
xor U4237 (N_4237,N_3880,N_2901);
or U4238 (N_4238,N_3799,N_3825);
or U4239 (N_4239,N_2926,N_2217);
xnor U4240 (N_4240,N_3395,N_2656);
nand U4241 (N_4241,N_2703,N_3170);
or U4242 (N_4242,N_3924,N_2865);
nor U4243 (N_4243,N_2389,N_2476);
and U4244 (N_4244,N_2619,N_2546);
nand U4245 (N_4245,N_2674,N_3859);
nand U4246 (N_4246,N_3396,N_3357);
nor U4247 (N_4247,N_3806,N_2455);
nand U4248 (N_4248,N_2328,N_3525);
nor U4249 (N_4249,N_2716,N_3330);
xor U4250 (N_4250,N_3965,N_2029);
nand U4251 (N_4251,N_3178,N_3754);
nand U4252 (N_4252,N_2163,N_2083);
and U4253 (N_4253,N_2620,N_2490);
nor U4254 (N_4254,N_3000,N_3344);
or U4255 (N_4255,N_3215,N_3456);
nor U4256 (N_4256,N_2019,N_2349);
nor U4257 (N_4257,N_2096,N_2912);
nand U4258 (N_4258,N_3546,N_3981);
nor U4259 (N_4259,N_3166,N_3064);
xor U4260 (N_4260,N_3024,N_2799);
nor U4261 (N_4261,N_3894,N_2404);
xnor U4262 (N_4262,N_2097,N_3630);
or U4263 (N_4263,N_3672,N_2675);
xor U4264 (N_4264,N_3358,N_2802);
nand U4265 (N_4265,N_2010,N_3629);
xnor U4266 (N_4266,N_2161,N_3966);
or U4267 (N_4267,N_2532,N_3001);
and U4268 (N_4268,N_3545,N_3882);
or U4269 (N_4269,N_2078,N_3817);
nand U4270 (N_4270,N_3491,N_3379);
and U4271 (N_4271,N_3012,N_2325);
and U4272 (N_4272,N_2090,N_2070);
or U4273 (N_4273,N_3400,N_3549);
xnor U4274 (N_4274,N_2135,N_3952);
or U4275 (N_4275,N_2858,N_2555);
and U4276 (N_4276,N_2397,N_2981);
nand U4277 (N_4277,N_3242,N_2978);
nor U4278 (N_4278,N_2493,N_3470);
nand U4279 (N_4279,N_3938,N_2298);
or U4280 (N_4280,N_3131,N_2343);
or U4281 (N_4281,N_3120,N_3524);
or U4282 (N_4282,N_3855,N_3829);
nor U4283 (N_4283,N_3983,N_2540);
or U4284 (N_4284,N_2923,N_3074);
xnor U4285 (N_4285,N_2456,N_2807);
xor U4286 (N_4286,N_3595,N_3171);
or U4287 (N_4287,N_3579,N_2966);
xnor U4288 (N_4288,N_2672,N_3289);
or U4289 (N_4289,N_3469,N_3415);
and U4290 (N_4290,N_3959,N_2333);
or U4291 (N_4291,N_3100,N_3901);
nor U4292 (N_4292,N_3134,N_2053);
xnor U4293 (N_4293,N_2034,N_3389);
or U4294 (N_4294,N_3371,N_2579);
and U4295 (N_4295,N_2682,N_3257);
and U4296 (N_4296,N_2953,N_3951);
and U4297 (N_4297,N_3536,N_2549);
and U4298 (N_4298,N_2467,N_2424);
or U4299 (N_4299,N_3557,N_3791);
xnor U4300 (N_4300,N_3282,N_2934);
nand U4301 (N_4301,N_2450,N_3427);
and U4302 (N_4302,N_2082,N_2792);
xor U4303 (N_4303,N_3724,N_2929);
nor U4304 (N_4304,N_2039,N_3332);
xnor U4305 (N_4305,N_2995,N_2685);
and U4306 (N_4306,N_3347,N_2441);
and U4307 (N_4307,N_2759,N_3658);
nor U4308 (N_4308,N_2909,N_2024);
and U4309 (N_4309,N_2773,N_2248);
and U4310 (N_4310,N_2958,N_3188);
nor U4311 (N_4311,N_3961,N_3158);
and U4312 (N_4312,N_2851,N_2204);
and U4313 (N_4313,N_2335,N_3167);
nor U4314 (N_4314,N_3950,N_2017);
nand U4315 (N_4315,N_2324,N_2501);
xor U4316 (N_4316,N_3733,N_3753);
xor U4317 (N_4317,N_2885,N_3173);
nand U4318 (N_4318,N_2410,N_2568);
nor U4319 (N_4319,N_3448,N_3848);
and U4320 (N_4320,N_2015,N_2877);
xor U4321 (N_4321,N_3297,N_2692);
nor U4322 (N_4322,N_2863,N_3986);
or U4323 (N_4323,N_2360,N_2895);
nor U4324 (N_4324,N_3944,N_2813);
or U4325 (N_4325,N_3836,N_2847);
nand U4326 (N_4326,N_3928,N_2528);
nand U4327 (N_4327,N_2839,N_3782);
nand U4328 (N_4328,N_2527,N_3975);
or U4329 (N_4329,N_2353,N_3190);
or U4330 (N_4330,N_2679,N_3014);
nor U4331 (N_4331,N_2394,N_3509);
nand U4332 (N_4332,N_2159,N_3380);
xnor U4333 (N_4333,N_3677,N_2092);
xnor U4334 (N_4334,N_2545,N_3093);
nand U4335 (N_4335,N_2075,N_2388);
or U4336 (N_4336,N_2383,N_3552);
nor U4337 (N_4337,N_2704,N_2275);
nor U4338 (N_4338,N_3693,N_3810);
nand U4339 (N_4339,N_2318,N_2293);
and U4340 (N_4340,N_3619,N_2761);
or U4341 (N_4341,N_3660,N_3097);
and U4342 (N_4342,N_2591,N_2067);
and U4343 (N_4343,N_2086,N_2835);
xor U4344 (N_4344,N_3554,N_3905);
nor U4345 (N_4345,N_3176,N_2431);
xnor U4346 (N_4346,N_2818,N_3706);
xor U4347 (N_4347,N_2697,N_3570);
and U4348 (N_4348,N_3893,N_2970);
xnor U4349 (N_4349,N_2196,N_2706);
and U4350 (N_4350,N_3261,N_2374);
xor U4351 (N_4351,N_2058,N_2635);
xor U4352 (N_4352,N_2271,N_2624);
and U4353 (N_4353,N_3115,N_2193);
nand U4354 (N_4354,N_3860,N_2173);
nand U4355 (N_4355,N_3465,N_3884);
nand U4356 (N_4356,N_2907,N_3172);
or U4357 (N_4357,N_2031,N_3770);
nand U4358 (N_4358,N_2420,N_3087);
nand U4359 (N_4359,N_3751,N_2273);
or U4360 (N_4360,N_3157,N_2984);
xnor U4361 (N_4361,N_3175,N_2562);
and U4362 (N_4362,N_3626,N_3224);
nor U4363 (N_4363,N_2409,N_3383);
or U4364 (N_4364,N_2502,N_2744);
nand U4365 (N_4365,N_2057,N_2479);
xor U4366 (N_4366,N_2860,N_2913);
xor U4367 (N_4367,N_2997,N_2602);
xor U4368 (N_4368,N_3988,N_2942);
or U4369 (N_4369,N_2866,N_3634);
or U4370 (N_4370,N_3287,N_3967);
nor U4371 (N_4371,N_2018,N_3438);
and U4372 (N_4372,N_3079,N_3199);
and U4373 (N_4373,N_3698,N_2812);
or U4374 (N_4374,N_3642,N_3312);
nand U4375 (N_4375,N_2195,N_2531);
and U4376 (N_4376,N_3877,N_2752);
xnor U4377 (N_4377,N_2985,N_3486);
nand U4378 (N_4378,N_3687,N_2180);
nand U4379 (N_4379,N_2683,N_2518);
or U4380 (N_4380,N_3083,N_3374);
or U4381 (N_4381,N_2473,N_3426);
and U4382 (N_4382,N_2345,N_3168);
or U4383 (N_4383,N_3850,N_2059);
xor U4384 (N_4384,N_3311,N_2254);
or U4385 (N_4385,N_3519,N_3459);
or U4386 (N_4386,N_3653,N_2227);
nor U4387 (N_4387,N_3290,N_2416);
or U4388 (N_4388,N_3558,N_2401);
and U4389 (N_4389,N_2140,N_2076);
nand U4390 (N_4390,N_3141,N_2557);
or U4391 (N_4391,N_2249,N_2150);
or U4392 (N_4392,N_2662,N_3604);
nand U4393 (N_4393,N_3406,N_2319);
and U4394 (N_4394,N_3887,N_3046);
xnor U4395 (N_4395,N_2162,N_2543);
nor U4396 (N_4396,N_2973,N_2370);
and U4397 (N_4397,N_2507,N_3099);
xnor U4398 (N_4398,N_3113,N_2646);
nand U4399 (N_4399,N_3645,N_2890);
and U4400 (N_4400,N_2534,N_3403);
xor U4401 (N_4401,N_2267,N_2288);
or U4402 (N_4402,N_2874,N_3649);
nand U4403 (N_4403,N_3270,N_2265);
nand U4404 (N_4404,N_2998,N_3112);
or U4405 (N_4405,N_2650,N_2725);
nand U4406 (N_4406,N_3902,N_3589);
xor U4407 (N_4407,N_3695,N_2172);
xor U4408 (N_4408,N_2027,N_3256);
nor U4409 (N_4409,N_3375,N_3129);
nor U4410 (N_4410,N_2481,N_3241);
nand U4411 (N_4411,N_2253,N_3135);
nor U4412 (N_4412,N_3429,N_3432);
nand U4413 (N_4413,N_3225,N_2242);
xnor U4414 (N_4414,N_2509,N_2355);
and U4415 (N_4415,N_2047,N_3229);
xor U4416 (N_4416,N_2746,N_3086);
or U4417 (N_4417,N_2004,N_2904);
nor U4418 (N_4418,N_3907,N_3946);
xor U4419 (N_4419,N_3906,N_2064);
and U4420 (N_4420,N_3710,N_2940);
xor U4421 (N_4421,N_2859,N_3310);
nand U4422 (N_4422,N_3165,N_2045);
and U4423 (N_4423,N_3193,N_3597);
or U4424 (N_4424,N_2084,N_3184);
or U4425 (N_4425,N_2841,N_2880);
nor U4426 (N_4426,N_2544,N_2002);
or U4427 (N_4427,N_3610,N_2151);
nor U4428 (N_4428,N_2089,N_3245);
nor U4429 (N_4429,N_3321,N_2411);
nand U4430 (N_4430,N_2263,N_3852);
nand U4431 (N_4431,N_2910,N_3286);
nand U4432 (N_4432,N_2898,N_3990);
nand U4433 (N_4433,N_2344,N_3895);
nand U4434 (N_4434,N_3707,N_2449);
and U4435 (N_4435,N_2062,N_2779);
nand U4436 (N_4436,N_2931,N_3370);
nand U4437 (N_4437,N_2690,N_2351);
or U4438 (N_4438,N_2782,N_3373);
nand U4439 (N_4439,N_2126,N_2768);
nor U4440 (N_4440,N_3237,N_2575);
or U4441 (N_4441,N_3164,N_3790);
or U4442 (N_4442,N_3211,N_2384);
or U4443 (N_4443,N_3730,N_3306);
xnor U4444 (N_4444,N_2051,N_2520);
xnor U4445 (N_4445,N_2765,N_3484);
nand U4446 (N_4446,N_3898,N_3159);
nand U4447 (N_4447,N_3654,N_3302);
xnor U4448 (N_4448,N_3865,N_2709);
nor U4449 (N_4449,N_2471,N_3124);
nor U4450 (N_4450,N_3466,N_2379);
nand U4451 (N_4451,N_3890,N_3916);
nand U4452 (N_4452,N_2021,N_3005);
nand U4453 (N_4453,N_2515,N_2695);
nor U4454 (N_4454,N_3757,N_2432);
and U4455 (N_4455,N_2244,N_3161);
nand U4456 (N_4456,N_2133,N_2559);
or U4457 (N_4457,N_2016,N_3451);
xor U4458 (N_4458,N_2505,N_2157);
and U4459 (N_4459,N_2330,N_3060);
and U4460 (N_4460,N_2368,N_2447);
xnor U4461 (N_4461,N_3278,N_2367);
nand U4462 (N_4462,N_2849,N_3700);
or U4463 (N_4463,N_3659,N_2130);
or U4464 (N_4464,N_2784,N_3249);
and U4465 (N_4465,N_3781,N_2939);
and U4466 (N_4466,N_2811,N_2128);
and U4467 (N_4467,N_3873,N_3016);
nand U4468 (N_4468,N_3433,N_3195);
or U4469 (N_4469,N_3542,N_3639);
xnor U4470 (N_4470,N_3078,N_2079);
and U4471 (N_4471,N_3027,N_3372);
xnor U4472 (N_4472,N_3384,N_2737);
xor U4473 (N_4473,N_3734,N_3253);
xor U4474 (N_4474,N_3367,N_2956);
nor U4475 (N_4475,N_3299,N_2442);
or U4476 (N_4476,N_2526,N_2102);
xor U4477 (N_4477,N_2614,N_2440);
xnor U4478 (N_4478,N_2071,N_2190);
nand U4479 (N_4479,N_3541,N_3010);
nor U4480 (N_4480,N_3073,N_3923);
and U4481 (N_4481,N_2310,N_3336);
nor U4482 (N_4482,N_3119,N_3210);
nand U4483 (N_4483,N_3737,N_3273);
nor U4484 (N_4484,N_2061,N_2831);
or U4485 (N_4485,N_2595,N_3600);
nand U4486 (N_4486,N_2395,N_3132);
nor U4487 (N_4487,N_3985,N_3566);
xor U4488 (N_4488,N_2109,N_3691);
nor U4489 (N_4489,N_3879,N_2419);
or U4490 (N_4490,N_2063,N_2982);
and U4491 (N_4491,N_2482,N_3382);
and U4492 (N_4492,N_2702,N_2804);
and U4493 (N_4493,N_3381,N_2080);
or U4494 (N_4494,N_3169,N_3259);
nor U4495 (N_4495,N_3017,N_2376);
and U4496 (N_4496,N_2663,N_2950);
and U4497 (N_4497,N_2590,N_3670);
nor U4498 (N_4498,N_3300,N_2776);
or U4499 (N_4499,N_2030,N_2582);
or U4500 (N_4500,N_3155,N_3341);
and U4501 (N_4501,N_3878,N_3162);
and U4502 (N_4502,N_2435,N_2764);
nor U4503 (N_4503,N_2669,N_2220);
nor U4504 (N_4504,N_2478,N_2572);
nand U4505 (N_4505,N_3666,N_2236);
nand U4506 (N_4506,N_3182,N_3363);
or U4507 (N_4507,N_3218,N_3387);
and U4508 (N_4508,N_3821,N_2127);
xnor U4509 (N_4509,N_2511,N_2727);
nand U4510 (N_4510,N_2312,N_2928);
and U4511 (N_4511,N_3538,N_3811);
or U4512 (N_4512,N_3077,N_3272);
or U4513 (N_4513,N_3833,N_2289);
nor U4514 (N_4514,N_2299,N_3831);
or U4515 (N_4515,N_3627,N_3468);
nor U4516 (N_4516,N_3805,N_3492);
xnor U4517 (N_4517,N_2320,N_2418);
nor U4518 (N_4518,N_2922,N_2185);
nor U4519 (N_4519,N_2038,N_2232);
or U4520 (N_4520,N_2941,N_2085);
nand U4521 (N_4521,N_3517,N_2547);
nand U4522 (N_4522,N_2219,N_3937);
and U4523 (N_4523,N_2487,N_3230);
and U4524 (N_4524,N_3777,N_2772);
or U4525 (N_4525,N_3264,N_2771);
or U4526 (N_4526,N_2612,N_2639);
or U4527 (N_4527,N_2974,N_3703);
or U4528 (N_4528,N_2303,N_2357);
nand U4529 (N_4529,N_3291,N_2352);
and U4530 (N_4530,N_3090,N_3739);
xor U4531 (N_4531,N_2609,N_3673);
nor U4532 (N_4532,N_3578,N_2747);
and U4533 (N_4533,N_3766,N_3819);
nor U4534 (N_4534,N_2323,N_3789);
or U4535 (N_4535,N_2040,N_3785);
or U4536 (N_4536,N_2170,N_3216);
and U4537 (N_4537,N_2732,N_2574);
xor U4538 (N_4538,N_3294,N_2247);
nand U4539 (N_4539,N_2044,N_3954);
xor U4540 (N_4540,N_2055,N_3128);
and U4541 (N_4541,N_2305,N_2188);
nor U4542 (N_4542,N_3885,N_3255);
xor U4543 (N_4543,N_3783,N_3052);
xnor U4544 (N_4544,N_2100,N_3399);
xnor U4545 (N_4545,N_2211,N_2917);
nor U4546 (N_4546,N_3471,N_2403);
nor U4547 (N_4547,N_3793,N_3243);
or U4548 (N_4548,N_3727,N_3711);
nor U4549 (N_4549,N_2668,N_2667);
nor U4550 (N_4550,N_3301,N_2987);
or U4551 (N_4551,N_2065,N_2808);
xor U4552 (N_4552,N_3127,N_2252);
nor U4553 (N_4553,N_2905,N_3562);
nor U4554 (N_4554,N_3065,N_2637);
xor U4555 (N_4555,N_3576,N_3362);
xor U4556 (N_4556,N_2302,N_2787);
and U4557 (N_4557,N_2492,N_2915);
nor U4558 (N_4558,N_2116,N_2142);
and U4559 (N_4559,N_3464,N_2514);
xor U4560 (N_4560,N_2426,N_3200);
and U4561 (N_4561,N_3420,N_3240);
and U4562 (N_4562,N_3174,N_2816);
nand U4563 (N_4563,N_3813,N_2696);
nor U4564 (N_4564,N_3254,N_3945);
xor U4565 (N_4565,N_3233,N_3251);
nor U4566 (N_4566,N_2226,N_3244);
nor U4567 (N_4567,N_2028,N_2183);
nand U4568 (N_4568,N_2286,N_2472);
xnor U4569 (N_4569,N_3338,N_3036);
xor U4570 (N_4570,N_2967,N_2499);
nor U4571 (N_4571,N_3667,N_2838);
or U4572 (N_4572,N_3922,N_2304);
and U4573 (N_4573,N_2077,N_3478);
nand U4574 (N_4574,N_3031,N_2645);
nor U4575 (N_4575,N_2801,N_3671);
nand U4576 (N_4576,N_3247,N_2138);
and U4577 (N_4577,N_2510,N_3020);
nor U4578 (N_4578,N_2245,N_3871);
xnor U4579 (N_4579,N_2870,N_3822);
and U4580 (N_4580,N_2486,N_3392);
or U4581 (N_4581,N_3535,N_2475);
and U4582 (N_4582,N_2933,N_2670);
or U4583 (N_4583,N_3992,N_2007);
nand U4584 (N_4584,N_2046,N_2415);
nand U4585 (N_4585,N_3968,N_2001);
nor U4586 (N_4586,N_2189,N_2777);
nor U4587 (N_4587,N_2201,N_3933);
nor U4588 (N_4588,N_3023,N_3656);
nor U4589 (N_4589,N_3354,N_2806);
nand U4590 (N_4590,N_3641,N_3553);
nand U4591 (N_4591,N_3435,N_3189);
or U4592 (N_4592,N_3431,N_3682);
xor U4593 (N_4593,N_3752,N_3602);
nor U4594 (N_4594,N_2175,N_2932);
nor U4595 (N_4595,N_3071,N_2337);
xor U4596 (N_4596,N_3476,N_2147);
nand U4597 (N_4597,N_3276,N_2093);
nor U4598 (N_4598,N_2000,N_2212);
and U4599 (N_4599,N_3883,N_3996);
and U4600 (N_4600,N_2118,N_3318);
nand U4601 (N_4601,N_3876,N_3828);
or U4602 (N_4602,N_3436,N_2489);
or U4603 (N_4603,N_2108,N_3963);
xnor U4604 (N_4604,N_2274,N_2268);
or U4605 (N_4605,N_3609,N_2991);
xnor U4606 (N_4606,N_2412,N_3317);
xnor U4607 (N_4607,N_2257,N_3868);
xor U4608 (N_4608,N_2908,N_2629);
and U4609 (N_4609,N_3927,N_2205);
nand U4610 (N_4610,N_2994,N_3544);
xor U4611 (N_4611,N_2042,N_3628);
and U4612 (N_4612,N_3376,N_2224);
or U4613 (N_4613,N_3705,N_2276);
and U4614 (N_4614,N_2250,N_2644);
nand U4615 (N_4615,N_3181,N_2504);
xor U4616 (N_4616,N_2608,N_3248);
or U4617 (N_4617,N_3694,N_3013);
nand U4618 (N_4618,N_2327,N_3692);
and U4619 (N_4619,N_3689,N_3108);
nor U4620 (N_4620,N_2964,N_2548);
nor U4621 (N_4621,N_2889,N_2853);
xnor U4622 (N_4622,N_3279,N_3572);
xnor U4623 (N_4623,N_3559,N_2798);
or U4624 (N_4624,N_3768,N_2154);
or U4625 (N_4625,N_2826,N_3152);
and U4626 (N_4626,N_3908,N_3140);
nand U4627 (N_4627,N_3615,N_2103);
nor U4628 (N_4628,N_3504,N_3832);
nand U4629 (N_4629,N_3220,N_2491);
or U4630 (N_4630,N_3019,N_2972);
or U4631 (N_4631,N_3035,N_3102);
or U4632 (N_4632,N_2073,N_3488);
or U4633 (N_4633,N_2182,N_2091);
and U4634 (N_4634,N_3925,N_3949);
xor U4635 (N_4635,N_3897,N_3274);
nor U4636 (N_4636,N_3280,N_2748);
nand U4637 (N_4637,N_3057,N_3919);
nand U4638 (N_4638,N_3846,N_3307);
or U4639 (N_4639,N_2883,N_3054);
nor U4640 (N_4640,N_2944,N_3939);
and U4641 (N_4641,N_3704,N_3092);
or U4642 (N_4642,N_3886,N_2198);
nand U4643 (N_4643,N_3936,N_3581);
and U4644 (N_4644,N_3417,N_2048);
xor U4645 (N_4645,N_2186,N_3238);
or U4646 (N_4646,N_3430,N_3062);
and U4647 (N_4647,N_3444,N_2169);
or U4648 (N_4648,N_2965,N_3139);
and U4649 (N_4649,N_3664,N_2136);
nand U4650 (N_4650,N_3365,N_3095);
or U4651 (N_4651,N_3030,N_3041);
nor U4652 (N_4652,N_3755,N_2392);
and U4653 (N_4653,N_3228,N_2803);
nor U4654 (N_4654,N_3473,N_2539);
nand U4655 (N_4655,N_3889,N_2167);
nor U4656 (N_4656,N_2336,N_3098);
nand U4657 (N_4657,N_3767,N_3040);
and U4658 (N_4658,N_3143,N_3970);
or U4659 (N_4659,N_3059,N_2281);
nand U4660 (N_4660,N_2237,N_3437);
nand U4661 (N_4661,N_2375,N_3479);
and U4662 (N_4662,N_3516,N_3839);
nor U4663 (N_4663,N_2707,N_3826);
nand U4664 (N_4664,N_2580,N_2900);
nor U4665 (N_4665,N_3298,N_2758);
nor U4666 (N_4666,N_3285,N_2542);
xnor U4667 (N_4667,N_3385,N_3820);
nor U4668 (N_4668,N_2210,N_3361);
or U4669 (N_4669,N_3047,N_3640);
or U4670 (N_4670,N_2463,N_2246);
nor U4671 (N_4671,N_2398,N_3006);
nor U4672 (N_4672,N_2745,N_2969);
xnor U4673 (N_4673,N_3861,N_3055);
and U4674 (N_4674,N_3475,N_3114);
nor U4675 (N_4675,N_2495,N_3960);
or U4676 (N_4676,N_3930,N_3364);
and U4677 (N_4677,N_2652,N_3713);
and U4678 (N_4678,N_2719,N_3386);
xor U4679 (N_4679,N_3636,N_2943);
nand U4680 (N_4680,N_2717,N_2731);
nand U4681 (N_4681,N_2269,N_2506);
nor U4682 (N_4682,N_2322,N_3971);
xnor U4683 (N_4683,N_2647,N_2176);
xor U4684 (N_4684,N_3109,N_2809);
or U4685 (N_4685,N_3145,N_3223);
and U4686 (N_4686,N_3910,N_3771);
and U4687 (N_4687,N_2054,N_2962);
or U4688 (N_4688,N_2980,N_2023);
or U4689 (N_4689,N_2222,N_2976);
nor U4690 (N_4690,N_3325,N_2443);
nor U4691 (N_4691,N_2445,N_2413);
nor U4692 (N_4692,N_3909,N_2465);
nand U4693 (N_4693,N_2778,N_2677);
or U4694 (N_4694,N_2300,N_2191);
or U4695 (N_4695,N_2270,N_3567);
nor U4696 (N_4696,N_2068,N_2309);
xnor U4697 (N_4697,N_2400,N_2894);
nor U4698 (N_4698,N_3758,N_3976);
xor U4699 (N_4699,N_2448,N_2417);
nor U4700 (N_4700,N_2868,N_3750);
and U4701 (N_4701,N_3726,N_3413);
xnor U4702 (N_4702,N_2421,N_2234);
or U4703 (N_4703,N_2640,N_3563);
nor U4704 (N_4704,N_3292,N_3717);
xnor U4705 (N_4705,N_2711,N_3393);
or U4706 (N_4706,N_3760,N_3746);
xor U4707 (N_4707,N_2373,N_2718);
nand U4708 (N_4708,N_3843,N_3611);
nand U4709 (N_4709,N_2598,N_3222);
xor U4710 (N_4710,N_3246,N_2840);
nor U4711 (N_4711,N_3101,N_2203);
nor U4712 (N_4712,N_3648,N_3360);
nand U4713 (N_4713,N_3787,N_3904);
nand U4714 (N_4714,N_3674,N_2990);
and U4715 (N_4715,N_2230,N_2561);
and U4716 (N_4716,N_3732,N_3323);
nand U4717 (N_4717,N_2041,N_2050);
and U4718 (N_4718,N_3410,N_2066);
nor U4719 (N_4719,N_3761,N_3522);
nand U4720 (N_4720,N_2622,N_3773);
nor U4721 (N_4721,N_2938,N_2272);
nand U4722 (N_4722,N_3551,N_3351);
or U4723 (N_4723,N_3457,N_3842);
nor U4724 (N_4724,N_3943,N_3953);
and U4725 (N_4725,N_2567,N_3487);
or U4726 (N_4726,N_2488,N_3830);
nand U4727 (N_4727,N_2262,N_3314);
nor U4728 (N_4728,N_2020,N_3588);
nand U4729 (N_4729,N_2494,N_2095);
nand U4730 (N_4730,N_2229,N_2615);
or U4731 (N_4731,N_3568,N_2155);
nor U4732 (N_4732,N_3185,N_2238);
xnor U4733 (N_4733,N_2197,N_3252);
nand U4734 (N_4734,N_2611,N_2239);
and U4735 (N_4735,N_2878,N_3574);
xnor U4736 (N_4736,N_2314,N_3296);
and U4737 (N_4737,N_2145,N_2513);
or U4738 (N_4738,N_3935,N_2975);
nand U4739 (N_4739,N_3605,N_3091);
nor U4740 (N_4740,N_3607,N_3697);
and U4741 (N_4741,N_2060,N_3792);
xor U4742 (N_4742,N_2283,N_2671);
xor U4743 (N_4743,N_3824,N_3449);
xor U4744 (N_4744,N_2508,N_2535);
and U4745 (N_4745,N_2714,N_3823);
and U4746 (N_4746,N_3721,N_2563);
or U4747 (N_4747,N_3133,N_3585);
nor U4748 (N_4748,N_3460,N_3663);
nor U4749 (N_4749,N_3150,N_3026);
and U4750 (N_4750,N_3932,N_2845);
nand U4751 (N_4751,N_3177,N_3368);
and U4752 (N_4752,N_3915,N_3434);
and U4753 (N_4753,N_3748,N_3350);
nor U4754 (N_4754,N_3201,N_2775);
nor U4755 (N_4755,N_3123,N_3142);
xor U4756 (N_4756,N_3575,N_3226);
and U4757 (N_4757,N_3866,N_3816);
and U4758 (N_4758,N_2893,N_2632);
nor U4759 (N_4759,N_3015,N_3962);
or U4760 (N_4760,N_3447,N_2951);
and U4761 (N_4761,N_2341,N_2623);
or U4762 (N_4762,N_2599,N_2875);
xor U4763 (N_4763,N_2119,N_2658);
nor U4764 (N_4764,N_3198,N_3353);
or U4765 (N_4765,N_3508,N_3918);
nor U4766 (N_4766,N_2887,N_2999);
or U4767 (N_4767,N_3309,N_3854);
nand U4768 (N_4768,N_2503,N_2720);
or U4769 (N_4769,N_3411,N_2342);
xor U4770 (N_4770,N_2594,N_3043);
xnor U4771 (N_4771,N_3756,N_3723);
and U4772 (N_4772,N_2628,N_2573);
nand U4773 (N_4773,N_2184,N_2221);
and U4774 (N_4774,N_2935,N_3499);
xnor U4775 (N_4775,N_2606,N_3657);
and U4776 (N_4776,N_2517,N_3284);
and U4777 (N_4777,N_3053,N_3560);
and U4778 (N_4778,N_2597,N_2536);
and U4779 (N_4779,N_2948,N_2797);
xor U4780 (N_4780,N_2634,N_3616);
nand U4781 (N_4781,N_2613,N_2474);
xor U4782 (N_4782,N_3402,N_3529);
nand U4783 (N_4783,N_2115,N_2153);
xnor U4784 (N_4784,N_2824,N_2660);
and U4785 (N_4785,N_2256,N_2105);
nand U4786 (N_4786,N_2788,N_3424);
or U4787 (N_4787,N_3872,N_3268);
xor U4788 (N_4788,N_2553,N_3837);
or U4789 (N_4789,N_2453,N_3075);
xnor U4790 (N_4790,N_3144,N_3678);
nor U4791 (N_4791,N_2920,N_3582);
and U4792 (N_4792,N_3683,N_2329);
or U4793 (N_4793,N_3827,N_2306);
or U4794 (N_4794,N_2819,N_3138);
nor U4795 (N_4795,N_2382,N_3763);
or U4796 (N_4796,N_3421,N_2560);
xor U4797 (N_4797,N_2570,N_2364);
nand U4798 (N_4798,N_3369,N_3116);
and U4799 (N_4799,N_3512,N_2171);
xnor U4800 (N_4800,N_3978,N_3784);
xor U4801 (N_4801,N_2721,N_3275);
or U4802 (N_4802,N_2630,N_2134);
xnor U4803 (N_4803,N_3920,N_3891);
or U4804 (N_4804,N_2209,N_2856);
nand U4805 (N_4805,N_2156,N_3738);
or U4806 (N_4806,N_2583,N_3989);
nand U4807 (N_4807,N_3494,N_2919);
or U4808 (N_4808,N_3798,N_3735);
nor U4809 (N_4809,N_2052,N_3148);
nand U4810 (N_4810,N_2386,N_2107);
and U4811 (N_4811,N_3676,N_3701);
nor U4812 (N_4812,N_3979,N_3740);
or U4813 (N_4813,N_3359,N_2346);
nor U4814 (N_4814,N_2049,N_2708);
xor U4815 (N_4815,N_3715,N_2793);
xnor U4816 (N_4816,N_2833,N_2625);
nand U4817 (N_4817,N_3685,N_3580);
or U4818 (N_4818,N_2117,N_2521);
and U4819 (N_4819,N_2363,N_2427);
and U4820 (N_4820,N_3614,N_3489);
nand U4821 (N_4821,N_3463,N_2321);
and U4822 (N_4822,N_3858,N_2408);
xor U4823 (N_4823,N_2168,N_3523);
xnor U4824 (N_4824,N_2604,N_2937);
xor U4825 (N_4825,N_2821,N_3809);
and U4826 (N_4826,N_2767,N_2177);
and U4827 (N_4827,N_3453,N_2331);
or U4828 (N_4828,N_2223,N_2805);
or U4829 (N_4829,N_2618,N_3234);
xor U4830 (N_4830,N_2655,N_2631);
and U4831 (N_4831,N_3775,N_3366);
xnor U4832 (N_4832,N_3440,N_3455);
or U4833 (N_4833,N_2918,N_2056);
nand U4834 (N_4834,N_3800,N_3009);
xnor U4835 (N_4835,N_2861,N_2387);
nand U4836 (N_4836,N_3788,N_2607);
nand U4837 (N_4837,N_3271,N_2850);
nand U4838 (N_4838,N_3926,N_2693);
or U4839 (N_4839,N_3862,N_2366);
and U4840 (N_4840,N_3921,N_3801);
nor U4841 (N_4841,N_3714,N_3042);
nand U4842 (N_4842,N_2661,N_3940);
nand U4843 (N_4843,N_3056,N_3931);
or U4844 (N_4844,N_2600,N_2869);
and U4845 (N_4845,N_2279,N_3875);
xor U4846 (N_4846,N_2009,N_2785);
nor U4847 (N_4847,N_3481,N_3022);
nor U4848 (N_4848,N_3845,N_3690);
and U4849 (N_4849,N_2844,N_3331);
nand U4850 (N_4850,N_3450,N_3728);
xor U4851 (N_4851,N_3621,N_3122);
and U4852 (N_4852,N_2786,N_2433);
or U4853 (N_4853,N_3067,N_2113);
and U4854 (N_4854,N_2446,N_2936);
xor U4855 (N_4855,N_2243,N_3929);
or U4856 (N_4856,N_2666,N_3419);
nand U4857 (N_4857,N_2149,N_3340);
nand U4858 (N_4858,N_3232,N_3587);
and U4859 (N_4859,N_3807,N_2459);
xor U4860 (N_4860,N_2830,N_3900);
xor U4861 (N_4861,N_2843,N_2313);
xor U4862 (N_4862,N_2678,N_2899);
or U4863 (N_4863,N_3964,N_3665);
nor U4864 (N_4864,N_3316,N_2402);
nand U4865 (N_4865,N_2033,N_2285);
nand U4866 (N_4866,N_2266,N_2022);
or U4867 (N_4867,N_2519,N_3565);
and U4868 (N_4868,N_3510,N_3995);
nand U4869 (N_4869,N_3503,N_2729);
and U4870 (N_4870,N_2523,N_3987);
xnor U4871 (N_4871,N_3335,N_2665);
nand U4872 (N_4872,N_3025,N_2347);
or U4873 (N_4873,N_3068,N_2114);
nor U4874 (N_4874,N_3500,N_2371);
nor U4875 (N_4875,N_2651,N_3661);
or U4876 (N_4876,N_3160,N_2642);
nand U4877 (N_4877,N_2992,N_3250);
and U4878 (N_4878,N_2228,N_2554);
nor U4879 (N_4879,N_3594,N_3586);
or U4880 (N_4880,N_2477,N_3391);
nand U4881 (N_4881,N_3474,N_3146);
and U4882 (N_4882,N_2872,N_3957);
or U4883 (N_4883,N_2565,N_3028);
nand U4884 (N_4884,N_3573,N_3183);
nand U4885 (N_4885,N_2945,N_3111);
nor U4886 (N_4886,N_3633,N_2700);
or U4887 (N_4887,N_2385,N_2829);
xor U4888 (N_4888,N_3295,N_3407);
and U4889 (N_4889,N_2452,N_3319);
or U4890 (N_4890,N_3796,N_2200);
xnor U4891 (N_4891,N_2848,N_3911);
or U4892 (N_4892,N_3794,N_2377);
xnor U4893 (N_4893,N_2751,N_3029);
or U4894 (N_4894,N_3485,N_3105);
nand U4895 (N_4895,N_3388,N_3622);
xnor U4896 (N_4896,N_3729,N_3207);
nand U4897 (N_4897,N_3853,N_2617);
nor U4898 (N_4898,N_3505,N_2735);
xnor U4899 (N_4899,N_2968,N_3749);
nand U4900 (N_4900,N_3094,N_3003);
nand U4901 (N_4901,N_2485,N_2790);
nor U4902 (N_4902,N_2814,N_2292);
nand U4903 (N_4903,N_3326,N_3533);
or U4904 (N_4904,N_2470,N_2876);
or U4905 (N_4905,N_3599,N_3593);
or U4906 (N_4906,N_3841,N_3398);
nor U4907 (N_4907,N_3334,N_2451);
and U4908 (N_4908,N_2564,N_2740);
xnor U4909 (N_4909,N_2712,N_3722);
nand U4910 (N_4910,N_2952,N_2896);
nor U4911 (N_4911,N_3958,N_2444);
and U4912 (N_4912,N_3452,N_3018);
xnor U4913 (N_4913,N_3089,N_3345);
or U4914 (N_4914,N_3149,N_2483);
xnor U4915 (N_4915,N_2927,N_2769);
xor U4916 (N_4916,N_3515,N_2846);
or U4917 (N_4917,N_2069,N_2199);
nand U4918 (N_4918,N_2955,N_3892);
nor U4919 (N_4919,N_2123,N_3004);
nor U4920 (N_4920,N_2362,N_2206);
nand U4921 (N_4921,N_2873,N_2522);
nor U4922 (N_4922,N_3265,N_2208);
and U4923 (N_4923,N_2011,N_2961);
and U4924 (N_4924,N_3840,N_3258);
nand U4925 (N_4925,N_2977,N_2255);
or U4926 (N_4926,N_2308,N_2466);
nor U4927 (N_4927,N_2921,N_2165);
nor U4928 (N_4928,N_2233,N_2121);
and U4929 (N_4929,N_2152,N_2429);
nand U4930 (N_4930,N_2691,N_3002);
nand U4931 (N_4931,N_2551,N_3534);
and U4932 (N_4932,N_2399,N_2596);
or U4933 (N_4933,N_3263,N_3038);
or U4934 (N_4934,N_2774,N_3262);
or U4935 (N_4935,N_3021,N_2348);
or U4936 (N_4936,N_3804,N_3635);
nand U4937 (N_4937,N_3045,N_2202);
xor U4938 (N_4938,N_2014,N_3103);
or U4939 (N_4939,N_3179,N_3675);
nor U4940 (N_4940,N_3708,N_2137);
xnor U4941 (N_4941,N_2592,N_2705);
nor U4942 (N_4942,N_2194,N_3942);
nor U4943 (N_4943,N_2989,N_2755);
xor U4944 (N_4944,N_3769,N_3864);
and U4945 (N_4945,N_3277,N_3982);
nand U4946 (N_4946,N_3069,N_3493);
or U4947 (N_4947,N_2578,N_2214);
nand U4948 (N_4948,N_2756,N_3390);
and U4949 (N_4949,N_2098,N_2524);
or U4950 (N_4950,N_2132,N_2129);
nor U4951 (N_4951,N_2657,N_3702);
or U4952 (N_4952,N_3835,N_3686);
nand U4953 (N_4953,N_3556,N_2770);
nand U4954 (N_4954,N_2741,N_3498);
nand U4955 (N_4955,N_3208,N_3096);
xor U4956 (N_4956,N_3356,N_3322);
xor U4957 (N_4957,N_3669,N_3812);
nand U4958 (N_4958,N_3917,N_2359);
and U4959 (N_4959,N_3776,N_2291);
nor U4960 (N_4960,N_3681,N_3206);
nand U4961 (N_4961,N_3507,N_3778);
or U4962 (N_4962,N_2550,N_2781);
or U4963 (N_4963,N_2827,N_3780);
or U4964 (N_4964,N_2911,N_2006);
xor U4965 (N_4965,N_2538,N_3526);
and U4966 (N_4966,N_2605,N_2842);
xnor U4967 (N_4967,N_3446,N_3725);
xor U4968 (N_4968,N_3106,N_3221);
nor U4969 (N_4969,N_3977,N_2641);
nor U4970 (N_4970,N_2689,N_3577);
or U4971 (N_4971,N_2822,N_3747);
or U4972 (N_4972,N_2855,N_3644);
or U4973 (N_4973,N_3304,N_2857);
xor U4974 (N_4974,N_3818,N_3313);
nand U4975 (N_4975,N_3647,N_2577);
and U4976 (N_4976,N_2380,N_3743);
or U4977 (N_4977,N_2730,N_3084);
nor U4978 (N_4978,N_2125,N_3765);
nand U4979 (N_4979,N_3912,N_3888);
nor U4980 (N_4980,N_3994,N_3461);
and U4981 (N_4981,N_3051,N_3213);
nor U4982 (N_4982,N_3655,N_2654);
and U4983 (N_4983,N_2148,N_2480);
or U4984 (N_4984,N_2795,N_3652);
and U4985 (N_4985,N_2791,N_3088);
nor U4986 (N_4986,N_3984,N_2428);
xor U4987 (N_4987,N_2817,N_2372);
xor U4988 (N_4988,N_2516,N_2930);
and U4989 (N_4989,N_3874,N_3646);
nor U4990 (N_4990,N_3518,N_2468);
xor U4991 (N_4991,N_3997,N_3881);
nor U4992 (N_4992,N_3625,N_3482);
nor U4993 (N_4993,N_2680,N_2626);
nor U4994 (N_4994,N_2260,N_2627);
or U4995 (N_4995,N_2498,N_3442);
or U4996 (N_4996,N_3543,N_2035);
and U4997 (N_4997,N_2946,N_2954);
or U4998 (N_4998,N_3072,N_2924);
nor U4999 (N_4999,N_3329,N_2749);
nand U5000 (N_5000,N_3909,N_3291);
nand U5001 (N_5001,N_2605,N_2424);
or U5002 (N_5002,N_2678,N_2071);
nor U5003 (N_5003,N_2121,N_3089);
and U5004 (N_5004,N_3055,N_3404);
and U5005 (N_5005,N_2847,N_2914);
xor U5006 (N_5006,N_2589,N_2850);
nor U5007 (N_5007,N_2250,N_3284);
or U5008 (N_5008,N_3643,N_2137);
nor U5009 (N_5009,N_3146,N_2572);
nor U5010 (N_5010,N_3751,N_3267);
or U5011 (N_5011,N_2197,N_3232);
and U5012 (N_5012,N_3747,N_2904);
nor U5013 (N_5013,N_3905,N_2005);
and U5014 (N_5014,N_3718,N_2376);
or U5015 (N_5015,N_3221,N_2219);
nor U5016 (N_5016,N_2782,N_3064);
nor U5017 (N_5017,N_3746,N_3108);
or U5018 (N_5018,N_2600,N_3405);
xor U5019 (N_5019,N_2614,N_2033);
or U5020 (N_5020,N_3308,N_3765);
nor U5021 (N_5021,N_3539,N_2850);
nor U5022 (N_5022,N_2074,N_3449);
nand U5023 (N_5023,N_2761,N_2453);
or U5024 (N_5024,N_3514,N_3299);
or U5025 (N_5025,N_2356,N_2862);
or U5026 (N_5026,N_2426,N_3529);
nand U5027 (N_5027,N_2420,N_3876);
xnor U5028 (N_5028,N_3961,N_3527);
xnor U5029 (N_5029,N_3593,N_3988);
nor U5030 (N_5030,N_3715,N_2920);
xnor U5031 (N_5031,N_3649,N_2237);
nand U5032 (N_5032,N_3245,N_2985);
xnor U5033 (N_5033,N_2069,N_3580);
and U5034 (N_5034,N_3063,N_2970);
nor U5035 (N_5035,N_3647,N_2015);
nor U5036 (N_5036,N_2274,N_3212);
nor U5037 (N_5037,N_2682,N_2252);
nand U5038 (N_5038,N_3011,N_2919);
and U5039 (N_5039,N_3067,N_2654);
nand U5040 (N_5040,N_2231,N_2275);
or U5041 (N_5041,N_3040,N_3343);
or U5042 (N_5042,N_2038,N_2306);
or U5043 (N_5043,N_3339,N_2566);
nand U5044 (N_5044,N_2027,N_2695);
or U5045 (N_5045,N_2505,N_2600);
or U5046 (N_5046,N_2053,N_3585);
nor U5047 (N_5047,N_3131,N_2653);
nor U5048 (N_5048,N_3378,N_2955);
xnor U5049 (N_5049,N_3203,N_3128);
nor U5050 (N_5050,N_2326,N_2687);
nor U5051 (N_5051,N_3104,N_3410);
and U5052 (N_5052,N_3542,N_2710);
and U5053 (N_5053,N_2399,N_2848);
nor U5054 (N_5054,N_2446,N_3797);
nor U5055 (N_5055,N_2286,N_2878);
xnor U5056 (N_5056,N_3765,N_3183);
nor U5057 (N_5057,N_2042,N_3274);
or U5058 (N_5058,N_3119,N_3415);
nand U5059 (N_5059,N_3301,N_3318);
nor U5060 (N_5060,N_3009,N_3542);
xor U5061 (N_5061,N_3304,N_3782);
nand U5062 (N_5062,N_3768,N_2327);
xor U5063 (N_5063,N_2497,N_3607);
xor U5064 (N_5064,N_2070,N_2341);
or U5065 (N_5065,N_3695,N_3711);
nand U5066 (N_5066,N_2952,N_2989);
nor U5067 (N_5067,N_3397,N_2523);
nor U5068 (N_5068,N_2374,N_3881);
nand U5069 (N_5069,N_2566,N_2509);
nor U5070 (N_5070,N_3105,N_2724);
xnor U5071 (N_5071,N_3659,N_3342);
xnor U5072 (N_5072,N_3308,N_3405);
xor U5073 (N_5073,N_2001,N_2689);
xnor U5074 (N_5074,N_3907,N_3460);
nand U5075 (N_5075,N_3309,N_3398);
xor U5076 (N_5076,N_2476,N_2322);
xor U5077 (N_5077,N_3743,N_3893);
nand U5078 (N_5078,N_3974,N_3124);
and U5079 (N_5079,N_3806,N_2261);
xnor U5080 (N_5080,N_3111,N_2607);
nor U5081 (N_5081,N_3554,N_3560);
and U5082 (N_5082,N_3117,N_3049);
nand U5083 (N_5083,N_2783,N_3623);
nand U5084 (N_5084,N_3747,N_2258);
nand U5085 (N_5085,N_3034,N_2086);
nand U5086 (N_5086,N_2752,N_3791);
or U5087 (N_5087,N_3055,N_3082);
xnor U5088 (N_5088,N_3387,N_3383);
and U5089 (N_5089,N_2346,N_2188);
nand U5090 (N_5090,N_3106,N_3060);
xnor U5091 (N_5091,N_3537,N_2607);
nor U5092 (N_5092,N_3427,N_3088);
xnor U5093 (N_5093,N_2650,N_2096);
or U5094 (N_5094,N_3701,N_3996);
xnor U5095 (N_5095,N_2834,N_2737);
nor U5096 (N_5096,N_2234,N_3593);
and U5097 (N_5097,N_3861,N_3781);
and U5098 (N_5098,N_2278,N_2280);
nand U5099 (N_5099,N_2204,N_2029);
nor U5100 (N_5100,N_3944,N_3393);
or U5101 (N_5101,N_2288,N_2131);
and U5102 (N_5102,N_2309,N_3979);
nor U5103 (N_5103,N_2049,N_2322);
and U5104 (N_5104,N_3059,N_3834);
and U5105 (N_5105,N_2743,N_2182);
xnor U5106 (N_5106,N_2001,N_3997);
xor U5107 (N_5107,N_2813,N_2423);
xor U5108 (N_5108,N_2071,N_2809);
xnor U5109 (N_5109,N_3595,N_2628);
xnor U5110 (N_5110,N_3912,N_2910);
and U5111 (N_5111,N_3617,N_2722);
xor U5112 (N_5112,N_3366,N_2237);
xor U5113 (N_5113,N_3488,N_3394);
nand U5114 (N_5114,N_3479,N_3705);
or U5115 (N_5115,N_3741,N_3877);
nand U5116 (N_5116,N_2040,N_3215);
xnor U5117 (N_5117,N_3808,N_2259);
xnor U5118 (N_5118,N_2260,N_2314);
or U5119 (N_5119,N_3673,N_3047);
or U5120 (N_5120,N_3573,N_2134);
xor U5121 (N_5121,N_3529,N_3594);
or U5122 (N_5122,N_2777,N_2628);
nand U5123 (N_5123,N_2484,N_3123);
and U5124 (N_5124,N_2317,N_3666);
and U5125 (N_5125,N_3515,N_3358);
xor U5126 (N_5126,N_2283,N_2266);
and U5127 (N_5127,N_2914,N_3469);
nand U5128 (N_5128,N_3212,N_3649);
nor U5129 (N_5129,N_2861,N_2668);
or U5130 (N_5130,N_2671,N_3732);
xor U5131 (N_5131,N_3344,N_2650);
xnor U5132 (N_5132,N_2132,N_3374);
xnor U5133 (N_5133,N_2576,N_3155);
or U5134 (N_5134,N_2573,N_2942);
and U5135 (N_5135,N_3338,N_3872);
nand U5136 (N_5136,N_2251,N_3238);
nor U5137 (N_5137,N_2655,N_3505);
nor U5138 (N_5138,N_3265,N_2998);
or U5139 (N_5139,N_2061,N_3391);
nor U5140 (N_5140,N_3122,N_2664);
or U5141 (N_5141,N_2378,N_2037);
nand U5142 (N_5142,N_3715,N_2392);
or U5143 (N_5143,N_3415,N_3315);
nor U5144 (N_5144,N_2531,N_3808);
and U5145 (N_5145,N_2311,N_2931);
nor U5146 (N_5146,N_3515,N_3796);
and U5147 (N_5147,N_2082,N_3152);
xnor U5148 (N_5148,N_3851,N_2239);
nor U5149 (N_5149,N_2989,N_2367);
nand U5150 (N_5150,N_2269,N_3576);
nand U5151 (N_5151,N_3105,N_2621);
nor U5152 (N_5152,N_2740,N_3224);
nor U5153 (N_5153,N_2213,N_2005);
nand U5154 (N_5154,N_3046,N_3302);
or U5155 (N_5155,N_2494,N_2419);
nand U5156 (N_5156,N_3707,N_2711);
nor U5157 (N_5157,N_2953,N_2981);
and U5158 (N_5158,N_3223,N_2950);
nand U5159 (N_5159,N_3029,N_3567);
nor U5160 (N_5160,N_3152,N_2725);
xor U5161 (N_5161,N_2038,N_3073);
and U5162 (N_5162,N_3846,N_3131);
or U5163 (N_5163,N_3565,N_2410);
and U5164 (N_5164,N_3069,N_2125);
nor U5165 (N_5165,N_2006,N_3831);
or U5166 (N_5166,N_2395,N_3578);
nor U5167 (N_5167,N_2321,N_3236);
nand U5168 (N_5168,N_2055,N_2081);
or U5169 (N_5169,N_3331,N_3600);
and U5170 (N_5170,N_3831,N_2799);
and U5171 (N_5171,N_3131,N_2997);
or U5172 (N_5172,N_3407,N_2562);
and U5173 (N_5173,N_3655,N_2451);
nor U5174 (N_5174,N_3369,N_3451);
nand U5175 (N_5175,N_3608,N_2728);
xnor U5176 (N_5176,N_3053,N_3199);
or U5177 (N_5177,N_3859,N_2456);
nand U5178 (N_5178,N_3764,N_2551);
and U5179 (N_5179,N_2573,N_3111);
and U5180 (N_5180,N_3420,N_2408);
nand U5181 (N_5181,N_3207,N_2075);
nand U5182 (N_5182,N_3419,N_2280);
nor U5183 (N_5183,N_2623,N_2218);
xnor U5184 (N_5184,N_2583,N_3644);
nor U5185 (N_5185,N_2127,N_3530);
xnor U5186 (N_5186,N_3790,N_3068);
and U5187 (N_5187,N_2156,N_2480);
xor U5188 (N_5188,N_3709,N_2075);
xor U5189 (N_5189,N_2511,N_3014);
and U5190 (N_5190,N_2349,N_3876);
xor U5191 (N_5191,N_3569,N_2796);
or U5192 (N_5192,N_2760,N_2991);
and U5193 (N_5193,N_3663,N_3432);
nand U5194 (N_5194,N_3374,N_3475);
xor U5195 (N_5195,N_3405,N_3828);
or U5196 (N_5196,N_2350,N_3851);
or U5197 (N_5197,N_3487,N_2825);
nor U5198 (N_5198,N_3144,N_3008);
xnor U5199 (N_5199,N_3195,N_2038);
nand U5200 (N_5200,N_2709,N_2331);
and U5201 (N_5201,N_2900,N_2088);
xor U5202 (N_5202,N_3451,N_3788);
xnor U5203 (N_5203,N_2954,N_2044);
nor U5204 (N_5204,N_3193,N_2112);
nand U5205 (N_5205,N_2284,N_3362);
nor U5206 (N_5206,N_3230,N_3157);
or U5207 (N_5207,N_3447,N_3085);
nand U5208 (N_5208,N_3031,N_3932);
xnor U5209 (N_5209,N_3892,N_3697);
nand U5210 (N_5210,N_3451,N_2130);
nor U5211 (N_5211,N_3026,N_2119);
or U5212 (N_5212,N_2651,N_3791);
nor U5213 (N_5213,N_3106,N_3188);
nand U5214 (N_5214,N_2208,N_2321);
xor U5215 (N_5215,N_3854,N_2097);
and U5216 (N_5216,N_2015,N_3848);
nor U5217 (N_5217,N_3802,N_3914);
and U5218 (N_5218,N_2637,N_2010);
and U5219 (N_5219,N_2468,N_3418);
xnor U5220 (N_5220,N_2332,N_3491);
nand U5221 (N_5221,N_2848,N_3099);
and U5222 (N_5222,N_3912,N_3275);
nor U5223 (N_5223,N_2482,N_2223);
or U5224 (N_5224,N_3658,N_3555);
and U5225 (N_5225,N_2447,N_3865);
nand U5226 (N_5226,N_3066,N_2652);
or U5227 (N_5227,N_2179,N_3499);
xor U5228 (N_5228,N_3744,N_3024);
or U5229 (N_5229,N_3610,N_2287);
nand U5230 (N_5230,N_2220,N_3654);
nand U5231 (N_5231,N_3914,N_2313);
xor U5232 (N_5232,N_3111,N_2932);
and U5233 (N_5233,N_2031,N_2662);
xor U5234 (N_5234,N_3033,N_3077);
nand U5235 (N_5235,N_3454,N_3913);
xor U5236 (N_5236,N_3430,N_2507);
nand U5237 (N_5237,N_3619,N_3775);
xor U5238 (N_5238,N_3039,N_3595);
xnor U5239 (N_5239,N_2711,N_3870);
and U5240 (N_5240,N_3123,N_2968);
and U5241 (N_5241,N_2274,N_2032);
nor U5242 (N_5242,N_3007,N_3174);
nand U5243 (N_5243,N_2722,N_3211);
nor U5244 (N_5244,N_2234,N_3677);
and U5245 (N_5245,N_2115,N_2748);
nand U5246 (N_5246,N_3375,N_3519);
or U5247 (N_5247,N_3742,N_2324);
xor U5248 (N_5248,N_2071,N_2202);
xnor U5249 (N_5249,N_2576,N_3477);
nor U5250 (N_5250,N_3806,N_3641);
nor U5251 (N_5251,N_3741,N_2857);
nand U5252 (N_5252,N_3320,N_3633);
nor U5253 (N_5253,N_3846,N_3964);
and U5254 (N_5254,N_2770,N_3704);
nor U5255 (N_5255,N_3492,N_2808);
and U5256 (N_5256,N_3078,N_2169);
or U5257 (N_5257,N_3798,N_2401);
or U5258 (N_5258,N_3049,N_3915);
and U5259 (N_5259,N_3470,N_3161);
xnor U5260 (N_5260,N_3685,N_3328);
xnor U5261 (N_5261,N_3675,N_2804);
or U5262 (N_5262,N_2130,N_3471);
nand U5263 (N_5263,N_2900,N_2823);
or U5264 (N_5264,N_3903,N_2929);
nor U5265 (N_5265,N_2627,N_3622);
nand U5266 (N_5266,N_3624,N_3690);
nor U5267 (N_5267,N_2442,N_3168);
xnor U5268 (N_5268,N_2284,N_2476);
nand U5269 (N_5269,N_3309,N_3344);
or U5270 (N_5270,N_2564,N_2784);
xor U5271 (N_5271,N_2826,N_2108);
nor U5272 (N_5272,N_3102,N_2500);
nand U5273 (N_5273,N_3232,N_3940);
nor U5274 (N_5274,N_2650,N_3589);
and U5275 (N_5275,N_3158,N_3201);
xnor U5276 (N_5276,N_3287,N_2959);
nand U5277 (N_5277,N_2813,N_2917);
xnor U5278 (N_5278,N_2032,N_2024);
or U5279 (N_5279,N_2553,N_2116);
nand U5280 (N_5280,N_3718,N_3768);
or U5281 (N_5281,N_3529,N_2290);
or U5282 (N_5282,N_2526,N_3698);
or U5283 (N_5283,N_2546,N_2507);
and U5284 (N_5284,N_3955,N_3840);
nand U5285 (N_5285,N_2485,N_3795);
nand U5286 (N_5286,N_2803,N_3283);
or U5287 (N_5287,N_2956,N_2039);
or U5288 (N_5288,N_3078,N_3051);
and U5289 (N_5289,N_2146,N_3386);
xor U5290 (N_5290,N_2345,N_2064);
or U5291 (N_5291,N_3313,N_3497);
nand U5292 (N_5292,N_2050,N_3729);
or U5293 (N_5293,N_2689,N_3470);
or U5294 (N_5294,N_2547,N_3018);
nand U5295 (N_5295,N_3598,N_3409);
nor U5296 (N_5296,N_2553,N_2987);
nor U5297 (N_5297,N_2769,N_2514);
nor U5298 (N_5298,N_2535,N_3094);
nor U5299 (N_5299,N_3461,N_2313);
and U5300 (N_5300,N_2057,N_2149);
and U5301 (N_5301,N_2556,N_2717);
or U5302 (N_5302,N_3598,N_2992);
xor U5303 (N_5303,N_2369,N_2777);
or U5304 (N_5304,N_2475,N_2611);
nand U5305 (N_5305,N_2490,N_3308);
xor U5306 (N_5306,N_2158,N_2907);
or U5307 (N_5307,N_3878,N_3237);
nand U5308 (N_5308,N_2540,N_3606);
nand U5309 (N_5309,N_2668,N_3241);
nor U5310 (N_5310,N_3657,N_3883);
xnor U5311 (N_5311,N_2285,N_2260);
nand U5312 (N_5312,N_2539,N_3375);
nand U5313 (N_5313,N_3204,N_2495);
or U5314 (N_5314,N_2426,N_2953);
nand U5315 (N_5315,N_3695,N_2119);
or U5316 (N_5316,N_3442,N_2810);
xor U5317 (N_5317,N_2168,N_2581);
and U5318 (N_5318,N_3242,N_3157);
or U5319 (N_5319,N_2238,N_2563);
and U5320 (N_5320,N_2035,N_3188);
nor U5321 (N_5321,N_2090,N_3365);
nand U5322 (N_5322,N_3897,N_3969);
and U5323 (N_5323,N_2482,N_2940);
or U5324 (N_5324,N_3884,N_3086);
and U5325 (N_5325,N_2946,N_3120);
nor U5326 (N_5326,N_3749,N_3213);
xnor U5327 (N_5327,N_2267,N_2899);
nand U5328 (N_5328,N_2509,N_3899);
nand U5329 (N_5329,N_3103,N_2258);
nor U5330 (N_5330,N_3764,N_3825);
and U5331 (N_5331,N_3369,N_2637);
nor U5332 (N_5332,N_3375,N_2920);
xor U5333 (N_5333,N_3327,N_3039);
or U5334 (N_5334,N_2555,N_2299);
or U5335 (N_5335,N_2756,N_3310);
xnor U5336 (N_5336,N_2066,N_2666);
xor U5337 (N_5337,N_2092,N_3300);
or U5338 (N_5338,N_3694,N_3098);
or U5339 (N_5339,N_3269,N_2188);
and U5340 (N_5340,N_3517,N_2679);
and U5341 (N_5341,N_3657,N_2620);
nand U5342 (N_5342,N_2328,N_2041);
nand U5343 (N_5343,N_2471,N_3232);
nand U5344 (N_5344,N_3495,N_3147);
and U5345 (N_5345,N_3832,N_2790);
or U5346 (N_5346,N_3036,N_3914);
xnor U5347 (N_5347,N_2911,N_2079);
and U5348 (N_5348,N_3919,N_2123);
nor U5349 (N_5349,N_2865,N_2262);
nor U5350 (N_5350,N_2485,N_2618);
nand U5351 (N_5351,N_3292,N_3556);
xnor U5352 (N_5352,N_2217,N_2024);
nand U5353 (N_5353,N_2925,N_2581);
nor U5354 (N_5354,N_3571,N_2813);
and U5355 (N_5355,N_3345,N_3353);
or U5356 (N_5356,N_2375,N_3210);
or U5357 (N_5357,N_3756,N_3773);
xor U5358 (N_5358,N_3124,N_2138);
nor U5359 (N_5359,N_3837,N_3901);
and U5360 (N_5360,N_3795,N_3261);
and U5361 (N_5361,N_2055,N_3578);
or U5362 (N_5362,N_2610,N_2062);
nor U5363 (N_5363,N_3113,N_3343);
and U5364 (N_5364,N_2719,N_2969);
nor U5365 (N_5365,N_3874,N_2376);
nor U5366 (N_5366,N_2074,N_3368);
nor U5367 (N_5367,N_3668,N_2252);
nor U5368 (N_5368,N_2053,N_2657);
and U5369 (N_5369,N_3571,N_3665);
or U5370 (N_5370,N_2028,N_2200);
nor U5371 (N_5371,N_3040,N_2150);
or U5372 (N_5372,N_2812,N_2252);
nand U5373 (N_5373,N_2988,N_2514);
nor U5374 (N_5374,N_2471,N_2113);
nand U5375 (N_5375,N_2116,N_2587);
nand U5376 (N_5376,N_3980,N_2636);
and U5377 (N_5377,N_3376,N_3031);
nor U5378 (N_5378,N_2014,N_3126);
nand U5379 (N_5379,N_3246,N_2797);
xor U5380 (N_5380,N_2003,N_3469);
nand U5381 (N_5381,N_2963,N_3422);
or U5382 (N_5382,N_3020,N_3746);
nand U5383 (N_5383,N_3759,N_3717);
or U5384 (N_5384,N_3039,N_2512);
or U5385 (N_5385,N_3268,N_3597);
or U5386 (N_5386,N_2511,N_2022);
nor U5387 (N_5387,N_2102,N_2635);
nor U5388 (N_5388,N_3317,N_3957);
nand U5389 (N_5389,N_2849,N_3004);
nor U5390 (N_5390,N_3182,N_3380);
xnor U5391 (N_5391,N_2636,N_2451);
nand U5392 (N_5392,N_3529,N_2634);
nand U5393 (N_5393,N_2114,N_3634);
or U5394 (N_5394,N_3524,N_3500);
nor U5395 (N_5395,N_3553,N_3346);
and U5396 (N_5396,N_3780,N_3686);
nand U5397 (N_5397,N_3003,N_3656);
nor U5398 (N_5398,N_3555,N_2709);
or U5399 (N_5399,N_3080,N_3546);
xor U5400 (N_5400,N_3013,N_3582);
nand U5401 (N_5401,N_3461,N_2092);
and U5402 (N_5402,N_3186,N_3680);
and U5403 (N_5403,N_3033,N_3768);
or U5404 (N_5404,N_3950,N_2540);
xor U5405 (N_5405,N_3650,N_2376);
xnor U5406 (N_5406,N_3614,N_3056);
or U5407 (N_5407,N_2933,N_2411);
or U5408 (N_5408,N_3800,N_3704);
nor U5409 (N_5409,N_2620,N_3010);
or U5410 (N_5410,N_2635,N_3950);
or U5411 (N_5411,N_2575,N_2876);
or U5412 (N_5412,N_3826,N_2523);
xnor U5413 (N_5413,N_3169,N_2493);
nor U5414 (N_5414,N_2255,N_2665);
or U5415 (N_5415,N_2395,N_2457);
and U5416 (N_5416,N_3752,N_3710);
or U5417 (N_5417,N_3561,N_3212);
nor U5418 (N_5418,N_3532,N_2060);
nand U5419 (N_5419,N_3264,N_3541);
nand U5420 (N_5420,N_2719,N_2034);
nor U5421 (N_5421,N_2644,N_3704);
nor U5422 (N_5422,N_2616,N_3123);
nand U5423 (N_5423,N_2078,N_3178);
nand U5424 (N_5424,N_3996,N_3065);
nor U5425 (N_5425,N_3278,N_2549);
xnor U5426 (N_5426,N_2218,N_2367);
xnor U5427 (N_5427,N_3258,N_2479);
nand U5428 (N_5428,N_2212,N_2495);
and U5429 (N_5429,N_3327,N_2716);
nor U5430 (N_5430,N_3057,N_3047);
or U5431 (N_5431,N_2710,N_3007);
nor U5432 (N_5432,N_3434,N_2050);
nand U5433 (N_5433,N_2644,N_3530);
nor U5434 (N_5434,N_2076,N_2888);
nor U5435 (N_5435,N_2332,N_3948);
nand U5436 (N_5436,N_3196,N_2312);
xnor U5437 (N_5437,N_2819,N_2269);
xnor U5438 (N_5438,N_3543,N_3110);
and U5439 (N_5439,N_3295,N_3375);
and U5440 (N_5440,N_3057,N_3292);
nor U5441 (N_5441,N_3255,N_2343);
nand U5442 (N_5442,N_2270,N_3373);
nand U5443 (N_5443,N_2576,N_3299);
xor U5444 (N_5444,N_2781,N_2582);
and U5445 (N_5445,N_2509,N_3554);
and U5446 (N_5446,N_2506,N_3347);
nor U5447 (N_5447,N_3634,N_2804);
xor U5448 (N_5448,N_2828,N_2150);
or U5449 (N_5449,N_2108,N_3365);
xnor U5450 (N_5450,N_2877,N_2493);
nand U5451 (N_5451,N_2027,N_3895);
nand U5452 (N_5452,N_2292,N_3331);
and U5453 (N_5453,N_2564,N_2833);
or U5454 (N_5454,N_2287,N_2996);
and U5455 (N_5455,N_3199,N_2072);
or U5456 (N_5456,N_3778,N_3849);
or U5457 (N_5457,N_3742,N_2680);
nor U5458 (N_5458,N_2965,N_3581);
xnor U5459 (N_5459,N_2822,N_3444);
or U5460 (N_5460,N_3730,N_2393);
and U5461 (N_5461,N_2508,N_2485);
nand U5462 (N_5462,N_3100,N_2261);
nor U5463 (N_5463,N_2480,N_3438);
nor U5464 (N_5464,N_3113,N_3298);
or U5465 (N_5465,N_2136,N_2429);
xnor U5466 (N_5466,N_2814,N_2183);
or U5467 (N_5467,N_2788,N_2678);
nand U5468 (N_5468,N_2982,N_2689);
nor U5469 (N_5469,N_3052,N_3276);
nand U5470 (N_5470,N_3291,N_2946);
or U5471 (N_5471,N_2171,N_2701);
xor U5472 (N_5472,N_3004,N_3009);
xnor U5473 (N_5473,N_2525,N_3381);
and U5474 (N_5474,N_2846,N_3252);
nor U5475 (N_5475,N_2494,N_3446);
and U5476 (N_5476,N_2995,N_3537);
nand U5477 (N_5477,N_3301,N_2434);
nor U5478 (N_5478,N_3495,N_2008);
xnor U5479 (N_5479,N_3453,N_3790);
nor U5480 (N_5480,N_2067,N_3703);
nand U5481 (N_5481,N_2044,N_3936);
xor U5482 (N_5482,N_3436,N_2239);
nand U5483 (N_5483,N_2380,N_3595);
or U5484 (N_5484,N_3149,N_2036);
nor U5485 (N_5485,N_2707,N_3075);
and U5486 (N_5486,N_3880,N_3660);
nand U5487 (N_5487,N_3536,N_3226);
nor U5488 (N_5488,N_2816,N_2070);
nor U5489 (N_5489,N_2847,N_3016);
xor U5490 (N_5490,N_3329,N_3074);
or U5491 (N_5491,N_3476,N_3077);
nor U5492 (N_5492,N_3422,N_2768);
and U5493 (N_5493,N_3927,N_2915);
nand U5494 (N_5494,N_3582,N_2245);
xor U5495 (N_5495,N_3530,N_2573);
xnor U5496 (N_5496,N_3605,N_3009);
nor U5497 (N_5497,N_2905,N_3684);
nand U5498 (N_5498,N_2923,N_3847);
nand U5499 (N_5499,N_2754,N_2427);
or U5500 (N_5500,N_3462,N_3949);
xor U5501 (N_5501,N_2323,N_3811);
nand U5502 (N_5502,N_3945,N_3161);
nand U5503 (N_5503,N_2273,N_2691);
or U5504 (N_5504,N_3856,N_2949);
and U5505 (N_5505,N_3888,N_2346);
or U5506 (N_5506,N_2269,N_3991);
nand U5507 (N_5507,N_2522,N_3956);
xor U5508 (N_5508,N_3036,N_2789);
xor U5509 (N_5509,N_3689,N_2388);
xnor U5510 (N_5510,N_2879,N_3355);
nand U5511 (N_5511,N_2411,N_3928);
nand U5512 (N_5512,N_3379,N_3283);
nor U5513 (N_5513,N_2504,N_2675);
nor U5514 (N_5514,N_3127,N_3328);
xnor U5515 (N_5515,N_3496,N_3605);
xor U5516 (N_5516,N_2417,N_3654);
nor U5517 (N_5517,N_2190,N_3978);
and U5518 (N_5518,N_2370,N_2987);
xnor U5519 (N_5519,N_2471,N_3219);
xor U5520 (N_5520,N_3717,N_2995);
xor U5521 (N_5521,N_2162,N_2650);
nand U5522 (N_5522,N_2536,N_3133);
xnor U5523 (N_5523,N_3863,N_2151);
nor U5524 (N_5524,N_3254,N_2572);
or U5525 (N_5525,N_3813,N_3750);
xor U5526 (N_5526,N_3050,N_2117);
or U5527 (N_5527,N_3473,N_2736);
xnor U5528 (N_5528,N_3382,N_3432);
and U5529 (N_5529,N_2483,N_2746);
xor U5530 (N_5530,N_2474,N_2621);
and U5531 (N_5531,N_3488,N_3887);
and U5532 (N_5532,N_2592,N_2103);
and U5533 (N_5533,N_3794,N_3407);
nor U5534 (N_5534,N_2745,N_3148);
nand U5535 (N_5535,N_3895,N_3222);
nand U5536 (N_5536,N_2740,N_2686);
nor U5537 (N_5537,N_2225,N_2194);
or U5538 (N_5538,N_3817,N_3677);
or U5539 (N_5539,N_3486,N_3106);
or U5540 (N_5540,N_3930,N_3850);
nor U5541 (N_5541,N_3394,N_2761);
and U5542 (N_5542,N_2926,N_3460);
nand U5543 (N_5543,N_2298,N_2864);
or U5544 (N_5544,N_3296,N_2009);
nor U5545 (N_5545,N_2483,N_2138);
or U5546 (N_5546,N_3856,N_2513);
nand U5547 (N_5547,N_2297,N_2647);
and U5548 (N_5548,N_3548,N_3411);
and U5549 (N_5549,N_2467,N_2604);
xor U5550 (N_5550,N_2244,N_2465);
nand U5551 (N_5551,N_3392,N_3620);
nand U5552 (N_5552,N_2175,N_2811);
xnor U5553 (N_5553,N_2282,N_2261);
or U5554 (N_5554,N_2535,N_3596);
and U5555 (N_5555,N_2945,N_2221);
xor U5556 (N_5556,N_3513,N_3983);
and U5557 (N_5557,N_2991,N_2279);
nand U5558 (N_5558,N_2249,N_2572);
nor U5559 (N_5559,N_3288,N_3187);
nand U5560 (N_5560,N_3219,N_3661);
xor U5561 (N_5561,N_2061,N_3721);
and U5562 (N_5562,N_3398,N_3270);
nor U5563 (N_5563,N_2993,N_2485);
and U5564 (N_5564,N_2549,N_2006);
nand U5565 (N_5565,N_2248,N_2242);
or U5566 (N_5566,N_2616,N_3731);
and U5567 (N_5567,N_2547,N_2738);
and U5568 (N_5568,N_3321,N_3311);
nor U5569 (N_5569,N_3651,N_2187);
nor U5570 (N_5570,N_3264,N_3462);
and U5571 (N_5571,N_2278,N_3586);
or U5572 (N_5572,N_2519,N_2859);
and U5573 (N_5573,N_3221,N_3134);
nor U5574 (N_5574,N_2438,N_3732);
xnor U5575 (N_5575,N_3250,N_2392);
xnor U5576 (N_5576,N_3661,N_3851);
or U5577 (N_5577,N_3809,N_2798);
xor U5578 (N_5578,N_2814,N_2378);
or U5579 (N_5579,N_2983,N_3882);
and U5580 (N_5580,N_3648,N_2907);
nand U5581 (N_5581,N_2497,N_3865);
nor U5582 (N_5582,N_2011,N_2096);
and U5583 (N_5583,N_3873,N_2373);
xnor U5584 (N_5584,N_2501,N_2356);
xnor U5585 (N_5585,N_2212,N_3024);
nor U5586 (N_5586,N_3430,N_3280);
and U5587 (N_5587,N_3175,N_3546);
and U5588 (N_5588,N_3790,N_2475);
or U5589 (N_5589,N_3079,N_2989);
nand U5590 (N_5590,N_2382,N_2490);
and U5591 (N_5591,N_3154,N_2395);
nand U5592 (N_5592,N_3428,N_3074);
and U5593 (N_5593,N_2740,N_3400);
or U5594 (N_5594,N_3398,N_3902);
and U5595 (N_5595,N_2182,N_3111);
xnor U5596 (N_5596,N_2357,N_2491);
nor U5597 (N_5597,N_2651,N_3905);
nor U5598 (N_5598,N_3465,N_2438);
xor U5599 (N_5599,N_2700,N_2172);
and U5600 (N_5600,N_3872,N_2575);
and U5601 (N_5601,N_3805,N_2365);
nor U5602 (N_5602,N_2806,N_2766);
nand U5603 (N_5603,N_2096,N_2214);
and U5604 (N_5604,N_3692,N_3179);
or U5605 (N_5605,N_3780,N_2332);
xnor U5606 (N_5606,N_2043,N_2391);
xnor U5607 (N_5607,N_2920,N_3150);
nor U5608 (N_5608,N_3424,N_2926);
or U5609 (N_5609,N_2043,N_2028);
nor U5610 (N_5610,N_2900,N_2601);
or U5611 (N_5611,N_3527,N_3285);
or U5612 (N_5612,N_2932,N_3903);
nand U5613 (N_5613,N_3489,N_3145);
and U5614 (N_5614,N_2345,N_3051);
xor U5615 (N_5615,N_3246,N_2833);
xor U5616 (N_5616,N_3908,N_3289);
nor U5617 (N_5617,N_2443,N_2711);
nand U5618 (N_5618,N_2647,N_2079);
and U5619 (N_5619,N_2352,N_2778);
nand U5620 (N_5620,N_2237,N_2692);
and U5621 (N_5621,N_3275,N_3075);
or U5622 (N_5622,N_2759,N_3909);
nor U5623 (N_5623,N_3952,N_2724);
or U5624 (N_5624,N_3739,N_2632);
or U5625 (N_5625,N_3839,N_2690);
and U5626 (N_5626,N_3957,N_3102);
nor U5627 (N_5627,N_3038,N_2672);
xnor U5628 (N_5628,N_2549,N_3857);
nand U5629 (N_5629,N_3212,N_2537);
and U5630 (N_5630,N_3988,N_3940);
nor U5631 (N_5631,N_3160,N_2555);
nand U5632 (N_5632,N_2105,N_3173);
nor U5633 (N_5633,N_2053,N_2442);
or U5634 (N_5634,N_2186,N_2958);
xor U5635 (N_5635,N_2271,N_2154);
xor U5636 (N_5636,N_2307,N_3743);
nor U5637 (N_5637,N_3535,N_3653);
xnor U5638 (N_5638,N_2932,N_2023);
nor U5639 (N_5639,N_2038,N_2063);
nand U5640 (N_5640,N_2810,N_2575);
xor U5641 (N_5641,N_2830,N_2645);
xnor U5642 (N_5642,N_3465,N_3571);
xnor U5643 (N_5643,N_3930,N_3165);
xnor U5644 (N_5644,N_3747,N_2869);
or U5645 (N_5645,N_2956,N_2341);
and U5646 (N_5646,N_3624,N_3628);
nor U5647 (N_5647,N_2951,N_3362);
or U5648 (N_5648,N_2039,N_2191);
xnor U5649 (N_5649,N_3562,N_3431);
nand U5650 (N_5650,N_2182,N_3523);
nand U5651 (N_5651,N_2612,N_2608);
and U5652 (N_5652,N_3714,N_3207);
nor U5653 (N_5653,N_3221,N_3351);
xor U5654 (N_5654,N_2609,N_3609);
xor U5655 (N_5655,N_3918,N_3471);
xnor U5656 (N_5656,N_3284,N_2745);
or U5657 (N_5657,N_2634,N_3282);
or U5658 (N_5658,N_2859,N_2103);
nand U5659 (N_5659,N_3672,N_3434);
xnor U5660 (N_5660,N_2124,N_3055);
and U5661 (N_5661,N_2606,N_3111);
xnor U5662 (N_5662,N_2847,N_3296);
xor U5663 (N_5663,N_3465,N_3569);
and U5664 (N_5664,N_3288,N_3396);
or U5665 (N_5665,N_3826,N_3854);
nor U5666 (N_5666,N_3573,N_2386);
xnor U5667 (N_5667,N_3616,N_3068);
and U5668 (N_5668,N_2054,N_2306);
nor U5669 (N_5669,N_2954,N_3990);
or U5670 (N_5670,N_3892,N_3078);
and U5671 (N_5671,N_2120,N_3181);
and U5672 (N_5672,N_3101,N_2979);
xor U5673 (N_5673,N_2078,N_3395);
xnor U5674 (N_5674,N_2791,N_2354);
and U5675 (N_5675,N_2702,N_3565);
nor U5676 (N_5676,N_2298,N_3818);
or U5677 (N_5677,N_2933,N_2242);
xnor U5678 (N_5678,N_2398,N_3763);
and U5679 (N_5679,N_3516,N_3991);
nand U5680 (N_5680,N_3336,N_2095);
xnor U5681 (N_5681,N_2134,N_3899);
and U5682 (N_5682,N_2084,N_2194);
xor U5683 (N_5683,N_3273,N_3949);
and U5684 (N_5684,N_3036,N_3101);
nor U5685 (N_5685,N_3872,N_2098);
or U5686 (N_5686,N_3000,N_2871);
or U5687 (N_5687,N_3423,N_2547);
xor U5688 (N_5688,N_3940,N_3312);
nand U5689 (N_5689,N_2759,N_3099);
nand U5690 (N_5690,N_3751,N_2815);
nor U5691 (N_5691,N_3448,N_2501);
or U5692 (N_5692,N_2300,N_2342);
xnor U5693 (N_5693,N_2961,N_2821);
xnor U5694 (N_5694,N_3596,N_2363);
nand U5695 (N_5695,N_3920,N_2239);
xor U5696 (N_5696,N_2230,N_3310);
xor U5697 (N_5697,N_2267,N_3966);
xor U5698 (N_5698,N_3520,N_3735);
or U5699 (N_5699,N_3645,N_2592);
xor U5700 (N_5700,N_3492,N_2565);
and U5701 (N_5701,N_3583,N_3386);
nand U5702 (N_5702,N_3381,N_3584);
or U5703 (N_5703,N_2976,N_2583);
nor U5704 (N_5704,N_2179,N_3926);
xor U5705 (N_5705,N_3477,N_3626);
nand U5706 (N_5706,N_2853,N_2477);
and U5707 (N_5707,N_3925,N_3081);
nand U5708 (N_5708,N_3474,N_3959);
and U5709 (N_5709,N_3092,N_2895);
nor U5710 (N_5710,N_3284,N_2953);
or U5711 (N_5711,N_2470,N_2560);
nor U5712 (N_5712,N_3990,N_2353);
nand U5713 (N_5713,N_3806,N_3344);
and U5714 (N_5714,N_3022,N_3624);
or U5715 (N_5715,N_3412,N_3572);
nor U5716 (N_5716,N_2530,N_2502);
or U5717 (N_5717,N_3158,N_2990);
xnor U5718 (N_5718,N_3044,N_2890);
xnor U5719 (N_5719,N_2380,N_2839);
nand U5720 (N_5720,N_3201,N_2984);
and U5721 (N_5721,N_3275,N_3902);
and U5722 (N_5722,N_2963,N_2648);
nand U5723 (N_5723,N_3916,N_2741);
or U5724 (N_5724,N_3160,N_2443);
or U5725 (N_5725,N_3284,N_3275);
and U5726 (N_5726,N_2893,N_2773);
nand U5727 (N_5727,N_2112,N_3752);
or U5728 (N_5728,N_3616,N_3605);
and U5729 (N_5729,N_3435,N_3111);
nand U5730 (N_5730,N_2490,N_2410);
xnor U5731 (N_5731,N_2477,N_2777);
nand U5732 (N_5732,N_3004,N_2931);
and U5733 (N_5733,N_3007,N_2989);
and U5734 (N_5734,N_2804,N_2736);
or U5735 (N_5735,N_3283,N_2608);
and U5736 (N_5736,N_2099,N_2382);
nor U5737 (N_5737,N_2172,N_3221);
nand U5738 (N_5738,N_2928,N_2946);
or U5739 (N_5739,N_2592,N_3743);
or U5740 (N_5740,N_2104,N_2033);
nand U5741 (N_5741,N_2897,N_3047);
nand U5742 (N_5742,N_3379,N_3649);
nor U5743 (N_5743,N_3922,N_3963);
xor U5744 (N_5744,N_3057,N_2764);
and U5745 (N_5745,N_2282,N_3276);
nand U5746 (N_5746,N_2872,N_3746);
xor U5747 (N_5747,N_3742,N_3459);
or U5748 (N_5748,N_3719,N_2838);
xor U5749 (N_5749,N_3423,N_2400);
or U5750 (N_5750,N_2196,N_2078);
nand U5751 (N_5751,N_3274,N_3562);
xor U5752 (N_5752,N_3629,N_2346);
or U5753 (N_5753,N_2795,N_2519);
and U5754 (N_5754,N_2365,N_2449);
nand U5755 (N_5755,N_2554,N_3259);
xnor U5756 (N_5756,N_3390,N_2459);
nor U5757 (N_5757,N_3670,N_2807);
and U5758 (N_5758,N_3842,N_2520);
xor U5759 (N_5759,N_2133,N_2734);
and U5760 (N_5760,N_2590,N_3080);
or U5761 (N_5761,N_2502,N_3028);
and U5762 (N_5762,N_3343,N_2498);
xnor U5763 (N_5763,N_2234,N_3772);
and U5764 (N_5764,N_3336,N_2186);
or U5765 (N_5765,N_3458,N_2628);
xor U5766 (N_5766,N_3291,N_2839);
nand U5767 (N_5767,N_3911,N_3051);
xnor U5768 (N_5768,N_2479,N_3464);
or U5769 (N_5769,N_2190,N_3039);
or U5770 (N_5770,N_3396,N_2333);
nand U5771 (N_5771,N_2080,N_2028);
nand U5772 (N_5772,N_2730,N_2295);
xor U5773 (N_5773,N_3189,N_3490);
and U5774 (N_5774,N_3494,N_2015);
nand U5775 (N_5775,N_2884,N_3919);
nor U5776 (N_5776,N_2618,N_3290);
xnor U5777 (N_5777,N_2158,N_2487);
and U5778 (N_5778,N_3594,N_3580);
and U5779 (N_5779,N_2437,N_2622);
or U5780 (N_5780,N_2431,N_3334);
or U5781 (N_5781,N_2782,N_3307);
nand U5782 (N_5782,N_3928,N_2184);
or U5783 (N_5783,N_2094,N_3794);
or U5784 (N_5784,N_2024,N_2448);
nor U5785 (N_5785,N_3573,N_2006);
and U5786 (N_5786,N_2061,N_3169);
or U5787 (N_5787,N_2916,N_3234);
nand U5788 (N_5788,N_2255,N_2409);
or U5789 (N_5789,N_3202,N_2562);
xnor U5790 (N_5790,N_3770,N_3439);
nand U5791 (N_5791,N_3028,N_2364);
and U5792 (N_5792,N_2863,N_3763);
and U5793 (N_5793,N_3538,N_3544);
nand U5794 (N_5794,N_2697,N_2590);
nand U5795 (N_5795,N_2783,N_2614);
nor U5796 (N_5796,N_2244,N_3612);
xnor U5797 (N_5797,N_2653,N_3413);
nand U5798 (N_5798,N_3116,N_2975);
nor U5799 (N_5799,N_2788,N_2192);
nand U5800 (N_5800,N_2091,N_3831);
or U5801 (N_5801,N_3918,N_2664);
and U5802 (N_5802,N_3491,N_3390);
and U5803 (N_5803,N_2202,N_2564);
xnor U5804 (N_5804,N_3684,N_3254);
and U5805 (N_5805,N_3960,N_3356);
or U5806 (N_5806,N_3390,N_3861);
or U5807 (N_5807,N_2852,N_3536);
xor U5808 (N_5808,N_2409,N_3298);
nand U5809 (N_5809,N_2394,N_2047);
nand U5810 (N_5810,N_2925,N_3700);
and U5811 (N_5811,N_3479,N_2928);
nor U5812 (N_5812,N_3158,N_3054);
or U5813 (N_5813,N_3778,N_3863);
nor U5814 (N_5814,N_3901,N_2852);
nand U5815 (N_5815,N_2719,N_3239);
xor U5816 (N_5816,N_2687,N_3226);
and U5817 (N_5817,N_3201,N_2117);
and U5818 (N_5818,N_3215,N_3900);
nand U5819 (N_5819,N_3605,N_2877);
xnor U5820 (N_5820,N_2715,N_3057);
nand U5821 (N_5821,N_2045,N_3174);
or U5822 (N_5822,N_2941,N_3934);
nand U5823 (N_5823,N_3875,N_2369);
and U5824 (N_5824,N_2021,N_2755);
nand U5825 (N_5825,N_2472,N_3480);
xor U5826 (N_5826,N_3649,N_2040);
nor U5827 (N_5827,N_3639,N_2498);
nor U5828 (N_5828,N_2318,N_3712);
nand U5829 (N_5829,N_3237,N_3416);
xnor U5830 (N_5830,N_3922,N_2726);
xor U5831 (N_5831,N_2981,N_2765);
and U5832 (N_5832,N_3700,N_3711);
or U5833 (N_5833,N_2382,N_3748);
nor U5834 (N_5834,N_2498,N_2220);
and U5835 (N_5835,N_2443,N_3882);
or U5836 (N_5836,N_3369,N_3351);
nor U5837 (N_5837,N_3471,N_2212);
or U5838 (N_5838,N_3583,N_2996);
xnor U5839 (N_5839,N_2420,N_2458);
xor U5840 (N_5840,N_3263,N_3077);
or U5841 (N_5841,N_3513,N_3653);
xor U5842 (N_5842,N_2064,N_2948);
nand U5843 (N_5843,N_2502,N_2001);
xnor U5844 (N_5844,N_2292,N_2454);
or U5845 (N_5845,N_3958,N_2894);
nand U5846 (N_5846,N_2440,N_2009);
xor U5847 (N_5847,N_2933,N_2649);
nand U5848 (N_5848,N_2168,N_3825);
and U5849 (N_5849,N_2752,N_2787);
nand U5850 (N_5850,N_3812,N_3653);
nor U5851 (N_5851,N_2463,N_3023);
or U5852 (N_5852,N_3945,N_2883);
xnor U5853 (N_5853,N_3174,N_3934);
xnor U5854 (N_5854,N_3532,N_3203);
nand U5855 (N_5855,N_3236,N_3589);
nor U5856 (N_5856,N_3197,N_3504);
xor U5857 (N_5857,N_3934,N_3746);
nor U5858 (N_5858,N_3585,N_2617);
nand U5859 (N_5859,N_2638,N_3097);
nand U5860 (N_5860,N_2523,N_2520);
xnor U5861 (N_5861,N_2185,N_3692);
nor U5862 (N_5862,N_3248,N_2844);
and U5863 (N_5863,N_3594,N_3058);
nand U5864 (N_5864,N_2644,N_3767);
nand U5865 (N_5865,N_3099,N_2054);
xnor U5866 (N_5866,N_3979,N_3481);
and U5867 (N_5867,N_2017,N_3673);
or U5868 (N_5868,N_2384,N_3745);
xor U5869 (N_5869,N_3850,N_2135);
nor U5870 (N_5870,N_2513,N_3996);
and U5871 (N_5871,N_3168,N_2240);
nand U5872 (N_5872,N_3807,N_2840);
or U5873 (N_5873,N_3815,N_2451);
and U5874 (N_5874,N_3256,N_3609);
nand U5875 (N_5875,N_2419,N_3578);
nor U5876 (N_5876,N_3324,N_3315);
or U5877 (N_5877,N_3775,N_2534);
xnor U5878 (N_5878,N_2033,N_2535);
nor U5879 (N_5879,N_3923,N_3982);
or U5880 (N_5880,N_3132,N_3983);
nor U5881 (N_5881,N_3684,N_3182);
nand U5882 (N_5882,N_3782,N_3485);
or U5883 (N_5883,N_2390,N_3838);
nor U5884 (N_5884,N_2444,N_3635);
and U5885 (N_5885,N_2652,N_3333);
nor U5886 (N_5886,N_3638,N_3311);
and U5887 (N_5887,N_2487,N_2657);
and U5888 (N_5888,N_3620,N_2130);
nand U5889 (N_5889,N_3078,N_3168);
and U5890 (N_5890,N_2776,N_3439);
and U5891 (N_5891,N_2407,N_2627);
or U5892 (N_5892,N_3208,N_3196);
or U5893 (N_5893,N_3027,N_2309);
and U5894 (N_5894,N_2542,N_2350);
or U5895 (N_5895,N_2325,N_2888);
and U5896 (N_5896,N_2518,N_2250);
nand U5897 (N_5897,N_2896,N_3527);
and U5898 (N_5898,N_3302,N_2667);
nor U5899 (N_5899,N_2647,N_3844);
nor U5900 (N_5900,N_3761,N_2665);
and U5901 (N_5901,N_3366,N_3905);
xnor U5902 (N_5902,N_2964,N_3668);
nor U5903 (N_5903,N_2306,N_2237);
or U5904 (N_5904,N_3864,N_3079);
nor U5905 (N_5905,N_3437,N_3913);
nor U5906 (N_5906,N_2719,N_2396);
nor U5907 (N_5907,N_3313,N_3448);
and U5908 (N_5908,N_2396,N_2693);
nand U5909 (N_5909,N_3600,N_3096);
nand U5910 (N_5910,N_2216,N_2291);
nand U5911 (N_5911,N_3826,N_3208);
nand U5912 (N_5912,N_3796,N_3755);
or U5913 (N_5913,N_3131,N_2219);
xor U5914 (N_5914,N_2174,N_2440);
or U5915 (N_5915,N_2136,N_2008);
nand U5916 (N_5916,N_2656,N_2276);
nor U5917 (N_5917,N_3435,N_3416);
xnor U5918 (N_5918,N_2438,N_3801);
nor U5919 (N_5919,N_3035,N_3232);
nand U5920 (N_5920,N_3971,N_2727);
nor U5921 (N_5921,N_3005,N_2985);
or U5922 (N_5922,N_2100,N_2535);
or U5923 (N_5923,N_2854,N_3638);
nand U5924 (N_5924,N_3314,N_2127);
or U5925 (N_5925,N_2091,N_3652);
and U5926 (N_5926,N_2943,N_3667);
xor U5927 (N_5927,N_2051,N_3984);
or U5928 (N_5928,N_3730,N_2307);
xor U5929 (N_5929,N_3014,N_3168);
and U5930 (N_5930,N_3134,N_3156);
and U5931 (N_5931,N_2863,N_3710);
xnor U5932 (N_5932,N_2552,N_3339);
nand U5933 (N_5933,N_2633,N_3984);
or U5934 (N_5934,N_3734,N_3848);
and U5935 (N_5935,N_2801,N_3984);
nand U5936 (N_5936,N_2478,N_2715);
nand U5937 (N_5937,N_2559,N_2966);
nand U5938 (N_5938,N_3753,N_3804);
nor U5939 (N_5939,N_3820,N_2395);
and U5940 (N_5940,N_3739,N_2599);
nor U5941 (N_5941,N_3551,N_3971);
xnor U5942 (N_5942,N_3964,N_3502);
nor U5943 (N_5943,N_2606,N_2751);
xnor U5944 (N_5944,N_3177,N_2831);
and U5945 (N_5945,N_3551,N_3021);
or U5946 (N_5946,N_3261,N_2024);
and U5947 (N_5947,N_3025,N_2690);
xor U5948 (N_5948,N_3842,N_2584);
xnor U5949 (N_5949,N_3182,N_3674);
or U5950 (N_5950,N_3819,N_3180);
nor U5951 (N_5951,N_2046,N_3368);
xor U5952 (N_5952,N_3659,N_3875);
xor U5953 (N_5953,N_2869,N_2887);
nor U5954 (N_5954,N_3667,N_2881);
xnor U5955 (N_5955,N_3037,N_2613);
and U5956 (N_5956,N_3973,N_2957);
nor U5957 (N_5957,N_2531,N_2831);
nor U5958 (N_5958,N_3433,N_3276);
nor U5959 (N_5959,N_3750,N_2149);
nor U5960 (N_5960,N_2422,N_3173);
nand U5961 (N_5961,N_2633,N_2193);
and U5962 (N_5962,N_3432,N_2489);
nand U5963 (N_5963,N_2033,N_2512);
nor U5964 (N_5964,N_2013,N_3117);
nand U5965 (N_5965,N_2199,N_3653);
or U5966 (N_5966,N_2808,N_2194);
nand U5967 (N_5967,N_3599,N_3970);
or U5968 (N_5968,N_2486,N_3837);
xor U5969 (N_5969,N_3777,N_3740);
xor U5970 (N_5970,N_2972,N_2599);
and U5971 (N_5971,N_2778,N_3109);
and U5972 (N_5972,N_3330,N_2179);
nor U5973 (N_5973,N_2497,N_2590);
and U5974 (N_5974,N_3674,N_3243);
and U5975 (N_5975,N_2757,N_2035);
xnor U5976 (N_5976,N_2578,N_2736);
nand U5977 (N_5977,N_2014,N_2321);
or U5978 (N_5978,N_3299,N_2972);
or U5979 (N_5979,N_3474,N_2396);
or U5980 (N_5980,N_3785,N_2541);
and U5981 (N_5981,N_2620,N_3334);
and U5982 (N_5982,N_3139,N_2031);
nand U5983 (N_5983,N_3646,N_3006);
nand U5984 (N_5984,N_2829,N_3249);
nor U5985 (N_5985,N_3829,N_2026);
or U5986 (N_5986,N_3145,N_2130);
xnor U5987 (N_5987,N_2847,N_3430);
or U5988 (N_5988,N_2930,N_3576);
xnor U5989 (N_5989,N_3695,N_3497);
nand U5990 (N_5990,N_2776,N_2947);
and U5991 (N_5991,N_3016,N_3152);
nand U5992 (N_5992,N_3066,N_2910);
nor U5993 (N_5993,N_2384,N_2760);
nand U5994 (N_5994,N_2757,N_2660);
xor U5995 (N_5995,N_2477,N_2197);
xor U5996 (N_5996,N_3203,N_3019);
nand U5997 (N_5997,N_3170,N_3539);
xor U5998 (N_5998,N_2367,N_2025);
or U5999 (N_5999,N_2857,N_3223);
nand U6000 (N_6000,N_4753,N_5481);
xnor U6001 (N_6001,N_5974,N_5894);
or U6002 (N_6002,N_4744,N_5678);
xnor U6003 (N_6003,N_4961,N_5211);
xor U6004 (N_6004,N_5278,N_5970);
and U6005 (N_6005,N_5059,N_5545);
and U6006 (N_6006,N_5418,N_4708);
nand U6007 (N_6007,N_5298,N_4728);
and U6008 (N_6008,N_4691,N_5792);
and U6009 (N_6009,N_5800,N_5687);
nand U6010 (N_6010,N_5683,N_4944);
nand U6011 (N_6011,N_5198,N_5540);
xor U6012 (N_6012,N_4342,N_4401);
xnor U6013 (N_6013,N_4509,N_4531);
nor U6014 (N_6014,N_5812,N_4384);
xnor U6015 (N_6015,N_5062,N_4975);
or U6016 (N_6016,N_4520,N_5315);
or U6017 (N_6017,N_4832,N_5959);
and U6018 (N_6018,N_4328,N_4900);
and U6019 (N_6019,N_4184,N_5684);
xnor U6020 (N_6020,N_4624,N_4171);
nor U6021 (N_6021,N_5669,N_4415);
xor U6022 (N_6022,N_4776,N_5564);
and U6023 (N_6023,N_4994,N_4080);
nand U6024 (N_6024,N_5875,N_4262);
or U6025 (N_6025,N_4715,N_5563);
nand U6026 (N_6026,N_5578,N_4949);
and U6027 (N_6027,N_4867,N_5907);
xor U6028 (N_6028,N_4897,N_5229);
xnor U6029 (N_6029,N_5554,N_5317);
and U6030 (N_6030,N_5865,N_4990);
nand U6031 (N_6031,N_4942,N_4124);
or U6032 (N_6032,N_4878,N_5045);
nand U6033 (N_6033,N_4089,N_4306);
nor U6034 (N_6034,N_4781,N_5797);
nand U6035 (N_6035,N_4159,N_4847);
nand U6036 (N_6036,N_5848,N_5770);
nand U6037 (N_6037,N_4206,N_5453);
xnor U6038 (N_6038,N_5880,N_5326);
nand U6039 (N_6039,N_5719,N_5555);
xor U6040 (N_6040,N_5726,N_4120);
xnor U6041 (N_6041,N_5526,N_4037);
nand U6042 (N_6042,N_4570,N_5460);
and U6043 (N_6043,N_4511,N_5051);
nor U6044 (N_6044,N_4060,N_5333);
or U6045 (N_6045,N_5834,N_5471);
xnor U6046 (N_6046,N_4759,N_5001);
nand U6047 (N_6047,N_4811,N_4219);
and U6048 (N_6048,N_4739,N_5356);
nor U6049 (N_6049,N_5506,N_5842);
or U6050 (N_6050,N_5435,N_4272);
and U6051 (N_6051,N_5112,N_4191);
nor U6052 (N_6052,N_5942,N_5273);
nand U6053 (N_6053,N_5941,N_5514);
or U6054 (N_6054,N_4221,N_5632);
nand U6055 (N_6055,N_4676,N_4620);
and U6056 (N_6056,N_5360,N_5499);
or U6057 (N_6057,N_4018,N_4843);
nor U6058 (N_6058,N_4631,N_5204);
or U6059 (N_6059,N_5151,N_4924);
and U6060 (N_6060,N_5937,N_4253);
nor U6061 (N_6061,N_5302,N_5288);
and U6062 (N_6062,N_4889,N_5818);
nor U6063 (N_6063,N_5420,N_5348);
or U6064 (N_6064,N_5919,N_4472);
nor U6065 (N_6065,N_4464,N_4877);
xnor U6066 (N_6066,N_4748,N_5616);
nor U6067 (N_6067,N_5203,N_5598);
nor U6068 (N_6068,N_4855,N_4083);
and U6069 (N_6069,N_4114,N_5659);
and U6070 (N_6070,N_5399,N_5237);
nor U6071 (N_6071,N_4972,N_4983);
or U6072 (N_6072,N_4864,N_5864);
xor U6073 (N_6073,N_5331,N_4394);
and U6074 (N_6074,N_4167,N_5600);
nor U6075 (N_6075,N_4872,N_5218);
xnor U6076 (N_6076,N_5674,N_4455);
or U6077 (N_6077,N_4140,N_5162);
nand U6078 (N_6078,N_5649,N_4984);
nor U6079 (N_6079,N_5831,N_4977);
and U6080 (N_6080,N_5964,N_4073);
or U6081 (N_6081,N_4956,N_4786);
xor U6082 (N_6082,N_5790,N_4849);
xnor U6083 (N_6083,N_5508,N_5383);
xnor U6084 (N_6084,N_5989,N_5101);
nor U6085 (N_6085,N_5259,N_4906);
nor U6086 (N_6086,N_4603,N_4071);
xnor U6087 (N_6087,N_5558,N_4022);
xnor U6088 (N_6088,N_5718,N_5784);
and U6089 (N_6089,N_4696,N_5207);
nand U6090 (N_6090,N_4226,N_4376);
and U6091 (N_6091,N_5780,N_5365);
and U6092 (N_6092,N_4233,N_4638);
xor U6093 (N_6093,N_5705,N_4103);
nand U6094 (N_6094,N_4870,N_5260);
nand U6095 (N_6095,N_4264,N_5978);
nor U6096 (N_6096,N_5954,N_4907);
and U6097 (N_6097,N_4367,N_4178);
or U6098 (N_6098,N_5244,N_5591);
xnor U6099 (N_6099,N_4935,N_5149);
or U6100 (N_6100,N_4225,N_4590);
nand U6101 (N_6101,N_5484,N_5923);
nor U6102 (N_6102,N_5374,N_4452);
or U6103 (N_6103,N_4719,N_5282);
and U6104 (N_6104,N_4816,N_4417);
nand U6105 (N_6105,N_5932,N_4170);
nand U6106 (N_6106,N_5988,N_5291);
or U6107 (N_6107,N_5118,N_5078);
xnor U6108 (N_6108,N_5336,N_5058);
xnor U6109 (N_6109,N_5998,N_4668);
and U6110 (N_6110,N_5666,N_4543);
nor U6111 (N_6111,N_5549,N_5061);
nor U6112 (N_6112,N_4941,N_4657);
xnor U6113 (N_6113,N_4617,N_4831);
xnor U6114 (N_6114,N_5593,N_5290);
nand U6115 (N_6115,N_5945,N_4003);
or U6116 (N_6116,N_5936,N_5769);
and U6117 (N_6117,N_5929,N_5410);
nor U6118 (N_6118,N_4495,N_4914);
and U6119 (N_6119,N_5210,N_4197);
or U6120 (N_6120,N_4322,N_4350);
xor U6121 (N_6121,N_5829,N_4583);
and U6122 (N_6122,N_5807,N_5573);
nor U6123 (N_6123,N_5537,N_4788);
and U6124 (N_6124,N_4693,N_4218);
or U6125 (N_6125,N_4020,N_4228);
nand U6126 (N_6126,N_5429,N_4694);
nand U6127 (N_6127,N_5405,N_4319);
xor U6128 (N_6128,N_4345,N_5841);
and U6129 (N_6129,N_5178,N_4658);
xor U6130 (N_6130,N_5685,N_5092);
nor U6131 (N_6131,N_5142,N_4069);
xnor U6132 (N_6132,N_5156,N_5525);
nor U6133 (N_6133,N_4666,N_5147);
nand U6134 (N_6134,N_5909,N_4176);
nor U6135 (N_6135,N_5764,N_4490);
nand U6136 (N_6136,N_4485,N_5888);
xnor U6137 (N_6137,N_4614,N_5991);
or U6138 (N_6138,N_5010,N_4783);
xnor U6139 (N_6139,N_4584,N_4749);
and U6140 (N_6140,N_4048,N_5856);
nand U6141 (N_6141,N_5778,N_5454);
nor U6142 (N_6142,N_4789,N_4599);
and U6143 (N_6143,N_4287,N_5032);
nor U6144 (N_6144,N_5358,N_4669);
and U6145 (N_6145,N_5762,N_4834);
xor U6146 (N_6146,N_4899,N_5050);
xor U6147 (N_6147,N_4143,N_4454);
and U6148 (N_6148,N_4099,N_5971);
xnor U6149 (N_6149,N_4213,N_5712);
nor U6150 (N_6150,N_4436,N_4161);
and U6151 (N_6151,N_4241,N_5274);
nand U6152 (N_6152,N_5761,N_5128);
or U6153 (N_6153,N_5592,N_5706);
or U6154 (N_6154,N_4510,N_4526);
or U6155 (N_6155,N_4200,N_5212);
xor U6156 (N_6156,N_5100,N_5601);
and U6157 (N_6157,N_4553,N_5975);
or U6158 (N_6158,N_4360,N_4644);
or U6159 (N_6159,N_5375,N_5347);
or U6160 (N_6160,N_5148,N_5739);
or U6161 (N_6161,N_4090,N_4959);
nor U6162 (N_6162,N_4162,N_5235);
xor U6163 (N_6163,N_5895,N_4671);
nor U6164 (N_6164,N_4762,N_5673);
nand U6165 (N_6165,N_4466,N_4109);
xnor U6166 (N_6166,N_4461,N_4030);
and U6167 (N_6167,N_5993,N_5720);
nor U6168 (N_6168,N_5610,N_4371);
nor U6169 (N_6169,N_5625,N_4954);
nor U6170 (N_6170,N_4738,N_4398);
or U6171 (N_6171,N_4246,N_4192);
and U6172 (N_6172,N_4933,N_4175);
nand U6173 (N_6173,N_4016,N_5741);
nor U6174 (N_6174,N_5734,N_5900);
or U6175 (N_6175,N_4836,N_5028);
nor U6176 (N_6176,N_5703,N_4137);
and U6177 (N_6177,N_4767,N_5485);
or U6178 (N_6178,N_5376,N_4157);
or U6179 (N_6179,N_4416,N_4431);
xnor U6180 (N_6180,N_5055,N_4164);
xor U6181 (N_6181,N_5414,N_5258);
xor U6182 (N_6182,N_4641,N_5081);
nand U6183 (N_6183,N_4479,N_5921);
nor U6184 (N_6184,N_4174,N_4546);
xnor U6185 (N_6185,N_5751,N_4707);
and U6186 (N_6186,N_4790,N_5738);
nand U6187 (N_6187,N_4547,N_5876);
and U6188 (N_6188,N_4411,N_5247);
and U6189 (N_6189,N_4727,N_5427);
or U6190 (N_6190,N_5576,N_4600);
nand U6191 (N_6191,N_5199,N_5392);
xnor U6192 (N_6192,N_5049,N_4647);
nor U6193 (N_6193,N_5456,N_5323);
or U6194 (N_6194,N_5773,N_4275);
nand U6195 (N_6195,N_5469,N_5445);
and U6196 (N_6196,N_4078,N_4395);
nor U6197 (N_6197,N_4268,N_4009);
or U6198 (N_6198,N_4427,N_4247);
xor U6199 (N_6199,N_5835,N_5458);
or U6200 (N_6200,N_4375,N_4697);
xor U6201 (N_6201,N_4356,N_5440);
nor U6202 (N_6202,N_5353,N_4895);
and U6203 (N_6203,N_4913,N_5691);
nor U6204 (N_6204,N_4243,N_4751);
nand U6205 (N_6205,N_5385,N_4709);
xor U6206 (N_6206,N_5587,N_4894);
or U6207 (N_6207,N_4640,N_5479);
or U6208 (N_6208,N_4491,N_4134);
nor U6209 (N_6209,N_4716,N_5184);
or U6210 (N_6210,N_5823,N_4541);
and U6211 (N_6211,N_4361,N_4551);
or U6212 (N_6212,N_4566,N_5815);
xnor U6213 (N_6213,N_4985,N_5568);
nor U6214 (N_6214,N_5103,N_4252);
nand U6215 (N_6215,N_5188,N_4166);
xor U6216 (N_6216,N_5953,N_4880);
nand U6217 (N_6217,N_5475,N_4105);
nor U6218 (N_6218,N_5722,N_5949);
or U6219 (N_6219,N_4629,N_4679);
nand U6220 (N_6220,N_5567,N_4632);
xor U6221 (N_6221,N_4592,N_5642);
and U6222 (N_6222,N_4766,N_5527);
xnor U6223 (N_6223,N_4795,N_5735);
nor U6224 (N_6224,N_4468,N_4742);
xor U6225 (N_6225,N_4554,N_4172);
and U6226 (N_6226,N_4712,N_5871);
nor U6227 (N_6227,N_5717,N_5849);
xor U6228 (N_6228,N_5168,N_4634);
nand U6229 (N_6229,N_5551,N_4049);
or U6230 (N_6230,N_5132,N_5619);
and U6231 (N_6231,N_4093,N_5867);
nor U6232 (N_6232,N_4156,N_5655);
and U6233 (N_6233,N_5373,N_5544);
xnor U6234 (N_6234,N_5756,N_5585);
and U6235 (N_6235,N_4958,N_5808);
and U6236 (N_6236,N_4672,N_5745);
or U6237 (N_6237,N_4119,N_4380);
and U6238 (N_6238,N_5434,N_4733);
or U6239 (N_6239,N_4571,N_5082);
xnor U6240 (N_6240,N_4095,N_5711);
nor U6241 (N_6241,N_4014,N_4024);
nand U6242 (N_6242,N_4273,N_4098);
nor U6243 (N_6243,N_4806,N_4128);
xnor U6244 (N_6244,N_4338,N_5119);
or U6245 (N_6245,N_5847,N_5425);
xor U6246 (N_6246,N_5490,N_5093);
and U6247 (N_6247,N_4248,N_4195);
nor U6248 (N_6248,N_5981,N_4819);
nor U6249 (N_6249,N_5825,N_4965);
xnor U6250 (N_6250,N_5589,N_4800);
nand U6251 (N_6251,N_4758,N_4550);
nor U6252 (N_6252,N_4528,N_4936);
and U6253 (N_6253,N_4298,N_4011);
xor U6254 (N_6254,N_5289,N_4276);
xor U6255 (N_6255,N_4177,N_5438);
nor U6256 (N_6256,N_4928,N_5505);
xnor U6257 (N_6257,N_4269,N_5268);
xnor U6258 (N_6258,N_4987,N_5166);
xor U6259 (N_6259,N_4721,N_5897);
nor U6260 (N_6260,N_5636,N_5368);
nor U6261 (N_6261,N_4106,N_4854);
and U6262 (N_6262,N_5521,N_5417);
nand U6263 (N_6263,N_5760,N_5217);
nor U6264 (N_6264,N_4068,N_4734);
and U6265 (N_6265,N_5707,N_4862);
and U6266 (N_6266,N_5401,N_4756);
nand U6267 (N_6267,N_4187,N_5874);
nor U6268 (N_6268,N_4331,N_4459);
or U6269 (N_6269,N_5306,N_5861);
or U6270 (N_6270,N_5209,N_4940);
and U6271 (N_6271,N_4997,N_5415);
or U6272 (N_6272,N_5520,N_4821);
or U6273 (N_6273,N_5457,N_4136);
nand U6274 (N_6274,N_4008,N_4007);
nand U6275 (N_6275,N_5304,N_5744);
nand U6276 (N_6276,N_5623,N_5901);
nand U6277 (N_6277,N_4702,N_5968);
xor U6278 (N_6278,N_4879,N_4916);
xor U6279 (N_6279,N_4768,N_5114);
and U6280 (N_6280,N_5023,N_4835);
and U6281 (N_6281,N_5271,N_4652);
xnor U6282 (N_6282,N_4239,N_4004);
nor U6283 (N_6283,N_4317,N_4056);
xor U6284 (N_6284,N_5191,N_4462);
xnor U6285 (N_6285,N_4092,N_5432);
nand U6286 (N_6286,N_5795,N_4608);
nand U6287 (N_6287,N_5441,N_4607);
xnor U6288 (N_6288,N_4683,N_4122);
or U6289 (N_6289,N_5608,N_5657);
and U6290 (N_6290,N_4237,N_5651);
or U6291 (N_6291,N_4160,N_5590);
and U6292 (N_6292,N_4355,N_4998);
xor U6293 (N_6293,N_4978,N_5817);
or U6294 (N_6294,N_5254,N_5701);
nand U6295 (N_6295,N_4082,N_5556);
xnor U6296 (N_6296,N_5866,N_4075);
nand U6297 (N_6297,N_4434,N_4278);
nand U6298 (N_6298,N_4882,N_5472);
and U6299 (N_6299,N_5339,N_5528);
nor U6300 (N_6300,N_4812,N_4687);
or U6301 (N_6301,N_5240,N_5287);
nor U6302 (N_6302,N_4070,N_4424);
or U6303 (N_6303,N_4163,N_4285);
nand U6304 (N_6304,N_5295,N_5190);
and U6305 (N_6305,N_4369,N_5223);
or U6306 (N_6306,N_5488,N_5077);
or U6307 (N_6307,N_5020,N_4094);
xnor U6308 (N_6308,N_4044,N_5197);
xor U6309 (N_6309,N_4667,N_5292);
nand U6310 (N_6310,N_5785,N_5136);
nor U6311 (N_6311,N_5412,N_5068);
nand U6312 (N_6312,N_4148,N_5477);
nor U6313 (N_6313,N_4792,N_5272);
nor U6314 (N_6314,N_4690,N_4304);
and U6315 (N_6315,N_4204,N_5962);
and U6316 (N_6316,N_5776,N_5017);
and U6317 (N_6317,N_5213,N_4893);
and U6318 (N_6318,N_4433,N_5022);
and U6319 (N_6319,N_4582,N_4596);
and U6320 (N_6320,N_5318,N_5882);
nor U6321 (N_6321,N_4006,N_4587);
nand U6322 (N_6322,N_4651,N_5896);
nor U6323 (N_6323,N_4308,N_4976);
or U6324 (N_6324,N_4934,N_5566);
nor U6325 (N_6325,N_5480,N_5535);
and U6326 (N_6326,N_5952,N_5884);
or U6327 (N_6327,N_4445,N_4868);
or U6328 (N_6328,N_5447,N_4488);
or U6329 (N_6329,N_4005,N_4680);
nor U6330 (N_6330,N_5987,N_5519);
xnor U6331 (N_6331,N_4519,N_5653);
nor U6332 (N_6332,N_4723,N_5473);
nor U6333 (N_6333,N_5428,N_4327);
or U6334 (N_6334,N_4798,N_5543);
nor U6335 (N_6335,N_5225,N_5003);
nor U6336 (N_6336,N_5740,N_5546);
or U6337 (N_6337,N_4027,N_5413);
nand U6338 (N_6338,N_4257,N_5965);
nor U6339 (N_6339,N_4557,N_5538);
nand U6340 (N_6340,N_5997,N_5056);
nor U6341 (N_6341,N_5513,N_5227);
or U6342 (N_6342,N_4747,N_4025);
and U6343 (N_6343,N_5926,N_4904);
nor U6344 (N_6344,N_4419,N_5046);
nand U6345 (N_6345,N_5140,N_4100);
nand U6346 (N_6346,N_5437,N_4310);
and U6347 (N_6347,N_5245,N_5973);
or U6348 (N_6348,N_4621,N_5588);
and U6349 (N_6349,N_5097,N_5325);
or U6350 (N_6350,N_5179,N_5782);
and U6351 (N_6351,N_4903,N_5877);
or U6352 (N_6352,N_5214,N_4223);
or U6353 (N_6353,N_5363,N_5943);
nor U6354 (N_6354,N_5367,N_5221);
and U6355 (N_6355,N_5379,N_5886);
and U6356 (N_6356,N_5448,N_5562);
xnor U6357 (N_6357,N_5135,N_4351);
xor U6358 (N_6358,N_5332,N_4947);
nand U6359 (N_6359,N_5487,N_5710);
nor U6360 (N_6360,N_4481,N_5904);
nor U6361 (N_6361,N_4493,N_4293);
or U6362 (N_6362,N_5638,N_4289);
nand U6363 (N_6363,N_5595,N_4780);
nand U6364 (N_6364,N_5123,N_4274);
or U6365 (N_6365,N_4181,N_4923);
nand U6366 (N_6366,N_4840,N_5681);
xor U6367 (N_6367,N_4421,N_4589);
nand U6368 (N_6368,N_4530,N_4898);
nand U6369 (N_6369,N_5580,N_4067);
nor U6370 (N_6370,N_5422,N_4318);
nor U6371 (N_6371,N_4457,N_4609);
nand U6372 (N_6372,N_4453,N_5646);
xor U6373 (N_6373,N_5950,N_4850);
and U6374 (N_6374,N_4785,N_5899);
or U6375 (N_6375,N_5430,N_5648);
and U6376 (N_6376,N_5881,N_4912);
and U6377 (N_6377,N_4333,N_4591);
nor U6378 (N_6378,N_5976,N_4061);
xnor U6379 (N_6379,N_4623,N_5352);
nand U6380 (N_6380,N_5724,N_4532);
and U6381 (N_6381,N_4238,N_4704);
xor U6382 (N_6382,N_5073,N_5700);
nor U6383 (N_6383,N_4188,N_4505);
nor U6384 (N_6384,N_5033,N_5215);
nor U6385 (N_6385,N_4874,N_5967);
nand U6386 (N_6386,N_4168,N_5624);
nand U6387 (N_6387,N_5721,N_4929);
xnor U6388 (N_6388,N_4833,N_5277);
nor U6389 (N_6389,N_4803,N_4993);
nor U6390 (N_6390,N_5181,N_5803);
xor U6391 (N_6391,N_5249,N_5862);
or U6392 (N_6392,N_4736,N_4130);
and U6393 (N_6393,N_4258,N_5164);
nor U6394 (N_6394,N_5502,N_5079);
or U6395 (N_6395,N_5671,N_4699);
nor U6396 (N_6396,N_4866,N_4569);
xor U6397 (N_6397,N_4203,N_4981);
or U6398 (N_6398,N_5708,N_4724);
or U6399 (N_6399,N_4408,N_5024);
xnor U6400 (N_6400,N_4277,N_5411);
nand U6401 (N_6401,N_5736,N_4391);
nor U6402 (N_6402,N_4000,N_4209);
and U6403 (N_6403,N_4649,N_4718);
and U6404 (N_6404,N_5634,N_5228);
or U6405 (N_6405,N_4227,N_4079);
and U6406 (N_6406,N_4881,N_5388);
nand U6407 (N_6407,N_5660,N_4922);
or U6408 (N_6408,N_5765,N_4999);
nand U6409 (N_6409,N_5006,N_5827);
nor U6410 (N_6410,N_4901,N_5534);
xor U6411 (N_6411,N_4217,N_5618);
and U6412 (N_6412,N_5391,N_4052);
xor U6413 (N_6413,N_5637,N_4829);
xnor U6414 (N_6414,N_4905,N_4026);
nor U6415 (N_6415,N_4556,N_5222);
and U6416 (N_6416,N_4324,N_4146);
or U6417 (N_6417,N_4741,N_4635);
or U6418 (N_6418,N_4793,N_4291);
or U6419 (N_6419,N_4957,N_4501);
nor U6420 (N_6420,N_5938,N_5493);
or U6421 (N_6421,N_4085,N_4522);
or U6422 (N_6422,N_5074,N_4810);
xnor U6423 (N_6423,N_4336,N_5497);
nand U6424 (N_6424,N_5672,N_4368);
or U6425 (N_6425,N_5072,N_5934);
and U6426 (N_6426,N_4787,N_5531);
and U6427 (N_6427,N_5643,N_4397);
xnor U6428 (N_6428,N_5947,N_4117);
xnor U6429 (N_6429,N_4193,N_4364);
and U6430 (N_6430,N_5366,N_4982);
nor U6431 (N_6431,N_4299,N_4951);
nor U6432 (N_6432,N_5029,N_5335);
nor U6433 (N_6433,N_5912,N_5138);
xor U6434 (N_6434,N_4626,N_4107);
nand U6435 (N_6435,N_5844,N_5878);
xor U6436 (N_6436,N_5163,N_4077);
and U6437 (N_6437,N_5308,N_5316);
or U6438 (N_6438,N_5639,N_5057);
nor U6439 (N_6439,N_5983,N_4469);
and U6440 (N_6440,N_5791,N_4886);
xor U6441 (N_6441,N_5731,N_4875);
xnor U6442 (N_6442,N_5826,N_4654);
or U6443 (N_6443,N_5115,N_4633);
or U6444 (N_6444,N_4055,N_5483);
nor U6445 (N_6445,N_5085,N_5768);
nand U6446 (N_6446,N_5297,N_4910);
nand U6447 (N_6447,N_5898,N_5153);
nor U6448 (N_6448,N_5071,N_5913);
and U6449 (N_6449,N_5944,N_4432);
or U6450 (N_6450,N_4118,N_4320);
or U6451 (N_6451,N_5130,N_5570);
xnor U6452 (N_6452,N_5005,N_5014);
nand U6453 (N_6453,N_5381,N_5522);
nor U6454 (N_6454,N_4363,N_5796);
nor U6455 (N_6455,N_5609,N_4205);
xnor U6456 (N_6456,N_4021,N_5433);
nor U6457 (N_6457,N_4678,N_5110);
xor U6458 (N_6458,N_5402,N_5195);
nand U6459 (N_6459,N_4474,N_4670);
or U6460 (N_6460,N_4516,N_5129);
or U6461 (N_6461,N_4013,N_4636);
xnor U6462 (N_6462,N_5183,N_4774);
xnor U6463 (N_6463,N_4279,N_4396);
nor U6464 (N_6464,N_5781,N_5786);
nand U6465 (N_6465,N_4244,N_4815);
nand U6466 (N_6466,N_4038,N_5507);
nor U6467 (N_6467,N_5094,N_4820);
and U6468 (N_6468,N_4955,N_4404);
xnor U6469 (N_6469,N_5342,N_5202);
xnor U6470 (N_6470,N_4964,N_5654);
nor U6471 (N_6471,N_5126,N_5980);
and U6472 (N_6472,N_5533,N_5927);
nor U6473 (N_6473,N_4471,N_5467);
and U6474 (N_6474,N_5969,N_4032);
or U6475 (N_6475,N_5424,N_5495);
or U6476 (N_6476,N_4435,N_5357);
or U6477 (N_6477,N_4525,N_5696);
or U6478 (N_6478,N_4418,N_5173);
and U6479 (N_6479,N_4451,N_4845);
nor U6480 (N_6480,N_5180,N_5139);
nand U6481 (N_6481,N_4659,N_5852);
nand U6482 (N_6482,N_5378,N_5713);
and U6483 (N_6483,N_5963,N_5037);
nor U6484 (N_6484,N_5594,N_5892);
or U6485 (N_6485,N_5120,N_4151);
or U6486 (N_6486,N_5958,N_4414);
nand U6487 (N_6487,N_4805,N_4830);
xor U6488 (N_6488,N_4732,N_5423);
xnor U6489 (N_6489,N_4131,N_5990);
or U6490 (N_6490,N_5501,N_4487);
or U6491 (N_6491,N_4033,N_4627);
and U6492 (N_6492,N_4392,N_4648);
nor U6493 (N_6493,N_4270,N_5075);
xnor U6494 (N_6494,N_4797,N_4284);
or U6495 (N_6495,N_5930,N_5801);
nor U6496 (N_6496,N_5048,N_4051);
xnor U6497 (N_6497,N_5270,N_4017);
or U6498 (N_6498,N_4735,N_4529);
nor U6499 (N_6499,N_4945,N_5830);
nand U6500 (N_6500,N_4559,N_4325);
xnor U6501 (N_6501,N_4564,N_5992);
nor U6502 (N_6502,N_4212,N_4307);
and U6503 (N_6503,N_4498,N_4602);
or U6504 (N_6504,N_4823,N_5088);
nand U6505 (N_6505,N_5515,N_5668);
nand U6506 (N_6506,N_4572,N_4674);
nand U6507 (N_6507,N_5906,N_4731);
nand U6508 (N_6508,N_4154,N_4261);
and U6509 (N_6509,N_4925,N_5098);
xnor U6510 (N_6510,N_5577,N_5102);
nor U6511 (N_6511,N_4066,N_4001);
nand U6512 (N_6512,N_5109,N_5465);
or U6513 (N_6513,N_4851,N_4996);
nor U6514 (N_6514,N_5868,N_5879);
and U6515 (N_6515,N_5474,N_4483);
or U6516 (N_6516,N_4286,N_4235);
nor U6517 (N_6517,N_5994,N_5084);
and U6518 (N_6518,N_4379,N_4655);
xor U6519 (N_6519,N_5676,N_5283);
and U6520 (N_6520,N_4852,N_4086);
xnor U6521 (N_6521,N_5285,N_4777);
xnor U6522 (N_6522,N_4442,N_5305);
or U6523 (N_6523,N_4339,N_5565);
or U6524 (N_6524,N_5746,N_5840);
xnor U6525 (N_6525,N_4220,N_4939);
xnor U6526 (N_6526,N_5063,N_4062);
and U6527 (N_6527,N_5920,N_4214);
nand U6528 (N_6528,N_4950,N_4064);
nand U6529 (N_6529,N_4967,N_4365);
xnor U6530 (N_6530,N_4297,N_4230);
nand U6531 (N_6531,N_4980,N_4344);
and U6532 (N_6532,N_5652,N_5859);
or U6533 (N_6533,N_4927,N_5394);
or U6534 (N_6534,N_5960,N_5451);
or U6535 (N_6535,N_5903,N_4865);
xor U6536 (N_6536,N_4673,N_5337);
nor U6537 (N_6537,N_4703,N_5171);
nor U6538 (N_6538,N_5013,N_5733);
xor U6539 (N_6539,N_5887,N_4335);
xnor U6540 (N_6540,N_5915,N_5758);
and U6541 (N_6541,N_4545,N_5052);
and U6542 (N_6542,N_5154,N_4377);
nor U6543 (N_6543,N_4314,N_5299);
xor U6544 (N_6544,N_4822,N_5832);
nor U6545 (N_6545,N_5729,N_4628);
nor U6546 (N_6546,N_4249,N_4698);
xor U6547 (N_6547,N_5890,N_4639);
nor U6548 (N_6548,N_4296,N_4358);
nor U6549 (N_6549,N_5523,N_4720);
or U6550 (N_6550,N_4475,N_4773);
nand U6551 (N_6551,N_4450,N_5267);
nand U6552 (N_6552,N_5313,N_4650);
nand U6553 (N_6553,N_4102,N_4222);
nand U6554 (N_6554,N_4372,N_5647);
or U6555 (N_6555,N_5397,N_5820);
xor U6556 (N_6556,N_5843,N_4588);
and U6557 (N_6557,N_4441,N_5819);
or U6558 (N_6558,N_4685,N_4825);
and U6559 (N_6559,N_5341,N_5170);
and U6560 (N_6560,N_4381,N_4323);
xor U6561 (N_6561,N_5253,N_4725);
xor U6562 (N_6562,N_4745,N_5182);
nor U6563 (N_6563,N_5622,N_4084);
nor U6564 (N_6564,N_5787,N_4841);
xnor U6565 (N_6565,N_5091,N_4711);
nor U6566 (N_6566,N_4514,N_5806);
xnor U6567 (N_6567,N_4574,N_4521);
and U6568 (N_6568,N_5737,N_4710);
and U6569 (N_6569,N_4796,N_5759);
and U6570 (N_6570,N_5265,N_5813);
nor U6571 (N_6571,N_4871,N_4207);
and U6572 (N_6572,N_5455,N_5349);
xnor U6573 (N_6573,N_5070,N_4625);
xor U6574 (N_6574,N_5836,N_5105);
xor U6575 (N_6575,N_5799,N_5606);
xor U6576 (N_6576,N_4653,N_5095);
xor U6577 (N_6577,N_5011,N_5851);
xnor U6578 (N_6578,N_4858,N_4771);
or U6579 (N_6579,N_5810,N_4046);
xnor U6580 (N_6580,N_5870,N_4410);
or U6581 (N_6581,N_4458,N_4036);
nor U6582 (N_6582,N_5688,N_5951);
nand U6583 (N_6583,N_5134,N_5498);
or U6584 (N_6584,N_4232,N_4429);
or U6585 (N_6585,N_5236,N_4357);
or U6586 (N_6586,N_5775,N_4240);
nand U6587 (N_6587,N_4029,N_5539);
and U6588 (N_6588,N_4266,N_5504);
nor U6589 (N_6589,N_5146,N_4309);
or U6590 (N_6590,N_4091,N_5106);
or U6591 (N_6591,N_4448,N_4689);
xor U6592 (N_6592,N_4210,N_5917);
and U6593 (N_6593,N_5409,N_5152);
nor U6594 (N_6594,N_5065,N_5312);
nand U6595 (N_6595,N_5404,N_5319);
or U6596 (N_6596,N_5257,N_4932);
and U6597 (N_6597,N_4594,N_5869);
and U6598 (N_6598,N_5863,N_5044);
and U6599 (N_6599,N_5697,N_5416);
nor U6600 (N_6600,N_5155,N_4552);
nand U6601 (N_6601,N_4963,N_5518);
xor U6602 (N_6602,N_4549,N_4202);
or U6603 (N_6603,N_4568,N_4754);
nor U6604 (N_6604,N_5234,N_5066);
and U6605 (N_6605,N_4743,N_4115);
nor U6606 (N_6606,N_5747,N_5444);
nand U6607 (N_6607,N_4775,N_4348);
nor U6608 (N_6608,N_5407,N_4502);
or U6609 (N_6609,N_4383,N_5030);
nor U6610 (N_6610,N_4111,N_4042);
nand U6611 (N_6611,N_4544,N_5113);
nor U6612 (N_6612,N_4260,N_4534);
nand U6613 (N_6613,N_5275,N_5346);
xor U6614 (N_6614,N_5661,N_5814);
and U6615 (N_6615,N_4489,N_4681);
nand U6616 (N_6616,N_5370,N_5732);
nor U6617 (N_6617,N_4863,N_5431);
and U6618 (N_6618,N_5226,N_4058);
xnor U6619 (N_6619,N_4467,N_4180);
or U6620 (N_6620,N_5276,N_4536);
nand U6621 (N_6621,N_4141,N_5611);
xnor U6622 (N_6622,N_4612,N_5167);
nor U6623 (N_6623,N_4619,N_4799);
xnor U6624 (N_6624,N_5334,N_5255);
nor U6625 (N_6625,N_4598,N_5984);
or U6626 (N_6626,N_5955,N_5575);
nand U6627 (N_6627,N_4560,N_5557);
nand U6628 (N_6628,N_5583,N_5193);
xnor U6629 (N_6629,N_5007,N_4665);
nor U6630 (N_6630,N_5667,N_5794);
and U6631 (N_6631,N_4326,N_4808);
nand U6632 (N_6632,N_5536,N_5386);
nand U6633 (N_6633,N_4354,N_5384);
and U6634 (N_6634,N_5344,N_5828);
nor U6635 (N_6635,N_4848,N_4034);
and U6636 (N_6636,N_4595,N_4028);
and U6637 (N_6637,N_4824,N_4885);
and U6638 (N_6638,N_5928,N_5406);
and U6639 (N_6639,N_4373,N_4890);
and U6640 (N_6640,N_5220,N_5086);
or U6641 (N_6641,N_4705,N_5311);
nor U6642 (N_6642,N_4856,N_4884);
and U6643 (N_6643,N_5749,N_5280);
nand U6644 (N_6644,N_4616,N_4353);
nand U6645 (N_6645,N_5727,N_5470);
or U6646 (N_6646,N_5607,N_4891);
nand U6647 (N_6647,N_5584,N_5121);
xor U6648 (N_6648,N_5946,N_5925);
nor U6649 (N_6649,N_5145,N_5626);
nor U6650 (N_6650,N_5995,N_4087);
or U6651 (N_6651,N_5329,N_5940);
nor U6652 (N_6652,N_4892,N_4460);
and U6653 (N_6653,N_4992,N_5256);
nor U6654 (N_6654,N_5169,N_4902);
xor U6655 (N_6655,N_4507,N_4446);
xor U6656 (N_6656,N_4422,N_5716);
or U6657 (N_6657,N_5205,N_4818);
and U6658 (N_6658,N_5599,N_5060);
xor U6659 (N_6659,N_4801,N_5266);
and U6660 (N_6660,N_4578,N_5459);
nand U6661 (N_6661,N_5579,N_5125);
nor U6662 (N_6662,N_5403,N_4765);
or U6663 (N_6663,N_5016,N_5857);
and U6664 (N_6664,N_5400,N_4015);
or U6665 (N_6665,N_4402,N_4147);
nor U6666 (N_6666,N_5380,N_4953);
or U6667 (N_6667,N_4919,N_5620);
and U6668 (N_6668,N_5748,N_5779);
nor U6669 (N_6669,N_5038,N_5574);
or U6670 (N_6670,N_4135,N_4412);
xor U6671 (N_6671,N_5977,N_4423);
nand U6672 (N_6672,N_4646,N_4769);
and U6673 (N_6673,N_5723,N_5393);
nand U6674 (N_6674,N_4389,N_4280);
or U6675 (N_6675,N_4837,N_5702);
or U6676 (N_6676,N_5369,N_5160);
or U6677 (N_6677,N_4125,N_4970);
and U6678 (N_6678,N_5511,N_5439);
xor U6679 (N_6679,N_5241,N_5054);
xor U6680 (N_6680,N_4784,N_4150);
and U6681 (N_6681,N_4562,N_5628);
and U6682 (N_6682,N_5371,N_5450);
nor U6683 (N_6683,N_5133,N_4908);
xor U6684 (N_6684,N_5027,N_5644);
or U6685 (N_6685,N_4610,N_5468);
or U6686 (N_6686,N_5948,N_4449);
and U6687 (N_6687,N_5850,N_5548);
nor U6688 (N_6688,N_4340,N_4618);
xor U6689 (N_6689,N_4791,N_4035);
nand U6690 (N_6690,N_4508,N_4012);
nand U6691 (N_6691,N_5679,N_4597);
nand U6692 (N_6692,N_5924,N_4142);
xor U6693 (N_6693,N_4660,N_5206);
nor U6694 (N_6694,N_5122,N_4645);
nor U6695 (N_6695,N_5986,N_5462);
nand U6696 (N_6696,N_5036,N_4039);
xor U6697 (N_6697,N_4265,N_5665);
or U6698 (N_6698,N_5552,N_5656);
or U6699 (N_6699,N_5922,N_4031);
xor U6700 (N_6700,N_5284,N_4752);
xor U6701 (N_6701,N_4523,N_5251);
or U6702 (N_6702,N_5489,N_5503);
nor U6703 (N_6703,N_4701,N_5390);
and U6704 (N_6704,N_5269,N_5144);
nor U6705 (N_6705,N_5127,N_4763);
xor U6706 (N_6706,N_4931,N_4229);
nor U6707 (N_6707,N_4138,N_4496);
nand U6708 (N_6708,N_4688,N_5242);
and U6709 (N_6709,N_5043,N_5883);
and U6710 (N_6710,N_4730,N_5307);
and U6711 (N_6711,N_4316,N_5187);
and U6712 (N_6712,N_5961,N_5314);
and U6713 (N_6713,N_5561,N_5177);
xnor U6714 (N_6714,N_4047,N_4382);
nor U6715 (N_6715,N_5686,N_4662);
nor U6716 (N_6716,N_4330,N_5026);
and U6717 (N_6717,N_5008,N_4132);
nor U6718 (N_6718,N_4456,N_5798);
and U6719 (N_6719,N_4236,N_4183);
and U6720 (N_6720,N_5777,N_5766);
or U6721 (N_6721,N_4642,N_4189);
nand U6722 (N_6722,N_4245,N_4362);
xnor U6723 (N_6723,N_4503,N_4430);
xor U6724 (N_6724,N_5783,N_5124);
or U6725 (N_6725,N_4746,N_5640);
nor U6726 (N_6726,N_5999,N_5693);
or U6727 (N_6727,N_5893,N_4860);
nor U6728 (N_6728,N_5757,N_4492);
nor U6729 (N_6729,N_5377,N_5463);
xor U6730 (N_6730,N_5571,N_5099);
nor U6731 (N_6731,N_4973,N_4387);
nor U6732 (N_6732,N_5042,N_4722);
nor U6733 (N_6733,N_4231,N_5621);
or U6734 (N_6734,N_4185,N_5449);
nor U6735 (N_6735,N_4542,N_4760);
nor U6736 (N_6736,N_5902,N_5617);
or U6737 (N_6737,N_5677,N_4772);
and U6738 (N_6738,N_5243,N_5279);
nor U6739 (N_6739,N_5572,N_5931);
or U6740 (N_6740,N_5252,N_5547);
xnor U6741 (N_6741,N_5224,N_4186);
nand U6742 (N_6742,N_4321,N_5704);
xnor U6743 (N_6743,N_4989,N_4349);
and U6744 (N_6744,N_4282,N_5309);
xor U6745 (N_6745,N_4540,N_5004);
nor U6746 (N_6746,N_5532,N_4347);
or U6747 (N_6747,N_5117,N_5755);
and U6748 (N_6748,N_4169,N_4063);
and U6749 (N_6749,N_4606,N_5345);
or U6750 (N_6750,N_5492,N_5550);
nor U6751 (N_6751,N_4312,N_4630);
and U6752 (N_6752,N_5631,N_5263);
or U6753 (N_6753,N_4440,N_5569);
nand U6754 (N_6754,N_5966,N_4294);
nor U6755 (N_6755,N_4986,N_5104);
and U6756 (N_6756,N_5730,N_4952);
or U6757 (N_6757,N_4804,N_5320);
xnor U6758 (N_6758,N_5194,N_4555);
xor U6759 (N_6759,N_4473,N_5087);
and U6760 (N_6760,N_4613,N_5192);
nand U6761 (N_6761,N_5452,N_5630);
nor U6762 (N_6762,N_4611,N_4991);
nand U6763 (N_6763,N_4465,N_5137);
nor U6764 (N_6764,N_4390,N_4129);
xnor U6765 (N_6765,N_5559,N_4827);
and U6766 (N_6766,N_5090,N_5159);
and U6767 (N_6767,N_5421,N_4943);
xor U6768 (N_6768,N_5031,N_5286);
and U6769 (N_6769,N_4828,N_4437);
or U6770 (N_6770,N_4575,N_4301);
xor U6771 (N_6771,N_4938,N_5633);
nor U6772 (N_6772,N_4915,N_4909);
nor U6773 (N_6773,N_4764,N_5699);
nor U6774 (N_6774,N_4968,N_4300);
and U6775 (N_6775,N_4517,N_4057);
nor U6776 (N_6776,N_4267,N_4663);
or U6777 (N_6777,N_4182,N_5083);
nand U6778 (N_6778,N_4332,N_5586);
xnor U6779 (N_6779,N_5694,N_5581);
nand U6780 (N_6780,N_5839,N_4370);
nand U6781 (N_6781,N_4873,N_5131);
nand U6782 (N_6782,N_4778,N_5597);
and U6783 (N_6783,N_5530,N_5047);
xnor U6784 (N_6784,N_4443,N_5854);
nor U6785 (N_6785,N_5039,N_5709);
and U6786 (N_6786,N_5246,N_4406);
or U6787 (N_6787,N_4428,N_5264);
or U6788 (N_6788,N_5714,N_5443);
nor U6789 (N_6789,N_5476,N_4196);
nand U6790 (N_6790,N_4315,N_5396);
and U6791 (N_6791,N_5604,N_4040);
or U6792 (N_6792,N_4615,N_4604);
or U6793 (N_6793,N_4158,N_4144);
or U6794 (N_6794,N_4023,N_5692);
and U6795 (N_6795,N_5015,N_5294);
or U6796 (N_6796,N_4930,N_4208);
nor U6797 (N_6797,N_5116,N_5500);
nor U6798 (N_6798,N_4378,N_5753);
nor U6799 (N_6799,N_5466,N_4499);
and U6800 (N_6800,N_4802,N_5324);
nor U6801 (N_6801,N_4385,N_4426);
nor U6802 (N_6802,N_5069,N_4779);
nor U6803 (N_6803,N_4576,N_5804);
nand U6804 (N_6804,N_5025,N_4692);
nor U6805 (N_6805,N_4656,N_4911);
nand U6806 (N_6806,N_5629,N_4484);
nor U6807 (N_6807,N_5635,N_5918);
nand U6808 (N_6808,N_5664,N_4838);
or U6809 (N_6809,N_5860,N_4292);
nand U6810 (N_6810,N_5248,N_4110);
xnor U6811 (N_6811,N_5165,N_5605);
nor U6812 (N_6812,N_5690,N_4149);
or U6813 (N_6813,N_4346,N_4123);
xor U6814 (N_6814,N_5012,N_4341);
nand U6815 (N_6815,N_4179,N_5529);
or U6816 (N_6816,N_5239,N_5771);
or U6817 (N_6817,N_4366,N_5833);
nor U6818 (N_6818,N_4420,N_5189);
nor U6819 (N_6819,N_4190,N_5512);
nor U6820 (N_6820,N_5000,N_5645);
or U6821 (N_6821,N_5542,N_5281);
nand U6822 (N_6822,N_4887,N_5080);
or U6823 (N_6823,N_4463,N_5321);
or U6824 (N_6824,N_4859,N_4041);
xor U6825 (N_6825,N_4303,N_4476);
nor U6826 (N_6826,N_5196,N_5034);
xnor U6827 (N_6827,N_4255,N_4165);
and U6828 (N_6828,N_5613,N_4586);
nor U6829 (N_6829,N_5096,N_5201);
or U6830 (N_6830,N_4794,N_4513);
nor U6831 (N_6831,N_5805,N_5161);
or U6832 (N_6832,N_4043,N_4413);
or U6833 (N_6833,N_5612,N_4407);
xnor U6834 (N_6834,N_5233,N_4403);
nand U6835 (N_6835,N_4121,N_4948);
or U6836 (N_6836,N_5905,N_4974);
nor U6837 (N_6837,N_5824,N_4995);
and U6838 (N_6838,N_4920,N_4605);
xnor U6839 (N_6839,N_4234,N_5510);
xnor U6840 (N_6840,N_5262,N_4533);
or U6841 (N_6841,N_5985,N_4104);
and U6842 (N_6842,N_5364,N_4661);
or U6843 (N_6843,N_4888,N_5509);
or U6844 (N_6844,N_5395,N_5935);
or U6845 (N_6845,N_5675,N_5663);
and U6846 (N_6846,N_4447,N_5752);
or U6847 (N_6847,N_5763,N_5979);
and U6848 (N_6848,N_4271,N_5372);
or U6849 (N_6849,N_5362,N_4478);
nor U6850 (N_6850,N_5009,N_4477);
xor U6851 (N_6851,N_5107,N_5728);
or U6852 (N_6852,N_4500,N_5464);
xor U6853 (N_6853,N_5614,N_5956);
or U6854 (N_6854,N_4088,N_5742);
and U6855 (N_6855,N_4224,N_4439);
and U6856 (N_6856,N_5750,N_4677);
and U6857 (N_6857,N_5772,N_4399);
nor U6858 (N_6858,N_5670,N_4548);
nor U6859 (N_6859,N_5873,N_5143);
nand U6860 (N_6860,N_4695,N_4538);
nand U6861 (N_6861,N_5064,N_5774);
or U6862 (N_6862,N_5018,N_5793);
nor U6863 (N_6863,N_5340,N_5914);
nor U6864 (N_6864,N_5641,N_5157);
nor U6865 (N_6865,N_4921,N_4717);
nand U6866 (N_6866,N_5698,N_5872);
nand U6867 (N_6867,N_4918,N_5767);
xor U6868 (N_6868,N_5908,N_5446);
nor U6869 (N_6869,N_4486,N_4101);
xnor U6870 (N_6870,N_4565,N_5682);
and U6871 (N_6871,N_5560,N_4494);
nor U6872 (N_6872,N_4295,N_4539);
xnor U6873 (N_6873,N_5351,N_4515);
nor U6874 (N_6874,N_5910,N_5846);
nand U6875 (N_6875,N_5111,N_4857);
xor U6876 (N_6876,N_5361,N_4283);
nand U6877 (N_6877,N_5387,N_4664);
or U6878 (N_6878,N_4313,N_4581);
and U6879 (N_6879,N_5426,N_5382);
or U6880 (N_6880,N_4112,N_4506);
nor U6881 (N_6881,N_4352,N_4844);
nand U6882 (N_6882,N_5658,N_4861);
or U6883 (N_6883,N_4757,N_5939);
nand U6884 (N_6884,N_5809,N_5261);
and U6885 (N_6885,N_4438,N_4917);
and U6886 (N_6886,N_5041,N_4601);
or U6887 (N_6887,N_4682,N_4152);
xnor U6888 (N_6888,N_4081,N_4577);
nand U6889 (N_6889,N_4194,N_4561);
xor U6890 (N_6890,N_4962,N_4761);
nand U6891 (N_6891,N_5174,N_5019);
and U6892 (N_6892,N_4585,N_4700);
or U6893 (N_6893,N_5596,N_5436);
nor U6894 (N_6894,N_4400,N_5603);
and U6895 (N_6895,N_5816,N_4216);
nor U6896 (N_6896,N_5482,N_5408);
or U6897 (N_6897,N_4393,N_5517);
xnor U6898 (N_6898,N_5855,N_5186);
xnor U6899 (N_6899,N_4139,N_5496);
nand U6900 (N_6900,N_5582,N_4643);
nor U6901 (N_6901,N_5553,N_4343);
nand U6902 (N_6902,N_4713,N_4675);
nor U6903 (N_6903,N_5419,N_5359);
nor U6904 (N_6904,N_5788,N_5141);
nand U6905 (N_6905,N_4966,N_5172);
or U6906 (N_6906,N_4242,N_5150);
or U6907 (N_6907,N_4988,N_5821);
or U6908 (N_6908,N_5301,N_4215);
nand U6909 (N_6909,N_5478,N_5461);
xor U6910 (N_6910,N_4126,N_4305);
or U6911 (N_6911,N_4527,N_5208);
xor U6912 (N_6912,N_4573,N_4074);
and U6913 (N_6913,N_4053,N_5524);
or U6914 (N_6914,N_4896,N_5303);
and U6915 (N_6915,N_4072,N_5627);
nor U6916 (N_6916,N_4290,N_5389);
or U6917 (N_6917,N_5845,N_5982);
or U6918 (N_6918,N_5002,N_4563);
nor U6919 (N_6919,N_5754,N_5327);
xor U6920 (N_6920,N_4686,N_5040);
or U6921 (N_6921,N_4579,N_4524);
or U6922 (N_6922,N_4960,N_4637);
nand U6923 (N_6923,N_5615,N_4518);
and U6924 (N_6924,N_4470,N_5802);
nand U6925 (N_6925,N_5602,N_4740);
nand U6926 (N_6926,N_4173,N_4045);
nor U6927 (N_6927,N_4755,N_5021);
nand U6928 (N_6928,N_5996,N_5695);
nand U6929 (N_6929,N_4782,N_5300);
or U6930 (N_6930,N_4019,N_4946);
and U6931 (N_6931,N_4869,N_4684);
nor U6932 (N_6932,N_5885,N_4482);
nand U6933 (N_6933,N_4388,N_4480);
xor U6934 (N_6934,N_5067,N_4002);
xor U6935 (N_6935,N_4311,N_4113);
nand U6936 (N_6936,N_4558,N_4839);
xnor U6937 (N_6937,N_4979,N_5176);
nand U6938 (N_6938,N_4145,N_5822);
or U6939 (N_6939,N_5089,N_4714);
and U6940 (N_6940,N_4405,N_4807);
and U6941 (N_6941,N_5108,N_4097);
nand U6942 (N_6942,N_4842,N_4969);
or U6943 (N_6943,N_5491,N_4127);
xor U6944 (N_6944,N_5354,N_4359);
nand U6945 (N_6945,N_5916,N_5541);
xor U6946 (N_6946,N_4334,N_4706);
xnor U6947 (N_6947,N_5715,N_4876);
or U6948 (N_6948,N_4813,N_4010);
nor U6949 (N_6949,N_5853,N_5680);
nand U6950 (N_6950,N_5350,N_5330);
nor U6951 (N_6951,N_5355,N_4512);
and U6952 (N_6952,N_4729,N_5293);
xor U6953 (N_6953,N_5516,N_5053);
and U6954 (N_6954,N_4256,N_4826);
nand U6955 (N_6955,N_4814,N_4770);
nand U6956 (N_6956,N_4726,N_5238);
xnor U6957 (N_6957,N_4065,N_4198);
and U6958 (N_6958,N_4567,N_5322);
nand U6959 (N_6959,N_4883,N_5838);
nand U6960 (N_6960,N_5911,N_4497);
nand U6961 (N_6961,N_4076,N_5858);
nor U6962 (N_6962,N_4817,N_5789);
and U6963 (N_6963,N_5957,N_5486);
nor U6964 (N_6964,N_4288,N_4535);
nor U6965 (N_6965,N_5328,N_4108);
nor U6966 (N_6966,N_4622,N_5972);
nor U6967 (N_6967,N_4444,N_4251);
nor U6968 (N_6968,N_4409,N_5933);
nand U6969 (N_6969,N_5230,N_5232);
nor U6970 (N_6970,N_5231,N_5076);
xor U6971 (N_6971,N_4155,N_4386);
or U6972 (N_6972,N_5442,N_4211);
nand U6973 (N_6973,N_5662,N_4201);
nand U6974 (N_6974,N_4337,N_4199);
and U6975 (N_6975,N_5200,N_5175);
or U6976 (N_6976,N_5891,N_4937);
nand U6977 (N_6977,N_4059,N_5250);
and U6978 (N_6978,N_5185,N_4263);
or U6979 (N_6979,N_4926,N_5338);
nand U6980 (N_6980,N_4593,N_5811);
and U6981 (N_6981,N_5837,N_5216);
or U6982 (N_6982,N_4971,N_5725);
xor U6983 (N_6983,N_4116,N_4750);
xor U6984 (N_6984,N_5310,N_4096);
xnor U6985 (N_6985,N_4153,N_4329);
and U6986 (N_6986,N_5889,N_5296);
xor U6987 (N_6987,N_4281,N_5743);
and U6988 (N_6988,N_5219,N_4133);
nand U6989 (N_6989,N_4846,N_4537);
and U6990 (N_6990,N_5343,N_5158);
xor U6991 (N_6991,N_4580,N_5398);
nand U6992 (N_6992,N_4259,N_5689);
nor U6993 (N_6993,N_4054,N_5035);
nor U6994 (N_6994,N_4302,N_4425);
xnor U6995 (N_6995,N_5650,N_4254);
nor U6996 (N_6996,N_4374,N_4250);
nor U6997 (N_6997,N_4737,N_4853);
nor U6998 (N_6998,N_4050,N_4809);
nand U6999 (N_6999,N_4504,N_5494);
nor U7000 (N_7000,N_5792,N_5121);
nand U7001 (N_7001,N_4478,N_5359);
nor U7002 (N_7002,N_4845,N_5039);
and U7003 (N_7003,N_4389,N_4024);
or U7004 (N_7004,N_4687,N_5808);
nand U7005 (N_7005,N_4754,N_4606);
and U7006 (N_7006,N_4695,N_4072);
and U7007 (N_7007,N_4444,N_4318);
nand U7008 (N_7008,N_4073,N_4760);
and U7009 (N_7009,N_4659,N_4656);
nand U7010 (N_7010,N_4497,N_5104);
xor U7011 (N_7011,N_5450,N_4906);
xor U7012 (N_7012,N_5516,N_4296);
and U7013 (N_7013,N_5051,N_4873);
xnor U7014 (N_7014,N_5389,N_5447);
or U7015 (N_7015,N_5161,N_4853);
and U7016 (N_7016,N_4943,N_4503);
nor U7017 (N_7017,N_5910,N_5397);
or U7018 (N_7018,N_5203,N_5008);
xnor U7019 (N_7019,N_4303,N_4586);
xor U7020 (N_7020,N_4873,N_5630);
xnor U7021 (N_7021,N_5281,N_5822);
or U7022 (N_7022,N_4092,N_4280);
nand U7023 (N_7023,N_5564,N_5637);
nor U7024 (N_7024,N_5312,N_5486);
nor U7025 (N_7025,N_4457,N_5931);
xor U7026 (N_7026,N_4752,N_5738);
nand U7027 (N_7027,N_4751,N_4328);
xor U7028 (N_7028,N_4461,N_5794);
nand U7029 (N_7029,N_5853,N_5502);
and U7030 (N_7030,N_5683,N_4264);
and U7031 (N_7031,N_5256,N_5297);
or U7032 (N_7032,N_4804,N_5243);
and U7033 (N_7033,N_5599,N_5493);
and U7034 (N_7034,N_5083,N_4279);
nand U7035 (N_7035,N_4734,N_5112);
nand U7036 (N_7036,N_4047,N_5163);
nor U7037 (N_7037,N_4833,N_5602);
or U7038 (N_7038,N_4858,N_5487);
and U7039 (N_7039,N_5886,N_4377);
and U7040 (N_7040,N_4467,N_5246);
xnor U7041 (N_7041,N_5713,N_4052);
and U7042 (N_7042,N_5222,N_4742);
and U7043 (N_7043,N_5819,N_4348);
nor U7044 (N_7044,N_5142,N_5174);
xor U7045 (N_7045,N_5563,N_4434);
nor U7046 (N_7046,N_4948,N_5750);
and U7047 (N_7047,N_5342,N_5203);
nor U7048 (N_7048,N_5436,N_4225);
and U7049 (N_7049,N_5513,N_5230);
nand U7050 (N_7050,N_4781,N_4026);
and U7051 (N_7051,N_5438,N_5023);
xnor U7052 (N_7052,N_4736,N_4218);
or U7053 (N_7053,N_4606,N_4628);
nand U7054 (N_7054,N_4940,N_4581);
nand U7055 (N_7055,N_4324,N_5442);
nor U7056 (N_7056,N_4236,N_5151);
nor U7057 (N_7057,N_5743,N_4075);
nor U7058 (N_7058,N_4896,N_4911);
nand U7059 (N_7059,N_5657,N_4903);
nor U7060 (N_7060,N_5552,N_5180);
and U7061 (N_7061,N_4053,N_5468);
nor U7062 (N_7062,N_4101,N_4292);
xor U7063 (N_7063,N_4024,N_4739);
nand U7064 (N_7064,N_5005,N_4618);
nand U7065 (N_7065,N_4956,N_4097);
or U7066 (N_7066,N_5842,N_4732);
nor U7067 (N_7067,N_5596,N_5769);
and U7068 (N_7068,N_4616,N_4279);
xnor U7069 (N_7069,N_4346,N_4326);
nand U7070 (N_7070,N_5752,N_5189);
nand U7071 (N_7071,N_5729,N_4010);
or U7072 (N_7072,N_4046,N_5739);
nand U7073 (N_7073,N_5619,N_4780);
and U7074 (N_7074,N_4989,N_5384);
or U7075 (N_7075,N_4030,N_4659);
nor U7076 (N_7076,N_4139,N_5803);
and U7077 (N_7077,N_4394,N_4685);
nand U7078 (N_7078,N_5682,N_5103);
nand U7079 (N_7079,N_5759,N_4404);
and U7080 (N_7080,N_4585,N_5302);
nand U7081 (N_7081,N_5295,N_5590);
xor U7082 (N_7082,N_5476,N_4954);
nor U7083 (N_7083,N_4987,N_5721);
and U7084 (N_7084,N_4307,N_5885);
or U7085 (N_7085,N_5116,N_5579);
nor U7086 (N_7086,N_5246,N_5710);
and U7087 (N_7087,N_4079,N_5527);
nor U7088 (N_7088,N_4837,N_5164);
xnor U7089 (N_7089,N_5113,N_5485);
or U7090 (N_7090,N_4669,N_5178);
and U7091 (N_7091,N_5488,N_4234);
nor U7092 (N_7092,N_4429,N_5588);
nand U7093 (N_7093,N_5207,N_5979);
xor U7094 (N_7094,N_5196,N_4081);
xor U7095 (N_7095,N_5582,N_4221);
nand U7096 (N_7096,N_4749,N_4797);
and U7097 (N_7097,N_5813,N_4883);
xnor U7098 (N_7098,N_4701,N_5099);
and U7099 (N_7099,N_4411,N_4140);
xor U7100 (N_7100,N_4227,N_5639);
nand U7101 (N_7101,N_4189,N_5576);
nor U7102 (N_7102,N_5752,N_5131);
and U7103 (N_7103,N_5898,N_5923);
xnor U7104 (N_7104,N_4932,N_5259);
or U7105 (N_7105,N_4113,N_5716);
or U7106 (N_7106,N_4655,N_4123);
nand U7107 (N_7107,N_5089,N_4027);
nor U7108 (N_7108,N_4637,N_5775);
or U7109 (N_7109,N_5587,N_4434);
or U7110 (N_7110,N_4804,N_4707);
xor U7111 (N_7111,N_4857,N_5702);
nand U7112 (N_7112,N_5927,N_5223);
and U7113 (N_7113,N_5577,N_4933);
xor U7114 (N_7114,N_5785,N_5810);
xor U7115 (N_7115,N_5394,N_4834);
and U7116 (N_7116,N_5426,N_5120);
nand U7117 (N_7117,N_5313,N_4103);
or U7118 (N_7118,N_5123,N_4582);
nor U7119 (N_7119,N_5553,N_4903);
or U7120 (N_7120,N_5120,N_5444);
and U7121 (N_7121,N_5819,N_5300);
or U7122 (N_7122,N_5832,N_4911);
or U7123 (N_7123,N_4130,N_5656);
and U7124 (N_7124,N_5351,N_5011);
nor U7125 (N_7125,N_4303,N_4468);
and U7126 (N_7126,N_5210,N_4138);
or U7127 (N_7127,N_4173,N_5103);
xor U7128 (N_7128,N_5620,N_5349);
nor U7129 (N_7129,N_4895,N_5469);
xor U7130 (N_7130,N_5568,N_4518);
xnor U7131 (N_7131,N_5188,N_4032);
nor U7132 (N_7132,N_4129,N_4795);
or U7133 (N_7133,N_5327,N_5187);
nand U7134 (N_7134,N_5808,N_4108);
xor U7135 (N_7135,N_4800,N_4494);
and U7136 (N_7136,N_4629,N_5800);
nand U7137 (N_7137,N_5379,N_4895);
xor U7138 (N_7138,N_5919,N_5952);
and U7139 (N_7139,N_4472,N_5462);
nor U7140 (N_7140,N_5248,N_4427);
and U7141 (N_7141,N_4040,N_5070);
nand U7142 (N_7142,N_5561,N_5535);
or U7143 (N_7143,N_4953,N_4763);
xnor U7144 (N_7144,N_5052,N_5888);
and U7145 (N_7145,N_5122,N_5061);
nor U7146 (N_7146,N_5828,N_4085);
xor U7147 (N_7147,N_4355,N_4917);
nand U7148 (N_7148,N_4227,N_5582);
xor U7149 (N_7149,N_5960,N_4828);
and U7150 (N_7150,N_4829,N_5606);
nand U7151 (N_7151,N_5642,N_4281);
nor U7152 (N_7152,N_4903,N_5819);
or U7153 (N_7153,N_5608,N_4627);
xor U7154 (N_7154,N_5264,N_5354);
or U7155 (N_7155,N_5955,N_4711);
and U7156 (N_7156,N_5172,N_4891);
nand U7157 (N_7157,N_5696,N_4077);
and U7158 (N_7158,N_4851,N_5138);
and U7159 (N_7159,N_5656,N_4247);
nand U7160 (N_7160,N_4892,N_5225);
or U7161 (N_7161,N_5051,N_5534);
nand U7162 (N_7162,N_4122,N_5996);
xnor U7163 (N_7163,N_4304,N_4720);
nor U7164 (N_7164,N_5091,N_4009);
xor U7165 (N_7165,N_4519,N_5569);
and U7166 (N_7166,N_4632,N_4899);
and U7167 (N_7167,N_4713,N_4578);
xor U7168 (N_7168,N_4560,N_4729);
nand U7169 (N_7169,N_5013,N_5188);
or U7170 (N_7170,N_4880,N_4607);
nand U7171 (N_7171,N_4972,N_4847);
nor U7172 (N_7172,N_5108,N_4486);
nor U7173 (N_7173,N_4204,N_5212);
or U7174 (N_7174,N_4658,N_5098);
nor U7175 (N_7175,N_4610,N_4467);
nor U7176 (N_7176,N_4437,N_5327);
or U7177 (N_7177,N_5765,N_4033);
nor U7178 (N_7178,N_4279,N_4115);
nor U7179 (N_7179,N_5735,N_5669);
nand U7180 (N_7180,N_4438,N_5521);
nand U7181 (N_7181,N_5515,N_4640);
nor U7182 (N_7182,N_5270,N_4841);
nand U7183 (N_7183,N_4421,N_5468);
or U7184 (N_7184,N_4455,N_5162);
xor U7185 (N_7185,N_4650,N_4588);
nor U7186 (N_7186,N_5541,N_5118);
and U7187 (N_7187,N_5216,N_5151);
or U7188 (N_7188,N_5848,N_4892);
nand U7189 (N_7189,N_5186,N_4433);
nor U7190 (N_7190,N_5567,N_4454);
nand U7191 (N_7191,N_5935,N_4958);
or U7192 (N_7192,N_4279,N_4267);
and U7193 (N_7193,N_5492,N_5667);
nand U7194 (N_7194,N_4054,N_4937);
nand U7195 (N_7195,N_5618,N_4771);
and U7196 (N_7196,N_5219,N_4172);
nand U7197 (N_7197,N_5648,N_5912);
and U7198 (N_7198,N_5998,N_4707);
or U7199 (N_7199,N_4005,N_5252);
nor U7200 (N_7200,N_5523,N_4339);
and U7201 (N_7201,N_5333,N_5109);
nand U7202 (N_7202,N_4700,N_4791);
and U7203 (N_7203,N_5923,N_4769);
and U7204 (N_7204,N_4264,N_5332);
or U7205 (N_7205,N_5675,N_4591);
nor U7206 (N_7206,N_4652,N_4468);
nor U7207 (N_7207,N_4437,N_5578);
or U7208 (N_7208,N_4046,N_5078);
nand U7209 (N_7209,N_4754,N_4629);
xor U7210 (N_7210,N_5185,N_5370);
and U7211 (N_7211,N_4701,N_4006);
and U7212 (N_7212,N_4578,N_5877);
nor U7213 (N_7213,N_5430,N_4415);
and U7214 (N_7214,N_4758,N_4815);
or U7215 (N_7215,N_4890,N_4770);
xnor U7216 (N_7216,N_4808,N_5987);
nand U7217 (N_7217,N_5287,N_5226);
and U7218 (N_7218,N_5882,N_4412);
and U7219 (N_7219,N_5074,N_4842);
or U7220 (N_7220,N_4219,N_4190);
nor U7221 (N_7221,N_4628,N_4305);
nor U7222 (N_7222,N_4467,N_4379);
xor U7223 (N_7223,N_4133,N_5521);
and U7224 (N_7224,N_5551,N_5112);
nor U7225 (N_7225,N_4368,N_5101);
nor U7226 (N_7226,N_4971,N_5205);
nor U7227 (N_7227,N_4026,N_4765);
nand U7228 (N_7228,N_5881,N_4030);
nand U7229 (N_7229,N_4930,N_5682);
nor U7230 (N_7230,N_5435,N_4719);
nor U7231 (N_7231,N_4680,N_4727);
and U7232 (N_7232,N_4977,N_4663);
nand U7233 (N_7233,N_5957,N_5993);
nand U7234 (N_7234,N_4451,N_5774);
or U7235 (N_7235,N_4325,N_5058);
xor U7236 (N_7236,N_5771,N_5110);
nor U7237 (N_7237,N_4516,N_4922);
or U7238 (N_7238,N_4579,N_5339);
or U7239 (N_7239,N_5438,N_4756);
and U7240 (N_7240,N_5912,N_5088);
nand U7241 (N_7241,N_4139,N_5003);
and U7242 (N_7242,N_4361,N_4356);
xnor U7243 (N_7243,N_4749,N_5735);
or U7244 (N_7244,N_5773,N_5265);
or U7245 (N_7245,N_4935,N_4393);
or U7246 (N_7246,N_5093,N_4934);
and U7247 (N_7247,N_5605,N_4363);
or U7248 (N_7248,N_5607,N_4456);
xnor U7249 (N_7249,N_4929,N_5294);
nor U7250 (N_7250,N_5460,N_4559);
and U7251 (N_7251,N_5867,N_5029);
nand U7252 (N_7252,N_5173,N_5782);
and U7253 (N_7253,N_5174,N_5821);
and U7254 (N_7254,N_4875,N_4843);
xnor U7255 (N_7255,N_5092,N_4029);
nand U7256 (N_7256,N_4336,N_4563);
xnor U7257 (N_7257,N_4866,N_5426);
and U7258 (N_7258,N_4735,N_5769);
xor U7259 (N_7259,N_4901,N_4217);
nor U7260 (N_7260,N_5790,N_5125);
nand U7261 (N_7261,N_4891,N_4948);
nand U7262 (N_7262,N_5247,N_5457);
nor U7263 (N_7263,N_4165,N_5557);
xor U7264 (N_7264,N_5899,N_4310);
and U7265 (N_7265,N_5760,N_5428);
or U7266 (N_7266,N_4695,N_5379);
and U7267 (N_7267,N_5453,N_5444);
and U7268 (N_7268,N_4400,N_5027);
xnor U7269 (N_7269,N_5844,N_4493);
nor U7270 (N_7270,N_4748,N_4807);
or U7271 (N_7271,N_5693,N_5878);
or U7272 (N_7272,N_5889,N_4470);
nor U7273 (N_7273,N_4079,N_4974);
nor U7274 (N_7274,N_4568,N_5490);
or U7275 (N_7275,N_5653,N_4536);
xor U7276 (N_7276,N_4677,N_5920);
xor U7277 (N_7277,N_4092,N_4847);
or U7278 (N_7278,N_5243,N_5320);
or U7279 (N_7279,N_4379,N_5486);
or U7280 (N_7280,N_5517,N_4351);
and U7281 (N_7281,N_4401,N_4697);
or U7282 (N_7282,N_5678,N_4799);
and U7283 (N_7283,N_4012,N_4354);
nor U7284 (N_7284,N_4864,N_5890);
nand U7285 (N_7285,N_5593,N_5247);
xor U7286 (N_7286,N_4818,N_4247);
nand U7287 (N_7287,N_5608,N_4278);
nor U7288 (N_7288,N_5001,N_5730);
nand U7289 (N_7289,N_4057,N_5837);
or U7290 (N_7290,N_4360,N_4698);
or U7291 (N_7291,N_4376,N_4780);
nor U7292 (N_7292,N_5180,N_4191);
or U7293 (N_7293,N_5494,N_5325);
xor U7294 (N_7294,N_4250,N_4267);
nand U7295 (N_7295,N_4143,N_5645);
nor U7296 (N_7296,N_5457,N_4923);
xor U7297 (N_7297,N_4525,N_4924);
or U7298 (N_7298,N_4955,N_4452);
or U7299 (N_7299,N_4412,N_4742);
and U7300 (N_7300,N_4634,N_4933);
nor U7301 (N_7301,N_5745,N_5501);
and U7302 (N_7302,N_5035,N_5916);
xnor U7303 (N_7303,N_5509,N_5821);
nor U7304 (N_7304,N_5594,N_4397);
and U7305 (N_7305,N_4556,N_5619);
nand U7306 (N_7306,N_5537,N_4623);
or U7307 (N_7307,N_5893,N_4826);
nor U7308 (N_7308,N_4878,N_5412);
or U7309 (N_7309,N_5724,N_4596);
or U7310 (N_7310,N_5256,N_4301);
nand U7311 (N_7311,N_4151,N_5090);
and U7312 (N_7312,N_5753,N_4200);
nor U7313 (N_7313,N_5218,N_4883);
xor U7314 (N_7314,N_4545,N_5318);
and U7315 (N_7315,N_5383,N_4225);
nand U7316 (N_7316,N_4934,N_4368);
and U7317 (N_7317,N_5795,N_5070);
xnor U7318 (N_7318,N_4874,N_5621);
nand U7319 (N_7319,N_4857,N_4591);
xor U7320 (N_7320,N_5718,N_4404);
nor U7321 (N_7321,N_5003,N_5342);
nor U7322 (N_7322,N_4999,N_5284);
nand U7323 (N_7323,N_5222,N_5255);
and U7324 (N_7324,N_5938,N_4455);
and U7325 (N_7325,N_5130,N_5611);
and U7326 (N_7326,N_4151,N_4129);
or U7327 (N_7327,N_5228,N_5720);
nand U7328 (N_7328,N_5695,N_4580);
nor U7329 (N_7329,N_5786,N_5083);
or U7330 (N_7330,N_4614,N_4304);
nand U7331 (N_7331,N_4766,N_4170);
nand U7332 (N_7332,N_5671,N_5593);
nor U7333 (N_7333,N_5049,N_5293);
nand U7334 (N_7334,N_5041,N_4406);
and U7335 (N_7335,N_5310,N_4228);
or U7336 (N_7336,N_5823,N_4733);
xnor U7337 (N_7337,N_4235,N_4873);
nor U7338 (N_7338,N_5000,N_5551);
nor U7339 (N_7339,N_4079,N_4020);
nor U7340 (N_7340,N_4776,N_4593);
nand U7341 (N_7341,N_5124,N_4146);
or U7342 (N_7342,N_5419,N_4229);
or U7343 (N_7343,N_4482,N_5632);
xor U7344 (N_7344,N_4655,N_5942);
xnor U7345 (N_7345,N_5391,N_5724);
and U7346 (N_7346,N_4139,N_4659);
nor U7347 (N_7347,N_4836,N_4967);
or U7348 (N_7348,N_5424,N_5388);
nand U7349 (N_7349,N_4015,N_5008);
nand U7350 (N_7350,N_4626,N_5269);
nor U7351 (N_7351,N_5426,N_5396);
and U7352 (N_7352,N_4043,N_4251);
nand U7353 (N_7353,N_4077,N_5473);
xor U7354 (N_7354,N_4130,N_5665);
and U7355 (N_7355,N_4090,N_4214);
nor U7356 (N_7356,N_4176,N_5776);
or U7357 (N_7357,N_5957,N_5740);
xor U7358 (N_7358,N_5302,N_4860);
and U7359 (N_7359,N_5019,N_5592);
or U7360 (N_7360,N_4711,N_4387);
xor U7361 (N_7361,N_4934,N_5160);
nor U7362 (N_7362,N_5126,N_4157);
nand U7363 (N_7363,N_5977,N_4191);
or U7364 (N_7364,N_4040,N_5240);
nand U7365 (N_7365,N_5932,N_5136);
xnor U7366 (N_7366,N_5362,N_5006);
or U7367 (N_7367,N_4987,N_4085);
nand U7368 (N_7368,N_4565,N_4320);
xor U7369 (N_7369,N_5626,N_5461);
and U7370 (N_7370,N_4857,N_5441);
and U7371 (N_7371,N_4304,N_5081);
xnor U7372 (N_7372,N_4171,N_4100);
or U7373 (N_7373,N_4233,N_4503);
xnor U7374 (N_7374,N_5820,N_4507);
or U7375 (N_7375,N_4551,N_4773);
nor U7376 (N_7376,N_4209,N_5797);
or U7377 (N_7377,N_4851,N_5862);
nor U7378 (N_7378,N_4770,N_4011);
xor U7379 (N_7379,N_5894,N_4479);
nand U7380 (N_7380,N_5737,N_5825);
and U7381 (N_7381,N_4700,N_4566);
nor U7382 (N_7382,N_4451,N_5694);
nand U7383 (N_7383,N_5944,N_4973);
nand U7384 (N_7384,N_5233,N_4561);
xnor U7385 (N_7385,N_4769,N_4757);
or U7386 (N_7386,N_4756,N_4706);
nand U7387 (N_7387,N_5327,N_5400);
nor U7388 (N_7388,N_4014,N_5969);
and U7389 (N_7389,N_4657,N_5520);
nand U7390 (N_7390,N_4025,N_4751);
and U7391 (N_7391,N_5772,N_5207);
nand U7392 (N_7392,N_5754,N_5495);
or U7393 (N_7393,N_5557,N_4962);
and U7394 (N_7394,N_5109,N_5307);
nand U7395 (N_7395,N_5246,N_4378);
nor U7396 (N_7396,N_5189,N_4533);
nor U7397 (N_7397,N_4492,N_4632);
nand U7398 (N_7398,N_4740,N_4300);
nor U7399 (N_7399,N_4921,N_5057);
and U7400 (N_7400,N_5503,N_4826);
and U7401 (N_7401,N_4574,N_5267);
nor U7402 (N_7402,N_5102,N_4235);
nand U7403 (N_7403,N_4071,N_5286);
nand U7404 (N_7404,N_4062,N_5936);
nor U7405 (N_7405,N_5337,N_4141);
nand U7406 (N_7406,N_5544,N_4075);
nor U7407 (N_7407,N_4793,N_4470);
or U7408 (N_7408,N_5956,N_4273);
nor U7409 (N_7409,N_4084,N_4707);
or U7410 (N_7410,N_5120,N_5198);
xnor U7411 (N_7411,N_5219,N_5258);
or U7412 (N_7412,N_4350,N_5413);
xnor U7413 (N_7413,N_5268,N_5628);
nor U7414 (N_7414,N_5223,N_5538);
and U7415 (N_7415,N_5615,N_4026);
nand U7416 (N_7416,N_5210,N_5780);
nand U7417 (N_7417,N_5148,N_5032);
nand U7418 (N_7418,N_4155,N_4767);
and U7419 (N_7419,N_5237,N_5551);
xor U7420 (N_7420,N_5876,N_4182);
or U7421 (N_7421,N_4129,N_5030);
nand U7422 (N_7422,N_5493,N_4050);
nor U7423 (N_7423,N_5858,N_5056);
nor U7424 (N_7424,N_4723,N_5962);
and U7425 (N_7425,N_5584,N_5733);
or U7426 (N_7426,N_5894,N_4996);
xor U7427 (N_7427,N_4360,N_4440);
and U7428 (N_7428,N_4346,N_4650);
xor U7429 (N_7429,N_4904,N_4599);
or U7430 (N_7430,N_5764,N_5665);
and U7431 (N_7431,N_4350,N_5368);
nand U7432 (N_7432,N_4579,N_4361);
and U7433 (N_7433,N_4797,N_4375);
nor U7434 (N_7434,N_4397,N_5421);
xnor U7435 (N_7435,N_5151,N_4896);
nor U7436 (N_7436,N_4882,N_5859);
and U7437 (N_7437,N_4343,N_4342);
nand U7438 (N_7438,N_4343,N_4159);
and U7439 (N_7439,N_5648,N_4592);
xor U7440 (N_7440,N_5410,N_5261);
or U7441 (N_7441,N_5418,N_5117);
and U7442 (N_7442,N_4021,N_5919);
nand U7443 (N_7443,N_4325,N_5911);
xor U7444 (N_7444,N_5567,N_4905);
and U7445 (N_7445,N_5636,N_5016);
nor U7446 (N_7446,N_4392,N_5661);
xor U7447 (N_7447,N_4009,N_4202);
xnor U7448 (N_7448,N_4894,N_4814);
and U7449 (N_7449,N_5387,N_5664);
nand U7450 (N_7450,N_4992,N_5757);
nand U7451 (N_7451,N_4714,N_4870);
nor U7452 (N_7452,N_5616,N_5841);
and U7453 (N_7453,N_4814,N_5269);
or U7454 (N_7454,N_5408,N_5176);
nor U7455 (N_7455,N_4595,N_5714);
and U7456 (N_7456,N_4597,N_5684);
and U7457 (N_7457,N_5500,N_5743);
nand U7458 (N_7458,N_4807,N_4234);
xor U7459 (N_7459,N_4411,N_4306);
nand U7460 (N_7460,N_4643,N_5514);
xor U7461 (N_7461,N_5686,N_5023);
xnor U7462 (N_7462,N_4114,N_4012);
or U7463 (N_7463,N_5189,N_5221);
or U7464 (N_7464,N_5520,N_4977);
and U7465 (N_7465,N_5486,N_4937);
nor U7466 (N_7466,N_4954,N_4129);
or U7467 (N_7467,N_4822,N_4906);
xor U7468 (N_7468,N_4388,N_5769);
and U7469 (N_7469,N_5649,N_5675);
and U7470 (N_7470,N_5333,N_5743);
nand U7471 (N_7471,N_4919,N_5622);
nand U7472 (N_7472,N_5609,N_5949);
nand U7473 (N_7473,N_4980,N_4520);
nand U7474 (N_7474,N_4967,N_4302);
and U7475 (N_7475,N_4235,N_4154);
nand U7476 (N_7476,N_4532,N_4977);
nor U7477 (N_7477,N_4508,N_4998);
nand U7478 (N_7478,N_4925,N_4513);
and U7479 (N_7479,N_5235,N_5265);
xor U7480 (N_7480,N_4052,N_4541);
nand U7481 (N_7481,N_5200,N_4119);
and U7482 (N_7482,N_5022,N_4719);
and U7483 (N_7483,N_4886,N_4687);
nor U7484 (N_7484,N_4027,N_5431);
xor U7485 (N_7485,N_4780,N_5926);
nand U7486 (N_7486,N_4545,N_4314);
nor U7487 (N_7487,N_5900,N_5408);
and U7488 (N_7488,N_4724,N_4878);
or U7489 (N_7489,N_5976,N_5435);
nor U7490 (N_7490,N_5305,N_5693);
nor U7491 (N_7491,N_4065,N_4109);
or U7492 (N_7492,N_4546,N_4265);
nand U7493 (N_7493,N_4389,N_5951);
nor U7494 (N_7494,N_5742,N_5619);
xnor U7495 (N_7495,N_4346,N_5197);
and U7496 (N_7496,N_4562,N_4324);
xor U7497 (N_7497,N_4528,N_4040);
and U7498 (N_7498,N_5456,N_5265);
xor U7499 (N_7499,N_4205,N_5347);
or U7500 (N_7500,N_5187,N_5722);
and U7501 (N_7501,N_5582,N_4737);
nand U7502 (N_7502,N_5525,N_5825);
xnor U7503 (N_7503,N_4069,N_4056);
xnor U7504 (N_7504,N_5045,N_4533);
nor U7505 (N_7505,N_5313,N_5964);
nand U7506 (N_7506,N_5645,N_5535);
nor U7507 (N_7507,N_5186,N_5379);
or U7508 (N_7508,N_5225,N_4787);
xor U7509 (N_7509,N_4324,N_5048);
nor U7510 (N_7510,N_5459,N_5209);
xor U7511 (N_7511,N_5801,N_5490);
and U7512 (N_7512,N_5744,N_4419);
nand U7513 (N_7513,N_5930,N_4768);
xnor U7514 (N_7514,N_5298,N_5460);
xor U7515 (N_7515,N_4362,N_5365);
nand U7516 (N_7516,N_5556,N_5100);
or U7517 (N_7517,N_4381,N_4833);
xnor U7518 (N_7518,N_5167,N_5332);
or U7519 (N_7519,N_4219,N_4582);
xnor U7520 (N_7520,N_4359,N_5337);
and U7521 (N_7521,N_5851,N_5462);
nand U7522 (N_7522,N_5457,N_4022);
nor U7523 (N_7523,N_5486,N_4223);
or U7524 (N_7524,N_5383,N_5438);
or U7525 (N_7525,N_5343,N_5112);
nand U7526 (N_7526,N_4678,N_4253);
or U7527 (N_7527,N_4781,N_5772);
xor U7528 (N_7528,N_5068,N_4862);
and U7529 (N_7529,N_4634,N_5859);
nor U7530 (N_7530,N_5051,N_5050);
nor U7531 (N_7531,N_5764,N_4721);
or U7532 (N_7532,N_4766,N_4773);
xnor U7533 (N_7533,N_5709,N_5486);
xnor U7534 (N_7534,N_4296,N_4064);
or U7535 (N_7535,N_4575,N_4543);
nor U7536 (N_7536,N_4443,N_4764);
nand U7537 (N_7537,N_5956,N_5734);
nor U7538 (N_7538,N_5339,N_4777);
or U7539 (N_7539,N_4022,N_4365);
nand U7540 (N_7540,N_4689,N_4670);
and U7541 (N_7541,N_4549,N_4115);
or U7542 (N_7542,N_5365,N_4934);
nor U7543 (N_7543,N_5161,N_5800);
nor U7544 (N_7544,N_5437,N_4535);
and U7545 (N_7545,N_4571,N_4156);
or U7546 (N_7546,N_4271,N_5178);
nand U7547 (N_7547,N_4624,N_5559);
nand U7548 (N_7548,N_4768,N_5251);
nand U7549 (N_7549,N_4616,N_4178);
or U7550 (N_7550,N_5268,N_4791);
or U7551 (N_7551,N_5975,N_5827);
nor U7552 (N_7552,N_4758,N_5291);
or U7553 (N_7553,N_4789,N_5080);
nand U7554 (N_7554,N_5242,N_4917);
xor U7555 (N_7555,N_4175,N_4038);
xor U7556 (N_7556,N_5715,N_4303);
nand U7557 (N_7557,N_4949,N_5094);
and U7558 (N_7558,N_5609,N_5639);
and U7559 (N_7559,N_4640,N_4546);
nor U7560 (N_7560,N_5043,N_4831);
nand U7561 (N_7561,N_4556,N_4808);
or U7562 (N_7562,N_4739,N_5789);
and U7563 (N_7563,N_4074,N_4002);
nor U7564 (N_7564,N_4348,N_4134);
nor U7565 (N_7565,N_5696,N_4613);
nand U7566 (N_7566,N_5053,N_4954);
and U7567 (N_7567,N_5696,N_5654);
nand U7568 (N_7568,N_5829,N_5080);
xnor U7569 (N_7569,N_5034,N_5421);
xor U7570 (N_7570,N_5243,N_4298);
nor U7571 (N_7571,N_4706,N_4273);
nand U7572 (N_7572,N_5670,N_4983);
xor U7573 (N_7573,N_4897,N_5354);
xor U7574 (N_7574,N_5534,N_5444);
nor U7575 (N_7575,N_5115,N_4837);
and U7576 (N_7576,N_4122,N_5185);
xor U7577 (N_7577,N_4307,N_4988);
nand U7578 (N_7578,N_4557,N_5927);
xor U7579 (N_7579,N_5009,N_5602);
and U7580 (N_7580,N_4353,N_5439);
xnor U7581 (N_7581,N_5947,N_4236);
xnor U7582 (N_7582,N_5934,N_4066);
nor U7583 (N_7583,N_5120,N_4500);
xnor U7584 (N_7584,N_5350,N_5848);
xor U7585 (N_7585,N_4908,N_5476);
nand U7586 (N_7586,N_4987,N_4976);
nor U7587 (N_7587,N_4877,N_5414);
nor U7588 (N_7588,N_5644,N_5244);
nor U7589 (N_7589,N_4087,N_5188);
nor U7590 (N_7590,N_5396,N_4704);
nor U7591 (N_7591,N_5024,N_4258);
and U7592 (N_7592,N_4712,N_4783);
nand U7593 (N_7593,N_5097,N_5866);
and U7594 (N_7594,N_5095,N_4167);
or U7595 (N_7595,N_4786,N_5650);
xnor U7596 (N_7596,N_4685,N_5584);
nand U7597 (N_7597,N_4979,N_4596);
xor U7598 (N_7598,N_5424,N_4989);
and U7599 (N_7599,N_4016,N_5722);
or U7600 (N_7600,N_4868,N_5727);
nand U7601 (N_7601,N_5727,N_4652);
nor U7602 (N_7602,N_4788,N_5319);
nand U7603 (N_7603,N_5126,N_5780);
xor U7604 (N_7604,N_5670,N_4343);
nand U7605 (N_7605,N_4793,N_4269);
nor U7606 (N_7606,N_5464,N_4206);
or U7607 (N_7607,N_5362,N_5169);
nor U7608 (N_7608,N_5648,N_5560);
nand U7609 (N_7609,N_4646,N_4203);
and U7610 (N_7610,N_4389,N_4961);
nand U7611 (N_7611,N_4665,N_4536);
or U7612 (N_7612,N_4638,N_5893);
nand U7613 (N_7613,N_5305,N_5548);
and U7614 (N_7614,N_5673,N_5124);
nor U7615 (N_7615,N_5272,N_4506);
nand U7616 (N_7616,N_4114,N_4737);
xnor U7617 (N_7617,N_4253,N_5079);
xnor U7618 (N_7618,N_5018,N_5543);
and U7619 (N_7619,N_4505,N_5648);
nor U7620 (N_7620,N_5003,N_5448);
nand U7621 (N_7621,N_4275,N_4779);
nor U7622 (N_7622,N_4944,N_5378);
and U7623 (N_7623,N_5424,N_5993);
nand U7624 (N_7624,N_4881,N_5494);
xor U7625 (N_7625,N_4833,N_4317);
xor U7626 (N_7626,N_5805,N_4362);
nand U7627 (N_7627,N_4636,N_5621);
and U7628 (N_7628,N_4445,N_4103);
or U7629 (N_7629,N_5328,N_4125);
and U7630 (N_7630,N_5805,N_5548);
and U7631 (N_7631,N_4987,N_4703);
and U7632 (N_7632,N_5514,N_4540);
nor U7633 (N_7633,N_5884,N_4448);
or U7634 (N_7634,N_5462,N_5643);
nor U7635 (N_7635,N_5233,N_5195);
and U7636 (N_7636,N_4980,N_5963);
xnor U7637 (N_7637,N_5000,N_5344);
or U7638 (N_7638,N_4104,N_5640);
and U7639 (N_7639,N_4362,N_5101);
nand U7640 (N_7640,N_4151,N_5877);
nor U7641 (N_7641,N_5281,N_5408);
nand U7642 (N_7642,N_5430,N_5731);
nor U7643 (N_7643,N_5418,N_4495);
nor U7644 (N_7644,N_4857,N_5614);
or U7645 (N_7645,N_5886,N_4041);
or U7646 (N_7646,N_4203,N_5103);
nand U7647 (N_7647,N_4907,N_5005);
nand U7648 (N_7648,N_5837,N_4706);
and U7649 (N_7649,N_5768,N_5558);
or U7650 (N_7650,N_5611,N_5896);
nor U7651 (N_7651,N_4904,N_5124);
and U7652 (N_7652,N_5798,N_5957);
nor U7653 (N_7653,N_5448,N_4938);
or U7654 (N_7654,N_4715,N_4000);
and U7655 (N_7655,N_4352,N_5923);
or U7656 (N_7656,N_5923,N_4899);
and U7657 (N_7657,N_5389,N_4497);
nand U7658 (N_7658,N_5862,N_5709);
nand U7659 (N_7659,N_4454,N_5018);
nor U7660 (N_7660,N_4231,N_5261);
nand U7661 (N_7661,N_4968,N_4838);
and U7662 (N_7662,N_4829,N_5510);
nand U7663 (N_7663,N_4563,N_4335);
nand U7664 (N_7664,N_4287,N_5832);
xnor U7665 (N_7665,N_4288,N_5195);
nand U7666 (N_7666,N_5349,N_4888);
and U7667 (N_7667,N_5109,N_4031);
and U7668 (N_7668,N_5307,N_4133);
or U7669 (N_7669,N_5779,N_5174);
and U7670 (N_7670,N_4326,N_4200);
and U7671 (N_7671,N_4042,N_4698);
xor U7672 (N_7672,N_4413,N_4278);
and U7673 (N_7673,N_5483,N_4998);
nand U7674 (N_7674,N_5695,N_4677);
nor U7675 (N_7675,N_4287,N_4522);
and U7676 (N_7676,N_5320,N_5636);
and U7677 (N_7677,N_4254,N_4754);
xnor U7678 (N_7678,N_5844,N_5027);
and U7679 (N_7679,N_5294,N_4435);
nand U7680 (N_7680,N_5994,N_5496);
or U7681 (N_7681,N_5573,N_5097);
or U7682 (N_7682,N_4283,N_4298);
or U7683 (N_7683,N_5643,N_4091);
or U7684 (N_7684,N_4503,N_4704);
or U7685 (N_7685,N_4354,N_5508);
nor U7686 (N_7686,N_4036,N_5272);
and U7687 (N_7687,N_5726,N_5034);
nand U7688 (N_7688,N_5354,N_5307);
nand U7689 (N_7689,N_5904,N_4268);
nand U7690 (N_7690,N_5670,N_5104);
xnor U7691 (N_7691,N_4116,N_4707);
xor U7692 (N_7692,N_4257,N_5031);
nand U7693 (N_7693,N_4636,N_5264);
xor U7694 (N_7694,N_5725,N_5707);
xor U7695 (N_7695,N_5447,N_4560);
xnor U7696 (N_7696,N_5689,N_5959);
and U7697 (N_7697,N_4547,N_5384);
xnor U7698 (N_7698,N_4269,N_5980);
and U7699 (N_7699,N_4467,N_4417);
nand U7700 (N_7700,N_4349,N_4608);
or U7701 (N_7701,N_4102,N_4336);
xnor U7702 (N_7702,N_4015,N_4302);
nor U7703 (N_7703,N_5993,N_5550);
and U7704 (N_7704,N_4938,N_5686);
or U7705 (N_7705,N_4351,N_5657);
or U7706 (N_7706,N_5727,N_4384);
or U7707 (N_7707,N_5743,N_5718);
xnor U7708 (N_7708,N_4369,N_5744);
nor U7709 (N_7709,N_5883,N_5762);
and U7710 (N_7710,N_4117,N_4616);
and U7711 (N_7711,N_4972,N_5567);
nor U7712 (N_7712,N_5980,N_5743);
nor U7713 (N_7713,N_4238,N_5667);
nor U7714 (N_7714,N_5977,N_5798);
xor U7715 (N_7715,N_4403,N_4901);
nor U7716 (N_7716,N_4765,N_5299);
xnor U7717 (N_7717,N_5874,N_4905);
or U7718 (N_7718,N_4092,N_4774);
xor U7719 (N_7719,N_4306,N_4294);
nand U7720 (N_7720,N_5170,N_5052);
nor U7721 (N_7721,N_5831,N_4346);
xnor U7722 (N_7722,N_4268,N_4496);
or U7723 (N_7723,N_4781,N_4208);
xor U7724 (N_7724,N_4485,N_4099);
xnor U7725 (N_7725,N_4930,N_5171);
nand U7726 (N_7726,N_4921,N_4722);
nor U7727 (N_7727,N_4381,N_4506);
or U7728 (N_7728,N_4182,N_4609);
nor U7729 (N_7729,N_5407,N_5240);
nand U7730 (N_7730,N_4556,N_4670);
and U7731 (N_7731,N_4586,N_5727);
and U7732 (N_7732,N_4577,N_5351);
or U7733 (N_7733,N_5665,N_5481);
nand U7734 (N_7734,N_4988,N_4710);
nor U7735 (N_7735,N_5221,N_4140);
and U7736 (N_7736,N_4392,N_4474);
and U7737 (N_7737,N_5105,N_4939);
nor U7738 (N_7738,N_5324,N_4688);
or U7739 (N_7739,N_5638,N_4654);
xor U7740 (N_7740,N_5872,N_5039);
and U7741 (N_7741,N_5524,N_4063);
or U7742 (N_7742,N_5361,N_5362);
or U7743 (N_7743,N_4539,N_4556);
nor U7744 (N_7744,N_5034,N_5022);
xor U7745 (N_7745,N_5777,N_5448);
nand U7746 (N_7746,N_4021,N_5224);
and U7747 (N_7747,N_5345,N_5195);
or U7748 (N_7748,N_5730,N_4092);
and U7749 (N_7749,N_4120,N_4883);
nor U7750 (N_7750,N_4579,N_4262);
xor U7751 (N_7751,N_4858,N_5693);
xor U7752 (N_7752,N_5847,N_4594);
xor U7753 (N_7753,N_4385,N_5331);
and U7754 (N_7754,N_5315,N_5457);
or U7755 (N_7755,N_4034,N_4178);
nand U7756 (N_7756,N_5989,N_4130);
nor U7757 (N_7757,N_5379,N_4630);
nor U7758 (N_7758,N_4918,N_5655);
nand U7759 (N_7759,N_5743,N_5106);
nand U7760 (N_7760,N_4691,N_5205);
and U7761 (N_7761,N_5706,N_5940);
or U7762 (N_7762,N_5889,N_5382);
and U7763 (N_7763,N_4335,N_4573);
xnor U7764 (N_7764,N_5979,N_5155);
nor U7765 (N_7765,N_5155,N_4897);
or U7766 (N_7766,N_5373,N_5735);
and U7767 (N_7767,N_5930,N_4044);
nand U7768 (N_7768,N_5394,N_5430);
nor U7769 (N_7769,N_5317,N_4206);
or U7770 (N_7770,N_5172,N_4134);
or U7771 (N_7771,N_4030,N_5808);
nor U7772 (N_7772,N_4321,N_4818);
or U7773 (N_7773,N_5437,N_5282);
nand U7774 (N_7774,N_5373,N_4472);
or U7775 (N_7775,N_5108,N_4729);
and U7776 (N_7776,N_5852,N_5568);
or U7777 (N_7777,N_4240,N_5060);
and U7778 (N_7778,N_4284,N_5532);
nor U7779 (N_7779,N_5693,N_4867);
or U7780 (N_7780,N_4847,N_4177);
xnor U7781 (N_7781,N_4342,N_5040);
nand U7782 (N_7782,N_5705,N_5356);
nor U7783 (N_7783,N_5379,N_4153);
xnor U7784 (N_7784,N_4728,N_5242);
nor U7785 (N_7785,N_5143,N_5614);
or U7786 (N_7786,N_4357,N_4065);
nor U7787 (N_7787,N_5270,N_4801);
or U7788 (N_7788,N_4977,N_5864);
nor U7789 (N_7789,N_5773,N_5069);
xnor U7790 (N_7790,N_4124,N_4625);
nor U7791 (N_7791,N_4084,N_5400);
nand U7792 (N_7792,N_5139,N_4364);
or U7793 (N_7793,N_5202,N_5144);
or U7794 (N_7794,N_5879,N_4816);
or U7795 (N_7795,N_5362,N_4135);
nor U7796 (N_7796,N_5726,N_4691);
xnor U7797 (N_7797,N_4599,N_4204);
or U7798 (N_7798,N_4890,N_4478);
and U7799 (N_7799,N_4770,N_5445);
and U7800 (N_7800,N_4504,N_5532);
or U7801 (N_7801,N_4873,N_5544);
xor U7802 (N_7802,N_4495,N_5235);
nor U7803 (N_7803,N_5267,N_5892);
nor U7804 (N_7804,N_4498,N_4949);
nand U7805 (N_7805,N_5311,N_4114);
or U7806 (N_7806,N_5280,N_5358);
and U7807 (N_7807,N_4206,N_4678);
or U7808 (N_7808,N_4433,N_4396);
and U7809 (N_7809,N_5950,N_4099);
and U7810 (N_7810,N_5802,N_4095);
nand U7811 (N_7811,N_5583,N_4505);
and U7812 (N_7812,N_5258,N_4410);
nor U7813 (N_7813,N_5447,N_4024);
xor U7814 (N_7814,N_4297,N_5997);
or U7815 (N_7815,N_4388,N_4862);
nor U7816 (N_7816,N_4222,N_4417);
or U7817 (N_7817,N_5735,N_4265);
and U7818 (N_7818,N_4642,N_5336);
nand U7819 (N_7819,N_5434,N_4835);
nor U7820 (N_7820,N_4062,N_5830);
nand U7821 (N_7821,N_4107,N_5395);
nand U7822 (N_7822,N_5080,N_5848);
xnor U7823 (N_7823,N_5190,N_4984);
xnor U7824 (N_7824,N_5279,N_4524);
xor U7825 (N_7825,N_5440,N_4405);
nor U7826 (N_7826,N_4534,N_5174);
nand U7827 (N_7827,N_5415,N_4323);
xnor U7828 (N_7828,N_4958,N_5327);
nor U7829 (N_7829,N_5977,N_4674);
xnor U7830 (N_7830,N_5337,N_4430);
or U7831 (N_7831,N_5904,N_5438);
nand U7832 (N_7832,N_4683,N_5789);
nand U7833 (N_7833,N_5435,N_5772);
nor U7834 (N_7834,N_5280,N_4380);
or U7835 (N_7835,N_4470,N_5720);
or U7836 (N_7836,N_4330,N_5174);
xnor U7837 (N_7837,N_5969,N_5491);
or U7838 (N_7838,N_5160,N_4553);
nor U7839 (N_7839,N_5783,N_4324);
nand U7840 (N_7840,N_4636,N_5906);
or U7841 (N_7841,N_4423,N_4300);
nand U7842 (N_7842,N_4486,N_4533);
xnor U7843 (N_7843,N_5965,N_4265);
and U7844 (N_7844,N_5704,N_5504);
or U7845 (N_7845,N_5894,N_4229);
or U7846 (N_7846,N_4944,N_5783);
and U7847 (N_7847,N_5664,N_5491);
nand U7848 (N_7848,N_4168,N_5160);
and U7849 (N_7849,N_4401,N_5933);
or U7850 (N_7850,N_5700,N_5669);
xor U7851 (N_7851,N_5581,N_4201);
and U7852 (N_7852,N_4050,N_4968);
nand U7853 (N_7853,N_4622,N_4052);
and U7854 (N_7854,N_4263,N_5991);
or U7855 (N_7855,N_5557,N_5915);
or U7856 (N_7856,N_5976,N_5320);
nor U7857 (N_7857,N_5149,N_5002);
xnor U7858 (N_7858,N_4893,N_5085);
or U7859 (N_7859,N_5186,N_4356);
or U7860 (N_7860,N_5105,N_4926);
xor U7861 (N_7861,N_4160,N_4516);
nand U7862 (N_7862,N_5639,N_4243);
or U7863 (N_7863,N_5007,N_5756);
nor U7864 (N_7864,N_5965,N_4240);
xnor U7865 (N_7865,N_5089,N_4300);
xor U7866 (N_7866,N_5621,N_5772);
and U7867 (N_7867,N_5976,N_5784);
or U7868 (N_7868,N_4628,N_5969);
and U7869 (N_7869,N_5914,N_5070);
nand U7870 (N_7870,N_4281,N_4359);
nor U7871 (N_7871,N_4225,N_4393);
or U7872 (N_7872,N_5803,N_4667);
nor U7873 (N_7873,N_4526,N_5346);
or U7874 (N_7874,N_4216,N_5102);
nand U7875 (N_7875,N_5438,N_4240);
nor U7876 (N_7876,N_4691,N_4328);
xor U7877 (N_7877,N_4701,N_4287);
or U7878 (N_7878,N_5673,N_4548);
nor U7879 (N_7879,N_4795,N_4174);
and U7880 (N_7880,N_5837,N_5813);
nor U7881 (N_7881,N_5236,N_5291);
and U7882 (N_7882,N_5912,N_4418);
nor U7883 (N_7883,N_4647,N_5950);
nand U7884 (N_7884,N_4205,N_5666);
or U7885 (N_7885,N_4974,N_4791);
nor U7886 (N_7886,N_4478,N_5568);
nand U7887 (N_7887,N_4581,N_4158);
nor U7888 (N_7888,N_5419,N_5122);
xor U7889 (N_7889,N_5661,N_5529);
and U7890 (N_7890,N_4652,N_4513);
nand U7891 (N_7891,N_4655,N_4112);
and U7892 (N_7892,N_4688,N_5194);
nand U7893 (N_7893,N_5668,N_5103);
xnor U7894 (N_7894,N_4519,N_5056);
nor U7895 (N_7895,N_5177,N_5985);
or U7896 (N_7896,N_5518,N_4101);
nor U7897 (N_7897,N_4293,N_5755);
nand U7898 (N_7898,N_4357,N_4544);
and U7899 (N_7899,N_5305,N_5737);
or U7900 (N_7900,N_4139,N_5661);
and U7901 (N_7901,N_5737,N_4726);
nand U7902 (N_7902,N_4907,N_5119);
nand U7903 (N_7903,N_4797,N_4038);
xor U7904 (N_7904,N_4642,N_4312);
nor U7905 (N_7905,N_5017,N_5313);
nand U7906 (N_7906,N_4859,N_4872);
or U7907 (N_7907,N_4009,N_4241);
xnor U7908 (N_7908,N_5763,N_5749);
or U7909 (N_7909,N_5812,N_4130);
and U7910 (N_7910,N_5653,N_4627);
nand U7911 (N_7911,N_4946,N_5752);
nor U7912 (N_7912,N_4983,N_4866);
or U7913 (N_7913,N_5228,N_5592);
nand U7914 (N_7914,N_4360,N_4917);
nor U7915 (N_7915,N_4379,N_4382);
nor U7916 (N_7916,N_4100,N_5824);
and U7917 (N_7917,N_5577,N_4207);
nor U7918 (N_7918,N_5682,N_5075);
xnor U7919 (N_7919,N_5172,N_5793);
and U7920 (N_7920,N_4688,N_5875);
nand U7921 (N_7921,N_4423,N_4214);
nor U7922 (N_7922,N_4065,N_5505);
nor U7923 (N_7923,N_4223,N_5732);
nand U7924 (N_7924,N_5145,N_4339);
nand U7925 (N_7925,N_4760,N_4292);
nand U7926 (N_7926,N_4350,N_4739);
and U7927 (N_7927,N_4303,N_5129);
or U7928 (N_7928,N_5228,N_5643);
nand U7929 (N_7929,N_4459,N_5379);
xnor U7930 (N_7930,N_4938,N_5495);
or U7931 (N_7931,N_5484,N_4179);
nand U7932 (N_7932,N_4545,N_4713);
nor U7933 (N_7933,N_4172,N_5608);
nand U7934 (N_7934,N_5646,N_4803);
or U7935 (N_7935,N_4082,N_5733);
nor U7936 (N_7936,N_4896,N_5720);
xor U7937 (N_7937,N_4310,N_4247);
or U7938 (N_7938,N_4802,N_4591);
nor U7939 (N_7939,N_4125,N_4880);
xnor U7940 (N_7940,N_5530,N_4746);
xnor U7941 (N_7941,N_5914,N_4486);
nand U7942 (N_7942,N_5158,N_5987);
or U7943 (N_7943,N_5212,N_5231);
or U7944 (N_7944,N_5739,N_4509);
and U7945 (N_7945,N_5648,N_4733);
nand U7946 (N_7946,N_4168,N_4895);
and U7947 (N_7947,N_5207,N_5309);
nor U7948 (N_7948,N_4548,N_4818);
xor U7949 (N_7949,N_5392,N_4974);
nor U7950 (N_7950,N_4424,N_5410);
nor U7951 (N_7951,N_5156,N_5026);
nor U7952 (N_7952,N_5386,N_4775);
nand U7953 (N_7953,N_4104,N_4488);
nand U7954 (N_7954,N_5795,N_4589);
or U7955 (N_7955,N_4935,N_5701);
nor U7956 (N_7956,N_4098,N_4093);
xor U7957 (N_7957,N_4412,N_4185);
and U7958 (N_7958,N_4074,N_5169);
nor U7959 (N_7959,N_4037,N_4885);
xnor U7960 (N_7960,N_4327,N_4244);
or U7961 (N_7961,N_5774,N_4962);
xnor U7962 (N_7962,N_4025,N_5550);
or U7963 (N_7963,N_4122,N_4534);
and U7964 (N_7964,N_4809,N_5488);
and U7965 (N_7965,N_5384,N_5016);
nor U7966 (N_7966,N_4194,N_5436);
xor U7967 (N_7967,N_4973,N_4809);
nand U7968 (N_7968,N_4332,N_5652);
or U7969 (N_7969,N_4108,N_5311);
and U7970 (N_7970,N_4376,N_4940);
nor U7971 (N_7971,N_5014,N_5423);
nor U7972 (N_7972,N_4112,N_5731);
nor U7973 (N_7973,N_5990,N_5948);
and U7974 (N_7974,N_4572,N_4705);
xnor U7975 (N_7975,N_5255,N_5686);
nor U7976 (N_7976,N_5958,N_5768);
and U7977 (N_7977,N_4801,N_4430);
nor U7978 (N_7978,N_4287,N_4311);
and U7979 (N_7979,N_5679,N_4022);
nand U7980 (N_7980,N_4902,N_4104);
or U7981 (N_7981,N_5650,N_4844);
xnor U7982 (N_7982,N_4533,N_5938);
and U7983 (N_7983,N_5417,N_5146);
nand U7984 (N_7984,N_5624,N_5630);
nand U7985 (N_7985,N_4318,N_4961);
xor U7986 (N_7986,N_4033,N_4338);
nand U7987 (N_7987,N_4346,N_4749);
xnor U7988 (N_7988,N_5258,N_5689);
and U7989 (N_7989,N_4286,N_5008);
and U7990 (N_7990,N_4071,N_5685);
xnor U7991 (N_7991,N_5197,N_5215);
or U7992 (N_7992,N_5408,N_4779);
nand U7993 (N_7993,N_5895,N_5058);
and U7994 (N_7994,N_5965,N_5981);
and U7995 (N_7995,N_5633,N_5253);
xor U7996 (N_7996,N_4441,N_4311);
or U7997 (N_7997,N_4280,N_4361);
nand U7998 (N_7998,N_5303,N_5601);
xor U7999 (N_7999,N_5194,N_5060);
and U8000 (N_8000,N_7250,N_6335);
nand U8001 (N_8001,N_7965,N_7600);
or U8002 (N_8002,N_6956,N_6122);
and U8003 (N_8003,N_6561,N_7426);
or U8004 (N_8004,N_7184,N_7593);
or U8005 (N_8005,N_6011,N_6704);
nor U8006 (N_8006,N_6052,N_6054);
or U8007 (N_8007,N_6450,N_6237);
xnor U8008 (N_8008,N_6766,N_7298);
nor U8009 (N_8009,N_6026,N_6400);
nor U8010 (N_8010,N_6253,N_6777);
nor U8011 (N_8011,N_6048,N_6735);
and U8012 (N_8012,N_7626,N_7098);
xnor U8013 (N_8013,N_6648,N_6817);
and U8014 (N_8014,N_6062,N_7716);
nand U8015 (N_8015,N_6476,N_7677);
nand U8016 (N_8016,N_7427,N_6964);
xnor U8017 (N_8017,N_7378,N_6812);
nor U8018 (N_8018,N_6258,N_7203);
nor U8019 (N_8019,N_6886,N_7934);
nor U8020 (N_8020,N_6053,N_6774);
and U8021 (N_8021,N_7812,N_6613);
nand U8022 (N_8022,N_6734,N_7731);
xor U8023 (N_8023,N_7562,N_7108);
or U8024 (N_8024,N_7324,N_6304);
nand U8025 (N_8025,N_7929,N_7846);
and U8026 (N_8026,N_6203,N_6342);
nor U8027 (N_8027,N_7615,N_7864);
nor U8028 (N_8028,N_7199,N_6222);
nor U8029 (N_8029,N_6155,N_7560);
xnor U8030 (N_8030,N_6263,N_7419);
and U8031 (N_8031,N_7479,N_6978);
nand U8032 (N_8032,N_6290,N_6680);
nor U8033 (N_8033,N_7340,N_7890);
xnor U8034 (N_8034,N_6971,N_7939);
nand U8035 (N_8035,N_6835,N_7636);
or U8036 (N_8036,N_7178,N_6439);
nor U8037 (N_8037,N_7473,N_6230);
nand U8038 (N_8038,N_6841,N_7102);
nand U8039 (N_8039,N_7577,N_6514);
or U8040 (N_8040,N_7829,N_7551);
nor U8041 (N_8041,N_6204,N_6435);
xor U8042 (N_8042,N_7632,N_6621);
nor U8043 (N_8043,N_7573,N_6034);
and U8044 (N_8044,N_7281,N_7079);
nor U8045 (N_8045,N_7580,N_7943);
xor U8046 (N_8046,N_6536,N_6483);
or U8047 (N_8047,N_6152,N_7645);
nor U8048 (N_8048,N_7305,N_6270);
nand U8049 (N_8049,N_7141,N_7416);
nand U8050 (N_8050,N_7706,N_6803);
nor U8051 (N_8051,N_6606,N_6518);
nor U8052 (N_8052,N_6816,N_7388);
xnor U8053 (N_8053,N_7154,N_7819);
and U8054 (N_8054,N_7086,N_7741);
or U8055 (N_8055,N_6714,N_6516);
or U8056 (N_8056,N_6453,N_6138);
nand U8057 (N_8057,N_7055,N_7208);
nor U8058 (N_8058,N_6020,N_7485);
or U8059 (N_8059,N_6460,N_7041);
nor U8060 (N_8060,N_6437,N_7885);
and U8061 (N_8061,N_6392,N_6854);
xnor U8062 (N_8062,N_7631,N_7163);
nor U8063 (N_8063,N_7268,N_6616);
and U8064 (N_8064,N_6467,N_6194);
nor U8065 (N_8065,N_7630,N_7145);
xnor U8066 (N_8066,N_7902,N_7985);
and U8067 (N_8067,N_6883,N_7285);
nand U8068 (N_8068,N_6355,N_6209);
xor U8069 (N_8069,N_7288,N_7532);
nor U8070 (N_8070,N_7494,N_6749);
nand U8071 (N_8071,N_6170,N_7231);
nand U8072 (N_8072,N_7164,N_7724);
nand U8073 (N_8073,N_6889,N_6504);
xor U8074 (N_8074,N_7100,N_7151);
nor U8075 (N_8075,N_7865,N_6140);
xor U8076 (N_8076,N_6281,N_6119);
nand U8077 (N_8077,N_6753,N_6544);
xnor U8078 (N_8078,N_6456,N_6583);
xor U8079 (N_8079,N_7161,N_6895);
or U8080 (N_8080,N_6452,N_6855);
or U8081 (N_8081,N_7099,N_6322);
nor U8082 (N_8082,N_7065,N_7085);
nor U8083 (N_8083,N_6389,N_7059);
nand U8084 (N_8084,N_7362,N_7693);
and U8085 (N_8085,N_6490,N_7404);
nand U8086 (N_8086,N_6401,N_7802);
xor U8087 (N_8087,N_7094,N_6495);
or U8088 (N_8088,N_6842,N_6655);
and U8089 (N_8089,N_7245,N_7444);
or U8090 (N_8090,N_6343,N_7173);
nor U8091 (N_8091,N_6684,N_7591);
nor U8092 (N_8092,N_7522,N_7465);
nand U8093 (N_8093,N_6614,N_7612);
xnor U8094 (N_8094,N_7247,N_7189);
nand U8095 (N_8095,N_7538,N_7990);
xor U8096 (N_8096,N_7499,N_7243);
xor U8097 (N_8097,N_6876,N_7110);
or U8098 (N_8098,N_6185,N_7228);
or U8099 (N_8099,N_6254,N_7824);
or U8100 (N_8100,N_6158,N_6031);
nand U8101 (N_8101,N_7949,N_7814);
nand U8102 (N_8102,N_6033,N_6162);
and U8103 (N_8103,N_7654,N_7042);
xnor U8104 (N_8104,N_6782,N_7491);
nor U8105 (N_8105,N_6550,N_7563);
nor U8106 (N_8106,N_7413,N_7169);
nor U8107 (N_8107,N_7549,N_6967);
nor U8108 (N_8108,N_7239,N_6791);
xnor U8109 (N_8109,N_6719,N_7862);
nand U8110 (N_8110,N_6920,N_6353);
or U8111 (N_8111,N_7174,N_7816);
or U8112 (N_8112,N_7686,N_7472);
nand U8113 (N_8113,N_6507,N_7193);
nand U8114 (N_8114,N_7194,N_6294);
or U8115 (N_8115,N_7223,N_6288);
nor U8116 (N_8116,N_6933,N_7260);
nor U8117 (N_8117,N_7953,N_6756);
nor U8118 (N_8118,N_7477,N_7035);
nand U8119 (N_8119,N_6136,N_7519);
nand U8120 (N_8120,N_6412,N_6298);
nor U8121 (N_8121,N_7070,N_7253);
xnor U8122 (N_8122,N_7905,N_7221);
or U8123 (N_8123,N_6528,N_7502);
nor U8124 (N_8124,N_7906,N_7021);
and U8125 (N_8125,N_7635,N_7157);
xnor U8126 (N_8126,N_7980,N_7928);
xor U8127 (N_8127,N_6218,N_6983);
nand U8128 (N_8128,N_7412,N_7304);
xnor U8129 (N_8129,N_6320,N_6084);
and U8130 (N_8130,N_6403,N_6159);
nor U8131 (N_8131,N_6906,N_7515);
or U8132 (N_8132,N_6571,N_6407);
and U8133 (N_8133,N_6718,N_7770);
and U8134 (N_8134,N_7020,N_7651);
nand U8135 (N_8135,N_7040,N_6010);
and U8136 (N_8136,N_7841,N_7940);
xnor U8137 (N_8137,N_7698,N_7667);
and U8138 (N_8138,N_6941,N_6307);
or U8139 (N_8139,N_6458,N_6802);
and U8140 (N_8140,N_7227,N_7782);
or U8141 (N_8141,N_7142,N_7136);
and U8142 (N_8142,N_7387,N_7637);
or U8143 (N_8143,N_7492,N_6018);
xor U8144 (N_8144,N_6709,N_6293);
xor U8145 (N_8145,N_6757,N_7312);
and U8146 (N_8146,N_7742,N_7868);
and U8147 (N_8147,N_6447,N_7808);
or U8148 (N_8148,N_6511,N_6787);
nand U8149 (N_8149,N_6679,N_6029);
or U8150 (N_8150,N_6661,N_6969);
xnor U8151 (N_8151,N_6847,N_6068);
xnor U8152 (N_8152,N_7175,N_6283);
xor U8153 (N_8153,N_7694,N_6313);
nand U8154 (N_8154,N_7728,N_7118);
nand U8155 (N_8155,N_7353,N_6006);
and U8156 (N_8156,N_6897,N_7555);
nor U8157 (N_8157,N_7652,N_6934);
and U8158 (N_8158,N_6344,N_7537);
or U8159 (N_8159,N_7323,N_6760);
nor U8160 (N_8160,N_6585,N_6821);
nor U8161 (N_8161,N_6903,N_6094);
or U8162 (N_8162,N_7454,N_7279);
xor U8163 (N_8163,N_6824,N_6347);
xnor U8164 (N_8164,N_7955,N_7958);
or U8165 (N_8165,N_7548,N_6475);
and U8166 (N_8166,N_6594,N_7254);
nor U8167 (N_8167,N_7013,N_6994);
nand U8168 (N_8168,N_7893,N_6051);
xnor U8169 (N_8169,N_6697,N_6144);
and U8170 (N_8170,N_6852,N_6239);
or U8171 (N_8171,N_6043,N_6190);
nor U8172 (N_8172,N_6484,N_7750);
or U8173 (N_8173,N_7986,N_7536);
and U8174 (N_8174,N_6323,N_7030);
xnor U8175 (N_8175,N_7096,N_6589);
and U8176 (N_8176,N_7503,N_7213);
nor U8177 (N_8177,N_6394,N_7963);
xor U8178 (N_8178,N_7500,N_7382);
and U8179 (N_8179,N_7753,N_7345);
xor U8180 (N_8180,N_7371,N_7606);
xor U8181 (N_8181,N_7639,N_7291);
xnor U8182 (N_8182,N_6701,N_6745);
xnor U8183 (N_8183,N_6037,N_6692);
and U8184 (N_8184,N_7735,N_7439);
or U8185 (N_8185,N_6512,N_7521);
nand U8186 (N_8186,N_7048,N_7874);
xnor U8187 (N_8187,N_6539,N_7861);
nor U8188 (N_8188,N_6527,N_6337);
or U8189 (N_8189,N_6302,N_7379);
nor U8190 (N_8190,N_7188,N_6038);
and U8191 (N_8191,N_6195,N_7396);
xnor U8192 (N_8192,N_6091,N_7331);
or U8193 (N_8193,N_7398,N_6861);
nand U8194 (N_8194,N_6169,N_7924);
or U8195 (N_8195,N_6954,N_7621);
xnor U8196 (N_8196,N_7091,N_6417);
and U8197 (N_8197,N_6461,N_7729);
or U8198 (N_8198,N_6397,N_7341);
nor U8199 (N_8199,N_7681,N_7229);
nand U8200 (N_8200,N_6063,N_6265);
or U8201 (N_8201,N_7003,N_7389);
nand U8202 (N_8202,N_7689,N_6117);
and U8203 (N_8203,N_7329,N_7992);
nor U8204 (N_8204,N_6945,N_6455);
and U8205 (N_8205,N_6255,N_7124);
and U8206 (N_8206,N_6911,N_6665);
nor U8207 (N_8207,N_7273,N_6578);
xnor U8208 (N_8208,N_6459,N_6794);
nor U8209 (N_8209,N_7881,N_7008);
xor U8210 (N_8210,N_7895,N_7987);
or U8211 (N_8211,N_6433,N_6211);
nand U8212 (N_8212,N_7400,N_6910);
nor U8213 (N_8213,N_7438,N_6348);
xnor U8214 (N_8214,N_7374,N_7025);
and U8215 (N_8215,N_7226,N_7550);
xnor U8216 (N_8216,N_7925,N_6380);
nand U8217 (N_8217,N_6815,N_7220);
xor U8218 (N_8218,N_6001,N_7872);
nand U8219 (N_8219,N_6295,N_7642);
xor U8220 (N_8220,N_7166,N_7710);
or U8221 (N_8221,N_7453,N_7797);
xnor U8222 (N_8222,N_6378,N_6105);
and U8223 (N_8223,N_7669,N_7431);
and U8224 (N_8224,N_7837,N_6073);
or U8225 (N_8225,N_6558,N_6365);
nor U8226 (N_8226,N_7113,N_6810);
nor U8227 (N_8227,N_6305,N_7576);
xnor U8228 (N_8228,N_7763,N_7531);
or U8229 (N_8229,N_7878,N_6932);
or U8230 (N_8230,N_6332,N_7259);
or U8231 (N_8231,N_7185,N_7355);
nand U8232 (N_8232,N_7687,N_6915);
or U8233 (N_8233,N_7338,N_7311);
xor U8234 (N_8234,N_6425,N_7719);
xnor U8235 (N_8235,N_7903,N_6390);
nand U8236 (N_8236,N_6501,N_6268);
and U8237 (N_8237,N_6864,N_6765);
and U8238 (N_8238,N_6838,N_7931);
nor U8239 (N_8239,N_6940,N_6074);
nand U8240 (N_8240,N_7832,N_7232);
and U8241 (N_8241,N_6731,N_6723);
and U8242 (N_8242,N_7659,N_6752);
and U8243 (N_8243,N_6232,N_7927);
nand U8244 (N_8244,N_6272,N_7590);
and U8245 (N_8245,N_7230,N_7700);
nor U8246 (N_8246,N_7442,N_7557);
or U8247 (N_8247,N_7073,N_6900);
or U8248 (N_8248,N_7033,N_6115);
nand U8249 (N_8249,N_6381,N_7678);
nor U8250 (N_8250,N_7249,N_7801);
nor U8251 (N_8251,N_7083,N_6975);
or U8252 (N_8252,N_6354,N_6212);
xor U8253 (N_8253,N_6167,N_7684);
nand U8254 (N_8254,N_6958,N_7674);
nor U8255 (N_8255,N_7514,N_6896);
or U8256 (N_8256,N_7045,N_7209);
and U8257 (N_8257,N_7775,N_7322);
xnor U8258 (N_8258,N_7219,N_6179);
xor U8259 (N_8259,N_7214,N_6286);
nor U8260 (N_8260,N_7391,N_7395);
nor U8261 (N_8261,N_7655,N_7968);
nor U8262 (N_8262,N_6235,N_6375);
or U8263 (N_8263,N_6667,N_6617);
xor U8264 (N_8264,N_7607,N_6454);
xor U8265 (N_8265,N_7506,N_7961);
and U8266 (N_8266,N_6541,N_6545);
nor U8267 (N_8267,N_7583,N_6582);
nand U8268 (N_8268,N_6083,N_6681);
and U8269 (N_8269,N_7195,N_6446);
or U8270 (N_8270,N_6049,N_6846);
xnor U8271 (N_8271,N_6493,N_6537);
nand U8272 (N_8272,N_7559,N_6654);
nor U8273 (N_8273,N_6013,N_7647);
and U8274 (N_8274,N_7957,N_6187);
and U8275 (N_8275,N_6893,N_7392);
or U8276 (N_8276,N_6248,N_7445);
or U8277 (N_8277,N_6421,N_7476);
nand U8278 (N_8278,N_6892,N_7262);
or U8279 (N_8279,N_6784,N_7661);
nand U8280 (N_8280,N_6832,N_6371);
nand U8281 (N_8281,N_6019,N_7777);
nand U8282 (N_8282,N_6826,N_7205);
xor U8283 (N_8283,N_6620,N_7211);
nand U8284 (N_8284,N_7464,N_6132);
xor U8285 (N_8285,N_6009,N_7682);
nand U8286 (N_8286,N_6464,N_7386);
nor U8287 (N_8287,N_7196,N_7662);
or U8288 (N_8288,N_6638,N_7437);
xnor U8289 (N_8289,N_7520,N_6126);
or U8290 (N_8290,N_6676,N_7999);
or U8291 (N_8291,N_7200,N_7191);
and U8292 (N_8292,N_7857,N_7349);
or U8293 (N_8293,N_6773,N_7352);
xor U8294 (N_8294,N_7384,N_7921);
nand U8295 (N_8295,N_7923,N_7450);
or U8296 (N_8296,N_6274,N_6267);
nor U8297 (N_8297,N_7628,N_7892);
nand U8298 (N_8298,N_7054,N_7779);
nor U8299 (N_8299,N_7276,N_6482);
nand U8300 (N_8300,N_6651,N_7081);
or U8301 (N_8301,N_7704,N_6739);
xnor U8302 (N_8302,N_6199,N_6828);
xor U8303 (N_8303,N_7361,N_6761);
nor U8304 (N_8304,N_7150,N_6890);
nor U8305 (N_8305,N_7316,N_7571);
and U8306 (N_8306,N_6592,N_7758);
xnor U8307 (N_8307,N_7475,N_7942);
xor U8308 (N_8308,N_6625,N_6759);
xor U8309 (N_8309,N_7051,N_6266);
xnor U8310 (N_8310,N_7293,N_7498);
and U8311 (N_8311,N_6003,N_6134);
nand U8312 (N_8312,N_6725,N_6823);
nand U8313 (N_8313,N_6377,N_6329);
nand U8314 (N_8314,N_6525,N_6226);
nand U8315 (N_8315,N_7605,N_6491);
and U8316 (N_8316,N_6521,N_7556);
or U8317 (N_8317,N_6840,N_6624);
nand U8318 (N_8318,N_7901,N_7844);
nand U8319 (N_8319,N_7567,N_7886);
xor U8320 (N_8320,N_6240,N_7019);
nand U8321 (N_8321,N_7032,N_7617);
nor U8322 (N_8322,N_6168,N_7240);
nor U8323 (N_8323,N_7014,N_6260);
or U8324 (N_8324,N_7405,N_6445);
nor U8325 (N_8325,N_6936,N_6747);
and U8326 (N_8326,N_6970,N_7015);
nand U8327 (N_8327,N_7176,N_6577);
nor U8328 (N_8328,N_6646,N_7598);
xnor U8329 (N_8329,N_7482,N_7767);
and U8330 (N_8330,N_6279,N_6002);
nor U8331 (N_8331,N_6131,N_7097);
or U8332 (N_8332,N_6150,N_7139);
nor U8333 (N_8333,N_7795,N_6742);
and U8334 (N_8334,N_7725,N_7991);
xnor U8335 (N_8335,N_6399,N_7317);
nand U8336 (N_8336,N_7351,N_7734);
xor U8337 (N_8337,N_7971,N_7319);
nand U8338 (N_8338,N_6573,N_7757);
nand U8339 (N_8339,N_7241,N_6127);
or U8340 (N_8340,N_6022,N_6384);
xnor U8341 (N_8341,N_6477,N_6386);
xor U8342 (N_8342,N_6411,N_6919);
xnor U8343 (N_8343,N_7806,N_7720);
xor U8344 (N_8344,N_7418,N_7640);
nand U8345 (N_8345,N_6652,N_6542);
xor U8346 (N_8346,N_7034,N_6809);
and U8347 (N_8347,N_6398,N_7303);
or U8348 (N_8348,N_7016,N_7899);
or U8349 (N_8349,N_6818,N_7507);
and U8350 (N_8350,N_7544,N_7333);
xor U8351 (N_8351,N_6587,N_7410);
and U8352 (N_8352,N_7269,N_7737);
or U8353 (N_8353,N_6856,N_7540);
and U8354 (N_8354,N_6311,N_6479);
or U8355 (N_8355,N_6165,N_7554);
xor U8356 (N_8356,N_6137,N_7265);
and U8357 (N_8357,N_7120,N_7586);
and U8358 (N_8358,N_6976,N_7709);
or U8359 (N_8359,N_6028,N_7613);
nand U8360 (N_8360,N_6017,N_6979);
xnor U8361 (N_8361,N_6796,N_6595);
nand U8362 (N_8362,N_6713,N_7641);
or U8363 (N_8363,N_6331,N_6873);
or U8364 (N_8364,N_7134,N_7354);
or U8365 (N_8365,N_6942,N_7805);
nand U8366 (N_8366,N_7225,N_6007);
and U8367 (N_8367,N_6247,N_6515);
xor U8368 (N_8368,N_6552,N_6385);
nand U8369 (N_8369,N_6111,N_6677);
nor U8370 (N_8370,N_7287,N_6339);
or U8371 (N_8371,N_7318,N_7149);
and U8372 (N_8372,N_7346,N_7278);
and U8373 (N_8373,N_7622,N_6848);
nand U8374 (N_8374,N_6988,N_7634);
xor U8375 (N_8375,N_7952,N_7207);
nor U8376 (N_8376,N_6438,N_7668);
xor U8377 (N_8377,N_6813,N_6079);
nand U8378 (N_8378,N_7043,N_6327);
nor U8379 (N_8379,N_7435,N_6419);
nor U8380 (N_8380,N_6372,N_6277);
or U8381 (N_8381,N_7432,N_7888);
nor U8382 (N_8382,N_7603,N_6858);
and U8383 (N_8383,N_6871,N_7063);
nand U8384 (N_8384,N_7959,N_6310);
nand U8385 (N_8385,N_7452,N_7050);
nor U8386 (N_8386,N_7356,N_7123);
or U8387 (N_8387,N_6580,N_7024);
nand U8388 (N_8388,N_6030,N_6086);
nor U8389 (N_8389,N_6186,N_6325);
and U8390 (N_8390,N_6529,N_6080);
and U8391 (N_8391,N_7428,N_6285);
nand U8392 (N_8392,N_6935,N_7181);
nand U8393 (N_8393,N_7525,N_7029);
nor U8394 (N_8394,N_7712,N_6382);
nor U8395 (N_8395,N_6042,N_6219);
xnor U8396 (N_8396,N_7941,N_7994);
or U8397 (N_8397,N_6866,N_7242);
or U8398 (N_8398,N_7313,N_7462);
xor U8399 (N_8399,N_6814,N_6517);
xnor U8400 (N_8400,N_6188,N_7620);
nor U8401 (N_8401,N_6292,N_7408);
and U8402 (N_8402,N_7186,N_6748);
and U8403 (N_8403,N_6224,N_6869);
and U8404 (N_8404,N_6457,N_6324);
and U8405 (N_8405,N_6801,N_7052);
xor U8406 (N_8406,N_7798,N_7179);
nand U8407 (N_8407,N_7481,N_6472);
or U8408 (N_8408,N_6931,N_7810);
nand U8409 (N_8409,N_7553,N_6533);
nand U8410 (N_8410,N_7484,N_6733);
nor U8411 (N_8411,N_6644,N_7302);
nor U8412 (N_8412,N_7204,N_6901);
nand U8413 (N_8413,N_6877,N_7146);
or U8414 (N_8414,N_6543,N_6744);
nand U8415 (N_8415,N_7270,N_6963);
nand U8416 (N_8416,N_6563,N_6303);
nor U8417 (N_8417,N_6928,N_6671);
and U8418 (N_8418,N_7308,N_7380);
xor U8419 (N_8419,N_6768,N_7701);
and U8420 (N_8420,N_6147,N_7168);
nor U8421 (N_8421,N_6229,N_7789);
or U8422 (N_8422,N_7599,N_7524);
or U8423 (N_8423,N_7582,N_6182);
nand U8424 (N_8424,N_6716,N_7135);
xor U8425 (N_8425,N_6440,N_6973);
nand U8426 (N_8426,N_6430,N_7512);
xnor U8427 (N_8427,N_6291,N_6770);
nor U8428 (N_8428,N_7467,N_6647);
and U8429 (N_8429,N_7171,N_6639);
or U8430 (N_8430,N_7977,N_7255);
and U8431 (N_8431,N_6220,N_6462);
xnor U8432 (N_8432,N_6103,N_6358);
xor U8433 (N_8433,N_7296,N_6980);
xnor U8434 (N_8434,N_7561,N_6214);
nor U8435 (N_8435,N_7954,N_7088);
nor U8436 (N_8436,N_6952,N_6604);
or U8437 (N_8437,N_7080,N_7095);
nand U8438 (N_8438,N_6991,N_6530);
nand U8439 (N_8439,N_7960,N_6064);
nand U8440 (N_8440,N_6366,N_7342);
xor U8441 (N_8441,N_7162,N_6612);
xnor U8442 (N_8442,N_7746,N_6180);
or U8443 (N_8443,N_6231,N_6938);
xor U8444 (N_8444,N_6047,N_7595);
or U8445 (N_8445,N_6862,N_7696);
xnor U8446 (N_8446,N_7945,N_7290);
xnor U8447 (N_8447,N_7769,N_7830);
or U8448 (N_8448,N_6736,N_6039);
xnor U8449 (N_8449,N_7926,N_6758);
xnor U8450 (N_8450,N_6574,N_6586);
nand U8451 (N_8451,N_6395,N_6771);
nor U8452 (N_8452,N_7261,N_7334);
and U8453 (N_8453,N_6427,N_7660);
and U8454 (N_8454,N_6487,N_6707);
xor U8455 (N_8455,N_7126,N_6125);
xnor U8456 (N_8456,N_7448,N_6618);
nand U8457 (N_8457,N_6635,N_6104);
nor U8458 (N_8458,N_6157,N_7456);
nor U8459 (N_8459,N_7237,N_6363);
xor U8460 (N_8460,N_6474,N_7683);
nor U8461 (N_8461,N_7912,N_6118);
and U8462 (N_8462,N_6112,N_7616);
and U8463 (N_8463,N_7107,N_6508);
xor U8464 (N_8464,N_6743,N_6153);
nand U8465 (N_8465,N_6004,N_6560);
and U8466 (N_8466,N_7821,N_6334);
xor U8467 (N_8467,N_7028,N_6061);
xnor U8468 (N_8468,N_7320,N_6308);
nand U8469 (N_8469,N_6992,N_7880);
xor U8470 (N_8470,N_7546,N_6738);
or U8471 (N_8471,N_6196,N_7364);
and U8472 (N_8472,N_6879,N_7744);
and U8473 (N_8473,N_6172,N_7505);
nor U8474 (N_8474,N_6256,N_6576);
or U8475 (N_8475,N_6071,N_6424);
and U8476 (N_8476,N_6166,N_6227);
or U8477 (N_8477,N_6827,N_7768);
nor U8478 (N_8478,N_7564,N_6675);
and U8479 (N_8479,N_7871,N_7158);
and U8480 (N_8480,N_6340,N_6961);
nand U8481 (N_8481,N_7160,N_6968);
nand U8482 (N_8482,N_6510,N_7947);
xor U8483 (N_8483,N_6114,N_7264);
and U8484 (N_8484,N_6637,N_6522);
nor U8485 (N_8485,N_6184,N_7978);
or U8486 (N_8486,N_7982,N_6696);
and U8487 (N_8487,N_7523,N_7248);
xor U8488 (N_8488,N_6101,N_7534);
or U8489 (N_8489,N_6176,N_7238);
or U8490 (N_8490,N_7327,N_7854);
or U8491 (N_8491,N_6921,N_7529);
nor U8492 (N_8492,N_6409,N_7918);
xnor U8493 (N_8493,N_7057,N_7461);
and U8494 (N_8494,N_7778,N_7064);
and U8495 (N_8495,N_6622,N_6767);
nor U8496 (N_8496,N_7508,N_7068);
xor U8497 (N_8497,N_7000,N_6572);
or U8498 (N_8498,N_6820,N_7372);
or U8499 (N_8499,N_7053,N_6341);
nand U8500 (N_8500,N_6634,N_7309);
and U8501 (N_8501,N_7212,N_7022);
nand U8502 (N_8502,N_7688,N_7692);
and U8503 (N_8503,N_7664,N_6436);
or U8504 (N_8504,N_7913,N_7138);
and U8505 (N_8505,N_7321,N_6405);
nor U8506 (N_8506,N_6642,N_6406);
and U8507 (N_8507,N_6151,N_6420);
or U8508 (N_8508,N_6781,N_6628);
xor U8509 (N_8509,N_6496,N_6069);
or U8510 (N_8510,N_7663,N_6857);
or U8511 (N_8511,N_7974,N_7393);
or U8512 (N_8512,N_6005,N_6044);
nor U8513 (N_8513,N_6076,N_7695);
nand U8514 (N_8514,N_6884,N_6197);
xnor U8515 (N_8515,N_6362,N_7713);
xor U8516 (N_8516,N_7764,N_6908);
nand U8517 (N_8517,N_6492,N_7332);
nor U8518 (N_8518,N_6569,N_7755);
nor U8519 (N_8519,N_6805,N_6962);
xor U8520 (N_8520,N_6819,N_7409);
nor U8521 (N_8521,N_6502,N_7542);
nor U8522 (N_8522,N_6762,N_7715);
nor U8523 (N_8523,N_6727,N_6129);
xor U8524 (N_8524,N_7101,N_6376);
xor U8525 (N_8525,N_6627,N_6977);
or U8526 (N_8526,N_6706,N_6630);
xor U8527 (N_8527,N_6402,N_7851);
or U8528 (N_8528,N_6690,N_7277);
or U8529 (N_8529,N_6844,N_7938);
nor U8530 (N_8530,N_7128,N_7796);
nor U8531 (N_8531,N_6965,N_6687);
and U8532 (N_8532,N_7845,N_7807);
xor U8533 (N_8533,N_7062,N_6568);
nand U8534 (N_8534,N_6046,N_7039);
and U8535 (N_8535,N_7046,N_7765);
and U8536 (N_8536,N_7856,N_6025);
xnor U8537 (N_8537,N_6645,N_6123);
nor U8538 (N_8538,N_6000,N_7989);
nand U8539 (N_8539,N_6315,N_7483);
and U8540 (N_8540,N_6682,N_6633);
or U8541 (N_8541,N_7675,N_7565);
and U8542 (N_8542,N_6619,N_6146);
nand U8543 (N_8543,N_6729,N_6730);
or U8544 (N_8544,N_6839,N_7643);
xnor U8545 (N_8545,N_7718,N_6724);
nand U8546 (N_8546,N_7670,N_6643);
xnor U8547 (N_8547,N_7480,N_7049);
nand U8548 (N_8548,N_6524,N_6391);
xor U8549 (N_8549,N_6238,N_6357);
or U8550 (N_8550,N_7496,N_6444);
xor U8551 (N_8551,N_7263,N_6067);
xnor U8552 (N_8552,N_7917,N_7608);
nor U8553 (N_8553,N_6726,N_7853);
nand U8554 (N_8554,N_7672,N_7896);
or U8555 (N_8555,N_7180,N_6130);
nor U8556 (N_8556,N_6554,N_6722);
xor U8557 (N_8557,N_7103,N_7588);
or U8558 (N_8558,N_6189,N_6370);
nor U8559 (N_8559,N_6960,N_6008);
and U8560 (N_8560,N_7967,N_6786);
or U8561 (N_8561,N_6192,N_7474);
xor U8562 (N_8562,N_6178,N_6546);
xor U8563 (N_8563,N_7726,N_7817);
nor U8564 (N_8564,N_7315,N_7944);
nand U8565 (N_8565,N_6754,N_6615);
nor U8566 (N_8566,N_7156,N_6299);
xnor U8567 (N_8567,N_6163,N_6443);
or U8568 (N_8568,N_7882,N_6387);
and U8569 (N_8569,N_6691,N_6780);
and U8570 (N_8570,N_6997,N_7368);
xor U8571 (N_8571,N_7973,N_6865);
nor U8572 (N_8572,N_7936,N_6557);
nand U8573 (N_8573,N_7201,N_6090);
nor U8574 (N_8574,N_7449,N_7933);
and U8575 (N_8575,N_7838,N_6829);
and U8576 (N_8576,N_6653,N_7543);
and U8577 (N_8577,N_6108,N_7394);
and U8578 (N_8578,N_7828,N_7920);
and U8579 (N_8579,N_6319,N_6788);
and U8580 (N_8580,N_6463,N_6951);
nor U8581 (N_8581,N_7155,N_7092);
nor U8582 (N_8582,N_6359,N_7951);
and U8583 (N_8583,N_7714,N_7056);
or U8584 (N_8584,N_6085,N_7597);
nor U8585 (N_8585,N_6317,N_7883);
nand U8586 (N_8586,N_6778,N_7547);
nor U8587 (N_8587,N_7375,N_6250);
nor U8588 (N_8588,N_6280,N_6093);
nand U8589 (N_8589,N_6135,N_7633);
xnor U8590 (N_8590,N_7115,N_7897);
xor U8591 (N_8591,N_7385,N_7023);
xnor U8592 (N_8592,N_6629,N_7995);
nand U8593 (N_8593,N_7104,N_6688);
or U8594 (N_8594,N_7833,N_7078);
nand U8595 (N_8595,N_6987,N_7908);
or U8596 (N_8596,N_6287,N_7759);
xnor U8597 (N_8597,N_6570,N_6075);
or U8598 (N_8598,N_6202,N_6995);
nand U8599 (N_8599,N_7367,N_6711);
xnor U8600 (N_8600,N_6565,N_6695);
or U8601 (N_8601,N_7084,N_7601);
nor U8602 (N_8602,N_7119,N_7610);
or U8603 (N_8603,N_6338,N_7792);
and U8604 (N_8604,N_6024,N_7723);
xor U8605 (N_8605,N_7658,N_7964);
nor U8606 (N_8606,N_6686,N_7397);
nor U8607 (N_8607,N_6273,N_6702);
nor U8608 (N_8608,N_6205,N_6413);
xnor U8609 (N_8609,N_7510,N_7114);
and U8610 (N_8610,N_7568,N_6448);
and U8611 (N_8611,N_6225,N_6208);
nand U8612 (N_8612,N_7137,N_7167);
xnor U8613 (N_8613,N_7860,N_6837);
nand U8614 (N_8614,N_7962,N_7786);
and U8615 (N_8615,N_7850,N_6849);
nand U8616 (N_8616,N_6924,N_6321);
and U8617 (N_8617,N_7440,N_6996);
nor U8618 (N_8618,N_7673,N_7572);
xor U8619 (N_8619,N_7116,N_6081);
nand U8620 (N_8620,N_6831,N_6783);
and U8621 (N_8621,N_7089,N_6056);
and U8622 (N_8622,N_7708,N_7703);
and U8623 (N_8623,N_6887,N_7129);
or U8624 (N_8624,N_7847,N_7344);
nor U8625 (N_8625,N_7348,N_7266);
nor U8626 (N_8626,N_6850,N_7826);
nor U8627 (N_8627,N_6597,N_7602);
nor U8628 (N_8628,N_6429,N_7702);
xnor U8629 (N_8629,N_7441,N_7140);
xor U8630 (N_8630,N_7087,N_6593);
xnor U8631 (N_8631,N_7337,N_7552);
nand U8632 (N_8632,N_7206,N_7916);
and U8633 (N_8633,N_6909,N_6949);
nor U8634 (N_8634,N_6825,N_6469);
or U8635 (N_8635,N_6609,N_7190);
xor U8636 (N_8636,N_6882,N_6750);
nor U8637 (N_8637,N_6822,N_6548);
nor U8638 (N_8638,N_7310,N_6471);
nand U8639 (N_8639,N_6795,N_6442);
nand U8640 (N_8640,N_6473,N_6173);
and U8641 (N_8641,N_6703,N_7884);
or U8642 (N_8642,N_7284,N_6423);
and U8643 (N_8643,N_7898,N_7423);
or U8644 (N_8644,N_7748,N_7979);
or U8645 (N_8645,N_6252,N_7447);
nor U8646 (N_8646,N_7585,N_7222);
and U8647 (N_8647,N_6664,N_6036);
nand U8648 (N_8648,N_7533,N_7422);
nand U8649 (N_8649,N_7809,N_7326);
xnor U8650 (N_8650,N_6830,N_6660);
nor U8651 (N_8651,N_6917,N_7623);
xor U8652 (N_8652,N_7486,N_6318);
xnor U8653 (N_8653,N_7970,N_6016);
nor U8654 (N_8654,N_6870,N_7587);
or U8655 (N_8655,N_7272,N_6242);
nand U8656 (N_8656,N_6217,N_7370);
nand U8657 (N_8657,N_7800,N_7090);
xor U8658 (N_8658,N_7676,N_6947);
and U8659 (N_8659,N_6066,N_7697);
nand U8660 (N_8660,N_6116,N_6663);
nor U8661 (N_8661,N_6673,N_7112);
xnor U8662 (N_8662,N_7733,N_7044);
nor U8663 (N_8663,N_7575,N_7366);
nand U8664 (N_8664,N_6098,N_6345);
and U8665 (N_8665,N_7541,N_7932);
nor U8666 (N_8666,N_6836,N_7566);
xnor U8667 (N_8667,N_7417,N_7509);
or U8668 (N_8668,N_6284,N_7411);
nor U8669 (N_8669,N_6800,N_7373);
nand U8670 (N_8670,N_7490,N_6314);
and U8671 (N_8671,N_6301,N_6124);
nor U8672 (N_8672,N_7402,N_7988);
nand U8673 (N_8673,N_7732,N_6160);
xor U8674 (N_8674,N_7010,N_6041);
nand U8675 (N_8675,N_6181,N_6732);
nor U8676 (N_8676,N_6943,N_6710);
and U8677 (N_8677,N_7570,N_6564);
nor U8678 (N_8678,N_7984,N_7596);
nand U8679 (N_8679,N_6045,N_6434);
and U8680 (N_8680,N_6243,N_7075);
or U8681 (N_8681,N_7815,N_7842);
nand U8682 (N_8682,N_6177,N_6540);
xnor U8683 (N_8683,N_7147,N_6899);
nor U8684 (N_8684,N_7183,N_6953);
and U8685 (N_8685,N_6575,N_6278);
and U8686 (N_8686,N_6912,N_7859);
nand U8687 (N_8687,N_7956,N_7948);
nor U8688 (N_8688,N_6035,N_7458);
or U8689 (N_8689,N_6746,N_7466);
nor U8690 (N_8690,N_7001,N_7751);
xor U8691 (N_8691,N_7148,N_6259);
xor U8692 (N_8692,N_6388,N_7109);
or U8693 (N_8693,N_6600,N_7058);
nand U8694 (N_8694,N_7153,N_6966);
and U8695 (N_8695,N_7401,N_6121);
xnor U8696 (N_8696,N_7066,N_6021);
xor U8697 (N_8697,N_6367,N_6505);
or U8698 (N_8698,N_6902,N_7047);
nand U8699 (N_8699,N_6275,N_6658);
nor U8700 (N_8700,N_6404,N_7489);
nor U8701 (N_8701,N_6721,N_7604);
nand U8702 (N_8702,N_7406,N_7504);
xnor U8703 (N_8703,N_7497,N_6793);
nand U8704 (N_8704,N_7840,N_7656);
nor U8705 (N_8705,N_7192,N_7430);
xnor U8706 (N_8706,N_6333,N_6351);
nand U8707 (N_8707,N_7012,N_7125);
nand U8708 (N_8708,N_7609,N_7900);
nand U8709 (N_8709,N_7791,N_7771);
xor U8710 (N_8710,N_7535,N_7217);
xor U8711 (N_8711,N_6925,N_6981);
nand U8712 (N_8712,N_6171,N_7594);
xor U8713 (N_8713,N_6683,N_7772);
xnor U8714 (N_8714,N_6674,N_6120);
and U8715 (N_8715,N_7680,N_6060);
or U8716 (N_8716,N_6503,N_7252);
nand U8717 (N_8717,N_6957,N_6143);
nand U8718 (N_8718,N_6888,N_6095);
nor U8719 (N_8719,N_6164,N_7894);
nand U8720 (N_8720,N_7299,N_7117);
nor U8721 (N_8721,N_6361,N_7993);
or U8722 (N_8722,N_6100,N_6494);
nor U8723 (N_8723,N_6154,N_7143);
nor U8724 (N_8724,N_6602,N_7935);
and U8725 (N_8725,N_6509,N_6336);
xnor U8726 (N_8726,N_7705,N_6206);
nand U8727 (N_8727,N_7740,N_6269);
and U8728 (N_8728,N_7358,N_6559);
xnor U8729 (N_8729,N_7127,N_6944);
and U8730 (N_8730,N_6432,N_7843);
and U8731 (N_8731,N_6608,N_7420);
nor U8732 (N_8732,N_7074,N_7007);
xnor U8733 (N_8733,N_6422,N_7121);
nor U8734 (N_8734,N_6914,N_7848);
or U8735 (N_8735,N_7783,N_7468);
and U8736 (N_8736,N_7471,N_6918);
and U8737 (N_8737,N_6834,N_7152);
xor U8738 (N_8738,N_6929,N_7495);
xnor U8739 (N_8739,N_6089,N_6349);
nand U8740 (N_8740,N_6694,N_7106);
and U8741 (N_8741,N_6418,N_7745);
and U8742 (N_8742,N_7006,N_7295);
and U8743 (N_8743,N_6489,N_7584);
nand U8744 (N_8744,N_7067,N_6087);
xor U8745 (N_8745,N_6881,N_6072);
nand U8746 (N_8746,N_6531,N_7443);
and U8747 (N_8747,N_6110,N_7717);
nand U8748 (N_8748,N_6058,N_7785);
xnor U8749 (N_8749,N_7836,N_7363);
or U8750 (N_8750,N_6107,N_7627);
xor U8751 (N_8751,N_6070,N_6426);
xnor U8752 (N_8752,N_7328,N_7429);
or U8753 (N_8753,N_7407,N_6300);
or U8754 (N_8754,N_7624,N_7339);
xor U8755 (N_8755,N_7425,N_7257);
and U8756 (N_8756,N_6986,N_6596);
and U8757 (N_8757,N_6982,N_7914);
and U8758 (N_8758,N_6289,N_6328);
xor U8759 (N_8759,N_7823,N_7077);
xor U8760 (N_8760,N_7076,N_6346);
nor U8761 (N_8761,N_7790,N_7011);
and U8762 (N_8762,N_7638,N_6200);
nor U8763 (N_8763,N_6097,N_6868);
or U8764 (N_8764,N_6451,N_6763);
and U8765 (N_8765,N_6233,N_6373);
xnor U8766 (N_8766,N_6607,N_6312);
or U8767 (N_8767,N_6599,N_6649);
xnor U8768 (N_8768,N_6859,N_7280);
xnor U8769 (N_8769,N_6082,N_6145);
and U8770 (N_8770,N_7876,N_7762);
or U8771 (N_8771,N_6913,N_7799);
or U8772 (N_8772,N_7739,N_6465);
or U8773 (N_8773,N_6666,N_7335);
or U8774 (N_8774,N_6174,N_7975);
nand U8775 (N_8775,N_7072,N_6799);
nor U8776 (N_8776,N_7579,N_6769);
or U8777 (N_8777,N_7649,N_6396);
nor U8778 (N_8778,N_6497,N_6216);
xnor U8779 (N_8779,N_6360,N_7365);
nand U8780 (N_8780,N_7233,N_7347);
or U8781 (N_8781,N_6972,N_6498);
xor U8782 (N_8782,N_6985,N_7251);
nand U8783 (N_8783,N_7286,N_6414);
or U8784 (N_8784,N_7946,N_7460);
xnor U8785 (N_8785,N_6853,N_7528);
and U8786 (N_8786,N_7907,N_7215);
nor U8787 (N_8787,N_6415,N_7983);
nand U8788 (N_8788,N_7060,N_7399);
nand U8789 (N_8789,N_7998,N_7747);
and U8790 (N_8790,N_6562,N_7182);
and U8791 (N_8791,N_7210,N_7297);
xor U8792 (N_8792,N_7216,N_7172);
and U8793 (N_8793,N_7976,N_6215);
and U8794 (N_8794,N_6221,N_7825);
nand U8795 (N_8795,N_6798,N_7325);
nor U8796 (N_8796,N_7469,N_7699);
xor U8797 (N_8797,N_6712,N_7915);
xnor U8798 (N_8798,N_6109,N_7292);
and U8799 (N_8799,N_7256,N_7831);
and U8800 (N_8800,N_6662,N_7513);
nor U8801 (N_8801,N_6670,N_7170);
nand U8802 (N_8802,N_6183,N_6657);
and U8803 (N_8803,N_7390,N_6478);
or U8804 (N_8804,N_7690,N_6672);
nor U8805 (N_8805,N_7235,N_6551);
nand U8806 (N_8806,N_7743,N_7187);
or U8807 (N_8807,N_6930,N_6811);
nand U8808 (N_8808,N_7271,N_7736);
or U8809 (N_8809,N_6689,N_7177);
nor U8810 (N_8810,N_6974,N_6898);
nand U8811 (N_8811,N_7130,N_7224);
nand U8812 (N_8812,N_7657,N_7027);
nor U8813 (N_8813,N_6556,N_7997);
nand U8814 (N_8814,N_6393,N_7159);
or U8815 (N_8815,N_6640,N_7330);
nand U8816 (N_8816,N_6246,N_6092);
nor U8817 (N_8817,N_7501,N_6282);
nand U8818 (N_8818,N_6993,N_6927);
nand U8819 (N_8819,N_6598,N_7122);
nand U8820 (N_8820,N_6113,N_6990);
or U8821 (N_8821,N_6485,N_6705);
and U8822 (N_8822,N_6015,N_6156);
or U8823 (N_8823,N_7625,N_7644);
or U8824 (N_8824,N_7071,N_7530);
nor U8825 (N_8825,N_6984,N_7618);
and U8826 (N_8826,N_7436,N_7069);
or U8827 (N_8827,N_6715,N_7517);
or U8828 (N_8828,N_7037,N_6065);
xnor U8829 (N_8829,N_6040,N_7093);
or U8830 (N_8830,N_6441,N_6792);
and U8831 (N_8831,N_6428,N_7198);
and U8832 (N_8832,N_6698,N_7813);
xor U8833 (N_8833,N_7707,N_6650);
or U8834 (N_8834,N_7197,N_6601);
xor U8835 (N_8835,N_6833,N_6141);
or U8836 (N_8836,N_6669,N_6959);
or U8837 (N_8837,N_6567,N_6636);
nor U8838 (N_8838,N_6142,N_7930);
and U8839 (N_8839,N_6659,N_6885);
xnor U8840 (N_8840,N_7619,N_6519);
nor U8841 (N_8841,N_7357,N_6316);
or U8842 (N_8842,N_7578,N_7275);
nor U8843 (N_8843,N_7165,N_7005);
xor U8844 (N_8844,N_6605,N_6904);
nand U8845 (N_8845,N_7867,N_7966);
nor U8846 (N_8846,N_6106,N_6201);
xor U8847 (N_8847,N_6262,N_7359);
or U8848 (N_8848,N_6139,N_7306);
nor U8849 (N_8849,N_6875,N_7858);
nor U8850 (N_8850,N_6466,N_6449);
nor U8851 (N_8851,N_7470,N_7234);
xnor U8852 (N_8852,N_6891,N_6685);
nor U8853 (N_8853,N_7910,N_6059);
xnor U8854 (N_8854,N_6678,N_6500);
nor U8855 (N_8855,N_6526,N_6486);
and U8856 (N_8856,N_6631,N_6693);
nand U8857 (N_8857,N_7518,N_6860);
nand U8858 (N_8858,N_6480,N_6271);
or U8859 (N_8859,N_7589,N_6532);
or U8860 (N_8860,N_7350,N_7527);
xor U8861 (N_8861,N_6740,N_7574);
and U8862 (N_8862,N_6210,N_7614);
nor U8863 (N_8863,N_7463,N_6055);
nor U8864 (N_8864,N_6356,N_7877);
nand U8865 (N_8865,N_7202,N_6481);
nand U8866 (N_8866,N_6946,N_6717);
and U8867 (N_8867,N_7381,N_6755);
nor U8868 (N_8868,N_6102,N_6410);
xor U8869 (N_8869,N_7592,N_7679);
nand U8870 (N_8870,N_7031,N_7487);
xor U8871 (N_8871,N_6057,N_6534);
nor U8872 (N_8872,N_7377,N_7730);
xnor U8873 (N_8873,N_7774,N_6207);
and U8874 (N_8874,N_6379,N_7879);
nand U8875 (N_8875,N_7761,N_6513);
or U8876 (N_8876,N_7218,N_7434);
or U8877 (N_8877,N_7414,N_6872);
nand U8878 (N_8878,N_6077,N_7911);
and U8879 (N_8879,N_6133,N_7839);
or U8880 (N_8880,N_6306,N_6907);
nor U8881 (N_8881,N_6623,N_6584);
nand U8882 (N_8882,N_7820,N_7852);
nor U8883 (N_8883,N_6894,N_6149);
and U8884 (N_8884,N_6776,N_6128);
and U8885 (N_8885,N_6161,N_7722);
nand U8886 (N_8886,N_7760,N_7289);
nand U8887 (N_8887,N_6368,N_6352);
xor U8888 (N_8888,N_6236,N_6198);
nand U8889 (N_8889,N_6581,N_7009);
nand U8890 (N_8890,N_7827,N_7793);
nor U8891 (N_8891,N_6579,N_6549);
or U8892 (N_8892,N_7887,N_6488);
and U8893 (N_8893,N_7459,N_6014);
nor U8894 (N_8894,N_7873,N_7671);
and U8895 (N_8895,N_6641,N_6785);
nand U8896 (N_8896,N_7539,N_6245);
or U8897 (N_8897,N_6223,N_6905);
nor U8898 (N_8898,N_7246,N_7488);
xor U8899 (N_8899,N_7545,N_7511);
nor U8900 (N_8900,N_6012,N_7646);
or U8901 (N_8901,N_6023,N_6364);
nor U8902 (N_8902,N_7752,N_7132);
and U8903 (N_8903,N_6807,N_6922);
nor U8904 (N_8904,N_6553,N_6845);
xnor U8905 (N_8905,N_6523,N_6737);
or U8906 (N_8906,N_7360,N_7875);
or U8907 (N_8907,N_7516,N_6923);
xnor U8908 (N_8908,N_6632,N_6878);
xnor U8909 (N_8909,N_6779,N_6937);
xnor U8910 (N_8910,N_7919,N_6728);
and U8911 (N_8911,N_7274,N_6939);
and U8912 (N_8912,N_7650,N_6926);
xnor U8913 (N_8913,N_6251,N_7133);
and U8914 (N_8914,N_7950,N_6741);
or U8915 (N_8915,N_7611,N_6050);
or U8916 (N_8916,N_7629,N_7369);
nor U8917 (N_8917,N_7017,N_6499);
xnor U8918 (N_8918,N_6148,N_7788);
nand U8919 (N_8919,N_7818,N_7569);
nor U8920 (N_8920,N_7244,N_7749);
xor U8921 (N_8921,N_7314,N_6610);
nand U8922 (N_8922,N_6520,N_6751);
or U8923 (N_8923,N_6588,N_6175);
and U8924 (N_8924,N_6228,N_6096);
or U8925 (N_8925,N_7282,N_7424);
or U8926 (N_8926,N_6297,N_6948);
nor U8927 (N_8927,N_6591,N_7294);
nor U8928 (N_8928,N_7258,N_7665);
nor U8929 (N_8929,N_7781,N_7738);
nor U8930 (N_8930,N_6416,N_6626);
or U8931 (N_8931,N_7834,N_6566);
xnor U8932 (N_8932,N_6720,N_6851);
or U8933 (N_8933,N_6797,N_7403);
nand U8934 (N_8934,N_6383,N_6032);
nor U8935 (N_8935,N_6330,N_6249);
nand U8936 (N_8936,N_7061,N_7653);
xnor U8937 (N_8937,N_6027,N_6326);
or U8938 (N_8938,N_6538,N_7849);
nor U8939 (N_8939,N_7526,N_6309);
nor U8940 (N_8940,N_6874,N_6547);
or U8941 (N_8941,N_7794,N_7004);
nor U8942 (N_8942,N_6078,N_7648);
nor U8943 (N_8943,N_6700,N_7870);
nor U8944 (N_8944,N_7451,N_7766);
or U8945 (N_8945,N_6955,N_6506);
or U8946 (N_8946,N_7433,N_6989);
nand U8947 (N_8947,N_6191,N_6843);
xnor U8948 (N_8948,N_6264,N_7981);
nand U8949 (N_8949,N_7666,N_7082);
nor U8950 (N_8950,N_7909,N_6535);
or U8951 (N_8951,N_7869,N_7457);
xor U8952 (N_8952,N_7478,N_7780);
xor U8953 (N_8953,N_7889,N_7300);
nand U8954 (N_8954,N_7038,N_7144);
xnor U8955 (N_8955,N_7996,N_7336);
and U8956 (N_8956,N_7105,N_7493);
nand U8957 (N_8957,N_7455,N_6431);
xor U8958 (N_8958,N_7811,N_7581);
or U8959 (N_8959,N_6374,N_7131);
and U8960 (N_8960,N_6999,N_6468);
xnor U8961 (N_8961,N_6867,N_7891);
or U8962 (N_8962,N_6808,N_6276);
xor U8963 (N_8963,N_7026,N_6863);
and U8964 (N_8964,N_6804,N_7283);
and U8965 (N_8965,N_7969,N_7937);
nor U8966 (N_8966,N_7711,N_6998);
xor U8967 (N_8967,N_6088,N_7343);
or U8968 (N_8968,N_7267,N_6408);
nand U8969 (N_8969,N_7376,N_7922);
xor U8970 (N_8970,N_7773,N_6699);
and U8971 (N_8971,N_7558,N_6708);
nor U8972 (N_8972,N_6296,N_6261);
and U8973 (N_8973,N_7036,N_7822);
or U8974 (N_8974,N_7721,N_6789);
and U8975 (N_8975,N_7018,N_7776);
xnor U8976 (N_8976,N_7691,N_7236);
and U8977 (N_8977,N_6241,N_7866);
nor U8978 (N_8978,N_7972,N_6611);
nand U8979 (N_8979,N_6193,N_6244);
nand U8980 (N_8980,N_7002,N_7784);
and U8981 (N_8981,N_6668,N_6099);
nand U8982 (N_8982,N_6880,N_6257);
or U8983 (N_8983,N_6213,N_7754);
nand U8984 (N_8984,N_7787,N_6656);
or U8985 (N_8985,N_7415,N_6555);
xor U8986 (N_8986,N_7111,N_7301);
nor U8987 (N_8987,N_7421,N_7904);
and U8988 (N_8988,N_6470,N_6806);
and U8989 (N_8989,N_7307,N_7685);
and U8990 (N_8990,N_6772,N_7803);
xnor U8991 (N_8991,N_6234,N_6350);
nor U8992 (N_8992,N_7756,N_6590);
xnor U8993 (N_8993,N_6775,N_6369);
and U8994 (N_8994,N_7835,N_6950);
or U8995 (N_8995,N_6603,N_6764);
nand U8996 (N_8996,N_7383,N_7727);
or U8997 (N_8997,N_7804,N_6790);
xnor U8998 (N_8998,N_6916,N_7446);
nand U8999 (N_8999,N_7855,N_7863);
or U9000 (N_9000,N_7588,N_7792);
nand U9001 (N_9001,N_7951,N_6078);
and U9002 (N_9002,N_7358,N_6485);
and U9003 (N_9003,N_6496,N_7803);
xor U9004 (N_9004,N_7064,N_6759);
or U9005 (N_9005,N_6662,N_6531);
nor U9006 (N_9006,N_7986,N_7373);
or U9007 (N_9007,N_7883,N_7713);
nand U9008 (N_9008,N_6479,N_7592);
or U9009 (N_9009,N_6419,N_7992);
nor U9010 (N_9010,N_7668,N_6019);
or U9011 (N_9011,N_7837,N_7192);
nor U9012 (N_9012,N_6888,N_7760);
nor U9013 (N_9013,N_7158,N_7028);
and U9014 (N_9014,N_6420,N_6605);
nand U9015 (N_9015,N_7167,N_7876);
and U9016 (N_9016,N_6687,N_7445);
nor U9017 (N_9017,N_6328,N_7345);
nand U9018 (N_9018,N_6040,N_6374);
nor U9019 (N_9019,N_7812,N_6775);
nand U9020 (N_9020,N_6313,N_6258);
xnor U9021 (N_9021,N_7133,N_6792);
and U9022 (N_9022,N_6718,N_7477);
or U9023 (N_9023,N_6553,N_6757);
or U9024 (N_9024,N_7122,N_6459);
and U9025 (N_9025,N_6450,N_6740);
nor U9026 (N_9026,N_6667,N_6177);
and U9027 (N_9027,N_7669,N_7852);
and U9028 (N_9028,N_6524,N_6636);
or U9029 (N_9029,N_7983,N_7042);
and U9030 (N_9030,N_6729,N_6113);
nand U9031 (N_9031,N_6408,N_6748);
nand U9032 (N_9032,N_6305,N_7013);
nand U9033 (N_9033,N_6321,N_6790);
nor U9034 (N_9034,N_6077,N_6043);
and U9035 (N_9035,N_6365,N_6426);
and U9036 (N_9036,N_7307,N_6534);
and U9037 (N_9037,N_6517,N_6735);
and U9038 (N_9038,N_7363,N_6993);
xnor U9039 (N_9039,N_6430,N_6730);
nand U9040 (N_9040,N_7627,N_7621);
or U9041 (N_9041,N_7671,N_7515);
nand U9042 (N_9042,N_6579,N_6636);
and U9043 (N_9043,N_6026,N_7237);
nand U9044 (N_9044,N_6442,N_6320);
and U9045 (N_9045,N_6722,N_6343);
nor U9046 (N_9046,N_6787,N_7217);
nand U9047 (N_9047,N_6935,N_7320);
or U9048 (N_9048,N_7285,N_6378);
or U9049 (N_9049,N_6539,N_6408);
or U9050 (N_9050,N_6877,N_6450);
xnor U9051 (N_9051,N_7520,N_6426);
or U9052 (N_9052,N_6896,N_7812);
nand U9053 (N_9053,N_6166,N_6723);
nor U9054 (N_9054,N_7382,N_7600);
xor U9055 (N_9055,N_7340,N_7540);
nand U9056 (N_9056,N_7109,N_6570);
xnor U9057 (N_9057,N_6819,N_6102);
or U9058 (N_9058,N_6862,N_7674);
nor U9059 (N_9059,N_7754,N_6717);
nor U9060 (N_9060,N_6797,N_7760);
or U9061 (N_9061,N_6353,N_6255);
and U9062 (N_9062,N_7264,N_7636);
nand U9063 (N_9063,N_7367,N_6376);
or U9064 (N_9064,N_7921,N_7088);
and U9065 (N_9065,N_7301,N_6041);
or U9066 (N_9066,N_7553,N_6470);
xor U9067 (N_9067,N_6439,N_7793);
xor U9068 (N_9068,N_7120,N_6396);
xnor U9069 (N_9069,N_7661,N_6615);
nand U9070 (N_9070,N_6713,N_7833);
or U9071 (N_9071,N_7745,N_6035);
or U9072 (N_9072,N_6647,N_6050);
or U9073 (N_9073,N_7268,N_6793);
xnor U9074 (N_9074,N_6499,N_7549);
xnor U9075 (N_9075,N_7862,N_7092);
nand U9076 (N_9076,N_7938,N_7427);
nor U9077 (N_9077,N_6903,N_6347);
and U9078 (N_9078,N_6263,N_7716);
and U9079 (N_9079,N_7746,N_6619);
xor U9080 (N_9080,N_7575,N_7167);
xnor U9081 (N_9081,N_7626,N_6575);
nand U9082 (N_9082,N_7414,N_7236);
nand U9083 (N_9083,N_7179,N_6879);
or U9084 (N_9084,N_7929,N_7559);
nand U9085 (N_9085,N_6573,N_6504);
or U9086 (N_9086,N_7825,N_7022);
or U9087 (N_9087,N_6072,N_7642);
and U9088 (N_9088,N_7123,N_6169);
xnor U9089 (N_9089,N_7261,N_7893);
nand U9090 (N_9090,N_6919,N_7649);
nand U9091 (N_9091,N_7409,N_7956);
or U9092 (N_9092,N_6750,N_6151);
nor U9093 (N_9093,N_6722,N_6423);
and U9094 (N_9094,N_7164,N_6273);
and U9095 (N_9095,N_6555,N_7089);
or U9096 (N_9096,N_7694,N_7430);
or U9097 (N_9097,N_6817,N_6680);
or U9098 (N_9098,N_6531,N_6232);
nor U9099 (N_9099,N_7901,N_6333);
nor U9100 (N_9100,N_6656,N_6928);
nand U9101 (N_9101,N_7947,N_6814);
nand U9102 (N_9102,N_6105,N_6160);
nand U9103 (N_9103,N_7029,N_7893);
and U9104 (N_9104,N_7760,N_6767);
and U9105 (N_9105,N_7620,N_7680);
nor U9106 (N_9106,N_6176,N_6733);
xnor U9107 (N_9107,N_6325,N_6295);
nand U9108 (N_9108,N_6423,N_6578);
nand U9109 (N_9109,N_6066,N_6471);
xnor U9110 (N_9110,N_6916,N_7387);
or U9111 (N_9111,N_6079,N_7673);
xor U9112 (N_9112,N_6826,N_6569);
and U9113 (N_9113,N_7131,N_7871);
and U9114 (N_9114,N_7327,N_6191);
nand U9115 (N_9115,N_6999,N_7210);
nand U9116 (N_9116,N_7590,N_7495);
nor U9117 (N_9117,N_7883,N_6259);
and U9118 (N_9118,N_6982,N_6729);
xor U9119 (N_9119,N_7556,N_6216);
and U9120 (N_9120,N_7066,N_7036);
and U9121 (N_9121,N_7434,N_7579);
or U9122 (N_9122,N_6242,N_6939);
or U9123 (N_9123,N_7091,N_6043);
nand U9124 (N_9124,N_6600,N_6200);
or U9125 (N_9125,N_6083,N_7157);
xor U9126 (N_9126,N_7003,N_7817);
or U9127 (N_9127,N_6809,N_7763);
and U9128 (N_9128,N_7324,N_6890);
and U9129 (N_9129,N_7557,N_7872);
xnor U9130 (N_9130,N_6779,N_7059);
or U9131 (N_9131,N_7038,N_7135);
and U9132 (N_9132,N_6889,N_6800);
and U9133 (N_9133,N_6964,N_6887);
nor U9134 (N_9134,N_7884,N_7673);
nand U9135 (N_9135,N_6384,N_6052);
xor U9136 (N_9136,N_6144,N_6991);
nand U9137 (N_9137,N_6610,N_6802);
and U9138 (N_9138,N_6827,N_7003);
or U9139 (N_9139,N_7300,N_6448);
or U9140 (N_9140,N_6209,N_6430);
nand U9141 (N_9141,N_7884,N_7470);
nor U9142 (N_9142,N_7233,N_7037);
xnor U9143 (N_9143,N_7665,N_6968);
and U9144 (N_9144,N_7514,N_7730);
nand U9145 (N_9145,N_6849,N_6638);
and U9146 (N_9146,N_6297,N_7520);
nand U9147 (N_9147,N_7823,N_6969);
and U9148 (N_9148,N_7148,N_6079);
and U9149 (N_9149,N_6910,N_6791);
xnor U9150 (N_9150,N_7692,N_7655);
xor U9151 (N_9151,N_7059,N_7333);
xor U9152 (N_9152,N_6518,N_7748);
nand U9153 (N_9153,N_7832,N_7048);
xnor U9154 (N_9154,N_7414,N_6053);
nand U9155 (N_9155,N_6308,N_7274);
nand U9156 (N_9156,N_6302,N_6856);
nand U9157 (N_9157,N_6217,N_7323);
nor U9158 (N_9158,N_7792,N_6025);
xnor U9159 (N_9159,N_6486,N_6873);
nor U9160 (N_9160,N_7571,N_6455);
nand U9161 (N_9161,N_6075,N_7311);
nand U9162 (N_9162,N_7563,N_6868);
and U9163 (N_9163,N_6777,N_6942);
nor U9164 (N_9164,N_7715,N_7989);
or U9165 (N_9165,N_7310,N_7744);
xnor U9166 (N_9166,N_6901,N_6529);
nand U9167 (N_9167,N_6001,N_6614);
nor U9168 (N_9168,N_7035,N_7837);
or U9169 (N_9169,N_6852,N_7351);
nor U9170 (N_9170,N_7549,N_6989);
nand U9171 (N_9171,N_7387,N_7850);
and U9172 (N_9172,N_6203,N_7053);
nor U9173 (N_9173,N_6444,N_7623);
nor U9174 (N_9174,N_6850,N_7723);
nor U9175 (N_9175,N_6539,N_7871);
xor U9176 (N_9176,N_7038,N_6163);
nand U9177 (N_9177,N_7049,N_7951);
nor U9178 (N_9178,N_6336,N_6115);
nand U9179 (N_9179,N_6946,N_7823);
xnor U9180 (N_9180,N_7635,N_7025);
xnor U9181 (N_9181,N_7533,N_6145);
xnor U9182 (N_9182,N_6725,N_6722);
nand U9183 (N_9183,N_7416,N_6043);
xnor U9184 (N_9184,N_6540,N_6498);
nor U9185 (N_9185,N_7048,N_7658);
xnor U9186 (N_9186,N_6849,N_6578);
nand U9187 (N_9187,N_7047,N_6571);
nand U9188 (N_9188,N_6599,N_7380);
nor U9189 (N_9189,N_7202,N_7061);
and U9190 (N_9190,N_6544,N_6431);
and U9191 (N_9191,N_7072,N_7127);
nand U9192 (N_9192,N_7257,N_6726);
xnor U9193 (N_9193,N_6245,N_6326);
xnor U9194 (N_9194,N_7150,N_7864);
nor U9195 (N_9195,N_6967,N_6338);
and U9196 (N_9196,N_7150,N_6756);
nand U9197 (N_9197,N_7346,N_7882);
xor U9198 (N_9198,N_7245,N_7376);
or U9199 (N_9199,N_7208,N_7410);
and U9200 (N_9200,N_7700,N_6692);
nor U9201 (N_9201,N_6698,N_7844);
and U9202 (N_9202,N_6475,N_6251);
or U9203 (N_9203,N_7134,N_6904);
nand U9204 (N_9204,N_7462,N_6892);
nor U9205 (N_9205,N_6228,N_6918);
or U9206 (N_9206,N_6843,N_6366);
or U9207 (N_9207,N_6544,N_7436);
and U9208 (N_9208,N_7095,N_7982);
and U9209 (N_9209,N_6652,N_7402);
xor U9210 (N_9210,N_7514,N_6438);
xnor U9211 (N_9211,N_6076,N_6842);
nand U9212 (N_9212,N_6839,N_7176);
and U9213 (N_9213,N_7885,N_6135);
and U9214 (N_9214,N_7443,N_6913);
nand U9215 (N_9215,N_6545,N_6808);
xor U9216 (N_9216,N_7246,N_6756);
and U9217 (N_9217,N_6553,N_7617);
nor U9218 (N_9218,N_7077,N_7907);
xnor U9219 (N_9219,N_6100,N_6268);
and U9220 (N_9220,N_7448,N_6459);
or U9221 (N_9221,N_6002,N_7737);
and U9222 (N_9222,N_7999,N_7947);
nor U9223 (N_9223,N_7992,N_6354);
or U9224 (N_9224,N_7971,N_6064);
nor U9225 (N_9225,N_6621,N_7052);
and U9226 (N_9226,N_6075,N_6708);
xnor U9227 (N_9227,N_7497,N_6227);
and U9228 (N_9228,N_6163,N_7536);
xnor U9229 (N_9229,N_7823,N_7621);
and U9230 (N_9230,N_7259,N_7302);
nand U9231 (N_9231,N_7634,N_7760);
nand U9232 (N_9232,N_6083,N_6903);
nand U9233 (N_9233,N_7275,N_6090);
and U9234 (N_9234,N_7378,N_7662);
or U9235 (N_9235,N_7018,N_6637);
or U9236 (N_9236,N_6114,N_7786);
xor U9237 (N_9237,N_6906,N_6212);
nand U9238 (N_9238,N_7407,N_7093);
or U9239 (N_9239,N_6687,N_7230);
nor U9240 (N_9240,N_7177,N_6311);
xnor U9241 (N_9241,N_7610,N_7190);
or U9242 (N_9242,N_6416,N_6653);
and U9243 (N_9243,N_7027,N_6023);
nor U9244 (N_9244,N_7484,N_6640);
and U9245 (N_9245,N_6317,N_7684);
nor U9246 (N_9246,N_7679,N_7882);
or U9247 (N_9247,N_6246,N_7974);
nor U9248 (N_9248,N_7383,N_7828);
or U9249 (N_9249,N_7114,N_7346);
or U9250 (N_9250,N_6758,N_7913);
xor U9251 (N_9251,N_6232,N_6293);
nand U9252 (N_9252,N_7072,N_7844);
nor U9253 (N_9253,N_6416,N_6707);
xor U9254 (N_9254,N_7262,N_6646);
and U9255 (N_9255,N_7099,N_6357);
or U9256 (N_9256,N_7221,N_6357);
nor U9257 (N_9257,N_6596,N_6706);
nor U9258 (N_9258,N_7565,N_7480);
or U9259 (N_9259,N_7814,N_7959);
nand U9260 (N_9260,N_7943,N_7652);
xor U9261 (N_9261,N_7317,N_6668);
nand U9262 (N_9262,N_6312,N_6023);
nor U9263 (N_9263,N_6447,N_7226);
and U9264 (N_9264,N_7502,N_7620);
or U9265 (N_9265,N_7432,N_7050);
and U9266 (N_9266,N_6958,N_7115);
nand U9267 (N_9267,N_6808,N_6063);
nor U9268 (N_9268,N_7384,N_6556);
nand U9269 (N_9269,N_7514,N_7525);
and U9270 (N_9270,N_7243,N_7730);
nand U9271 (N_9271,N_7994,N_6909);
nand U9272 (N_9272,N_7566,N_6339);
nand U9273 (N_9273,N_6459,N_7743);
nor U9274 (N_9274,N_6550,N_7619);
nand U9275 (N_9275,N_6188,N_6787);
nand U9276 (N_9276,N_6997,N_7893);
xor U9277 (N_9277,N_7078,N_7800);
nand U9278 (N_9278,N_6483,N_7410);
nand U9279 (N_9279,N_7427,N_6013);
xnor U9280 (N_9280,N_6305,N_6523);
or U9281 (N_9281,N_6301,N_7382);
xnor U9282 (N_9282,N_7609,N_7183);
xor U9283 (N_9283,N_6628,N_7938);
nor U9284 (N_9284,N_6081,N_6925);
xor U9285 (N_9285,N_6144,N_6676);
nor U9286 (N_9286,N_6094,N_6468);
and U9287 (N_9287,N_6977,N_6898);
and U9288 (N_9288,N_7589,N_7406);
nor U9289 (N_9289,N_7217,N_7092);
nand U9290 (N_9290,N_6254,N_6859);
nor U9291 (N_9291,N_6229,N_6224);
and U9292 (N_9292,N_7252,N_7569);
and U9293 (N_9293,N_6360,N_7283);
or U9294 (N_9294,N_6360,N_7066);
and U9295 (N_9295,N_7234,N_7469);
nor U9296 (N_9296,N_6462,N_7707);
nand U9297 (N_9297,N_7519,N_6501);
nand U9298 (N_9298,N_7125,N_6787);
or U9299 (N_9299,N_6320,N_7517);
or U9300 (N_9300,N_7485,N_6278);
nand U9301 (N_9301,N_6159,N_6082);
nand U9302 (N_9302,N_7728,N_6454);
nor U9303 (N_9303,N_7415,N_7566);
xnor U9304 (N_9304,N_6851,N_6879);
xnor U9305 (N_9305,N_6285,N_7784);
or U9306 (N_9306,N_7551,N_7601);
nor U9307 (N_9307,N_7635,N_7902);
xor U9308 (N_9308,N_7354,N_7361);
or U9309 (N_9309,N_6677,N_6819);
and U9310 (N_9310,N_6108,N_7164);
nand U9311 (N_9311,N_6346,N_7557);
xnor U9312 (N_9312,N_7902,N_7354);
nand U9313 (N_9313,N_7260,N_6980);
and U9314 (N_9314,N_7204,N_6467);
xnor U9315 (N_9315,N_7983,N_7227);
xnor U9316 (N_9316,N_6038,N_7562);
and U9317 (N_9317,N_7515,N_7146);
nor U9318 (N_9318,N_6191,N_7982);
nor U9319 (N_9319,N_6709,N_6787);
or U9320 (N_9320,N_6294,N_7496);
or U9321 (N_9321,N_6368,N_6026);
xor U9322 (N_9322,N_6952,N_6995);
nand U9323 (N_9323,N_6806,N_6746);
and U9324 (N_9324,N_7474,N_6409);
and U9325 (N_9325,N_6745,N_7281);
xor U9326 (N_9326,N_7807,N_6597);
or U9327 (N_9327,N_6569,N_6181);
xor U9328 (N_9328,N_7575,N_6960);
and U9329 (N_9329,N_6760,N_7468);
xor U9330 (N_9330,N_6699,N_7480);
or U9331 (N_9331,N_6542,N_7896);
or U9332 (N_9332,N_6312,N_7766);
nor U9333 (N_9333,N_7357,N_6365);
and U9334 (N_9334,N_7018,N_6464);
and U9335 (N_9335,N_6920,N_6976);
xnor U9336 (N_9336,N_6154,N_6028);
xnor U9337 (N_9337,N_6609,N_7226);
or U9338 (N_9338,N_7914,N_7502);
and U9339 (N_9339,N_7409,N_7771);
or U9340 (N_9340,N_7882,N_6169);
xnor U9341 (N_9341,N_6764,N_6087);
or U9342 (N_9342,N_7330,N_7836);
nor U9343 (N_9343,N_7399,N_6280);
xnor U9344 (N_9344,N_7306,N_7842);
xnor U9345 (N_9345,N_6287,N_6744);
or U9346 (N_9346,N_6860,N_7274);
or U9347 (N_9347,N_6415,N_6100);
nand U9348 (N_9348,N_7068,N_6322);
nor U9349 (N_9349,N_7949,N_7035);
or U9350 (N_9350,N_6453,N_7873);
xnor U9351 (N_9351,N_6586,N_6723);
nand U9352 (N_9352,N_7059,N_6961);
and U9353 (N_9353,N_7781,N_6736);
and U9354 (N_9354,N_7077,N_7889);
or U9355 (N_9355,N_7302,N_7141);
xor U9356 (N_9356,N_7827,N_7055);
nor U9357 (N_9357,N_7736,N_6616);
nor U9358 (N_9358,N_7458,N_6100);
nand U9359 (N_9359,N_7717,N_7671);
or U9360 (N_9360,N_7244,N_7282);
xnor U9361 (N_9361,N_7589,N_7291);
or U9362 (N_9362,N_6880,N_7672);
xor U9363 (N_9363,N_7615,N_6751);
or U9364 (N_9364,N_7772,N_6458);
xor U9365 (N_9365,N_7099,N_6325);
nor U9366 (N_9366,N_7854,N_6188);
xnor U9367 (N_9367,N_7143,N_6243);
xnor U9368 (N_9368,N_7784,N_7891);
nor U9369 (N_9369,N_6311,N_7897);
nand U9370 (N_9370,N_7386,N_7393);
and U9371 (N_9371,N_6085,N_6609);
nor U9372 (N_9372,N_7633,N_6268);
nor U9373 (N_9373,N_7853,N_7742);
xnor U9374 (N_9374,N_6548,N_7282);
or U9375 (N_9375,N_7182,N_6481);
nand U9376 (N_9376,N_6957,N_6471);
nor U9377 (N_9377,N_6055,N_6429);
or U9378 (N_9378,N_7994,N_7380);
and U9379 (N_9379,N_6047,N_7111);
and U9380 (N_9380,N_7769,N_7527);
or U9381 (N_9381,N_6580,N_6745);
nand U9382 (N_9382,N_6830,N_6701);
nand U9383 (N_9383,N_7648,N_6766);
nand U9384 (N_9384,N_6929,N_6275);
and U9385 (N_9385,N_6145,N_7124);
nand U9386 (N_9386,N_6444,N_6638);
xnor U9387 (N_9387,N_7160,N_7182);
xnor U9388 (N_9388,N_6546,N_6239);
nor U9389 (N_9389,N_6094,N_6258);
and U9390 (N_9390,N_7513,N_6846);
nor U9391 (N_9391,N_6433,N_6962);
and U9392 (N_9392,N_7047,N_6421);
xor U9393 (N_9393,N_6930,N_7311);
xor U9394 (N_9394,N_6843,N_7054);
and U9395 (N_9395,N_6647,N_7261);
nand U9396 (N_9396,N_7962,N_7552);
or U9397 (N_9397,N_6113,N_6956);
xor U9398 (N_9398,N_6352,N_7337);
xnor U9399 (N_9399,N_7106,N_6760);
nor U9400 (N_9400,N_6962,N_7039);
xor U9401 (N_9401,N_7966,N_6167);
and U9402 (N_9402,N_6678,N_7834);
nand U9403 (N_9403,N_6294,N_7668);
xnor U9404 (N_9404,N_7316,N_7330);
nor U9405 (N_9405,N_6100,N_6361);
and U9406 (N_9406,N_7247,N_7767);
nor U9407 (N_9407,N_7959,N_7612);
or U9408 (N_9408,N_7154,N_7561);
nor U9409 (N_9409,N_6463,N_6804);
xor U9410 (N_9410,N_6604,N_7490);
nor U9411 (N_9411,N_6284,N_6632);
nor U9412 (N_9412,N_7004,N_7841);
nand U9413 (N_9413,N_7623,N_6469);
nor U9414 (N_9414,N_7877,N_7298);
nand U9415 (N_9415,N_6186,N_7242);
nor U9416 (N_9416,N_6742,N_6284);
xnor U9417 (N_9417,N_6162,N_6672);
xor U9418 (N_9418,N_6517,N_7771);
and U9419 (N_9419,N_6665,N_7350);
or U9420 (N_9420,N_6730,N_7641);
nand U9421 (N_9421,N_6186,N_6390);
nand U9422 (N_9422,N_6892,N_6299);
nor U9423 (N_9423,N_7885,N_6436);
xor U9424 (N_9424,N_7070,N_6021);
nand U9425 (N_9425,N_6215,N_6124);
nor U9426 (N_9426,N_7741,N_6382);
or U9427 (N_9427,N_6121,N_7871);
xor U9428 (N_9428,N_7200,N_6167);
xnor U9429 (N_9429,N_6056,N_6799);
and U9430 (N_9430,N_6120,N_6228);
nor U9431 (N_9431,N_7473,N_7133);
nand U9432 (N_9432,N_6132,N_6952);
xnor U9433 (N_9433,N_6989,N_7872);
and U9434 (N_9434,N_7415,N_6778);
or U9435 (N_9435,N_6727,N_6438);
nor U9436 (N_9436,N_6010,N_6239);
and U9437 (N_9437,N_6326,N_6491);
nor U9438 (N_9438,N_6130,N_7002);
and U9439 (N_9439,N_7462,N_6687);
or U9440 (N_9440,N_6066,N_7822);
and U9441 (N_9441,N_6200,N_7405);
or U9442 (N_9442,N_6515,N_7131);
xnor U9443 (N_9443,N_7547,N_7046);
xor U9444 (N_9444,N_6588,N_6561);
and U9445 (N_9445,N_7486,N_7606);
and U9446 (N_9446,N_6321,N_7685);
xor U9447 (N_9447,N_7329,N_6322);
nor U9448 (N_9448,N_7548,N_6787);
xor U9449 (N_9449,N_7620,N_6545);
or U9450 (N_9450,N_7414,N_7336);
nor U9451 (N_9451,N_7575,N_7423);
and U9452 (N_9452,N_6345,N_7222);
or U9453 (N_9453,N_7305,N_7406);
and U9454 (N_9454,N_7213,N_7173);
nand U9455 (N_9455,N_7472,N_6099);
or U9456 (N_9456,N_7979,N_6312);
or U9457 (N_9457,N_7127,N_7913);
and U9458 (N_9458,N_7369,N_7432);
or U9459 (N_9459,N_6632,N_7398);
or U9460 (N_9460,N_7130,N_7795);
xnor U9461 (N_9461,N_6842,N_7000);
nand U9462 (N_9462,N_7373,N_7729);
nor U9463 (N_9463,N_6985,N_6396);
or U9464 (N_9464,N_7070,N_6262);
nand U9465 (N_9465,N_6972,N_7123);
nor U9466 (N_9466,N_6181,N_6474);
or U9467 (N_9467,N_7517,N_6511);
and U9468 (N_9468,N_7306,N_7653);
or U9469 (N_9469,N_6645,N_7516);
nor U9470 (N_9470,N_7771,N_7147);
and U9471 (N_9471,N_6345,N_6352);
xnor U9472 (N_9472,N_6527,N_7435);
or U9473 (N_9473,N_6629,N_6992);
nand U9474 (N_9474,N_6439,N_7056);
nor U9475 (N_9475,N_7772,N_7167);
or U9476 (N_9476,N_6296,N_6295);
xor U9477 (N_9477,N_6328,N_7173);
xor U9478 (N_9478,N_6172,N_6541);
nand U9479 (N_9479,N_6645,N_6654);
and U9480 (N_9480,N_6472,N_6092);
nor U9481 (N_9481,N_7888,N_7974);
nand U9482 (N_9482,N_6656,N_6955);
nand U9483 (N_9483,N_6409,N_6332);
and U9484 (N_9484,N_7432,N_6139);
xor U9485 (N_9485,N_7517,N_7182);
xor U9486 (N_9486,N_7430,N_7529);
and U9487 (N_9487,N_7665,N_6044);
nor U9488 (N_9488,N_7557,N_6928);
nor U9489 (N_9489,N_7333,N_6944);
xnor U9490 (N_9490,N_6783,N_6564);
nor U9491 (N_9491,N_6394,N_7680);
or U9492 (N_9492,N_7867,N_6904);
nor U9493 (N_9493,N_6128,N_6221);
and U9494 (N_9494,N_7126,N_6934);
nor U9495 (N_9495,N_6361,N_6820);
xor U9496 (N_9496,N_7705,N_7117);
nand U9497 (N_9497,N_6740,N_7913);
nand U9498 (N_9498,N_6184,N_7383);
nand U9499 (N_9499,N_6713,N_6520);
nand U9500 (N_9500,N_6533,N_7063);
or U9501 (N_9501,N_7187,N_6629);
nand U9502 (N_9502,N_7145,N_7316);
nor U9503 (N_9503,N_6594,N_6322);
or U9504 (N_9504,N_6200,N_7511);
nor U9505 (N_9505,N_7359,N_6209);
and U9506 (N_9506,N_7522,N_6010);
nand U9507 (N_9507,N_6007,N_6323);
nor U9508 (N_9508,N_6836,N_6544);
or U9509 (N_9509,N_6977,N_7092);
and U9510 (N_9510,N_7583,N_7157);
and U9511 (N_9511,N_7963,N_7396);
nand U9512 (N_9512,N_7305,N_6121);
nand U9513 (N_9513,N_7946,N_6826);
and U9514 (N_9514,N_7634,N_6707);
xor U9515 (N_9515,N_7588,N_7168);
nor U9516 (N_9516,N_6653,N_6467);
and U9517 (N_9517,N_7420,N_7130);
nand U9518 (N_9518,N_7783,N_6721);
nand U9519 (N_9519,N_6556,N_7475);
nor U9520 (N_9520,N_7909,N_7008);
nor U9521 (N_9521,N_6510,N_7232);
nor U9522 (N_9522,N_7878,N_6117);
nor U9523 (N_9523,N_6937,N_6980);
or U9524 (N_9524,N_7313,N_6761);
and U9525 (N_9525,N_7656,N_6147);
or U9526 (N_9526,N_7782,N_6765);
and U9527 (N_9527,N_6085,N_7819);
nand U9528 (N_9528,N_6634,N_6830);
xnor U9529 (N_9529,N_6302,N_6674);
nor U9530 (N_9530,N_7300,N_6065);
or U9531 (N_9531,N_6796,N_6912);
or U9532 (N_9532,N_6138,N_6655);
xnor U9533 (N_9533,N_6108,N_7578);
xnor U9534 (N_9534,N_6165,N_7180);
and U9535 (N_9535,N_6353,N_7991);
nor U9536 (N_9536,N_7308,N_7572);
or U9537 (N_9537,N_6659,N_7143);
nand U9538 (N_9538,N_6143,N_6724);
nand U9539 (N_9539,N_7620,N_7535);
and U9540 (N_9540,N_6558,N_6985);
nand U9541 (N_9541,N_6429,N_7473);
nor U9542 (N_9542,N_6037,N_7245);
and U9543 (N_9543,N_6500,N_7568);
nor U9544 (N_9544,N_6058,N_6629);
nand U9545 (N_9545,N_7546,N_6741);
xnor U9546 (N_9546,N_7178,N_6384);
or U9547 (N_9547,N_6568,N_6997);
and U9548 (N_9548,N_7658,N_6859);
nor U9549 (N_9549,N_7676,N_7531);
or U9550 (N_9550,N_7782,N_7199);
and U9551 (N_9551,N_7630,N_7887);
and U9552 (N_9552,N_6319,N_7217);
or U9553 (N_9553,N_6224,N_6968);
nand U9554 (N_9554,N_6151,N_6964);
nor U9555 (N_9555,N_6637,N_6902);
nor U9556 (N_9556,N_6146,N_6676);
and U9557 (N_9557,N_6278,N_7688);
nor U9558 (N_9558,N_7467,N_6726);
nand U9559 (N_9559,N_6454,N_7336);
nand U9560 (N_9560,N_7491,N_7206);
nand U9561 (N_9561,N_6027,N_7466);
or U9562 (N_9562,N_7039,N_6887);
nand U9563 (N_9563,N_7443,N_6737);
and U9564 (N_9564,N_7416,N_6097);
nand U9565 (N_9565,N_7172,N_6810);
nor U9566 (N_9566,N_6630,N_7094);
nor U9567 (N_9567,N_6181,N_6477);
nand U9568 (N_9568,N_7358,N_6240);
or U9569 (N_9569,N_6031,N_6834);
nand U9570 (N_9570,N_6441,N_7322);
nor U9571 (N_9571,N_6369,N_7293);
or U9572 (N_9572,N_7193,N_6879);
nor U9573 (N_9573,N_7410,N_7853);
or U9574 (N_9574,N_6820,N_6011);
nand U9575 (N_9575,N_6941,N_6963);
nor U9576 (N_9576,N_6984,N_7619);
or U9577 (N_9577,N_6270,N_6390);
and U9578 (N_9578,N_6732,N_7634);
and U9579 (N_9579,N_6458,N_6809);
or U9580 (N_9580,N_7326,N_7990);
or U9581 (N_9581,N_7131,N_7972);
nor U9582 (N_9582,N_6219,N_7292);
or U9583 (N_9583,N_6622,N_7623);
nor U9584 (N_9584,N_6255,N_6302);
nor U9585 (N_9585,N_7388,N_6034);
nand U9586 (N_9586,N_7606,N_6726);
xor U9587 (N_9587,N_6952,N_6756);
xnor U9588 (N_9588,N_6279,N_6541);
nor U9589 (N_9589,N_6364,N_7055);
nand U9590 (N_9590,N_7108,N_6713);
nor U9591 (N_9591,N_6943,N_7822);
nor U9592 (N_9592,N_6458,N_7209);
nand U9593 (N_9593,N_6608,N_6332);
nand U9594 (N_9594,N_7408,N_7108);
xor U9595 (N_9595,N_6494,N_7879);
and U9596 (N_9596,N_7449,N_6666);
xnor U9597 (N_9597,N_6895,N_6650);
and U9598 (N_9598,N_6978,N_6491);
nand U9599 (N_9599,N_7815,N_7145);
xnor U9600 (N_9600,N_6494,N_6912);
nand U9601 (N_9601,N_6831,N_6414);
nor U9602 (N_9602,N_6048,N_7263);
and U9603 (N_9603,N_7879,N_6286);
nor U9604 (N_9604,N_7926,N_7277);
nor U9605 (N_9605,N_6853,N_6710);
nand U9606 (N_9606,N_6193,N_7611);
xor U9607 (N_9607,N_7972,N_7494);
nand U9608 (N_9608,N_7222,N_7053);
xnor U9609 (N_9609,N_7415,N_7085);
nand U9610 (N_9610,N_6960,N_6849);
xor U9611 (N_9611,N_7226,N_7250);
nand U9612 (N_9612,N_7461,N_7484);
or U9613 (N_9613,N_6748,N_6450);
nor U9614 (N_9614,N_6071,N_7901);
and U9615 (N_9615,N_6016,N_6487);
nor U9616 (N_9616,N_6564,N_6604);
nand U9617 (N_9617,N_7617,N_7198);
nor U9618 (N_9618,N_7779,N_6718);
and U9619 (N_9619,N_6899,N_7258);
and U9620 (N_9620,N_7715,N_7113);
xor U9621 (N_9621,N_7551,N_6993);
or U9622 (N_9622,N_7932,N_7258);
nor U9623 (N_9623,N_6183,N_6379);
nor U9624 (N_9624,N_6546,N_7183);
and U9625 (N_9625,N_7467,N_7381);
nand U9626 (N_9626,N_7559,N_7417);
and U9627 (N_9627,N_7692,N_6817);
or U9628 (N_9628,N_6396,N_7114);
or U9629 (N_9629,N_6891,N_7438);
and U9630 (N_9630,N_6592,N_6681);
and U9631 (N_9631,N_6319,N_7357);
nor U9632 (N_9632,N_7806,N_7919);
xnor U9633 (N_9633,N_6736,N_6587);
and U9634 (N_9634,N_7415,N_7287);
or U9635 (N_9635,N_6978,N_7380);
and U9636 (N_9636,N_7206,N_7485);
nor U9637 (N_9637,N_7452,N_7527);
or U9638 (N_9638,N_7719,N_7955);
nand U9639 (N_9639,N_7686,N_7723);
or U9640 (N_9640,N_7269,N_7796);
and U9641 (N_9641,N_6759,N_7778);
and U9642 (N_9642,N_6445,N_6227);
and U9643 (N_9643,N_6798,N_6606);
nor U9644 (N_9644,N_7939,N_7351);
or U9645 (N_9645,N_7972,N_7097);
xor U9646 (N_9646,N_7149,N_6920);
or U9647 (N_9647,N_6695,N_7078);
xnor U9648 (N_9648,N_6166,N_7475);
and U9649 (N_9649,N_7395,N_7709);
or U9650 (N_9650,N_6667,N_6091);
nand U9651 (N_9651,N_6560,N_6566);
nor U9652 (N_9652,N_7034,N_6106);
and U9653 (N_9653,N_7500,N_7153);
nor U9654 (N_9654,N_7772,N_7435);
and U9655 (N_9655,N_6002,N_6612);
or U9656 (N_9656,N_7359,N_6308);
nor U9657 (N_9657,N_7260,N_7140);
nor U9658 (N_9658,N_7627,N_7120);
or U9659 (N_9659,N_6199,N_7728);
nand U9660 (N_9660,N_7482,N_6324);
nand U9661 (N_9661,N_6950,N_7853);
or U9662 (N_9662,N_7887,N_7272);
or U9663 (N_9663,N_7023,N_7015);
nor U9664 (N_9664,N_6617,N_7792);
nand U9665 (N_9665,N_6162,N_6630);
nor U9666 (N_9666,N_6303,N_6578);
or U9667 (N_9667,N_6792,N_6382);
or U9668 (N_9668,N_6477,N_6694);
nand U9669 (N_9669,N_6050,N_7981);
or U9670 (N_9670,N_6540,N_6338);
nor U9671 (N_9671,N_7951,N_6864);
xor U9672 (N_9672,N_6653,N_6620);
and U9673 (N_9673,N_6211,N_6435);
nor U9674 (N_9674,N_7182,N_7957);
and U9675 (N_9675,N_6352,N_7946);
and U9676 (N_9676,N_6490,N_6116);
nor U9677 (N_9677,N_7578,N_6519);
and U9678 (N_9678,N_6528,N_6449);
nor U9679 (N_9679,N_7196,N_7143);
or U9680 (N_9680,N_7732,N_7961);
nor U9681 (N_9681,N_7246,N_6478);
xnor U9682 (N_9682,N_6101,N_7577);
or U9683 (N_9683,N_7765,N_7154);
or U9684 (N_9684,N_7382,N_7724);
xor U9685 (N_9685,N_6345,N_6210);
xnor U9686 (N_9686,N_6533,N_7993);
or U9687 (N_9687,N_6726,N_7315);
xor U9688 (N_9688,N_7104,N_7480);
xnor U9689 (N_9689,N_7076,N_7113);
and U9690 (N_9690,N_6622,N_6427);
and U9691 (N_9691,N_6029,N_7806);
nand U9692 (N_9692,N_6446,N_7441);
or U9693 (N_9693,N_6844,N_7264);
or U9694 (N_9694,N_7580,N_6753);
and U9695 (N_9695,N_6133,N_6925);
or U9696 (N_9696,N_7927,N_7487);
xor U9697 (N_9697,N_7741,N_6969);
and U9698 (N_9698,N_7847,N_6672);
nand U9699 (N_9699,N_7798,N_6160);
xnor U9700 (N_9700,N_7477,N_6007);
or U9701 (N_9701,N_7620,N_7840);
nand U9702 (N_9702,N_6644,N_7867);
nor U9703 (N_9703,N_6109,N_6954);
or U9704 (N_9704,N_6734,N_7468);
and U9705 (N_9705,N_6454,N_6033);
nand U9706 (N_9706,N_6164,N_7676);
nor U9707 (N_9707,N_7407,N_7028);
and U9708 (N_9708,N_6714,N_7665);
nand U9709 (N_9709,N_6934,N_6340);
xor U9710 (N_9710,N_6059,N_6860);
nand U9711 (N_9711,N_6065,N_6932);
or U9712 (N_9712,N_7997,N_6388);
xnor U9713 (N_9713,N_7547,N_7886);
xor U9714 (N_9714,N_7315,N_7219);
nand U9715 (N_9715,N_7112,N_7638);
xnor U9716 (N_9716,N_7370,N_7273);
or U9717 (N_9717,N_6295,N_6116);
or U9718 (N_9718,N_7797,N_7762);
nor U9719 (N_9719,N_6278,N_6049);
nor U9720 (N_9720,N_7648,N_6322);
and U9721 (N_9721,N_7016,N_7850);
or U9722 (N_9722,N_6225,N_7389);
nand U9723 (N_9723,N_7644,N_7807);
or U9724 (N_9724,N_7371,N_7675);
or U9725 (N_9725,N_7471,N_6837);
and U9726 (N_9726,N_7349,N_7135);
or U9727 (N_9727,N_6569,N_7514);
and U9728 (N_9728,N_7883,N_6116);
nor U9729 (N_9729,N_7491,N_7443);
or U9730 (N_9730,N_6922,N_6706);
and U9731 (N_9731,N_7869,N_7262);
nor U9732 (N_9732,N_6867,N_7885);
nand U9733 (N_9733,N_6075,N_6325);
nor U9734 (N_9734,N_7934,N_6239);
xor U9735 (N_9735,N_6893,N_6871);
nand U9736 (N_9736,N_7665,N_7075);
and U9737 (N_9737,N_7172,N_6175);
nor U9738 (N_9738,N_7781,N_7580);
xnor U9739 (N_9739,N_7069,N_7895);
nor U9740 (N_9740,N_6026,N_7719);
and U9741 (N_9741,N_6121,N_6963);
and U9742 (N_9742,N_7847,N_7442);
or U9743 (N_9743,N_7908,N_7609);
nand U9744 (N_9744,N_7741,N_6013);
nor U9745 (N_9745,N_6099,N_7009);
or U9746 (N_9746,N_6748,N_7502);
nor U9747 (N_9747,N_7577,N_6413);
xor U9748 (N_9748,N_7066,N_6485);
or U9749 (N_9749,N_7421,N_7039);
nor U9750 (N_9750,N_6860,N_7979);
nor U9751 (N_9751,N_6148,N_7930);
xnor U9752 (N_9752,N_7831,N_7155);
and U9753 (N_9753,N_7597,N_7115);
nand U9754 (N_9754,N_7611,N_6741);
xor U9755 (N_9755,N_7555,N_7955);
nand U9756 (N_9756,N_6094,N_7118);
xnor U9757 (N_9757,N_6367,N_6495);
or U9758 (N_9758,N_7595,N_7172);
nor U9759 (N_9759,N_7175,N_6767);
nand U9760 (N_9760,N_7950,N_7264);
nor U9761 (N_9761,N_6154,N_6235);
nor U9762 (N_9762,N_7052,N_7231);
nand U9763 (N_9763,N_7247,N_7539);
and U9764 (N_9764,N_7258,N_6049);
nor U9765 (N_9765,N_7204,N_7582);
xnor U9766 (N_9766,N_6475,N_7444);
nor U9767 (N_9767,N_7119,N_7020);
or U9768 (N_9768,N_7186,N_6137);
and U9769 (N_9769,N_7601,N_6275);
and U9770 (N_9770,N_7497,N_6570);
xnor U9771 (N_9771,N_7438,N_6948);
nand U9772 (N_9772,N_7679,N_7906);
nand U9773 (N_9773,N_7289,N_7785);
or U9774 (N_9774,N_6654,N_6284);
nor U9775 (N_9775,N_7997,N_6050);
nor U9776 (N_9776,N_7271,N_6170);
xor U9777 (N_9777,N_6410,N_6392);
and U9778 (N_9778,N_7337,N_6796);
nor U9779 (N_9779,N_7979,N_7493);
nand U9780 (N_9780,N_7411,N_7508);
xnor U9781 (N_9781,N_7667,N_6951);
or U9782 (N_9782,N_6779,N_6940);
xnor U9783 (N_9783,N_6971,N_6192);
and U9784 (N_9784,N_7761,N_7610);
nand U9785 (N_9785,N_6170,N_6204);
nor U9786 (N_9786,N_6255,N_7709);
and U9787 (N_9787,N_7461,N_6551);
or U9788 (N_9788,N_6933,N_6790);
nor U9789 (N_9789,N_6855,N_7248);
nor U9790 (N_9790,N_6577,N_7989);
and U9791 (N_9791,N_7241,N_6638);
and U9792 (N_9792,N_7732,N_7108);
or U9793 (N_9793,N_6656,N_6016);
nor U9794 (N_9794,N_7521,N_7438);
xnor U9795 (N_9795,N_7402,N_6412);
nor U9796 (N_9796,N_7929,N_7855);
xnor U9797 (N_9797,N_7447,N_7569);
or U9798 (N_9798,N_7145,N_6464);
xnor U9799 (N_9799,N_7615,N_6750);
nand U9800 (N_9800,N_6300,N_7964);
nor U9801 (N_9801,N_7288,N_7406);
nand U9802 (N_9802,N_7812,N_7045);
nand U9803 (N_9803,N_7460,N_6923);
nand U9804 (N_9804,N_7704,N_6579);
nor U9805 (N_9805,N_7220,N_6241);
or U9806 (N_9806,N_7168,N_7229);
and U9807 (N_9807,N_7372,N_6840);
xor U9808 (N_9808,N_6762,N_7227);
nand U9809 (N_9809,N_6834,N_6060);
nor U9810 (N_9810,N_6932,N_6210);
xor U9811 (N_9811,N_6510,N_6650);
and U9812 (N_9812,N_7123,N_6503);
or U9813 (N_9813,N_7574,N_7186);
nand U9814 (N_9814,N_6913,N_6917);
nand U9815 (N_9815,N_7607,N_7365);
nand U9816 (N_9816,N_6218,N_6369);
and U9817 (N_9817,N_6441,N_7628);
nor U9818 (N_9818,N_6350,N_6808);
or U9819 (N_9819,N_7504,N_6874);
and U9820 (N_9820,N_6390,N_7092);
xnor U9821 (N_9821,N_6730,N_6887);
xor U9822 (N_9822,N_6142,N_6869);
and U9823 (N_9823,N_6932,N_7483);
or U9824 (N_9824,N_6572,N_7427);
or U9825 (N_9825,N_6199,N_7027);
and U9826 (N_9826,N_6433,N_6746);
and U9827 (N_9827,N_7754,N_6414);
nand U9828 (N_9828,N_6277,N_6383);
and U9829 (N_9829,N_7383,N_7358);
xor U9830 (N_9830,N_6414,N_6894);
xor U9831 (N_9831,N_7468,N_6883);
nor U9832 (N_9832,N_7542,N_6724);
nor U9833 (N_9833,N_6780,N_6110);
and U9834 (N_9834,N_7050,N_7501);
nor U9835 (N_9835,N_6876,N_6234);
nand U9836 (N_9836,N_6060,N_6683);
xnor U9837 (N_9837,N_7327,N_6733);
and U9838 (N_9838,N_7449,N_6179);
nand U9839 (N_9839,N_6173,N_6635);
nor U9840 (N_9840,N_7653,N_6793);
nor U9841 (N_9841,N_7754,N_7254);
xnor U9842 (N_9842,N_6803,N_6163);
xnor U9843 (N_9843,N_6116,N_7765);
nor U9844 (N_9844,N_6920,N_7765);
xor U9845 (N_9845,N_6040,N_6660);
or U9846 (N_9846,N_6593,N_6102);
xor U9847 (N_9847,N_7095,N_7607);
and U9848 (N_9848,N_7667,N_7357);
xor U9849 (N_9849,N_6931,N_6302);
nand U9850 (N_9850,N_7510,N_6015);
nor U9851 (N_9851,N_6156,N_6332);
or U9852 (N_9852,N_7347,N_6016);
xor U9853 (N_9853,N_6707,N_6636);
and U9854 (N_9854,N_6475,N_6663);
nor U9855 (N_9855,N_7787,N_6847);
and U9856 (N_9856,N_7679,N_6994);
nand U9857 (N_9857,N_6875,N_6453);
nand U9858 (N_9858,N_6468,N_6569);
nor U9859 (N_9859,N_7429,N_6318);
or U9860 (N_9860,N_7847,N_7828);
xor U9861 (N_9861,N_6300,N_6747);
and U9862 (N_9862,N_6449,N_6880);
nand U9863 (N_9863,N_7968,N_7620);
or U9864 (N_9864,N_6624,N_6241);
xnor U9865 (N_9865,N_7803,N_6169);
xor U9866 (N_9866,N_7652,N_7012);
nor U9867 (N_9867,N_6008,N_7393);
nor U9868 (N_9868,N_6233,N_6488);
nand U9869 (N_9869,N_7083,N_6871);
and U9870 (N_9870,N_6715,N_6081);
or U9871 (N_9871,N_6106,N_7468);
or U9872 (N_9872,N_7268,N_7622);
nand U9873 (N_9873,N_7963,N_6990);
or U9874 (N_9874,N_6624,N_6449);
nand U9875 (N_9875,N_7981,N_7151);
and U9876 (N_9876,N_6209,N_6058);
nor U9877 (N_9877,N_7884,N_6961);
nor U9878 (N_9878,N_7540,N_6393);
and U9879 (N_9879,N_6866,N_7588);
or U9880 (N_9880,N_6144,N_7160);
xor U9881 (N_9881,N_6216,N_7434);
and U9882 (N_9882,N_6205,N_7121);
xnor U9883 (N_9883,N_7972,N_6102);
nor U9884 (N_9884,N_6050,N_6579);
nand U9885 (N_9885,N_7331,N_6273);
xnor U9886 (N_9886,N_7613,N_6760);
and U9887 (N_9887,N_6862,N_6480);
xnor U9888 (N_9888,N_7014,N_6944);
xnor U9889 (N_9889,N_6519,N_7518);
xnor U9890 (N_9890,N_6687,N_7003);
nand U9891 (N_9891,N_6292,N_7998);
and U9892 (N_9892,N_6671,N_6482);
nor U9893 (N_9893,N_7525,N_7990);
nor U9894 (N_9894,N_7355,N_6477);
or U9895 (N_9895,N_6202,N_7875);
xor U9896 (N_9896,N_7360,N_7284);
xnor U9897 (N_9897,N_7255,N_6592);
nand U9898 (N_9898,N_7847,N_7620);
nor U9899 (N_9899,N_6007,N_6409);
xnor U9900 (N_9900,N_6194,N_6238);
and U9901 (N_9901,N_7886,N_6654);
nor U9902 (N_9902,N_7864,N_6560);
xor U9903 (N_9903,N_7979,N_7366);
nor U9904 (N_9904,N_6961,N_6524);
xnor U9905 (N_9905,N_7633,N_6121);
nand U9906 (N_9906,N_7569,N_7383);
or U9907 (N_9907,N_6706,N_7829);
or U9908 (N_9908,N_6521,N_7873);
or U9909 (N_9909,N_7435,N_6154);
nor U9910 (N_9910,N_6308,N_6893);
nor U9911 (N_9911,N_6605,N_7651);
xnor U9912 (N_9912,N_6534,N_6033);
nor U9913 (N_9913,N_6392,N_7708);
nor U9914 (N_9914,N_6225,N_7635);
nand U9915 (N_9915,N_7895,N_6730);
or U9916 (N_9916,N_7695,N_6571);
and U9917 (N_9917,N_7402,N_6962);
or U9918 (N_9918,N_6358,N_6101);
nand U9919 (N_9919,N_7668,N_7378);
nor U9920 (N_9920,N_7657,N_7926);
xnor U9921 (N_9921,N_7047,N_7170);
nand U9922 (N_9922,N_6617,N_7021);
xor U9923 (N_9923,N_6729,N_7988);
nor U9924 (N_9924,N_6560,N_6234);
nand U9925 (N_9925,N_7735,N_6498);
and U9926 (N_9926,N_6083,N_6889);
xor U9927 (N_9927,N_6358,N_6960);
xor U9928 (N_9928,N_6133,N_7697);
xor U9929 (N_9929,N_6456,N_6827);
xnor U9930 (N_9930,N_6845,N_7067);
or U9931 (N_9931,N_6021,N_6866);
nor U9932 (N_9932,N_7324,N_7113);
nand U9933 (N_9933,N_7801,N_7394);
nor U9934 (N_9934,N_7782,N_6776);
or U9935 (N_9935,N_6962,N_7448);
or U9936 (N_9936,N_6408,N_7904);
or U9937 (N_9937,N_6994,N_6404);
nand U9938 (N_9938,N_7617,N_6312);
xor U9939 (N_9939,N_6443,N_7447);
nand U9940 (N_9940,N_6968,N_6074);
nand U9941 (N_9941,N_6343,N_6257);
nor U9942 (N_9942,N_6530,N_7180);
and U9943 (N_9943,N_7380,N_6315);
and U9944 (N_9944,N_7222,N_7559);
xor U9945 (N_9945,N_6372,N_6725);
nand U9946 (N_9946,N_6498,N_6670);
xnor U9947 (N_9947,N_6438,N_6781);
and U9948 (N_9948,N_7718,N_7850);
xnor U9949 (N_9949,N_6537,N_7336);
and U9950 (N_9950,N_6406,N_7403);
nand U9951 (N_9951,N_7966,N_7238);
nor U9952 (N_9952,N_7994,N_6011);
and U9953 (N_9953,N_7562,N_6847);
xnor U9954 (N_9954,N_7992,N_6377);
nand U9955 (N_9955,N_7206,N_7709);
and U9956 (N_9956,N_6478,N_7528);
nor U9957 (N_9957,N_6617,N_7024);
xnor U9958 (N_9958,N_7146,N_6728);
xnor U9959 (N_9959,N_7663,N_6070);
or U9960 (N_9960,N_6069,N_7747);
nand U9961 (N_9961,N_7897,N_6226);
or U9962 (N_9962,N_6945,N_6100);
or U9963 (N_9963,N_7681,N_6504);
or U9964 (N_9964,N_7766,N_6577);
xor U9965 (N_9965,N_7939,N_6061);
and U9966 (N_9966,N_7220,N_7076);
nand U9967 (N_9967,N_6511,N_6429);
or U9968 (N_9968,N_7334,N_7524);
or U9969 (N_9969,N_6363,N_7521);
nand U9970 (N_9970,N_7704,N_6629);
xor U9971 (N_9971,N_7334,N_7106);
or U9972 (N_9972,N_6509,N_6404);
or U9973 (N_9973,N_6692,N_6714);
nand U9974 (N_9974,N_7861,N_6429);
or U9975 (N_9975,N_6796,N_7516);
nand U9976 (N_9976,N_7410,N_6660);
nor U9977 (N_9977,N_6850,N_6196);
xor U9978 (N_9978,N_7716,N_6300);
and U9979 (N_9979,N_7280,N_6748);
xor U9980 (N_9980,N_6857,N_7781);
xnor U9981 (N_9981,N_7974,N_6838);
nor U9982 (N_9982,N_7706,N_6404);
nand U9983 (N_9983,N_7994,N_6240);
xnor U9984 (N_9984,N_6374,N_7390);
nand U9985 (N_9985,N_6207,N_6962);
nor U9986 (N_9986,N_6965,N_7877);
and U9987 (N_9987,N_7942,N_6240);
or U9988 (N_9988,N_6581,N_7519);
nor U9989 (N_9989,N_7877,N_6587);
xnor U9990 (N_9990,N_6789,N_6267);
nand U9991 (N_9991,N_7950,N_7135);
or U9992 (N_9992,N_7650,N_6536);
or U9993 (N_9993,N_7671,N_6379);
xor U9994 (N_9994,N_6862,N_7954);
nor U9995 (N_9995,N_6174,N_7825);
and U9996 (N_9996,N_7237,N_6865);
or U9997 (N_9997,N_6188,N_7123);
xor U9998 (N_9998,N_6555,N_6966);
or U9999 (N_9999,N_7678,N_6555);
nor U10000 (N_10000,N_9902,N_8618);
and U10001 (N_10001,N_9969,N_8539);
or U10002 (N_10002,N_9550,N_9838);
nor U10003 (N_10003,N_8706,N_8547);
or U10004 (N_10004,N_8005,N_9579);
xnor U10005 (N_10005,N_8336,N_8074);
or U10006 (N_10006,N_8368,N_9340);
or U10007 (N_10007,N_9193,N_8669);
nor U10008 (N_10008,N_9758,N_8117);
xnor U10009 (N_10009,N_9986,N_9745);
nand U10010 (N_10010,N_9393,N_9091);
or U10011 (N_10011,N_9649,N_8762);
nand U10012 (N_10012,N_9822,N_8974);
nand U10013 (N_10013,N_8955,N_8533);
xnor U10014 (N_10014,N_8782,N_9026);
and U10015 (N_10015,N_8876,N_8361);
and U10016 (N_10016,N_9118,N_8788);
nor U10017 (N_10017,N_8932,N_9061);
or U10018 (N_10018,N_8779,N_8888);
nand U10019 (N_10019,N_8075,N_9709);
or U10020 (N_10020,N_9071,N_9212);
or U10021 (N_10021,N_9789,N_8123);
nand U10022 (N_10022,N_9763,N_8459);
nor U10023 (N_10023,N_8844,N_9820);
nor U10024 (N_10024,N_9366,N_9946);
nor U10025 (N_10025,N_9547,N_9596);
nor U10026 (N_10026,N_9689,N_9405);
nand U10027 (N_10027,N_8715,N_9055);
nor U10028 (N_10028,N_8236,N_8068);
or U10029 (N_10029,N_8081,N_8319);
xnor U10030 (N_10030,N_9330,N_9487);
and U10031 (N_10031,N_9600,N_8880);
xor U10032 (N_10032,N_8770,N_8713);
nand U10033 (N_10033,N_8949,N_9185);
and U10034 (N_10034,N_9623,N_9300);
nand U10035 (N_10035,N_9034,N_9577);
nor U10036 (N_10036,N_8550,N_8785);
nor U10037 (N_10037,N_8507,N_8842);
xor U10038 (N_10038,N_8857,N_8233);
and U10039 (N_10039,N_9461,N_8093);
nand U10040 (N_10040,N_8742,N_8559);
or U10041 (N_10041,N_9933,N_8743);
xor U10042 (N_10042,N_9908,N_9270);
xnor U10043 (N_10043,N_8920,N_8603);
xnor U10044 (N_10044,N_9096,N_8396);
or U10045 (N_10045,N_9180,N_8486);
nor U10046 (N_10046,N_8029,N_9925);
nand U10047 (N_10047,N_8951,N_8690);
xor U10048 (N_10048,N_8724,N_9500);
and U10049 (N_10049,N_9204,N_9712);
nand U10050 (N_10050,N_8196,N_9168);
and U10051 (N_10051,N_9081,N_8247);
nand U10052 (N_10052,N_9602,N_9291);
nand U10053 (N_10053,N_9837,N_8449);
nand U10054 (N_10054,N_9974,N_9617);
and U10055 (N_10055,N_9786,N_8398);
xnor U10056 (N_10056,N_9785,N_9738);
or U10057 (N_10057,N_8381,N_8269);
or U10058 (N_10058,N_9750,N_8731);
nand U10059 (N_10059,N_8586,N_9509);
xor U10060 (N_10060,N_9188,N_8552);
nand U10061 (N_10061,N_9276,N_9422);
and U10062 (N_10062,N_8481,N_8971);
nand U10063 (N_10063,N_9201,N_8327);
nand U10064 (N_10064,N_9778,N_8546);
or U10065 (N_10065,N_9231,N_8443);
nand U10066 (N_10066,N_9216,N_8866);
nor U10067 (N_10067,N_8549,N_9351);
and U10068 (N_10068,N_8227,N_9961);
nor U10069 (N_10069,N_8088,N_8197);
and U10070 (N_10070,N_8085,N_8184);
or U10071 (N_10071,N_8030,N_9977);
nand U10072 (N_10072,N_8044,N_8835);
or U10073 (N_10073,N_9542,N_9251);
nand U10074 (N_10074,N_9315,N_8491);
xnor U10075 (N_10075,N_9691,N_8171);
xnor U10076 (N_10076,N_9962,N_9545);
xor U10077 (N_10077,N_9480,N_9981);
nor U10078 (N_10078,N_8682,N_9540);
nand U10079 (N_10079,N_9511,N_9283);
xor U10080 (N_10080,N_9620,N_9978);
nor U10081 (N_10081,N_9899,N_8947);
nand U10082 (N_10082,N_8066,N_8192);
or U10083 (N_10083,N_8148,N_8836);
nor U10084 (N_10084,N_8019,N_9896);
nor U10085 (N_10085,N_8011,N_8786);
and U10086 (N_10086,N_8458,N_9830);
xnor U10087 (N_10087,N_9581,N_9998);
nand U10088 (N_10088,N_8651,N_8598);
nand U10089 (N_10089,N_9433,N_9211);
or U10090 (N_10090,N_8521,N_8940);
nor U10091 (N_10091,N_8166,N_8277);
nor U10092 (N_10092,N_9816,N_8714);
nor U10093 (N_10093,N_9407,N_9895);
nand U10094 (N_10094,N_9713,N_8037);
or U10095 (N_10095,N_8446,N_8581);
xor U10096 (N_10096,N_9943,N_8245);
nor U10097 (N_10097,N_9373,N_8001);
and U10098 (N_10098,N_8622,N_8226);
nand U10099 (N_10099,N_8594,N_8606);
or U10100 (N_10100,N_8664,N_8772);
or U10101 (N_10101,N_8749,N_9170);
nor U10102 (N_10102,N_8004,N_8903);
and U10103 (N_10103,N_9099,N_8204);
nand U10104 (N_10104,N_9489,N_8878);
or U10105 (N_10105,N_9704,N_8364);
xnor U10106 (N_10106,N_8248,N_9095);
nor U10107 (N_10107,N_9406,N_8809);
nor U10108 (N_10108,N_8829,N_9834);
or U10109 (N_10109,N_9358,N_8355);
nor U10110 (N_10110,N_8700,N_9595);
and U10111 (N_10111,N_8806,N_9906);
xnor U10112 (N_10112,N_9606,N_8092);
nand U10113 (N_10113,N_9403,N_9225);
and U10114 (N_10114,N_8203,N_9284);
nor U10115 (N_10115,N_8211,N_9715);
xor U10116 (N_10116,N_9524,N_9835);
nor U10117 (N_10117,N_9268,N_9803);
and U10118 (N_10118,N_8988,N_8627);
nor U10119 (N_10119,N_8286,N_9131);
nor U10120 (N_10120,N_8031,N_9360);
and U10121 (N_10121,N_8432,N_8079);
nand U10122 (N_10122,N_9323,N_8576);
xnor U10123 (N_10123,N_9440,N_9828);
nand U10124 (N_10124,N_8597,N_8165);
nor U10125 (N_10125,N_9862,N_9458);
nand U10126 (N_10126,N_9066,N_9872);
xor U10127 (N_10127,N_9918,N_8214);
nor U10128 (N_10128,N_8383,N_8754);
xnor U10129 (N_10129,N_8050,N_9467);
nor U10130 (N_10130,N_9674,N_9367);
and U10131 (N_10131,N_8387,N_8474);
and U10132 (N_10132,N_9074,N_9381);
nor U10133 (N_10133,N_9516,N_9255);
nand U10134 (N_10134,N_9249,N_8267);
nor U10135 (N_10135,N_8264,N_8045);
xor U10136 (N_10136,N_9355,N_9448);
or U10137 (N_10137,N_9636,N_9028);
nand U10138 (N_10138,N_9339,N_8747);
xnor U10139 (N_10139,N_8262,N_8290);
or U10140 (N_10140,N_8385,N_8401);
xnor U10141 (N_10141,N_9648,N_9389);
and U10142 (N_10142,N_9451,N_8761);
and U10143 (N_10143,N_9000,N_9885);
and U10144 (N_10144,N_9285,N_8116);
xor U10145 (N_10145,N_9082,N_8944);
or U10146 (N_10146,N_9863,N_8450);
nand U10147 (N_10147,N_9025,N_8934);
and U10148 (N_10148,N_8232,N_9727);
xor U10149 (N_10149,N_8753,N_9097);
or U10150 (N_10150,N_8078,N_9804);
nand U10151 (N_10151,N_9894,N_9496);
nor U10152 (N_10152,N_8055,N_8198);
and U10153 (N_10153,N_8511,N_9575);
xor U10154 (N_10154,N_9236,N_8111);
or U10155 (N_10155,N_9200,N_8456);
nand U10156 (N_10156,N_8331,N_9569);
nor U10157 (N_10157,N_9703,N_8989);
or U10158 (N_10158,N_9277,N_8154);
or U10159 (N_10159,N_9769,N_9777);
xor U10160 (N_10160,N_8482,N_8362);
or U10161 (N_10161,N_8419,N_8624);
nor U10162 (N_10162,N_8140,N_9821);
nand U10163 (N_10163,N_8833,N_9077);
xor U10164 (N_10164,N_8811,N_8457);
xnor U10165 (N_10165,N_8418,N_8750);
and U10166 (N_10166,N_9207,N_8670);
nor U10167 (N_10167,N_8129,N_8689);
or U10168 (N_10168,N_8153,N_9714);
and U10169 (N_10169,N_9658,N_8912);
nor U10170 (N_10170,N_8984,N_9797);
and U10171 (N_10171,N_9528,N_9701);
xor U10172 (N_10172,N_9049,N_8515);
or U10173 (N_10173,N_9047,N_9673);
nand U10174 (N_10174,N_8483,N_8508);
nor U10175 (N_10175,N_9829,N_8900);
nand U10176 (N_10176,N_9603,N_8520);
nor U10177 (N_10177,N_9419,N_8643);
xor U10178 (N_10178,N_9431,N_9149);
nor U10179 (N_10179,N_8239,N_8122);
and U10180 (N_10180,N_8144,N_8592);
and U10181 (N_10181,N_9337,N_9555);
or U10182 (N_10182,N_8720,N_8869);
xnor U10183 (N_10183,N_8544,N_8615);
or U10184 (N_10184,N_8370,N_8015);
and U10185 (N_10185,N_9332,N_8366);
or U10186 (N_10186,N_8193,N_9811);
or U10187 (N_10187,N_9352,N_9086);
nand U10188 (N_10188,N_9967,N_8047);
and U10189 (N_10189,N_9481,N_8565);
nor U10190 (N_10190,N_8571,N_8677);
nand U10191 (N_10191,N_9983,N_8250);
and U10192 (N_10192,N_8188,N_9772);
xor U10193 (N_10193,N_8879,N_9436);
xnor U10194 (N_10194,N_8617,N_9464);
nand U10195 (N_10195,N_9274,N_9048);
or U10196 (N_10196,N_8616,N_8463);
or U10197 (N_10197,N_8475,N_9767);
xnor U10198 (N_10198,N_9995,N_9073);
and U10199 (N_10199,N_9333,N_8796);
xor U10200 (N_10200,N_8126,N_9080);
or U10201 (N_10201,N_8252,N_9697);
or U10202 (N_10202,N_9587,N_9956);
and U10203 (N_10203,N_8119,N_8444);
nor U10204 (N_10204,N_8378,N_8426);
xnor U10205 (N_10205,N_8234,N_8964);
nor U10206 (N_10206,N_9369,N_8910);
nand U10207 (N_10207,N_8337,N_8212);
nor U10208 (N_10208,N_9809,N_9425);
xor U10209 (N_10209,N_8229,N_8591);
nor U10210 (N_10210,N_9243,N_8114);
or U10211 (N_10211,N_8404,N_8816);
nor U10212 (N_10212,N_9378,N_8678);
or U10213 (N_10213,N_8914,N_9105);
nor U10214 (N_10214,N_8377,N_8014);
and U10215 (N_10215,N_8696,N_8871);
nor U10216 (N_10216,N_9363,N_8864);
nor U10217 (N_10217,N_9331,N_8175);
xor U10218 (N_10218,N_9043,N_8656);
nand U10219 (N_10219,N_8469,N_9666);
or U10220 (N_10220,N_8408,N_9794);
or U10221 (N_10221,N_9904,N_9326);
xnor U10222 (N_10222,N_8840,N_8342);
or U10223 (N_10223,N_8798,N_9447);
nor U10224 (N_10224,N_9039,N_9860);
nor U10225 (N_10225,N_8961,N_8261);
or U10226 (N_10226,N_8440,N_9650);
and U10227 (N_10227,N_8256,N_8106);
nor U10228 (N_10228,N_9841,N_8025);
xnor U10229 (N_10229,N_9934,N_9221);
and U10230 (N_10230,N_9508,N_8919);
or U10231 (N_10231,N_8219,N_8978);
or U10232 (N_10232,N_8650,N_9759);
xnor U10233 (N_10233,N_9898,N_8332);
nor U10234 (N_10234,N_9825,N_8548);
xnor U10235 (N_10235,N_9571,N_8825);
or U10236 (N_10236,N_8411,N_8545);
xor U10237 (N_10237,N_8688,N_9965);
xor U10238 (N_10238,N_8722,N_8453);
nor U10239 (N_10239,N_8202,N_8858);
nor U10240 (N_10240,N_9659,N_8136);
and U10241 (N_10241,N_8455,N_8213);
nor U10242 (N_10242,N_9215,N_9226);
nor U10243 (N_10243,N_9321,N_8557);
and U10244 (N_10244,N_8841,N_9779);
nand U10245 (N_10245,N_8354,N_8846);
or U10246 (N_10246,N_8767,N_9046);
and U10247 (N_10247,N_8413,N_9134);
nor U10248 (N_10248,N_8287,N_8847);
nor U10249 (N_10249,N_8200,N_9390);
nor U10250 (N_10250,N_8069,N_9817);
nand U10251 (N_10251,N_8205,N_9948);
or U10252 (N_10252,N_9437,N_9783);
nand U10253 (N_10253,N_8317,N_8296);
xnor U10254 (N_10254,N_9229,N_8537);
xor U10255 (N_10255,N_8107,N_8610);
xnor U10256 (N_10256,N_9669,N_8735);
nand U10257 (N_10257,N_8938,N_8304);
and U10258 (N_10258,N_8054,N_8830);
nor U10259 (N_10259,N_8963,N_8372);
and U10260 (N_10260,N_9409,N_8705);
nor U10261 (N_10261,N_9526,N_9824);
nand U10262 (N_10262,N_8771,N_8348);
nand U10263 (N_10263,N_9143,N_9865);
or U10264 (N_10264,N_8099,N_8283);
xnor U10265 (N_10265,N_8943,N_9755);
or U10266 (N_10266,N_9850,N_9734);
or U10267 (N_10267,N_9963,N_9970);
or U10268 (N_10268,N_8409,N_8693);
xnor U10269 (N_10269,N_9051,N_8240);
and U10270 (N_10270,N_9334,N_9890);
nor U10271 (N_10271,N_8431,N_9724);
or U10272 (N_10272,N_9147,N_9338);
and U10273 (N_10273,N_9175,N_8745);
xor U10274 (N_10274,N_8983,N_8913);
nand U10275 (N_10275,N_9470,N_9126);
nand U10276 (N_10276,N_9722,N_8080);
or U10277 (N_10277,N_8769,N_8422);
or U10278 (N_10278,N_8959,N_8895);
nand U10279 (N_10279,N_8863,N_8502);
nand U10280 (N_10280,N_8764,N_9123);
and U10281 (N_10281,N_9905,N_8230);
and U10282 (N_10282,N_8568,N_8077);
or U10283 (N_10283,N_8330,N_9146);
nand U10284 (N_10284,N_8916,N_9459);
and U10285 (N_10285,N_9917,N_9937);
nor U10286 (N_10286,N_8562,N_8575);
xnor U10287 (N_10287,N_8326,N_8967);
xor U10288 (N_10288,N_9991,N_9417);
and U10289 (N_10289,N_8733,N_9197);
and U10290 (N_10290,N_8393,N_9566);
xnor U10291 (N_10291,N_8340,N_8254);
xnor U10292 (N_10292,N_9973,N_9442);
xnor U10293 (N_10293,N_8942,N_8495);
xnor U10294 (N_10294,N_9657,N_9923);
xnor U10295 (N_10295,N_9029,N_9434);
or U10296 (N_10296,N_9324,N_9064);
or U10297 (N_10297,N_9031,N_8740);
xor U10298 (N_10298,N_9130,N_9719);
and U10299 (N_10299,N_9079,N_9490);
xnor U10300 (N_10300,N_9716,N_9241);
and U10301 (N_10301,N_8890,N_8135);
nand U10302 (N_10302,N_9612,N_9423);
nor U10303 (N_10303,N_8347,N_9037);
and U10304 (N_10304,N_8746,N_8633);
or U10305 (N_10305,N_8259,N_9747);
or U10306 (N_10306,N_8852,N_8896);
and U10307 (N_10307,N_8324,N_9676);
or U10308 (N_10308,N_8636,N_8341);
nand U10309 (N_10309,N_9058,N_9370);
xor U10310 (N_10310,N_8087,N_8773);
nor U10311 (N_10311,N_9445,N_9296);
nand U10312 (N_10312,N_9594,N_8725);
nor U10313 (N_10313,N_8002,N_8020);
nor U10314 (N_10314,N_8373,N_8108);
nand U10315 (N_10315,N_9760,N_9158);
nor U10316 (N_10316,N_9012,N_9304);
xor U10317 (N_10317,N_9202,N_9021);
nor U10318 (N_10318,N_8501,N_9678);
nor U10319 (N_10319,N_8777,N_9242);
xnor U10320 (N_10320,N_8139,N_8886);
or U10321 (N_10321,N_8569,N_9013);
or U10322 (N_10322,N_9735,N_9743);
nor U10323 (N_10323,N_9667,N_8194);
or U10324 (N_10324,N_8101,N_9223);
xor U10325 (N_10325,N_8338,N_8875);
nand U10326 (N_10326,N_9893,N_8307);
or U10327 (N_10327,N_9926,N_9533);
xor U10328 (N_10328,N_9640,N_8026);
xnor U10329 (N_10329,N_8975,N_9279);
and U10330 (N_10330,N_9465,N_8648);
nand U10331 (N_10331,N_8371,N_9394);
nor U10332 (N_10332,N_8487,N_8414);
nor U10333 (N_10333,N_9848,N_8589);
nand U10334 (N_10334,N_9087,N_8803);
xnor U10335 (N_10335,N_9989,N_9380);
xor U10336 (N_10336,N_9644,N_8007);
or U10337 (N_10337,N_8588,N_9260);
or U10338 (N_10338,N_8388,N_9453);
or U10339 (N_10339,N_8865,N_8113);
xor U10340 (N_10340,N_9883,N_9607);
xnor U10341 (N_10341,N_8496,N_8358);
nand U10342 (N_10342,N_8110,N_8590);
and U10343 (N_10343,N_9843,N_9628);
and U10344 (N_10344,N_8350,N_9611);
or U10345 (N_10345,N_9294,N_8845);
and U10346 (N_10346,N_8468,N_9597);
or U10347 (N_10347,N_8512,N_9368);
and U10348 (N_10348,N_9144,N_8436);
xnor U10349 (N_10349,N_9990,N_8536);
nand U10350 (N_10350,N_8018,N_8904);
and U10351 (N_10351,N_9022,N_8191);
nor U10352 (N_10352,N_9686,N_8780);
nand U10353 (N_10353,N_9664,N_9397);
xnor U10354 (N_10354,N_8817,N_9011);
xnor U10355 (N_10355,N_8893,N_9371);
nor U10356 (N_10356,N_8685,N_9094);
nor U10357 (N_10357,N_9795,N_8478);
nand U10358 (N_10358,N_9780,N_9477);
nor U10359 (N_10359,N_8323,N_8022);
nand U10360 (N_10360,N_9941,N_8125);
nand U10361 (N_10361,N_8021,N_8936);
nand U10362 (N_10362,N_8161,N_9139);
and U10363 (N_10363,N_8497,N_9135);
xnor U10364 (N_10364,N_9377,N_8861);
and U10365 (N_10365,N_9398,N_9015);
and U10366 (N_10366,N_9627,N_8853);
and U10367 (N_10367,N_9151,N_9230);
nand U10368 (N_10368,N_9093,N_8281);
and U10369 (N_10369,N_9732,N_9023);
nand U10370 (N_10370,N_9936,N_8570);
nor U10371 (N_10371,N_8527,N_8902);
xnor U10372 (N_10372,N_8711,N_9375);
nand U10373 (N_10373,N_8352,N_9960);
and U10374 (N_10374,N_8519,N_8666);
nand U10375 (N_10375,N_9815,N_8472);
or U10376 (N_10376,N_8003,N_9953);
or U10377 (N_10377,N_9773,N_8158);
and U10378 (N_10378,N_9810,N_8579);
or U10379 (N_10379,N_9726,N_9537);
nor U10380 (N_10380,N_8132,N_8027);
nor U10381 (N_10381,N_9444,N_8578);
and U10382 (N_10382,N_8676,N_9827);
xnor U10383 (N_10383,N_9741,N_9859);
xor U10384 (N_10384,N_8400,N_8278);
nor U10385 (N_10385,N_8048,N_8702);
xnor U10386 (N_10386,N_9928,N_8553);
xnor U10387 (N_10387,N_9036,N_8784);
nand U10388 (N_10388,N_8929,N_9114);
xnor U10389 (N_10389,N_8433,N_9387);
nor U10390 (N_10390,N_9009,N_8577);
or U10391 (N_10391,N_8775,N_8424);
nor U10392 (N_10392,N_8216,N_9038);
or U10393 (N_10393,N_9104,N_9210);
and U10394 (N_10394,N_9040,N_9111);
and U10395 (N_10395,N_9832,N_9452);
nand U10396 (N_10396,N_8270,N_8966);
or U10397 (N_10397,N_9167,N_9984);
nand U10398 (N_10398,N_9125,N_9997);
or U10399 (N_10399,N_9016,N_9282);
or U10400 (N_10400,N_9247,N_8405);
nor U10401 (N_10401,N_8768,N_9632);
or U10402 (N_10402,N_9532,N_8941);
or U10403 (N_10403,N_8612,N_9462);
or U10404 (N_10404,N_8462,N_9761);
xor U10405 (N_10405,N_9224,N_9610);
or U10406 (N_10406,N_9162,N_9754);
nand U10407 (N_10407,N_9505,N_9115);
and U10408 (N_10408,N_9705,N_9749);
and U10409 (N_10409,N_9148,N_9349);
nand U10410 (N_10410,N_9090,N_9002);
and U10411 (N_10411,N_8672,N_8661);
or U10412 (N_10412,N_9866,N_8112);
and U10413 (N_10413,N_9313,N_8905);
xnor U10414 (N_10414,N_8391,N_9631);
nor U10415 (N_10415,N_8976,N_9519);
nor U10416 (N_10416,N_9121,N_8346);
nand U10417 (N_10417,N_8009,N_9529);
and U10418 (N_10418,N_8542,N_8675);
and U10419 (N_10419,N_9565,N_8421);
xnor U10420 (N_10420,N_9518,N_8345);
or U10421 (N_10421,N_9350,N_8505);
nand U10422 (N_10422,N_8320,N_9306);
nand U10423 (N_10423,N_9858,N_8309);
nor U10424 (N_10424,N_8339,N_8827);
or U10425 (N_10425,N_8314,N_9302);
nand U10426 (N_10426,N_9538,N_8266);
nor U10427 (N_10427,N_9557,N_8255);
and U10428 (N_10428,N_8102,N_9141);
xnor U10429 (N_10429,N_8429,N_9515);
nor U10430 (N_10430,N_9062,N_8222);
nand U10431 (N_10431,N_9930,N_9473);
or U10432 (N_10432,N_8856,N_9307);
or U10433 (N_10433,N_9235,N_8170);
xor U10434 (N_10434,N_8103,N_8611);
nand U10435 (N_10435,N_8086,N_9053);
or U10436 (N_10436,N_9922,N_8057);
and U10437 (N_10437,N_9567,N_8820);
nor U10438 (N_10438,N_8684,N_8221);
nor U10439 (N_10439,N_8146,N_8982);
and U10440 (N_10440,N_8084,N_9110);
nand U10441 (N_10441,N_9027,N_9041);
nor U10442 (N_10442,N_9892,N_8766);
xor U10443 (N_10443,N_9101,N_9554);
or U10444 (N_10444,N_9897,N_8822);
or U10445 (N_10445,N_8038,N_8891);
nor U10446 (N_10446,N_8168,N_9488);
or U10447 (N_10447,N_9695,N_8757);
nor U10448 (N_10448,N_9033,N_9067);
xor U10449 (N_10449,N_9539,N_9069);
nor U10450 (N_10450,N_9868,N_8185);
xor U10451 (N_10451,N_8187,N_8156);
and U10452 (N_10452,N_9228,N_9399);
and U10453 (N_10453,N_9152,N_8774);
or U10454 (N_10454,N_8778,N_8793);
or U10455 (N_10455,N_8489,N_9171);
or U10456 (N_10456,N_8376,N_9248);
nor U10457 (N_10457,N_9740,N_9849);
nor U10458 (N_10458,N_8253,N_9641);
nand U10459 (N_10459,N_8637,N_9684);
nand U10460 (N_10460,N_9173,N_8040);
nor U10461 (N_10461,N_8127,N_8737);
nor U10462 (N_10462,N_8169,N_9454);
xor U10463 (N_10463,N_9214,N_9254);
nor U10464 (N_10464,N_9308,N_9138);
or U10465 (N_10465,N_8076,N_8873);
xor U10466 (N_10466,N_9559,N_9757);
or U10467 (N_10467,N_9878,N_8210);
or U10468 (N_10468,N_8041,N_8760);
nor U10469 (N_10469,N_8979,N_8884);
nand U10470 (N_10470,N_9006,N_8924);
nand U10471 (N_10471,N_9840,N_8867);
and U10472 (N_10472,N_9874,N_9700);
nor U10473 (N_10473,N_9548,N_9955);
and U10474 (N_10474,N_9831,N_9233);
xor U10475 (N_10475,N_9971,N_8284);
and U10476 (N_10476,N_8524,N_9792);
nor U10477 (N_10477,N_9927,N_8329);
or U10478 (N_10478,N_8823,N_9347);
nand U10479 (N_10479,N_8131,N_9359);
xnor U10480 (N_10480,N_8560,N_8805);
or U10481 (N_10481,N_9169,N_8176);
nand U10482 (N_10482,N_9301,N_9106);
nand U10483 (N_10483,N_8096,N_8687);
and U10484 (N_10484,N_8667,N_8901);
xnor U10485 (N_10485,N_8375,N_9471);
xor U10486 (N_10486,N_8128,N_8937);
nand U10487 (N_10487,N_8473,N_9784);
and U10488 (N_10488,N_8763,N_8639);
nand U10489 (N_10489,N_8091,N_8289);
nand U10490 (N_10490,N_8625,N_8503);
and U10491 (N_10491,N_8062,N_8889);
xor U10492 (N_10492,N_9531,N_8972);
nand U10493 (N_10493,N_9160,N_9671);
nor U10494 (N_10494,N_8417,N_8855);
nor U10495 (N_10495,N_9271,N_9706);
nand U10496 (N_10496,N_8958,N_8072);
and U10497 (N_10497,N_8828,N_9942);
or U10498 (N_10498,N_9589,N_9463);
xor U10499 (N_10499,N_9314,N_9245);
nor U10500 (N_10500,N_9309,N_8596);
or U10501 (N_10501,N_9582,N_9154);
xnor U10502 (N_10502,N_8199,N_9357);
and U10503 (N_10503,N_9267,N_9564);
and U10504 (N_10504,N_9818,N_8065);
xnor U10505 (N_10505,N_9621,N_8752);
and U10506 (N_10506,N_9469,N_9072);
and U10507 (N_10507,N_9092,N_9573);
xnor U10508 (N_10508,N_8147,N_8490);
or U10509 (N_10509,N_8160,N_8999);
and U10510 (N_10510,N_8063,N_8881);
nor U10511 (N_10511,N_9497,N_8797);
and U10512 (N_10512,N_8945,N_9568);
xnor U10513 (N_10513,N_9208,N_8023);
nand U10514 (N_10514,N_8668,N_8427);
nand U10515 (N_10515,N_8298,N_9317);
nor U10516 (N_10516,N_9864,N_8406);
xor U10517 (N_10517,N_9003,N_9551);
and U10518 (N_10518,N_9278,N_8950);
nand U10519 (N_10519,N_9781,N_9753);
or U10520 (N_10520,N_9875,N_9052);
xnor U10521 (N_10521,N_9698,N_9172);
or U10522 (N_10522,N_9520,N_9661);
and U10523 (N_10523,N_9484,N_8118);
nand U10524 (N_10524,N_9685,N_8271);
and U10525 (N_10525,N_8172,N_8470);
nor U10526 (N_10526,N_8815,N_9512);
and U10527 (N_10527,N_9263,N_8629);
nand U10528 (N_10528,N_8654,N_9570);
xnor U10529 (N_10529,N_9506,N_8741);
and U10530 (N_10530,N_9530,N_8514);
nor U10531 (N_10531,N_8862,N_8303);
or U10532 (N_10532,N_9476,N_8053);
or U10533 (N_10533,N_9861,N_9702);
or U10534 (N_10534,N_8516,N_9999);
or U10535 (N_10535,N_9889,N_9654);
xor U10536 (N_10536,N_9075,N_8585);
and U10537 (N_10537,N_8328,N_8969);
or U10538 (N_10538,N_8981,N_8476);
or U10539 (N_10539,N_9576,N_8268);
or U10540 (N_10540,N_8732,N_9288);
or U10541 (N_10541,N_9915,N_9157);
and U10542 (N_10542,N_9909,N_9517);
nand U10543 (N_10543,N_8995,N_9468);
nor U10544 (N_10544,N_8821,N_9653);
or U10545 (N_10545,N_9482,N_9968);
nand U10546 (N_10546,N_9731,N_9402);
xor U10547 (N_10547,N_9376,N_8532);
or U10548 (N_10548,N_9218,N_9017);
xnor U10549 (N_10549,N_9266,N_9007);
and U10550 (N_10550,N_9498,N_9592);
and U10551 (N_10551,N_8035,N_9494);
xor U10552 (N_10552,N_9382,N_9787);
and U10553 (N_10553,N_9608,N_9639);
nand U10554 (N_10554,N_8697,N_9790);
xor U10555 (N_10555,N_8386,N_9624);
nand U10556 (N_10556,N_9992,N_8311);
or U10557 (N_10557,N_8305,N_8282);
and U10558 (N_10558,N_9944,N_9156);
xor U10559 (N_10559,N_9305,N_9299);
nand U10560 (N_10560,N_8095,N_9921);
nand U10561 (N_10561,N_8294,N_8564);
and U10562 (N_10562,N_9290,N_9558);
xnor U10563 (N_10563,N_9578,N_9253);
nor U10564 (N_10564,N_9356,N_9165);
or U10565 (N_10565,N_8641,N_8343);
nor U10566 (N_10566,N_9931,N_9109);
nand U10567 (N_10567,N_9042,N_8471);
nor U10568 (N_10568,N_8201,N_8538);
xnor U10569 (N_10569,N_9122,N_9774);
nand U10570 (N_10570,N_8179,N_8794);
and U10571 (N_10571,N_9766,N_8703);
or U10572 (N_10572,N_8365,N_8083);
or U10573 (N_10573,N_8935,N_9396);
nor U10574 (N_10574,N_8051,N_8952);
xor U10575 (N_10575,N_9670,N_9525);
and U10576 (N_10576,N_9113,N_8789);
xor U10577 (N_10577,N_8619,N_9384);
xor U10578 (N_10578,N_9854,N_8334);
xor U10579 (N_10579,N_8605,N_8556);
and U10580 (N_10580,N_9812,N_8157);
or U10581 (N_10581,N_9107,N_8885);
nand U10582 (N_10582,N_9174,N_9708);
xor U10583 (N_10583,N_9823,N_8504);
nand U10584 (N_10584,N_8056,N_8887);
xnor U10585 (N_10585,N_9262,N_9329);
xnor U10586 (N_10586,N_8407,N_8509);
nand U10587 (N_10587,N_9456,N_8759);
nand U10588 (N_10588,N_9450,N_9327);
and U10589 (N_10589,N_8518,N_8241);
nor U10590 (N_10590,N_9259,N_8645);
or U10591 (N_10591,N_8224,N_8839);
or U10592 (N_10592,N_8279,N_9001);
xnor U10593 (N_10593,N_8838,N_8189);
or U10594 (N_10594,N_8244,N_9879);
or U10595 (N_10595,N_9428,N_9421);
and U10596 (N_10596,N_9510,N_9916);
or U10597 (N_10597,N_8206,N_8640);
xor U10598 (N_10598,N_9945,N_9386);
nor U10599 (N_10599,N_9045,N_8464);
and U10600 (N_10600,N_8799,N_8583);
or U10601 (N_10601,N_8379,N_8218);
and U10602 (N_10602,N_9063,N_9054);
nor U10603 (N_10603,N_9742,N_9756);
nand U10604 (N_10604,N_9637,N_8164);
and U10605 (N_10605,N_8691,N_9178);
nand U10606 (N_10606,N_9070,N_9935);
nor U10607 (N_10607,N_8899,N_8089);
xnor U10608 (N_10608,N_9388,N_9788);
nand U10609 (N_10609,N_9762,N_8874);
or U10610 (N_10610,N_8238,N_8563);
and U10611 (N_10611,N_9361,N_8181);
and U10612 (N_10612,N_8990,N_8609);
nand U10613 (N_10613,N_8356,N_9663);
and U10614 (N_10614,N_9681,N_9613);
nor U10615 (N_10615,N_9993,N_8061);
nand U10616 (N_10616,N_8526,N_9826);
xnor U10617 (N_10617,N_9884,N_8921);
and U10618 (N_10618,N_9994,N_9867);
nand U10619 (N_10619,N_9257,N_9598);
or U10620 (N_10620,N_9083,N_8868);
xnor U10621 (N_10621,N_9982,N_8993);
or U10622 (N_10622,N_9181,N_8152);
nand U10623 (N_10623,N_9322,N_8996);
and U10624 (N_10624,N_8987,N_9707);
nand U10625 (N_10625,N_8712,N_8814);
nand U10626 (N_10626,N_9415,N_8783);
xnor U10627 (N_10627,N_9808,N_9239);
nand U10628 (N_10628,N_9354,N_8228);
xnor U10629 (N_10629,N_8930,N_8756);
and U10630 (N_10630,N_8382,N_9493);
and U10631 (N_10631,N_9298,N_9920);
nor U10632 (N_10632,N_9699,N_9438);
nor U10633 (N_10633,N_9882,N_9544);
nand U10634 (N_10634,N_9910,N_8448);
or U10635 (N_10635,N_9183,N_9335);
nand U10636 (N_10636,N_9507,N_8800);
or U10637 (N_10637,N_9374,N_8953);
xnor U10638 (N_10638,N_9744,N_9987);
xnor U10639 (N_10639,N_9005,N_9751);
nand U10640 (N_10640,N_8802,N_8430);
nor U10641 (N_10641,N_9234,N_8215);
or U10642 (N_10642,N_8595,N_8465);
or U10643 (N_10643,N_8225,N_9057);
and U10644 (N_10644,N_8810,N_9552);
nand U10645 (N_10645,N_9629,N_8727);
nor U10646 (N_10646,N_8531,N_9084);
nor U10647 (N_10647,N_8998,N_9127);
xnor U10648 (N_10648,N_8917,N_9219);
nand U10649 (N_10649,N_8291,N_9264);
nand U10650 (N_10650,N_8566,N_9913);
xor U10651 (N_10651,N_8173,N_8402);
xor U10652 (N_10652,N_8860,N_9010);
or U10653 (N_10653,N_9736,N_9919);
nor U10654 (N_10654,N_8297,N_9668);
nor U10655 (N_10655,N_8109,N_8790);
xor U10656 (N_10656,N_8986,N_8190);
nand U10657 (N_10657,N_8013,N_9474);
and U10658 (N_10658,N_9646,N_8658);
xor U10659 (N_10659,N_9833,N_9227);
and U10660 (N_10660,N_9441,N_8321);
or U10661 (N_10661,N_8500,N_9205);
nor U10662 (N_10662,N_9996,N_8620);
nand U10663 (N_10663,N_9887,N_8049);
or U10664 (N_10664,N_8384,N_9630);
nand U10665 (N_10665,N_8447,N_9798);
nor U10666 (N_10666,N_9728,N_8580);
or U10667 (N_10667,N_9591,N_9720);
and U10668 (N_10668,N_9710,N_8416);
or U10669 (N_10669,N_8831,N_8686);
or U10670 (N_10670,N_9546,N_8601);
xnor U10671 (N_10671,N_9572,N_8985);
and U10672 (N_10672,N_8104,N_9198);
nand U10673 (N_10673,N_9807,N_8363);
xor U10674 (N_10674,N_9588,N_8755);
nand U10675 (N_10675,N_8392,N_9609);
and U10676 (N_10676,N_9599,N_8349);
nand U10677 (N_10677,N_8679,N_9319);
nand U10678 (N_10678,N_8058,N_9132);
or U10679 (N_10679,N_8607,N_8442);
or U10680 (N_10680,N_9343,N_9404);
or U10681 (N_10681,N_8602,N_8306);
nor U10682 (N_10682,N_9059,N_9411);
nand U10683 (N_10683,N_8723,N_8425);
xnor U10684 (N_10684,N_9232,N_8302);
nor U10685 (N_10685,N_9966,N_9583);
xnor U10686 (N_10686,N_8274,N_9238);
and U10687 (N_10687,N_9163,N_8150);
xor U10688 (N_10688,N_8510,N_8142);
nand U10689 (N_10689,N_9793,N_9656);
or U10690 (N_10690,N_9903,N_8374);
nor U10691 (N_10691,N_8626,N_9503);
nor U10692 (N_10692,N_9137,N_8134);
and U10693 (N_10693,N_9643,N_8397);
nand U10694 (N_10694,N_9203,N_9900);
nor U10695 (N_10695,N_8813,N_9586);
and U10696 (N_10696,N_9342,N_9891);
nor U10697 (N_10697,N_9975,N_9379);
or U10698 (N_10698,N_9362,N_8801);
nand U10699 (N_10699,N_8217,N_9292);
and U10700 (N_10700,N_9618,N_8968);
and U10701 (N_10701,N_8410,N_8299);
nor U10702 (N_10702,N_9561,N_8451);
or U10703 (N_10703,N_9801,N_8265);
nand U10704 (N_10704,N_9439,N_9957);
and U10705 (N_10705,N_8992,N_8632);
xor U10706 (N_10706,N_8739,N_9950);
nand U10707 (N_10707,N_9182,N_8659);
nand U10708 (N_10708,N_9929,N_8698);
nand U10709 (N_10709,N_8517,N_9240);
nand U10710 (N_10710,N_8412,N_8071);
nand U10711 (N_10711,N_8848,N_8804);
nand U10712 (N_10712,N_8043,N_8906);
xnor U10713 (N_10713,N_9014,N_8059);
nand U10714 (N_10714,N_8671,N_9938);
xor U10715 (N_10715,N_9189,N_9341);
or U10716 (N_10716,N_8353,N_8621);
xor U10717 (N_10717,N_8843,N_9281);
nor U10718 (N_10718,N_9881,N_8965);
xnor U10719 (N_10719,N_9112,N_8033);
nand U10720 (N_10720,N_9847,N_8623);
nand U10721 (N_10721,N_9626,N_9196);
nand U10722 (N_10722,N_8008,N_8631);
nor U10723 (N_10723,N_8420,N_9024);
nand U10724 (N_10724,N_9056,N_9652);
nand U10725 (N_10725,N_9870,N_8060);
or U10726 (N_10726,N_8155,N_8434);
nor U10727 (N_10727,N_8115,N_9293);
nand U10728 (N_10728,N_9222,N_8994);
xnor U10729 (N_10729,N_8728,N_9019);
xor U10730 (N_10730,N_8390,N_9844);
and U10731 (N_10731,N_8251,N_9845);
nand U10732 (N_10732,N_9802,N_9513);
nand U10733 (N_10733,N_8380,N_8834);
and U10734 (N_10734,N_9244,N_9395);
or U10735 (N_10735,N_8898,N_9269);
xnor U10736 (N_10736,N_8660,N_8477);
xor U10737 (N_10737,N_9680,N_8918);
xor U10738 (N_10738,N_9392,N_9187);
and U10739 (N_10739,N_8243,N_9076);
nand U10740 (N_10740,N_9190,N_8644);
nor U10741 (N_10741,N_8663,N_8138);
nand U10742 (N_10742,N_9871,N_9102);
nor U10743 (N_10743,N_8012,N_9964);
nand U10744 (N_10744,N_8024,N_8911);
nor U10745 (N_10745,N_8467,N_9721);
or U10746 (N_10746,N_9690,N_8067);
nor U10747 (N_10747,N_9100,N_9297);
and U10748 (N_10748,N_8017,N_8105);
nor U10749 (N_10749,N_9796,N_9195);
nand U10750 (N_10750,N_9560,N_8708);
xnor U10751 (N_10751,N_8883,N_9348);
nand U10752 (N_10752,N_9687,N_9806);
nor U10753 (N_10753,N_9932,N_9336);
xnor U10754 (N_10754,N_8599,N_8870);
xor U10755 (N_10755,N_9289,N_9764);
nand U10756 (N_10756,N_8555,N_8130);
or U10757 (N_10757,N_9514,N_8534);
nand U10758 (N_10758,N_9725,N_8716);
and U10759 (N_10759,N_9672,N_9768);
xnor U10760 (N_10760,N_8275,N_9880);
nand U10761 (N_10761,N_8293,N_8795);
nand U10762 (N_10762,N_8032,N_8541);
nand U10763 (N_10763,N_9574,N_9344);
xor U10764 (N_10764,N_9770,N_8614);
or U10765 (N_10765,N_9692,N_9273);
and U10766 (N_10766,N_9030,N_9694);
or U10767 (N_10767,N_8628,N_8312);
nor U10768 (N_10768,N_8454,N_9638);
and U10769 (N_10769,N_9886,N_8121);
and U10770 (N_10770,N_9791,N_9541);
nor U10771 (N_10771,N_8039,N_8133);
nand U10772 (N_10772,N_9733,N_9522);
or U10773 (N_10773,N_9133,N_8479);
nand U10774 (N_10774,N_9217,N_8167);
xnor U10775 (N_10775,N_9136,N_8235);
xor U10776 (N_10776,N_8638,N_9988);
or U10777 (N_10777,N_9472,N_8832);
or U10778 (N_10778,N_8791,N_8034);
or U10779 (N_10779,N_9128,N_9819);
and U10780 (N_10780,N_8540,N_8681);
nor U10781 (N_10781,N_8183,N_8273);
nor U10782 (N_10782,N_9947,N_8719);
xor U10783 (N_10783,N_8090,N_8851);
xor U10784 (N_10784,N_9958,N_8600);
nand U10785 (N_10785,N_8389,N_9287);
and U10786 (N_10786,N_8246,N_8701);
and U10787 (N_10787,N_9914,N_9479);
nand U10788 (N_10788,N_8792,N_9166);
nand U10789 (N_10789,N_8933,N_8776);
or U10790 (N_10790,N_9979,N_8915);
and U10791 (N_10791,N_8494,N_9486);
nand U10792 (N_10792,N_8461,N_8073);
or U10793 (N_10793,N_9853,N_9584);
xnor U10794 (N_10794,N_9176,N_9846);
nand U10795 (N_10795,N_9206,N_8525);
and U10796 (N_10796,N_9145,N_9408);
nand U10797 (N_10797,N_8751,N_8124);
or U10798 (N_10798,N_8907,N_8649);
or U10799 (N_10799,N_9718,N_9655);
nand U10800 (N_10800,N_9625,N_9549);
and U10801 (N_10801,N_9164,N_8530);
and U10802 (N_10802,N_8635,N_9590);
nor U10803 (N_10803,N_8209,N_9466);
nand U10804 (N_10804,N_8322,N_9103);
or U10805 (N_10805,N_8946,N_9085);
xor U10806 (N_10806,N_8100,N_8908);
nor U10807 (N_10807,N_9677,N_9616);
nand U10808 (N_10808,N_9739,N_9800);
or U10809 (N_10809,N_9060,N_8046);
xor U10810 (N_10810,N_8439,N_8973);
nand U10811 (N_10811,N_8826,N_8182);
xor U10812 (N_10812,N_8535,N_8954);
and U10813 (N_10813,N_8894,N_9427);
xnor U10814 (N_10814,N_9907,N_8149);
nor U10815 (N_10815,N_9534,N_9593);
and U10816 (N_10816,N_8094,N_9153);
nand U10817 (N_10817,N_9924,N_8926);
nand U10818 (N_10818,N_9199,N_9839);
xor U10819 (N_10819,N_9499,N_9633);
nand U10820 (N_10820,N_9035,N_8333);
xor U10821 (N_10821,N_9604,N_9478);
and U10822 (N_10822,N_9852,N_8849);
nand U10823 (N_10823,N_9446,N_8765);
nand U10824 (N_10824,N_9065,N_9413);
nor U10825 (N_10825,N_8683,N_9008);
or U10826 (N_10826,N_9246,N_9855);
xor U10827 (N_10827,N_8781,N_8036);
or U10828 (N_10828,N_8415,N_8403);
or U10829 (N_10829,N_9457,N_9120);
nor U10830 (N_10830,N_9108,N_9688);
and U10831 (N_10831,N_8258,N_9443);
and U10832 (N_10832,N_9737,N_8498);
xnor U10833 (N_10833,N_9265,N_8445);
nand U10834 (N_10834,N_9683,N_9495);
nand U10835 (N_10835,N_9432,N_9295);
nand U10836 (N_10836,N_9435,N_8977);
nor U10837 (N_10837,N_8276,N_8151);
xor U10838 (N_10838,N_9536,N_9050);
nand U10839 (N_10839,N_8016,N_8163);
nand U10840 (N_10840,N_8939,N_9004);
xor U10841 (N_10841,N_9475,N_9418);
nor U10842 (N_10842,N_9353,N_8082);
nand U10843 (N_10843,N_8647,N_9799);
xor U10844 (N_10844,N_8423,N_9192);
and U10845 (N_10845,N_9078,N_9972);
nor U10846 (N_10846,N_8042,N_9400);
nand U10847 (N_10847,N_8543,N_8980);
and U10848 (N_10848,N_8485,N_8308);
xnor U10849 (N_10849,N_8070,N_9776);
xor U10850 (N_10850,N_8730,N_9275);
nand U10851 (N_10851,N_9385,N_8316);
xnor U10852 (N_10852,N_9044,N_9068);
or U10853 (N_10853,N_8351,N_9954);
and U10854 (N_10854,N_8242,N_8285);
nand U10855 (N_10855,N_8220,N_9679);
nor U10856 (N_10856,N_8877,N_8707);
nand U10857 (N_10857,N_8923,N_9696);
and U10858 (N_10858,N_9911,N_9980);
nor U10859 (N_10859,N_8301,N_8499);
or U10860 (N_10860,N_8177,N_9771);
nand U10861 (N_10861,N_9032,N_8710);
nor U10862 (N_10862,N_9647,N_9585);
xor U10863 (N_10863,N_8850,N_8726);
and U10864 (N_10864,N_9098,N_8582);
and U10865 (N_10865,N_9645,N_8295);
nand U10866 (N_10866,N_8748,N_8231);
xnor U10867 (N_10867,N_8604,N_8584);
xor U10868 (N_10868,N_9634,N_9746);
and U10869 (N_10869,N_9730,N_9316);
and U10870 (N_10870,N_8897,N_8699);
or U10871 (N_10871,N_9191,N_8466);
nand U10872 (N_10872,N_8962,N_8662);
nand U10873 (N_10873,N_9901,N_8709);
or U10874 (N_10874,N_8787,N_8642);
nand U10875 (N_10875,N_9876,N_9580);
nand U10876 (N_10876,N_8310,N_9449);
xnor U10877 (N_10877,N_9426,N_9455);
nor U10878 (N_10878,N_8927,N_9401);
xor U10879 (N_10879,N_8704,N_9420);
and U10880 (N_10880,N_9543,N_9345);
nand U10881 (N_10881,N_9250,N_8249);
or U10882 (N_10882,N_9416,N_8159);
xor U10883 (N_10883,N_8280,N_8523);
xnor U10884 (N_10884,N_8052,N_9310);
nand U10885 (N_10885,N_9765,N_9563);
nor U10886 (N_10886,N_9959,N_9912);
xor U10887 (N_10887,N_8186,N_9635);
nor U10888 (N_10888,N_8925,N_8695);
nand U10889 (N_10889,N_8292,N_8344);
nor U10890 (N_10890,N_8028,N_9985);
nor U10891 (N_10891,N_9142,N_9364);
xor U10892 (N_10892,N_8854,N_8572);
and U10893 (N_10893,N_9949,N_8484);
or U10894 (N_10894,N_8812,N_8325);
and U10895 (N_10895,N_8573,N_8970);
xnor U10896 (N_10896,N_8394,N_8437);
nor U10897 (N_10897,N_8064,N_8593);
or U10898 (N_10898,N_8729,N_9615);
xnor U10899 (N_10899,N_9527,N_8652);
or U10900 (N_10900,N_9662,N_9723);
or U10901 (N_10901,N_8438,N_8692);
and U10902 (N_10902,N_9280,N_9140);
and U10903 (N_10903,N_9124,N_9501);
or U10904 (N_10904,N_9020,N_9752);
or U10905 (N_10905,N_9129,N_8721);
or U10906 (N_10906,N_9256,N_9491);
or U10907 (N_10907,N_9492,N_8718);
nor U10908 (N_10908,N_8882,N_9325);
nor U10909 (N_10909,N_8097,N_9018);
nor U10910 (N_10910,N_9311,N_8460);
nor U10911 (N_10911,N_9729,N_9535);
xnor U10912 (N_10912,N_8006,N_8997);
and U10913 (N_10913,N_9430,N_8957);
and U10914 (N_10914,N_9089,N_8808);
xor U10915 (N_10915,N_9150,N_9318);
and U10916 (N_10916,N_9682,N_9814);
xnor U10917 (N_10917,N_9424,N_8807);
or U10918 (N_10918,N_9888,N_9877);
or U10919 (N_10919,N_8928,N_8960);
xnor U10920 (N_10920,N_9873,N_8435);
and U10921 (N_10921,N_8357,N_9504);
and U10922 (N_10922,N_8528,N_8657);
nor U10923 (N_10923,N_9951,N_9605);
xnor U10924 (N_10924,N_8288,N_8318);
or U10925 (N_10925,N_8892,N_9088);
nor U10926 (N_10926,N_8208,N_9601);
nor U10927 (N_10927,N_8480,N_8207);
xnor U10928 (N_10928,N_8137,N_8263);
xnor U10929 (N_10929,N_8143,N_8694);
or U10930 (N_10930,N_8673,N_9272);
nor U10931 (N_10931,N_9328,N_9976);
xor U10932 (N_10932,N_8315,N_9320);
nor U10933 (N_10933,N_8313,N_8837);
and U10934 (N_10934,N_8665,N_9258);
or U10935 (N_10935,N_8680,N_8162);
nor U10936 (N_10936,N_9521,N_9412);
xnor U10937 (N_10937,N_8738,N_9414);
nor U10938 (N_10938,N_9651,N_8819);
xor U10939 (N_10939,N_9303,N_9119);
nor U10940 (N_10940,N_9952,N_8367);
nand U10941 (N_10941,N_8872,N_9161);
or U10942 (N_10942,N_9748,N_9940);
nor U10943 (N_10943,N_9159,N_8141);
or U10944 (N_10944,N_9857,N_8567);
and U10945 (N_10945,N_9116,N_8174);
nand U10946 (N_10946,N_8195,N_8634);
xnor U10947 (N_10947,N_9553,N_8506);
xnor U10948 (N_10948,N_9775,N_9179);
nor U10949 (N_10949,N_9220,N_9642);
nand U10950 (N_10950,N_8574,N_8561);
or U10951 (N_10951,N_8646,N_8145);
and U10952 (N_10952,N_9213,N_9665);
nor U10953 (N_10953,N_8000,N_8513);
nand U10954 (N_10954,N_8824,N_8488);
and U10955 (N_10955,N_8441,N_9562);
nand U10956 (N_10956,N_9460,N_8948);
and U10957 (N_10957,N_8744,N_9391);
nand U10958 (N_10958,N_8758,N_9660);
nor U10959 (N_10959,N_9194,N_9117);
and U10960 (N_10960,N_9252,N_9836);
nand U10961 (N_10961,N_9856,N_8587);
nand U10962 (N_10962,N_8956,N_8608);
nor U10963 (N_10963,N_9556,N_8734);
nand U10964 (N_10964,N_8359,N_9614);
nand U10965 (N_10965,N_9851,N_8223);
nand U10966 (N_10966,N_9523,N_8395);
nor U10967 (N_10967,N_8630,N_9237);
nor U10968 (N_10968,N_9429,N_8674);
nor U10969 (N_10969,N_8717,N_8529);
nand U10970 (N_10970,N_9622,N_9483);
and U10971 (N_10971,N_9261,N_8452);
xor U10972 (N_10972,N_9485,N_9782);
nor U10973 (N_10973,N_9693,N_9869);
nand U10974 (N_10974,N_8428,N_8300);
nand U10975 (N_10975,N_9383,N_9410);
or U10976 (N_10976,N_8399,N_9155);
xor U10977 (N_10977,N_8010,N_9372);
nand U10978 (N_10978,N_8492,N_8613);
xnor U10979 (N_10979,N_9346,N_8522);
nor U10980 (N_10980,N_9286,N_9209);
nor U10981 (N_10981,N_9675,N_9939);
or U10982 (N_10982,N_8909,N_9186);
or U10983 (N_10983,N_8493,N_8554);
nor U10984 (N_10984,N_8859,N_8178);
xor U10985 (N_10985,N_8922,N_8260);
and U10986 (N_10986,N_9717,N_9184);
nand U10987 (N_10987,N_9711,N_9177);
nand U10988 (N_10988,N_8655,N_8360);
nor U10989 (N_10989,N_8931,N_9813);
and U10990 (N_10990,N_8180,N_9805);
nand U10991 (N_10991,N_8551,N_8818);
xor U10992 (N_10992,N_8558,N_8653);
and U10993 (N_10993,N_8098,N_8257);
or U10994 (N_10994,N_8120,N_8991);
and U10995 (N_10995,N_9619,N_9365);
and U10996 (N_10996,N_8335,N_8237);
nand U10997 (N_10997,N_8736,N_8369);
nand U10998 (N_10998,N_9842,N_8272);
nand U10999 (N_10999,N_9312,N_9502);
nand U11000 (N_11000,N_9945,N_9270);
nand U11001 (N_11001,N_8323,N_8804);
nor U11002 (N_11002,N_8532,N_8967);
xor U11003 (N_11003,N_8354,N_9571);
or U11004 (N_11004,N_8143,N_8233);
nand U11005 (N_11005,N_8104,N_9844);
or U11006 (N_11006,N_9848,N_9010);
nor U11007 (N_11007,N_8888,N_9246);
xor U11008 (N_11008,N_9347,N_9993);
nor U11009 (N_11009,N_8208,N_9082);
and U11010 (N_11010,N_8759,N_9609);
and U11011 (N_11011,N_9491,N_8008);
xnor U11012 (N_11012,N_8756,N_9447);
or U11013 (N_11013,N_8559,N_8321);
nor U11014 (N_11014,N_8888,N_9249);
or U11015 (N_11015,N_8480,N_9973);
or U11016 (N_11016,N_9795,N_9262);
and U11017 (N_11017,N_8862,N_8446);
and U11018 (N_11018,N_8269,N_8222);
and U11019 (N_11019,N_8050,N_9355);
nand U11020 (N_11020,N_8507,N_8908);
xor U11021 (N_11021,N_8911,N_8441);
nor U11022 (N_11022,N_8844,N_8712);
nor U11023 (N_11023,N_8064,N_9604);
nand U11024 (N_11024,N_9153,N_9651);
nand U11025 (N_11025,N_9288,N_9089);
or U11026 (N_11026,N_9950,N_8312);
nor U11027 (N_11027,N_8368,N_8791);
xor U11028 (N_11028,N_8130,N_8509);
nor U11029 (N_11029,N_8163,N_8980);
nor U11030 (N_11030,N_8416,N_8120);
and U11031 (N_11031,N_9412,N_9948);
nand U11032 (N_11032,N_9354,N_9397);
nand U11033 (N_11033,N_9266,N_9622);
xor U11034 (N_11034,N_9681,N_9052);
or U11035 (N_11035,N_8453,N_8868);
xor U11036 (N_11036,N_9083,N_9148);
nor U11037 (N_11037,N_8073,N_8476);
nand U11038 (N_11038,N_9608,N_9688);
and U11039 (N_11039,N_9752,N_8226);
or U11040 (N_11040,N_8641,N_9294);
nor U11041 (N_11041,N_9633,N_9677);
xor U11042 (N_11042,N_8788,N_9086);
xnor U11043 (N_11043,N_9843,N_8606);
and U11044 (N_11044,N_8245,N_9485);
nor U11045 (N_11045,N_8894,N_8501);
and U11046 (N_11046,N_8817,N_9127);
xor U11047 (N_11047,N_9055,N_9880);
nor U11048 (N_11048,N_8197,N_9071);
and U11049 (N_11049,N_9688,N_9786);
and U11050 (N_11050,N_9555,N_8204);
nor U11051 (N_11051,N_8411,N_9039);
nand U11052 (N_11052,N_9560,N_8501);
or U11053 (N_11053,N_9144,N_8170);
xor U11054 (N_11054,N_8866,N_9830);
xor U11055 (N_11055,N_8770,N_9068);
xor U11056 (N_11056,N_9690,N_9752);
nor U11057 (N_11057,N_9942,N_8115);
nor U11058 (N_11058,N_9106,N_9208);
nor U11059 (N_11059,N_8749,N_9815);
nor U11060 (N_11060,N_9217,N_9416);
nor U11061 (N_11061,N_8616,N_9290);
xnor U11062 (N_11062,N_8229,N_9044);
nor U11063 (N_11063,N_8248,N_9217);
xor U11064 (N_11064,N_8928,N_8796);
nand U11065 (N_11065,N_9983,N_8090);
nor U11066 (N_11066,N_8520,N_8811);
nand U11067 (N_11067,N_9631,N_9868);
nor U11068 (N_11068,N_8327,N_9670);
nor U11069 (N_11069,N_8812,N_8080);
and U11070 (N_11070,N_8993,N_9330);
and U11071 (N_11071,N_8643,N_9997);
nand U11072 (N_11072,N_9079,N_8871);
and U11073 (N_11073,N_8588,N_9121);
xor U11074 (N_11074,N_8383,N_9766);
xnor U11075 (N_11075,N_8051,N_8948);
or U11076 (N_11076,N_9277,N_9597);
or U11077 (N_11077,N_9133,N_8102);
nand U11078 (N_11078,N_8686,N_8666);
nand U11079 (N_11079,N_9575,N_8866);
nand U11080 (N_11080,N_8191,N_8090);
xor U11081 (N_11081,N_9583,N_9705);
and U11082 (N_11082,N_9193,N_9339);
and U11083 (N_11083,N_9638,N_9109);
nand U11084 (N_11084,N_9506,N_8948);
and U11085 (N_11085,N_9464,N_8062);
and U11086 (N_11086,N_8868,N_9488);
and U11087 (N_11087,N_8970,N_9367);
nand U11088 (N_11088,N_9080,N_9159);
and U11089 (N_11089,N_9184,N_9149);
xnor U11090 (N_11090,N_9232,N_9727);
and U11091 (N_11091,N_9262,N_8740);
and U11092 (N_11092,N_9449,N_8273);
or U11093 (N_11093,N_8603,N_8891);
xor U11094 (N_11094,N_8551,N_9164);
nor U11095 (N_11095,N_9915,N_8711);
nor U11096 (N_11096,N_9696,N_9190);
nand U11097 (N_11097,N_9025,N_9009);
nand U11098 (N_11098,N_8069,N_8751);
and U11099 (N_11099,N_8398,N_9992);
and U11100 (N_11100,N_8696,N_8675);
and U11101 (N_11101,N_9201,N_9354);
nand U11102 (N_11102,N_8360,N_9240);
xor U11103 (N_11103,N_8149,N_8745);
or U11104 (N_11104,N_8544,N_9946);
xor U11105 (N_11105,N_9064,N_8443);
nor U11106 (N_11106,N_9437,N_8121);
or U11107 (N_11107,N_8176,N_9650);
nand U11108 (N_11108,N_9712,N_9368);
or U11109 (N_11109,N_9233,N_8376);
nand U11110 (N_11110,N_8924,N_8826);
or U11111 (N_11111,N_9238,N_9754);
nor U11112 (N_11112,N_8806,N_8776);
nand U11113 (N_11113,N_9982,N_8182);
or U11114 (N_11114,N_9905,N_9212);
and U11115 (N_11115,N_9766,N_9793);
or U11116 (N_11116,N_9476,N_9250);
xor U11117 (N_11117,N_9870,N_8479);
xor U11118 (N_11118,N_8135,N_9168);
nand U11119 (N_11119,N_8514,N_8248);
xnor U11120 (N_11120,N_8064,N_9665);
nand U11121 (N_11121,N_8641,N_8894);
xnor U11122 (N_11122,N_9295,N_8447);
xor U11123 (N_11123,N_9787,N_9302);
xor U11124 (N_11124,N_8032,N_9320);
xnor U11125 (N_11125,N_9281,N_9772);
xor U11126 (N_11126,N_8633,N_8037);
or U11127 (N_11127,N_8783,N_8636);
nor U11128 (N_11128,N_8001,N_9705);
nor U11129 (N_11129,N_8027,N_9861);
nand U11130 (N_11130,N_8099,N_9481);
nor U11131 (N_11131,N_9067,N_8349);
xor U11132 (N_11132,N_9184,N_9641);
nand U11133 (N_11133,N_8238,N_8395);
nand U11134 (N_11134,N_8678,N_9108);
nor U11135 (N_11135,N_9970,N_8802);
and U11136 (N_11136,N_8066,N_8088);
nor U11137 (N_11137,N_8918,N_9051);
or U11138 (N_11138,N_9674,N_9498);
nor U11139 (N_11139,N_9998,N_8854);
and U11140 (N_11140,N_8401,N_8950);
nand U11141 (N_11141,N_8836,N_9329);
or U11142 (N_11142,N_8359,N_9909);
nand U11143 (N_11143,N_8529,N_8718);
or U11144 (N_11144,N_8383,N_8556);
and U11145 (N_11145,N_9863,N_9708);
and U11146 (N_11146,N_8787,N_9624);
xnor U11147 (N_11147,N_9593,N_8990);
xnor U11148 (N_11148,N_9041,N_8054);
and U11149 (N_11149,N_8320,N_8293);
nor U11150 (N_11150,N_8403,N_9830);
and U11151 (N_11151,N_9241,N_8695);
nor U11152 (N_11152,N_8781,N_9463);
xor U11153 (N_11153,N_8090,N_8742);
nor U11154 (N_11154,N_8685,N_9092);
nor U11155 (N_11155,N_8853,N_8918);
nand U11156 (N_11156,N_9377,N_8103);
or U11157 (N_11157,N_9028,N_9441);
nor U11158 (N_11158,N_8635,N_8655);
and U11159 (N_11159,N_8549,N_8878);
and U11160 (N_11160,N_9489,N_9527);
xnor U11161 (N_11161,N_8547,N_8068);
or U11162 (N_11162,N_9717,N_8174);
nor U11163 (N_11163,N_8787,N_9714);
nand U11164 (N_11164,N_8550,N_9833);
xor U11165 (N_11165,N_9366,N_9900);
xnor U11166 (N_11166,N_9807,N_8623);
xor U11167 (N_11167,N_9684,N_8469);
nand U11168 (N_11168,N_8251,N_9020);
xnor U11169 (N_11169,N_9545,N_8535);
xor U11170 (N_11170,N_9475,N_9976);
xnor U11171 (N_11171,N_8406,N_9694);
xor U11172 (N_11172,N_8349,N_9639);
nand U11173 (N_11173,N_8730,N_8674);
nand U11174 (N_11174,N_8009,N_8378);
xnor U11175 (N_11175,N_8222,N_9838);
xnor U11176 (N_11176,N_8464,N_9463);
and U11177 (N_11177,N_8608,N_8069);
or U11178 (N_11178,N_8048,N_8127);
or U11179 (N_11179,N_9239,N_9763);
xnor U11180 (N_11180,N_8389,N_8917);
and U11181 (N_11181,N_8574,N_8458);
nand U11182 (N_11182,N_9400,N_8782);
or U11183 (N_11183,N_8851,N_9426);
nor U11184 (N_11184,N_9252,N_9221);
and U11185 (N_11185,N_9214,N_9807);
and U11186 (N_11186,N_8065,N_9678);
nor U11187 (N_11187,N_8462,N_8902);
or U11188 (N_11188,N_9237,N_9921);
xnor U11189 (N_11189,N_8319,N_8687);
nand U11190 (N_11190,N_8116,N_8453);
and U11191 (N_11191,N_9488,N_8296);
nor U11192 (N_11192,N_8479,N_8386);
or U11193 (N_11193,N_8446,N_9124);
nand U11194 (N_11194,N_9372,N_8197);
xnor U11195 (N_11195,N_9927,N_9379);
nand U11196 (N_11196,N_9280,N_8762);
xor U11197 (N_11197,N_9152,N_8832);
nand U11198 (N_11198,N_9795,N_9859);
nor U11199 (N_11199,N_9480,N_8694);
or U11200 (N_11200,N_9036,N_8874);
or U11201 (N_11201,N_9727,N_8126);
nand U11202 (N_11202,N_8293,N_8350);
nand U11203 (N_11203,N_9050,N_9935);
xnor U11204 (N_11204,N_9240,N_9733);
nor U11205 (N_11205,N_9642,N_8192);
or U11206 (N_11206,N_9842,N_8602);
or U11207 (N_11207,N_9430,N_9110);
nand U11208 (N_11208,N_9352,N_9790);
and U11209 (N_11209,N_9073,N_8707);
nor U11210 (N_11210,N_8154,N_9974);
and U11211 (N_11211,N_9486,N_8560);
or U11212 (N_11212,N_9910,N_9840);
and U11213 (N_11213,N_8154,N_8982);
nor U11214 (N_11214,N_9175,N_9010);
xor U11215 (N_11215,N_8233,N_9168);
nor U11216 (N_11216,N_8852,N_8944);
xnor U11217 (N_11217,N_9789,N_8720);
and U11218 (N_11218,N_8484,N_8347);
xor U11219 (N_11219,N_8810,N_9716);
and U11220 (N_11220,N_8960,N_9127);
xor U11221 (N_11221,N_9597,N_8503);
nand U11222 (N_11222,N_9759,N_8202);
or U11223 (N_11223,N_8663,N_8017);
xnor U11224 (N_11224,N_8214,N_8236);
nand U11225 (N_11225,N_8275,N_9904);
or U11226 (N_11226,N_8130,N_8303);
nor U11227 (N_11227,N_8424,N_8781);
and U11228 (N_11228,N_8455,N_9738);
and U11229 (N_11229,N_8060,N_8481);
or U11230 (N_11230,N_8534,N_9304);
or U11231 (N_11231,N_9702,N_9934);
and U11232 (N_11232,N_9389,N_9912);
or U11233 (N_11233,N_8026,N_9871);
nand U11234 (N_11234,N_9537,N_9268);
nand U11235 (N_11235,N_8565,N_9478);
or U11236 (N_11236,N_9986,N_9221);
and U11237 (N_11237,N_8858,N_9145);
nor U11238 (N_11238,N_9799,N_8887);
and U11239 (N_11239,N_8874,N_9982);
nand U11240 (N_11240,N_9008,N_8061);
and U11241 (N_11241,N_9046,N_9806);
nand U11242 (N_11242,N_8834,N_9902);
and U11243 (N_11243,N_8576,N_9006);
and U11244 (N_11244,N_9648,N_8552);
nor U11245 (N_11245,N_9292,N_9293);
or U11246 (N_11246,N_9148,N_9460);
xor U11247 (N_11247,N_8985,N_8454);
nor U11248 (N_11248,N_9744,N_9524);
xnor U11249 (N_11249,N_8479,N_8732);
and U11250 (N_11250,N_9401,N_8161);
nor U11251 (N_11251,N_8870,N_9593);
nor U11252 (N_11252,N_9302,N_9678);
nand U11253 (N_11253,N_9786,N_9035);
xnor U11254 (N_11254,N_8050,N_8831);
xor U11255 (N_11255,N_9952,N_8520);
nor U11256 (N_11256,N_8743,N_9629);
nand U11257 (N_11257,N_8181,N_8233);
and U11258 (N_11258,N_8332,N_9782);
xnor U11259 (N_11259,N_9591,N_8931);
or U11260 (N_11260,N_8808,N_9962);
and U11261 (N_11261,N_8350,N_9985);
and U11262 (N_11262,N_8296,N_9325);
xnor U11263 (N_11263,N_9652,N_9265);
nand U11264 (N_11264,N_8691,N_9868);
or U11265 (N_11265,N_9736,N_8488);
and U11266 (N_11266,N_8314,N_9465);
or U11267 (N_11267,N_9210,N_8132);
and U11268 (N_11268,N_9442,N_9818);
or U11269 (N_11269,N_9681,N_9713);
or U11270 (N_11270,N_8385,N_9532);
xnor U11271 (N_11271,N_9241,N_8084);
or U11272 (N_11272,N_8272,N_9623);
nor U11273 (N_11273,N_9863,N_9293);
or U11274 (N_11274,N_8782,N_9372);
nand U11275 (N_11275,N_8491,N_9912);
nor U11276 (N_11276,N_9659,N_9689);
nor U11277 (N_11277,N_8558,N_8571);
nor U11278 (N_11278,N_8729,N_9541);
nor U11279 (N_11279,N_9652,N_9846);
or U11280 (N_11280,N_9575,N_8820);
or U11281 (N_11281,N_8731,N_9644);
xor U11282 (N_11282,N_8939,N_9752);
nor U11283 (N_11283,N_8895,N_8810);
and U11284 (N_11284,N_9812,N_9601);
nand U11285 (N_11285,N_8738,N_9413);
or U11286 (N_11286,N_8740,N_8789);
or U11287 (N_11287,N_9670,N_9226);
or U11288 (N_11288,N_8962,N_8837);
nor U11289 (N_11289,N_9451,N_9136);
and U11290 (N_11290,N_9663,N_9912);
xor U11291 (N_11291,N_8724,N_8548);
nand U11292 (N_11292,N_9967,N_9356);
or U11293 (N_11293,N_9523,N_9063);
nand U11294 (N_11294,N_9255,N_8822);
and U11295 (N_11295,N_9760,N_9286);
and U11296 (N_11296,N_8948,N_8439);
nand U11297 (N_11297,N_8605,N_9139);
or U11298 (N_11298,N_9924,N_9270);
or U11299 (N_11299,N_8161,N_8501);
or U11300 (N_11300,N_9017,N_8850);
or U11301 (N_11301,N_9324,N_8124);
xor U11302 (N_11302,N_8814,N_8500);
or U11303 (N_11303,N_8075,N_9203);
xor U11304 (N_11304,N_9614,N_8361);
xor U11305 (N_11305,N_9368,N_9522);
or U11306 (N_11306,N_9979,N_8483);
nor U11307 (N_11307,N_9062,N_9114);
nor U11308 (N_11308,N_9672,N_9352);
xor U11309 (N_11309,N_9277,N_9955);
nor U11310 (N_11310,N_9983,N_9971);
nor U11311 (N_11311,N_9715,N_9893);
and U11312 (N_11312,N_9289,N_8772);
nand U11313 (N_11313,N_9577,N_8395);
nor U11314 (N_11314,N_8110,N_9502);
or U11315 (N_11315,N_8763,N_8238);
nor U11316 (N_11316,N_8946,N_9950);
or U11317 (N_11317,N_9697,N_9046);
or U11318 (N_11318,N_9411,N_8121);
nand U11319 (N_11319,N_9783,N_8488);
nand U11320 (N_11320,N_9320,N_9097);
and U11321 (N_11321,N_8920,N_8839);
and U11322 (N_11322,N_9332,N_9606);
and U11323 (N_11323,N_8103,N_8937);
or U11324 (N_11324,N_9704,N_8326);
xnor U11325 (N_11325,N_9371,N_9785);
nor U11326 (N_11326,N_8060,N_8888);
xnor U11327 (N_11327,N_9501,N_8138);
xor U11328 (N_11328,N_8243,N_9340);
nor U11329 (N_11329,N_9721,N_9519);
nor U11330 (N_11330,N_9042,N_8827);
or U11331 (N_11331,N_9571,N_8657);
or U11332 (N_11332,N_9759,N_8803);
and U11333 (N_11333,N_9516,N_8108);
xor U11334 (N_11334,N_8264,N_9461);
and U11335 (N_11335,N_9466,N_9867);
and U11336 (N_11336,N_9146,N_9813);
nor U11337 (N_11337,N_9485,N_9217);
and U11338 (N_11338,N_9130,N_9071);
or U11339 (N_11339,N_8166,N_9789);
or U11340 (N_11340,N_9901,N_9467);
nand U11341 (N_11341,N_8568,N_9871);
xnor U11342 (N_11342,N_9401,N_8125);
or U11343 (N_11343,N_8651,N_8329);
xnor U11344 (N_11344,N_9765,N_8910);
xnor U11345 (N_11345,N_8198,N_9288);
and U11346 (N_11346,N_8627,N_9864);
and U11347 (N_11347,N_8405,N_9948);
xnor U11348 (N_11348,N_8309,N_9682);
xnor U11349 (N_11349,N_8668,N_9825);
or U11350 (N_11350,N_9109,N_9138);
or U11351 (N_11351,N_9933,N_8518);
nand U11352 (N_11352,N_9627,N_8248);
or U11353 (N_11353,N_8630,N_9306);
nor U11354 (N_11354,N_8900,N_9221);
xor U11355 (N_11355,N_8084,N_9944);
or U11356 (N_11356,N_8223,N_8404);
xor U11357 (N_11357,N_8764,N_8229);
and U11358 (N_11358,N_9427,N_8818);
xnor U11359 (N_11359,N_8725,N_8921);
xnor U11360 (N_11360,N_9124,N_9980);
nand U11361 (N_11361,N_9506,N_8092);
xnor U11362 (N_11362,N_9860,N_9720);
nand U11363 (N_11363,N_9402,N_9177);
xor U11364 (N_11364,N_8619,N_9786);
nand U11365 (N_11365,N_8759,N_9610);
xor U11366 (N_11366,N_9402,N_9204);
and U11367 (N_11367,N_9955,N_9306);
and U11368 (N_11368,N_8626,N_8081);
nor U11369 (N_11369,N_8393,N_9229);
xor U11370 (N_11370,N_8289,N_9479);
or U11371 (N_11371,N_9915,N_8380);
nand U11372 (N_11372,N_9515,N_8339);
nand U11373 (N_11373,N_8773,N_8313);
or U11374 (N_11374,N_8115,N_8650);
nor U11375 (N_11375,N_9524,N_8506);
nand U11376 (N_11376,N_8875,N_8535);
and U11377 (N_11377,N_9171,N_9609);
nor U11378 (N_11378,N_8001,N_8435);
and U11379 (N_11379,N_8761,N_8989);
and U11380 (N_11380,N_8352,N_9833);
and U11381 (N_11381,N_9645,N_8260);
xnor U11382 (N_11382,N_8984,N_9865);
xor U11383 (N_11383,N_9472,N_8091);
nor U11384 (N_11384,N_9261,N_8776);
nor U11385 (N_11385,N_8108,N_9318);
and U11386 (N_11386,N_8760,N_9750);
nor U11387 (N_11387,N_8984,N_8555);
and U11388 (N_11388,N_9587,N_8298);
or U11389 (N_11389,N_8621,N_9415);
nand U11390 (N_11390,N_9444,N_9664);
nor U11391 (N_11391,N_9490,N_9401);
and U11392 (N_11392,N_8792,N_9533);
nor U11393 (N_11393,N_8337,N_8330);
nand U11394 (N_11394,N_8802,N_8970);
nand U11395 (N_11395,N_8128,N_8713);
and U11396 (N_11396,N_9585,N_8452);
nand U11397 (N_11397,N_9118,N_9304);
and U11398 (N_11398,N_9431,N_9942);
nor U11399 (N_11399,N_8650,N_9792);
or U11400 (N_11400,N_8187,N_8997);
or U11401 (N_11401,N_9529,N_8953);
and U11402 (N_11402,N_9928,N_9293);
nor U11403 (N_11403,N_8059,N_9999);
xor U11404 (N_11404,N_8680,N_8886);
nand U11405 (N_11405,N_8043,N_8238);
or U11406 (N_11406,N_8636,N_8395);
or U11407 (N_11407,N_8839,N_8502);
xnor U11408 (N_11408,N_9993,N_9419);
nand U11409 (N_11409,N_9273,N_9746);
and U11410 (N_11410,N_8444,N_9229);
nand U11411 (N_11411,N_8934,N_9893);
and U11412 (N_11412,N_9102,N_9290);
nor U11413 (N_11413,N_9965,N_9439);
xor U11414 (N_11414,N_8985,N_8157);
or U11415 (N_11415,N_8222,N_9670);
nand U11416 (N_11416,N_8031,N_9515);
and U11417 (N_11417,N_9978,N_9119);
or U11418 (N_11418,N_8928,N_8167);
nand U11419 (N_11419,N_8635,N_8896);
and U11420 (N_11420,N_8697,N_8673);
xor U11421 (N_11421,N_9577,N_8756);
nand U11422 (N_11422,N_8302,N_8000);
and U11423 (N_11423,N_9926,N_8822);
or U11424 (N_11424,N_8973,N_9880);
nand U11425 (N_11425,N_9688,N_9236);
nand U11426 (N_11426,N_8245,N_8847);
nand U11427 (N_11427,N_8875,N_9171);
xor U11428 (N_11428,N_9173,N_9704);
or U11429 (N_11429,N_9450,N_8082);
xnor U11430 (N_11430,N_9518,N_8105);
xnor U11431 (N_11431,N_9654,N_9916);
and U11432 (N_11432,N_9366,N_8141);
and U11433 (N_11433,N_9800,N_8583);
nor U11434 (N_11434,N_9495,N_8426);
and U11435 (N_11435,N_8396,N_9496);
or U11436 (N_11436,N_8148,N_9232);
and U11437 (N_11437,N_8325,N_9495);
nand U11438 (N_11438,N_9713,N_8590);
nand U11439 (N_11439,N_9027,N_9594);
nand U11440 (N_11440,N_8587,N_8871);
nor U11441 (N_11441,N_8846,N_8357);
xor U11442 (N_11442,N_8317,N_8213);
and U11443 (N_11443,N_8894,N_8180);
nand U11444 (N_11444,N_8275,N_8164);
nor U11445 (N_11445,N_9089,N_8035);
or U11446 (N_11446,N_8848,N_8574);
or U11447 (N_11447,N_9340,N_8813);
nor U11448 (N_11448,N_8569,N_8239);
or U11449 (N_11449,N_9953,N_9491);
nor U11450 (N_11450,N_8223,N_8306);
and U11451 (N_11451,N_8151,N_8133);
xor U11452 (N_11452,N_9406,N_9219);
nand U11453 (N_11453,N_9303,N_8078);
xor U11454 (N_11454,N_8997,N_8663);
nand U11455 (N_11455,N_9950,N_9808);
and U11456 (N_11456,N_9370,N_9481);
and U11457 (N_11457,N_8627,N_8087);
nor U11458 (N_11458,N_9215,N_8522);
or U11459 (N_11459,N_9115,N_9733);
xor U11460 (N_11460,N_9079,N_9753);
nand U11461 (N_11461,N_9126,N_8910);
xnor U11462 (N_11462,N_8575,N_9515);
nand U11463 (N_11463,N_8131,N_8425);
xor U11464 (N_11464,N_8695,N_9664);
or U11465 (N_11465,N_8646,N_8279);
and U11466 (N_11466,N_9133,N_8677);
xnor U11467 (N_11467,N_8772,N_9832);
xor U11468 (N_11468,N_9250,N_9288);
or U11469 (N_11469,N_9918,N_8303);
nor U11470 (N_11470,N_8377,N_9304);
and U11471 (N_11471,N_9490,N_8484);
xor U11472 (N_11472,N_9012,N_8437);
nand U11473 (N_11473,N_9717,N_8992);
nand U11474 (N_11474,N_9593,N_8633);
xnor U11475 (N_11475,N_9956,N_8657);
and U11476 (N_11476,N_9174,N_8925);
or U11477 (N_11477,N_9127,N_9062);
nor U11478 (N_11478,N_8748,N_9255);
xor U11479 (N_11479,N_8228,N_8758);
xnor U11480 (N_11480,N_9593,N_8677);
nand U11481 (N_11481,N_9790,N_9890);
nor U11482 (N_11482,N_9937,N_9057);
and U11483 (N_11483,N_8083,N_9179);
xor U11484 (N_11484,N_9163,N_9392);
or U11485 (N_11485,N_8002,N_9021);
xnor U11486 (N_11486,N_9588,N_9461);
nand U11487 (N_11487,N_8946,N_8995);
xnor U11488 (N_11488,N_8916,N_8481);
nor U11489 (N_11489,N_9690,N_9460);
xnor U11490 (N_11490,N_8815,N_8555);
xor U11491 (N_11491,N_9916,N_9873);
and U11492 (N_11492,N_9644,N_9461);
nor U11493 (N_11493,N_8415,N_8663);
nand U11494 (N_11494,N_8000,N_8539);
xnor U11495 (N_11495,N_9843,N_9083);
nand U11496 (N_11496,N_8559,N_8414);
nand U11497 (N_11497,N_8353,N_8326);
nand U11498 (N_11498,N_8622,N_8674);
nor U11499 (N_11499,N_8800,N_8915);
nand U11500 (N_11500,N_8214,N_8543);
nor U11501 (N_11501,N_8543,N_8444);
nand U11502 (N_11502,N_9233,N_8637);
and U11503 (N_11503,N_9434,N_8889);
and U11504 (N_11504,N_9537,N_9076);
or U11505 (N_11505,N_8175,N_8731);
or U11506 (N_11506,N_9098,N_8208);
or U11507 (N_11507,N_8801,N_8454);
and U11508 (N_11508,N_9111,N_8157);
nor U11509 (N_11509,N_8325,N_9467);
xnor U11510 (N_11510,N_9099,N_8645);
nand U11511 (N_11511,N_9358,N_9396);
or U11512 (N_11512,N_9061,N_9833);
xor U11513 (N_11513,N_9372,N_9441);
or U11514 (N_11514,N_9257,N_9581);
xor U11515 (N_11515,N_9304,N_8048);
and U11516 (N_11516,N_8538,N_8589);
nand U11517 (N_11517,N_9969,N_8362);
xnor U11518 (N_11518,N_8631,N_8431);
nand U11519 (N_11519,N_9519,N_9874);
xor U11520 (N_11520,N_8928,N_8684);
or U11521 (N_11521,N_8017,N_9038);
and U11522 (N_11522,N_9083,N_8845);
and U11523 (N_11523,N_8809,N_9535);
xor U11524 (N_11524,N_8978,N_8189);
or U11525 (N_11525,N_9650,N_8806);
or U11526 (N_11526,N_8086,N_8028);
nand U11527 (N_11527,N_8455,N_8632);
xnor U11528 (N_11528,N_8519,N_9412);
and U11529 (N_11529,N_9454,N_9216);
nand U11530 (N_11530,N_8967,N_9301);
or U11531 (N_11531,N_8056,N_8459);
or U11532 (N_11532,N_9140,N_9418);
nand U11533 (N_11533,N_8512,N_8308);
xor U11534 (N_11534,N_9812,N_8514);
nor U11535 (N_11535,N_9253,N_9541);
xnor U11536 (N_11536,N_9663,N_9147);
xnor U11537 (N_11537,N_9492,N_8361);
nand U11538 (N_11538,N_8867,N_9330);
xnor U11539 (N_11539,N_9095,N_9537);
nor U11540 (N_11540,N_8710,N_8121);
or U11541 (N_11541,N_8788,N_8518);
and U11542 (N_11542,N_8424,N_9575);
nand U11543 (N_11543,N_9085,N_8859);
nand U11544 (N_11544,N_8152,N_9335);
nand U11545 (N_11545,N_9115,N_8272);
nand U11546 (N_11546,N_8199,N_8015);
xnor U11547 (N_11547,N_9512,N_8119);
nand U11548 (N_11548,N_8558,N_9189);
or U11549 (N_11549,N_8230,N_8925);
or U11550 (N_11550,N_8677,N_8924);
nor U11551 (N_11551,N_9610,N_8908);
nor U11552 (N_11552,N_8757,N_8177);
xor U11553 (N_11553,N_8053,N_8447);
and U11554 (N_11554,N_8682,N_9508);
xnor U11555 (N_11555,N_9108,N_9791);
xnor U11556 (N_11556,N_9889,N_8644);
or U11557 (N_11557,N_9153,N_9733);
and U11558 (N_11558,N_8978,N_9716);
xnor U11559 (N_11559,N_8532,N_9451);
and U11560 (N_11560,N_8270,N_9526);
or U11561 (N_11561,N_8322,N_8190);
nor U11562 (N_11562,N_8873,N_8735);
nor U11563 (N_11563,N_9653,N_9850);
or U11564 (N_11564,N_9988,N_9926);
or U11565 (N_11565,N_8313,N_8379);
nand U11566 (N_11566,N_9537,N_8277);
xor U11567 (N_11567,N_8501,N_8025);
and U11568 (N_11568,N_8212,N_8712);
nand U11569 (N_11569,N_8280,N_8521);
nand U11570 (N_11570,N_9679,N_8158);
xor U11571 (N_11571,N_9829,N_8402);
nand U11572 (N_11572,N_9956,N_9112);
xnor U11573 (N_11573,N_9913,N_9665);
or U11574 (N_11574,N_9458,N_9388);
xnor U11575 (N_11575,N_8384,N_9977);
or U11576 (N_11576,N_9191,N_8196);
xnor U11577 (N_11577,N_8965,N_8503);
nand U11578 (N_11578,N_8263,N_8483);
nor U11579 (N_11579,N_8887,N_8576);
or U11580 (N_11580,N_8343,N_8921);
nand U11581 (N_11581,N_9112,N_9337);
and U11582 (N_11582,N_9527,N_9102);
xnor U11583 (N_11583,N_8330,N_9913);
xnor U11584 (N_11584,N_9931,N_8156);
and U11585 (N_11585,N_8001,N_9353);
or U11586 (N_11586,N_9707,N_8428);
nor U11587 (N_11587,N_8167,N_8694);
xor U11588 (N_11588,N_9321,N_8018);
nand U11589 (N_11589,N_8212,N_8356);
or U11590 (N_11590,N_9426,N_9845);
nand U11591 (N_11591,N_9607,N_9126);
nor U11592 (N_11592,N_9376,N_9904);
nand U11593 (N_11593,N_8978,N_9655);
xor U11594 (N_11594,N_8375,N_9690);
xor U11595 (N_11595,N_8340,N_9009);
nor U11596 (N_11596,N_8442,N_9268);
and U11597 (N_11597,N_8519,N_9910);
and U11598 (N_11598,N_9780,N_9175);
or U11599 (N_11599,N_8540,N_8727);
nand U11600 (N_11600,N_8555,N_9823);
nand U11601 (N_11601,N_9138,N_9370);
or U11602 (N_11602,N_9129,N_9930);
and U11603 (N_11603,N_8486,N_8796);
nand U11604 (N_11604,N_8540,N_8378);
xor U11605 (N_11605,N_9396,N_8920);
nor U11606 (N_11606,N_8817,N_9645);
nor U11607 (N_11607,N_8425,N_8159);
xor U11608 (N_11608,N_9645,N_8775);
or U11609 (N_11609,N_8937,N_8117);
and U11610 (N_11610,N_9364,N_8217);
xor U11611 (N_11611,N_9545,N_9015);
xor U11612 (N_11612,N_9739,N_9523);
or U11613 (N_11613,N_8871,N_9203);
xor U11614 (N_11614,N_9864,N_8654);
xor U11615 (N_11615,N_8679,N_8683);
nor U11616 (N_11616,N_9411,N_8753);
or U11617 (N_11617,N_8357,N_9641);
or U11618 (N_11618,N_8352,N_8757);
and U11619 (N_11619,N_9946,N_9309);
xnor U11620 (N_11620,N_8863,N_9750);
nor U11621 (N_11621,N_8397,N_9997);
nand U11622 (N_11622,N_8614,N_8019);
nand U11623 (N_11623,N_9444,N_9684);
or U11624 (N_11624,N_9513,N_9901);
or U11625 (N_11625,N_8034,N_8864);
xnor U11626 (N_11626,N_9849,N_8440);
and U11627 (N_11627,N_8222,N_8675);
and U11628 (N_11628,N_9598,N_9250);
nor U11629 (N_11629,N_8050,N_9965);
nor U11630 (N_11630,N_8664,N_8987);
xnor U11631 (N_11631,N_8516,N_8042);
or U11632 (N_11632,N_9680,N_8556);
and U11633 (N_11633,N_8693,N_9811);
xnor U11634 (N_11634,N_8405,N_8035);
and U11635 (N_11635,N_8077,N_8500);
nand U11636 (N_11636,N_9470,N_8946);
nor U11637 (N_11637,N_9883,N_8859);
or U11638 (N_11638,N_8653,N_8066);
or U11639 (N_11639,N_8174,N_8062);
and U11640 (N_11640,N_8050,N_9548);
or U11641 (N_11641,N_9604,N_8411);
and U11642 (N_11642,N_9462,N_9247);
or U11643 (N_11643,N_9712,N_9776);
xnor U11644 (N_11644,N_9998,N_9081);
or U11645 (N_11645,N_8132,N_9481);
or U11646 (N_11646,N_8755,N_9765);
nor U11647 (N_11647,N_8576,N_9357);
or U11648 (N_11648,N_8560,N_8405);
nand U11649 (N_11649,N_9144,N_8821);
or U11650 (N_11650,N_9739,N_8745);
xnor U11651 (N_11651,N_8036,N_8863);
and U11652 (N_11652,N_8075,N_8071);
and U11653 (N_11653,N_9667,N_9017);
xor U11654 (N_11654,N_8016,N_8052);
nand U11655 (N_11655,N_9195,N_9927);
nand U11656 (N_11656,N_9589,N_8344);
and U11657 (N_11657,N_9443,N_8893);
xor U11658 (N_11658,N_8144,N_9471);
or U11659 (N_11659,N_9676,N_9524);
xor U11660 (N_11660,N_8469,N_9839);
and U11661 (N_11661,N_8238,N_9892);
xor U11662 (N_11662,N_8769,N_9742);
nor U11663 (N_11663,N_9118,N_9700);
nand U11664 (N_11664,N_8097,N_9719);
nor U11665 (N_11665,N_9531,N_8150);
nand U11666 (N_11666,N_8361,N_8862);
xor U11667 (N_11667,N_8290,N_9028);
and U11668 (N_11668,N_8201,N_8175);
nor U11669 (N_11669,N_9871,N_9813);
nand U11670 (N_11670,N_8919,N_9994);
nand U11671 (N_11671,N_9135,N_8270);
and U11672 (N_11672,N_9355,N_9542);
xnor U11673 (N_11673,N_9502,N_8490);
or U11674 (N_11674,N_8646,N_8128);
xor U11675 (N_11675,N_8729,N_8000);
xor U11676 (N_11676,N_8953,N_8025);
or U11677 (N_11677,N_9418,N_8997);
nand U11678 (N_11678,N_9450,N_9238);
or U11679 (N_11679,N_9400,N_9252);
and U11680 (N_11680,N_9582,N_8057);
xor U11681 (N_11681,N_8539,N_8055);
nand U11682 (N_11682,N_9897,N_9413);
or U11683 (N_11683,N_8605,N_8757);
nor U11684 (N_11684,N_8922,N_8832);
and U11685 (N_11685,N_8058,N_9080);
nor U11686 (N_11686,N_9858,N_9377);
and U11687 (N_11687,N_8610,N_8272);
or U11688 (N_11688,N_8349,N_9406);
nor U11689 (N_11689,N_8844,N_8796);
and U11690 (N_11690,N_8727,N_9450);
xnor U11691 (N_11691,N_8782,N_9860);
or U11692 (N_11692,N_8081,N_8642);
nand U11693 (N_11693,N_8820,N_8445);
nor U11694 (N_11694,N_9423,N_9368);
or U11695 (N_11695,N_9895,N_8066);
xnor U11696 (N_11696,N_8716,N_9559);
xnor U11697 (N_11697,N_8072,N_8253);
nand U11698 (N_11698,N_9427,N_8240);
nand U11699 (N_11699,N_9790,N_9861);
or U11700 (N_11700,N_8474,N_8366);
nor U11701 (N_11701,N_9675,N_8909);
xnor U11702 (N_11702,N_9990,N_9179);
xor U11703 (N_11703,N_8800,N_8214);
nand U11704 (N_11704,N_8409,N_8183);
xor U11705 (N_11705,N_9823,N_8641);
nand U11706 (N_11706,N_8766,N_9255);
or U11707 (N_11707,N_8664,N_9569);
nor U11708 (N_11708,N_9308,N_8770);
and U11709 (N_11709,N_9226,N_8783);
nor U11710 (N_11710,N_8653,N_9955);
nand U11711 (N_11711,N_9831,N_8821);
nand U11712 (N_11712,N_8485,N_9125);
nor U11713 (N_11713,N_9379,N_8828);
nor U11714 (N_11714,N_9702,N_9679);
or U11715 (N_11715,N_9331,N_9540);
nand U11716 (N_11716,N_9991,N_9277);
nor U11717 (N_11717,N_8275,N_8162);
or U11718 (N_11718,N_9841,N_9165);
nor U11719 (N_11719,N_9602,N_9259);
nand U11720 (N_11720,N_9168,N_9955);
or U11721 (N_11721,N_8916,N_9861);
xor U11722 (N_11722,N_9585,N_9331);
nor U11723 (N_11723,N_9083,N_8989);
nor U11724 (N_11724,N_8060,N_8045);
xnor U11725 (N_11725,N_9848,N_8936);
xor U11726 (N_11726,N_8534,N_8098);
and U11727 (N_11727,N_9815,N_9500);
xnor U11728 (N_11728,N_8791,N_9294);
or U11729 (N_11729,N_8221,N_9293);
nand U11730 (N_11730,N_8811,N_8275);
and U11731 (N_11731,N_9873,N_8666);
nor U11732 (N_11732,N_8470,N_9303);
nor U11733 (N_11733,N_8579,N_8173);
nor U11734 (N_11734,N_9857,N_8847);
and U11735 (N_11735,N_9450,N_8293);
and U11736 (N_11736,N_9316,N_8677);
and U11737 (N_11737,N_9764,N_9275);
or U11738 (N_11738,N_9513,N_8038);
or U11739 (N_11739,N_9375,N_8044);
nand U11740 (N_11740,N_9838,N_8761);
nand U11741 (N_11741,N_8157,N_9542);
xor U11742 (N_11742,N_9179,N_8676);
nand U11743 (N_11743,N_9990,N_8495);
and U11744 (N_11744,N_8533,N_9510);
or U11745 (N_11745,N_9937,N_8853);
nand U11746 (N_11746,N_9235,N_9423);
or U11747 (N_11747,N_9218,N_9651);
nor U11748 (N_11748,N_9563,N_9130);
nor U11749 (N_11749,N_9012,N_8504);
nor U11750 (N_11750,N_8281,N_9148);
and U11751 (N_11751,N_9775,N_8175);
or U11752 (N_11752,N_9279,N_9818);
and U11753 (N_11753,N_8197,N_9016);
and U11754 (N_11754,N_9816,N_8802);
and U11755 (N_11755,N_9968,N_9006);
xnor U11756 (N_11756,N_8525,N_8937);
nand U11757 (N_11757,N_8637,N_8402);
and U11758 (N_11758,N_9735,N_9585);
or U11759 (N_11759,N_9384,N_9085);
and U11760 (N_11760,N_8765,N_8278);
or U11761 (N_11761,N_8835,N_9024);
and U11762 (N_11762,N_9988,N_9184);
and U11763 (N_11763,N_9118,N_9990);
or U11764 (N_11764,N_9613,N_8193);
nand U11765 (N_11765,N_8667,N_8183);
nand U11766 (N_11766,N_8195,N_8961);
nand U11767 (N_11767,N_8811,N_9878);
nand U11768 (N_11768,N_8347,N_9158);
and U11769 (N_11769,N_8681,N_8676);
nand U11770 (N_11770,N_8519,N_9475);
xor U11771 (N_11771,N_9009,N_9700);
and U11772 (N_11772,N_9258,N_8885);
or U11773 (N_11773,N_9909,N_8161);
nor U11774 (N_11774,N_9252,N_8988);
or U11775 (N_11775,N_8861,N_8639);
or U11776 (N_11776,N_8793,N_9308);
nor U11777 (N_11777,N_9053,N_8189);
nor U11778 (N_11778,N_9996,N_9433);
or U11779 (N_11779,N_8861,N_9774);
and U11780 (N_11780,N_8888,N_9919);
xnor U11781 (N_11781,N_9274,N_9352);
xnor U11782 (N_11782,N_9898,N_9440);
xnor U11783 (N_11783,N_8689,N_9427);
nor U11784 (N_11784,N_8783,N_9146);
xor U11785 (N_11785,N_9802,N_8283);
nor U11786 (N_11786,N_8386,N_8613);
or U11787 (N_11787,N_9136,N_9249);
nor U11788 (N_11788,N_9131,N_9145);
nand U11789 (N_11789,N_9071,N_9763);
nand U11790 (N_11790,N_8311,N_9683);
xor U11791 (N_11791,N_9011,N_9455);
nand U11792 (N_11792,N_8628,N_9444);
nor U11793 (N_11793,N_8881,N_9234);
xnor U11794 (N_11794,N_9957,N_8636);
or U11795 (N_11795,N_8382,N_9179);
xnor U11796 (N_11796,N_9486,N_8125);
xnor U11797 (N_11797,N_8030,N_9994);
nor U11798 (N_11798,N_9790,N_9959);
or U11799 (N_11799,N_9217,N_9809);
nand U11800 (N_11800,N_8764,N_9589);
xor U11801 (N_11801,N_9186,N_8054);
nor U11802 (N_11802,N_9564,N_8790);
nor U11803 (N_11803,N_9626,N_8325);
or U11804 (N_11804,N_8744,N_8622);
xnor U11805 (N_11805,N_9943,N_8626);
and U11806 (N_11806,N_9738,N_9884);
or U11807 (N_11807,N_8468,N_9037);
nand U11808 (N_11808,N_9058,N_8401);
and U11809 (N_11809,N_8750,N_9409);
xnor U11810 (N_11810,N_9669,N_9991);
nand U11811 (N_11811,N_8033,N_8928);
and U11812 (N_11812,N_8923,N_9618);
nor U11813 (N_11813,N_9489,N_8964);
nor U11814 (N_11814,N_9981,N_9452);
and U11815 (N_11815,N_9552,N_9541);
xor U11816 (N_11816,N_9200,N_8233);
nor U11817 (N_11817,N_9016,N_8795);
nand U11818 (N_11818,N_8019,N_9413);
and U11819 (N_11819,N_9638,N_8261);
nor U11820 (N_11820,N_9586,N_8279);
nor U11821 (N_11821,N_8978,N_8311);
or U11822 (N_11822,N_9252,N_8592);
or U11823 (N_11823,N_8234,N_8257);
xnor U11824 (N_11824,N_9465,N_9119);
or U11825 (N_11825,N_9318,N_9407);
and U11826 (N_11826,N_8536,N_8699);
xnor U11827 (N_11827,N_9752,N_8080);
or U11828 (N_11828,N_8022,N_8740);
nor U11829 (N_11829,N_8196,N_9094);
nor U11830 (N_11830,N_8172,N_8178);
nand U11831 (N_11831,N_9815,N_9045);
or U11832 (N_11832,N_9607,N_9898);
xor U11833 (N_11833,N_8423,N_8027);
nor U11834 (N_11834,N_8120,N_9816);
nand U11835 (N_11835,N_8502,N_9056);
xnor U11836 (N_11836,N_8718,N_9970);
and U11837 (N_11837,N_9113,N_8574);
and U11838 (N_11838,N_9876,N_8071);
nor U11839 (N_11839,N_8800,N_8743);
or U11840 (N_11840,N_9809,N_8543);
and U11841 (N_11841,N_8530,N_9270);
and U11842 (N_11842,N_8946,N_9561);
and U11843 (N_11843,N_8108,N_9691);
xnor U11844 (N_11844,N_8550,N_9189);
nor U11845 (N_11845,N_9421,N_9521);
and U11846 (N_11846,N_8184,N_9833);
xor U11847 (N_11847,N_9927,N_9531);
xor U11848 (N_11848,N_9772,N_9074);
or U11849 (N_11849,N_8395,N_8235);
or U11850 (N_11850,N_9658,N_9937);
or U11851 (N_11851,N_8728,N_8357);
and U11852 (N_11852,N_9785,N_9413);
xnor U11853 (N_11853,N_8901,N_9054);
or U11854 (N_11854,N_8105,N_8536);
nand U11855 (N_11855,N_8347,N_8016);
xnor U11856 (N_11856,N_9130,N_8628);
xor U11857 (N_11857,N_8971,N_8052);
and U11858 (N_11858,N_9237,N_9530);
or U11859 (N_11859,N_9638,N_8160);
xor U11860 (N_11860,N_9494,N_9516);
nor U11861 (N_11861,N_9965,N_9175);
or U11862 (N_11862,N_9162,N_8396);
nor U11863 (N_11863,N_8035,N_9190);
or U11864 (N_11864,N_9167,N_9418);
nand U11865 (N_11865,N_9971,N_9979);
nand U11866 (N_11866,N_9140,N_8174);
and U11867 (N_11867,N_8502,N_8984);
xor U11868 (N_11868,N_9504,N_8455);
nor U11869 (N_11869,N_9245,N_9269);
or U11870 (N_11870,N_8376,N_8321);
xnor U11871 (N_11871,N_8778,N_9826);
nand U11872 (N_11872,N_8215,N_8270);
xor U11873 (N_11873,N_9400,N_9016);
or U11874 (N_11874,N_8470,N_9585);
or U11875 (N_11875,N_8879,N_9578);
nor U11876 (N_11876,N_8020,N_8358);
nor U11877 (N_11877,N_8743,N_8948);
and U11878 (N_11878,N_8911,N_8661);
nor U11879 (N_11879,N_9242,N_8665);
and U11880 (N_11880,N_9892,N_9679);
or U11881 (N_11881,N_8881,N_8308);
and U11882 (N_11882,N_9400,N_8780);
xnor U11883 (N_11883,N_8948,N_9178);
and U11884 (N_11884,N_8041,N_9179);
nor U11885 (N_11885,N_9990,N_9768);
nor U11886 (N_11886,N_8928,N_8597);
and U11887 (N_11887,N_9779,N_9830);
or U11888 (N_11888,N_9409,N_8517);
and U11889 (N_11889,N_8305,N_8000);
nor U11890 (N_11890,N_9423,N_9146);
xnor U11891 (N_11891,N_8288,N_9252);
or U11892 (N_11892,N_9265,N_9266);
or U11893 (N_11893,N_9040,N_8282);
xnor U11894 (N_11894,N_8085,N_8819);
or U11895 (N_11895,N_8078,N_8624);
and U11896 (N_11896,N_8151,N_9256);
nand U11897 (N_11897,N_9622,N_8225);
or U11898 (N_11898,N_8660,N_8901);
nand U11899 (N_11899,N_8051,N_9265);
nand U11900 (N_11900,N_8308,N_8156);
nor U11901 (N_11901,N_8442,N_8274);
or U11902 (N_11902,N_8016,N_8054);
nand U11903 (N_11903,N_9497,N_9994);
xor U11904 (N_11904,N_8183,N_9855);
and U11905 (N_11905,N_9316,N_8200);
or U11906 (N_11906,N_9292,N_8552);
nand U11907 (N_11907,N_9679,N_9677);
xor U11908 (N_11908,N_9523,N_8380);
nor U11909 (N_11909,N_8453,N_8688);
nand U11910 (N_11910,N_8097,N_8748);
nor U11911 (N_11911,N_9181,N_8324);
and U11912 (N_11912,N_9359,N_9361);
xor U11913 (N_11913,N_8740,N_9304);
nand U11914 (N_11914,N_8953,N_8129);
nand U11915 (N_11915,N_9743,N_8071);
nand U11916 (N_11916,N_9512,N_9002);
and U11917 (N_11917,N_9192,N_9688);
or U11918 (N_11918,N_8426,N_9487);
xnor U11919 (N_11919,N_8861,N_8687);
and U11920 (N_11920,N_9546,N_9285);
nor U11921 (N_11921,N_9686,N_8144);
and U11922 (N_11922,N_8950,N_8784);
or U11923 (N_11923,N_9235,N_8011);
xnor U11924 (N_11924,N_8529,N_9016);
nor U11925 (N_11925,N_9951,N_8685);
xor U11926 (N_11926,N_8824,N_8778);
nor U11927 (N_11927,N_8403,N_9825);
or U11928 (N_11928,N_8247,N_9639);
nor U11929 (N_11929,N_8915,N_9363);
and U11930 (N_11930,N_9691,N_9304);
or U11931 (N_11931,N_9396,N_8341);
nand U11932 (N_11932,N_9126,N_9979);
xor U11933 (N_11933,N_8898,N_9011);
or U11934 (N_11934,N_8791,N_8958);
and U11935 (N_11935,N_8116,N_8877);
or U11936 (N_11936,N_9038,N_8673);
and U11937 (N_11937,N_9148,N_9171);
nand U11938 (N_11938,N_9347,N_9595);
xnor U11939 (N_11939,N_8927,N_9700);
or U11940 (N_11940,N_9830,N_9974);
and U11941 (N_11941,N_9059,N_9353);
nor U11942 (N_11942,N_9957,N_8969);
or U11943 (N_11943,N_8676,N_8289);
and U11944 (N_11944,N_8000,N_8269);
nand U11945 (N_11945,N_9043,N_8982);
nand U11946 (N_11946,N_8332,N_8357);
nor U11947 (N_11947,N_9729,N_8979);
nor U11948 (N_11948,N_9210,N_9447);
nor U11949 (N_11949,N_9687,N_8645);
nor U11950 (N_11950,N_9332,N_8043);
and U11951 (N_11951,N_8295,N_9453);
nor U11952 (N_11952,N_9086,N_8520);
xnor U11953 (N_11953,N_8876,N_9436);
nand U11954 (N_11954,N_8171,N_9594);
nor U11955 (N_11955,N_8683,N_9455);
or U11956 (N_11956,N_8286,N_9732);
and U11957 (N_11957,N_9799,N_9096);
and U11958 (N_11958,N_9670,N_9450);
and U11959 (N_11959,N_9936,N_8197);
nor U11960 (N_11960,N_9349,N_8350);
nand U11961 (N_11961,N_9108,N_9422);
or U11962 (N_11962,N_8258,N_8459);
or U11963 (N_11963,N_9530,N_9151);
nor U11964 (N_11964,N_9379,N_9294);
nor U11965 (N_11965,N_8941,N_9802);
nand U11966 (N_11966,N_9808,N_8179);
xnor U11967 (N_11967,N_8489,N_9629);
or U11968 (N_11968,N_8067,N_8338);
and U11969 (N_11969,N_9951,N_9889);
nand U11970 (N_11970,N_8842,N_9567);
nor U11971 (N_11971,N_8283,N_8435);
nand U11972 (N_11972,N_9876,N_9279);
xnor U11973 (N_11973,N_9310,N_9129);
or U11974 (N_11974,N_8055,N_9967);
nand U11975 (N_11975,N_9052,N_9590);
nand U11976 (N_11976,N_8167,N_8359);
or U11977 (N_11977,N_9397,N_9621);
or U11978 (N_11978,N_9079,N_9878);
nand U11979 (N_11979,N_9869,N_8416);
and U11980 (N_11980,N_9821,N_8308);
nor U11981 (N_11981,N_8896,N_8434);
nand U11982 (N_11982,N_8087,N_8846);
nand U11983 (N_11983,N_8306,N_8843);
nand U11984 (N_11984,N_9054,N_9934);
and U11985 (N_11985,N_8963,N_9296);
xnor U11986 (N_11986,N_8684,N_8094);
nor U11987 (N_11987,N_9757,N_8994);
xnor U11988 (N_11988,N_9472,N_9214);
or U11989 (N_11989,N_9766,N_9699);
and U11990 (N_11990,N_8908,N_9873);
and U11991 (N_11991,N_8914,N_8575);
nand U11992 (N_11992,N_8546,N_9504);
nand U11993 (N_11993,N_9314,N_8543);
xnor U11994 (N_11994,N_9127,N_8117);
nor U11995 (N_11995,N_8713,N_9268);
xnor U11996 (N_11996,N_9900,N_9567);
or U11997 (N_11997,N_8674,N_8722);
nor U11998 (N_11998,N_9568,N_8567);
nand U11999 (N_11999,N_8469,N_9425);
or U12000 (N_12000,N_11157,N_11924);
xor U12001 (N_12001,N_10095,N_10931);
xnor U12002 (N_12002,N_11758,N_10282);
nand U12003 (N_12003,N_11147,N_11543);
nand U12004 (N_12004,N_10425,N_11304);
xnor U12005 (N_12005,N_11876,N_11711);
and U12006 (N_12006,N_10779,N_10768);
nor U12007 (N_12007,N_10819,N_10423);
xnor U12008 (N_12008,N_10316,N_11978);
xor U12009 (N_12009,N_10939,N_10869);
nor U12010 (N_12010,N_10688,N_10146);
nor U12011 (N_12011,N_10693,N_11313);
nor U12012 (N_12012,N_11700,N_11937);
xnor U12013 (N_12013,N_11424,N_10786);
xnor U12014 (N_12014,N_11547,N_10604);
nand U12015 (N_12015,N_10626,N_11176);
xnor U12016 (N_12016,N_11976,N_11838);
nor U12017 (N_12017,N_10789,N_10589);
xnor U12018 (N_12018,N_11315,N_11303);
or U12019 (N_12019,N_11829,N_11845);
nor U12020 (N_12020,N_11423,N_10974);
or U12021 (N_12021,N_10962,N_10635);
nor U12022 (N_12022,N_10273,N_10806);
nand U12023 (N_12023,N_11098,N_11478);
nor U12024 (N_12024,N_11030,N_10812);
or U12025 (N_12025,N_10992,N_11609);
xnor U12026 (N_12026,N_10845,N_11942);
nand U12027 (N_12027,N_11750,N_10192);
and U12028 (N_12028,N_10526,N_11379);
xor U12029 (N_12029,N_10313,N_10734);
nor U12030 (N_12030,N_10096,N_11902);
or U12031 (N_12031,N_11244,N_10361);
nand U12032 (N_12032,N_10994,N_11367);
or U12033 (N_12033,N_11742,N_10108);
nor U12034 (N_12034,N_11192,N_11506);
and U12035 (N_12035,N_11767,N_11272);
xnor U12036 (N_12036,N_10385,N_11975);
nand U12037 (N_12037,N_11327,N_11910);
nor U12038 (N_12038,N_10023,N_11453);
or U12039 (N_12039,N_10272,N_11687);
nor U12040 (N_12040,N_11649,N_11065);
nor U12041 (N_12041,N_10623,N_10215);
xnor U12042 (N_12042,N_11961,N_10340);
xnor U12043 (N_12043,N_10548,N_11761);
nor U12044 (N_12044,N_10290,N_10824);
or U12045 (N_12045,N_11685,N_10403);
or U12046 (N_12046,N_10762,N_10190);
nand U12047 (N_12047,N_10339,N_11029);
nand U12048 (N_12048,N_10102,N_11209);
xnor U12049 (N_12049,N_11677,N_10666);
xor U12050 (N_12050,N_10119,N_11397);
nor U12051 (N_12051,N_11476,N_10266);
or U12052 (N_12052,N_11214,N_10223);
nand U12053 (N_12053,N_10764,N_11222);
or U12054 (N_12054,N_10249,N_10797);
nor U12055 (N_12055,N_11593,N_11396);
or U12056 (N_12056,N_11336,N_10694);
nand U12057 (N_12057,N_10957,N_11915);
nor U12058 (N_12058,N_10835,N_10245);
nor U12059 (N_12059,N_10205,N_11469);
and U12060 (N_12060,N_10391,N_11159);
and U12061 (N_12061,N_11969,N_10871);
xnor U12062 (N_12062,N_11354,N_11884);
nor U12063 (N_12063,N_11046,N_11300);
nand U12064 (N_12064,N_10073,N_10438);
xnor U12065 (N_12065,N_11514,N_11095);
nor U12066 (N_12066,N_11950,N_10528);
nand U12067 (N_12067,N_10332,N_11972);
xnor U12068 (N_12068,N_11109,N_10236);
nor U12069 (N_12069,N_10879,N_11001);
or U12070 (N_12070,N_11979,N_11099);
xnor U12071 (N_12071,N_10706,N_10109);
or U12072 (N_12072,N_10222,N_10252);
and U12073 (N_12073,N_10996,N_10759);
nor U12074 (N_12074,N_11253,N_10043);
or U12075 (N_12075,N_10560,N_10349);
or U12076 (N_12076,N_10711,N_11306);
xnor U12077 (N_12077,N_11079,N_11971);
and U12078 (N_12078,N_10959,N_11289);
and U12079 (N_12079,N_11102,N_11734);
nor U12080 (N_12080,N_10207,N_11169);
nor U12081 (N_12081,N_10611,N_10941);
nand U12082 (N_12082,N_11994,N_11977);
and U12083 (N_12083,N_10794,N_11509);
nand U12084 (N_12084,N_11954,N_11682);
nor U12085 (N_12085,N_11923,N_11404);
or U12086 (N_12086,N_10322,N_11556);
xnor U12087 (N_12087,N_11648,N_11513);
xnor U12088 (N_12088,N_10531,N_11817);
nor U12089 (N_12089,N_11004,N_11066);
or U12090 (N_12090,N_11140,N_11533);
nand U12091 (N_12091,N_10174,N_10851);
nor U12092 (N_12092,N_10828,N_11394);
or U12093 (N_12093,N_10659,N_10866);
and U12094 (N_12094,N_11588,N_10596);
and U12095 (N_12095,N_11285,N_11550);
nand U12096 (N_12096,N_10757,N_11167);
nand U12097 (N_12097,N_11049,N_10776);
nand U12098 (N_12098,N_10480,N_11803);
nand U12099 (N_12099,N_11365,N_10540);
xnor U12100 (N_12100,N_11928,N_11026);
and U12101 (N_12101,N_11230,N_11567);
nand U12102 (N_12102,N_10088,N_10750);
nand U12103 (N_12103,N_10612,N_10760);
nand U12104 (N_12104,N_10907,N_11097);
and U12105 (N_12105,N_11843,N_11060);
xor U12106 (N_12106,N_10614,N_10294);
or U12107 (N_12107,N_11538,N_11265);
and U12108 (N_12108,N_10892,N_10360);
or U12109 (N_12109,N_10353,N_10581);
nand U12110 (N_12110,N_11481,N_11431);
nand U12111 (N_12111,N_11105,N_11227);
xnor U12112 (N_12112,N_10297,N_10124);
xor U12113 (N_12113,N_11589,N_10695);
nand U12114 (N_12114,N_11773,N_11061);
or U12115 (N_12115,N_10747,N_11717);
and U12116 (N_12116,N_10071,N_11670);
and U12117 (N_12117,N_10004,N_11186);
nor U12118 (N_12118,N_11775,N_11744);
and U12119 (N_12119,N_10140,N_10860);
nand U12120 (N_12120,N_10191,N_10459);
nand U12121 (N_12121,N_11467,N_11395);
nor U12122 (N_12122,N_10737,N_11881);
and U12123 (N_12123,N_10868,N_10795);
nand U12124 (N_12124,N_11247,N_11207);
xor U12125 (N_12125,N_10769,N_10479);
nor U12126 (N_12126,N_10415,N_11319);
nor U12127 (N_12127,N_11444,N_11410);
nor U12128 (N_12128,N_10699,N_10705);
or U12129 (N_12129,N_11009,N_10743);
and U12130 (N_12130,N_11739,N_10771);
xnor U12131 (N_12131,N_10514,N_11204);
or U12132 (N_12132,N_10037,N_11804);
xnor U12133 (N_12133,N_11528,N_10638);
xnor U12134 (N_12134,N_10168,N_11993);
or U12135 (N_12135,N_10572,N_11400);
or U12136 (N_12136,N_11020,N_10450);
nand U12137 (N_12137,N_11816,N_11155);
or U12138 (N_12138,N_11032,N_11388);
or U12139 (N_12139,N_10928,N_11890);
nand U12140 (N_12140,N_10905,N_10390);
or U12141 (N_12141,N_10404,N_10110);
or U12142 (N_12142,N_10075,N_10571);
nand U12143 (N_12143,N_10656,N_10151);
nor U12144 (N_12144,N_10617,N_11715);
nand U12145 (N_12145,N_10212,N_10722);
xor U12146 (N_12146,N_10891,N_11495);
and U12147 (N_12147,N_11859,N_10251);
or U12148 (N_12148,N_10847,N_10984);
xor U12149 (N_12149,N_11196,N_10086);
or U12150 (N_12150,N_11836,N_10320);
xor U12151 (N_12151,N_10577,N_11219);
or U12152 (N_12152,N_10317,N_10723);
nand U12153 (N_12153,N_11323,N_11357);
nor U12154 (N_12154,N_11276,N_11137);
nor U12155 (N_12155,N_11943,N_11282);
and U12156 (N_12156,N_11963,N_11312);
and U12157 (N_12157,N_11248,N_10104);
nor U12158 (N_12158,N_10661,N_10053);
xnor U12159 (N_12159,N_11339,N_11027);
nand U12160 (N_12160,N_11221,N_11828);
xnor U12161 (N_12161,N_10621,N_10180);
and U12162 (N_12162,N_11091,N_10940);
and U12163 (N_12163,N_10630,N_11175);
nand U12164 (N_12164,N_11525,N_11059);
nor U12165 (N_12165,N_11008,N_11151);
and U12166 (N_12166,N_11659,N_11656);
or U12167 (N_12167,N_11755,N_10484);
and U12168 (N_12168,N_11714,N_10965);
nor U12169 (N_12169,N_11555,N_10858);
nor U12170 (N_12170,N_10001,N_11406);
nor U12171 (N_12171,N_10998,N_10502);
or U12172 (N_12172,N_11621,N_11889);
or U12173 (N_12173,N_11358,N_10232);
xnor U12174 (N_12174,N_10202,N_11895);
or U12175 (N_12175,N_10503,N_11540);
nor U12176 (N_12176,N_10886,N_11421);
xnor U12177 (N_12177,N_10123,N_11922);
nand U12178 (N_12178,N_10544,N_11238);
and U12179 (N_12179,N_10432,N_11645);
and U12180 (N_12180,N_11044,N_11047);
nor U12181 (N_12181,N_10641,N_11986);
xnor U12182 (N_12182,N_10289,N_11128);
nand U12183 (N_12183,N_11642,N_10643);
xnor U12184 (N_12184,N_10020,N_11921);
and U12185 (N_12185,N_10061,N_11661);
nand U12186 (N_12186,N_11749,N_10377);
nor U12187 (N_12187,N_10394,N_11329);
xor U12188 (N_12188,N_11662,N_11795);
and U12189 (N_12189,N_10118,N_11295);
and U12190 (N_12190,N_10523,N_10622);
xnor U12191 (N_12191,N_11366,N_10872);
and U12192 (N_12192,N_10777,N_10628);
or U12193 (N_12193,N_11628,N_11441);
or U12194 (N_12194,N_11006,N_11852);
nor U12195 (N_12195,N_11442,N_10665);
or U12196 (N_12196,N_10605,N_10285);
and U12197 (N_12197,N_11636,N_11330);
xor U12198 (N_12198,N_11402,N_10172);
xor U12199 (N_12199,N_10233,N_10591);
and U12200 (N_12200,N_11806,N_10738);
and U12201 (N_12201,N_11765,N_10983);
and U12202 (N_12202,N_11084,N_10034);
nand U12203 (N_12203,N_10700,N_11604);
xor U12204 (N_12204,N_11232,N_10530);
and U12205 (N_12205,N_10507,N_10056);
xnor U12206 (N_12206,N_10100,N_11987);
nor U12207 (N_12207,N_11624,N_10539);
and U12208 (N_12208,N_10298,N_10739);
xnor U12209 (N_12209,N_11871,N_11194);
or U12210 (N_12210,N_10896,N_10303);
nand U12211 (N_12211,N_11158,N_10167);
nor U12212 (N_12212,N_10668,N_10097);
nand U12213 (N_12213,N_10434,N_10411);
xor U12214 (N_12214,N_10427,N_10127);
nand U12215 (N_12215,N_11531,N_10400);
or U12216 (N_12216,N_10302,N_11119);
nor U12217 (N_12217,N_11800,N_11374);
nand U12218 (N_12218,N_11595,N_10068);
xnor U12219 (N_12219,N_11732,N_10890);
nor U12220 (N_12220,N_10066,N_10898);
or U12221 (N_12221,N_10836,N_11428);
nor U12222 (N_12222,N_10510,N_10966);
xnor U12223 (N_12223,N_11722,N_11055);
and U12224 (N_12224,N_10846,N_10913);
nor U12225 (N_12225,N_10923,N_10365);
nor U12226 (N_12226,N_11599,N_10970);
and U12227 (N_12227,N_10562,N_10185);
xor U12228 (N_12228,N_10359,N_11445);
and U12229 (N_12229,N_10449,N_11991);
nor U12230 (N_12230,N_11335,N_10608);
or U12231 (N_12231,N_11759,N_10454);
nor U12232 (N_12232,N_11848,N_10206);
nand U12233 (N_12233,N_10173,N_11063);
or U12234 (N_12234,N_11602,N_10052);
nor U12235 (N_12235,N_10894,N_11641);
or U12236 (N_12236,N_11252,N_10158);
xor U12237 (N_12237,N_10328,N_10569);
nor U12238 (N_12238,N_10991,N_11258);
nand U12239 (N_12239,N_10565,N_11608);
and U12240 (N_12240,N_10152,N_10187);
or U12241 (N_12241,N_10224,N_11138);
nor U12242 (N_12242,N_11663,N_11437);
and U12243 (N_12243,N_11919,N_11373);
or U12244 (N_12244,N_11139,N_11016);
or U12245 (N_12245,N_10006,N_10545);
nor U12246 (N_12246,N_10417,N_10646);
nor U12247 (N_12247,N_10463,N_11746);
xor U12248 (N_12248,N_10080,N_10935);
and U12249 (N_12249,N_11815,N_10269);
and U12250 (N_12250,N_10199,N_10128);
xnor U12251 (N_12251,N_10946,N_11764);
or U12252 (N_12252,N_10193,N_10064);
or U12253 (N_12253,N_11766,N_10798);
nand U12254 (N_12254,N_11713,N_11771);
and U12255 (N_12255,N_11107,N_10257);
nor U12256 (N_12256,N_11679,N_10519);
and U12257 (N_12257,N_10270,N_10312);
or U12258 (N_12258,N_11652,N_11712);
and U12259 (N_12259,N_10234,N_10660);
xor U12260 (N_12260,N_10163,N_10465);
xor U12261 (N_12261,N_10329,N_11302);
xnor U12262 (N_12262,N_10765,N_11945);
xor U12263 (N_12263,N_11702,N_10889);
nand U12264 (N_12264,N_11242,N_10542);
nor U12265 (N_12265,N_10363,N_11832);
or U12266 (N_12266,N_10731,N_10599);
nand U12267 (N_12267,N_11786,N_11962);
and U12268 (N_12268,N_11743,N_11703);
and U12269 (N_12269,N_11925,N_11796);
xnor U12270 (N_12270,N_10337,N_11825);
xor U12271 (N_12271,N_11484,N_10107);
nand U12272 (N_12272,N_11847,N_10262);
nand U12273 (N_12273,N_10787,N_11283);
and U12274 (N_12274,N_10586,N_10216);
or U12275 (N_12275,N_10408,N_11983);
nor U12276 (N_12276,N_11043,N_10231);
and U12277 (N_12277,N_10755,N_11607);
xor U12278 (N_12278,N_11747,N_11673);
nor U12279 (N_12279,N_10135,N_10247);
nand U12280 (N_12280,N_10585,N_11681);
nor U12281 (N_12281,N_10387,N_10116);
and U12282 (N_12282,N_10520,N_10000);
nand U12283 (N_12283,N_11637,N_11705);
and U12284 (N_12284,N_11948,N_11998);
xnor U12285 (N_12285,N_10943,N_10371);
or U12286 (N_12286,N_10547,N_11081);
nand U12287 (N_12287,N_11146,N_11532);
or U12288 (N_12288,N_11579,N_10553);
nor U12289 (N_12289,N_10239,N_11856);
nand U12290 (N_12290,N_11892,N_10632);
nor U12291 (N_12291,N_10782,N_11572);
and U12292 (N_12292,N_10876,N_11949);
nand U12293 (N_12293,N_10451,N_10942);
or U12294 (N_12294,N_10673,N_11728);
nor U12295 (N_12295,N_11777,N_10505);
or U12296 (N_12296,N_11181,N_11267);
nand U12297 (N_12297,N_11472,N_11028);
nand U12298 (N_12298,N_10308,N_10726);
or U12299 (N_12299,N_10671,N_10494);
xnor U12300 (N_12300,N_11088,N_10587);
nor U12301 (N_12301,N_10284,N_10568);
xor U12302 (N_12302,N_10022,N_10240);
nand U12303 (N_12303,N_11310,N_11344);
and U12304 (N_12304,N_10278,N_10575);
nand U12305 (N_12305,N_10573,N_11036);
nand U12306 (N_12306,N_11582,N_10336);
or U12307 (N_12307,N_10470,N_10161);
nor U12308 (N_12308,N_11570,N_10335);
or U12309 (N_12309,N_11121,N_11501);
nor U12310 (N_12310,N_10979,N_11477);
nor U12311 (N_12311,N_10951,N_10813);
and U12312 (N_12312,N_11292,N_10355);
xnor U12313 (N_12313,N_11314,N_10685);
nor U12314 (N_12314,N_11808,N_11187);
and U12315 (N_12315,N_11518,N_10477);
nand U12316 (N_12316,N_11503,N_11692);
nand U12317 (N_12317,N_11510,N_11671);
xnor U12318 (N_12318,N_11398,N_10033);
xor U12319 (N_12319,N_11855,N_11149);
nor U12320 (N_12320,N_11075,N_11970);
nor U12321 (N_12321,N_10620,N_10720);
nand U12322 (N_12322,N_10971,N_11288);
nor U12323 (N_12323,N_11311,N_11350);
and U12324 (N_12324,N_10319,N_11229);
or U12325 (N_12325,N_10143,N_10595);
xnor U12326 (N_12326,N_10352,N_10842);
nor U12327 (N_12327,N_11737,N_10198);
nand U12328 (N_12328,N_10792,N_11080);
xor U12329 (N_12329,N_10334,N_10950);
and U12330 (N_12330,N_11814,N_10330);
and U12331 (N_12331,N_10549,N_10716);
nand U12332 (N_12332,N_10713,N_10025);
xor U12333 (N_12333,N_10343,N_11507);
nand U12334 (N_12334,N_11264,N_11522);
and U12335 (N_12335,N_11240,N_10036);
nor U12336 (N_12336,N_10160,N_10535);
nor U12337 (N_12337,N_11150,N_11638);
or U12338 (N_12338,N_10537,N_11721);
and U12339 (N_12339,N_10594,N_10799);
and U12340 (N_12340,N_11658,N_11590);
and U12341 (N_12341,N_10396,N_11526);
and U12342 (N_12342,N_11130,N_10429);
xnor U12343 (N_12343,N_10578,N_11197);
or U12344 (N_12344,N_11184,N_11045);
nand U12345 (N_12345,N_10372,N_10238);
or U12346 (N_12346,N_11701,N_11529);
or U12347 (N_12347,N_10389,N_10274);
or U12348 (N_12348,N_10142,N_11015);
and U12349 (N_12349,N_11465,N_10296);
or U12350 (N_12350,N_11504,N_11408);
and U12351 (N_12351,N_11340,N_10702);
xor U12352 (N_12352,N_10949,N_10496);
xor U12353 (N_12353,N_10624,N_10730);
xnor U12354 (N_12354,N_10111,N_11752);
nor U12355 (N_12355,N_11826,N_11947);
and U12356 (N_12356,N_11573,N_10379);
or U12357 (N_12357,N_11633,N_10267);
nand U12358 (N_12358,N_10552,N_10444);
xnor U12359 (N_12359,N_10131,N_10639);
nor U12360 (N_12360,N_10501,N_11770);
xor U12361 (N_12361,N_11191,N_11818);
nor U12362 (N_12362,N_11654,N_11446);
nor U12363 (N_12363,N_10024,N_10002);
nor U12364 (N_12364,N_10684,N_11216);
nand U12365 (N_12365,N_10409,N_10839);
nand U12366 (N_12366,N_10855,N_10026);
nand U12367 (N_12367,N_11498,N_11324);
and U12368 (N_12368,N_11390,N_10556);
nor U12369 (N_12369,N_11085,N_11708);
nor U12370 (N_12370,N_10579,N_10155);
or U12371 (N_12371,N_11268,N_11941);
or U12372 (N_12372,N_10832,N_10288);
xor U12373 (N_12373,N_10165,N_11985);
nor U12374 (N_12374,N_10516,N_10376);
nand U12375 (N_12375,N_10546,N_11841);
xor U12376 (N_12376,N_10490,N_10509);
nand U12377 (N_12377,N_11564,N_11912);
nor U12378 (N_12378,N_10810,N_11762);
nand U12379 (N_12379,N_10159,N_11180);
or U12380 (N_12380,N_10933,N_10072);
nor U12381 (N_12381,N_11234,N_10341);
xnor U12382 (N_12382,N_10114,N_10783);
xnor U12383 (N_12383,N_11166,N_11486);
or U12384 (N_12384,N_11291,N_10647);
and U12385 (N_12385,N_10582,N_11988);
and U12386 (N_12386,N_10823,N_10048);
nor U12387 (N_12387,N_11603,N_11791);
nor U12388 (N_12388,N_10362,N_11792);
and U12389 (N_12389,N_11592,N_10382);
nand U12390 (N_12390,N_10597,N_10864);
nor U12391 (N_12391,N_11413,N_11464);
nor U12392 (N_12392,N_10791,N_11083);
and U12393 (N_12393,N_10144,N_10261);
and U12394 (N_12394,N_10541,N_10770);
or U12395 (N_12395,N_10197,N_10993);
nand U12396 (N_12396,N_11202,N_11041);
or U12397 (N_12397,N_10670,N_10725);
xor U12398 (N_12398,N_11290,N_11675);
and U12399 (N_12399,N_10865,N_10854);
and U12400 (N_12400,N_10050,N_11430);
or U12401 (N_12401,N_11165,N_11274);
nand U12402 (N_12402,N_11474,N_11322);
and U12403 (N_12403,N_10606,N_10976);
and U12404 (N_12404,N_11013,N_10089);
or U12405 (N_12405,N_11778,N_11647);
nor U12406 (N_12406,N_11223,N_10051);
and U12407 (N_12407,N_11886,N_10271);
xnor U12408 (N_12408,N_10076,N_10042);
and U12409 (N_12409,N_10712,N_10662);
xor U12410 (N_12410,N_10978,N_10139);
xnor U12411 (N_12411,N_11087,N_10714);
and U12412 (N_12412,N_10074,N_10990);
or U12413 (N_12413,N_10848,N_11460);
nor U12414 (N_12414,N_10914,N_11042);
or U12415 (N_12415,N_11096,N_10543);
nor U12416 (N_12416,N_11364,N_11756);
nand U12417 (N_12417,N_11519,N_11585);
nand U12418 (N_12418,N_11391,N_11414);
and U12419 (N_12419,N_11092,N_11735);
nor U12420 (N_12420,N_11280,N_11461);
nor U12421 (N_12421,N_10486,N_10276);
or U12422 (N_12422,N_11868,N_11751);
nand U12423 (N_12423,N_10602,N_10021);
nand U12424 (N_12424,N_11376,N_11776);
or U12425 (N_12425,N_10210,N_10658);
xor U12426 (N_12426,N_11035,N_10751);
and U12427 (N_12427,N_10069,N_10310);
nor U12428 (N_12428,N_11918,N_11784);
or U12429 (N_12429,N_11680,N_10259);
nand U12430 (N_12430,N_10398,N_11073);
nor U12431 (N_12431,N_10358,N_10012);
and U12432 (N_12432,N_11990,N_10081);
xnor U12433 (N_12433,N_11299,N_11823);
nand U12434 (N_12434,N_10487,N_11683);
or U12435 (N_12435,N_10164,N_11089);
xor U12436 (N_12436,N_11710,N_11014);
xor U12437 (N_12437,N_11386,N_10475);
or U12438 (N_12438,N_11611,N_11877);
and U12439 (N_12439,N_11499,N_11380);
and U12440 (N_12440,N_11862,N_11185);
nand U12441 (N_12441,N_10557,N_11309);
nor U12442 (N_12442,N_10149,N_11135);
and U12443 (N_12443,N_10669,N_10888);
nor U12444 (N_12444,N_11034,N_11141);
nand U12445 (N_12445,N_10532,N_11940);
or U12446 (N_12446,N_10478,N_11007);
and U12447 (N_12447,N_11872,N_10280);
xor U12448 (N_12448,N_11480,N_11551);
and U12449 (N_12449,N_11651,N_11368);
nor U12450 (N_12450,N_10126,N_11409);
or U12451 (N_12451,N_10129,N_10536);
or U12452 (N_12452,N_11557,N_10645);
nor U12453 (N_12453,N_10920,N_10038);
or U12454 (N_12454,N_10644,N_11057);
and U12455 (N_12455,N_11269,N_10982);
xnor U12456 (N_12456,N_10761,N_10469);
xnor U12457 (N_12457,N_10227,N_10584);
nand U12458 (N_12458,N_10137,N_11490);
or U12459 (N_12459,N_10682,N_10495);
or U12460 (N_12460,N_10837,N_11419);
xnor U12461 (N_12461,N_11050,N_10301);
nor U12462 (N_12462,N_11351,N_11783);
nand U12463 (N_12463,N_10318,N_10115);
or U12464 (N_12464,N_10452,N_10566);
or U12465 (N_12465,N_11270,N_11342);
and U12466 (N_12466,N_10679,N_11875);
nor U12467 (N_12467,N_11438,N_11415);
nor U12468 (N_12468,N_10182,N_10286);
nor U12469 (N_12469,N_11182,N_10229);
nor U12470 (N_12470,N_11716,N_11691);
xor U12471 (N_12471,N_10815,N_11577);
nand U12472 (N_12472,N_11296,N_11953);
nand U12473 (N_12473,N_11120,N_10435);
and U12474 (N_12474,N_10032,N_10281);
nand U12475 (N_12475,N_11853,N_11213);
nor U12476 (N_12476,N_10030,N_10748);
and U12477 (N_12477,N_10194,N_10347);
xor U12478 (N_12478,N_10521,N_11500);
or U12479 (N_12479,N_10058,N_10098);
or U12480 (N_12480,N_11473,N_11878);
and U12481 (N_12481,N_11596,N_10431);
or U12482 (N_12482,N_11417,N_11610);
nand U12483 (N_12483,N_11471,N_11900);
or U12484 (N_12484,N_10040,N_11173);
nand U12485 (N_12485,N_11082,N_10084);
nand U12486 (N_12486,N_11888,N_11880);
or U12487 (N_12487,N_11201,N_11846);
nor U12488 (N_12488,N_10458,N_11600);
and U12489 (N_12489,N_10652,N_11172);
xnor U12490 (N_12490,N_11443,N_11346);
xnor U12491 (N_12491,N_11866,N_10323);
or U12492 (N_12492,N_10321,N_10986);
or U12493 (N_12493,N_10255,N_10834);
nor U12494 (N_12494,N_10181,N_11479);
xnor U12495 (N_12495,N_10916,N_10356);
nor U12496 (N_12496,N_10011,N_11699);
xnor U12497 (N_12497,N_10524,N_11858);
and U12498 (N_12498,N_11174,N_10041);
or U12499 (N_12499,N_11427,N_10753);
nor U12500 (N_12500,N_11025,N_10567);
and U12501 (N_12501,N_11545,N_11226);
nand U12502 (N_12502,N_10900,N_10386);
xor U12503 (N_12503,N_11726,N_10985);
nor U12504 (N_12504,N_11553,N_10870);
nand U12505 (N_12505,N_11466,N_10518);
or U12506 (N_12506,N_10195,N_10246);
xor U12507 (N_12507,N_11831,N_10395);
nor U12508 (N_12508,N_11644,N_11523);
or U12509 (N_12509,N_11076,N_10627);
xnor U12510 (N_12510,N_10440,N_10856);
and U12511 (N_12511,N_10374,N_10456);
or U12512 (N_12512,N_10576,N_11615);
nand U12513 (N_12513,N_10844,N_10326);
nand U12514 (N_12514,N_10826,N_10250);
and U12515 (N_12515,N_11170,N_11005);
xor U12516 (N_12516,N_11134,N_10121);
nand U12517 (N_12517,N_10821,N_11781);
or U12518 (N_12518,N_10461,N_10800);
nor U12519 (N_12519,N_10258,N_10903);
nor U12520 (N_12520,N_10055,N_11362);
and U12521 (N_12521,N_10707,N_11439);
or U12522 (N_12522,N_10825,N_11799);
or U12523 (N_12523,N_10275,N_10784);
xor U12524 (N_12524,N_10925,N_11114);
nor U12525 (N_12525,N_11530,N_11021);
xor U12526 (N_12526,N_10721,N_10200);
and U12527 (N_12527,N_10367,N_11927);
and U12528 (N_12528,N_11863,N_11920);
and U12529 (N_12529,N_10369,N_10906);
and U12530 (N_12530,N_11320,N_10439);
xnor U12531 (N_12531,N_11729,N_10752);
nand U12532 (N_12532,N_11999,N_10633);
nor U12533 (N_12533,N_10176,N_10696);
and U12534 (N_12534,N_10090,N_10774);
xnor U12535 (N_12535,N_11256,N_10065);
nand U12536 (N_12536,N_11497,N_11332);
xor U12537 (N_12537,N_11904,N_11665);
or U12538 (N_12538,N_10917,N_11730);
and U12539 (N_12539,N_10392,N_11617);
nand U12540 (N_12540,N_11622,N_11597);
and U12541 (N_12541,N_11215,N_10324);
nor U12542 (N_12542,N_10915,N_11436);
and U12543 (N_12543,N_10106,N_10981);
or U12544 (N_12544,N_10674,N_11403);
or U12545 (N_12545,N_11206,N_10999);
and U12546 (N_12546,N_10989,N_11951);
or U12547 (N_12547,N_10987,N_11787);
or U12548 (N_12548,N_11676,N_11966);
xnor U12549 (N_12549,N_11782,N_10551);
or U12550 (N_12550,N_10952,N_11891);
xor U12551 (N_12551,N_11132,N_11483);
or U12552 (N_12552,N_10049,N_10263);
xor U12553 (N_12553,N_10029,N_11024);
nand U12554 (N_12554,N_10350,N_11797);
or U12555 (N_12555,N_11809,N_10555);
xor U12556 (N_12556,N_10327,N_11512);
nor U12557 (N_12557,N_10831,N_10691);
xor U12558 (N_12558,N_11505,N_10201);
nand U12559 (N_12559,N_11537,N_10863);
xor U12560 (N_12560,N_11156,N_10083);
xor U12561 (N_12561,N_11997,N_11271);
xnor U12562 (N_12562,N_10527,N_11982);
nand U12563 (N_12563,N_10945,N_10874);
xnor U12564 (N_12564,N_11040,N_11359);
nand U12565 (N_12565,N_10457,N_10746);
xor U12566 (N_12566,N_11574,N_11934);
nor U12567 (N_12567,N_11763,N_11640);
xnor U12568 (N_12568,N_11217,N_11334);
nand U12569 (N_12569,N_11392,N_11416);
or U12570 (N_12570,N_11278,N_10468);
xor U12571 (N_12571,N_10122,N_11907);
nor U12572 (N_12572,N_10592,N_11992);
or U12573 (N_12573,N_11494,N_10046);
xnor U12574 (N_12574,N_11284,N_10840);
nand U12575 (N_12575,N_11914,N_11375);
or U12576 (N_12576,N_10063,N_11152);
or U12577 (N_12577,N_10428,N_10895);
xor U12578 (N_12578,N_11581,N_10099);
or U12579 (N_12579,N_11623,N_11245);
nand U12580 (N_12580,N_11874,N_10342);
nor U12581 (N_12581,N_10663,N_11338);
xnor U12582 (N_12582,N_11606,N_10817);
nand U12583 (N_12583,N_11885,N_10057);
and U12584 (N_12584,N_10675,N_11546);
nand U12585 (N_12585,N_11697,N_10681);
or U12586 (N_12586,N_10756,N_10728);
nor U12587 (N_12587,N_10028,N_10655);
xnor U12588 (N_12588,N_11432,N_10701);
nand U12589 (N_12589,N_11801,N_10472);
or U12590 (N_12590,N_11345,N_10314);
or U12591 (N_12591,N_10132,N_10930);
or U12592 (N_12592,N_10859,N_11361);
and U12593 (N_12593,N_11405,N_10593);
or U12594 (N_12594,N_10841,N_11542);
or U12595 (N_12595,N_11451,N_11709);
or U12596 (N_12596,N_11113,N_11565);
nor U12597 (N_12597,N_10583,N_10625);
xor U12598 (N_12598,N_10710,N_11377);
and U12599 (N_12599,N_10977,N_10649);
nor U12600 (N_12600,N_11811,N_11101);
or U12601 (N_12601,N_10785,N_11093);
nor U12602 (N_12602,N_10171,N_10538);
nor U12603 (N_12603,N_10947,N_10862);
nand U12604 (N_12604,N_10960,N_11870);
xor U12605 (N_12605,N_10226,N_11189);
xor U12606 (N_12606,N_10574,N_10448);
nand U12607 (N_12607,N_11496,N_10689);
nor U12608 (N_12608,N_10513,N_10816);
or U12609 (N_12609,N_11143,N_11667);
nor U12610 (N_12610,N_10901,N_10453);
nand U12611 (N_12611,N_11321,N_10085);
and U12612 (N_12612,N_11448,N_11629);
xor U12613 (N_12613,N_11205,N_10447);
xor U12614 (N_12614,N_10506,N_11901);
nor U12615 (N_12615,N_10204,N_11154);
or U12616 (N_12616,N_11694,N_11646);
or U12617 (N_12617,N_11381,N_11887);
or U12618 (N_12618,N_11821,N_11266);
or U12619 (N_12619,N_10283,N_11297);
or U12620 (N_12620,N_11981,N_11672);
and U12621 (N_12621,N_10508,N_10969);
and U12622 (N_12622,N_10936,N_10550);
and U12623 (N_12623,N_10166,N_11929);
and U12624 (N_12624,N_11627,N_11657);
nand U12625 (N_12625,N_10062,N_10995);
nor U12626 (N_12626,N_11177,N_10443);
nand U12627 (N_12627,N_11110,N_11789);
nand U12628 (N_12628,N_11719,N_10922);
or U12629 (N_12629,N_11161,N_11179);
xnor U12630 (N_12630,N_10818,N_11864);
and U12631 (N_12631,N_10601,N_10610);
xnor U12632 (N_12632,N_10926,N_11944);
and U12633 (N_12633,N_10934,N_10039);
nand U12634 (N_12634,N_11989,N_10887);
or U12635 (N_12635,N_10932,N_11360);
or U12636 (N_12636,N_11632,N_11903);
or U12637 (N_12637,N_11980,N_11485);
or U12638 (N_12638,N_11273,N_10492);
nor U12639 (N_12639,N_11246,N_10311);
nand U12640 (N_12640,N_10878,N_11536);
xnor U12641 (N_12641,N_11562,N_10677);
or U12642 (N_12642,N_11078,N_11251);
xor U12643 (N_12643,N_11286,N_11356);
or U12644 (N_12644,N_11544,N_10489);
nor U12645 (N_12645,N_10406,N_11023);
nand U12646 (N_12646,N_10912,N_11865);
xnor U12647 (N_12647,N_11489,N_10134);
nand U12648 (N_12648,N_10838,N_11183);
and U12649 (N_12649,N_10154,N_11840);
nand U12650 (N_12650,N_11849,N_11631);
or U12651 (N_12651,N_10885,N_10580);
nor U12652 (N_12652,N_11475,N_11517);
xor U12653 (N_12653,N_11720,N_10801);
nor U12654 (N_12654,N_11793,N_11487);
or U12655 (N_12655,N_10474,N_11822);
xnor U12656 (N_12656,N_10125,N_10153);
or U12657 (N_12657,N_10220,N_11837);
nand U12658 (N_12658,N_10338,N_11974);
xor U12659 (N_12659,N_10268,N_10418);
nor U12660 (N_12660,N_11435,N_11958);
or U12661 (N_12661,N_10664,N_10893);
nand U12662 (N_12662,N_10619,N_11839);
and U12663 (N_12663,N_11349,N_11188);
nand U12664 (N_12664,N_11521,N_10007);
nand U12665 (N_12665,N_10016,N_11195);
and U12666 (N_12666,N_11372,N_10909);
or U12667 (N_12667,N_11630,N_10483);
and U12668 (N_12668,N_11779,N_11249);
nor U12669 (N_12669,N_10631,N_10598);
xor U12670 (N_12670,N_10150,N_11539);
or U12671 (N_12671,N_10758,N_11239);
or U12672 (N_12672,N_11813,N_10228);
or U12673 (N_12673,N_10802,N_10031);
or U12674 (N_12674,N_11136,N_10929);
and U12675 (N_12675,N_11854,N_11468);
nand U12676 (N_12676,N_11898,N_10958);
xor U12677 (N_12677,N_10218,N_11541);
and U12678 (N_12678,N_10875,N_10348);
or U12679 (N_12679,N_11769,N_11457);
and U12680 (N_12680,N_11401,N_10005);
nand U12681 (N_12681,N_10307,N_10412);
xnor U12682 (N_12682,N_11583,N_11869);
xnor U12683 (N_12683,N_10809,N_11690);
and U12684 (N_12684,N_11162,N_10277);
nor U12685 (N_12685,N_11810,N_10497);
and U12686 (N_12686,N_10704,N_11287);
xnor U12687 (N_12687,N_10178,N_10441);
or U12688 (N_12688,N_10749,N_11452);
and U12689 (N_12689,N_10600,N_10476);
nor U12690 (N_12690,N_11458,N_10830);
and U12691 (N_12691,N_11851,N_10130);
nor U12692 (N_12692,N_11038,N_11411);
and U12693 (N_12693,N_11163,N_10745);
nor U12694 (N_12694,N_10687,N_11873);
nor U12695 (N_12695,N_10775,N_11964);
or U12696 (N_12696,N_10708,N_10241);
nor U12697 (N_12697,N_11723,N_11011);
and U12698 (N_12698,N_11434,N_11936);
xnor U12699 (N_12699,N_10609,N_10481);
nor U12700 (N_12700,N_11301,N_10243);
or U12701 (N_12701,N_10804,N_11100);
or U12702 (N_12702,N_10189,N_10260);
and U12703 (N_12703,N_10325,N_10380);
or U12704 (N_12704,N_10157,N_10287);
nand U12705 (N_12705,N_11054,N_10117);
nor U12706 (N_12706,N_11412,N_10442);
nor U12707 (N_12707,N_10690,N_11224);
nor U12708 (N_12708,N_11605,N_11559);
and U12709 (N_12709,N_10672,N_10653);
or U12710 (N_12710,N_10333,N_11200);
nor U12711 (N_12711,N_11754,N_10402);
and U12712 (N_12712,N_10732,N_10010);
xnor U12713 (N_12713,N_11067,N_10018);
or U12714 (N_12714,N_10955,N_11598);
xnor U12715 (N_12715,N_10822,N_10735);
and U12716 (N_12716,N_11867,N_11666);
and U12717 (N_12717,N_10796,N_11785);
xor U12718 (N_12718,N_10741,N_11698);
nand U12719 (N_12719,N_10686,N_10401);
nand U12720 (N_12720,N_11171,N_11956);
nand U12721 (N_12721,N_10908,N_10615);
nand U12722 (N_12722,N_10517,N_10754);
or U12723 (N_12723,N_10375,N_11212);
or U12724 (N_12724,N_11220,N_11456);
nor U12725 (N_12725,N_11508,N_11674);
and U12726 (N_12726,N_10911,N_10667);
or U12727 (N_12727,N_10805,N_10680);
and U12728 (N_12728,N_10253,N_10345);
nor U12729 (N_12729,N_11086,N_11429);
xnor U12730 (N_12730,N_10742,N_11211);
nor U12731 (N_12731,N_11635,N_11824);
or U12732 (N_12732,N_10729,N_11706);
nand U12733 (N_12733,N_11738,N_10156);
nand U12734 (N_12734,N_11684,N_10235);
nor U12735 (N_12735,N_11462,N_10419);
nor U12736 (N_12736,N_10044,N_11516);
nand U12737 (N_12737,N_10522,N_11352);
xor U12738 (N_12738,N_11420,N_11440);
and U12739 (N_12739,N_10880,N_11736);
xnor U12740 (N_12740,N_11807,N_11757);
nand U12741 (N_12741,N_11326,N_11639);
and U12742 (N_12742,N_11235,N_11935);
nor U12743 (N_12743,N_10388,N_11492);
xor U12744 (N_12744,N_10867,N_10640);
nor U12745 (N_12745,N_10420,N_11425);
nor U12746 (N_12746,N_10937,N_11255);
nand U12747 (N_12747,N_10709,N_10534);
nand U12748 (N_12748,N_11580,N_11835);
or U12749 (N_12749,N_11601,N_11144);
or U12750 (N_12750,N_10698,N_10603);
xor U12751 (N_12751,N_10368,N_11741);
nand U12752 (N_12752,N_10293,N_11363);
xor U12753 (N_12753,N_11190,N_11834);
nand U12754 (N_12754,N_10740,N_11074);
or U12755 (N_12755,N_10963,N_10373);
xnor U12756 (N_12756,N_11894,N_11422);
nor U12757 (N_12757,N_10422,N_10188);
and U12758 (N_12758,N_11072,N_11316);
nor U12759 (N_12759,N_11693,N_11909);
nand U12760 (N_12760,N_11064,N_10421);
nand U12761 (N_12761,N_10629,N_11277);
or U12762 (N_12762,N_11257,N_10727);
nor U12763 (N_12763,N_11660,N_11571);
and U12764 (N_12764,N_10047,N_11355);
nor U12765 (N_12765,N_10533,N_11017);
or U12766 (N_12766,N_11389,N_11261);
xnor U12767 (N_12767,N_11090,N_10808);
xor U12768 (N_12768,N_11328,N_11558);
nor U12769 (N_12769,N_11298,N_11696);
and U12770 (N_12770,N_10811,N_11447);
and U12771 (N_12771,N_11619,N_10485);
and U12772 (N_12772,N_10471,N_10570);
nand U12773 (N_12773,N_10070,N_11833);
and U12774 (N_12774,N_10054,N_10924);
and U12775 (N_12775,N_11104,N_10697);
xnor U12776 (N_12776,N_10997,N_10133);
or U12777 (N_12777,N_10183,N_10413);
xor U12778 (N_12778,N_10820,N_10416);
nor U12779 (N_12779,N_11384,N_10103);
nand U12780 (N_12780,N_11407,N_10790);
or U12781 (N_12781,N_11768,N_10703);
xnor U12782 (N_12782,N_11650,N_11908);
nor U12783 (N_12783,N_10651,N_10186);
and U12784 (N_12784,N_11382,N_10778);
nand U12785 (N_12785,N_11861,N_11225);
and U12786 (N_12786,N_10718,N_10692);
and U12787 (N_12787,N_10019,N_11996);
and U12788 (N_12788,N_11724,N_11449);
or U12789 (N_12789,N_10113,N_11399);
xnor U12790 (N_12790,N_11178,N_11370);
xnor U12791 (N_12791,N_11616,N_11788);
and U12792 (N_12792,N_11231,N_10426);
and U12793 (N_12793,N_11686,N_11926);
xnor U12794 (N_12794,N_10590,N_11198);
and U12795 (N_12795,N_11037,N_10724);
xnor U12796 (N_12796,N_10265,N_11844);
and U12797 (N_12797,N_10512,N_11482);
xor U12798 (N_12798,N_11378,N_10292);
nor U12799 (N_12799,N_10511,N_11893);
nor U12800 (N_12800,N_10766,N_11010);
nor U12801 (N_12801,N_10291,N_10482);
nor U12802 (N_12802,N_10975,N_11718);
xnor U12803 (N_12803,N_10882,N_10861);
and U12804 (N_12804,N_11493,N_10264);
or U12805 (N_12805,N_10364,N_10145);
xor U12806 (N_12806,N_11860,N_10944);
and U12807 (N_12807,N_11033,N_11812);
nor U12808 (N_12808,N_11678,N_10613);
or U12809 (N_12809,N_11905,N_10466);
xnor U12810 (N_12810,N_11655,N_10460);
and U12811 (N_12811,N_10383,N_10209);
xnor U12812 (N_12812,N_11210,N_10078);
xnor U12813 (N_12813,N_10500,N_10014);
or U12814 (N_12814,N_10462,N_10491);
and U12815 (N_12815,N_11689,N_11618);
or U12816 (N_12816,N_11454,N_10964);
nand U12817 (N_12817,N_10961,N_11727);
and U12818 (N_12818,N_10921,N_10676);
xor U12819 (N_12819,N_11554,N_11058);
nor U12820 (N_12820,N_11108,N_11960);
nor U12821 (N_12821,N_11731,N_11911);
nand U12822 (N_12822,N_11068,N_10967);
nand U12823 (N_12823,N_10954,N_10225);
and U12824 (N_12824,N_10304,N_11383);
or U12825 (N_12825,N_11668,N_10504);
xor U12826 (N_12826,N_11056,N_11984);
nand U12827 (N_12827,N_11000,N_11906);
and U12828 (N_12828,N_10393,N_11070);
xnor U12829 (N_12829,N_10857,N_11353);
xnor U12830 (N_12830,N_10525,N_11325);
xnor U12831 (N_12831,N_11535,N_11126);
nor U12832 (N_12832,N_11664,N_11587);
xor U12833 (N_12833,N_10059,N_10315);
nand U12834 (N_12834,N_10008,N_11307);
nor U12835 (N_12835,N_11748,N_10493);
nor U12836 (N_12836,N_10833,N_11111);
xnor U12837 (N_12837,N_10715,N_11802);
and U12838 (N_12838,N_11116,N_10763);
and U12839 (N_12839,N_11281,N_10035);
xor U12840 (N_12840,N_11827,N_11450);
nor U12841 (N_12841,N_10366,N_10244);
nor U12842 (N_12842,N_10331,N_10618);
xor U12843 (N_12843,N_11341,N_11053);
and U12844 (N_12844,N_10467,N_11563);
xor U12845 (N_12845,N_10295,N_10254);
xor U12846 (N_12846,N_11347,N_10093);
nor U12847 (N_12847,N_10242,N_10060);
or U12848 (N_12848,N_10827,N_11048);
and U12849 (N_12849,N_10424,N_11103);
or U12850 (N_12850,N_10414,N_11077);
or U12851 (N_12851,N_11586,N_11193);
or U12852 (N_12852,N_10436,N_10843);
and U12853 (N_12853,N_11549,N_11952);
or U12854 (N_12854,N_11002,N_10803);
xnor U12855 (N_12855,N_11275,N_11153);
or U12856 (N_12856,N_10919,N_10306);
nor U12857 (N_12857,N_10744,N_10559);
xor U12858 (N_12858,N_10169,N_11233);
nor U12859 (N_12859,N_10221,N_11968);
nor U12860 (N_12860,N_11333,N_10980);
nand U12861 (N_12861,N_11745,N_11527);
and U12862 (N_12862,N_11123,N_10904);
and U12863 (N_12863,N_11798,N_11263);
nand U12864 (N_12864,N_11118,N_10211);
and U12865 (N_12865,N_10499,N_11643);
or U12866 (N_12866,N_11218,N_10299);
and U12867 (N_12867,N_11208,N_11125);
nand U12868 (N_12868,N_10237,N_10654);
or U12869 (N_12869,N_11133,N_10883);
xor U12870 (N_12870,N_10430,N_11260);
nand U12871 (N_12871,N_11243,N_11688);
and U12872 (N_12872,N_11228,N_11348);
nor U12873 (N_12873,N_11052,N_11241);
and U12874 (N_12874,N_10248,N_11669);
nor U12875 (N_12875,N_11933,N_10938);
nor U12876 (N_12876,N_10849,N_10045);
and U12877 (N_12877,N_11820,N_10607);
xor U12878 (N_12878,N_11946,N_10927);
nor U12879 (N_12879,N_11897,N_10378);
or U12880 (N_12880,N_11850,N_11071);
nor U12881 (N_12881,N_10956,N_11857);
nor U12882 (N_12882,N_10564,N_11145);
nor U12883 (N_12883,N_11620,N_11566);
nand U12884 (N_12884,N_11882,N_11051);
xnor U12885 (N_12885,N_10918,N_11124);
nand U12886 (N_12886,N_11305,N_11279);
and U12887 (N_12887,N_10455,N_10717);
nor U12888 (N_12888,N_11790,N_10850);
xnor U12889 (N_12889,N_11488,N_10445);
xor U12890 (N_12890,N_10357,N_11199);
or U12891 (N_12891,N_10988,N_11142);
or U12892 (N_12892,N_11575,N_10563);
and U12893 (N_12893,N_10162,N_10184);
nand U12894 (N_12894,N_11704,N_10300);
xnor U12895 (N_12895,N_10973,N_11117);
and U12896 (N_12896,N_11613,N_10136);
nor U12897 (N_12897,N_11369,N_11393);
or U12898 (N_12898,N_11250,N_10558);
xnor U12899 (N_12899,N_11955,N_10410);
xnor U12900 (N_12900,N_10853,N_11931);
or U12901 (N_12901,N_10807,N_10616);
nand U12902 (N_12902,N_10354,N_10105);
or U12903 (N_12903,N_11259,N_11883);
or U12904 (N_12904,N_11237,N_11842);
xor U12905 (N_12905,N_10147,N_10003);
nor U12906 (N_12906,N_10177,N_10148);
nand U12907 (N_12907,N_11106,N_10736);
nand U12908 (N_12908,N_11973,N_11733);
nand U12909 (N_12909,N_10829,N_11653);
nor U12910 (N_12910,N_11031,N_11725);
and U12911 (N_12911,N_10902,N_10678);
nand U12912 (N_12912,N_10910,N_10498);
or U12913 (N_12913,N_11018,N_11560);
nor U12914 (N_12914,N_11772,N_10079);
nand U12915 (N_12915,N_10138,N_11131);
or U12916 (N_12916,N_11879,N_11548);
nor U12917 (N_12917,N_11115,N_11418);
and U12918 (N_12918,N_10488,N_10230);
xnor U12919 (N_12919,N_10170,N_10015);
and U12920 (N_12920,N_10092,N_11433);
or U12921 (N_12921,N_10344,N_10881);
or U12922 (N_12922,N_11830,N_11774);
and U12923 (N_12923,N_10256,N_11794);
xnor U12924 (N_12924,N_10781,N_10948);
or U12925 (N_12925,N_11236,N_10120);
and U12926 (N_12926,N_11819,N_10208);
nor U12927 (N_12927,N_11203,N_11780);
nor U12928 (N_12928,N_11939,N_11917);
nor U12929 (N_12929,N_10650,N_11957);
nor U12930 (N_12930,N_10529,N_11426);
nand U12931 (N_12931,N_10683,N_10446);
or U12932 (N_12932,N_11760,N_11069);
or U12933 (N_12933,N_11318,N_11561);
nand U12934 (N_12934,N_11938,N_10094);
nand U12935 (N_12935,N_11967,N_10464);
nor U12936 (N_12936,N_10968,N_11343);
or U12937 (N_12937,N_11552,N_10384);
or U12938 (N_12938,N_11502,N_10877);
nand U12939 (N_12939,N_11127,N_11932);
nand U12940 (N_12940,N_10399,N_11019);
or U12941 (N_12941,N_11899,N_10793);
and U12942 (N_12942,N_11625,N_11916);
nand U12943 (N_12943,N_10733,N_10407);
and U12944 (N_12944,N_10433,N_11317);
nand U12945 (N_12945,N_11959,N_11387);
and U12946 (N_12946,N_10101,N_10719);
nand U12947 (N_12947,N_10219,N_10346);
xnor U12948 (N_12948,N_11634,N_11695);
nand U12949 (N_12949,N_10873,N_11262);
nand U12950 (N_12950,N_11470,N_11062);
or U12951 (N_12951,N_11520,N_11164);
nand U12952 (N_12952,N_10972,N_10899);
nor U12953 (N_12953,N_10217,N_11591);
nor U12954 (N_12954,N_10780,N_10309);
nor U12955 (N_12955,N_11455,N_11168);
nor U12956 (N_12956,N_11293,N_11491);
xor U12957 (N_12957,N_10397,N_10203);
nand U12958 (N_12958,N_10657,N_11459);
nand U12959 (N_12959,N_11003,N_10852);
or U12960 (N_12960,N_11022,N_11294);
or U12961 (N_12961,N_10279,N_10897);
or U12962 (N_12962,N_10515,N_10561);
nand U12963 (N_12963,N_10370,N_10637);
xor U12964 (N_12964,N_10017,N_10588);
nand U12965 (N_12965,N_10351,N_11569);
nand U12966 (N_12966,N_10141,N_10067);
xnor U12967 (N_12967,N_11148,N_11707);
or U12968 (N_12968,N_10175,N_11337);
or U12969 (N_12969,N_10767,N_10196);
xnor U12970 (N_12970,N_10473,N_10077);
and U12971 (N_12971,N_10953,N_11371);
and U12972 (N_12972,N_11594,N_11896);
xnor U12973 (N_12973,N_11331,N_10437);
nand U12974 (N_12974,N_11385,N_11568);
nand U12975 (N_12975,N_11740,N_11122);
xor U12976 (N_12976,N_11511,N_10814);
xnor U12977 (N_12977,N_11930,N_11578);
nand U12978 (N_12978,N_11584,N_11995);
xnor U12979 (N_12979,N_10112,N_11094);
nand U12980 (N_12980,N_11160,N_10013);
nand U12981 (N_12981,N_11612,N_10082);
or U12982 (N_12982,N_10788,N_10634);
nor U12983 (N_12983,N_11039,N_11515);
or U12984 (N_12984,N_10009,N_11626);
xor U12985 (N_12985,N_10405,N_11965);
nor U12986 (N_12986,N_10305,N_11308);
nor U12987 (N_12987,N_11254,N_11805);
and U12988 (N_12988,N_10636,N_11112);
or U12989 (N_12989,N_11614,N_11524);
xnor U12990 (N_12990,N_11576,N_10027);
and U12991 (N_12991,N_11753,N_11463);
xnor U12992 (N_12992,N_11129,N_11913);
xnor U12993 (N_12993,N_10773,N_10213);
and U12994 (N_12994,N_10884,N_10087);
nor U12995 (N_12995,N_11534,N_11012);
nor U12996 (N_12996,N_10554,N_10381);
xnor U12997 (N_12997,N_10648,N_10772);
nand U12998 (N_12998,N_10642,N_10179);
xnor U12999 (N_12999,N_10214,N_10091);
or U13000 (N_13000,N_11359,N_10012);
nor U13001 (N_13001,N_11049,N_11420);
nand U13002 (N_13002,N_11238,N_11216);
and U13003 (N_13003,N_11693,N_10738);
nor U13004 (N_13004,N_11440,N_10265);
xor U13005 (N_13005,N_10583,N_11090);
nand U13006 (N_13006,N_10879,N_11017);
nor U13007 (N_13007,N_10265,N_10378);
or U13008 (N_13008,N_11823,N_11467);
xnor U13009 (N_13009,N_11416,N_10023);
or U13010 (N_13010,N_10345,N_11795);
nand U13011 (N_13011,N_11541,N_11236);
nand U13012 (N_13012,N_11433,N_11763);
nor U13013 (N_13013,N_10557,N_10216);
or U13014 (N_13014,N_10060,N_11422);
nand U13015 (N_13015,N_10988,N_10201);
or U13016 (N_13016,N_11733,N_10632);
or U13017 (N_13017,N_11219,N_10036);
nor U13018 (N_13018,N_11141,N_11567);
xnor U13019 (N_13019,N_10115,N_11021);
nor U13020 (N_13020,N_10172,N_11204);
and U13021 (N_13021,N_11381,N_11661);
and U13022 (N_13022,N_11231,N_10922);
or U13023 (N_13023,N_11255,N_10269);
xnor U13024 (N_13024,N_10912,N_10982);
nor U13025 (N_13025,N_11455,N_11434);
xnor U13026 (N_13026,N_10564,N_10654);
or U13027 (N_13027,N_10145,N_11443);
nand U13028 (N_13028,N_11797,N_10590);
xnor U13029 (N_13029,N_11931,N_10493);
and U13030 (N_13030,N_11617,N_11325);
and U13031 (N_13031,N_11543,N_11701);
nand U13032 (N_13032,N_10637,N_11636);
or U13033 (N_13033,N_10900,N_11327);
and U13034 (N_13034,N_10537,N_11819);
nand U13035 (N_13035,N_10424,N_11475);
or U13036 (N_13036,N_10681,N_10033);
and U13037 (N_13037,N_11868,N_11266);
xnor U13038 (N_13038,N_10739,N_11897);
nor U13039 (N_13039,N_10528,N_10467);
and U13040 (N_13040,N_10979,N_10234);
or U13041 (N_13041,N_10395,N_11830);
nor U13042 (N_13042,N_11980,N_11585);
and U13043 (N_13043,N_10226,N_11480);
nor U13044 (N_13044,N_10346,N_10565);
xnor U13045 (N_13045,N_11984,N_10541);
xor U13046 (N_13046,N_11914,N_10008);
or U13047 (N_13047,N_10999,N_10540);
xor U13048 (N_13048,N_10447,N_11387);
nor U13049 (N_13049,N_11490,N_10598);
nor U13050 (N_13050,N_10043,N_10737);
or U13051 (N_13051,N_10251,N_11665);
and U13052 (N_13052,N_11285,N_10211);
and U13053 (N_13053,N_11317,N_11816);
nand U13054 (N_13054,N_11194,N_10231);
xnor U13055 (N_13055,N_10671,N_11610);
and U13056 (N_13056,N_11982,N_10928);
nand U13057 (N_13057,N_10904,N_11048);
and U13058 (N_13058,N_10062,N_11077);
or U13059 (N_13059,N_11808,N_10361);
or U13060 (N_13060,N_11612,N_10974);
or U13061 (N_13061,N_11686,N_11352);
or U13062 (N_13062,N_11160,N_10448);
or U13063 (N_13063,N_11929,N_10172);
and U13064 (N_13064,N_11565,N_11454);
or U13065 (N_13065,N_10640,N_10716);
nand U13066 (N_13066,N_10496,N_10741);
or U13067 (N_13067,N_10166,N_11539);
xor U13068 (N_13068,N_10126,N_10106);
and U13069 (N_13069,N_10677,N_10322);
and U13070 (N_13070,N_10830,N_11998);
nor U13071 (N_13071,N_11184,N_11193);
and U13072 (N_13072,N_10975,N_11406);
nand U13073 (N_13073,N_11103,N_10188);
nor U13074 (N_13074,N_10240,N_11523);
xor U13075 (N_13075,N_10139,N_11053);
xnor U13076 (N_13076,N_11960,N_10424);
and U13077 (N_13077,N_10139,N_11043);
nor U13078 (N_13078,N_10727,N_10952);
and U13079 (N_13079,N_11545,N_11162);
xor U13080 (N_13080,N_10330,N_10001);
or U13081 (N_13081,N_10238,N_11297);
nor U13082 (N_13082,N_11149,N_10894);
xor U13083 (N_13083,N_10794,N_10549);
and U13084 (N_13084,N_11066,N_11854);
nor U13085 (N_13085,N_10007,N_10582);
and U13086 (N_13086,N_11223,N_10058);
and U13087 (N_13087,N_11910,N_10176);
xor U13088 (N_13088,N_11415,N_11980);
xnor U13089 (N_13089,N_10790,N_10114);
xnor U13090 (N_13090,N_11847,N_10061);
and U13091 (N_13091,N_11538,N_10839);
and U13092 (N_13092,N_10981,N_10945);
or U13093 (N_13093,N_10786,N_11714);
nand U13094 (N_13094,N_11984,N_10853);
xor U13095 (N_13095,N_11325,N_10028);
nor U13096 (N_13096,N_11631,N_11525);
and U13097 (N_13097,N_10202,N_10319);
nand U13098 (N_13098,N_10340,N_10654);
xnor U13099 (N_13099,N_10605,N_10615);
and U13100 (N_13100,N_10723,N_10888);
nor U13101 (N_13101,N_11800,N_10477);
xor U13102 (N_13102,N_10156,N_11468);
xor U13103 (N_13103,N_11895,N_11696);
xor U13104 (N_13104,N_10384,N_10345);
and U13105 (N_13105,N_10967,N_11005);
xnor U13106 (N_13106,N_10634,N_11885);
or U13107 (N_13107,N_10204,N_10624);
xnor U13108 (N_13108,N_10366,N_10783);
nor U13109 (N_13109,N_10450,N_10897);
and U13110 (N_13110,N_10672,N_11039);
and U13111 (N_13111,N_10461,N_10178);
nand U13112 (N_13112,N_10384,N_10640);
nor U13113 (N_13113,N_11274,N_10100);
xor U13114 (N_13114,N_11502,N_11995);
nor U13115 (N_13115,N_10310,N_11347);
xor U13116 (N_13116,N_10453,N_11529);
nor U13117 (N_13117,N_10690,N_10502);
nor U13118 (N_13118,N_10072,N_11876);
xnor U13119 (N_13119,N_10997,N_11492);
xnor U13120 (N_13120,N_10181,N_11676);
xnor U13121 (N_13121,N_11065,N_10171);
and U13122 (N_13122,N_10807,N_10025);
and U13123 (N_13123,N_10996,N_11964);
and U13124 (N_13124,N_11865,N_11092);
xnor U13125 (N_13125,N_11014,N_10146);
or U13126 (N_13126,N_10709,N_11383);
nor U13127 (N_13127,N_11144,N_11986);
or U13128 (N_13128,N_10469,N_11334);
or U13129 (N_13129,N_10608,N_10562);
nand U13130 (N_13130,N_10003,N_11770);
and U13131 (N_13131,N_11687,N_10859);
or U13132 (N_13132,N_10366,N_10021);
xor U13133 (N_13133,N_10731,N_11697);
or U13134 (N_13134,N_10150,N_11662);
or U13135 (N_13135,N_10601,N_11623);
nor U13136 (N_13136,N_10485,N_11705);
and U13137 (N_13137,N_10404,N_11297);
nor U13138 (N_13138,N_10419,N_11768);
nor U13139 (N_13139,N_10138,N_10565);
nor U13140 (N_13140,N_10671,N_10573);
and U13141 (N_13141,N_10259,N_10470);
or U13142 (N_13142,N_11391,N_10921);
nand U13143 (N_13143,N_11597,N_10615);
nor U13144 (N_13144,N_11572,N_10792);
nand U13145 (N_13145,N_11572,N_11907);
or U13146 (N_13146,N_11322,N_10135);
and U13147 (N_13147,N_10765,N_11189);
nand U13148 (N_13148,N_11593,N_11688);
and U13149 (N_13149,N_11052,N_11224);
or U13150 (N_13150,N_11987,N_11409);
or U13151 (N_13151,N_11685,N_10264);
xor U13152 (N_13152,N_10959,N_11840);
and U13153 (N_13153,N_11726,N_11913);
xnor U13154 (N_13154,N_10136,N_10252);
nor U13155 (N_13155,N_11500,N_10509);
or U13156 (N_13156,N_11502,N_11572);
and U13157 (N_13157,N_11739,N_11353);
and U13158 (N_13158,N_10708,N_10292);
nand U13159 (N_13159,N_10947,N_10618);
nand U13160 (N_13160,N_10555,N_10305);
nand U13161 (N_13161,N_10048,N_11413);
and U13162 (N_13162,N_10536,N_10616);
nand U13163 (N_13163,N_10353,N_10414);
nand U13164 (N_13164,N_11636,N_10502);
xnor U13165 (N_13165,N_10692,N_11652);
or U13166 (N_13166,N_10552,N_10001);
nor U13167 (N_13167,N_11445,N_10860);
and U13168 (N_13168,N_10931,N_11873);
and U13169 (N_13169,N_11950,N_11992);
nor U13170 (N_13170,N_10142,N_10163);
xnor U13171 (N_13171,N_10187,N_11762);
nand U13172 (N_13172,N_11243,N_10083);
nor U13173 (N_13173,N_11764,N_11700);
and U13174 (N_13174,N_11160,N_11512);
or U13175 (N_13175,N_11471,N_10177);
nand U13176 (N_13176,N_10188,N_11502);
nor U13177 (N_13177,N_10847,N_10254);
nor U13178 (N_13178,N_10944,N_10008);
xor U13179 (N_13179,N_10498,N_10549);
xor U13180 (N_13180,N_10739,N_11795);
nand U13181 (N_13181,N_10660,N_10023);
xor U13182 (N_13182,N_10172,N_11838);
xor U13183 (N_13183,N_10818,N_11176);
nor U13184 (N_13184,N_10095,N_10414);
or U13185 (N_13185,N_10652,N_10424);
and U13186 (N_13186,N_11251,N_10042);
or U13187 (N_13187,N_11510,N_11880);
nand U13188 (N_13188,N_10518,N_11311);
and U13189 (N_13189,N_11822,N_11845);
nor U13190 (N_13190,N_10918,N_11122);
nor U13191 (N_13191,N_11789,N_11638);
or U13192 (N_13192,N_11705,N_11579);
or U13193 (N_13193,N_10483,N_10600);
and U13194 (N_13194,N_11272,N_10848);
or U13195 (N_13195,N_10830,N_11373);
nand U13196 (N_13196,N_10260,N_11793);
or U13197 (N_13197,N_11570,N_10074);
xor U13198 (N_13198,N_11557,N_10221);
and U13199 (N_13199,N_11256,N_10310);
and U13200 (N_13200,N_11237,N_10891);
and U13201 (N_13201,N_11236,N_10541);
xnor U13202 (N_13202,N_11982,N_10384);
nand U13203 (N_13203,N_11558,N_10097);
xor U13204 (N_13204,N_11955,N_10453);
nand U13205 (N_13205,N_11874,N_10839);
xnor U13206 (N_13206,N_10537,N_11281);
xor U13207 (N_13207,N_11116,N_11461);
nor U13208 (N_13208,N_11191,N_11402);
nor U13209 (N_13209,N_10668,N_10612);
nand U13210 (N_13210,N_11409,N_10542);
nor U13211 (N_13211,N_11197,N_11122);
nor U13212 (N_13212,N_11835,N_10252);
nor U13213 (N_13213,N_11203,N_11028);
nand U13214 (N_13214,N_10637,N_10406);
nand U13215 (N_13215,N_11064,N_10245);
and U13216 (N_13216,N_10469,N_10367);
nand U13217 (N_13217,N_11083,N_11504);
and U13218 (N_13218,N_10421,N_11167);
or U13219 (N_13219,N_11146,N_10945);
xor U13220 (N_13220,N_11847,N_10826);
or U13221 (N_13221,N_11100,N_10190);
or U13222 (N_13222,N_10624,N_10326);
nand U13223 (N_13223,N_11491,N_10369);
and U13224 (N_13224,N_10974,N_11649);
nor U13225 (N_13225,N_10064,N_11024);
and U13226 (N_13226,N_10429,N_10325);
or U13227 (N_13227,N_11280,N_11269);
or U13228 (N_13228,N_10488,N_11909);
or U13229 (N_13229,N_10523,N_10069);
and U13230 (N_13230,N_11100,N_11379);
and U13231 (N_13231,N_11114,N_10626);
and U13232 (N_13232,N_10418,N_11164);
and U13233 (N_13233,N_10116,N_10555);
nor U13234 (N_13234,N_11305,N_11899);
nor U13235 (N_13235,N_11802,N_11257);
nor U13236 (N_13236,N_11557,N_11062);
nand U13237 (N_13237,N_10810,N_10656);
or U13238 (N_13238,N_11507,N_10423);
and U13239 (N_13239,N_11724,N_10795);
nor U13240 (N_13240,N_11446,N_10229);
and U13241 (N_13241,N_11446,N_10128);
nor U13242 (N_13242,N_10033,N_10043);
or U13243 (N_13243,N_10847,N_10549);
and U13244 (N_13244,N_11248,N_11633);
nand U13245 (N_13245,N_10260,N_10350);
and U13246 (N_13246,N_10461,N_10159);
or U13247 (N_13247,N_10855,N_11799);
xor U13248 (N_13248,N_10323,N_10225);
nor U13249 (N_13249,N_11938,N_11550);
or U13250 (N_13250,N_10926,N_11664);
or U13251 (N_13251,N_10805,N_10027);
xnor U13252 (N_13252,N_10329,N_11497);
xnor U13253 (N_13253,N_11576,N_10683);
and U13254 (N_13254,N_10752,N_11288);
nor U13255 (N_13255,N_11111,N_11877);
or U13256 (N_13256,N_11923,N_10436);
nand U13257 (N_13257,N_10240,N_10160);
nor U13258 (N_13258,N_10561,N_11576);
xnor U13259 (N_13259,N_11654,N_10703);
nand U13260 (N_13260,N_10163,N_11274);
and U13261 (N_13261,N_10629,N_11208);
xnor U13262 (N_13262,N_11762,N_11034);
xnor U13263 (N_13263,N_10094,N_11736);
and U13264 (N_13264,N_11573,N_10195);
nand U13265 (N_13265,N_10651,N_10922);
or U13266 (N_13266,N_11327,N_10309);
or U13267 (N_13267,N_10744,N_10045);
or U13268 (N_13268,N_10436,N_11160);
nor U13269 (N_13269,N_11319,N_11190);
nor U13270 (N_13270,N_11244,N_10431);
and U13271 (N_13271,N_11373,N_11473);
xnor U13272 (N_13272,N_10699,N_11111);
nor U13273 (N_13273,N_11565,N_11212);
or U13274 (N_13274,N_11542,N_11152);
or U13275 (N_13275,N_10225,N_11173);
nand U13276 (N_13276,N_11286,N_11259);
nand U13277 (N_13277,N_10680,N_11042);
or U13278 (N_13278,N_11357,N_11294);
nor U13279 (N_13279,N_11588,N_10410);
nand U13280 (N_13280,N_10169,N_10245);
nand U13281 (N_13281,N_11338,N_11905);
xnor U13282 (N_13282,N_11088,N_11569);
or U13283 (N_13283,N_10251,N_11997);
and U13284 (N_13284,N_10393,N_10856);
xor U13285 (N_13285,N_11228,N_11356);
xnor U13286 (N_13286,N_10042,N_11114);
or U13287 (N_13287,N_10120,N_11314);
or U13288 (N_13288,N_10795,N_10192);
nor U13289 (N_13289,N_11469,N_11905);
nor U13290 (N_13290,N_10229,N_10069);
or U13291 (N_13291,N_11839,N_10561);
xnor U13292 (N_13292,N_11647,N_10249);
nand U13293 (N_13293,N_11315,N_11515);
or U13294 (N_13294,N_10973,N_11455);
or U13295 (N_13295,N_11499,N_10802);
and U13296 (N_13296,N_10787,N_11979);
nand U13297 (N_13297,N_10219,N_10762);
nor U13298 (N_13298,N_10771,N_10455);
nor U13299 (N_13299,N_10802,N_11804);
or U13300 (N_13300,N_11736,N_11624);
nor U13301 (N_13301,N_10465,N_11895);
xor U13302 (N_13302,N_11536,N_10467);
nand U13303 (N_13303,N_11939,N_11300);
nor U13304 (N_13304,N_11324,N_10193);
and U13305 (N_13305,N_11442,N_11542);
nand U13306 (N_13306,N_10702,N_11553);
nand U13307 (N_13307,N_11476,N_11413);
nor U13308 (N_13308,N_10890,N_11483);
or U13309 (N_13309,N_10512,N_11952);
xor U13310 (N_13310,N_10579,N_11187);
nor U13311 (N_13311,N_11064,N_11060);
nand U13312 (N_13312,N_11706,N_11081);
and U13313 (N_13313,N_10045,N_11499);
nor U13314 (N_13314,N_10891,N_11211);
nand U13315 (N_13315,N_10063,N_10571);
nor U13316 (N_13316,N_11535,N_11046);
xnor U13317 (N_13317,N_11423,N_10529);
nand U13318 (N_13318,N_10519,N_10028);
xnor U13319 (N_13319,N_10709,N_10125);
or U13320 (N_13320,N_11907,N_10300);
nand U13321 (N_13321,N_10453,N_10235);
nand U13322 (N_13322,N_10569,N_11339);
nor U13323 (N_13323,N_10487,N_10060);
xnor U13324 (N_13324,N_10302,N_10597);
xor U13325 (N_13325,N_11450,N_11697);
nand U13326 (N_13326,N_10358,N_10406);
nand U13327 (N_13327,N_10735,N_10325);
nand U13328 (N_13328,N_10737,N_11622);
xor U13329 (N_13329,N_11680,N_11496);
and U13330 (N_13330,N_11447,N_11935);
nand U13331 (N_13331,N_11310,N_11486);
and U13332 (N_13332,N_11427,N_11433);
xnor U13333 (N_13333,N_10332,N_11292);
nor U13334 (N_13334,N_11304,N_11052);
and U13335 (N_13335,N_10389,N_11056);
nor U13336 (N_13336,N_10606,N_10982);
and U13337 (N_13337,N_11137,N_11535);
nor U13338 (N_13338,N_10907,N_10837);
xor U13339 (N_13339,N_10340,N_11544);
nor U13340 (N_13340,N_11105,N_10067);
nor U13341 (N_13341,N_10342,N_11798);
or U13342 (N_13342,N_10280,N_11578);
nor U13343 (N_13343,N_10134,N_10485);
or U13344 (N_13344,N_10428,N_11940);
nand U13345 (N_13345,N_11813,N_11853);
nor U13346 (N_13346,N_10946,N_10537);
or U13347 (N_13347,N_10863,N_10150);
xnor U13348 (N_13348,N_11749,N_11514);
nand U13349 (N_13349,N_10037,N_11435);
nand U13350 (N_13350,N_10850,N_10679);
nor U13351 (N_13351,N_11460,N_10681);
or U13352 (N_13352,N_11326,N_11542);
and U13353 (N_13353,N_10351,N_11577);
nor U13354 (N_13354,N_10696,N_10535);
nor U13355 (N_13355,N_11797,N_10636);
xnor U13356 (N_13356,N_11496,N_10291);
and U13357 (N_13357,N_11680,N_10850);
xor U13358 (N_13358,N_11400,N_10281);
and U13359 (N_13359,N_11835,N_10938);
or U13360 (N_13360,N_11660,N_10762);
and U13361 (N_13361,N_11385,N_10513);
nor U13362 (N_13362,N_11280,N_10091);
nand U13363 (N_13363,N_10387,N_11411);
and U13364 (N_13364,N_11872,N_11237);
xnor U13365 (N_13365,N_11864,N_11950);
and U13366 (N_13366,N_11477,N_11678);
and U13367 (N_13367,N_11018,N_10719);
and U13368 (N_13368,N_10133,N_11438);
nor U13369 (N_13369,N_11517,N_11015);
and U13370 (N_13370,N_10530,N_10005);
or U13371 (N_13371,N_11175,N_10493);
nor U13372 (N_13372,N_11200,N_11999);
or U13373 (N_13373,N_10267,N_11841);
or U13374 (N_13374,N_11768,N_11303);
and U13375 (N_13375,N_10223,N_11468);
xor U13376 (N_13376,N_11964,N_11259);
and U13377 (N_13377,N_11220,N_11124);
nor U13378 (N_13378,N_11213,N_10350);
nor U13379 (N_13379,N_11909,N_11498);
nor U13380 (N_13380,N_11594,N_10840);
xor U13381 (N_13381,N_11920,N_10211);
nand U13382 (N_13382,N_11646,N_10628);
or U13383 (N_13383,N_10837,N_11992);
nand U13384 (N_13384,N_11094,N_11639);
nor U13385 (N_13385,N_10951,N_11786);
xnor U13386 (N_13386,N_10291,N_10656);
nor U13387 (N_13387,N_11524,N_10465);
xnor U13388 (N_13388,N_10130,N_10096);
nor U13389 (N_13389,N_11605,N_11575);
and U13390 (N_13390,N_10385,N_10906);
and U13391 (N_13391,N_10158,N_10347);
nor U13392 (N_13392,N_11043,N_10932);
and U13393 (N_13393,N_11223,N_10805);
nor U13394 (N_13394,N_10988,N_10790);
xor U13395 (N_13395,N_11479,N_10635);
nor U13396 (N_13396,N_11982,N_10616);
nor U13397 (N_13397,N_11162,N_11988);
nor U13398 (N_13398,N_11851,N_11708);
nor U13399 (N_13399,N_11013,N_10114);
nand U13400 (N_13400,N_11882,N_11323);
xnor U13401 (N_13401,N_11794,N_11469);
nand U13402 (N_13402,N_10075,N_10683);
and U13403 (N_13403,N_11304,N_11663);
and U13404 (N_13404,N_11976,N_11793);
or U13405 (N_13405,N_11390,N_10779);
or U13406 (N_13406,N_11063,N_11040);
or U13407 (N_13407,N_10463,N_10621);
nor U13408 (N_13408,N_10070,N_11501);
and U13409 (N_13409,N_11187,N_10628);
nor U13410 (N_13410,N_10511,N_10860);
xnor U13411 (N_13411,N_11792,N_10968);
xor U13412 (N_13412,N_11909,N_11383);
xnor U13413 (N_13413,N_11639,N_10807);
and U13414 (N_13414,N_11376,N_11218);
nand U13415 (N_13415,N_10101,N_11299);
nand U13416 (N_13416,N_11973,N_10202);
xnor U13417 (N_13417,N_11857,N_11677);
nor U13418 (N_13418,N_10397,N_10635);
nor U13419 (N_13419,N_10904,N_10718);
or U13420 (N_13420,N_11007,N_11322);
or U13421 (N_13421,N_10775,N_10453);
or U13422 (N_13422,N_10031,N_10085);
xor U13423 (N_13423,N_10562,N_11907);
and U13424 (N_13424,N_11613,N_11602);
nand U13425 (N_13425,N_11813,N_10438);
nand U13426 (N_13426,N_11635,N_10317);
or U13427 (N_13427,N_10665,N_10825);
xor U13428 (N_13428,N_11621,N_11917);
or U13429 (N_13429,N_10618,N_11662);
or U13430 (N_13430,N_10760,N_11731);
and U13431 (N_13431,N_11777,N_11766);
nor U13432 (N_13432,N_11265,N_11933);
xnor U13433 (N_13433,N_10965,N_10302);
and U13434 (N_13434,N_11675,N_10562);
nand U13435 (N_13435,N_10398,N_11030);
nand U13436 (N_13436,N_10766,N_10136);
and U13437 (N_13437,N_11405,N_11919);
and U13438 (N_13438,N_10271,N_10177);
or U13439 (N_13439,N_11838,N_11880);
or U13440 (N_13440,N_11197,N_10469);
nand U13441 (N_13441,N_10380,N_11559);
and U13442 (N_13442,N_11039,N_11934);
nor U13443 (N_13443,N_11030,N_11067);
and U13444 (N_13444,N_10052,N_11054);
nand U13445 (N_13445,N_10689,N_10299);
xnor U13446 (N_13446,N_11552,N_10045);
or U13447 (N_13447,N_11968,N_11146);
or U13448 (N_13448,N_11048,N_11977);
or U13449 (N_13449,N_11173,N_11409);
nor U13450 (N_13450,N_10383,N_11338);
nand U13451 (N_13451,N_10952,N_10313);
xnor U13452 (N_13452,N_11897,N_10054);
nand U13453 (N_13453,N_11185,N_10794);
and U13454 (N_13454,N_10187,N_10630);
or U13455 (N_13455,N_11745,N_10696);
and U13456 (N_13456,N_10068,N_11706);
or U13457 (N_13457,N_10947,N_10228);
nor U13458 (N_13458,N_11449,N_11161);
or U13459 (N_13459,N_10511,N_11491);
xor U13460 (N_13460,N_11422,N_10274);
nand U13461 (N_13461,N_11414,N_11010);
nor U13462 (N_13462,N_10628,N_11308);
nand U13463 (N_13463,N_11258,N_11587);
or U13464 (N_13464,N_11837,N_10852);
or U13465 (N_13465,N_10838,N_10251);
and U13466 (N_13466,N_11904,N_10368);
nor U13467 (N_13467,N_11871,N_11093);
xor U13468 (N_13468,N_10584,N_11437);
nand U13469 (N_13469,N_11161,N_10392);
nor U13470 (N_13470,N_11215,N_11018);
and U13471 (N_13471,N_10935,N_10543);
nor U13472 (N_13472,N_10161,N_10090);
nor U13473 (N_13473,N_10721,N_10632);
nand U13474 (N_13474,N_11183,N_11684);
nand U13475 (N_13475,N_11848,N_11733);
nor U13476 (N_13476,N_10761,N_10838);
xor U13477 (N_13477,N_11682,N_11732);
nor U13478 (N_13478,N_10130,N_11444);
and U13479 (N_13479,N_11047,N_11287);
nand U13480 (N_13480,N_10645,N_10309);
xnor U13481 (N_13481,N_10748,N_10788);
xor U13482 (N_13482,N_10597,N_11759);
xor U13483 (N_13483,N_10804,N_11083);
and U13484 (N_13484,N_11346,N_10015);
and U13485 (N_13485,N_10036,N_10597);
and U13486 (N_13486,N_10765,N_10826);
nor U13487 (N_13487,N_11247,N_11192);
xnor U13488 (N_13488,N_10179,N_10111);
nand U13489 (N_13489,N_11281,N_10155);
nand U13490 (N_13490,N_11770,N_10648);
and U13491 (N_13491,N_10318,N_10131);
xor U13492 (N_13492,N_10842,N_11623);
nor U13493 (N_13493,N_11566,N_11963);
nor U13494 (N_13494,N_10347,N_10773);
nand U13495 (N_13495,N_10152,N_11212);
or U13496 (N_13496,N_10540,N_11935);
and U13497 (N_13497,N_10791,N_10782);
and U13498 (N_13498,N_11912,N_11071);
nor U13499 (N_13499,N_11982,N_10534);
and U13500 (N_13500,N_11043,N_11670);
nand U13501 (N_13501,N_11872,N_10319);
xor U13502 (N_13502,N_11336,N_11158);
nand U13503 (N_13503,N_11637,N_11608);
and U13504 (N_13504,N_11431,N_10655);
or U13505 (N_13505,N_10060,N_10386);
and U13506 (N_13506,N_10318,N_11897);
nor U13507 (N_13507,N_10241,N_11266);
xor U13508 (N_13508,N_10186,N_10844);
or U13509 (N_13509,N_11143,N_11473);
or U13510 (N_13510,N_10929,N_10975);
nand U13511 (N_13511,N_10105,N_11553);
or U13512 (N_13512,N_10957,N_11769);
or U13513 (N_13513,N_11539,N_11810);
nand U13514 (N_13514,N_11407,N_11876);
nor U13515 (N_13515,N_11902,N_10755);
xor U13516 (N_13516,N_11291,N_10300);
xnor U13517 (N_13517,N_10585,N_10425);
nand U13518 (N_13518,N_10116,N_10850);
nor U13519 (N_13519,N_10377,N_11503);
nand U13520 (N_13520,N_10848,N_11831);
nand U13521 (N_13521,N_10277,N_11718);
nor U13522 (N_13522,N_11175,N_10649);
nor U13523 (N_13523,N_10508,N_11922);
nor U13524 (N_13524,N_10244,N_11081);
xor U13525 (N_13525,N_10633,N_10540);
xor U13526 (N_13526,N_11708,N_10063);
nor U13527 (N_13527,N_11020,N_11425);
xor U13528 (N_13528,N_10510,N_11701);
and U13529 (N_13529,N_11346,N_11321);
nor U13530 (N_13530,N_11664,N_11529);
nor U13531 (N_13531,N_10505,N_10236);
nor U13532 (N_13532,N_11874,N_10140);
nor U13533 (N_13533,N_11387,N_10234);
xnor U13534 (N_13534,N_11082,N_11201);
nor U13535 (N_13535,N_10268,N_11154);
xnor U13536 (N_13536,N_10460,N_11907);
xor U13537 (N_13537,N_11667,N_10026);
and U13538 (N_13538,N_11346,N_11827);
nand U13539 (N_13539,N_10918,N_11098);
or U13540 (N_13540,N_10389,N_10503);
or U13541 (N_13541,N_10934,N_11564);
or U13542 (N_13542,N_10415,N_11750);
nand U13543 (N_13543,N_11923,N_11906);
nor U13544 (N_13544,N_11426,N_10354);
nor U13545 (N_13545,N_11045,N_11292);
xor U13546 (N_13546,N_10009,N_11889);
and U13547 (N_13547,N_11218,N_10338);
nand U13548 (N_13548,N_10081,N_10384);
xor U13549 (N_13549,N_11163,N_11447);
or U13550 (N_13550,N_10278,N_11560);
nand U13551 (N_13551,N_11307,N_10095);
nor U13552 (N_13552,N_10744,N_10180);
xnor U13553 (N_13553,N_11322,N_11820);
xnor U13554 (N_13554,N_10261,N_10595);
nand U13555 (N_13555,N_10765,N_11589);
or U13556 (N_13556,N_11913,N_11886);
or U13557 (N_13557,N_10736,N_11145);
xnor U13558 (N_13558,N_10328,N_10234);
or U13559 (N_13559,N_10864,N_11878);
nand U13560 (N_13560,N_11956,N_10432);
and U13561 (N_13561,N_10266,N_10901);
xor U13562 (N_13562,N_10981,N_11762);
xor U13563 (N_13563,N_10265,N_10669);
nor U13564 (N_13564,N_11546,N_10478);
nor U13565 (N_13565,N_11085,N_11137);
and U13566 (N_13566,N_11970,N_11652);
xor U13567 (N_13567,N_10413,N_11026);
and U13568 (N_13568,N_10836,N_10846);
nand U13569 (N_13569,N_10927,N_10525);
or U13570 (N_13570,N_11431,N_11455);
and U13571 (N_13571,N_10242,N_10911);
nor U13572 (N_13572,N_10750,N_11879);
xor U13573 (N_13573,N_10267,N_11989);
or U13574 (N_13574,N_10569,N_11676);
nand U13575 (N_13575,N_11958,N_11581);
nor U13576 (N_13576,N_10251,N_11763);
nand U13577 (N_13577,N_11185,N_10371);
xor U13578 (N_13578,N_10383,N_11248);
nor U13579 (N_13579,N_11051,N_11247);
or U13580 (N_13580,N_10806,N_10559);
nand U13581 (N_13581,N_11828,N_11946);
or U13582 (N_13582,N_10780,N_10958);
or U13583 (N_13583,N_10646,N_11807);
and U13584 (N_13584,N_10577,N_11210);
nand U13585 (N_13585,N_10792,N_11619);
or U13586 (N_13586,N_11470,N_10744);
or U13587 (N_13587,N_10652,N_10657);
nand U13588 (N_13588,N_11663,N_10497);
nor U13589 (N_13589,N_11709,N_11632);
or U13590 (N_13590,N_11733,N_10414);
nand U13591 (N_13591,N_11665,N_10177);
xnor U13592 (N_13592,N_10844,N_11169);
or U13593 (N_13593,N_11029,N_10975);
xor U13594 (N_13594,N_11580,N_10910);
nor U13595 (N_13595,N_10113,N_11910);
nand U13596 (N_13596,N_10695,N_10566);
and U13597 (N_13597,N_11768,N_10122);
or U13598 (N_13598,N_10873,N_11667);
or U13599 (N_13599,N_11576,N_10818);
and U13600 (N_13600,N_10857,N_11443);
and U13601 (N_13601,N_10645,N_10873);
nand U13602 (N_13602,N_11151,N_11092);
or U13603 (N_13603,N_10225,N_11060);
nor U13604 (N_13604,N_11021,N_10668);
nand U13605 (N_13605,N_10038,N_10312);
or U13606 (N_13606,N_10419,N_10397);
and U13607 (N_13607,N_11303,N_11458);
and U13608 (N_13608,N_11028,N_10190);
nor U13609 (N_13609,N_11510,N_11709);
xor U13610 (N_13610,N_11950,N_11523);
nand U13611 (N_13611,N_11750,N_11384);
nor U13612 (N_13612,N_11635,N_10748);
nor U13613 (N_13613,N_10632,N_10306);
and U13614 (N_13614,N_11527,N_10991);
nand U13615 (N_13615,N_11941,N_11551);
and U13616 (N_13616,N_10718,N_11326);
nand U13617 (N_13617,N_11630,N_11117);
nor U13618 (N_13618,N_11931,N_10435);
nand U13619 (N_13619,N_11369,N_10723);
nor U13620 (N_13620,N_11798,N_10142);
nand U13621 (N_13621,N_11697,N_10412);
or U13622 (N_13622,N_10827,N_11060);
nor U13623 (N_13623,N_10659,N_11384);
xnor U13624 (N_13624,N_10944,N_11588);
nor U13625 (N_13625,N_11678,N_10133);
and U13626 (N_13626,N_11601,N_10652);
nor U13627 (N_13627,N_10912,N_10435);
nand U13628 (N_13628,N_11703,N_10664);
nand U13629 (N_13629,N_11233,N_10616);
and U13630 (N_13630,N_11450,N_10882);
nand U13631 (N_13631,N_11523,N_10785);
nor U13632 (N_13632,N_11563,N_10342);
or U13633 (N_13633,N_10199,N_11901);
nor U13634 (N_13634,N_10159,N_11834);
nor U13635 (N_13635,N_10827,N_11616);
or U13636 (N_13636,N_11379,N_11137);
and U13637 (N_13637,N_11771,N_11973);
and U13638 (N_13638,N_11110,N_10810);
or U13639 (N_13639,N_10351,N_11059);
xnor U13640 (N_13640,N_10978,N_10609);
xor U13641 (N_13641,N_10170,N_11463);
nor U13642 (N_13642,N_10279,N_11256);
or U13643 (N_13643,N_10003,N_10439);
or U13644 (N_13644,N_11567,N_11285);
and U13645 (N_13645,N_10037,N_10848);
xnor U13646 (N_13646,N_11795,N_10990);
or U13647 (N_13647,N_10443,N_10706);
or U13648 (N_13648,N_10182,N_10849);
xnor U13649 (N_13649,N_10907,N_10858);
or U13650 (N_13650,N_10870,N_11257);
or U13651 (N_13651,N_10961,N_11995);
and U13652 (N_13652,N_11205,N_11305);
or U13653 (N_13653,N_10732,N_10642);
and U13654 (N_13654,N_10954,N_11079);
or U13655 (N_13655,N_11750,N_11838);
nand U13656 (N_13656,N_10523,N_11437);
or U13657 (N_13657,N_11546,N_10029);
xor U13658 (N_13658,N_10857,N_11211);
and U13659 (N_13659,N_10054,N_11399);
or U13660 (N_13660,N_11624,N_11017);
or U13661 (N_13661,N_10119,N_11721);
and U13662 (N_13662,N_10561,N_10639);
or U13663 (N_13663,N_10821,N_11879);
nand U13664 (N_13664,N_10359,N_11662);
or U13665 (N_13665,N_11283,N_10366);
nor U13666 (N_13666,N_11358,N_10903);
nor U13667 (N_13667,N_11295,N_10414);
or U13668 (N_13668,N_11476,N_10292);
nand U13669 (N_13669,N_10348,N_10955);
nor U13670 (N_13670,N_11107,N_11791);
nand U13671 (N_13671,N_10899,N_11463);
nand U13672 (N_13672,N_11764,N_10287);
nor U13673 (N_13673,N_10443,N_10914);
nand U13674 (N_13674,N_11446,N_10428);
and U13675 (N_13675,N_11228,N_11760);
or U13676 (N_13676,N_11971,N_10472);
xnor U13677 (N_13677,N_10657,N_10896);
nor U13678 (N_13678,N_11535,N_10976);
or U13679 (N_13679,N_10010,N_11136);
or U13680 (N_13680,N_11386,N_11507);
nand U13681 (N_13681,N_10163,N_10890);
xor U13682 (N_13682,N_10275,N_11365);
and U13683 (N_13683,N_11791,N_10527);
nor U13684 (N_13684,N_10689,N_10930);
xor U13685 (N_13685,N_11728,N_11720);
nand U13686 (N_13686,N_11558,N_10961);
xor U13687 (N_13687,N_10095,N_11452);
nand U13688 (N_13688,N_11641,N_11566);
xnor U13689 (N_13689,N_10810,N_10247);
and U13690 (N_13690,N_11804,N_10774);
nor U13691 (N_13691,N_10322,N_10511);
and U13692 (N_13692,N_11513,N_10269);
nand U13693 (N_13693,N_10113,N_10269);
xor U13694 (N_13694,N_10447,N_11210);
and U13695 (N_13695,N_11400,N_11770);
xnor U13696 (N_13696,N_11253,N_10984);
nor U13697 (N_13697,N_10026,N_10694);
or U13698 (N_13698,N_10808,N_10963);
or U13699 (N_13699,N_11679,N_11196);
or U13700 (N_13700,N_10353,N_11520);
or U13701 (N_13701,N_10905,N_11605);
or U13702 (N_13702,N_10140,N_11323);
nand U13703 (N_13703,N_10591,N_11681);
and U13704 (N_13704,N_10998,N_10643);
or U13705 (N_13705,N_10820,N_10422);
xor U13706 (N_13706,N_11123,N_10645);
and U13707 (N_13707,N_10598,N_11101);
and U13708 (N_13708,N_11683,N_11179);
and U13709 (N_13709,N_10697,N_11540);
nor U13710 (N_13710,N_11884,N_11827);
nor U13711 (N_13711,N_10109,N_10203);
and U13712 (N_13712,N_10100,N_10787);
nor U13713 (N_13713,N_10693,N_10271);
or U13714 (N_13714,N_10472,N_11007);
xnor U13715 (N_13715,N_10966,N_10499);
nand U13716 (N_13716,N_11114,N_11983);
or U13717 (N_13717,N_10032,N_10732);
xnor U13718 (N_13718,N_11159,N_10583);
or U13719 (N_13719,N_10370,N_10070);
xor U13720 (N_13720,N_11288,N_11479);
xnor U13721 (N_13721,N_10133,N_11826);
and U13722 (N_13722,N_11611,N_10113);
xor U13723 (N_13723,N_11794,N_10607);
nor U13724 (N_13724,N_10949,N_10548);
and U13725 (N_13725,N_10768,N_11834);
nand U13726 (N_13726,N_10781,N_11003);
nand U13727 (N_13727,N_11640,N_10526);
nand U13728 (N_13728,N_11860,N_10529);
xor U13729 (N_13729,N_11991,N_10628);
or U13730 (N_13730,N_10380,N_10035);
nand U13731 (N_13731,N_11935,N_10330);
xor U13732 (N_13732,N_11096,N_11883);
or U13733 (N_13733,N_11367,N_11957);
and U13734 (N_13734,N_10248,N_11602);
and U13735 (N_13735,N_10050,N_11054);
nor U13736 (N_13736,N_10156,N_10114);
xnor U13737 (N_13737,N_11254,N_11659);
nand U13738 (N_13738,N_10224,N_10774);
xnor U13739 (N_13739,N_10919,N_10879);
nor U13740 (N_13740,N_10106,N_10828);
xor U13741 (N_13741,N_10093,N_10096);
or U13742 (N_13742,N_10330,N_10409);
or U13743 (N_13743,N_10224,N_10561);
and U13744 (N_13744,N_11868,N_11336);
nand U13745 (N_13745,N_10574,N_11309);
xor U13746 (N_13746,N_11561,N_10818);
and U13747 (N_13747,N_10666,N_10746);
nor U13748 (N_13748,N_11663,N_10444);
or U13749 (N_13749,N_10454,N_11306);
xnor U13750 (N_13750,N_10450,N_11166);
nor U13751 (N_13751,N_11017,N_11332);
nor U13752 (N_13752,N_11363,N_10378);
nand U13753 (N_13753,N_10699,N_11691);
or U13754 (N_13754,N_10237,N_11754);
or U13755 (N_13755,N_11429,N_11459);
xnor U13756 (N_13756,N_11665,N_11569);
and U13757 (N_13757,N_11550,N_11669);
or U13758 (N_13758,N_10664,N_11402);
and U13759 (N_13759,N_11745,N_11009);
xor U13760 (N_13760,N_11824,N_10699);
xnor U13761 (N_13761,N_11437,N_10298);
nand U13762 (N_13762,N_11747,N_10800);
nand U13763 (N_13763,N_10361,N_10038);
and U13764 (N_13764,N_10652,N_11419);
nor U13765 (N_13765,N_10846,N_11971);
nor U13766 (N_13766,N_11765,N_10685);
xnor U13767 (N_13767,N_11691,N_10308);
and U13768 (N_13768,N_11150,N_10326);
xnor U13769 (N_13769,N_11269,N_11807);
nor U13770 (N_13770,N_11203,N_11461);
nand U13771 (N_13771,N_10626,N_11577);
or U13772 (N_13772,N_11668,N_10657);
or U13773 (N_13773,N_10020,N_10228);
nand U13774 (N_13774,N_11039,N_10645);
xor U13775 (N_13775,N_11701,N_10668);
xnor U13776 (N_13776,N_11476,N_10078);
nand U13777 (N_13777,N_10766,N_11540);
or U13778 (N_13778,N_11414,N_10826);
nand U13779 (N_13779,N_10566,N_10121);
xor U13780 (N_13780,N_10787,N_10718);
and U13781 (N_13781,N_10433,N_10679);
xnor U13782 (N_13782,N_10879,N_10263);
and U13783 (N_13783,N_11147,N_10227);
nand U13784 (N_13784,N_10112,N_11874);
or U13785 (N_13785,N_10087,N_11076);
xnor U13786 (N_13786,N_11589,N_11439);
or U13787 (N_13787,N_10170,N_11876);
xor U13788 (N_13788,N_11330,N_10608);
nor U13789 (N_13789,N_10594,N_10346);
nand U13790 (N_13790,N_10397,N_10104);
or U13791 (N_13791,N_10397,N_10218);
xnor U13792 (N_13792,N_10752,N_11949);
xnor U13793 (N_13793,N_10782,N_10308);
xor U13794 (N_13794,N_10638,N_11847);
or U13795 (N_13795,N_11316,N_11931);
and U13796 (N_13796,N_10552,N_10449);
nor U13797 (N_13797,N_11493,N_11468);
or U13798 (N_13798,N_10823,N_11708);
or U13799 (N_13799,N_10529,N_11978);
nor U13800 (N_13800,N_10013,N_10809);
or U13801 (N_13801,N_11976,N_11297);
and U13802 (N_13802,N_11420,N_11479);
nor U13803 (N_13803,N_11881,N_10963);
nor U13804 (N_13804,N_10170,N_10086);
xnor U13805 (N_13805,N_11206,N_11021);
and U13806 (N_13806,N_11952,N_10064);
nor U13807 (N_13807,N_10301,N_10481);
xnor U13808 (N_13808,N_11787,N_11944);
or U13809 (N_13809,N_10517,N_10330);
or U13810 (N_13810,N_10043,N_10479);
or U13811 (N_13811,N_10856,N_10259);
nand U13812 (N_13812,N_11282,N_10747);
nor U13813 (N_13813,N_10775,N_10591);
nand U13814 (N_13814,N_10084,N_10676);
nor U13815 (N_13815,N_11432,N_11301);
nand U13816 (N_13816,N_11640,N_10958);
xnor U13817 (N_13817,N_10161,N_10264);
xor U13818 (N_13818,N_11231,N_10642);
or U13819 (N_13819,N_11028,N_10476);
and U13820 (N_13820,N_10810,N_10161);
nand U13821 (N_13821,N_11484,N_11955);
and U13822 (N_13822,N_11838,N_11201);
nor U13823 (N_13823,N_10242,N_10463);
nand U13824 (N_13824,N_10145,N_10796);
nor U13825 (N_13825,N_11457,N_11602);
nor U13826 (N_13826,N_11057,N_11555);
xor U13827 (N_13827,N_11030,N_10711);
nand U13828 (N_13828,N_10049,N_11898);
and U13829 (N_13829,N_10377,N_11114);
or U13830 (N_13830,N_10273,N_10518);
nor U13831 (N_13831,N_10693,N_11746);
nor U13832 (N_13832,N_10494,N_10793);
or U13833 (N_13833,N_11025,N_10575);
or U13834 (N_13834,N_11689,N_10528);
and U13835 (N_13835,N_10640,N_10839);
or U13836 (N_13836,N_10208,N_11554);
or U13837 (N_13837,N_10891,N_10021);
nor U13838 (N_13838,N_11293,N_10657);
or U13839 (N_13839,N_11518,N_10375);
nand U13840 (N_13840,N_10825,N_11071);
nand U13841 (N_13841,N_11287,N_11505);
nand U13842 (N_13842,N_11774,N_10418);
nor U13843 (N_13843,N_10907,N_11383);
xor U13844 (N_13844,N_10625,N_10258);
nor U13845 (N_13845,N_10121,N_10434);
and U13846 (N_13846,N_10421,N_10265);
nor U13847 (N_13847,N_10173,N_11690);
nand U13848 (N_13848,N_10768,N_10693);
and U13849 (N_13849,N_10189,N_10612);
or U13850 (N_13850,N_10151,N_10281);
nand U13851 (N_13851,N_10790,N_10802);
xor U13852 (N_13852,N_11652,N_10073);
nor U13853 (N_13853,N_11988,N_10952);
or U13854 (N_13854,N_11124,N_11741);
and U13855 (N_13855,N_10135,N_11540);
nor U13856 (N_13856,N_10712,N_10647);
and U13857 (N_13857,N_11139,N_10386);
xnor U13858 (N_13858,N_11591,N_11624);
xor U13859 (N_13859,N_11160,N_11963);
nor U13860 (N_13860,N_10863,N_10734);
and U13861 (N_13861,N_10765,N_10442);
or U13862 (N_13862,N_10150,N_11163);
or U13863 (N_13863,N_11280,N_10669);
xnor U13864 (N_13864,N_11633,N_11474);
xor U13865 (N_13865,N_11126,N_10360);
nand U13866 (N_13866,N_10166,N_10148);
xnor U13867 (N_13867,N_10670,N_11931);
or U13868 (N_13868,N_11558,N_10730);
nand U13869 (N_13869,N_11424,N_11595);
and U13870 (N_13870,N_10139,N_11228);
nand U13871 (N_13871,N_11450,N_10459);
and U13872 (N_13872,N_10550,N_10609);
xnor U13873 (N_13873,N_10579,N_10096);
xor U13874 (N_13874,N_10477,N_11227);
xnor U13875 (N_13875,N_10207,N_10068);
xor U13876 (N_13876,N_11656,N_11890);
xor U13877 (N_13877,N_11500,N_10094);
and U13878 (N_13878,N_10006,N_10175);
xor U13879 (N_13879,N_11560,N_10710);
nor U13880 (N_13880,N_10713,N_10929);
xnor U13881 (N_13881,N_11491,N_11178);
nand U13882 (N_13882,N_10421,N_11030);
or U13883 (N_13883,N_11249,N_10124);
or U13884 (N_13884,N_10451,N_11320);
or U13885 (N_13885,N_11592,N_10373);
and U13886 (N_13886,N_11541,N_11438);
nor U13887 (N_13887,N_10242,N_10502);
xor U13888 (N_13888,N_11817,N_10269);
nor U13889 (N_13889,N_11877,N_11715);
and U13890 (N_13890,N_10625,N_10682);
and U13891 (N_13891,N_10716,N_11994);
nor U13892 (N_13892,N_10087,N_11321);
xnor U13893 (N_13893,N_11884,N_10948);
nor U13894 (N_13894,N_10777,N_10500);
nor U13895 (N_13895,N_10655,N_11084);
or U13896 (N_13896,N_11157,N_10671);
or U13897 (N_13897,N_10918,N_10945);
and U13898 (N_13898,N_10543,N_11803);
xor U13899 (N_13899,N_11557,N_10569);
or U13900 (N_13900,N_11250,N_10145);
and U13901 (N_13901,N_11153,N_10630);
or U13902 (N_13902,N_10333,N_10935);
nor U13903 (N_13903,N_10149,N_10490);
nor U13904 (N_13904,N_11078,N_11126);
xnor U13905 (N_13905,N_11665,N_11009);
or U13906 (N_13906,N_10898,N_11221);
xnor U13907 (N_13907,N_10800,N_11229);
xnor U13908 (N_13908,N_11678,N_10375);
or U13909 (N_13909,N_11366,N_11432);
nand U13910 (N_13910,N_11531,N_11155);
and U13911 (N_13911,N_10934,N_11590);
xnor U13912 (N_13912,N_11285,N_10226);
or U13913 (N_13913,N_10803,N_10070);
and U13914 (N_13914,N_11175,N_11238);
or U13915 (N_13915,N_10063,N_10261);
or U13916 (N_13916,N_11690,N_10599);
xor U13917 (N_13917,N_11017,N_11834);
and U13918 (N_13918,N_11912,N_11962);
and U13919 (N_13919,N_10321,N_10683);
or U13920 (N_13920,N_10707,N_10115);
xnor U13921 (N_13921,N_11516,N_11880);
or U13922 (N_13922,N_11758,N_10217);
xnor U13923 (N_13923,N_11570,N_11404);
nand U13924 (N_13924,N_10659,N_11801);
nand U13925 (N_13925,N_11365,N_10013);
nor U13926 (N_13926,N_10132,N_10078);
nor U13927 (N_13927,N_11958,N_10379);
nand U13928 (N_13928,N_11151,N_10769);
nand U13929 (N_13929,N_10068,N_11268);
nor U13930 (N_13930,N_10850,N_10834);
and U13931 (N_13931,N_11896,N_11344);
xnor U13932 (N_13932,N_11892,N_10250);
xor U13933 (N_13933,N_11318,N_10161);
or U13934 (N_13934,N_10717,N_10998);
and U13935 (N_13935,N_10756,N_11324);
xor U13936 (N_13936,N_11275,N_11150);
or U13937 (N_13937,N_11640,N_10542);
nor U13938 (N_13938,N_10421,N_10137);
or U13939 (N_13939,N_10838,N_10193);
xor U13940 (N_13940,N_10647,N_11858);
nor U13941 (N_13941,N_11032,N_10745);
and U13942 (N_13942,N_11383,N_11735);
nand U13943 (N_13943,N_10448,N_11260);
nand U13944 (N_13944,N_10126,N_10770);
and U13945 (N_13945,N_11253,N_10411);
or U13946 (N_13946,N_11451,N_10848);
nor U13947 (N_13947,N_11281,N_11067);
nand U13948 (N_13948,N_10305,N_10043);
xor U13949 (N_13949,N_11780,N_11582);
xor U13950 (N_13950,N_11695,N_11887);
xnor U13951 (N_13951,N_11063,N_10841);
and U13952 (N_13952,N_10662,N_11607);
and U13953 (N_13953,N_10212,N_10259);
nor U13954 (N_13954,N_11914,N_10768);
or U13955 (N_13955,N_10553,N_11314);
nor U13956 (N_13956,N_11749,N_11518);
xor U13957 (N_13957,N_10139,N_11936);
and U13958 (N_13958,N_11217,N_10662);
nand U13959 (N_13959,N_10525,N_10344);
nand U13960 (N_13960,N_11979,N_11972);
xor U13961 (N_13961,N_10015,N_11513);
and U13962 (N_13962,N_10342,N_11606);
nand U13963 (N_13963,N_10870,N_11253);
nor U13964 (N_13964,N_11428,N_11831);
nor U13965 (N_13965,N_10428,N_10244);
nor U13966 (N_13966,N_10301,N_11129);
xor U13967 (N_13967,N_10448,N_11244);
nand U13968 (N_13968,N_10236,N_11806);
nand U13969 (N_13969,N_11715,N_10638);
nor U13970 (N_13970,N_11118,N_11285);
and U13971 (N_13971,N_10976,N_10286);
nor U13972 (N_13972,N_11301,N_10020);
nand U13973 (N_13973,N_11203,N_10981);
xor U13974 (N_13974,N_10510,N_10847);
nand U13975 (N_13975,N_11224,N_10602);
nand U13976 (N_13976,N_10563,N_10053);
or U13977 (N_13977,N_11040,N_11412);
or U13978 (N_13978,N_10940,N_10043);
nor U13979 (N_13979,N_11648,N_10181);
or U13980 (N_13980,N_11614,N_10599);
nand U13981 (N_13981,N_11199,N_11413);
or U13982 (N_13982,N_11803,N_11485);
nor U13983 (N_13983,N_11845,N_10012);
xor U13984 (N_13984,N_10997,N_11049);
xnor U13985 (N_13985,N_10644,N_10298);
nand U13986 (N_13986,N_10451,N_10432);
xnor U13987 (N_13987,N_11081,N_11379);
xnor U13988 (N_13988,N_11527,N_11549);
nand U13989 (N_13989,N_10736,N_10996);
xor U13990 (N_13990,N_10360,N_10269);
and U13991 (N_13991,N_11356,N_10977);
nor U13992 (N_13992,N_11672,N_10122);
or U13993 (N_13993,N_11173,N_11666);
and U13994 (N_13994,N_10326,N_11118);
xor U13995 (N_13995,N_11084,N_11429);
nand U13996 (N_13996,N_11871,N_10840);
or U13997 (N_13997,N_10596,N_11720);
nor U13998 (N_13998,N_10391,N_11913);
nand U13999 (N_13999,N_10679,N_10719);
or U14000 (N_14000,N_13598,N_13243);
and U14001 (N_14001,N_12908,N_12670);
xor U14002 (N_14002,N_13068,N_12888);
nor U14003 (N_14003,N_12357,N_12366);
nor U14004 (N_14004,N_13400,N_13135);
or U14005 (N_14005,N_13700,N_12781);
and U14006 (N_14006,N_12803,N_12764);
nor U14007 (N_14007,N_12875,N_13547);
nor U14008 (N_14008,N_12899,N_12337);
xnor U14009 (N_14009,N_13620,N_12805);
or U14010 (N_14010,N_13444,N_12237);
xnor U14011 (N_14011,N_12240,N_13744);
nor U14012 (N_14012,N_12647,N_13080);
and U14013 (N_14013,N_12548,N_12308);
nor U14014 (N_14014,N_12198,N_13706);
and U14015 (N_14015,N_13174,N_13915);
nand U14016 (N_14016,N_12913,N_12189);
nand U14017 (N_14017,N_13719,N_12173);
or U14018 (N_14018,N_13951,N_12649);
xnor U14019 (N_14019,N_12638,N_12207);
or U14020 (N_14020,N_12511,N_12686);
nor U14021 (N_14021,N_13750,N_12613);
nor U14022 (N_14022,N_13844,N_13156);
xor U14023 (N_14023,N_12313,N_12573);
or U14024 (N_14024,N_12767,N_12364);
nand U14025 (N_14025,N_13064,N_12255);
nand U14026 (N_14026,N_13587,N_13989);
or U14027 (N_14027,N_13786,N_13623);
or U14028 (N_14028,N_12377,N_12397);
and U14029 (N_14029,N_12598,N_12792);
xnor U14030 (N_14030,N_12859,N_12137);
nand U14031 (N_14031,N_12810,N_12201);
or U14032 (N_14032,N_13026,N_12321);
and U14033 (N_14033,N_13416,N_13000);
nand U14034 (N_14034,N_13248,N_12244);
nor U14035 (N_14035,N_13987,N_12095);
and U14036 (N_14036,N_12532,N_13297);
and U14037 (N_14037,N_13211,N_12685);
xnor U14038 (N_14038,N_12303,N_13647);
or U14039 (N_14039,N_13874,N_13943);
or U14040 (N_14040,N_12170,N_13290);
nor U14041 (N_14041,N_12442,N_12980);
or U14042 (N_14042,N_13770,N_13425);
nand U14043 (N_14043,N_12657,N_12790);
and U14044 (N_14044,N_13670,N_12746);
xnor U14045 (N_14045,N_13338,N_12640);
nor U14046 (N_14046,N_13690,N_13116);
nor U14047 (N_14047,N_13194,N_12384);
and U14048 (N_14048,N_13346,N_13776);
or U14049 (N_14049,N_12452,N_13573);
xnor U14050 (N_14050,N_13809,N_13308);
nand U14051 (N_14051,N_12334,N_13845);
or U14052 (N_14052,N_12236,N_13823);
or U14053 (N_14053,N_12493,N_13164);
and U14054 (N_14054,N_13457,N_12820);
or U14055 (N_14055,N_13489,N_13223);
nand U14056 (N_14056,N_12969,N_12411);
or U14057 (N_14057,N_12560,N_12759);
and U14058 (N_14058,N_12542,N_12033);
or U14059 (N_14059,N_13752,N_13885);
nor U14060 (N_14060,N_12512,N_13315);
xnor U14061 (N_14061,N_12341,N_13998);
and U14062 (N_14062,N_13610,N_13274);
nor U14063 (N_14063,N_12077,N_12645);
xor U14064 (N_14064,N_12401,N_13242);
and U14065 (N_14065,N_13258,N_12043);
nand U14066 (N_14066,N_13749,N_12571);
and U14067 (N_14067,N_13143,N_13863);
and U14068 (N_14068,N_12580,N_13394);
nor U14069 (N_14069,N_12404,N_12449);
nor U14070 (N_14070,N_13365,N_13353);
and U14071 (N_14071,N_13238,N_12656);
xor U14072 (N_14072,N_13603,N_12249);
and U14073 (N_14073,N_13890,N_13284);
nor U14074 (N_14074,N_13761,N_12338);
xnor U14075 (N_14075,N_13254,N_12842);
or U14076 (N_14076,N_13453,N_12831);
nand U14077 (N_14077,N_12241,N_12109);
xor U14078 (N_14078,N_13138,N_12713);
or U14079 (N_14079,N_12959,N_12729);
and U14080 (N_14080,N_13569,N_13664);
and U14081 (N_14081,N_13282,N_13960);
nand U14082 (N_14082,N_12434,N_12763);
or U14083 (N_14083,N_13168,N_13491);
or U14084 (N_14084,N_12912,N_13183);
or U14085 (N_14085,N_12127,N_12565);
or U14086 (N_14086,N_12497,N_13411);
xnor U14087 (N_14087,N_12001,N_13437);
and U14088 (N_14088,N_13165,N_12163);
and U14089 (N_14089,N_12932,N_12225);
nor U14090 (N_14090,N_13972,N_12678);
nand U14091 (N_14091,N_13013,N_12925);
xnor U14092 (N_14092,N_13436,N_13538);
xor U14093 (N_14093,N_13182,N_13339);
nor U14094 (N_14094,N_12305,N_12957);
and U14095 (N_14095,N_12426,N_12011);
and U14096 (N_14096,N_12361,N_12048);
nand U14097 (N_14097,N_12468,N_12438);
or U14098 (N_14098,N_13644,N_13358);
xor U14099 (N_14099,N_13060,N_13025);
nand U14100 (N_14100,N_13144,N_13604);
and U14101 (N_14101,N_12292,N_12075);
xor U14102 (N_14102,N_12986,N_12193);
xnor U14103 (N_14103,N_12360,N_13220);
or U14104 (N_14104,N_12020,N_13506);
xor U14105 (N_14105,N_12607,N_12226);
nand U14106 (N_14106,N_13551,N_12402);
nor U14107 (N_14107,N_12262,N_12787);
nand U14108 (N_14108,N_12427,N_12687);
nand U14109 (N_14109,N_12435,N_13558);
and U14110 (N_14110,N_13628,N_13084);
nand U14111 (N_14111,N_13104,N_13663);
nor U14112 (N_14112,N_12168,N_13775);
nand U14113 (N_14113,N_13218,N_13379);
nand U14114 (N_14114,N_12002,N_13130);
nor U14115 (N_14115,N_13800,N_13682);
nor U14116 (N_14116,N_13197,N_12040);
xor U14117 (N_14117,N_13591,N_13709);
or U14118 (N_14118,N_12692,N_13461);
or U14119 (N_14119,N_13643,N_12393);
or U14120 (N_14120,N_12926,N_13513);
nor U14121 (N_14121,N_12467,N_12280);
nand U14122 (N_14122,N_13203,N_12462);
or U14123 (N_14123,N_12381,N_13237);
xnor U14124 (N_14124,N_13184,N_12806);
and U14125 (N_14125,N_13853,N_12794);
or U14126 (N_14126,N_13291,N_12761);
xnor U14127 (N_14127,N_13917,N_12741);
xnor U14128 (N_14128,N_12348,N_12501);
nor U14129 (N_14129,N_13110,N_12588);
and U14130 (N_14130,N_12725,N_12443);
and U14131 (N_14131,N_12190,N_12116);
nand U14132 (N_14132,N_12715,N_12504);
and U14133 (N_14133,N_12601,N_13925);
nor U14134 (N_14134,N_12674,N_13902);
nand U14135 (N_14135,N_12537,N_13503);
and U14136 (N_14136,N_13128,N_12391);
or U14137 (N_14137,N_13153,N_13313);
and U14138 (N_14138,N_12574,N_12703);
xor U14139 (N_14139,N_13798,N_12306);
and U14140 (N_14140,N_12895,N_12138);
xnor U14141 (N_14141,N_12429,N_12486);
nor U14142 (N_14142,N_13751,N_12967);
nor U14143 (N_14143,N_12270,N_12707);
nand U14144 (N_14144,N_13772,N_12133);
or U14145 (N_14145,N_13660,N_12775);
xnor U14146 (N_14146,N_12835,N_12094);
or U14147 (N_14147,N_12883,N_12463);
xor U14148 (N_14148,N_12609,N_12708);
or U14149 (N_14149,N_12086,N_13518);
or U14150 (N_14150,N_13426,N_12330);
nor U14151 (N_14151,N_12832,N_12227);
or U14152 (N_14152,N_13970,N_13947);
xnor U14153 (N_14153,N_12522,N_13012);
and U14154 (N_14154,N_12526,N_13460);
nand U14155 (N_14155,N_13697,N_13415);
nor U14156 (N_14156,N_13973,N_12785);
or U14157 (N_14157,N_12375,N_12917);
nand U14158 (N_14158,N_13650,N_12057);
and U14159 (N_14159,N_12331,N_12887);
or U14160 (N_14160,N_13961,N_12242);
nor U14161 (N_14161,N_13901,N_13119);
nand U14162 (N_14162,N_12166,N_13510);
or U14163 (N_14163,N_12160,N_12049);
xor U14164 (N_14164,N_13967,N_12065);
nor U14165 (N_14165,N_12108,N_13031);
xor U14166 (N_14166,N_12010,N_12762);
xor U14167 (N_14167,N_12815,N_13757);
nand U14168 (N_14168,N_12705,N_13954);
xor U14169 (N_14169,N_12460,N_13819);
nand U14170 (N_14170,N_13993,N_12162);
and U14171 (N_14171,N_13482,N_13364);
nor U14172 (N_14172,N_13396,N_13142);
nand U14173 (N_14173,N_13196,N_12555);
and U14174 (N_14174,N_12490,N_12045);
xnor U14175 (N_14175,N_13523,N_13913);
nand U14176 (N_14176,N_13790,N_12218);
xor U14177 (N_14177,N_12431,N_13803);
and U14178 (N_14178,N_13494,N_13198);
nor U14179 (N_14179,N_13893,N_13383);
nor U14180 (N_14180,N_13377,N_12952);
and U14181 (N_14181,N_13011,N_12693);
or U14182 (N_14182,N_13410,N_13115);
nor U14183 (N_14183,N_13386,N_12389);
and U14184 (N_14184,N_12216,N_13492);
and U14185 (N_14185,N_13337,N_13134);
xnor U14186 (N_14186,N_12791,N_13016);
or U14187 (N_14187,N_12250,N_13382);
nor U14188 (N_14188,N_12689,N_12720);
nand U14189 (N_14189,N_12266,N_12437);
and U14190 (N_14190,N_13795,N_12985);
nor U14191 (N_14191,N_13361,N_13695);
nand U14192 (N_14192,N_12727,N_13428);
or U14193 (N_14193,N_12646,N_12372);
xnor U14194 (N_14194,N_12850,N_13722);
and U14195 (N_14195,N_12854,N_13368);
xor U14196 (N_14196,N_13009,N_13688);
or U14197 (N_14197,N_13317,N_13930);
or U14198 (N_14198,N_13300,N_13816);
or U14199 (N_14199,N_13859,N_12386);
xor U14200 (N_14200,N_12058,N_13497);
or U14201 (N_14201,N_13720,N_13662);
nand U14202 (N_14202,N_12596,N_13945);
nor U14203 (N_14203,N_12891,N_13439);
and U14204 (N_14204,N_12824,N_12695);
nand U14205 (N_14205,N_12398,N_12996);
or U14206 (N_14206,N_12858,N_13575);
nor U14207 (N_14207,N_13570,N_12873);
and U14208 (N_14208,N_13637,N_12484);
or U14209 (N_14209,N_12079,N_12205);
xor U14210 (N_14210,N_12871,N_13023);
nor U14211 (N_14211,N_13981,N_13600);
and U14212 (N_14212,N_13306,N_13672);
nand U14213 (N_14213,N_12740,N_12317);
nand U14214 (N_14214,N_13081,N_12325);
xor U14215 (N_14215,N_13057,N_12071);
and U14216 (N_14216,N_12901,N_12737);
nand U14217 (N_14217,N_12167,N_13092);
xor U14218 (N_14218,N_12634,N_13824);
xor U14219 (N_14219,N_12903,N_13431);
and U14220 (N_14220,N_12704,N_13043);
and U14221 (N_14221,N_12714,N_12298);
nand U14222 (N_14222,N_13543,N_12149);
or U14223 (N_14223,N_13735,N_13154);
and U14224 (N_14224,N_13272,N_13122);
xnor U14225 (N_14225,N_13384,N_12852);
or U14226 (N_14226,N_13319,N_13469);
or U14227 (N_14227,N_12754,N_13742);
xnor U14228 (N_14228,N_12320,N_12099);
xnor U14229 (N_14229,N_12874,N_13424);
and U14230 (N_14230,N_12973,N_13657);
nor U14231 (N_14231,N_13381,N_13454);
nand U14232 (N_14232,N_13818,N_13283);
nand U14233 (N_14233,N_13030,N_12157);
or U14234 (N_14234,N_13099,N_12845);
xnor U14235 (N_14235,N_12736,N_12184);
nand U14236 (N_14236,N_12476,N_13159);
nor U14237 (N_14237,N_12159,N_12546);
nand U14238 (N_14238,N_13162,N_13160);
xor U14239 (N_14239,N_13208,N_12788);
and U14240 (N_14240,N_13257,N_12808);
xnor U14241 (N_14241,N_12374,N_12644);
or U14242 (N_14242,N_13225,N_13783);
and U14243 (N_14243,N_12827,N_13810);
nand U14244 (N_14244,N_13926,N_13785);
xor U14245 (N_14245,N_12456,N_13251);
nor U14246 (N_14246,N_12698,N_12963);
nand U14247 (N_14247,N_13033,N_13204);
or U14248 (N_14248,N_12822,N_12572);
and U14249 (N_14249,N_13347,N_12067);
xor U14250 (N_14250,N_12515,N_12648);
or U14251 (N_14251,N_12395,N_12194);
or U14252 (N_14252,N_12221,N_13541);
or U14253 (N_14253,N_12091,N_13330);
and U14254 (N_14254,N_13141,N_12552);
nand U14255 (N_14255,N_13509,N_13342);
and U14256 (N_14256,N_12628,N_13875);
xor U14257 (N_14257,N_12641,N_13679);
and U14258 (N_14258,N_13597,N_13774);
nand U14259 (N_14259,N_12039,N_12481);
and U14260 (N_14260,N_13638,N_12651);
xor U14261 (N_14261,N_13071,N_13360);
or U14262 (N_14262,N_12230,N_13487);
xnor U14263 (N_14263,N_13617,N_12951);
xnor U14264 (N_14264,N_12088,N_12066);
nor U14265 (N_14265,N_12614,N_13350);
and U14266 (N_14266,N_13027,N_12448);
nor U14267 (N_14267,N_12921,N_12885);
xor U14268 (N_14268,N_12283,N_13864);
and U14269 (N_14269,N_12502,N_13440);
and U14270 (N_14270,N_12367,N_13892);
and U14271 (N_14271,N_13498,N_12282);
and U14272 (N_14272,N_13354,N_12399);
and U14273 (N_14273,N_13086,N_12096);
and U14274 (N_14274,N_13515,N_12639);
and U14275 (N_14275,N_13804,N_12724);
xor U14276 (N_14276,N_12275,N_13255);
nand U14277 (N_14277,N_13937,N_12626);
nor U14278 (N_14278,N_12751,N_12735);
and U14279 (N_14279,N_12121,N_12022);
or U14280 (N_14280,N_12425,N_13029);
or U14281 (N_14281,N_13769,N_13979);
xnor U14282 (N_14282,N_13574,N_12749);
nor U14283 (N_14283,N_12106,N_12709);
nand U14284 (N_14284,N_12793,N_12405);
and U14285 (N_14285,N_12879,N_13992);
xnor U14286 (N_14286,N_12999,N_13516);
or U14287 (N_14287,N_13070,N_13019);
nand U14288 (N_14288,N_13352,N_12018);
or U14289 (N_14289,N_13699,N_13152);
or U14290 (N_14290,N_12529,N_13626);
nor U14291 (N_14291,N_13234,N_12107);
and U14292 (N_14292,N_13097,N_12451);
and U14293 (N_14293,N_13676,N_12445);
xnor U14294 (N_14294,N_13921,N_13683);
nor U14295 (N_14295,N_13422,N_13727);
nor U14296 (N_14296,N_13959,N_13613);
xnor U14297 (N_14297,N_12606,N_13734);
xor U14298 (N_14298,N_13999,N_12310);
or U14299 (N_14299,N_13402,N_12930);
nor U14300 (N_14300,N_12368,N_13414);
and U14301 (N_14301,N_12281,N_12929);
nand U14302 (N_14302,N_13273,N_13805);
or U14303 (N_14303,N_13256,N_12579);
nand U14304 (N_14304,N_13554,N_13519);
nor U14305 (N_14305,N_12217,N_12302);
nand U14306 (N_14306,N_12347,N_12892);
xnor U14307 (N_14307,N_13227,N_13836);
xor U14308 (N_14308,N_12365,N_12800);
nand U14309 (N_14309,N_13903,N_13696);
or U14310 (N_14310,N_13589,N_12524);
or U14311 (N_14311,N_13166,N_13567);
nand U14312 (N_14312,N_12956,N_12510);
xnor U14313 (N_14313,N_13686,N_12474);
nand U14314 (N_14314,N_12072,N_13262);
nand U14315 (N_14315,N_12514,N_12717);
nor U14316 (N_14316,N_12436,N_13828);
nor U14317 (N_14317,N_12680,N_13740);
nand U14318 (N_14318,N_12506,N_13525);
or U14319 (N_14319,N_13843,N_13899);
nor U14320 (N_14320,N_13149,N_13034);
nand U14321 (N_14321,N_12177,N_12642);
or U14322 (N_14322,N_12706,N_12097);
xnor U14323 (N_14323,N_13991,N_12183);
nand U14324 (N_14324,N_13546,N_13118);
or U14325 (N_14325,N_13045,N_12046);
nand U14326 (N_14326,N_12587,N_12654);
or U14327 (N_14327,N_12721,N_13674);
nor U14328 (N_14328,N_12556,N_12830);
xor U14329 (N_14329,N_13145,N_12605);
xor U14330 (N_14330,N_13172,N_13213);
xor U14331 (N_14331,N_13565,N_13148);
nor U14332 (N_14332,N_12770,N_13181);
nor U14333 (N_14333,N_13348,N_12599);
nor U14334 (N_14334,N_12156,N_13260);
nor U14335 (N_14335,N_13655,N_13830);
nand U14336 (N_14336,N_13106,N_13847);
xor U14337 (N_14337,N_12344,N_13754);
and U14338 (N_14338,N_13388,N_13420);
nand U14339 (N_14339,N_13759,N_13421);
or U14340 (N_14340,N_13015,N_13710);
and U14341 (N_14341,N_13579,N_13002);
and U14342 (N_14342,N_12152,N_13179);
xor U14343 (N_14343,N_13356,N_13187);
and U14344 (N_14344,N_13840,N_13867);
and U14345 (N_14345,N_13656,N_12894);
and U14346 (N_14346,N_13233,N_12898);
or U14347 (N_14347,N_12134,N_13708);
and U14348 (N_14348,N_12979,N_13292);
nor U14349 (N_14349,N_12471,N_13821);
nand U14350 (N_14350,N_13933,N_13661);
or U14351 (N_14351,N_13521,N_13778);
nand U14352 (N_14352,N_12119,N_13059);
xor U14353 (N_14353,N_13528,N_12944);
or U14354 (N_14354,N_13268,N_13161);
xnor U14355 (N_14355,N_12487,N_12750);
or U14356 (N_14356,N_13044,N_13500);
nand U14357 (N_14357,N_12329,N_13533);
or U14358 (N_14358,N_12976,N_12795);
and U14359 (N_14359,N_13773,N_13985);
nor U14360 (N_14360,N_13441,N_13111);
nand U14361 (N_14361,N_12450,N_12440);
xor U14362 (N_14362,N_13607,N_13802);
or U14363 (N_14363,N_12652,N_12323);
and U14364 (N_14364,N_12379,N_12410);
nor U14365 (N_14365,N_12991,N_12618);
or U14366 (N_14366,N_13455,N_13737);
nand U14367 (N_14367,N_12439,N_12733);
nor U14368 (N_14368,N_12132,N_12297);
or U14369 (N_14369,N_12195,N_13814);
xnor U14370 (N_14370,N_12843,N_13698);
nor U14371 (N_14371,N_13053,N_12837);
nand U14372 (N_14372,N_12286,N_13990);
and U14373 (N_14373,N_12783,N_12161);
xor U14374 (N_14374,N_13689,N_13561);
or U14375 (N_14375,N_13239,N_13496);
or U14376 (N_14376,N_13910,N_12600);
xnor U14377 (N_14377,N_12235,N_13493);
and U14378 (N_14378,N_13288,N_12307);
or U14379 (N_14379,N_13630,N_12044);
xor U14380 (N_14380,N_13555,N_12905);
nand U14381 (N_14381,N_13862,N_13878);
xnor U14382 (N_14382,N_12359,N_13355);
nor U14383 (N_14383,N_12014,N_13595);
and U14384 (N_14384,N_12472,N_13854);
nand U14385 (N_14385,N_13395,N_13851);
nor U14386 (N_14386,N_12219,N_13247);
xor U14387 (N_14387,N_12540,N_12718);
xor U14388 (N_14388,N_12016,N_13488);
or U14389 (N_14389,N_12535,N_12103);
nor U14390 (N_14390,N_12866,N_12061);
xnor U14391 (N_14391,N_12910,N_13711);
and U14392 (N_14392,N_12145,N_13504);
or U14393 (N_14393,N_12355,N_12690);
nor U14394 (N_14394,N_12861,N_13564);
or U14395 (N_14395,N_12592,N_12433);
nor U14396 (N_14396,N_13340,N_13462);
and U14397 (N_14397,N_13940,N_12615);
xor U14398 (N_14398,N_12576,N_12153);
xor U14399 (N_14399,N_13559,N_12259);
xor U14400 (N_14400,N_13185,N_13036);
nor U14401 (N_14401,N_13124,N_13920);
or U14402 (N_14402,N_12475,N_13612);
xor U14403 (N_14403,N_12739,N_12455);
nor U14404 (N_14404,N_12804,N_12878);
nor U14405 (N_14405,N_13922,N_13642);
and U14406 (N_14406,N_12661,N_12796);
and U14407 (N_14407,N_13017,N_13052);
xor U14408 (N_14408,N_13797,N_12684);
nor U14409 (N_14409,N_13677,N_13884);
or U14410 (N_14410,N_13404,N_12319);
nand U14411 (N_14411,N_13877,N_13965);
xor U14412 (N_14412,N_12035,N_12446);
xor U14413 (N_14413,N_13267,N_13614);
or U14414 (N_14414,N_12054,N_13950);
nand U14415 (N_14415,N_13067,N_12557);
nand U14416 (N_14416,N_13850,N_13812);
or U14417 (N_14417,N_12937,N_12232);
and U14418 (N_14418,N_13310,N_12336);
or U14419 (N_14419,N_12383,N_13536);
or U14420 (N_14420,N_13083,N_12350);
and U14421 (N_14421,N_12594,N_13856);
xnor U14422 (N_14422,N_13007,N_12243);
xnor U14423 (N_14423,N_12568,N_13409);
or U14424 (N_14424,N_13188,N_12773);
xnor U14425 (N_14425,N_12478,N_13611);
nand U14426 (N_14426,N_13280,N_12738);
nor U14427 (N_14427,N_13594,N_13327);
xor U14428 (N_14428,N_13584,N_12853);
xor U14429 (N_14429,N_12882,N_13171);
nor U14430 (N_14430,N_13216,N_12073);
xor U14431 (N_14431,N_13934,N_13219);
and U14432 (N_14432,N_13517,N_13433);
or U14433 (N_14433,N_13667,N_12633);
and U14434 (N_14434,N_12087,N_13351);
nor U14435 (N_14435,N_13540,N_12730);
nand U14436 (N_14436,N_13235,N_13296);
or U14437 (N_14437,N_12516,N_13881);
nand U14438 (N_14438,N_13527,N_12978);
and U14439 (N_14439,N_12688,N_12696);
or U14440 (N_14440,N_12060,N_12616);
nor U14441 (N_14441,N_13429,N_13393);
and U14442 (N_14442,N_12766,N_13833);
nor U14443 (N_14443,N_13855,N_13944);
xnor U14444 (N_14444,N_12977,N_12051);
xor U14445 (N_14445,N_12777,N_13784);
nor U14446 (N_14446,N_13245,N_12483);
nor U14447 (N_14447,N_13467,N_12176);
nor U14448 (N_14448,N_12821,N_13984);
xnor U14449 (N_14449,N_12916,N_13037);
nand U14450 (N_14450,N_12256,N_13003);
and U14451 (N_14451,N_13852,N_13725);
nor U14452 (N_14452,N_12954,N_13051);
or U14453 (N_14453,N_12291,N_12264);
nand U14454 (N_14454,N_13914,N_13969);
nor U14455 (N_14455,N_12682,N_13311);
and U14456 (N_14456,N_13675,N_13841);
nand U14457 (N_14457,N_13544,N_13743);
nor U14458 (N_14458,N_12407,N_13471);
and U14459 (N_14459,N_13507,N_13103);
xor U14460 (N_14460,N_12254,N_12631);
nand U14461 (N_14461,N_12037,N_13021);
or U14462 (N_14462,N_13294,N_13264);
and U14463 (N_14463,N_12945,N_13609);
and U14464 (N_14464,N_12353,N_13250);
and U14465 (N_14465,N_12265,N_12672);
nor U14466 (N_14466,N_13636,N_13349);
and U14467 (N_14467,N_13834,N_12617);
and U14468 (N_14468,N_13745,N_12007);
or U14469 (N_14469,N_12786,N_13842);
nor U14470 (N_14470,N_12948,N_13562);
nor U14471 (N_14471,N_13090,N_13287);
nand U14472 (N_14472,N_12082,N_13793);
and U14473 (N_14473,N_12697,N_13501);
nand U14474 (N_14474,N_13894,N_12258);
or U14475 (N_14475,N_12525,N_12855);
and U14476 (N_14476,N_13694,N_12581);
xnor U14477 (N_14477,N_12995,N_12612);
nand U14478 (N_14478,N_12050,N_13946);
or U14479 (N_14479,N_13701,N_12671);
and U14480 (N_14480,N_12416,N_12120);
nand U14481 (N_14481,N_12828,N_12135);
and U14482 (N_14482,N_12760,N_12335);
nor U14483 (N_14483,N_13207,N_12424);
or U14484 (N_14484,N_13906,N_12518);
nor U14485 (N_14485,N_13646,N_13397);
and U14486 (N_14486,N_12964,N_12919);
or U14487 (N_14487,N_12772,N_13158);
or U14488 (N_14488,N_12798,N_12807);
xor U14489 (N_14489,N_12447,N_13781);
nand U14490 (N_14490,N_13687,N_12834);
and U14491 (N_14491,N_12140,N_12036);
nor U14492 (N_14492,N_12659,N_13407);
xor U14493 (N_14493,N_13935,N_12743);
nand U14494 (N_14494,N_13163,N_12131);
or U14495 (N_14495,N_13839,N_12358);
and U14496 (N_14496,N_13596,N_12199);
nor U14497 (N_14497,N_13486,N_13018);
nor U14498 (N_14498,N_13210,N_12711);
and U14499 (N_14499,N_12753,N_12078);
xnor U14500 (N_14500,N_12829,N_13837);
nor U14501 (N_14501,N_13801,N_12893);
nand U14502 (N_14502,N_12210,N_13633);
nand U14503 (N_14503,N_13055,N_12034);
nor U14504 (N_14504,N_13120,N_12586);
or U14505 (N_14505,N_12248,N_13712);
and U14506 (N_14506,N_13089,N_13072);
or U14507 (N_14507,N_13733,N_13963);
nand U14508 (N_14508,N_13514,N_13100);
or U14509 (N_14509,N_13063,N_12295);
nor U14510 (N_14510,N_12273,N_12059);
and U14511 (N_14511,N_13189,N_12547);
nand U14512 (N_14512,N_13654,N_13581);
nor U14513 (N_14513,N_12623,N_13316);
nand U14514 (N_14514,N_12083,N_13741);
nand U14515 (N_14515,N_13465,N_13868);
nor U14516 (N_14516,N_12403,N_13281);
xnor U14517 (N_14517,N_12569,N_13576);
nor U14518 (N_14518,N_12019,N_13490);
nor U14519 (N_14519,N_13094,N_12716);
xnor U14520 (N_14520,N_13448,N_13205);
xnor U14521 (N_14521,N_12585,N_13253);
xnor U14522 (N_14522,N_13117,N_12158);
or U14523 (N_14523,N_13333,N_12745);
nand U14524 (N_14524,N_13703,N_12006);
nor U14525 (N_14525,N_12257,N_13035);
nand U14526 (N_14526,N_13459,N_12562);
nand U14527 (N_14527,N_13826,N_12126);
xor U14528 (N_14528,N_13641,N_13779);
or U14529 (N_14529,N_13322,N_12987);
nor U14530 (N_14530,N_13997,N_13511);
and U14531 (N_14531,N_13178,N_13304);
xnor U14532 (N_14532,N_13666,N_13222);
or U14533 (N_14533,N_13983,N_13639);
nand U14534 (N_14534,N_12492,N_13362);
and U14535 (N_14535,N_12143,N_12268);
xnor U14536 (N_14536,N_12998,N_12550);
and U14537 (N_14537,N_13132,N_12527);
and U14538 (N_14538,N_12363,N_12234);
or U14539 (N_14539,N_12473,N_12400);
nor U14540 (N_14540,N_12136,N_13765);
nor U14541 (N_14541,N_12577,N_13872);
and U14542 (N_14542,N_12994,N_13049);
xor U14543 (N_14543,N_13066,N_12971);
xnor U14544 (N_14544,N_12085,N_13593);
or U14545 (N_14545,N_12064,N_13085);
xnor U14546 (N_14546,N_12710,N_13275);
xor U14547 (N_14547,N_13427,N_13592);
and U14548 (N_14548,N_13476,N_13345);
xor U14549 (N_14549,N_13807,N_13535);
nor U14550 (N_14550,N_13456,N_12351);
nand U14551 (N_14551,N_12677,N_12387);
xnor U14552 (N_14552,N_12142,N_13401);
xnor U14553 (N_14553,N_13209,N_13746);
nor U14554 (N_14554,N_12876,N_13056);
or U14555 (N_14555,N_12862,N_13146);
or U14556 (N_14556,N_13024,N_13726);
and U14557 (N_14557,N_12909,N_12174);
nor U14558 (N_14558,N_12857,N_13366);
xnor U14559 (N_14559,N_13048,N_12936);
xor U14560 (N_14560,N_12371,N_12069);
nand U14561 (N_14561,N_13039,N_13229);
xor U14562 (N_14562,N_13040,N_12274);
xor U14563 (N_14563,N_13096,N_12520);
or U14564 (N_14564,N_13539,N_13125);
or U14565 (N_14565,N_13109,N_13240);
and U14566 (N_14566,N_12604,N_12966);
xor U14567 (N_14567,N_12922,N_13403);
nand U14568 (N_14568,N_13825,N_12239);
xnor U14569 (N_14569,N_13820,N_13114);
nand U14570 (N_14570,N_13047,N_12042);
nor U14571 (N_14571,N_12498,N_13151);
xor U14572 (N_14572,N_13756,N_13879);
or U14573 (N_14573,N_12012,N_13615);
and U14574 (N_14574,N_13838,N_13718);
and U14575 (N_14575,N_12544,N_12856);
nor U14576 (N_14576,N_13640,N_13417);
or U14577 (N_14577,N_12277,N_13653);
or U14578 (N_14578,N_12884,N_12380);
or U14579 (N_14579,N_13483,N_12454);
and U14580 (N_14580,N_12499,N_12890);
xor U14581 (N_14581,N_12582,N_13739);
nor U14582 (N_14582,N_13897,N_12333);
xnor U14583 (N_14583,N_12208,N_12222);
or U14584 (N_14584,N_13378,N_13704);
or U14585 (N_14585,N_12940,N_13962);
and U14586 (N_14586,N_13318,N_13113);
nand U14587 (N_14587,N_13762,N_12396);
nor U14588 (N_14588,N_13276,N_13550);
nor U14589 (N_14589,N_12982,N_13298);
or U14590 (N_14590,N_12643,N_13723);
or U14591 (N_14591,N_13508,N_12927);
nand U14592 (N_14592,N_12461,N_13087);
or U14593 (N_14593,N_13767,N_13485);
and U14594 (N_14594,N_13680,N_13061);
or U14595 (N_14595,N_13957,N_12683);
xnor U14596 (N_14596,N_13811,N_13214);
nand U14597 (N_14597,N_13714,N_13974);
or U14598 (N_14598,N_13450,N_12742);
and U14599 (N_14599,N_12997,N_12287);
nor U14600 (N_14600,N_12863,N_12595);
xor U14601 (N_14601,N_13452,N_12968);
nor U14602 (N_14602,N_12056,N_13732);
or U14603 (N_14603,N_13758,N_12008);
or U14604 (N_14604,N_12147,N_13446);
xnor U14605 (N_14605,N_12326,N_13095);
nor U14606 (N_14606,N_12343,N_13817);
and U14607 (N_14607,N_13369,N_12825);
nand U14608 (N_14608,N_13705,N_13918);
and U14609 (N_14609,N_12110,N_12203);
xnor U14610 (N_14610,N_12345,N_12151);
nor U14611 (N_14611,N_13577,N_13129);
or U14612 (N_14612,N_12252,N_13911);
xnor U14613 (N_14613,N_13966,N_12053);
nor U14614 (N_14614,N_12267,N_12299);
xnor U14615 (N_14615,N_13167,N_13101);
nand U14616 (N_14616,N_12765,N_13848);
or U14617 (N_14617,N_13495,N_13470);
and U14618 (N_14618,N_12175,N_12315);
and U14619 (N_14619,N_12591,N_12611);
nor U14620 (N_14620,N_12939,N_13075);
nand U14621 (N_14621,N_12062,N_13619);
and U14622 (N_14622,N_12747,N_12112);
nor U14623 (N_14623,N_13370,N_12279);
nor U14624 (N_14624,N_13193,N_12289);
xnor U14625 (N_14625,N_13869,N_13108);
and U14626 (N_14626,N_13062,N_12839);
nor U14627 (N_14627,N_13367,N_13763);
and U14628 (N_14628,N_13731,N_13659);
nand U14629 (N_14629,N_13898,N_12660);
and U14630 (N_14630,N_12676,N_12503);
and U14631 (N_14631,N_12171,N_13190);
nand U14632 (N_14632,N_13618,N_12340);
xnor U14633 (N_14633,N_13212,N_13215);
xor U14634 (N_14634,N_12826,N_13230);
and U14635 (N_14635,N_12271,N_12477);
nand U14636 (N_14636,N_12179,N_12118);
and U14637 (N_14637,N_13861,N_13079);
xor U14638 (N_14638,N_12318,N_13375);
nor U14639 (N_14639,N_12665,N_12673);
nand U14640 (N_14640,N_12622,N_13590);
and U14641 (N_14641,N_13419,N_13932);
and U14642 (N_14642,N_13988,N_13312);
nand U14643 (N_14643,N_13912,N_12983);
and U14644 (N_14644,N_13232,N_12920);
nor U14645 (N_14645,N_12115,N_13112);
xnor U14646 (N_14646,N_12459,N_13464);
or U14647 (N_14647,N_12489,N_13293);
or U14648 (N_14648,N_12768,N_12004);
xnor U14649 (N_14649,N_13578,N_13948);
nor U14650 (N_14650,N_13526,N_13883);
nor U14651 (N_14651,N_12974,N_13996);
nor U14652 (N_14652,N_12491,N_13994);
and U14653 (N_14653,N_13792,N_13445);
nor U14654 (N_14654,N_12990,N_13952);
or U14655 (N_14655,N_12780,N_12933);
xnor U14656 (N_14656,N_12458,N_12993);
and U14657 (N_14657,N_12105,N_12196);
xnor U14658 (N_14658,N_13329,N_13246);
nor U14659 (N_14659,N_12774,N_12975);
or U14660 (N_14660,N_13557,N_13014);
or U14661 (N_14661,N_13608,N_12949);
and U14662 (N_14662,N_12970,N_13673);
or U14663 (N_14663,N_12833,N_13399);
nor U14664 (N_14664,N_13616,N_12164);
nand U14665 (N_14665,N_12950,N_13259);
and U14666 (N_14666,N_13054,N_13279);
nand U14667 (N_14667,N_13556,N_13269);
xor U14668 (N_14668,N_13363,N_12288);
nor U14669 (N_14669,N_13729,N_12052);
and U14670 (N_14670,N_13468,N_13466);
nor U14671 (N_14671,N_12584,N_12352);
or U14672 (N_14672,N_12013,N_13668);
nand U14673 (N_14673,N_13334,N_12414);
nor U14674 (N_14674,N_13001,N_13721);
nor U14675 (N_14675,N_12789,N_12811);
nand U14676 (N_14676,N_13479,N_13321);
and U14677 (N_14677,N_12566,N_12769);
xnor U14678 (N_14678,N_12531,N_12027);
nand U14679 (N_14679,N_12943,N_13941);
or U14680 (N_14680,N_12860,N_12734);
xnor U14681 (N_14681,N_13571,N_12263);
xnor U14682 (N_14682,N_13813,N_12146);
or U14683 (N_14683,N_12186,N_12509);
or U14684 (N_14684,N_12346,N_12938);
or U14685 (N_14685,N_12896,N_12675);
nand U14686 (N_14686,N_12712,N_12278);
xor U14687 (N_14687,N_12958,N_12003);
and U14688 (N_14688,N_13206,N_13789);
nand U14689 (N_14689,N_12629,N_13499);
and U14690 (N_14690,N_13076,N_13412);
or U14691 (N_14691,N_12955,N_12494);
nand U14692 (N_14692,N_12627,N_12480);
or U14693 (N_14693,N_13069,N_13908);
nand U14694 (N_14694,N_12369,N_12251);
and U14695 (N_14695,N_13563,N_12191);
nand U14696 (N_14696,N_12851,N_12632);
nand U14697 (N_14697,N_13568,N_12444);
nor U14698 (N_14698,N_12941,N_13627);
nor U14699 (N_14699,N_13738,N_12508);
xor U14700 (N_14700,N_12102,N_12026);
nor U14701 (N_14701,N_13606,N_12385);
xor U14702 (N_14702,N_12918,N_12394);
or U14703 (N_14703,N_13413,N_13583);
xnor U14704 (N_14704,N_12284,N_12390);
nand U14705 (N_14705,N_13782,N_12453);
nor U14706 (N_14706,N_13586,N_12185);
and U14707 (N_14707,N_12523,N_12100);
or U14708 (N_14708,N_13484,N_13387);
nor U14709 (N_14709,N_13359,N_13865);
xor U14710 (N_14710,N_12621,N_13938);
xor U14711 (N_14711,N_13956,N_12864);
and U14712 (N_14712,N_12561,N_13435);
xnor U14713 (N_14713,N_13093,N_13566);
nor U14714 (N_14714,N_13671,N_12942);
xnor U14715 (N_14715,N_13907,N_13748);
nand U14716 (N_14716,N_12965,N_13270);
nand U14717 (N_14717,N_13126,N_12015);
or U14718 (N_14718,N_13502,N_12801);
and U14719 (N_14719,N_13858,N_12519);
nand U14720 (N_14720,N_12902,N_13978);
xor U14721 (N_14721,N_12200,N_12211);
or U14722 (N_14722,N_13301,N_13022);
nand U14723 (N_14723,N_13980,N_12479);
xor U14724 (N_14724,N_13221,N_12567);
or U14725 (N_14725,N_12469,N_12005);
nand U14726 (N_14726,N_13923,N_12691);
xor U14727 (N_14727,N_12700,N_13860);
nor U14728 (N_14728,N_13693,N_12590);
nor U14729 (N_14729,N_13684,N_13545);
nand U14730 (N_14730,N_12841,N_12719);
xor U14731 (N_14731,N_12823,N_13648);
or U14732 (N_14732,N_12294,N_12418);
nand U14733 (N_14733,N_12517,N_12417);
nor U14734 (N_14734,N_12541,N_13681);
or U14735 (N_14735,N_13082,N_12701);
or U14736 (N_14736,N_12797,N_12597);
nor U14737 (N_14737,N_13028,N_13685);
xor U14738 (N_14738,N_13916,N_12496);
and U14739 (N_14739,N_12017,N_13451);
nand U14740 (N_14740,N_13224,N_12228);
nor U14741 (N_14741,N_13261,N_12327);
and U14742 (N_14742,N_12229,N_13176);
nand U14743 (N_14743,N_13195,N_13389);
xor U14744 (N_14744,N_12148,N_13091);
or U14745 (N_14745,N_12869,N_13217);
nor U14746 (N_14746,N_12972,N_12055);
or U14747 (N_14747,N_13423,N_12081);
xor U14748 (N_14748,N_12182,N_12914);
xnor U14749 (N_14749,N_13191,N_12507);
xor U14750 (N_14750,N_13582,N_12322);
nand U14751 (N_14751,N_12513,N_12880);
nor U14752 (N_14752,N_12495,N_13651);
xor U14753 (N_14753,N_12799,N_13534);
or U14754 (N_14754,N_12482,N_12224);
xor U14755 (N_14755,N_13249,N_13046);
and U14756 (N_14756,N_12233,N_13252);
and U14757 (N_14757,N_12877,N_12209);
xor U14758 (N_14758,N_13927,N_13314);
nand U14759 (N_14759,N_12881,N_12187);
xor U14760 (N_14760,N_13580,N_12028);
or U14761 (N_14761,N_12551,N_12430);
nor U14762 (N_14762,N_12530,N_13438);
or U14763 (N_14763,N_12408,N_13532);
nor U14764 (N_14764,N_13768,N_13553);
nand U14765 (N_14765,N_13891,N_12589);
nand U14766 (N_14766,N_13531,N_13876);
nand U14767 (N_14767,N_13186,N_13244);
nand U14768 (N_14768,N_12731,N_13900);
xnor U14769 (N_14769,N_12663,N_12865);
nor U14770 (N_14770,N_12776,N_12549);
nor U14771 (N_14771,N_13635,N_12812);
and U14772 (N_14772,N_13102,N_13669);
nor U14773 (N_14773,N_13939,N_12293);
nand U14774 (N_14774,N_12583,N_13777);
xor U14775 (N_14775,N_13886,N_13849);
or U14776 (N_14776,N_13766,N_13228);
nand U14777 (N_14777,N_12470,N_12231);
nor U14778 (N_14778,N_13226,N_12699);
xor U14779 (N_14779,N_13524,N_12935);
and U14780 (N_14780,N_13008,N_12758);
xnor U14781 (N_14781,N_13077,N_13588);
xor U14782 (N_14782,N_13472,N_13286);
and U14783 (N_14783,N_12354,N_13392);
and U14784 (N_14784,N_12063,N_12031);
or U14785 (N_14785,N_13736,N_12269);
nor U14786 (N_14786,N_12603,N_13831);
and U14787 (N_14787,N_12924,N_13150);
and U14788 (N_14788,N_12637,N_12602);
xnor U14789 (N_14789,N_12886,N_12907);
xor U14790 (N_14790,N_13624,N_13432);
nor U14791 (N_14791,N_12847,N_12953);
xor U14792 (N_14792,N_12370,N_13241);
or U14793 (N_14793,N_12285,N_12900);
xor U14794 (N_14794,N_12030,N_12276);
or U14795 (N_14795,N_13010,N_13631);
nor U14796 (N_14796,N_12533,N_12070);
nor U14797 (N_14797,N_13976,N_13265);
or U14798 (N_14798,N_13078,N_13691);
xnor U14799 (N_14799,N_12388,N_13857);
nor U14800 (N_14800,N_13665,N_12619);
nor U14801 (N_14801,N_12076,N_12272);
and U14802 (N_14802,N_12624,N_12415);
nand U14803 (N_14803,N_12245,N_12578);
xor U14804 (N_14804,N_12261,N_12406);
xnor U14805 (N_14805,N_12024,N_12867);
or U14806 (N_14806,N_13303,N_13136);
nor U14807 (N_14807,N_12904,N_12197);
and U14808 (N_14808,N_12023,N_12349);
nand U14809 (N_14809,N_12563,N_13289);
nand U14810 (N_14810,N_13390,N_12169);
or U14811 (N_14811,N_12419,N_12981);
xor U14812 (N_14812,N_12155,N_12373);
or U14813 (N_14813,N_13827,N_12041);
or U14814 (N_14814,N_13909,N_13634);
xnor U14815 (N_14815,N_13192,N_12214);
or U14816 (N_14816,N_13505,N_12543);
and U14817 (N_14817,N_12124,N_12098);
nand U14818 (N_14818,N_13822,N_12553);
or U14819 (N_14819,N_12202,N_13231);
xor U14820 (N_14820,N_13716,N_13041);
xnor U14821 (N_14821,N_12356,N_12593);
and U14822 (N_14822,N_13808,N_13799);
nand U14823 (N_14823,N_12382,N_13343);
and U14824 (N_14824,N_12931,N_13328);
and U14825 (N_14825,N_13846,N_13602);
and U14826 (N_14826,N_12757,N_12457);
and U14827 (N_14827,N_13542,N_13326);
or U14828 (N_14828,N_13278,N_12068);
and U14829 (N_14829,N_12722,N_13601);
or U14830 (N_14830,N_12868,N_13305);
or U14831 (N_14831,N_13307,N_13715);
nand U14832 (N_14832,N_12755,N_13173);
xor U14833 (N_14833,N_12744,N_12778);
nand U14834 (N_14834,N_12111,N_12655);
nor U14835 (N_14835,N_13032,N_13477);
and U14836 (N_14836,N_13406,N_13949);
nor U14837 (N_14837,N_13806,N_12213);
xor U14838 (N_14838,N_12620,N_12779);
xor U14839 (N_14839,N_13678,N_13299);
nor U14840 (N_14840,N_13928,N_12653);
nand U14841 (N_14841,N_12771,N_12180);
and U14842 (N_14842,N_12934,N_12032);
nand U14843 (N_14843,N_13480,N_13964);
or U14844 (N_14844,N_12223,N_12246);
or U14845 (N_14845,N_12204,N_13832);
nor U14846 (N_14846,N_13105,N_12332);
nand U14847 (N_14847,N_13236,N_12212);
nand U14848 (N_14848,N_13873,N_13139);
xor U14849 (N_14849,N_13755,N_13692);
nor U14850 (N_14850,N_12150,N_13199);
or U14851 (N_14851,N_13552,N_12122);
nand U14852 (N_14852,N_13323,N_12608);
nor U14853 (N_14853,N_13202,N_13788);
or U14854 (N_14854,N_13127,N_13073);
xnor U14855 (N_14855,N_12311,N_12339);
xor U14856 (N_14856,N_13169,N_13549);
nor U14857 (N_14857,N_13131,N_13374);
xor U14858 (N_14858,N_13447,N_13295);
nor U14859 (N_14859,N_12409,N_13929);
xnor U14860 (N_14860,N_12422,N_12679);
and U14861 (N_14861,N_13309,N_13835);
or U14862 (N_14862,N_12814,N_12872);
and U14863 (N_14863,N_13919,N_12625);
nand U14864 (N_14864,N_12610,N_12188);
nand U14865 (N_14865,N_13357,N_13760);
nor U14866 (N_14866,N_13605,N_12215);
nand U14867 (N_14867,N_12089,N_13332);
nand U14868 (N_14868,N_13895,N_12984);
or U14869 (N_14869,N_13285,N_13622);
nor U14870 (N_14870,N_12911,N_12093);
nor U14871 (N_14871,N_13971,N_12816);
or U14872 (N_14872,N_12694,N_12314);
and U14873 (N_14873,N_12090,N_12342);
nor U14874 (N_14874,N_13385,N_13796);
nand U14875 (N_14875,N_13463,N_12130);
xnor U14876 (N_14876,N_12290,N_13088);
and U14877 (N_14877,N_13341,N_12992);
and U14878 (N_14878,N_12813,N_12906);
nand U14879 (N_14879,N_13530,N_13005);
or U14880 (N_14880,N_12238,N_12309);
nand U14881 (N_14881,N_12947,N_12485);
or U14882 (N_14882,N_12300,N_13905);
or U14883 (N_14883,N_12681,N_13140);
and U14884 (N_14884,N_13442,N_13336);
nor U14885 (N_14885,N_12923,N_12178);
nand U14886 (N_14886,N_12324,N_12782);
and U14887 (N_14887,N_12570,N_13815);
and U14888 (N_14888,N_13512,N_12838);
xnor U14889 (N_14889,N_12748,N_13020);
and U14890 (N_14890,N_12846,N_13006);
xor U14891 (N_14891,N_12554,N_12848);
nand U14892 (N_14892,N_12666,N_13133);
nand U14893 (N_14893,N_13373,N_13870);
nand U14894 (N_14894,N_12080,N_12114);
and U14895 (N_14895,N_13042,N_12849);
or U14896 (N_14896,N_12505,N_13728);
and U14897 (N_14897,N_13458,N_12558);
or U14898 (N_14898,N_13175,N_13408);
nand U14899 (N_14899,N_13889,N_13157);
nand U14900 (N_14900,N_12084,N_12669);
nor U14901 (N_14901,N_13585,N_12650);
and U14902 (N_14902,N_12726,N_13977);
or U14903 (N_14903,N_13320,N_13371);
nand U14904 (N_14904,N_12559,N_12538);
xnor U14905 (N_14905,N_13924,N_13050);
nand U14906 (N_14906,N_13107,N_13887);
nand U14907 (N_14907,N_12139,N_13529);
nor U14908 (N_14908,N_12988,N_13380);
nor U14909 (N_14909,N_13829,N_12296);
xor U14910 (N_14910,N_13871,N_12819);
nor U14911 (N_14911,N_12662,N_12528);
xor U14912 (N_14912,N_12304,N_13074);
and U14913 (N_14913,N_13038,N_13882);
and U14914 (N_14914,N_13880,N_13707);
xnor U14915 (N_14915,N_12412,N_12464);
nor U14916 (N_14916,N_12029,N_13621);
nand U14917 (N_14917,N_12465,N_13794);
and U14918 (N_14918,N_13147,N_12488);
and U14919 (N_14919,N_13520,N_12844);
and U14920 (N_14920,N_13481,N_13434);
and U14921 (N_14921,N_12144,N_13263);
nor U14922 (N_14922,N_12172,N_13764);
nand U14923 (N_14923,N_12636,N_12129);
or U14924 (N_14924,N_13942,N_12423);
nand U14925 (N_14925,N_13004,N_12260);
or U14926 (N_14926,N_12192,N_13418);
nor U14927 (N_14927,N_12840,N_13958);
nor U14928 (N_14928,N_12009,N_12000);
nand U14929 (N_14929,N_12421,N_12301);
nand U14930 (N_14930,N_13200,N_13787);
and U14931 (N_14931,N_12809,N_13098);
xor U14932 (N_14932,N_13645,N_13572);
or U14933 (N_14933,N_13271,N_13931);
xnor U14934 (N_14934,N_12432,N_12817);
and U14935 (N_14935,N_12915,N_13065);
or U14936 (N_14936,N_12092,N_13730);
nor U14937 (N_14937,N_12428,N_13936);
or U14938 (N_14938,N_13391,N_12818);
nand U14939 (N_14939,N_13995,N_12870);
and U14940 (N_14940,N_13702,N_12378);
nand U14941 (N_14941,N_12658,N_13398);
xor U14942 (N_14942,N_12312,N_13180);
nand U14943 (N_14943,N_12253,N_13123);
nand U14944 (N_14944,N_12536,N_12117);
nand U14945 (N_14945,N_12392,N_13474);
xor U14946 (N_14946,N_12220,N_13625);
nor U14947 (N_14947,N_13629,N_12466);
nand U14948 (N_14948,N_12113,N_13896);
nor U14949 (N_14949,N_12667,N_12128);
nand U14950 (N_14950,N_13121,N_13968);
xor U14951 (N_14951,N_12104,N_12802);
nor U14952 (N_14952,N_12664,N_12564);
or U14953 (N_14953,N_12125,N_13747);
nor U14954 (N_14954,N_13780,N_13632);
xor U14955 (N_14955,N_12101,N_13302);
xnor U14956 (N_14956,N_12575,N_12962);
or U14957 (N_14957,N_13137,N_12539);
and U14958 (N_14958,N_13324,N_13277);
nor U14959 (N_14959,N_12960,N_12441);
nand U14960 (N_14960,N_13888,N_13266);
nand U14961 (N_14961,N_13155,N_13449);
nor U14962 (N_14962,N_12784,N_12752);
nand U14963 (N_14963,N_12123,N_13713);
or U14964 (N_14964,N_13955,N_12316);
xor U14965 (N_14965,N_13335,N_13443);
nand U14966 (N_14966,N_12141,N_12165);
or U14967 (N_14967,N_12500,N_12702);
nand U14968 (N_14968,N_12021,N_13372);
nor U14969 (N_14969,N_12961,N_13331);
nor U14970 (N_14970,N_12047,N_13475);
or U14971 (N_14971,N_13177,N_13649);
nor U14972 (N_14972,N_13982,N_13658);
nand U14973 (N_14973,N_13904,N_13975);
or U14974 (N_14974,N_13170,N_12247);
and U14975 (N_14975,N_13405,N_13986);
xor U14976 (N_14976,N_12732,N_12362);
or U14977 (N_14977,N_13791,N_12181);
or U14978 (N_14978,N_12723,N_13548);
xnor U14979 (N_14979,N_13201,N_12038);
or U14980 (N_14980,N_13325,N_13473);
nand U14981 (N_14981,N_12756,N_12420);
and U14982 (N_14982,N_12946,N_12836);
nand U14983 (N_14983,N_13953,N_13430);
nor U14984 (N_14984,N_12635,N_12154);
or U14985 (N_14985,N_12989,N_12025);
and U14986 (N_14986,N_12889,N_13652);
or U14987 (N_14987,N_13771,N_13537);
xor U14988 (N_14988,N_12328,N_13058);
nand U14989 (N_14989,N_12728,N_13478);
xor U14990 (N_14990,N_12376,N_12074);
or U14991 (N_14991,N_13717,N_13522);
and U14992 (N_14992,N_13560,N_12206);
xor U14993 (N_14993,N_13724,N_12545);
xor U14994 (N_14994,N_13376,N_12521);
xor U14995 (N_14995,N_13866,N_13599);
or U14996 (N_14996,N_13753,N_12928);
and U14997 (N_14997,N_12897,N_12413);
nand U14998 (N_14998,N_12630,N_13344);
nand U14999 (N_14999,N_12534,N_12668);
or U15000 (N_15000,N_13818,N_12509);
nand U15001 (N_15001,N_12155,N_13201);
or U15002 (N_15002,N_12098,N_13573);
nand U15003 (N_15003,N_13479,N_12072);
xnor U15004 (N_15004,N_13666,N_13282);
nor U15005 (N_15005,N_12970,N_12206);
or U15006 (N_15006,N_13429,N_13445);
xnor U15007 (N_15007,N_13153,N_13499);
nand U15008 (N_15008,N_12963,N_12175);
nor U15009 (N_15009,N_12463,N_12911);
or U15010 (N_15010,N_12574,N_13387);
or U15011 (N_15011,N_12693,N_13820);
nand U15012 (N_15012,N_12237,N_13378);
nor U15013 (N_15013,N_12504,N_12492);
or U15014 (N_15014,N_13082,N_13467);
or U15015 (N_15015,N_12298,N_13120);
and U15016 (N_15016,N_13308,N_13616);
nor U15017 (N_15017,N_13651,N_12534);
or U15018 (N_15018,N_12220,N_12241);
and U15019 (N_15019,N_13702,N_13201);
xor U15020 (N_15020,N_13347,N_12381);
xnor U15021 (N_15021,N_13453,N_13870);
or U15022 (N_15022,N_13466,N_12469);
xnor U15023 (N_15023,N_13916,N_13328);
or U15024 (N_15024,N_12986,N_13096);
xor U15025 (N_15025,N_13932,N_13428);
nand U15026 (N_15026,N_13673,N_12939);
nand U15027 (N_15027,N_12384,N_12140);
nand U15028 (N_15028,N_12137,N_13075);
or U15029 (N_15029,N_13019,N_12165);
nand U15030 (N_15030,N_12686,N_12842);
nand U15031 (N_15031,N_13338,N_13005);
xnor U15032 (N_15032,N_12462,N_12195);
nor U15033 (N_15033,N_13523,N_12530);
nor U15034 (N_15034,N_12382,N_12965);
and U15035 (N_15035,N_13630,N_13452);
xnor U15036 (N_15036,N_13610,N_12442);
nand U15037 (N_15037,N_13645,N_13737);
and U15038 (N_15038,N_13593,N_13739);
nand U15039 (N_15039,N_12682,N_12831);
or U15040 (N_15040,N_13483,N_12696);
xor U15041 (N_15041,N_13845,N_13024);
nor U15042 (N_15042,N_12778,N_13857);
nor U15043 (N_15043,N_13348,N_13578);
xor U15044 (N_15044,N_12768,N_12487);
or U15045 (N_15045,N_12037,N_12465);
xnor U15046 (N_15046,N_13308,N_12333);
or U15047 (N_15047,N_12176,N_12606);
nor U15048 (N_15048,N_13290,N_13531);
nand U15049 (N_15049,N_13492,N_13418);
nand U15050 (N_15050,N_12646,N_12028);
nor U15051 (N_15051,N_13264,N_12485);
nor U15052 (N_15052,N_13215,N_13749);
or U15053 (N_15053,N_12271,N_12301);
nor U15054 (N_15054,N_12149,N_12677);
xor U15055 (N_15055,N_12911,N_12204);
xor U15056 (N_15056,N_12496,N_12683);
nand U15057 (N_15057,N_13918,N_12911);
and U15058 (N_15058,N_13986,N_13657);
or U15059 (N_15059,N_13939,N_12656);
and U15060 (N_15060,N_13456,N_13621);
and U15061 (N_15061,N_12831,N_12865);
nor U15062 (N_15062,N_12096,N_12743);
nand U15063 (N_15063,N_13124,N_13108);
xor U15064 (N_15064,N_12110,N_12259);
and U15065 (N_15065,N_12476,N_12818);
nand U15066 (N_15066,N_13342,N_13242);
nand U15067 (N_15067,N_12377,N_13951);
xor U15068 (N_15068,N_12895,N_12096);
or U15069 (N_15069,N_12159,N_13327);
nor U15070 (N_15070,N_13030,N_13316);
xor U15071 (N_15071,N_13132,N_13617);
and U15072 (N_15072,N_13661,N_12361);
and U15073 (N_15073,N_13577,N_12480);
xnor U15074 (N_15074,N_12766,N_12628);
and U15075 (N_15075,N_13443,N_12398);
and U15076 (N_15076,N_13109,N_12116);
nand U15077 (N_15077,N_12870,N_13301);
nor U15078 (N_15078,N_13195,N_13556);
or U15079 (N_15079,N_12349,N_13311);
nand U15080 (N_15080,N_13564,N_13088);
nand U15081 (N_15081,N_13704,N_12171);
or U15082 (N_15082,N_13450,N_13163);
nand U15083 (N_15083,N_13984,N_13199);
or U15084 (N_15084,N_13524,N_13390);
and U15085 (N_15085,N_13620,N_13480);
and U15086 (N_15086,N_12029,N_13074);
and U15087 (N_15087,N_12024,N_12144);
xor U15088 (N_15088,N_13825,N_13210);
and U15089 (N_15089,N_13184,N_12932);
nand U15090 (N_15090,N_12859,N_12797);
and U15091 (N_15091,N_12045,N_13617);
and U15092 (N_15092,N_12467,N_13702);
nand U15093 (N_15093,N_13244,N_13440);
nor U15094 (N_15094,N_12765,N_13728);
nor U15095 (N_15095,N_12390,N_12517);
and U15096 (N_15096,N_13673,N_13983);
nand U15097 (N_15097,N_12290,N_12864);
or U15098 (N_15098,N_13172,N_12651);
nor U15099 (N_15099,N_13662,N_12532);
and U15100 (N_15100,N_13429,N_13565);
nor U15101 (N_15101,N_13020,N_12438);
nand U15102 (N_15102,N_13270,N_12298);
or U15103 (N_15103,N_13140,N_12989);
and U15104 (N_15104,N_12633,N_12177);
nor U15105 (N_15105,N_13635,N_13998);
or U15106 (N_15106,N_13797,N_12225);
nor U15107 (N_15107,N_12133,N_12466);
nand U15108 (N_15108,N_13234,N_12119);
or U15109 (N_15109,N_12448,N_13061);
nand U15110 (N_15110,N_13108,N_13457);
nand U15111 (N_15111,N_12346,N_12323);
nand U15112 (N_15112,N_13438,N_13701);
nor U15113 (N_15113,N_12818,N_12541);
xnor U15114 (N_15114,N_13633,N_12811);
xor U15115 (N_15115,N_12003,N_13046);
nor U15116 (N_15116,N_12576,N_12156);
and U15117 (N_15117,N_12672,N_12160);
or U15118 (N_15118,N_13468,N_13387);
nand U15119 (N_15119,N_12534,N_13326);
nor U15120 (N_15120,N_13095,N_13979);
nor U15121 (N_15121,N_13040,N_13379);
nor U15122 (N_15122,N_13492,N_13244);
nand U15123 (N_15123,N_12298,N_12708);
nand U15124 (N_15124,N_13064,N_12092);
or U15125 (N_15125,N_13020,N_13487);
nand U15126 (N_15126,N_12936,N_12071);
and U15127 (N_15127,N_13668,N_12387);
nor U15128 (N_15128,N_12533,N_12314);
nand U15129 (N_15129,N_13756,N_13443);
and U15130 (N_15130,N_12231,N_13816);
nand U15131 (N_15131,N_12771,N_13410);
xor U15132 (N_15132,N_12374,N_12668);
nand U15133 (N_15133,N_12970,N_12405);
nor U15134 (N_15134,N_13909,N_12243);
xnor U15135 (N_15135,N_12150,N_12830);
nand U15136 (N_15136,N_13284,N_12319);
nand U15137 (N_15137,N_13895,N_12242);
nor U15138 (N_15138,N_13635,N_13652);
nor U15139 (N_15139,N_12864,N_13808);
xnor U15140 (N_15140,N_13378,N_13225);
or U15141 (N_15141,N_13410,N_12413);
xor U15142 (N_15142,N_13477,N_13570);
and U15143 (N_15143,N_12965,N_12509);
nor U15144 (N_15144,N_12173,N_13376);
xnor U15145 (N_15145,N_12443,N_13579);
or U15146 (N_15146,N_13259,N_13198);
nor U15147 (N_15147,N_12166,N_13731);
xnor U15148 (N_15148,N_12605,N_12292);
nor U15149 (N_15149,N_12923,N_12755);
and U15150 (N_15150,N_13907,N_13426);
xor U15151 (N_15151,N_13772,N_12878);
and U15152 (N_15152,N_12588,N_13671);
nor U15153 (N_15153,N_12786,N_13374);
nand U15154 (N_15154,N_12050,N_13691);
or U15155 (N_15155,N_13588,N_12658);
and U15156 (N_15156,N_12567,N_12442);
or U15157 (N_15157,N_12577,N_13465);
or U15158 (N_15158,N_12761,N_13757);
nand U15159 (N_15159,N_13221,N_12176);
xor U15160 (N_15160,N_12645,N_13838);
and U15161 (N_15161,N_13107,N_12147);
nand U15162 (N_15162,N_12862,N_12984);
or U15163 (N_15163,N_13118,N_12655);
nor U15164 (N_15164,N_13245,N_12534);
xor U15165 (N_15165,N_13931,N_13270);
xnor U15166 (N_15166,N_12793,N_13789);
nor U15167 (N_15167,N_12325,N_13421);
and U15168 (N_15168,N_13862,N_13100);
or U15169 (N_15169,N_12215,N_13069);
or U15170 (N_15170,N_13222,N_12217);
nand U15171 (N_15171,N_13830,N_12035);
nor U15172 (N_15172,N_13652,N_13333);
nand U15173 (N_15173,N_12818,N_12068);
nand U15174 (N_15174,N_13313,N_13260);
and U15175 (N_15175,N_12742,N_13600);
or U15176 (N_15176,N_12137,N_13630);
xnor U15177 (N_15177,N_12636,N_12761);
or U15178 (N_15178,N_13889,N_13607);
nand U15179 (N_15179,N_13352,N_12778);
nor U15180 (N_15180,N_13296,N_12974);
nand U15181 (N_15181,N_12223,N_12317);
xor U15182 (N_15182,N_13322,N_12907);
xor U15183 (N_15183,N_13392,N_12477);
xor U15184 (N_15184,N_12083,N_12280);
and U15185 (N_15185,N_12661,N_13018);
nand U15186 (N_15186,N_13582,N_12081);
or U15187 (N_15187,N_13335,N_13455);
and U15188 (N_15188,N_13178,N_13616);
or U15189 (N_15189,N_12661,N_12607);
or U15190 (N_15190,N_13077,N_12303);
and U15191 (N_15191,N_12231,N_12486);
and U15192 (N_15192,N_12501,N_12869);
or U15193 (N_15193,N_13557,N_13269);
nand U15194 (N_15194,N_12961,N_13194);
nor U15195 (N_15195,N_12240,N_13137);
nand U15196 (N_15196,N_13264,N_12985);
xor U15197 (N_15197,N_13590,N_13810);
nand U15198 (N_15198,N_13012,N_13262);
or U15199 (N_15199,N_12026,N_13631);
xor U15200 (N_15200,N_13672,N_12477);
xnor U15201 (N_15201,N_13617,N_13426);
nand U15202 (N_15202,N_13599,N_12102);
and U15203 (N_15203,N_12435,N_13687);
nand U15204 (N_15204,N_12238,N_13157);
or U15205 (N_15205,N_13768,N_13709);
and U15206 (N_15206,N_13858,N_12885);
nor U15207 (N_15207,N_12859,N_13335);
nor U15208 (N_15208,N_12574,N_13722);
and U15209 (N_15209,N_12759,N_12319);
nand U15210 (N_15210,N_13080,N_13214);
or U15211 (N_15211,N_13921,N_13242);
xnor U15212 (N_15212,N_12911,N_12576);
nand U15213 (N_15213,N_13869,N_13571);
or U15214 (N_15214,N_13274,N_12378);
or U15215 (N_15215,N_13828,N_12375);
xor U15216 (N_15216,N_13278,N_13517);
nand U15217 (N_15217,N_13840,N_13034);
and U15218 (N_15218,N_13353,N_13003);
nand U15219 (N_15219,N_13020,N_12424);
nor U15220 (N_15220,N_12316,N_12590);
or U15221 (N_15221,N_13948,N_12349);
or U15222 (N_15222,N_12161,N_12519);
nor U15223 (N_15223,N_12986,N_13221);
nand U15224 (N_15224,N_13297,N_13703);
or U15225 (N_15225,N_12354,N_13207);
and U15226 (N_15226,N_13270,N_12339);
xnor U15227 (N_15227,N_13940,N_13128);
xnor U15228 (N_15228,N_12822,N_12940);
or U15229 (N_15229,N_12666,N_13930);
nor U15230 (N_15230,N_12287,N_13956);
xor U15231 (N_15231,N_13307,N_13957);
nand U15232 (N_15232,N_12024,N_12775);
xor U15233 (N_15233,N_13912,N_13991);
nand U15234 (N_15234,N_13750,N_12905);
nor U15235 (N_15235,N_13206,N_12139);
xnor U15236 (N_15236,N_12703,N_12936);
or U15237 (N_15237,N_12063,N_13741);
nand U15238 (N_15238,N_12785,N_12014);
nor U15239 (N_15239,N_13146,N_12444);
nor U15240 (N_15240,N_13920,N_13722);
and U15241 (N_15241,N_13327,N_12248);
or U15242 (N_15242,N_12380,N_12314);
nor U15243 (N_15243,N_12373,N_12158);
or U15244 (N_15244,N_13966,N_13729);
xnor U15245 (N_15245,N_13457,N_13347);
nand U15246 (N_15246,N_12324,N_13813);
and U15247 (N_15247,N_13769,N_12901);
nand U15248 (N_15248,N_13400,N_12661);
and U15249 (N_15249,N_12876,N_12803);
and U15250 (N_15250,N_12176,N_13238);
and U15251 (N_15251,N_13641,N_12147);
nand U15252 (N_15252,N_13016,N_13352);
nor U15253 (N_15253,N_13604,N_12051);
nand U15254 (N_15254,N_12831,N_13850);
or U15255 (N_15255,N_12729,N_13173);
nor U15256 (N_15256,N_13108,N_12977);
xnor U15257 (N_15257,N_13039,N_13839);
or U15258 (N_15258,N_13995,N_13674);
nand U15259 (N_15259,N_13953,N_12338);
xnor U15260 (N_15260,N_12911,N_12887);
xor U15261 (N_15261,N_13783,N_13748);
or U15262 (N_15262,N_13434,N_12638);
nand U15263 (N_15263,N_12039,N_12264);
xor U15264 (N_15264,N_12012,N_13028);
xor U15265 (N_15265,N_13102,N_13653);
and U15266 (N_15266,N_13988,N_12399);
and U15267 (N_15267,N_13749,N_12528);
nor U15268 (N_15268,N_13162,N_13161);
nor U15269 (N_15269,N_13450,N_13112);
nor U15270 (N_15270,N_12218,N_13128);
nand U15271 (N_15271,N_13606,N_13799);
xor U15272 (N_15272,N_12832,N_12917);
nor U15273 (N_15273,N_12126,N_13628);
nand U15274 (N_15274,N_13554,N_12835);
and U15275 (N_15275,N_13376,N_12071);
nor U15276 (N_15276,N_12212,N_12485);
nand U15277 (N_15277,N_13531,N_13945);
and U15278 (N_15278,N_12779,N_12854);
or U15279 (N_15279,N_12211,N_12014);
xor U15280 (N_15280,N_13170,N_12404);
or U15281 (N_15281,N_13953,N_13169);
nand U15282 (N_15282,N_13565,N_12730);
and U15283 (N_15283,N_12174,N_12352);
xor U15284 (N_15284,N_13267,N_13165);
and U15285 (N_15285,N_12986,N_12913);
xor U15286 (N_15286,N_12020,N_12774);
nand U15287 (N_15287,N_12941,N_13073);
xnor U15288 (N_15288,N_13053,N_12271);
or U15289 (N_15289,N_12589,N_12904);
nor U15290 (N_15290,N_13802,N_13227);
xnor U15291 (N_15291,N_12877,N_13491);
or U15292 (N_15292,N_13272,N_13073);
and U15293 (N_15293,N_12784,N_13276);
xnor U15294 (N_15294,N_12138,N_12307);
nor U15295 (N_15295,N_12340,N_12358);
nor U15296 (N_15296,N_12041,N_13460);
xor U15297 (N_15297,N_13883,N_13283);
and U15298 (N_15298,N_13123,N_13809);
nor U15299 (N_15299,N_13844,N_12301);
or U15300 (N_15300,N_12988,N_13096);
or U15301 (N_15301,N_13876,N_12880);
nand U15302 (N_15302,N_13515,N_12753);
or U15303 (N_15303,N_13276,N_12058);
or U15304 (N_15304,N_13072,N_13223);
nor U15305 (N_15305,N_13437,N_12800);
nand U15306 (N_15306,N_12142,N_12961);
nand U15307 (N_15307,N_13018,N_13867);
xor U15308 (N_15308,N_13093,N_12607);
and U15309 (N_15309,N_12823,N_12648);
nor U15310 (N_15310,N_12843,N_12479);
xnor U15311 (N_15311,N_13859,N_12762);
nand U15312 (N_15312,N_12909,N_12354);
xnor U15313 (N_15313,N_13471,N_12032);
and U15314 (N_15314,N_13416,N_12217);
or U15315 (N_15315,N_12189,N_12151);
nand U15316 (N_15316,N_12689,N_13997);
nor U15317 (N_15317,N_13582,N_12803);
nand U15318 (N_15318,N_13304,N_12705);
or U15319 (N_15319,N_12893,N_13128);
or U15320 (N_15320,N_13960,N_12584);
xnor U15321 (N_15321,N_12017,N_13546);
nor U15322 (N_15322,N_13107,N_12452);
and U15323 (N_15323,N_13498,N_12113);
and U15324 (N_15324,N_12378,N_12080);
nand U15325 (N_15325,N_13000,N_13388);
or U15326 (N_15326,N_12385,N_12748);
and U15327 (N_15327,N_12691,N_13049);
xor U15328 (N_15328,N_13308,N_13668);
nand U15329 (N_15329,N_13298,N_12662);
or U15330 (N_15330,N_13357,N_13088);
and U15331 (N_15331,N_12963,N_13750);
or U15332 (N_15332,N_12695,N_12511);
xor U15333 (N_15333,N_12857,N_12715);
xor U15334 (N_15334,N_13992,N_13702);
nand U15335 (N_15335,N_12399,N_13552);
and U15336 (N_15336,N_12427,N_13561);
nand U15337 (N_15337,N_12927,N_13266);
xnor U15338 (N_15338,N_12307,N_13133);
or U15339 (N_15339,N_12395,N_12002);
xor U15340 (N_15340,N_12464,N_12786);
and U15341 (N_15341,N_12255,N_13590);
xnor U15342 (N_15342,N_12892,N_13423);
xor U15343 (N_15343,N_12744,N_12289);
and U15344 (N_15344,N_12778,N_13938);
nand U15345 (N_15345,N_12192,N_12440);
nand U15346 (N_15346,N_12454,N_12613);
xnor U15347 (N_15347,N_12625,N_13659);
or U15348 (N_15348,N_13930,N_12255);
nand U15349 (N_15349,N_13714,N_13619);
or U15350 (N_15350,N_12861,N_12474);
or U15351 (N_15351,N_13912,N_12431);
nor U15352 (N_15352,N_13960,N_13456);
and U15353 (N_15353,N_12800,N_13930);
nand U15354 (N_15354,N_12021,N_12062);
nand U15355 (N_15355,N_12568,N_13611);
nor U15356 (N_15356,N_13254,N_13878);
nor U15357 (N_15357,N_13924,N_13696);
or U15358 (N_15358,N_13251,N_13953);
nor U15359 (N_15359,N_13694,N_13262);
xor U15360 (N_15360,N_13066,N_12200);
nand U15361 (N_15361,N_12072,N_12024);
nor U15362 (N_15362,N_12376,N_12229);
xnor U15363 (N_15363,N_12289,N_12409);
nor U15364 (N_15364,N_13410,N_13751);
or U15365 (N_15365,N_12711,N_13554);
nor U15366 (N_15366,N_12417,N_12914);
xnor U15367 (N_15367,N_12893,N_12952);
or U15368 (N_15368,N_13865,N_13246);
nand U15369 (N_15369,N_12149,N_13767);
xnor U15370 (N_15370,N_13197,N_12806);
nand U15371 (N_15371,N_13161,N_12719);
nor U15372 (N_15372,N_13406,N_13343);
and U15373 (N_15373,N_12170,N_12196);
or U15374 (N_15374,N_13890,N_13368);
nand U15375 (N_15375,N_13284,N_12437);
and U15376 (N_15376,N_12848,N_13819);
and U15377 (N_15377,N_13931,N_13155);
xor U15378 (N_15378,N_12438,N_13439);
or U15379 (N_15379,N_12179,N_13599);
nand U15380 (N_15380,N_13606,N_13481);
nor U15381 (N_15381,N_13338,N_13984);
xnor U15382 (N_15382,N_13134,N_12365);
xnor U15383 (N_15383,N_13175,N_13184);
nand U15384 (N_15384,N_13481,N_12713);
or U15385 (N_15385,N_13493,N_13939);
nor U15386 (N_15386,N_12442,N_12278);
or U15387 (N_15387,N_12654,N_13035);
and U15388 (N_15388,N_13424,N_12815);
and U15389 (N_15389,N_13337,N_13941);
xor U15390 (N_15390,N_12976,N_12316);
nor U15391 (N_15391,N_13276,N_12747);
or U15392 (N_15392,N_12291,N_13150);
or U15393 (N_15393,N_13915,N_12864);
xor U15394 (N_15394,N_13961,N_12891);
nand U15395 (N_15395,N_13660,N_13038);
nand U15396 (N_15396,N_12566,N_13076);
and U15397 (N_15397,N_12778,N_12122);
nor U15398 (N_15398,N_12383,N_13608);
nand U15399 (N_15399,N_13743,N_12485);
xor U15400 (N_15400,N_12635,N_13290);
nand U15401 (N_15401,N_13041,N_12905);
xnor U15402 (N_15402,N_12432,N_13432);
nor U15403 (N_15403,N_12598,N_13111);
or U15404 (N_15404,N_13219,N_12928);
nand U15405 (N_15405,N_13528,N_12254);
nor U15406 (N_15406,N_12137,N_13791);
nand U15407 (N_15407,N_13137,N_12520);
xor U15408 (N_15408,N_12991,N_12037);
or U15409 (N_15409,N_12232,N_12277);
nand U15410 (N_15410,N_13051,N_12851);
xnor U15411 (N_15411,N_12665,N_12762);
or U15412 (N_15412,N_12111,N_13965);
xor U15413 (N_15413,N_12265,N_13014);
nor U15414 (N_15414,N_13634,N_12202);
and U15415 (N_15415,N_13219,N_13330);
nor U15416 (N_15416,N_13068,N_12462);
xnor U15417 (N_15417,N_13005,N_13939);
xnor U15418 (N_15418,N_12174,N_13970);
or U15419 (N_15419,N_12125,N_13982);
or U15420 (N_15420,N_12972,N_12440);
xnor U15421 (N_15421,N_12642,N_13293);
and U15422 (N_15422,N_13091,N_12510);
and U15423 (N_15423,N_12628,N_12521);
xor U15424 (N_15424,N_12313,N_12189);
nand U15425 (N_15425,N_13178,N_13579);
xor U15426 (N_15426,N_12665,N_12460);
or U15427 (N_15427,N_13900,N_13475);
and U15428 (N_15428,N_12367,N_12814);
nor U15429 (N_15429,N_13798,N_12248);
nand U15430 (N_15430,N_13546,N_13615);
nor U15431 (N_15431,N_13453,N_13563);
and U15432 (N_15432,N_12998,N_13763);
xnor U15433 (N_15433,N_13013,N_13645);
nand U15434 (N_15434,N_12952,N_12867);
or U15435 (N_15435,N_12181,N_13449);
nand U15436 (N_15436,N_12648,N_13229);
nand U15437 (N_15437,N_12651,N_13410);
xnor U15438 (N_15438,N_13918,N_13037);
nand U15439 (N_15439,N_13442,N_13369);
and U15440 (N_15440,N_12767,N_13438);
and U15441 (N_15441,N_13811,N_12394);
and U15442 (N_15442,N_12158,N_13189);
xnor U15443 (N_15443,N_12227,N_13228);
nand U15444 (N_15444,N_12735,N_12272);
nor U15445 (N_15445,N_13003,N_12665);
xor U15446 (N_15446,N_13335,N_13564);
nor U15447 (N_15447,N_12739,N_13531);
nor U15448 (N_15448,N_13282,N_13389);
nand U15449 (N_15449,N_13189,N_12616);
nand U15450 (N_15450,N_13011,N_13020);
xnor U15451 (N_15451,N_12186,N_12847);
and U15452 (N_15452,N_13616,N_12514);
nand U15453 (N_15453,N_12572,N_13790);
nand U15454 (N_15454,N_12623,N_13734);
nand U15455 (N_15455,N_12611,N_12694);
or U15456 (N_15456,N_13009,N_12850);
or U15457 (N_15457,N_12645,N_12342);
nor U15458 (N_15458,N_12499,N_13432);
nor U15459 (N_15459,N_12718,N_12789);
and U15460 (N_15460,N_13357,N_12264);
xor U15461 (N_15461,N_12103,N_12689);
and U15462 (N_15462,N_12149,N_13770);
nand U15463 (N_15463,N_12920,N_13959);
nor U15464 (N_15464,N_13045,N_13280);
nand U15465 (N_15465,N_13185,N_13353);
nand U15466 (N_15466,N_13362,N_13511);
nand U15467 (N_15467,N_13300,N_13262);
xor U15468 (N_15468,N_13263,N_13738);
nor U15469 (N_15469,N_12548,N_12495);
or U15470 (N_15470,N_13163,N_12082);
nand U15471 (N_15471,N_12095,N_12594);
nand U15472 (N_15472,N_12117,N_12545);
xor U15473 (N_15473,N_13350,N_12195);
nand U15474 (N_15474,N_12455,N_13517);
xnor U15475 (N_15475,N_13691,N_13823);
or U15476 (N_15476,N_13117,N_13710);
nor U15477 (N_15477,N_12316,N_13784);
xnor U15478 (N_15478,N_12968,N_13953);
or U15479 (N_15479,N_13646,N_13800);
and U15480 (N_15480,N_13095,N_13823);
and U15481 (N_15481,N_12566,N_13762);
xor U15482 (N_15482,N_12694,N_12655);
or U15483 (N_15483,N_13985,N_12300);
nor U15484 (N_15484,N_12120,N_13086);
nor U15485 (N_15485,N_12201,N_13974);
or U15486 (N_15486,N_13901,N_12173);
and U15487 (N_15487,N_13925,N_13330);
nand U15488 (N_15488,N_12350,N_12287);
xor U15489 (N_15489,N_13197,N_12043);
or U15490 (N_15490,N_12456,N_13893);
or U15491 (N_15491,N_12985,N_12243);
nor U15492 (N_15492,N_12976,N_12177);
and U15493 (N_15493,N_12560,N_12860);
xnor U15494 (N_15494,N_12277,N_13256);
or U15495 (N_15495,N_12427,N_12096);
xnor U15496 (N_15496,N_13843,N_12469);
and U15497 (N_15497,N_13961,N_13870);
or U15498 (N_15498,N_12569,N_12299);
nor U15499 (N_15499,N_13083,N_13453);
nand U15500 (N_15500,N_13378,N_12035);
nand U15501 (N_15501,N_12471,N_12497);
xnor U15502 (N_15502,N_12409,N_13587);
or U15503 (N_15503,N_12222,N_13759);
nor U15504 (N_15504,N_13516,N_13283);
xor U15505 (N_15505,N_13657,N_12631);
or U15506 (N_15506,N_13918,N_13112);
and U15507 (N_15507,N_13368,N_13288);
or U15508 (N_15508,N_12952,N_13641);
nand U15509 (N_15509,N_12852,N_13810);
and U15510 (N_15510,N_12902,N_13876);
or U15511 (N_15511,N_13989,N_12485);
or U15512 (N_15512,N_13855,N_13717);
xor U15513 (N_15513,N_13358,N_12324);
nor U15514 (N_15514,N_13606,N_12157);
nand U15515 (N_15515,N_13609,N_13921);
or U15516 (N_15516,N_13455,N_13552);
or U15517 (N_15517,N_12030,N_12710);
or U15518 (N_15518,N_13100,N_12617);
or U15519 (N_15519,N_13301,N_13289);
and U15520 (N_15520,N_12456,N_13822);
and U15521 (N_15521,N_13035,N_13273);
xnor U15522 (N_15522,N_12516,N_13994);
nand U15523 (N_15523,N_12156,N_13736);
xor U15524 (N_15524,N_13395,N_12397);
nand U15525 (N_15525,N_13406,N_12330);
and U15526 (N_15526,N_12334,N_13071);
or U15527 (N_15527,N_12108,N_13494);
nor U15528 (N_15528,N_12795,N_13280);
nand U15529 (N_15529,N_12059,N_13013);
or U15530 (N_15530,N_13043,N_13979);
nand U15531 (N_15531,N_13078,N_12069);
nand U15532 (N_15532,N_13813,N_13759);
xor U15533 (N_15533,N_12066,N_13275);
nor U15534 (N_15534,N_12542,N_13765);
nor U15535 (N_15535,N_13634,N_12125);
nor U15536 (N_15536,N_12298,N_13299);
or U15537 (N_15537,N_12025,N_13737);
and U15538 (N_15538,N_12796,N_12061);
or U15539 (N_15539,N_13930,N_13371);
xnor U15540 (N_15540,N_13169,N_13467);
xnor U15541 (N_15541,N_13992,N_13290);
xor U15542 (N_15542,N_13220,N_13109);
or U15543 (N_15543,N_12131,N_12980);
and U15544 (N_15544,N_12282,N_12815);
nor U15545 (N_15545,N_12655,N_12903);
or U15546 (N_15546,N_12746,N_13619);
nor U15547 (N_15547,N_13195,N_13545);
xnor U15548 (N_15548,N_12222,N_13870);
xor U15549 (N_15549,N_12160,N_12780);
xor U15550 (N_15550,N_12111,N_13822);
and U15551 (N_15551,N_13052,N_12179);
nor U15552 (N_15552,N_12082,N_13270);
xor U15553 (N_15553,N_12385,N_12289);
and U15554 (N_15554,N_12070,N_12342);
xnor U15555 (N_15555,N_12264,N_12404);
nand U15556 (N_15556,N_13990,N_13926);
or U15557 (N_15557,N_12360,N_12682);
nand U15558 (N_15558,N_12604,N_13973);
nand U15559 (N_15559,N_12661,N_12270);
xor U15560 (N_15560,N_13554,N_13489);
nor U15561 (N_15561,N_12975,N_13809);
xnor U15562 (N_15562,N_12152,N_12766);
nand U15563 (N_15563,N_13638,N_13536);
or U15564 (N_15564,N_12959,N_13410);
and U15565 (N_15565,N_13579,N_12586);
nand U15566 (N_15566,N_13956,N_13951);
nor U15567 (N_15567,N_13696,N_13169);
nor U15568 (N_15568,N_13115,N_12356);
or U15569 (N_15569,N_13506,N_13847);
or U15570 (N_15570,N_13930,N_12477);
or U15571 (N_15571,N_12638,N_13424);
or U15572 (N_15572,N_13358,N_12668);
and U15573 (N_15573,N_12363,N_12532);
nand U15574 (N_15574,N_12626,N_12500);
xnor U15575 (N_15575,N_12201,N_13863);
nor U15576 (N_15576,N_12713,N_13911);
nor U15577 (N_15577,N_12144,N_12904);
nand U15578 (N_15578,N_13111,N_13897);
and U15579 (N_15579,N_13227,N_13136);
or U15580 (N_15580,N_12945,N_13798);
and U15581 (N_15581,N_13394,N_12843);
or U15582 (N_15582,N_13466,N_12679);
or U15583 (N_15583,N_12504,N_13617);
nand U15584 (N_15584,N_12370,N_13287);
and U15585 (N_15585,N_13936,N_12967);
and U15586 (N_15586,N_13807,N_13639);
xnor U15587 (N_15587,N_12735,N_13983);
or U15588 (N_15588,N_13347,N_12961);
nor U15589 (N_15589,N_13713,N_12701);
nand U15590 (N_15590,N_12024,N_13605);
nand U15591 (N_15591,N_13638,N_12721);
or U15592 (N_15592,N_13187,N_13273);
nand U15593 (N_15593,N_13176,N_12146);
and U15594 (N_15594,N_13236,N_13800);
nand U15595 (N_15595,N_13855,N_13914);
and U15596 (N_15596,N_13684,N_13069);
nor U15597 (N_15597,N_12852,N_13969);
nor U15598 (N_15598,N_13593,N_12388);
nor U15599 (N_15599,N_13485,N_13130);
xor U15600 (N_15600,N_13435,N_13415);
or U15601 (N_15601,N_12556,N_12333);
xnor U15602 (N_15602,N_13301,N_12684);
nor U15603 (N_15603,N_13267,N_13529);
nor U15604 (N_15604,N_12915,N_12395);
and U15605 (N_15605,N_12872,N_13759);
or U15606 (N_15606,N_13661,N_13233);
nand U15607 (N_15607,N_13889,N_12366);
and U15608 (N_15608,N_12705,N_12018);
xor U15609 (N_15609,N_12148,N_12096);
or U15610 (N_15610,N_13618,N_12743);
xnor U15611 (N_15611,N_13271,N_13401);
and U15612 (N_15612,N_12814,N_12941);
or U15613 (N_15613,N_13925,N_13064);
or U15614 (N_15614,N_12243,N_12904);
xnor U15615 (N_15615,N_12772,N_13869);
nor U15616 (N_15616,N_12098,N_12357);
and U15617 (N_15617,N_13637,N_13086);
and U15618 (N_15618,N_12972,N_12254);
and U15619 (N_15619,N_13561,N_13340);
and U15620 (N_15620,N_12948,N_12481);
nand U15621 (N_15621,N_13621,N_12311);
or U15622 (N_15622,N_13342,N_13880);
or U15623 (N_15623,N_12432,N_13397);
or U15624 (N_15624,N_12193,N_12857);
and U15625 (N_15625,N_13862,N_13912);
nor U15626 (N_15626,N_13327,N_12156);
nor U15627 (N_15627,N_12424,N_12562);
and U15628 (N_15628,N_12654,N_12806);
or U15629 (N_15629,N_13798,N_13726);
or U15630 (N_15630,N_13916,N_13997);
xor U15631 (N_15631,N_13404,N_13392);
or U15632 (N_15632,N_13419,N_13524);
nor U15633 (N_15633,N_12810,N_12084);
xor U15634 (N_15634,N_13411,N_13892);
xor U15635 (N_15635,N_12048,N_12269);
nand U15636 (N_15636,N_12261,N_12130);
and U15637 (N_15637,N_12196,N_12919);
xnor U15638 (N_15638,N_13871,N_13821);
nor U15639 (N_15639,N_12119,N_12355);
nor U15640 (N_15640,N_12778,N_12211);
nor U15641 (N_15641,N_12617,N_12953);
xnor U15642 (N_15642,N_13457,N_13572);
nor U15643 (N_15643,N_13100,N_12499);
xnor U15644 (N_15644,N_13831,N_13101);
or U15645 (N_15645,N_12601,N_12174);
nand U15646 (N_15646,N_12914,N_12137);
and U15647 (N_15647,N_12594,N_12855);
nor U15648 (N_15648,N_13474,N_13121);
and U15649 (N_15649,N_13776,N_13277);
xnor U15650 (N_15650,N_13935,N_12655);
or U15651 (N_15651,N_13919,N_12205);
xor U15652 (N_15652,N_13586,N_12786);
and U15653 (N_15653,N_12517,N_12806);
nor U15654 (N_15654,N_12709,N_13090);
and U15655 (N_15655,N_13504,N_12984);
xnor U15656 (N_15656,N_13930,N_13761);
and U15657 (N_15657,N_13635,N_12217);
and U15658 (N_15658,N_13418,N_13505);
nor U15659 (N_15659,N_13236,N_12304);
or U15660 (N_15660,N_12022,N_13632);
or U15661 (N_15661,N_13938,N_12231);
xnor U15662 (N_15662,N_13740,N_13278);
nor U15663 (N_15663,N_12765,N_12343);
nand U15664 (N_15664,N_12857,N_13213);
nand U15665 (N_15665,N_13254,N_13357);
or U15666 (N_15666,N_12389,N_12360);
or U15667 (N_15667,N_13929,N_12652);
or U15668 (N_15668,N_13146,N_12928);
or U15669 (N_15669,N_13813,N_13534);
or U15670 (N_15670,N_12431,N_13689);
nand U15671 (N_15671,N_13234,N_12870);
nor U15672 (N_15672,N_12284,N_13248);
or U15673 (N_15673,N_12555,N_13537);
or U15674 (N_15674,N_12004,N_12725);
xor U15675 (N_15675,N_12567,N_13505);
nand U15676 (N_15676,N_12571,N_12433);
xor U15677 (N_15677,N_12506,N_13867);
nand U15678 (N_15678,N_12355,N_12552);
xnor U15679 (N_15679,N_12874,N_12384);
xnor U15680 (N_15680,N_13346,N_13737);
xnor U15681 (N_15681,N_13426,N_12251);
nor U15682 (N_15682,N_13953,N_13888);
and U15683 (N_15683,N_12982,N_12156);
and U15684 (N_15684,N_13939,N_12536);
nand U15685 (N_15685,N_12659,N_12552);
or U15686 (N_15686,N_12027,N_13404);
nand U15687 (N_15687,N_12465,N_13135);
nand U15688 (N_15688,N_12104,N_13186);
xnor U15689 (N_15689,N_13553,N_12022);
and U15690 (N_15690,N_12918,N_12738);
or U15691 (N_15691,N_12697,N_12046);
or U15692 (N_15692,N_13100,N_12242);
nand U15693 (N_15693,N_13943,N_13137);
and U15694 (N_15694,N_13335,N_12583);
and U15695 (N_15695,N_12369,N_12288);
or U15696 (N_15696,N_12882,N_12630);
nand U15697 (N_15697,N_13198,N_13383);
xnor U15698 (N_15698,N_13887,N_12572);
xnor U15699 (N_15699,N_13278,N_13143);
nor U15700 (N_15700,N_13936,N_12951);
nor U15701 (N_15701,N_12631,N_13438);
or U15702 (N_15702,N_13834,N_13789);
xnor U15703 (N_15703,N_13267,N_12823);
xnor U15704 (N_15704,N_12227,N_12726);
xnor U15705 (N_15705,N_13304,N_12313);
or U15706 (N_15706,N_12441,N_12715);
and U15707 (N_15707,N_12980,N_12147);
or U15708 (N_15708,N_12867,N_13141);
xor U15709 (N_15709,N_12006,N_12492);
nor U15710 (N_15710,N_13901,N_13389);
and U15711 (N_15711,N_12358,N_13015);
nor U15712 (N_15712,N_12394,N_13989);
or U15713 (N_15713,N_12523,N_13057);
or U15714 (N_15714,N_12977,N_13565);
and U15715 (N_15715,N_12367,N_12594);
nand U15716 (N_15716,N_13414,N_13330);
or U15717 (N_15717,N_12291,N_13191);
and U15718 (N_15718,N_12903,N_13118);
nand U15719 (N_15719,N_12473,N_12654);
and U15720 (N_15720,N_13028,N_12878);
nand U15721 (N_15721,N_13696,N_13271);
and U15722 (N_15722,N_12349,N_13731);
nor U15723 (N_15723,N_12108,N_13025);
and U15724 (N_15724,N_13895,N_13356);
nand U15725 (N_15725,N_12860,N_12975);
or U15726 (N_15726,N_12388,N_13159);
nand U15727 (N_15727,N_12759,N_12378);
nor U15728 (N_15728,N_12718,N_13275);
xor U15729 (N_15729,N_13919,N_12415);
or U15730 (N_15730,N_12854,N_13324);
nand U15731 (N_15731,N_13267,N_13712);
nor U15732 (N_15732,N_12730,N_13614);
nand U15733 (N_15733,N_13928,N_13520);
and U15734 (N_15734,N_12464,N_13472);
or U15735 (N_15735,N_12556,N_13167);
or U15736 (N_15736,N_13019,N_13760);
nand U15737 (N_15737,N_13883,N_12328);
nand U15738 (N_15738,N_12459,N_12691);
and U15739 (N_15739,N_13681,N_13472);
or U15740 (N_15740,N_13002,N_12154);
xor U15741 (N_15741,N_13921,N_13512);
nor U15742 (N_15742,N_12485,N_12910);
xnor U15743 (N_15743,N_13441,N_12434);
nand U15744 (N_15744,N_13252,N_13972);
xnor U15745 (N_15745,N_13786,N_12101);
and U15746 (N_15746,N_13911,N_13642);
and U15747 (N_15747,N_13586,N_13831);
xor U15748 (N_15748,N_12234,N_12417);
or U15749 (N_15749,N_12409,N_13020);
nand U15750 (N_15750,N_13049,N_12865);
xor U15751 (N_15751,N_12285,N_12715);
or U15752 (N_15752,N_13226,N_12384);
and U15753 (N_15753,N_13502,N_13525);
xor U15754 (N_15754,N_13445,N_13375);
nor U15755 (N_15755,N_12976,N_12216);
nor U15756 (N_15756,N_13829,N_12928);
nand U15757 (N_15757,N_12430,N_13875);
or U15758 (N_15758,N_12167,N_13141);
nor U15759 (N_15759,N_12739,N_12414);
nor U15760 (N_15760,N_12157,N_13675);
or U15761 (N_15761,N_13476,N_13074);
or U15762 (N_15762,N_13876,N_13099);
xnor U15763 (N_15763,N_12776,N_13356);
or U15764 (N_15764,N_12806,N_12084);
xnor U15765 (N_15765,N_12938,N_12207);
and U15766 (N_15766,N_12125,N_13969);
xnor U15767 (N_15767,N_13731,N_12561);
nor U15768 (N_15768,N_13536,N_12692);
xnor U15769 (N_15769,N_12554,N_13270);
xnor U15770 (N_15770,N_12890,N_13049);
or U15771 (N_15771,N_12371,N_13209);
nand U15772 (N_15772,N_12430,N_12041);
and U15773 (N_15773,N_13331,N_12359);
and U15774 (N_15774,N_12327,N_12136);
nor U15775 (N_15775,N_12458,N_12921);
nand U15776 (N_15776,N_13162,N_13501);
nor U15777 (N_15777,N_13473,N_13714);
or U15778 (N_15778,N_13630,N_13284);
nor U15779 (N_15779,N_13609,N_12106);
and U15780 (N_15780,N_12050,N_12850);
and U15781 (N_15781,N_13092,N_12406);
xnor U15782 (N_15782,N_12868,N_12036);
or U15783 (N_15783,N_12818,N_12205);
and U15784 (N_15784,N_13060,N_13955);
and U15785 (N_15785,N_13193,N_12595);
nor U15786 (N_15786,N_12437,N_12471);
or U15787 (N_15787,N_12611,N_13355);
or U15788 (N_15788,N_12972,N_13136);
and U15789 (N_15789,N_12498,N_12355);
nor U15790 (N_15790,N_13082,N_12534);
and U15791 (N_15791,N_13946,N_12659);
nor U15792 (N_15792,N_13386,N_12347);
nor U15793 (N_15793,N_13213,N_13554);
or U15794 (N_15794,N_12549,N_12975);
and U15795 (N_15795,N_12998,N_13228);
and U15796 (N_15796,N_13888,N_13490);
or U15797 (N_15797,N_13825,N_12270);
and U15798 (N_15798,N_12459,N_12003);
or U15799 (N_15799,N_12238,N_13788);
nand U15800 (N_15800,N_13927,N_12393);
and U15801 (N_15801,N_12351,N_13479);
nand U15802 (N_15802,N_13652,N_13222);
nand U15803 (N_15803,N_13256,N_13632);
nor U15804 (N_15804,N_12696,N_13353);
nand U15805 (N_15805,N_12617,N_13835);
xor U15806 (N_15806,N_12290,N_12443);
nor U15807 (N_15807,N_13433,N_13102);
and U15808 (N_15808,N_12514,N_12979);
and U15809 (N_15809,N_12079,N_13695);
nor U15810 (N_15810,N_12287,N_13735);
or U15811 (N_15811,N_13115,N_12523);
xnor U15812 (N_15812,N_12082,N_12969);
xor U15813 (N_15813,N_12096,N_13551);
nor U15814 (N_15814,N_12397,N_13312);
nor U15815 (N_15815,N_13615,N_13228);
or U15816 (N_15816,N_12165,N_13966);
nand U15817 (N_15817,N_13452,N_13618);
and U15818 (N_15818,N_13534,N_12311);
nor U15819 (N_15819,N_13158,N_12994);
nor U15820 (N_15820,N_12873,N_12865);
nand U15821 (N_15821,N_12779,N_13927);
nor U15822 (N_15822,N_12034,N_13345);
nand U15823 (N_15823,N_13411,N_12629);
xor U15824 (N_15824,N_12935,N_13687);
xnor U15825 (N_15825,N_12813,N_13240);
or U15826 (N_15826,N_13807,N_12550);
or U15827 (N_15827,N_13462,N_13400);
xnor U15828 (N_15828,N_13735,N_12676);
or U15829 (N_15829,N_12273,N_12859);
and U15830 (N_15830,N_13164,N_12147);
or U15831 (N_15831,N_12220,N_12665);
nand U15832 (N_15832,N_12046,N_12756);
and U15833 (N_15833,N_13114,N_13382);
or U15834 (N_15834,N_12478,N_12177);
xor U15835 (N_15835,N_13104,N_13291);
nand U15836 (N_15836,N_12130,N_12968);
or U15837 (N_15837,N_13457,N_13422);
xnor U15838 (N_15838,N_12498,N_12588);
nor U15839 (N_15839,N_13254,N_13897);
or U15840 (N_15840,N_12705,N_13374);
and U15841 (N_15841,N_12858,N_12282);
and U15842 (N_15842,N_13772,N_12715);
and U15843 (N_15843,N_13570,N_13325);
xnor U15844 (N_15844,N_13401,N_12326);
and U15845 (N_15845,N_12656,N_13361);
or U15846 (N_15846,N_13928,N_12803);
xnor U15847 (N_15847,N_13382,N_12769);
nor U15848 (N_15848,N_12028,N_13564);
nand U15849 (N_15849,N_13985,N_12626);
xnor U15850 (N_15850,N_13094,N_13606);
xnor U15851 (N_15851,N_12808,N_12458);
nand U15852 (N_15852,N_12533,N_12003);
nor U15853 (N_15853,N_13455,N_13505);
xnor U15854 (N_15854,N_13215,N_13130);
xor U15855 (N_15855,N_12562,N_12957);
and U15856 (N_15856,N_13122,N_13243);
nor U15857 (N_15857,N_13375,N_12616);
nand U15858 (N_15858,N_13364,N_12053);
or U15859 (N_15859,N_12116,N_12814);
nand U15860 (N_15860,N_13539,N_12097);
or U15861 (N_15861,N_13880,N_12873);
xnor U15862 (N_15862,N_12358,N_12198);
or U15863 (N_15863,N_13827,N_13654);
nor U15864 (N_15864,N_12847,N_13579);
or U15865 (N_15865,N_13218,N_13179);
and U15866 (N_15866,N_13332,N_12082);
or U15867 (N_15867,N_12879,N_13719);
or U15868 (N_15868,N_12562,N_13841);
and U15869 (N_15869,N_13742,N_13984);
nand U15870 (N_15870,N_13025,N_13148);
nor U15871 (N_15871,N_12307,N_12927);
nor U15872 (N_15872,N_13842,N_12625);
and U15873 (N_15873,N_13141,N_12986);
xnor U15874 (N_15874,N_13909,N_12507);
and U15875 (N_15875,N_12542,N_12827);
nand U15876 (N_15876,N_12171,N_13985);
and U15877 (N_15877,N_13603,N_13128);
or U15878 (N_15878,N_12937,N_12775);
nor U15879 (N_15879,N_13334,N_13243);
nand U15880 (N_15880,N_13528,N_12572);
xor U15881 (N_15881,N_13793,N_12756);
or U15882 (N_15882,N_13939,N_13416);
and U15883 (N_15883,N_12403,N_12071);
xnor U15884 (N_15884,N_12570,N_12696);
nor U15885 (N_15885,N_13435,N_13720);
nand U15886 (N_15886,N_12674,N_13428);
xor U15887 (N_15887,N_13673,N_12776);
and U15888 (N_15888,N_12172,N_13829);
xor U15889 (N_15889,N_12503,N_12787);
nand U15890 (N_15890,N_13045,N_13965);
xnor U15891 (N_15891,N_12351,N_13956);
or U15892 (N_15892,N_13036,N_13649);
and U15893 (N_15893,N_13588,N_12579);
xor U15894 (N_15894,N_12931,N_13567);
nor U15895 (N_15895,N_12274,N_12157);
xor U15896 (N_15896,N_12992,N_12505);
xnor U15897 (N_15897,N_12233,N_13222);
nand U15898 (N_15898,N_13067,N_13507);
xnor U15899 (N_15899,N_13534,N_12107);
xor U15900 (N_15900,N_13755,N_13830);
xnor U15901 (N_15901,N_13463,N_12282);
nand U15902 (N_15902,N_13694,N_13087);
nand U15903 (N_15903,N_12926,N_13702);
nor U15904 (N_15904,N_13804,N_13578);
nor U15905 (N_15905,N_13366,N_12530);
xor U15906 (N_15906,N_13017,N_13401);
or U15907 (N_15907,N_12840,N_13388);
or U15908 (N_15908,N_12704,N_12050);
or U15909 (N_15909,N_13911,N_13941);
or U15910 (N_15910,N_12321,N_13656);
and U15911 (N_15911,N_12314,N_13800);
and U15912 (N_15912,N_13242,N_12232);
xor U15913 (N_15913,N_12288,N_13710);
or U15914 (N_15914,N_12378,N_12782);
nor U15915 (N_15915,N_12923,N_12264);
and U15916 (N_15916,N_13008,N_13785);
nor U15917 (N_15917,N_12629,N_13420);
nor U15918 (N_15918,N_12656,N_12757);
xor U15919 (N_15919,N_13087,N_13189);
nand U15920 (N_15920,N_12186,N_13654);
nand U15921 (N_15921,N_13927,N_12455);
nand U15922 (N_15922,N_13247,N_12707);
or U15923 (N_15923,N_13513,N_12005);
nor U15924 (N_15924,N_12574,N_13687);
and U15925 (N_15925,N_12144,N_13521);
nor U15926 (N_15926,N_12717,N_13535);
or U15927 (N_15927,N_12057,N_12935);
nor U15928 (N_15928,N_12612,N_12023);
nor U15929 (N_15929,N_13342,N_12241);
nor U15930 (N_15930,N_13690,N_12182);
nand U15931 (N_15931,N_13069,N_12975);
nand U15932 (N_15932,N_12808,N_13305);
nor U15933 (N_15933,N_12184,N_13612);
and U15934 (N_15934,N_12750,N_12696);
xnor U15935 (N_15935,N_13801,N_13936);
nand U15936 (N_15936,N_12487,N_13585);
nand U15937 (N_15937,N_12779,N_12723);
xnor U15938 (N_15938,N_12481,N_13323);
nor U15939 (N_15939,N_13335,N_12457);
xor U15940 (N_15940,N_13891,N_12682);
nor U15941 (N_15941,N_13100,N_12800);
nor U15942 (N_15942,N_12191,N_12718);
nand U15943 (N_15943,N_13366,N_13642);
nand U15944 (N_15944,N_12839,N_12620);
and U15945 (N_15945,N_13182,N_12423);
nand U15946 (N_15946,N_12524,N_12217);
nor U15947 (N_15947,N_12830,N_12045);
nor U15948 (N_15948,N_13472,N_12007);
and U15949 (N_15949,N_12076,N_13010);
or U15950 (N_15950,N_13530,N_13700);
nor U15951 (N_15951,N_12729,N_12275);
or U15952 (N_15952,N_12654,N_12966);
xnor U15953 (N_15953,N_13859,N_12532);
or U15954 (N_15954,N_13153,N_12436);
nor U15955 (N_15955,N_12309,N_13471);
nand U15956 (N_15956,N_13409,N_13029);
nor U15957 (N_15957,N_12602,N_12859);
or U15958 (N_15958,N_12355,N_12974);
nor U15959 (N_15959,N_13125,N_12214);
xnor U15960 (N_15960,N_12869,N_13406);
or U15961 (N_15961,N_13721,N_13294);
xor U15962 (N_15962,N_12615,N_13771);
xor U15963 (N_15963,N_13097,N_13225);
nand U15964 (N_15964,N_13426,N_13685);
nand U15965 (N_15965,N_12222,N_13161);
and U15966 (N_15966,N_12516,N_12663);
xor U15967 (N_15967,N_13560,N_12801);
or U15968 (N_15968,N_13653,N_13349);
and U15969 (N_15969,N_12262,N_13372);
and U15970 (N_15970,N_13574,N_12576);
nand U15971 (N_15971,N_13345,N_12457);
nand U15972 (N_15972,N_12401,N_13848);
and U15973 (N_15973,N_13858,N_13742);
and U15974 (N_15974,N_12404,N_13402);
and U15975 (N_15975,N_12608,N_12768);
and U15976 (N_15976,N_13040,N_13100);
nor U15977 (N_15977,N_12858,N_13987);
nor U15978 (N_15978,N_12667,N_12739);
nand U15979 (N_15979,N_12342,N_12836);
or U15980 (N_15980,N_13480,N_12339);
or U15981 (N_15981,N_12259,N_12136);
xnor U15982 (N_15982,N_13906,N_13001);
nor U15983 (N_15983,N_13485,N_12134);
nand U15984 (N_15984,N_13170,N_12598);
or U15985 (N_15985,N_12503,N_12868);
nand U15986 (N_15986,N_12370,N_12926);
or U15987 (N_15987,N_13802,N_12652);
nor U15988 (N_15988,N_13032,N_13857);
nand U15989 (N_15989,N_12684,N_12626);
nor U15990 (N_15990,N_12632,N_13640);
nand U15991 (N_15991,N_13905,N_13264);
or U15992 (N_15992,N_13658,N_12804);
or U15993 (N_15993,N_12926,N_12003);
xnor U15994 (N_15994,N_12536,N_13385);
xnor U15995 (N_15995,N_13082,N_12725);
nand U15996 (N_15996,N_12807,N_13322);
nor U15997 (N_15997,N_12394,N_13066);
nand U15998 (N_15998,N_13512,N_12003);
or U15999 (N_15999,N_12603,N_13506);
nor U16000 (N_16000,N_14736,N_14143);
or U16001 (N_16001,N_15083,N_14251);
nor U16002 (N_16002,N_15450,N_14370);
nor U16003 (N_16003,N_15247,N_14089);
or U16004 (N_16004,N_14844,N_15966);
and U16005 (N_16005,N_14630,N_14620);
xor U16006 (N_16006,N_15105,N_14674);
xor U16007 (N_16007,N_15600,N_15315);
nor U16008 (N_16008,N_15778,N_14715);
xor U16009 (N_16009,N_15486,N_15972);
or U16010 (N_16010,N_15408,N_15789);
or U16011 (N_16011,N_15165,N_14946);
xnor U16012 (N_16012,N_15103,N_14778);
nor U16013 (N_16013,N_14903,N_14995);
nor U16014 (N_16014,N_14244,N_15442);
xor U16015 (N_16015,N_15380,N_15825);
nor U16016 (N_16016,N_15999,N_14781);
or U16017 (N_16017,N_14074,N_14739);
and U16018 (N_16018,N_15301,N_14261);
or U16019 (N_16019,N_15494,N_15181);
and U16020 (N_16020,N_14256,N_15582);
nor U16021 (N_16021,N_14317,N_15296);
nand U16022 (N_16022,N_15608,N_14327);
and U16023 (N_16023,N_15762,N_14664);
nor U16024 (N_16024,N_14455,N_15751);
or U16025 (N_16025,N_14612,N_14610);
nand U16026 (N_16026,N_15548,N_14889);
and U16027 (N_16027,N_14274,N_15655);
and U16028 (N_16028,N_14238,N_14449);
nor U16029 (N_16029,N_14085,N_14894);
nor U16030 (N_16030,N_14146,N_14094);
xor U16031 (N_16031,N_14058,N_14158);
or U16032 (N_16032,N_15903,N_14044);
nand U16033 (N_16033,N_14631,N_15588);
xor U16034 (N_16034,N_14341,N_14895);
nand U16035 (N_16035,N_14276,N_15962);
nand U16036 (N_16036,N_15777,N_14770);
and U16037 (N_16037,N_15914,N_14651);
nand U16038 (N_16038,N_15680,N_15506);
nor U16039 (N_16039,N_15458,N_14979);
nand U16040 (N_16040,N_15696,N_14281);
nor U16041 (N_16041,N_14694,N_15515);
xor U16042 (N_16042,N_15550,N_15091);
xnor U16043 (N_16043,N_14282,N_14371);
and U16044 (N_16044,N_14354,N_14452);
nand U16045 (N_16045,N_15078,N_14167);
nor U16046 (N_16046,N_15695,N_14078);
or U16047 (N_16047,N_15243,N_15362);
nand U16048 (N_16048,N_15415,N_15736);
or U16049 (N_16049,N_15421,N_14975);
or U16050 (N_16050,N_14788,N_15463);
and U16051 (N_16051,N_15743,N_14800);
nor U16052 (N_16052,N_15995,N_15270);
or U16053 (N_16053,N_15146,N_14734);
nor U16054 (N_16054,N_14666,N_15116);
xnor U16055 (N_16055,N_15724,N_15794);
nor U16056 (N_16056,N_14120,N_15395);
xnor U16057 (N_16057,N_14223,N_15709);
nand U16058 (N_16058,N_14291,N_14095);
nand U16059 (N_16059,N_14421,N_15788);
nand U16060 (N_16060,N_15213,N_15454);
nor U16061 (N_16061,N_15166,N_14220);
xnor U16062 (N_16062,N_14743,N_15882);
or U16063 (N_16063,N_14791,N_14575);
or U16064 (N_16064,N_14640,N_14320);
nand U16065 (N_16065,N_15446,N_14717);
xor U16066 (N_16066,N_14249,N_15796);
nand U16067 (N_16067,N_15005,N_14811);
and U16068 (N_16068,N_15341,N_15924);
nand U16069 (N_16069,N_15178,N_14346);
nor U16070 (N_16070,N_15244,N_14834);
xnor U16071 (N_16071,N_14269,N_15644);
nor U16072 (N_16072,N_14542,N_15417);
or U16073 (N_16073,N_14713,N_14657);
and U16074 (N_16074,N_15536,N_14339);
nor U16075 (N_16075,N_15209,N_15635);
nand U16076 (N_16076,N_14698,N_15858);
nand U16077 (N_16077,N_15441,N_15356);
and U16078 (N_16078,N_14672,N_14553);
nor U16079 (N_16079,N_15014,N_15856);
or U16080 (N_16080,N_15969,N_14797);
xnor U16081 (N_16081,N_15241,N_14295);
nor U16082 (N_16082,N_15823,N_14842);
and U16083 (N_16083,N_14121,N_15212);
and U16084 (N_16084,N_15674,N_15003);
and U16085 (N_16085,N_14932,N_15568);
and U16086 (N_16086,N_15854,N_15431);
or U16087 (N_16087,N_14767,N_14350);
xnor U16088 (N_16088,N_14031,N_15990);
nand U16089 (N_16089,N_14056,N_15697);
xor U16090 (N_16090,N_14192,N_14377);
and U16091 (N_16091,N_15836,N_14125);
xor U16092 (N_16092,N_15922,N_14447);
and U16093 (N_16093,N_15386,N_15714);
nor U16094 (N_16094,N_14272,N_14373);
or U16095 (N_16095,N_15394,N_15916);
nand U16096 (N_16096,N_15367,N_15612);
or U16097 (N_16097,N_15862,N_14827);
or U16098 (N_16098,N_14547,N_15991);
and U16099 (N_16099,N_14207,N_15671);
nand U16100 (N_16100,N_15578,N_14200);
nor U16101 (N_16101,N_14983,N_15346);
nand U16102 (N_16102,N_15797,N_14003);
or U16103 (N_16103,N_14599,N_15719);
and U16104 (N_16104,N_14073,N_14821);
nor U16105 (N_16105,N_14145,N_15487);
xor U16106 (N_16106,N_15867,N_15305);
or U16107 (N_16107,N_14904,N_14991);
and U16108 (N_16108,N_15514,N_15760);
or U16109 (N_16109,N_14805,N_14388);
nor U16110 (N_16110,N_14255,N_15511);
nor U16111 (N_16111,N_14619,N_15143);
nor U16112 (N_16112,N_14213,N_15370);
nand U16113 (N_16113,N_14087,N_14212);
nor U16114 (N_16114,N_14773,N_14488);
xnor U16115 (N_16115,N_14695,N_14460);
nand U16116 (N_16116,N_15616,N_14551);
and U16117 (N_16117,N_15598,N_15159);
nand U16118 (N_16118,N_15521,N_15574);
xnor U16119 (N_16119,N_14675,N_14835);
xnor U16120 (N_16120,N_15253,N_14337);
or U16121 (N_16121,N_14549,N_14825);
or U16122 (N_16122,N_15526,N_14495);
or U16123 (N_16123,N_14925,N_14755);
or U16124 (N_16124,N_14086,N_15054);
or U16125 (N_16125,N_15237,N_15012);
and U16126 (N_16126,N_14275,N_15281);
xor U16127 (N_16127,N_15733,N_14430);
and U16128 (N_16128,N_15145,N_14159);
nor U16129 (N_16129,N_14959,N_15002);
nand U16130 (N_16130,N_14182,N_14264);
and U16131 (N_16131,N_14434,N_15482);
nand U16132 (N_16132,N_14165,N_14497);
and U16133 (N_16133,N_14309,N_15438);
nand U16134 (N_16134,N_14909,N_14535);
nor U16135 (N_16135,N_14629,N_15325);
or U16136 (N_16136,N_14266,N_14113);
and U16137 (N_16137,N_15610,N_15814);
nand U16138 (N_16138,N_14027,N_14208);
nor U16139 (N_16139,N_14479,N_15950);
nor U16140 (N_16140,N_14768,N_14225);
nand U16141 (N_16141,N_14880,N_15898);
and U16142 (N_16142,N_15749,N_14418);
nor U16143 (N_16143,N_14559,N_14018);
xnor U16144 (N_16144,N_14877,N_14002);
nand U16145 (N_16145,N_14926,N_14428);
and U16146 (N_16146,N_15744,N_15713);
xor U16147 (N_16147,N_15586,N_15018);
or U16148 (N_16148,N_14246,N_14253);
xnor U16149 (N_16149,N_15066,N_15955);
and U16150 (N_16150,N_14798,N_14845);
or U16151 (N_16151,N_14234,N_14693);
nor U16152 (N_16152,N_14187,N_14221);
nand U16153 (N_16153,N_14908,N_14417);
xor U16154 (N_16154,N_14096,N_15040);
xor U16155 (N_16155,N_14149,N_15859);
and U16156 (N_16156,N_15741,N_15566);
xor U16157 (N_16157,N_15755,N_14928);
nand U16158 (N_16158,N_15177,N_15099);
or U16159 (N_16159,N_14127,N_15126);
xor U16160 (N_16160,N_14712,N_14386);
nor U16161 (N_16161,N_14750,N_14673);
xor U16162 (N_16162,N_15812,N_15223);
and U16163 (N_16163,N_15208,N_15071);
nand U16164 (N_16164,N_15001,N_15119);
nand U16165 (N_16165,N_15705,N_14494);
xnor U16166 (N_16166,N_15101,N_14725);
xnor U16167 (N_16167,N_14466,N_14563);
xor U16168 (N_16168,N_14705,N_15601);
and U16169 (N_16169,N_15140,N_14133);
nor U16170 (N_16170,N_15987,N_14911);
nand U16171 (N_16171,N_14037,N_15770);
nand U16172 (N_16172,N_15860,N_15011);
or U16173 (N_16173,N_15965,N_15915);
xor U16174 (N_16174,N_15492,N_14558);
xnor U16175 (N_16175,N_15411,N_14950);
xnor U16176 (N_16176,N_15469,N_14980);
nor U16177 (N_16177,N_14597,N_14526);
nand U16178 (N_16178,N_14544,N_15410);
xnor U16179 (N_16179,N_15470,N_14528);
nand U16180 (N_16180,N_14548,N_15874);
xor U16181 (N_16181,N_15352,N_14247);
xor U16182 (N_16182,N_15552,N_15210);
nand U16183 (N_16183,N_15654,N_15747);
and U16184 (N_16184,N_15803,N_15436);
and U16185 (N_16185,N_15685,N_14190);
nand U16186 (N_16186,N_15925,N_15282);
or U16187 (N_16187,N_14410,N_14570);
and U16188 (N_16188,N_14202,N_15382);
or U16189 (N_16189,N_14314,N_15134);
and U16190 (N_16190,N_15834,N_14571);
nor U16191 (N_16191,N_15535,N_15285);
or U16192 (N_16192,N_14878,N_14738);
nor U16193 (N_16193,N_15988,N_14016);
or U16194 (N_16194,N_15840,N_15052);
nor U16195 (N_16195,N_15712,N_15031);
nand U16196 (N_16196,N_14965,N_15848);
nor U16197 (N_16197,N_15636,N_15868);
or U16198 (N_16198,N_15483,N_15871);
nor U16199 (N_16199,N_14901,N_14652);
or U16200 (N_16200,N_14365,N_15656);
or U16201 (N_16201,N_14776,N_15093);
and U16202 (N_16202,N_14680,N_14049);
and U16203 (N_16203,N_14484,N_15553);
nor U16204 (N_16204,N_15043,N_14573);
and U16205 (N_16205,N_15985,N_14333);
or U16206 (N_16206,N_14179,N_14342);
nor U16207 (N_16207,N_14067,N_15219);
or U16208 (N_16208,N_15646,N_15484);
nand U16209 (N_16209,N_14432,N_15707);
nand U16210 (N_16210,N_14828,N_14013);
or U16211 (N_16211,N_15503,N_15038);
nor U16212 (N_16212,N_14440,N_15184);
nand U16213 (N_16213,N_14872,N_15288);
and U16214 (N_16214,N_14112,N_15102);
xor U16215 (N_16215,N_14870,N_15984);
and U16216 (N_16216,N_15114,N_14476);
and U16217 (N_16217,N_14357,N_15307);
or U16218 (N_16218,N_14458,N_14730);
nand U16219 (N_16219,N_14245,N_15308);
or U16220 (N_16220,N_14283,N_14316);
xnor U16221 (N_16221,N_15248,N_15306);
and U16222 (N_16222,N_15629,N_14775);
xor U16223 (N_16223,N_15355,N_15224);
and U16224 (N_16224,N_15400,N_14057);
xor U16225 (N_16225,N_15088,N_15993);
xnor U16226 (N_16226,N_14948,N_14010);
and U16227 (N_16227,N_15518,N_15785);
nand U16228 (N_16228,N_14136,N_14009);
nor U16229 (N_16229,N_15912,N_15827);
and U16230 (N_16230,N_15425,N_15662);
nor U16231 (N_16231,N_15734,N_15485);
xor U16232 (N_16232,N_14823,N_15832);
or U16233 (N_16233,N_15693,N_15667);
xnor U16234 (N_16234,N_14756,N_14638);
or U16235 (N_16235,N_15405,N_15268);
and U16236 (N_16236,N_14607,N_14682);
nor U16237 (N_16237,N_15849,N_15138);
or U16238 (N_16238,N_15387,N_14332);
and U16239 (N_16239,N_14546,N_14941);
nor U16240 (N_16240,N_14017,N_14684);
nor U16241 (N_16241,N_15948,N_15833);
xnor U16242 (N_16242,N_14838,N_14389);
or U16243 (N_16243,N_15754,N_15689);
or U16244 (N_16244,N_14012,N_15742);
nor U16245 (N_16245,N_14391,N_14669);
nand U16246 (N_16246,N_15516,N_15949);
or U16247 (N_16247,N_15549,N_15222);
and U16248 (N_16248,N_15678,N_15074);
or U16249 (N_16249,N_15732,N_15905);
or U16250 (N_16250,N_14881,N_15187);
nand U16251 (N_16251,N_14142,N_15221);
nand U16252 (N_16252,N_15179,N_15344);
or U16253 (N_16253,N_14581,N_15008);
xnor U16254 (N_16254,N_14232,N_14855);
xor U16255 (N_16255,N_15543,N_15909);
nor U16256 (N_16256,N_14867,N_14242);
xor U16257 (N_16257,N_14921,N_14171);
nor U16258 (N_16258,N_14169,N_15414);
nand U16259 (N_16259,N_14794,N_15716);
and U16260 (N_16260,N_15593,N_15933);
or U16261 (N_16261,N_14191,N_15190);
nand U16262 (N_16262,N_14996,N_15108);
nand U16263 (N_16263,N_14092,N_15959);
nor U16264 (N_16264,N_14345,N_14248);
or U16265 (N_16265,N_15401,N_14853);
or U16266 (N_16266,N_14961,N_14564);
nor U16267 (N_16267,N_15121,N_15261);
nor U16268 (N_16268,N_14971,N_14661);
or U16269 (N_16269,N_14071,N_15540);
xor U16270 (N_16270,N_14514,N_14303);
and U16271 (N_16271,N_15118,N_15837);
nand U16272 (N_16272,N_14968,N_15626);
or U16273 (N_16273,N_14183,N_14045);
and U16274 (N_16274,N_14829,N_15249);
xnor U16275 (N_16275,N_15453,N_14662);
xnor U16276 (N_16276,N_14601,N_15802);
and U16277 (N_16277,N_14425,N_15853);
and U16278 (N_16278,N_15756,N_15954);
nand U16279 (N_16279,N_15064,N_14235);
and U16280 (N_16280,N_15923,N_15900);
or U16281 (N_16281,N_15215,N_14026);
and U16282 (N_16282,N_15319,N_15191);
nor U16283 (N_16283,N_15894,N_14659);
or U16284 (N_16284,N_15133,N_15917);
and U16285 (N_16285,N_15891,N_14701);
or U16286 (N_16286,N_15943,N_14347);
xor U16287 (N_16287,N_14847,N_14602);
nor U16288 (N_16288,N_14069,N_15198);
nor U16289 (N_16289,N_15499,N_15456);
or U16290 (N_16290,N_14329,N_15496);
nor U16291 (N_16291,N_15846,N_14617);
or U16292 (N_16292,N_15533,N_15721);
nand U16293 (N_16293,N_15058,N_14006);
and U16294 (N_16294,N_15613,N_15371);
xor U16295 (N_16295,N_15967,N_15231);
or U16296 (N_16296,N_15799,N_15182);
and U16297 (N_16297,N_15498,N_15227);
or U16298 (N_16298,N_15297,N_15176);
and U16299 (N_16299,N_14066,N_14038);
xnor U16300 (N_16300,N_15065,N_14076);
xor U16301 (N_16301,N_14539,N_15207);
or U16302 (N_16302,N_15973,N_14955);
or U16303 (N_16303,N_15877,N_15952);
and U16304 (N_16304,N_15639,N_14592);
nor U16305 (N_16305,N_14993,N_15677);
xnor U16306 (N_16306,N_15337,N_15561);
nand U16307 (N_16307,N_14195,N_14913);
and U16308 (N_16308,N_15911,N_15232);
and U16309 (N_16309,N_14040,N_15274);
nor U16310 (N_16310,N_15766,N_14874);
xor U16311 (N_16311,N_14456,N_14536);
and U16312 (N_16312,N_15542,N_15383);
or U16313 (N_16313,N_15508,N_14920);
nor U16314 (N_16314,N_14740,N_15945);
and U16315 (N_16315,N_15528,N_15791);
nand U16316 (N_16316,N_14751,N_14288);
nand U16317 (N_16317,N_14140,N_14450);
or U16318 (N_16318,N_14972,N_15081);
nor U16319 (N_16319,N_15545,N_15365);
nand U16320 (N_16320,N_14344,N_14565);
or U16321 (N_16321,N_14296,N_15218);
or U16322 (N_16322,N_14826,N_14338);
or U16323 (N_16323,N_15230,N_15378);
nand U16324 (N_16324,N_15541,N_14519);
nor U16325 (N_16325,N_14749,N_14005);
nand U16326 (N_16326,N_14902,N_14268);
and U16327 (N_16327,N_15385,N_14884);
and U16328 (N_16328,N_15045,N_15000);
nor U16329 (N_16329,N_14439,N_15614);
nor U16330 (N_16330,N_15746,N_14441);
or U16331 (N_16331,N_14915,N_15435);
xor U16332 (N_16332,N_14442,N_14382);
nand U16333 (N_16333,N_14819,N_14645);
and U16334 (N_16334,N_14922,N_15587);
nand U16335 (N_16335,N_14887,N_14493);
nand U16336 (N_16336,N_14379,N_15523);
nor U16337 (N_16337,N_14356,N_15653);
or U16338 (N_16338,N_15750,N_15938);
and U16339 (N_16339,N_15022,N_15072);
or U16340 (N_16340,N_14735,N_15532);
or U16341 (N_16341,N_15956,N_14958);
xor U16342 (N_16342,N_15475,N_14104);
nor U16343 (N_16343,N_15495,N_15885);
nand U16344 (N_16344,N_14075,N_14898);
nand U16345 (N_16345,N_14999,N_15951);
or U16346 (N_16346,N_15971,N_14046);
nor U16347 (N_16347,N_14807,N_15838);
or U16348 (N_16348,N_15185,N_15947);
nor U16349 (N_16349,N_14864,N_14839);
or U16350 (N_16350,N_15334,N_15590);
xor U16351 (N_16351,N_15360,N_15046);
nand U16352 (N_16352,N_14331,N_15564);
nor U16353 (N_16353,N_15339,N_15330);
nor U16354 (N_16354,N_15781,N_15089);
or U16355 (N_16355,N_14405,N_14298);
nor U16356 (N_16356,N_15028,N_14041);
nand U16357 (N_16357,N_15726,N_14611);
nand U16358 (N_16358,N_14832,N_15807);
nor U16359 (N_16359,N_15842,N_14728);
nor U16360 (N_16360,N_15761,N_15350);
nand U16361 (N_16361,N_15472,N_14433);
nand U16362 (N_16362,N_14478,N_15638);
nand U16363 (N_16363,N_14907,N_14804);
and U16364 (N_16364,N_14194,N_14369);
nand U16365 (N_16365,N_15419,N_14929);
or U16366 (N_16366,N_14608,N_15896);
nand U16367 (N_16367,N_14541,N_14636);
xnor U16368 (N_16368,N_15529,N_14806);
nand U16369 (N_16369,N_14992,N_14173);
or U16370 (N_16370,N_15476,N_14783);
or U16371 (N_16371,N_14683,N_15835);
or U16372 (N_16372,N_15783,N_14093);
nor U16373 (N_16373,N_14131,N_15448);
and U16374 (N_16374,N_14933,N_15464);
and U16375 (N_16375,N_14101,N_14240);
nand U16376 (N_16376,N_15094,N_14982);
xor U16377 (N_16377,N_15666,N_15457);
nand U16378 (N_16378,N_14063,N_15620);
nand U16379 (N_16379,N_15324,N_15625);
and U16380 (N_16380,N_14474,N_15267);
nor U16381 (N_16381,N_15277,N_15937);
nor U16382 (N_16382,N_15170,N_14550);
xnor U16383 (N_16383,N_15188,N_14023);
xor U16384 (N_16384,N_14977,N_14792);
and U16385 (N_16385,N_14205,N_15429);
nand U16386 (N_16386,N_15399,N_15136);
xnor U16387 (N_16387,N_14162,N_14916);
nand U16388 (N_16388,N_14030,N_15275);
nor U16389 (N_16389,N_14668,N_14688);
nor U16390 (N_16390,N_14893,N_14181);
nand U16391 (N_16391,N_14480,N_15919);
nand U16392 (N_16392,N_14711,N_14944);
and U16393 (N_16393,N_14764,N_14833);
nand U16394 (N_16394,N_14754,N_15537);
nand U16395 (N_16395,N_15201,N_14831);
nor U16396 (N_16396,N_15481,N_15664);
or U16397 (N_16397,N_14355,N_15351);
nor U16398 (N_16398,N_14803,N_15690);
xor U16399 (N_16399,N_14856,N_15975);
or U16400 (N_16400,N_14567,N_15748);
and U16401 (N_16401,N_15688,N_14362);
or U16402 (N_16402,N_15617,N_15567);
and U16403 (N_16403,N_14822,N_14325);
or U16404 (N_16404,N_14021,N_15701);
xor U16405 (N_16405,N_15953,N_14670);
nor U16406 (N_16406,N_14448,N_15100);
xor U16407 (N_16407,N_14352,N_14020);
xor U16408 (N_16408,N_14801,N_14518);
and U16409 (N_16409,N_15725,N_15353);
nor U16410 (N_16410,N_14679,N_14118);
or U16411 (N_16411,N_15621,N_15648);
xnor U16412 (N_16412,N_14733,N_14392);
nor U16413 (N_16413,N_15708,N_15026);
xnor U16414 (N_16414,N_14888,N_14957);
nor U16415 (N_16415,N_14917,N_15137);
xor U16416 (N_16416,N_14796,N_15220);
nor U16417 (N_16417,N_14985,N_14084);
nor U16418 (N_16418,N_14361,N_15041);
nor U16419 (N_16419,N_15168,N_15944);
nand U16420 (N_16420,N_14290,N_15776);
and U16421 (N_16421,N_15359,N_15013);
nor U16422 (N_16422,N_14525,N_15645);
and U16423 (N_16423,N_14988,N_15265);
nor U16424 (N_16424,N_14380,N_15266);
nor U16425 (N_16425,N_14393,N_15085);
nand U16426 (N_16426,N_14262,N_14859);
or U16427 (N_16427,N_14237,N_15595);
and U16428 (N_16428,N_15009,N_15607);
xor U16429 (N_16429,N_15283,N_14224);
and U16430 (N_16430,N_15125,N_14818);
and U16431 (N_16431,N_15793,N_15461);
nor U16432 (N_16432,N_14789,N_14924);
and U16433 (N_16433,N_14947,N_15424);
or U16434 (N_16434,N_14981,N_14891);
xnor U16435 (N_16435,N_15234,N_15556);
nand U16436 (N_16436,N_14252,N_14487);
nand U16437 (N_16437,N_14919,N_14577);
nand U16438 (N_16438,N_15148,N_14397);
nand U16439 (N_16439,N_14503,N_14472);
and U16440 (N_16440,N_14854,N_15633);
nand U16441 (N_16441,N_15828,N_15815);
and U16442 (N_16442,N_14624,N_15852);
xor U16443 (N_16443,N_15331,N_15731);
nand U16444 (N_16444,N_14278,N_15455);
nor U16445 (N_16445,N_15321,N_15377);
nor U16446 (N_16446,N_15197,N_14720);
and U16447 (N_16447,N_14697,N_15106);
and U16448 (N_16448,N_14411,N_15997);
nor U16449 (N_16449,N_14782,N_14938);
or U16450 (N_16450,N_15488,N_15530);
nand U16451 (N_16451,N_14896,N_15702);
nand U16452 (N_16452,N_14241,N_15687);
xor U16453 (N_16453,N_15512,N_14270);
nor U16454 (N_16454,N_15162,N_15131);
and U16455 (N_16455,N_15418,N_14485);
nand U16456 (N_16456,N_14746,N_14257);
xnor U16457 (N_16457,N_14060,N_14414);
or U16458 (N_16458,N_15167,N_14407);
or U16459 (N_16459,N_15963,N_14481);
nor U16460 (N_16460,N_15310,N_15142);
nor U16461 (N_16461,N_14032,N_14967);
xor U16462 (N_16462,N_14025,N_15067);
nand U16463 (N_16463,N_15665,N_14340);
nand U16464 (N_16464,N_15024,N_15772);
or U16465 (N_16465,N_14203,N_14090);
nand U16466 (N_16466,N_14359,N_14696);
xor U16467 (N_16467,N_14966,N_14155);
or U16468 (N_16468,N_14065,N_14422);
xnor U16469 (N_16469,N_15704,N_15557);
nand U16470 (N_16470,N_14545,N_14300);
nand U16471 (N_16471,N_15311,N_15745);
and U16472 (N_16472,N_14050,N_14349);
nand U16473 (N_16473,N_15700,N_14530);
nor U16474 (N_16474,N_15520,N_14731);
nand U16475 (N_16475,N_14882,N_15059);
or U16476 (N_16476,N_14130,N_14489);
xor U16477 (N_16477,N_15942,N_15447);
xnor U16478 (N_16478,N_14008,N_14412);
and U16479 (N_16479,N_15109,N_14204);
xor U16480 (N_16480,N_14939,N_15768);
nand U16481 (N_16481,N_15316,N_14492);
nand U16482 (N_16482,N_15910,N_15752);
nor U16483 (N_16483,N_15547,N_14615);
xnor U16484 (N_16484,N_15077,N_14576);
nand U16485 (N_16485,N_15873,N_15294);
xor U16486 (N_16486,N_15606,N_15501);
or U16487 (N_16487,N_14054,N_15194);
and U16488 (N_16488,N_15117,N_15682);
xnor U16489 (N_16489,N_14160,N_14862);
nor U16490 (N_16490,N_15706,N_14216);
and U16491 (N_16491,N_14394,N_14633);
or U16492 (N_16492,N_15252,N_14523);
or U16493 (N_16493,N_14228,N_14072);
or U16494 (N_16494,N_15027,N_15340);
nand U16495 (N_16495,N_15670,N_14584);
or U16496 (N_16496,N_14088,N_14554);
nor U16497 (N_16497,N_15104,N_14036);
or U16498 (N_16498,N_15030,N_14001);
nor U16499 (N_16499,N_15864,N_15869);
nand U16500 (N_16500,N_15642,N_14444);
xnor U16501 (N_16501,N_15519,N_14419);
nand U16502 (N_16502,N_14866,N_15782);
xnor U16503 (N_16503,N_14691,N_14572);
and U16504 (N_16504,N_15392,N_15787);
nand U16505 (N_16505,N_15444,N_14978);
nor U16506 (N_16506,N_15251,N_14267);
xnor U16507 (N_16507,N_14729,N_15402);
and U16508 (N_16508,N_15160,N_14555);
nand U16509 (N_16509,N_15149,N_14153);
nand U16510 (N_16510,N_14138,N_15818);
nand U16511 (N_16511,N_15976,N_14185);
nand U16512 (N_16512,N_14043,N_15591);
and U16513 (N_16513,N_15899,N_14520);
and U16514 (N_16514,N_14372,N_14068);
nand U16515 (N_16515,N_14157,N_14752);
nand U16516 (N_16516,N_14653,N_15242);
xnor U16517 (N_16517,N_15847,N_14227);
xnor U16518 (N_16518,N_15711,N_14897);
nor U16519 (N_16519,N_14742,N_14614);
and U16520 (N_16520,N_15144,N_14912);
xnor U16521 (N_16521,N_14000,N_14384);
and U16522 (N_16522,N_14569,N_15683);
and U16523 (N_16523,N_14132,N_15245);
nor U16524 (N_16524,N_14533,N_15703);
or U16525 (N_16525,N_15630,N_14222);
xor U16526 (N_16526,N_14144,N_14004);
or U16527 (N_16527,N_15130,N_14330);
nand U16528 (N_16528,N_14151,N_14593);
nor U16529 (N_16529,N_14562,N_14126);
nor U16530 (N_16530,N_15060,N_15336);
and U16531 (N_16531,N_15907,N_15879);
or U16532 (N_16532,N_15260,N_14353);
or U16533 (N_16533,N_14174,N_15430);
xor U16534 (N_16534,N_14445,N_14218);
and U16535 (N_16535,N_14134,N_14973);
xnor U16536 (N_16536,N_15889,N_15391);
nor U16537 (N_16537,N_15017,N_15264);
and U16538 (N_16538,N_15679,N_15964);
nand U16539 (N_16539,N_14462,N_14632);
nand U16540 (N_16540,N_15809,N_15660);
xor U16541 (N_16541,N_15669,N_15372);
or U16542 (N_16542,N_15958,N_15299);
nor U16543 (N_16543,N_14292,N_15255);
or U16544 (N_16544,N_15489,N_15152);
nor U16545 (N_16545,N_15396,N_15819);
and U16546 (N_16546,N_15998,N_14033);
and U16547 (N_16547,N_15141,N_14840);
and U16548 (N_16548,N_15676,N_14294);
and U16549 (N_16549,N_15565,N_14590);
nor U16550 (N_16550,N_15328,N_15684);
xnor U16551 (N_16551,N_14015,N_14820);
nand U16552 (N_16552,N_15699,N_14461);
and U16553 (N_16553,N_14304,N_14501);
or U16554 (N_16554,N_14817,N_15581);
and U16555 (N_16555,N_15111,N_14103);
nand U16556 (N_16556,N_14102,N_14766);
or U16557 (N_16557,N_14616,N_15172);
or U16558 (N_16558,N_14574,N_14007);
nor U16559 (N_16559,N_15037,N_15280);
or U16560 (N_16560,N_15773,N_15135);
and U16561 (N_16561,N_15006,N_14164);
xor U16562 (N_16562,N_14873,N_15525);
nand U16563 (N_16563,N_14502,N_14217);
or U16564 (N_16564,N_14471,N_14358);
and U16565 (N_16565,N_14201,N_14374);
and U16566 (N_16566,N_15936,N_14685);
xnor U16567 (N_16567,N_15632,N_14512);
or U16568 (N_16568,N_14598,N_14306);
xnor U16569 (N_16569,N_14605,N_14189);
and U16570 (N_16570,N_14906,N_14692);
or U16571 (N_16571,N_15686,N_15107);
nor U16572 (N_16572,N_15186,N_15361);
or U16573 (N_16573,N_14719,N_14129);
xor U16574 (N_16574,N_15289,N_14343);
and U16575 (N_16575,N_15196,N_15895);
xnor U16576 (N_16576,N_15661,N_14047);
xor U16577 (N_16577,N_15364,N_15157);
nor U16578 (N_16578,N_14387,N_15961);
nand U16579 (N_16579,N_15426,N_15865);
or U16580 (N_16580,N_14515,N_15007);
and U16581 (N_16581,N_14028,N_14589);
and U16582 (N_16582,N_15211,N_14406);
or U16583 (N_16583,N_15075,N_15774);
xor U16584 (N_16584,N_14029,N_15981);
nor U16585 (N_16585,N_15611,N_14588);
xnor U16586 (N_16586,N_14263,N_15407);
xnor U16587 (N_16587,N_15977,N_15300);
nand U16588 (N_16588,N_14677,N_15855);
nor U16589 (N_16589,N_14110,N_14656);
xnor U16590 (N_16590,N_15158,N_15658);
or U16591 (N_16591,N_15575,N_14319);
or U16592 (N_16592,N_15663,N_14336);
xnor U16593 (N_16593,N_15171,N_14626);
and U16594 (N_16594,N_15810,N_14622);
or U16595 (N_16595,N_15403,N_15497);
nor U16596 (N_16596,N_15579,N_15082);
and U16597 (N_16597,N_15982,N_14024);
nand U16598 (N_16598,N_14521,N_14453);
xnor U16599 (N_16599,N_14658,N_15694);
xor U16600 (N_16600,N_15738,N_15189);
xor U16601 (N_16601,N_15278,N_15049);
or U16602 (N_16602,N_14560,N_15546);
xor U16603 (N_16603,N_14970,N_15490);
and U16604 (N_16604,N_15675,N_15333);
xor U16605 (N_16605,N_15845,N_14475);
and U16606 (N_16606,N_14335,N_15327);
or U16607 (N_16607,N_14595,N_15238);
or U16608 (N_16608,N_14532,N_14375);
xnor U16609 (N_16609,N_15539,N_15409);
and U16610 (N_16610,N_14585,N_15228);
or U16611 (N_16611,N_14211,N_15246);
and U16612 (N_16612,N_14875,N_14082);
nor U16613 (N_16613,N_15622,N_14259);
or U16614 (N_16614,N_14865,N_15460);
nand U16615 (N_16615,N_15628,N_14506);
or U16616 (N_16616,N_15439,N_14150);
or U16617 (N_16617,N_15816,N_15817);
nand U16618 (N_16618,N_14048,N_15412);
and U16619 (N_16619,N_14443,N_14774);
nand U16620 (N_16620,N_14315,N_15573);
and U16621 (N_16621,N_14814,N_15594);
xor U16622 (N_16622,N_14732,N_14505);
and U16623 (N_16623,N_15291,N_14869);
nand U16624 (N_16624,N_15051,N_15767);
nor U16625 (N_16625,N_14771,N_14312);
nor U16626 (N_16626,N_15163,N_14148);
and U16627 (N_16627,N_14236,N_15374);
nand U16628 (N_16628,N_14284,N_15585);
nand U16629 (N_16629,N_14918,N_14537);
or U16630 (N_16630,N_14100,N_15326);
xnor U16631 (N_16631,N_14199,N_15513);
nor U16632 (N_16632,N_15878,N_14931);
nor U16633 (N_16633,N_15432,N_15509);
nand U16634 (N_16634,N_14952,N_15926);
and U16635 (N_16635,N_15576,N_14923);
nand U16636 (N_16636,N_14052,N_14543);
or U16637 (N_16637,N_15124,N_15691);
nor U16638 (N_16638,N_14810,N_14124);
xnor U16639 (N_16639,N_15931,N_15129);
nand U16640 (N_16640,N_15522,N_14876);
or U16641 (N_16641,N_14285,N_15284);
or U16642 (N_16642,N_14566,N_14976);
and U16643 (N_16643,N_14299,N_15589);
xnor U16644 (N_16644,N_14634,N_15259);
or U16645 (N_16645,N_14604,N_15147);
and U16646 (N_16646,N_15164,N_14301);
nor U16647 (N_16647,N_14513,N_15531);
nor U16648 (N_16648,N_15467,N_15069);
nand U16649 (N_16649,N_14473,N_15042);
or U16650 (N_16650,N_15569,N_15718);
nand U16651 (N_16651,N_15004,N_14757);
nor U16652 (N_16652,N_14403,N_14324);
xnor U16653 (N_16653,N_15183,N_15563);
or U16654 (N_16654,N_15015,N_15025);
and U16655 (N_16655,N_15427,N_14863);
or U16656 (N_16656,N_15035,N_14042);
xnor U16657 (N_16657,N_15068,N_14135);
nor U16658 (N_16658,N_15398,N_15239);
nand U16659 (N_16659,N_14128,N_15132);
nand U16660 (N_16660,N_14233,N_15056);
xnor U16661 (N_16661,N_14381,N_15657);
nor U16662 (N_16662,N_14531,N_14107);
xnor U16663 (N_16663,N_14106,N_15086);
nand U16664 (N_16664,N_15139,N_14424);
xor U16665 (N_16665,N_15887,N_15303);
and U16666 (N_16666,N_14699,N_15771);
nand U16667 (N_16667,N_14254,N_15449);
xor U16668 (N_16668,N_14077,N_14180);
nand U16669 (N_16669,N_15122,N_14363);
nor U16670 (N_16670,N_14671,N_15200);
nor U16671 (N_16671,N_15505,N_14168);
xnor U16672 (N_16672,N_14215,N_14648);
nor U16673 (N_16673,N_15290,N_15792);
or U16674 (N_16674,N_15863,N_15927);
nand U16675 (N_16675,N_14663,N_14399);
nand U16676 (N_16676,N_15668,N_14594);
nor U16677 (N_16677,N_14943,N_15098);
or U16678 (N_16678,N_14022,N_14197);
nor U16679 (N_16679,N_15866,N_14824);
or U16680 (N_16680,N_15960,N_15806);
nor U16681 (N_16681,N_15154,N_14280);
and U16682 (N_16682,N_14446,N_15354);
nor U16683 (N_16683,N_14986,N_14609);
or U16684 (N_16684,N_15206,N_15287);
and U16685 (N_16685,N_15920,N_15551);
or U16686 (N_16686,N_15804,N_14498);
nand U16687 (N_16687,N_14848,N_15605);
or U16688 (N_16688,N_15019,N_14079);
nor U16689 (N_16689,N_15805,N_14250);
nor U16690 (N_16690,N_15292,N_14426);
xor U16691 (N_16691,N_14930,N_14960);
and U16692 (N_16692,N_15560,N_15650);
or U16693 (N_16693,N_14949,N_15113);
and U16694 (N_16694,N_15957,N_14643);
or U16695 (N_16695,N_14760,N_14623);
and U16696 (N_16696,N_14846,N_15468);
nand U16697 (N_16697,N_15886,N_15389);
or U16698 (N_16698,N_14378,N_14660);
and U16699 (N_16699,N_15940,N_15048);
nand U16700 (N_16700,N_15764,N_15715);
nor U16701 (N_16701,N_15554,N_15822);
xnor U16702 (N_16702,N_14385,N_14366);
nor U16703 (N_16703,N_14690,N_14606);
and U16704 (N_16704,N_15723,N_15571);
nor U16705 (N_16705,N_14328,N_14177);
and U16706 (N_16706,N_15240,N_14469);
nand U16707 (N_16707,N_14219,N_14689);
xor U16708 (N_16708,N_15763,N_14364);
or U16709 (N_16709,N_15730,N_14061);
xor U16710 (N_16710,N_15692,N_14477);
nor U16711 (N_16711,N_14322,N_15225);
or U16712 (N_16712,N_15902,N_15216);
xnor U16713 (N_16713,N_14307,N_15153);
or U16714 (N_16714,N_14686,N_14176);
and U16715 (N_16715,N_15602,N_15884);
nor U16716 (N_16716,N_14721,N_14708);
and U16717 (N_16717,N_15204,N_15659);
or U16718 (N_16718,N_15544,N_14230);
or U16719 (N_16719,N_14511,N_14885);
or U16720 (N_16720,N_15020,N_15624);
nand U16721 (N_16721,N_15451,N_14166);
nor U16722 (N_16722,N_15775,N_14116);
xnor U16723 (N_16723,N_15343,N_14650);
nand U16724 (N_16724,N_15538,N_15465);
nor U16725 (N_16725,N_15881,N_14527);
xor U16726 (N_16726,N_15558,N_14787);
xnor U16727 (N_16727,N_15366,N_14070);
or U16728 (N_16728,N_14454,N_14508);
nor U16729 (N_16729,N_14500,N_14748);
or U16730 (N_16730,N_15090,N_14702);
nor U16731 (N_16731,N_15079,N_15928);
xor U16732 (N_16732,N_15044,N_15076);
nand U16733 (N_16733,N_15720,N_15935);
nor U16734 (N_16734,N_14198,N_14871);
nor U16735 (N_16735,N_15478,N_15298);
and U16736 (N_16736,N_15480,N_15623);
nor U16737 (N_16737,N_14723,N_15236);
nand U16738 (N_16738,N_14360,N_14790);
or U16739 (N_16739,N_14786,N_15829);
nor U16740 (N_16740,N_14302,N_14318);
or U16741 (N_16741,N_15986,N_14091);
and U16742 (N_16742,N_15811,N_14408);
or U16743 (N_16743,N_15850,N_15397);
nor U16744 (N_16744,N_14785,N_14716);
nor U16745 (N_16745,N_14396,N_15110);
xor U16746 (N_16746,N_14780,N_14311);
nor U16747 (N_16747,N_14637,N_15314);
or U16748 (N_16748,N_14753,N_14765);
nor U16749 (N_16749,N_14984,N_15890);
xnor U16750 (N_16750,N_15820,N_15717);
or U16751 (N_16751,N_15180,N_14667);
or U16752 (N_16752,N_14310,N_14522);
nand U16753 (N_16753,N_15175,N_14809);
nor U16754 (N_16754,N_15983,N_14139);
xor U16755 (N_16755,N_15422,N_15758);
xor U16756 (N_16756,N_15619,N_14308);
and U16757 (N_16757,N_15780,N_15271);
nor U16758 (N_16758,N_14997,N_15870);
and U16759 (N_16759,N_14900,N_15474);
nor U16760 (N_16760,N_15363,N_15618);
nand U16761 (N_16761,N_14178,N_15272);
and U16762 (N_16762,N_15368,N_14193);
xor U16763 (N_16763,N_14772,N_15839);
nor U16764 (N_16764,N_15649,N_15445);
nand U16765 (N_16765,N_14808,N_14402);
xnor U16766 (N_16766,N_14297,N_14286);
and U16767 (N_16767,N_15462,N_15876);
and U16768 (N_16768,N_14260,N_15073);
nand U16769 (N_16769,N_15517,N_15729);
nand U16770 (N_16770,N_14184,N_15379);
nand U16771 (N_16771,N_15021,N_15123);
or U16772 (N_16772,N_15323,N_15369);
or U16773 (N_16773,N_14097,N_15095);
nand U16774 (N_16774,N_15504,N_15637);
nor U16775 (N_16775,N_14722,N_15084);
or U16776 (N_16776,N_14137,N_15348);
nand U16777 (N_16777,N_15440,N_15786);
nand U16778 (N_16778,N_14596,N_15698);
or U16779 (N_16779,N_14051,N_15273);
and U16780 (N_16780,N_14777,N_15279);
nor U16781 (N_16781,N_15737,N_15813);
and U16782 (N_16782,N_15583,N_15826);
or U16783 (N_16783,N_15641,N_14161);
xor U16784 (N_16784,N_15735,N_14390);
nor U16785 (N_16785,N_14348,N_14927);
xnor U16786 (N_16786,N_15562,N_14059);
nor U16787 (N_16787,N_15795,N_14579);
nor U16788 (N_16788,N_15534,N_14289);
nor U16789 (N_16789,N_15390,N_15974);
xor U16790 (N_16790,N_14890,N_14843);
and U16791 (N_16791,N_14816,N_15250);
or U16792 (N_16792,N_14415,N_14510);
or U16793 (N_16793,N_15824,N_15087);
or U16794 (N_16794,N_14490,N_14451);
nor U16795 (N_16795,N_14524,N_15727);
nor U16796 (N_16796,N_14998,N_15115);
xor U16797 (N_16797,N_15801,N_14613);
xnor U16798 (N_16798,N_14758,N_14726);
nor U16799 (N_16799,N_14628,N_14857);
nor U16800 (N_16800,N_15577,N_15790);
nand U16801 (N_16801,N_14279,N_14108);
or U16802 (N_16802,N_15254,N_15062);
and U16803 (N_16803,N_14034,N_14540);
or U16804 (N_16804,N_14850,N_15437);
or U16805 (N_16805,N_15169,N_15647);
nor U16806 (N_16806,N_14676,N_14083);
nor U16807 (N_16807,N_14147,N_14470);
nor U16808 (N_16808,N_14724,N_15443);
nand U16809 (N_16809,N_15304,N_14861);
nand U16810 (N_16810,N_15318,N_15681);
and U16811 (N_16811,N_14517,N_14431);
xnor U16812 (N_16812,N_14639,N_14744);
nand U16813 (N_16813,N_14175,N_14404);
nor U16814 (N_16814,N_14293,N_15373);
nor U16815 (N_16815,N_14111,N_15128);
nand U16816 (N_16816,N_15673,N_14641);
or U16817 (N_16817,N_15096,N_14987);
or U16818 (N_16818,N_14463,N_14457);
nand U16819 (N_16819,N_14769,N_15524);
nor U16820 (N_16820,N_15968,N_14644);
or U16821 (N_16821,N_15404,N_15994);
nor U16822 (N_16822,N_15798,N_14305);
xor U16823 (N_16823,N_14964,N_14621);
nand U16824 (N_16824,N_14851,N_14557);
nor U16825 (N_16825,N_14156,N_15193);
xnor U16826 (N_16826,N_14586,N_14114);
nor U16827 (N_16827,N_15332,N_15643);
xnor U16828 (N_16828,N_15800,N_14383);
or U16829 (N_16829,N_14516,N_15500);
and U16830 (N_16830,N_15672,N_15120);
or U16831 (N_16831,N_15070,N_15631);
nor U16832 (N_16832,N_15235,N_14231);
or U16833 (N_16833,N_14035,N_14761);
or U16834 (N_16834,N_14868,N_14323);
or U16835 (N_16835,N_14762,N_14914);
nor U16836 (N_16836,N_15913,N_14934);
xor U16837 (N_16837,N_15572,N_14935);
nor U16838 (N_16838,N_15921,N_14759);
nand U16839 (N_16839,N_15502,N_14649);
and U16840 (N_16840,N_14287,N_15627);
nand U16841 (N_16841,N_14956,N_14940);
nand U16842 (N_16842,N_15112,N_15901);
and U16843 (N_16843,N_14423,N_14556);
nor U16844 (N_16844,N_15821,N_15640);
xor U16845 (N_16845,N_15603,N_14080);
and U16846 (N_16846,N_14813,N_14603);
nor U16847 (N_16847,N_14963,N_15939);
xnor U16848 (N_16848,N_14141,N_14271);
or U16849 (N_16849,N_14491,N_15205);
or U16850 (N_16850,N_14496,N_14438);
nand U16851 (N_16851,N_15053,N_14265);
nor U16852 (N_16852,N_15452,N_14974);
nand U16853 (N_16853,N_14618,N_14600);
nand U16854 (N_16854,N_15428,N_15342);
or U16855 (N_16855,N_15097,N_15883);
nor U16856 (N_16856,N_15580,N_14062);
or U16857 (N_16857,N_15203,N_15345);
and U16858 (N_16858,N_14486,N_14627);
xnor U16859 (N_16859,N_14681,N_15029);
or U16860 (N_16860,N_15036,N_15904);
nand U16861 (N_16861,N_14799,N_14994);
and U16862 (N_16862,N_14886,N_15226);
nand U16863 (N_16863,N_14578,N_15929);
nor U16864 (N_16864,N_15423,N_15880);
nor U16865 (N_16865,N_15375,N_14945);
or U16866 (N_16866,N_15970,N_14647);
or U16867 (N_16867,N_15233,N_14852);
or U16868 (N_16868,N_15493,N_14587);
nand U16869 (N_16869,N_15384,N_15831);
or U16870 (N_16870,N_15652,N_15039);
nor U16871 (N_16871,N_15830,N_15150);
nand U16872 (N_16872,N_14154,N_15393);
nand U16873 (N_16873,N_15420,N_14568);
and U16874 (N_16874,N_14465,N_14435);
and U16875 (N_16875,N_15016,N_14170);
xnor U16876 (N_16876,N_15381,N_15559);
nand U16877 (N_16877,N_14784,N_15202);
nor U16878 (N_16878,N_14105,N_14499);
nor U16879 (N_16879,N_15841,N_15269);
xor U16880 (N_16880,N_15584,N_14714);
and U16881 (N_16881,N_14313,N_15413);
xnor U16882 (N_16882,N_15263,N_15312);
nor U16883 (N_16883,N_14534,N_14109);
xnor U16884 (N_16884,N_15286,N_15293);
nand U16885 (N_16885,N_14243,N_15335);
nor U16886 (N_16886,N_14582,N_14706);
or U16887 (N_16887,N_15570,N_15338);
nand U16888 (N_16888,N_15710,N_15597);
and U16889 (N_16889,N_14123,N_15893);
nand U16890 (N_16890,N_15908,N_14529);
nand U16891 (N_16891,N_15295,N_14561);
nor U16892 (N_16892,N_15888,N_15349);
nor U16893 (N_16893,N_15527,N_15199);
and U16894 (N_16894,N_14321,N_15861);
and U16895 (N_16895,N_15434,N_14954);
nand U16896 (N_16896,N_15061,N_15256);
and U16897 (N_16897,N_14942,N_15599);
and U16898 (N_16898,N_15262,N_15055);
nor U16899 (N_16899,N_14119,N_15808);
nand U16900 (N_16900,N_15156,N_15875);
or U16901 (N_16901,N_15918,N_15634);
nor U16902 (N_16902,N_14152,N_15857);
xor U16903 (N_16903,N_14115,N_15033);
nor U16904 (N_16904,N_14704,N_14625);
xnor U16905 (N_16905,N_14459,N_15376);
nor U16906 (N_16906,N_15322,N_14226);
nand U16907 (N_16907,N_15851,N_15047);
nand U16908 (N_16908,N_15127,N_15192);
nand U16909 (N_16909,N_14580,N_14055);
or U16910 (N_16910,N_15479,N_14483);
or U16911 (N_16911,N_15174,N_15161);
nor U16912 (N_16912,N_14014,N_14413);
nor U16913 (N_16913,N_15980,N_15173);
or U16914 (N_16914,N_14879,N_14718);
and U16915 (N_16915,N_15843,N_14395);
or U16916 (N_16916,N_14707,N_15510);
and U16917 (N_16917,N_15739,N_14188);
nor U16918 (N_16918,N_15872,N_14277);
nand U16919 (N_16919,N_14812,N_14509);
nand U16920 (N_16920,N_15329,N_15080);
or U16921 (N_16921,N_15258,N_14905);
xor U16922 (N_16922,N_14099,N_14745);
or U16923 (N_16923,N_15214,N_15765);
nor U16924 (N_16924,N_14122,N_14214);
or U16925 (N_16925,N_14892,N_15507);
or U16926 (N_16926,N_14635,N_14951);
xnor U16927 (N_16927,N_14700,N_14703);
or U16928 (N_16928,N_14793,N_14376);
nand U16929 (N_16929,N_14011,N_14841);
xnor U16930 (N_16930,N_14937,N_14468);
and U16931 (N_16931,N_14186,N_14229);
and U16932 (N_16932,N_15932,N_14482);
nor U16933 (N_16933,N_14368,N_14507);
or U16934 (N_16934,N_15769,N_14642);
or U16935 (N_16935,N_14858,N_15609);
nand U16936 (N_16936,N_14665,N_14936);
or U16937 (N_16937,N_15032,N_14436);
and U16938 (N_16938,N_14962,N_15057);
or U16939 (N_16939,N_14779,N_15433);
nand U16940 (N_16940,N_14538,N_14953);
xor U16941 (N_16941,N_15477,N_14464);
or U16942 (N_16942,N_14400,N_15615);
nor U16943 (N_16943,N_14210,N_14117);
nand U16944 (N_16944,N_14429,N_14504);
xor U16945 (N_16945,N_15941,N_15759);
and U16946 (N_16946,N_15596,N_14398);
and U16947 (N_16947,N_14258,N_15906);
nand U16948 (N_16948,N_15844,N_14583);
or U16949 (N_16949,N_14709,N_14039);
or U16950 (N_16950,N_15309,N_15989);
and U16951 (N_16951,N_15406,N_14836);
or U16952 (N_16952,N_14990,N_14591);
or U16953 (N_16953,N_15320,N_15946);
or U16954 (N_16954,N_15276,N_14081);
nor U16955 (N_16955,N_15416,N_15466);
nor U16956 (N_16956,N_14737,N_15313);
or U16957 (N_16957,N_15357,N_14910);
nand U16958 (N_16958,N_14467,N_14019);
nand U16959 (N_16959,N_15092,N_15555);
or U16960 (N_16960,N_15784,N_15388);
nand U16961 (N_16961,N_14795,N_15302);
nand U16962 (N_16962,N_14351,N_14989);
and U16963 (N_16963,N_15978,N_14802);
nand U16964 (N_16964,N_15897,N_14172);
nand U16965 (N_16965,N_14206,N_14860);
xor U16966 (N_16966,N_15722,N_15010);
nand U16967 (N_16967,N_14815,N_15740);
or U16968 (N_16968,N_14837,N_14367);
nor U16969 (N_16969,N_14098,N_14334);
nand U16970 (N_16970,N_15979,N_15996);
xnor U16971 (N_16971,N_14727,N_15358);
and U16972 (N_16972,N_15471,N_14678);
nor U16973 (N_16973,N_14710,N_14209);
nand U16974 (N_16974,N_14163,N_15151);
or U16975 (N_16975,N_15753,N_14053);
nand U16976 (N_16976,N_15317,N_14883);
or U16977 (N_16977,N_15023,N_15459);
nor U16978 (N_16978,N_14899,N_15651);
or U16979 (N_16979,N_14273,N_14747);
or U16980 (N_16980,N_15779,N_15757);
nor U16981 (N_16981,N_15892,N_15992);
xor U16982 (N_16982,N_14326,N_15347);
or U16983 (N_16983,N_14830,N_15604);
xnor U16984 (N_16984,N_15034,N_14763);
xnor U16985 (N_16985,N_15592,N_14401);
and U16986 (N_16986,N_14420,N_15491);
xnor U16987 (N_16987,N_15229,N_14416);
or U16988 (N_16988,N_14687,N_14239);
and U16989 (N_16989,N_15930,N_14646);
nor U16990 (N_16990,N_15050,N_15728);
nand U16991 (N_16991,N_14409,N_14969);
nand U16992 (N_16992,N_14552,N_15257);
nand U16993 (N_16993,N_15195,N_14064);
or U16994 (N_16994,N_14655,N_14741);
nor U16995 (N_16995,N_15217,N_15473);
nor U16996 (N_16996,N_14437,N_15155);
nand U16997 (N_16997,N_15934,N_15063);
and U16998 (N_16998,N_14196,N_14849);
or U16999 (N_16999,N_14427,N_14654);
or U17000 (N_17000,N_14695,N_15179);
and U17001 (N_17001,N_14545,N_14258);
nand U17002 (N_17002,N_14747,N_14400);
or U17003 (N_17003,N_15408,N_15071);
xnor U17004 (N_17004,N_14256,N_14933);
xnor U17005 (N_17005,N_15847,N_14493);
and U17006 (N_17006,N_14707,N_14584);
nor U17007 (N_17007,N_15276,N_14947);
nand U17008 (N_17008,N_15072,N_15466);
and U17009 (N_17009,N_14035,N_14433);
and U17010 (N_17010,N_15761,N_15016);
xnor U17011 (N_17011,N_14516,N_15697);
nand U17012 (N_17012,N_14483,N_15066);
nor U17013 (N_17013,N_14992,N_15441);
nor U17014 (N_17014,N_14947,N_15734);
nor U17015 (N_17015,N_14259,N_14114);
nor U17016 (N_17016,N_15485,N_14342);
nand U17017 (N_17017,N_15287,N_14200);
xnor U17018 (N_17018,N_14446,N_15456);
xnor U17019 (N_17019,N_14467,N_15305);
or U17020 (N_17020,N_15173,N_15544);
nor U17021 (N_17021,N_15376,N_15880);
nand U17022 (N_17022,N_14528,N_14951);
xnor U17023 (N_17023,N_14929,N_14463);
nand U17024 (N_17024,N_15181,N_14499);
nor U17025 (N_17025,N_15367,N_14769);
nand U17026 (N_17026,N_15929,N_15913);
nor U17027 (N_17027,N_14571,N_15694);
xor U17028 (N_17028,N_14036,N_15610);
xnor U17029 (N_17029,N_15892,N_15781);
xor U17030 (N_17030,N_14767,N_15660);
or U17031 (N_17031,N_15136,N_15841);
nor U17032 (N_17032,N_14253,N_14393);
and U17033 (N_17033,N_15966,N_15519);
and U17034 (N_17034,N_14749,N_14932);
nand U17035 (N_17035,N_14835,N_14935);
or U17036 (N_17036,N_15891,N_14441);
or U17037 (N_17037,N_14056,N_14041);
or U17038 (N_17038,N_15655,N_14958);
and U17039 (N_17039,N_14750,N_15284);
and U17040 (N_17040,N_15330,N_15055);
and U17041 (N_17041,N_14057,N_14888);
nor U17042 (N_17042,N_15300,N_14811);
and U17043 (N_17043,N_15173,N_15894);
xor U17044 (N_17044,N_14557,N_14381);
and U17045 (N_17045,N_14964,N_14261);
xnor U17046 (N_17046,N_15467,N_14466);
xnor U17047 (N_17047,N_15769,N_14115);
xnor U17048 (N_17048,N_15808,N_14983);
and U17049 (N_17049,N_14999,N_15825);
and U17050 (N_17050,N_15764,N_14161);
or U17051 (N_17051,N_15066,N_14305);
xor U17052 (N_17052,N_15965,N_15901);
nand U17053 (N_17053,N_14696,N_14769);
xor U17054 (N_17054,N_15601,N_14788);
nand U17055 (N_17055,N_15264,N_14306);
and U17056 (N_17056,N_14901,N_14341);
xor U17057 (N_17057,N_15727,N_14345);
nor U17058 (N_17058,N_14638,N_14166);
xnor U17059 (N_17059,N_15339,N_14485);
nand U17060 (N_17060,N_14912,N_14616);
or U17061 (N_17061,N_15669,N_14404);
nand U17062 (N_17062,N_14931,N_14921);
or U17063 (N_17063,N_15132,N_15021);
nor U17064 (N_17064,N_15480,N_14281);
xnor U17065 (N_17065,N_14650,N_14774);
xor U17066 (N_17066,N_14668,N_14028);
or U17067 (N_17067,N_14978,N_14513);
nand U17068 (N_17068,N_14570,N_15344);
xor U17069 (N_17069,N_14813,N_14184);
and U17070 (N_17070,N_14989,N_14016);
nand U17071 (N_17071,N_14302,N_14215);
or U17072 (N_17072,N_15397,N_15386);
xnor U17073 (N_17073,N_14254,N_14748);
and U17074 (N_17074,N_15843,N_14541);
xor U17075 (N_17075,N_15091,N_14010);
nor U17076 (N_17076,N_15655,N_14063);
nand U17077 (N_17077,N_15895,N_14503);
nand U17078 (N_17078,N_14855,N_15269);
xor U17079 (N_17079,N_14368,N_14688);
and U17080 (N_17080,N_15932,N_15598);
or U17081 (N_17081,N_15962,N_14041);
xor U17082 (N_17082,N_14700,N_14099);
nand U17083 (N_17083,N_14415,N_15924);
xor U17084 (N_17084,N_15702,N_14691);
and U17085 (N_17085,N_14868,N_14552);
nand U17086 (N_17086,N_14113,N_14598);
and U17087 (N_17087,N_15990,N_14927);
nand U17088 (N_17088,N_14688,N_14715);
or U17089 (N_17089,N_15988,N_14855);
and U17090 (N_17090,N_14665,N_15658);
or U17091 (N_17091,N_14975,N_15281);
nor U17092 (N_17092,N_14886,N_15380);
and U17093 (N_17093,N_15276,N_14149);
nor U17094 (N_17094,N_15204,N_15366);
and U17095 (N_17095,N_14907,N_15049);
nor U17096 (N_17096,N_14647,N_15673);
and U17097 (N_17097,N_14352,N_14117);
nor U17098 (N_17098,N_15984,N_14576);
xnor U17099 (N_17099,N_15749,N_14295);
and U17100 (N_17100,N_15228,N_15580);
or U17101 (N_17101,N_14163,N_15067);
xnor U17102 (N_17102,N_15410,N_15814);
xnor U17103 (N_17103,N_14758,N_15527);
xnor U17104 (N_17104,N_14779,N_14198);
xnor U17105 (N_17105,N_14887,N_15301);
nand U17106 (N_17106,N_15244,N_15434);
nor U17107 (N_17107,N_14692,N_14100);
xnor U17108 (N_17108,N_15633,N_15480);
or U17109 (N_17109,N_15179,N_14673);
nand U17110 (N_17110,N_14636,N_15217);
nand U17111 (N_17111,N_15380,N_14139);
and U17112 (N_17112,N_14157,N_15993);
nand U17113 (N_17113,N_14680,N_14601);
nand U17114 (N_17114,N_14487,N_14763);
xor U17115 (N_17115,N_15887,N_15590);
nand U17116 (N_17116,N_14171,N_15222);
nand U17117 (N_17117,N_14339,N_15304);
and U17118 (N_17118,N_14510,N_14898);
xor U17119 (N_17119,N_14067,N_14054);
nor U17120 (N_17120,N_15996,N_14737);
nand U17121 (N_17121,N_14146,N_15889);
and U17122 (N_17122,N_15514,N_15521);
xnor U17123 (N_17123,N_14986,N_15705);
xnor U17124 (N_17124,N_14310,N_15970);
xor U17125 (N_17125,N_15498,N_15548);
and U17126 (N_17126,N_14692,N_15792);
nand U17127 (N_17127,N_14547,N_15451);
and U17128 (N_17128,N_15844,N_14283);
xor U17129 (N_17129,N_15448,N_15148);
nand U17130 (N_17130,N_14591,N_14316);
nor U17131 (N_17131,N_15416,N_14620);
or U17132 (N_17132,N_14878,N_14807);
xor U17133 (N_17133,N_14927,N_15654);
or U17134 (N_17134,N_14154,N_15817);
nor U17135 (N_17135,N_14503,N_14932);
and U17136 (N_17136,N_14853,N_14637);
nor U17137 (N_17137,N_14100,N_14836);
nand U17138 (N_17138,N_14834,N_14390);
nor U17139 (N_17139,N_14765,N_15630);
nor U17140 (N_17140,N_14923,N_14448);
or U17141 (N_17141,N_15144,N_15432);
nand U17142 (N_17142,N_15959,N_15410);
nor U17143 (N_17143,N_14050,N_15435);
and U17144 (N_17144,N_15094,N_14283);
xnor U17145 (N_17145,N_15926,N_15623);
xnor U17146 (N_17146,N_14638,N_14997);
nor U17147 (N_17147,N_14764,N_15133);
and U17148 (N_17148,N_15761,N_14032);
and U17149 (N_17149,N_14926,N_14624);
or U17150 (N_17150,N_14518,N_15345);
and U17151 (N_17151,N_14475,N_15114);
or U17152 (N_17152,N_15318,N_15250);
nand U17153 (N_17153,N_14017,N_14151);
nor U17154 (N_17154,N_15426,N_14909);
nor U17155 (N_17155,N_15387,N_15452);
nor U17156 (N_17156,N_14574,N_14272);
nor U17157 (N_17157,N_15087,N_15411);
xnor U17158 (N_17158,N_15063,N_14744);
or U17159 (N_17159,N_15602,N_14678);
xor U17160 (N_17160,N_14336,N_15392);
or U17161 (N_17161,N_15914,N_14438);
or U17162 (N_17162,N_15704,N_14846);
or U17163 (N_17163,N_15021,N_14243);
nand U17164 (N_17164,N_15138,N_15404);
nor U17165 (N_17165,N_14009,N_14464);
and U17166 (N_17166,N_14416,N_14480);
and U17167 (N_17167,N_14909,N_14757);
xnor U17168 (N_17168,N_14853,N_15963);
nand U17169 (N_17169,N_14274,N_14458);
nor U17170 (N_17170,N_14108,N_14586);
or U17171 (N_17171,N_15728,N_15482);
nor U17172 (N_17172,N_14738,N_14319);
and U17173 (N_17173,N_14891,N_15199);
and U17174 (N_17174,N_14065,N_14166);
or U17175 (N_17175,N_15548,N_14785);
nand U17176 (N_17176,N_15700,N_14416);
xnor U17177 (N_17177,N_15038,N_14616);
and U17178 (N_17178,N_14850,N_15870);
or U17179 (N_17179,N_14251,N_15007);
xor U17180 (N_17180,N_15793,N_15889);
or U17181 (N_17181,N_15948,N_14099);
nor U17182 (N_17182,N_15759,N_15412);
nor U17183 (N_17183,N_14733,N_15261);
nor U17184 (N_17184,N_14937,N_15552);
and U17185 (N_17185,N_14532,N_15578);
and U17186 (N_17186,N_15118,N_14887);
nor U17187 (N_17187,N_15352,N_15905);
xor U17188 (N_17188,N_14162,N_14272);
xnor U17189 (N_17189,N_14713,N_14241);
nor U17190 (N_17190,N_15143,N_14969);
xor U17191 (N_17191,N_14292,N_14752);
xnor U17192 (N_17192,N_15115,N_14297);
nor U17193 (N_17193,N_15694,N_14350);
nor U17194 (N_17194,N_15143,N_15092);
nand U17195 (N_17195,N_14253,N_14367);
nand U17196 (N_17196,N_15882,N_14345);
nor U17197 (N_17197,N_15744,N_14175);
and U17198 (N_17198,N_14797,N_15472);
and U17199 (N_17199,N_14712,N_15789);
or U17200 (N_17200,N_14802,N_14235);
nor U17201 (N_17201,N_14677,N_15747);
or U17202 (N_17202,N_15968,N_14889);
xor U17203 (N_17203,N_14700,N_15051);
or U17204 (N_17204,N_15865,N_14396);
or U17205 (N_17205,N_15461,N_15082);
or U17206 (N_17206,N_14663,N_14735);
and U17207 (N_17207,N_14463,N_15283);
xnor U17208 (N_17208,N_14857,N_14407);
nand U17209 (N_17209,N_14880,N_14319);
nor U17210 (N_17210,N_14591,N_15991);
nand U17211 (N_17211,N_14615,N_15426);
and U17212 (N_17212,N_15436,N_14924);
nor U17213 (N_17213,N_15675,N_14805);
xnor U17214 (N_17214,N_15899,N_14107);
and U17215 (N_17215,N_14906,N_14152);
xor U17216 (N_17216,N_15116,N_15414);
and U17217 (N_17217,N_14285,N_14394);
xor U17218 (N_17218,N_14985,N_14576);
nand U17219 (N_17219,N_14234,N_14347);
and U17220 (N_17220,N_15374,N_14338);
xnor U17221 (N_17221,N_15190,N_15171);
nor U17222 (N_17222,N_14275,N_14805);
nand U17223 (N_17223,N_14784,N_15030);
or U17224 (N_17224,N_14891,N_14302);
or U17225 (N_17225,N_14451,N_15950);
or U17226 (N_17226,N_15609,N_14755);
or U17227 (N_17227,N_14901,N_15000);
xor U17228 (N_17228,N_15442,N_14980);
or U17229 (N_17229,N_14398,N_15425);
nand U17230 (N_17230,N_14030,N_15839);
and U17231 (N_17231,N_15482,N_14339);
and U17232 (N_17232,N_15282,N_14549);
nand U17233 (N_17233,N_14334,N_14469);
nand U17234 (N_17234,N_14626,N_14007);
or U17235 (N_17235,N_15674,N_15084);
nor U17236 (N_17236,N_14473,N_14344);
nor U17237 (N_17237,N_15398,N_14241);
nor U17238 (N_17238,N_15555,N_15209);
or U17239 (N_17239,N_14300,N_15905);
and U17240 (N_17240,N_14682,N_15722);
nor U17241 (N_17241,N_14672,N_15751);
nand U17242 (N_17242,N_15406,N_14208);
or U17243 (N_17243,N_14914,N_15822);
nor U17244 (N_17244,N_14887,N_14436);
or U17245 (N_17245,N_15818,N_14236);
or U17246 (N_17246,N_15082,N_14907);
nand U17247 (N_17247,N_15831,N_15770);
or U17248 (N_17248,N_14657,N_14932);
and U17249 (N_17249,N_14463,N_15517);
or U17250 (N_17250,N_14213,N_14483);
nor U17251 (N_17251,N_14296,N_15110);
nand U17252 (N_17252,N_14414,N_15476);
xnor U17253 (N_17253,N_15059,N_14161);
or U17254 (N_17254,N_14932,N_14461);
or U17255 (N_17255,N_15503,N_15833);
or U17256 (N_17256,N_15738,N_14457);
and U17257 (N_17257,N_14603,N_14818);
nor U17258 (N_17258,N_15707,N_14850);
nor U17259 (N_17259,N_15882,N_14128);
xor U17260 (N_17260,N_14964,N_15192);
or U17261 (N_17261,N_15260,N_14838);
xnor U17262 (N_17262,N_15035,N_15911);
nand U17263 (N_17263,N_15181,N_15739);
xor U17264 (N_17264,N_14319,N_15035);
nand U17265 (N_17265,N_15603,N_15231);
xnor U17266 (N_17266,N_15538,N_15238);
nand U17267 (N_17267,N_15545,N_14107);
and U17268 (N_17268,N_14428,N_14698);
and U17269 (N_17269,N_14683,N_15308);
or U17270 (N_17270,N_15293,N_14987);
nor U17271 (N_17271,N_14300,N_14404);
xnor U17272 (N_17272,N_15409,N_15281);
or U17273 (N_17273,N_14181,N_15542);
or U17274 (N_17274,N_14234,N_14461);
or U17275 (N_17275,N_14059,N_15354);
nand U17276 (N_17276,N_15036,N_14888);
and U17277 (N_17277,N_15206,N_14440);
and U17278 (N_17278,N_15770,N_15342);
nor U17279 (N_17279,N_15260,N_15213);
xor U17280 (N_17280,N_14626,N_15861);
nor U17281 (N_17281,N_14125,N_15873);
nor U17282 (N_17282,N_14313,N_14125);
or U17283 (N_17283,N_14004,N_15839);
nor U17284 (N_17284,N_15958,N_14227);
xor U17285 (N_17285,N_14044,N_14069);
nor U17286 (N_17286,N_15077,N_15779);
nor U17287 (N_17287,N_14959,N_14089);
xor U17288 (N_17288,N_14096,N_15520);
nor U17289 (N_17289,N_14216,N_14443);
nor U17290 (N_17290,N_14955,N_15496);
nand U17291 (N_17291,N_14471,N_14608);
nand U17292 (N_17292,N_14465,N_15316);
and U17293 (N_17293,N_14532,N_15633);
or U17294 (N_17294,N_14479,N_14671);
nand U17295 (N_17295,N_14581,N_14175);
xor U17296 (N_17296,N_14063,N_14738);
nand U17297 (N_17297,N_14182,N_14813);
xnor U17298 (N_17298,N_15910,N_14368);
nand U17299 (N_17299,N_14913,N_14592);
nand U17300 (N_17300,N_14769,N_15737);
xor U17301 (N_17301,N_14719,N_15378);
nor U17302 (N_17302,N_14074,N_14292);
and U17303 (N_17303,N_15180,N_14687);
xnor U17304 (N_17304,N_15094,N_14631);
nor U17305 (N_17305,N_14013,N_15748);
nor U17306 (N_17306,N_15226,N_15560);
nor U17307 (N_17307,N_14711,N_14050);
or U17308 (N_17308,N_15722,N_15061);
xnor U17309 (N_17309,N_15016,N_15912);
nand U17310 (N_17310,N_15308,N_15355);
xnor U17311 (N_17311,N_15785,N_14288);
and U17312 (N_17312,N_15102,N_15254);
nand U17313 (N_17313,N_14919,N_15647);
nor U17314 (N_17314,N_14855,N_15881);
nand U17315 (N_17315,N_14529,N_15660);
nor U17316 (N_17316,N_15137,N_15086);
nand U17317 (N_17317,N_15792,N_15876);
xnor U17318 (N_17318,N_15137,N_15028);
or U17319 (N_17319,N_15152,N_15406);
and U17320 (N_17320,N_15182,N_14309);
or U17321 (N_17321,N_14054,N_15225);
nand U17322 (N_17322,N_15170,N_15601);
xnor U17323 (N_17323,N_15097,N_15801);
nand U17324 (N_17324,N_14291,N_14895);
xor U17325 (N_17325,N_15674,N_15282);
or U17326 (N_17326,N_15667,N_14129);
xnor U17327 (N_17327,N_14536,N_15425);
or U17328 (N_17328,N_15869,N_15191);
xnor U17329 (N_17329,N_14472,N_14331);
or U17330 (N_17330,N_14502,N_14346);
nor U17331 (N_17331,N_15648,N_14271);
xor U17332 (N_17332,N_15341,N_15306);
nand U17333 (N_17333,N_14894,N_14255);
and U17334 (N_17334,N_14556,N_14478);
xor U17335 (N_17335,N_14060,N_15934);
nand U17336 (N_17336,N_14275,N_15077);
xor U17337 (N_17337,N_14657,N_14732);
or U17338 (N_17338,N_14252,N_14080);
or U17339 (N_17339,N_15805,N_15535);
and U17340 (N_17340,N_14732,N_14010);
xnor U17341 (N_17341,N_15980,N_14371);
and U17342 (N_17342,N_15497,N_15352);
nor U17343 (N_17343,N_14001,N_14164);
nand U17344 (N_17344,N_14062,N_14822);
or U17345 (N_17345,N_14559,N_15134);
and U17346 (N_17346,N_15272,N_14977);
xnor U17347 (N_17347,N_15487,N_15793);
and U17348 (N_17348,N_15412,N_14913);
or U17349 (N_17349,N_15665,N_15872);
nand U17350 (N_17350,N_14353,N_14588);
and U17351 (N_17351,N_14395,N_14871);
nor U17352 (N_17352,N_15433,N_15941);
xnor U17353 (N_17353,N_15690,N_15040);
or U17354 (N_17354,N_14425,N_15686);
nor U17355 (N_17355,N_14082,N_15784);
nor U17356 (N_17356,N_15093,N_15097);
or U17357 (N_17357,N_15989,N_15118);
nand U17358 (N_17358,N_14422,N_15468);
and U17359 (N_17359,N_15255,N_14557);
and U17360 (N_17360,N_15376,N_14576);
nand U17361 (N_17361,N_14148,N_15171);
nand U17362 (N_17362,N_14208,N_15980);
nand U17363 (N_17363,N_14948,N_15170);
xor U17364 (N_17364,N_14569,N_15436);
nand U17365 (N_17365,N_15837,N_15465);
xor U17366 (N_17366,N_14041,N_14364);
nand U17367 (N_17367,N_14070,N_15268);
nor U17368 (N_17368,N_15883,N_15564);
xnor U17369 (N_17369,N_14956,N_14078);
nor U17370 (N_17370,N_15440,N_14229);
or U17371 (N_17371,N_14846,N_14704);
xor U17372 (N_17372,N_14944,N_14437);
nand U17373 (N_17373,N_15678,N_14024);
and U17374 (N_17374,N_15005,N_14679);
xnor U17375 (N_17375,N_14452,N_14436);
xnor U17376 (N_17376,N_15449,N_14594);
or U17377 (N_17377,N_15661,N_15335);
nand U17378 (N_17378,N_15289,N_15497);
or U17379 (N_17379,N_15024,N_14860);
nor U17380 (N_17380,N_15357,N_15747);
xnor U17381 (N_17381,N_15146,N_14067);
nand U17382 (N_17382,N_15110,N_15821);
or U17383 (N_17383,N_14494,N_15122);
xnor U17384 (N_17384,N_14758,N_15445);
nor U17385 (N_17385,N_15966,N_15217);
xor U17386 (N_17386,N_14294,N_14982);
or U17387 (N_17387,N_15096,N_15215);
and U17388 (N_17388,N_15894,N_14553);
nand U17389 (N_17389,N_14599,N_14443);
xnor U17390 (N_17390,N_15125,N_14191);
nor U17391 (N_17391,N_14810,N_14998);
or U17392 (N_17392,N_15343,N_14359);
or U17393 (N_17393,N_14983,N_14908);
nor U17394 (N_17394,N_15215,N_15406);
and U17395 (N_17395,N_14867,N_14513);
nor U17396 (N_17396,N_14337,N_15784);
nor U17397 (N_17397,N_15357,N_15460);
and U17398 (N_17398,N_15911,N_15793);
nor U17399 (N_17399,N_15221,N_15383);
or U17400 (N_17400,N_15638,N_14901);
xnor U17401 (N_17401,N_15513,N_15082);
xor U17402 (N_17402,N_15645,N_15793);
or U17403 (N_17403,N_15203,N_15093);
xnor U17404 (N_17404,N_15625,N_15611);
nand U17405 (N_17405,N_15998,N_14715);
or U17406 (N_17406,N_15004,N_14967);
or U17407 (N_17407,N_14392,N_15994);
xor U17408 (N_17408,N_14373,N_15612);
and U17409 (N_17409,N_15771,N_15872);
nor U17410 (N_17410,N_15550,N_14474);
nor U17411 (N_17411,N_15640,N_15894);
xor U17412 (N_17412,N_14401,N_14676);
xor U17413 (N_17413,N_15008,N_14466);
nor U17414 (N_17414,N_14098,N_15465);
xnor U17415 (N_17415,N_14282,N_15649);
and U17416 (N_17416,N_15157,N_15545);
and U17417 (N_17417,N_15612,N_15153);
or U17418 (N_17418,N_14722,N_15647);
nor U17419 (N_17419,N_14769,N_14673);
nor U17420 (N_17420,N_15200,N_15535);
or U17421 (N_17421,N_15407,N_14781);
nand U17422 (N_17422,N_15052,N_14923);
or U17423 (N_17423,N_14482,N_14940);
and U17424 (N_17424,N_15922,N_14114);
and U17425 (N_17425,N_14251,N_15864);
xor U17426 (N_17426,N_15256,N_14321);
nor U17427 (N_17427,N_14302,N_14564);
nand U17428 (N_17428,N_14587,N_15118);
nor U17429 (N_17429,N_15193,N_15230);
nand U17430 (N_17430,N_15588,N_15994);
or U17431 (N_17431,N_15396,N_14745);
or U17432 (N_17432,N_15799,N_15046);
nor U17433 (N_17433,N_15855,N_15312);
nand U17434 (N_17434,N_15849,N_14370);
and U17435 (N_17435,N_15069,N_14751);
xor U17436 (N_17436,N_15147,N_15771);
and U17437 (N_17437,N_14652,N_14927);
nor U17438 (N_17438,N_14562,N_14954);
and U17439 (N_17439,N_15256,N_15479);
nand U17440 (N_17440,N_15471,N_15120);
and U17441 (N_17441,N_15467,N_15374);
nand U17442 (N_17442,N_14715,N_14821);
nand U17443 (N_17443,N_14156,N_15781);
or U17444 (N_17444,N_14608,N_14235);
and U17445 (N_17445,N_15797,N_14955);
and U17446 (N_17446,N_15544,N_15972);
or U17447 (N_17447,N_14287,N_15694);
nor U17448 (N_17448,N_15536,N_15027);
nand U17449 (N_17449,N_14378,N_15408);
nor U17450 (N_17450,N_15573,N_15921);
or U17451 (N_17451,N_14480,N_14384);
nand U17452 (N_17452,N_14220,N_14244);
nor U17453 (N_17453,N_15504,N_15934);
or U17454 (N_17454,N_15284,N_14538);
nor U17455 (N_17455,N_15597,N_14083);
and U17456 (N_17456,N_14392,N_14090);
xor U17457 (N_17457,N_15548,N_14118);
xor U17458 (N_17458,N_15442,N_15642);
and U17459 (N_17459,N_14863,N_14053);
xnor U17460 (N_17460,N_15031,N_14545);
and U17461 (N_17461,N_14898,N_14081);
and U17462 (N_17462,N_14051,N_15702);
nor U17463 (N_17463,N_15849,N_14214);
nor U17464 (N_17464,N_15125,N_15405);
or U17465 (N_17465,N_14906,N_15749);
or U17466 (N_17466,N_15975,N_14978);
nor U17467 (N_17467,N_15264,N_14430);
nor U17468 (N_17468,N_15334,N_14225);
and U17469 (N_17469,N_14599,N_15498);
xnor U17470 (N_17470,N_14270,N_14028);
nor U17471 (N_17471,N_15715,N_15562);
nand U17472 (N_17472,N_14357,N_15129);
and U17473 (N_17473,N_14797,N_15953);
nand U17474 (N_17474,N_15165,N_15538);
xnor U17475 (N_17475,N_14961,N_15347);
nand U17476 (N_17476,N_14227,N_14110);
or U17477 (N_17477,N_14061,N_15563);
nor U17478 (N_17478,N_15714,N_14030);
nor U17479 (N_17479,N_15409,N_15825);
or U17480 (N_17480,N_15643,N_14387);
nand U17481 (N_17481,N_15080,N_15682);
nor U17482 (N_17482,N_14678,N_15518);
nor U17483 (N_17483,N_14349,N_15439);
and U17484 (N_17484,N_15459,N_14295);
nand U17485 (N_17485,N_15599,N_14058);
nand U17486 (N_17486,N_14348,N_14661);
and U17487 (N_17487,N_15677,N_15168);
and U17488 (N_17488,N_15788,N_15685);
and U17489 (N_17489,N_15214,N_15239);
or U17490 (N_17490,N_15246,N_14805);
and U17491 (N_17491,N_15943,N_14897);
and U17492 (N_17492,N_15792,N_14742);
nor U17493 (N_17493,N_14313,N_14575);
or U17494 (N_17494,N_14097,N_14898);
nand U17495 (N_17495,N_14018,N_14183);
nor U17496 (N_17496,N_14887,N_15550);
or U17497 (N_17497,N_14509,N_14113);
nand U17498 (N_17498,N_14239,N_15684);
and U17499 (N_17499,N_15572,N_15271);
or U17500 (N_17500,N_14579,N_15714);
nand U17501 (N_17501,N_15774,N_14735);
or U17502 (N_17502,N_14464,N_14798);
and U17503 (N_17503,N_15774,N_14322);
or U17504 (N_17504,N_14761,N_14701);
or U17505 (N_17505,N_14883,N_15345);
or U17506 (N_17506,N_15921,N_15344);
and U17507 (N_17507,N_14390,N_14210);
xor U17508 (N_17508,N_14140,N_15198);
and U17509 (N_17509,N_14343,N_15877);
nand U17510 (N_17510,N_15970,N_14777);
and U17511 (N_17511,N_15157,N_14508);
xnor U17512 (N_17512,N_14941,N_14145);
xnor U17513 (N_17513,N_14999,N_15850);
nand U17514 (N_17514,N_14373,N_15210);
nor U17515 (N_17515,N_14021,N_14831);
or U17516 (N_17516,N_15190,N_14548);
or U17517 (N_17517,N_14727,N_15191);
xor U17518 (N_17518,N_14381,N_15856);
or U17519 (N_17519,N_14929,N_14896);
and U17520 (N_17520,N_15917,N_15200);
nor U17521 (N_17521,N_14252,N_15622);
and U17522 (N_17522,N_15872,N_15987);
and U17523 (N_17523,N_15962,N_15947);
xor U17524 (N_17524,N_15577,N_15262);
nor U17525 (N_17525,N_15843,N_14748);
nand U17526 (N_17526,N_14233,N_15086);
nand U17527 (N_17527,N_15586,N_14621);
or U17528 (N_17528,N_15436,N_14783);
or U17529 (N_17529,N_14583,N_14370);
xor U17530 (N_17530,N_15363,N_15595);
nor U17531 (N_17531,N_15350,N_14489);
nand U17532 (N_17532,N_15378,N_14370);
or U17533 (N_17533,N_14352,N_14555);
xor U17534 (N_17534,N_14744,N_15100);
or U17535 (N_17535,N_14555,N_15285);
xnor U17536 (N_17536,N_15661,N_15365);
or U17537 (N_17537,N_15312,N_14935);
nand U17538 (N_17538,N_15560,N_15322);
nor U17539 (N_17539,N_14369,N_14419);
nor U17540 (N_17540,N_14148,N_14283);
or U17541 (N_17541,N_14487,N_15115);
nor U17542 (N_17542,N_14974,N_15990);
nand U17543 (N_17543,N_15572,N_15479);
nand U17544 (N_17544,N_14605,N_15145);
or U17545 (N_17545,N_15121,N_14216);
xnor U17546 (N_17546,N_14013,N_14363);
nor U17547 (N_17547,N_14312,N_14263);
nor U17548 (N_17548,N_14445,N_15527);
or U17549 (N_17549,N_14090,N_14205);
nand U17550 (N_17550,N_15013,N_14097);
or U17551 (N_17551,N_14844,N_14482);
nor U17552 (N_17552,N_14983,N_14014);
or U17553 (N_17553,N_15827,N_14072);
nand U17554 (N_17554,N_14569,N_14014);
nor U17555 (N_17555,N_15400,N_15317);
xor U17556 (N_17556,N_15694,N_14256);
nand U17557 (N_17557,N_14811,N_14575);
and U17558 (N_17558,N_14213,N_15077);
nor U17559 (N_17559,N_14999,N_15969);
and U17560 (N_17560,N_15258,N_14785);
and U17561 (N_17561,N_14458,N_14644);
nand U17562 (N_17562,N_14968,N_14469);
nor U17563 (N_17563,N_15508,N_14540);
nand U17564 (N_17564,N_14306,N_15009);
nand U17565 (N_17565,N_15568,N_15818);
xor U17566 (N_17566,N_14357,N_14691);
nor U17567 (N_17567,N_15722,N_14574);
and U17568 (N_17568,N_15025,N_15634);
or U17569 (N_17569,N_15952,N_14480);
xnor U17570 (N_17570,N_14658,N_15588);
and U17571 (N_17571,N_14290,N_14447);
or U17572 (N_17572,N_15205,N_14052);
nand U17573 (N_17573,N_15407,N_14965);
or U17574 (N_17574,N_15270,N_15941);
nor U17575 (N_17575,N_14805,N_14441);
nand U17576 (N_17576,N_15023,N_14661);
xnor U17577 (N_17577,N_14597,N_15433);
or U17578 (N_17578,N_15293,N_14462);
and U17579 (N_17579,N_14156,N_15956);
nand U17580 (N_17580,N_15406,N_15662);
and U17581 (N_17581,N_14687,N_15657);
nand U17582 (N_17582,N_15922,N_15513);
nand U17583 (N_17583,N_14428,N_14806);
or U17584 (N_17584,N_14231,N_15107);
xor U17585 (N_17585,N_15446,N_14939);
xnor U17586 (N_17586,N_15026,N_15563);
nor U17587 (N_17587,N_15422,N_15299);
and U17588 (N_17588,N_14569,N_14784);
and U17589 (N_17589,N_14248,N_14928);
or U17590 (N_17590,N_14863,N_14260);
nor U17591 (N_17591,N_15064,N_15385);
nor U17592 (N_17592,N_15657,N_14481);
nand U17593 (N_17593,N_15350,N_15563);
nor U17594 (N_17594,N_15823,N_14610);
nand U17595 (N_17595,N_15707,N_14785);
xnor U17596 (N_17596,N_14075,N_15900);
nand U17597 (N_17597,N_15951,N_15515);
nand U17598 (N_17598,N_14898,N_15291);
nand U17599 (N_17599,N_14301,N_14473);
nand U17600 (N_17600,N_14171,N_14210);
or U17601 (N_17601,N_15403,N_15935);
or U17602 (N_17602,N_15728,N_15464);
and U17603 (N_17603,N_15875,N_15462);
xnor U17604 (N_17604,N_14729,N_15776);
nand U17605 (N_17605,N_14262,N_15412);
xnor U17606 (N_17606,N_14278,N_14375);
nand U17607 (N_17607,N_14719,N_15153);
nor U17608 (N_17608,N_15407,N_14287);
xnor U17609 (N_17609,N_14017,N_14978);
and U17610 (N_17610,N_15356,N_15606);
xnor U17611 (N_17611,N_15786,N_14343);
xnor U17612 (N_17612,N_15533,N_14687);
xor U17613 (N_17613,N_14965,N_15690);
and U17614 (N_17614,N_14402,N_14416);
or U17615 (N_17615,N_15768,N_15027);
nor U17616 (N_17616,N_14539,N_15794);
and U17617 (N_17617,N_15723,N_14675);
nand U17618 (N_17618,N_15194,N_14732);
or U17619 (N_17619,N_14336,N_14727);
nor U17620 (N_17620,N_15321,N_14525);
and U17621 (N_17621,N_15066,N_14224);
or U17622 (N_17622,N_15363,N_14641);
or U17623 (N_17623,N_14677,N_15301);
and U17624 (N_17624,N_15008,N_14585);
nand U17625 (N_17625,N_14698,N_15465);
xor U17626 (N_17626,N_15004,N_15443);
or U17627 (N_17627,N_14223,N_15828);
or U17628 (N_17628,N_15384,N_15361);
nand U17629 (N_17629,N_14371,N_15831);
nand U17630 (N_17630,N_14468,N_14244);
or U17631 (N_17631,N_14617,N_14946);
nand U17632 (N_17632,N_15392,N_15015);
nor U17633 (N_17633,N_15580,N_14224);
or U17634 (N_17634,N_15475,N_14502);
nor U17635 (N_17635,N_15765,N_15311);
nor U17636 (N_17636,N_15256,N_15963);
xor U17637 (N_17637,N_14825,N_14139);
or U17638 (N_17638,N_14749,N_14926);
nand U17639 (N_17639,N_14254,N_14372);
xor U17640 (N_17640,N_14059,N_14819);
nor U17641 (N_17641,N_15310,N_15320);
xor U17642 (N_17642,N_14016,N_15516);
xor U17643 (N_17643,N_14803,N_15959);
and U17644 (N_17644,N_15898,N_15428);
nand U17645 (N_17645,N_15514,N_15452);
or U17646 (N_17646,N_15279,N_15728);
and U17647 (N_17647,N_14873,N_15903);
or U17648 (N_17648,N_15441,N_15990);
nand U17649 (N_17649,N_15098,N_15855);
or U17650 (N_17650,N_14665,N_15308);
nand U17651 (N_17651,N_14743,N_14863);
nor U17652 (N_17652,N_15957,N_14282);
xor U17653 (N_17653,N_15852,N_15572);
nand U17654 (N_17654,N_15740,N_14443);
xor U17655 (N_17655,N_15184,N_14124);
or U17656 (N_17656,N_14665,N_15670);
and U17657 (N_17657,N_14883,N_15468);
and U17658 (N_17658,N_14075,N_14370);
nor U17659 (N_17659,N_15837,N_15963);
or U17660 (N_17660,N_14317,N_15183);
nand U17661 (N_17661,N_15586,N_15993);
or U17662 (N_17662,N_15419,N_14996);
xor U17663 (N_17663,N_15071,N_14760);
and U17664 (N_17664,N_15837,N_15189);
xnor U17665 (N_17665,N_15599,N_15091);
nor U17666 (N_17666,N_15661,N_15142);
xor U17667 (N_17667,N_15181,N_15389);
xnor U17668 (N_17668,N_15205,N_14988);
or U17669 (N_17669,N_14371,N_15915);
and U17670 (N_17670,N_14355,N_15650);
or U17671 (N_17671,N_14482,N_14825);
and U17672 (N_17672,N_15418,N_15285);
nand U17673 (N_17673,N_14320,N_15261);
xor U17674 (N_17674,N_14411,N_15923);
and U17675 (N_17675,N_15094,N_14011);
nor U17676 (N_17676,N_15345,N_15870);
xor U17677 (N_17677,N_15919,N_14864);
nor U17678 (N_17678,N_14976,N_15238);
nor U17679 (N_17679,N_15277,N_15087);
and U17680 (N_17680,N_14049,N_14001);
and U17681 (N_17681,N_15345,N_14522);
or U17682 (N_17682,N_14108,N_15205);
nor U17683 (N_17683,N_14883,N_15651);
or U17684 (N_17684,N_15998,N_14489);
nand U17685 (N_17685,N_15820,N_14684);
and U17686 (N_17686,N_15988,N_15602);
nor U17687 (N_17687,N_14233,N_14621);
nor U17688 (N_17688,N_14859,N_14156);
and U17689 (N_17689,N_14738,N_14818);
xor U17690 (N_17690,N_15493,N_15712);
nand U17691 (N_17691,N_14378,N_14324);
and U17692 (N_17692,N_14065,N_14865);
xor U17693 (N_17693,N_14443,N_14025);
xnor U17694 (N_17694,N_14132,N_15677);
xnor U17695 (N_17695,N_14837,N_15952);
and U17696 (N_17696,N_15743,N_15175);
xnor U17697 (N_17697,N_14008,N_14944);
nand U17698 (N_17698,N_14200,N_14400);
xnor U17699 (N_17699,N_14539,N_14019);
nor U17700 (N_17700,N_14013,N_15361);
nor U17701 (N_17701,N_14296,N_15688);
nor U17702 (N_17702,N_15396,N_14111);
and U17703 (N_17703,N_15932,N_14454);
xor U17704 (N_17704,N_15095,N_14031);
or U17705 (N_17705,N_15636,N_14985);
nand U17706 (N_17706,N_15393,N_15270);
nor U17707 (N_17707,N_14471,N_15771);
or U17708 (N_17708,N_15531,N_14902);
nand U17709 (N_17709,N_15953,N_15566);
nor U17710 (N_17710,N_14669,N_15631);
nand U17711 (N_17711,N_14335,N_15195);
nor U17712 (N_17712,N_15802,N_15166);
xnor U17713 (N_17713,N_14433,N_15019);
nor U17714 (N_17714,N_15347,N_14900);
and U17715 (N_17715,N_15555,N_14466);
and U17716 (N_17716,N_14818,N_15033);
nand U17717 (N_17717,N_15287,N_15047);
xnor U17718 (N_17718,N_15405,N_15379);
nand U17719 (N_17719,N_14015,N_14649);
and U17720 (N_17720,N_14221,N_14747);
and U17721 (N_17721,N_14454,N_15465);
and U17722 (N_17722,N_15067,N_14773);
or U17723 (N_17723,N_14847,N_14257);
or U17724 (N_17724,N_15062,N_14724);
and U17725 (N_17725,N_15988,N_15725);
or U17726 (N_17726,N_15435,N_15922);
nand U17727 (N_17727,N_15206,N_14296);
and U17728 (N_17728,N_15508,N_14207);
and U17729 (N_17729,N_15311,N_15460);
and U17730 (N_17730,N_15602,N_14425);
xor U17731 (N_17731,N_15162,N_15965);
nor U17732 (N_17732,N_15874,N_14256);
nor U17733 (N_17733,N_15923,N_14149);
nand U17734 (N_17734,N_15720,N_15410);
nand U17735 (N_17735,N_14636,N_14130);
or U17736 (N_17736,N_15947,N_14838);
nor U17737 (N_17737,N_14652,N_14502);
nand U17738 (N_17738,N_14497,N_14938);
or U17739 (N_17739,N_14857,N_15117);
or U17740 (N_17740,N_14755,N_14789);
nand U17741 (N_17741,N_14854,N_14549);
nand U17742 (N_17742,N_14469,N_14093);
xnor U17743 (N_17743,N_14686,N_15401);
nand U17744 (N_17744,N_14734,N_14573);
nor U17745 (N_17745,N_14961,N_14126);
or U17746 (N_17746,N_15521,N_15341);
nor U17747 (N_17747,N_14326,N_15716);
nand U17748 (N_17748,N_14429,N_14620);
nand U17749 (N_17749,N_15985,N_14807);
and U17750 (N_17750,N_14409,N_15675);
xor U17751 (N_17751,N_15296,N_14860);
nor U17752 (N_17752,N_14871,N_14553);
and U17753 (N_17753,N_14929,N_14753);
nand U17754 (N_17754,N_14025,N_14373);
and U17755 (N_17755,N_15945,N_15736);
or U17756 (N_17756,N_14165,N_15205);
and U17757 (N_17757,N_15223,N_14230);
nor U17758 (N_17758,N_15619,N_15336);
nor U17759 (N_17759,N_14662,N_15470);
and U17760 (N_17760,N_15495,N_15641);
nand U17761 (N_17761,N_15712,N_14813);
and U17762 (N_17762,N_14384,N_15137);
nor U17763 (N_17763,N_14335,N_15869);
nand U17764 (N_17764,N_15623,N_15984);
and U17765 (N_17765,N_14878,N_14999);
nor U17766 (N_17766,N_15720,N_14220);
xnor U17767 (N_17767,N_15307,N_15395);
nand U17768 (N_17768,N_14783,N_15079);
nand U17769 (N_17769,N_15154,N_15642);
nand U17770 (N_17770,N_14218,N_14567);
xor U17771 (N_17771,N_15479,N_15835);
nand U17772 (N_17772,N_14588,N_15565);
xor U17773 (N_17773,N_14511,N_14858);
xnor U17774 (N_17774,N_14029,N_14317);
nor U17775 (N_17775,N_15427,N_15452);
or U17776 (N_17776,N_14712,N_14592);
and U17777 (N_17777,N_14313,N_14470);
or U17778 (N_17778,N_14405,N_14656);
and U17779 (N_17779,N_15462,N_14368);
nand U17780 (N_17780,N_14828,N_15168);
nand U17781 (N_17781,N_15234,N_14439);
nand U17782 (N_17782,N_14393,N_14189);
or U17783 (N_17783,N_15214,N_14432);
or U17784 (N_17784,N_15217,N_14871);
nand U17785 (N_17785,N_14188,N_14490);
nand U17786 (N_17786,N_15775,N_14026);
and U17787 (N_17787,N_14084,N_15614);
xnor U17788 (N_17788,N_15802,N_15897);
xor U17789 (N_17789,N_15926,N_15485);
and U17790 (N_17790,N_15279,N_14301);
and U17791 (N_17791,N_15918,N_15037);
nand U17792 (N_17792,N_14764,N_14316);
xnor U17793 (N_17793,N_14397,N_14063);
and U17794 (N_17794,N_15869,N_14345);
or U17795 (N_17795,N_15353,N_14030);
xor U17796 (N_17796,N_14438,N_15531);
and U17797 (N_17797,N_15832,N_14190);
nand U17798 (N_17798,N_15047,N_14686);
nor U17799 (N_17799,N_15761,N_14677);
xor U17800 (N_17800,N_15196,N_14343);
and U17801 (N_17801,N_15219,N_14937);
xnor U17802 (N_17802,N_14481,N_15745);
and U17803 (N_17803,N_15468,N_15091);
or U17804 (N_17804,N_14622,N_15393);
or U17805 (N_17805,N_15609,N_14050);
nor U17806 (N_17806,N_14405,N_14062);
nand U17807 (N_17807,N_15567,N_14858);
nand U17808 (N_17808,N_14419,N_15622);
nor U17809 (N_17809,N_14935,N_14310);
nand U17810 (N_17810,N_14830,N_15080);
or U17811 (N_17811,N_15803,N_15430);
nand U17812 (N_17812,N_15393,N_14574);
nor U17813 (N_17813,N_14319,N_15657);
nand U17814 (N_17814,N_14268,N_14701);
nor U17815 (N_17815,N_15842,N_14889);
or U17816 (N_17816,N_15881,N_14175);
or U17817 (N_17817,N_14317,N_14955);
or U17818 (N_17818,N_14881,N_15615);
and U17819 (N_17819,N_15674,N_14271);
nand U17820 (N_17820,N_14121,N_15289);
or U17821 (N_17821,N_14049,N_15633);
xor U17822 (N_17822,N_15288,N_15225);
nor U17823 (N_17823,N_14335,N_15225);
and U17824 (N_17824,N_15692,N_14624);
xor U17825 (N_17825,N_14968,N_14293);
nand U17826 (N_17826,N_14105,N_14630);
nor U17827 (N_17827,N_14780,N_14223);
and U17828 (N_17828,N_14888,N_14909);
or U17829 (N_17829,N_14126,N_15928);
nand U17830 (N_17830,N_14298,N_15982);
nor U17831 (N_17831,N_15384,N_14229);
nand U17832 (N_17832,N_15119,N_15552);
and U17833 (N_17833,N_14899,N_14678);
nor U17834 (N_17834,N_14420,N_15904);
or U17835 (N_17835,N_14873,N_15498);
nor U17836 (N_17836,N_15938,N_14544);
xor U17837 (N_17837,N_15003,N_14400);
or U17838 (N_17838,N_14110,N_14178);
nand U17839 (N_17839,N_15049,N_15370);
nor U17840 (N_17840,N_15678,N_15054);
xor U17841 (N_17841,N_15466,N_14777);
and U17842 (N_17842,N_14540,N_15716);
xnor U17843 (N_17843,N_15266,N_14859);
and U17844 (N_17844,N_15967,N_15410);
xor U17845 (N_17845,N_15588,N_15922);
xor U17846 (N_17846,N_14031,N_14499);
xnor U17847 (N_17847,N_15807,N_15065);
xor U17848 (N_17848,N_15439,N_15019);
xnor U17849 (N_17849,N_15794,N_14637);
nor U17850 (N_17850,N_14787,N_14512);
or U17851 (N_17851,N_14100,N_14270);
and U17852 (N_17852,N_15672,N_14331);
xor U17853 (N_17853,N_15118,N_14379);
xnor U17854 (N_17854,N_15334,N_15811);
nor U17855 (N_17855,N_14794,N_14300);
nand U17856 (N_17856,N_14741,N_15628);
nand U17857 (N_17857,N_14990,N_14302);
nand U17858 (N_17858,N_14525,N_14713);
and U17859 (N_17859,N_15945,N_15345);
xnor U17860 (N_17860,N_14149,N_14249);
nand U17861 (N_17861,N_14384,N_14323);
nand U17862 (N_17862,N_14845,N_15689);
nand U17863 (N_17863,N_14980,N_15016);
nor U17864 (N_17864,N_14451,N_15801);
and U17865 (N_17865,N_15672,N_15069);
nand U17866 (N_17866,N_14208,N_14137);
xnor U17867 (N_17867,N_14463,N_14890);
xor U17868 (N_17868,N_14188,N_14645);
or U17869 (N_17869,N_15496,N_14302);
nor U17870 (N_17870,N_15044,N_14164);
and U17871 (N_17871,N_15075,N_14801);
and U17872 (N_17872,N_14221,N_15562);
nor U17873 (N_17873,N_15818,N_15193);
xnor U17874 (N_17874,N_15982,N_15113);
nor U17875 (N_17875,N_15329,N_14031);
xnor U17876 (N_17876,N_15942,N_14824);
nor U17877 (N_17877,N_14203,N_14002);
nand U17878 (N_17878,N_14127,N_14899);
nor U17879 (N_17879,N_14315,N_14537);
nor U17880 (N_17880,N_15448,N_15377);
or U17881 (N_17881,N_15809,N_15813);
xnor U17882 (N_17882,N_14302,N_15397);
and U17883 (N_17883,N_14101,N_14999);
nor U17884 (N_17884,N_15757,N_15356);
and U17885 (N_17885,N_14513,N_14350);
xnor U17886 (N_17886,N_14333,N_15897);
nor U17887 (N_17887,N_14799,N_14454);
or U17888 (N_17888,N_15653,N_15549);
xnor U17889 (N_17889,N_15933,N_15942);
nor U17890 (N_17890,N_15290,N_15607);
and U17891 (N_17891,N_14163,N_15403);
and U17892 (N_17892,N_14303,N_14540);
nand U17893 (N_17893,N_15445,N_14169);
xor U17894 (N_17894,N_14266,N_15827);
xnor U17895 (N_17895,N_14913,N_15358);
or U17896 (N_17896,N_14996,N_15001);
xor U17897 (N_17897,N_14606,N_14005);
xor U17898 (N_17898,N_14895,N_15637);
nor U17899 (N_17899,N_15188,N_15897);
and U17900 (N_17900,N_14619,N_15300);
or U17901 (N_17901,N_15998,N_15281);
and U17902 (N_17902,N_15763,N_15613);
nor U17903 (N_17903,N_14376,N_14537);
and U17904 (N_17904,N_14867,N_14021);
nand U17905 (N_17905,N_15111,N_14558);
and U17906 (N_17906,N_15124,N_15921);
and U17907 (N_17907,N_15390,N_14913);
or U17908 (N_17908,N_15061,N_15431);
nand U17909 (N_17909,N_14900,N_14223);
and U17910 (N_17910,N_15562,N_14069);
or U17911 (N_17911,N_15192,N_14372);
nor U17912 (N_17912,N_15878,N_14380);
nor U17913 (N_17913,N_15594,N_15234);
xor U17914 (N_17914,N_14631,N_15448);
or U17915 (N_17915,N_14081,N_15444);
xnor U17916 (N_17916,N_15503,N_14497);
and U17917 (N_17917,N_14709,N_15207);
xor U17918 (N_17918,N_15901,N_15229);
and U17919 (N_17919,N_14561,N_15761);
nand U17920 (N_17920,N_15040,N_14019);
nor U17921 (N_17921,N_15070,N_15701);
and U17922 (N_17922,N_15317,N_14582);
or U17923 (N_17923,N_14021,N_14816);
nor U17924 (N_17924,N_15929,N_15669);
nor U17925 (N_17925,N_14878,N_14761);
xnor U17926 (N_17926,N_15026,N_15682);
nor U17927 (N_17927,N_15305,N_15780);
xor U17928 (N_17928,N_14364,N_15614);
or U17929 (N_17929,N_14946,N_15589);
or U17930 (N_17930,N_15937,N_14370);
and U17931 (N_17931,N_14327,N_14073);
xor U17932 (N_17932,N_14147,N_14557);
nor U17933 (N_17933,N_14183,N_15784);
and U17934 (N_17934,N_15866,N_15389);
nand U17935 (N_17935,N_14924,N_15420);
xor U17936 (N_17936,N_15228,N_14348);
nor U17937 (N_17937,N_14020,N_14544);
or U17938 (N_17938,N_15103,N_15123);
xor U17939 (N_17939,N_14243,N_14800);
and U17940 (N_17940,N_15553,N_14691);
and U17941 (N_17941,N_14906,N_15450);
nor U17942 (N_17942,N_14629,N_14996);
nor U17943 (N_17943,N_14076,N_15260);
nand U17944 (N_17944,N_15355,N_14329);
or U17945 (N_17945,N_15790,N_15044);
xor U17946 (N_17946,N_15490,N_14034);
nand U17947 (N_17947,N_14398,N_15350);
or U17948 (N_17948,N_15512,N_14753);
xnor U17949 (N_17949,N_14243,N_15375);
or U17950 (N_17950,N_14783,N_14098);
or U17951 (N_17951,N_14641,N_15478);
nor U17952 (N_17952,N_14900,N_15241);
and U17953 (N_17953,N_14071,N_14271);
nor U17954 (N_17954,N_15168,N_14293);
nor U17955 (N_17955,N_14383,N_15923);
nand U17956 (N_17956,N_15970,N_15850);
nand U17957 (N_17957,N_15686,N_15120);
nor U17958 (N_17958,N_14754,N_15792);
nor U17959 (N_17959,N_14799,N_15652);
nor U17960 (N_17960,N_14558,N_14377);
nor U17961 (N_17961,N_15214,N_14814);
or U17962 (N_17962,N_14756,N_15912);
nor U17963 (N_17963,N_15279,N_15942);
and U17964 (N_17964,N_15905,N_15331);
and U17965 (N_17965,N_15419,N_15581);
nand U17966 (N_17966,N_14043,N_14267);
xor U17967 (N_17967,N_14181,N_14837);
xnor U17968 (N_17968,N_14818,N_15326);
nand U17969 (N_17969,N_14364,N_14439);
and U17970 (N_17970,N_14224,N_14079);
nor U17971 (N_17971,N_15269,N_15299);
or U17972 (N_17972,N_15148,N_15489);
nor U17973 (N_17973,N_14923,N_15631);
nand U17974 (N_17974,N_15885,N_15819);
nand U17975 (N_17975,N_14053,N_15227);
nand U17976 (N_17976,N_15312,N_14708);
or U17977 (N_17977,N_14589,N_14926);
nand U17978 (N_17978,N_15392,N_15110);
nand U17979 (N_17979,N_14342,N_14389);
nand U17980 (N_17980,N_14011,N_15434);
xnor U17981 (N_17981,N_15130,N_15438);
nand U17982 (N_17982,N_15689,N_14611);
nand U17983 (N_17983,N_15807,N_15068);
nand U17984 (N_17984,N_14003,N_15602);
or U17985 (N_17985,N_14609,N_14048);
or U17986 (N_17986,N_15962,N_14753);
and U17987 (N_17987,N_15733,N_14778);
xnor U17988 (N_17988,N_14553,N_15344);
or U17989 (N_17989,N_15667,N_15731);
nor U17990 (N_17990,N_14406,N_15088);
nor U17991 (N_17991,N_14930,N_14826);
nor U17992 (N_17992,N_14530,N_14169);
and U17993 (N_17993,N_15969,N_15175);
xor U17994 (N_17994,N_14754,N_14300);
nand U17995 (N_17995,N_15561,N_15386);
or U17996 (N_17996,N_14343,N_15689);
and U17997 (N_17997,N_14483,N_14623);
nand U17998 (N_17998,N_14379,N_14863);
and U17999 (N_17999,N_15941,N_14680);
and U18000 (N_18000,N_16381,N_17281);
or U18001 (N_18001,N_17709,N_16675);
or U18002 (N_18002,N_16110,N_16292);
nand U18003 (N_18003,N_17371,N_17559);
or U18004 (N_18004,N_16620,N_16617);
nor U18005 (N_18005,N_17380,N_16266);
and U18006 (N_18006,N_16809,N_17913);
nor U18007 (N_18007,N_17126,N_16562);
or U18008 (N_18008,N_16155,N_16277);
or U18009 (N_18009,N_16184,N_16237);
nor U18010 (N_18010,N_16076,N_16670);
nor U18011 (N_18011,N_16442,N_17908);
and U18012 (N_18012,N_16386,N_17675);
xnor U18013 (N_18013,N_17677,N_17504);
nand U18014 (N_18014,N_16420,N_17160);
nor U18015 (N_18015,N_16048,N_17657);
or U18016 (N_18016,N_16471,N_16289);
nor U18017 (N_18017,N_17074,N_17343);
nand U18018 (N_18018,N_16642,N_17886);
nor U18019 (N_18019,N_16456,N_17631);
and U18020 (N_18020,N_17237,N_16521);
nand U18021 (N_18021,N_17876,N_16597);
nor U18022 (N_18022,N_17097,N_17098);
nor U18023 (N_18023,N_17427,N_16802);
or U18024 (N_18024,N_17331,N_16206);
and U18025 (N_18025,N_16777,N_16779);
and U18026 (N_18026,N_16689,N_17565);
and U18027 (N_18027,N_17770,N_17285);
nand U18028 (N_18028,N_17139,N_16919);
and U18029 (N_18029,N_16781,N_16963);
nand U18030 (N_18030,N_16115,N_16545);
nor U18031 (N_18031,N_16969,N_16105);
xnor U18032 (N_18032,N_17884,N_16201);
xor U18033 (N_18033,N_17907,N_17665);
xor U18034 (N_18034,N_16463,N_17533);
xor U18035 (N_18035,N_17662,N_16715);
and U18036 (N_18036,N_17635,N_16189);
nand U18037 (N_18037,N_17523,N_17661);
nor U18038 (N_18038,N_16871,N_17682);
nand U18039 (N_18039,N_16719,N_17834);
and U18040 (N_18040,N_17353,N_17349);
or U18041 (N_18041,N_16122,N_16044);
or U18042 (N_18042,N_16150,N_17958);
xnor U18043 (N_18043,N_17182,N_17712);
nor U18044 (N_18044,N_16223,N_16556);
xnor U18045 (N_18045,N_16068,N_17015);
and U18046 (N_18046,N_16198,N_16078);
or U18047 (N_18047,N_17987,N_16708);
xor U18048 (N_18048,N_17377,N_16868);
nand U18049 (N_18049,N_16859,N_17871);
nor U18050 (N_18050,N_17835,N_17455);
xor U18051 (N_18051,N_17899,N_17608);
nor U18052 (N_18052,N_16728,N_16692);
nand U18053 (N_18053,N_17018,N_16782);
and U18054 (N_18054,N_17280,N_16563);
xnor U18055 (N_18055,N_16994,N_17529);
and U18056 (N_18056,N_17252,N_16844);
nand U18057 (N_18057,N_16209,N_16747);
xnor U18058 (N_18058,N_17865,N_16548);
nor U18059 (N_18059,N_16441,N_16251);
nor U18060 (N_18060,N_17292,N_17558);
xor U18061 (N_18061,N_17761,N_16338);
or U18062 (N_18062,N_16482,N_16389);
and U18063 (N_18063,N_16773,N_16108);
nand U18064 (N_18064,N_17467,N_16928);
nor U18065 (N_18065,N_17989,N_16662);
or U18066 (N_18066,N_17440,N_17161);
nand U18067 (N_18067,N_16646,N_17214);
xor U18068 (N_18068,N_16653,N_16351);
xor U18069 (N_18069,N_17069,N_17232);
xnor U18070 (N_18070,N_17119,N_16930);
nor U18071 (N_18071,N_17025,N_16881);
or U18072 (N_18072,N_16981,N_17612);
nand U18073 (N_18073,N_17852,N_17058);
xnor U18074 (N_18074,N_17585,N_16605);
or U18075 (N_18075,N_17159,N_16286);
xor U18076 (N_18076,N_17000,N_17127);
nand U18077 (N_18077,N_16226,N_16603);
and U18078 (N_18078,N_17187,N_17451);
and U18079 (N_18079,N_17370,N_16834);
nor U18080 (N_18080,N_16967,N_17554);
or U18081 (N_18081,N_17295,N_16455);
or U18082 (N_18082,N_16271,N_17879);
nand U18083 (N_18083,N_16248,N_16912);
xnor U18084 (N_18084,N_16904,N_17954);
nand U18085 (N_18085,N_16474,N_17569);
and U18086 (N_18086,N_17937,N_16811);
nand U18087 (N_18087,N_16353,N_16537);
nand U18088 (N_18088,N_16768,N_16475);
nor U18089 (N_18089,N_17962,N_17385);
and U18090 (N_18090,N_17875,N_16958);
and U18091 (N_18091,N_17438,N_17499);
nor U18092 (N_18092,N_17108,N_17810);
or U18093 (N_18093,N_17430,N_17955);
nand U18094 (N_18094,N_17124,N_16991);
nand U18095 (N_18095,N_16683,N_16152);
and U18096 (N_18096,N_16660,N_17563);
nor U18097 (N_18097,N_17723,N_16872);
or U18098 (N_18098,N_16318,N_16090);
xor U18099 (N_18099,N_17616,N_16933);
nand U18100 (N_18100,N_17691,N_17624);
nor U18101 (N_18101,N_17898,N_16553);
xor U18102 (N_18102,N_17830,N_17656);
nor U18103 (N_18103,N_16832,N_16737);
xnor U18104 (N_18104,N_17923,N_16778);
nand U18105 (N_18105,N_16842,N_16060);
nor U18106 (N_18106,N_17114,N_17732);
nor U18107 (N_18107,N_17200,N_17809);
or U18108 (N_18108,N_16494,N_17382);
nand U18109 (N_18109,N_16697,N_16400);
and U18110 (N_18110,N_17916,N_17474);
and U18111 (N_18111,N_17950,N_17328);
or U18112 (N_18112,N_16913,N_17432);
xnor U18113 (N_18113,N_17547,N_17488);
and U18114 (N_18114,N_16036,N_17995);
and U18115 (N_18115,N_16310,N_16448);
nor U18116 (N_18116,N_17170,N_17526);
nand U18117 (N_18117,N_16245,N_16290);
or U18118 (N_18118,N_16512,N_16945);
or U18119 (N_18119,N_16821,N_17372);
nand U18120 (N_18120,N_17306,N_16899);
nor U18121 (N_18121,N_17673,N_17644);
and U18122 (N_18122,N_17329,N_16723);
nor U18123 (N_18123,N_16657,N_17457);
and U18124 (N_18124,N_17763,N_16473);
nand U18125 (N_18125,N_16439,N_17773);
or U18126 (N_18126,N_17755,N_17615);
and U18127 (N_18127,N_17494,N_16787);
nor U18128 (N_18128,N_17690,N_17535);
nand U18129 (N_18129,N_17775,N_16328);
nor U18130 (N_18130,N_17304,N_17699);
and U18131 (N_18131,N_17376,N_16129);
xor U18132 (N_18132,N_16917,N_17392);
or U18133 (N_18133,N_17931,N_16363);
xnor U18134 (N_18134,N_16918,N_16072);
xnor U18135 (N_18135,N_17505,N_17593);
nand U18136 (N_18136,N_16826,N_17949);
nor U18137 (N_18137,N_17519,N_17525);
and U18138 (N_18138,N_17068,N_17713);
and U18139 (N_18139,N_17130,N_16644);
and U18140 (N_18140,N_16190,N_16648);
or U18141 (N_18141,N_16718,N_17356);
xor U18142 (N_18142,N_17277,N_16167);
or U18143 (N_18143,N_17599,N_17978);
nor U18144 (N_18144,N_16327,N_16238);
or U18145 (N_18145,N_17468,N_17191);
and U18146 (N_18146,N_17414,N_17296);
or U18147 (N_18147,N_17874,N_16793);
and U18148 (N_18148,N_17341,N_16024);
nor U18149 (N_18149,N_16572,N_16028);
and U18150 (N_18150,N_16931,N_16829);
and U18151 (N_18151,N_17495,N_16023);
nand U18152 (N_18152,N_17646,N_16416);
nor U18153 (N_18153,N_17754,N_16216);
nand U18154 (N_18154,N_16403,N_16336);
nand U18155 (N_18155,N_16458,N_17895);
xnor U18156 (N_18156,N_17185,N_16259);
and U18157 (N_18157,N_16584,N_17654);
and U18158 (N_18158,N_17625,N_17260);
or U18159 (N_18159,N_16602,N_16422);
nor U18160 (N_18160,N_16067,N_16618);
xor U18161 (N_18161,N_16951,N_16795);
nor U18162 (N_18162,N_16760,N_16668);
and U18163 (N_18163,N_16748,N_16295);
nand U18164 (N_18164,N_16695,N_16978);
or U18165 (N_18165,N_17019,N_16031);
nand U18166 (N_18166,N_16061,N_16733);
xor U18167 (N_18167,N_17597,N_16460);
and U18168 (N_18168,N_16095,N_17172);
nand U18169 (N_18169,N_16477,N_17075);
xor U18170 (N_18170,N_16262,N_16203);
or U18171 (N_18171,N_17373,N_17404);
nor U18172 (N_18172,N_17009,N_17708);
nor U18173 (N_18173,N_16616,N_16901);
or U18174 (N_18174,N_17818,N_16846);
nand U18175 (N_18175,N_17144,N_16267);
and U18176 (N_18176,N_17165,N_17155);
xor U18177 (N_18177,N_17660,N_17458);
or U18178 (N_18178,N_16008,N_17758);
nand U18179 (N_18179,N_17846,N_17463);
or U18180 (N_18180,N_16082,N_17143);
and U18181 (N_18181,N_17573,N_16232);
and U18182 (N_18182,N_16412,N_16828);
xor U18183 (N_18183,N_16869,N_16307);
or U18184 (N_18184,N_17636,N_17205);
or U18185 (N_18185,N_16891,N_16395);
or U18186 (N_18186,N_17626,N_17452);
nor U18187 (N_18187,N_16533,N_17218);
nor U18188 (N_18188,N_16924,N_17147);
and U18189 (N_18189,N_17350,N_16505);
nor U18190 (N_18190,N_17491,N_16106);
xor U18191 (N_18191,N_16797,N_16487);
nand U18192 (N_18192,N_16451,N_17222);
and U18193 (N_18193,N_16275,N_16630);
or U18194 (N_18194,N_17856,N_16995);
xor U18195 (N_18195,N_16217,N_17821);
nand U18196 (N_18196,N_16497,N_17294);
and U18197 (N_18197,N_16172,N_17084);
and U18198 (N_18198,N_16961,N_16698);
and U18199 (N_18199,N_17901,N_16624);
nor U18200 (N_18200,N_16043,N_17462);
or U18201 (N_18201,N_16037,N_16428);
or U18202 (N_18202,N_16069,N_16847);
nand U18203 (N_18203,N_17007,N_16625);
or U18204 (N_18204,N_17632,N_17738);
and U18205 (N_18205,N_16489,N_17053);
xnor U18206 (N_18206,N_17622,N_16765);
or U18207 (N_18207,N_16818,N_17028);
nor U18208 (N_18208,N_17305,N_16261);
xor U18209 (N_18209,N_16385,N_16601);
nand U18210 (N_18210,N_16210,N_16233);
nor U18211 (N_18211,N_17245,N_17092);
nor U18212 (N_18212,N_17426,N_16405);
nand U18213 (N_18213,N_17442,N_16394);
nor U18214 (N_18214,N_17859,N_16864);
xnor U18215 (N_18215,N_17518,N_17716);
nor U18216 (N_18216,N_17889,N_17687);
or U18217 (N_18217,N_16772,N_17515);
nand U18218 (N_18218,N_16895,N_16466);
nor U18219 (N_18219,N_17229,N_17006);
and U18220 (N_18220,N_16180,N_16374);
and U18221 (N_18221,N_17402,N_17105);
nand U18222 (N_18222,N_16691,N_16433);
and U18223 (N_18223,N_16702,N_17301);
nand U18224 (N_18224,N_17823,N_16656);
nand U18225 (N_18225,N_16304,N_17782);
xor U18226 (N_18226,N_17138,N_16462);
or U18227 (N_18227,N_17419,N_16287);
xor U18228 (N_18228,N_17539,N_16960);
xnor U18229 (N_18229,N_17102,N_16306);
xor U18230 (N_18230,N_17470,N_17976);
or U18231 (N_18231,N_17101,N_17694);
xnor U18232 (N_18232,N_17735,N_16929);
nand U18233 (N_18233,N_16707,N_17706);
nor U18234 (N_18234,N_17911,N_17647);
xor U18235 (N_18235,N_16352,N_17984);
and U18236 (N_18236,N_16089,N_16982);
and U18237 (N_18237,N_16454,N_16026);
and U18238 (N_18238,N_16360,N_16502);
or U18239 (N_18239,N_17060,N_17829);
xor U18240 (N_18240,N_17896,N_17737);
and U18241 (N_18241,N_17933,N_16199);
nor U18242 (N_18242,N_16212,N_17934);
nand U18243 (N_18243,N_16706,N_16119);
or U18244 (N_18244,N_17083,N_16231);
and U18245 (N_18245,N_16188,N_16301);
xor U18246 (N_18246,N_16335,N_16421);
nand U18247 (N_18247,N_16160,N_16468);
and U18248 (N_18248,N_16014,N_17339);
nand U18249 (N_18249,N_16839,N_16481);
xnor U18250 (N_18250,N_16264,N_17142);
nand U18251 (N_18251,N_16575,N_16075);
xnor U18252 (N_18252,N_17293,N_17578);
and U18253 (N_18253,N_17096,N_17960);
nand U18254 (N_18254,N_17831,N_17079);
nor U18255 (N_18255,N_17669,N_16571);
and U18256 (N_18256,N_17562,N_17759);
and U18257 (N_18257,N_17220,N_16732);
or U18258 (N_18258,N_16244,N_17845);
and U18259 (N_18259,N_17928,N_16058);
or U18260 (N_18260,N_16088,N_16558);
and U18261 (N_18261,N_17650,N_17259);
xnor U18262 (N_18262,N_16239,N_16032);
and U18263 (N_18263,N_17692,N_17134);
and U18264 (N_18264,N_16034,N_16125);
nand U18265 (N_18265,N_17965,N_17595);
xnor U18266 (N_18266,N_17374,N_17812);
or U18267 (N_18267,N_16956,N_17046);
xor U18268 (N_18268,N_17784,N_17327);
nand U18269 (N_18269,N_16638,N_17945);
nand U18270 (N_18270,N_17420,N_16260);
and U18271 (N_18271,N_16042,N_17925);
nor U18272 (N_18272,N_17781,N_16957);
and U18273 (N_18273,N_16138,N_16499);
and U18274 (N_18274,N_16170,N_16705);
nand U18275 (N_18275,N_17855,N_16440);
and U18276 (N_18276,N_16017,N_17930);
nand U18277 (N_18277,N_17072,N_17364);
nand U18278 (N_18278,N_16438,N_17583);
nand U18279 (N_18279,N_16763,N_17906);
and U18280 (N_18280,N_16128,N_16329);
nand U18281 (N_18281,N_16971,N_17645);
or U18282 (N_18282,N_17044,N_16399);
xnor U18283 (N_18283,N_16815,N_16012);
nor U18284 (N_18284,N_17666,N_16701);
or U18285 (N_18285,N_17902,N_16506);
nor U18286 (N_18286,N_17815,N_17177);
xnor U18287 (N_18287,N_17684,N_16908);
nand U18288 (N_18288,N_17238,N_17257);
or U18289 (N_18289,N_16741,N_17062);
or U18290 (N_18290,N_16814,N_16970);
nand U18291 (N_18291,N_16002,N_17552);
nand U18292 (N_18292,N_16051,N_16746);
and U18293 (N_18293,N_17571,N_16993);
nand U18294 (N_18294,N_16279,N_16907);
xnor U18295 (N_18295,N_16643,N_17514);
or U18296 (N_18296,N_16984,N_16446);
nand U18297 (N_18297,N_17592,N_16528);
or U18298 (N_18298,N_17825,N_17566);
nor U18299 (N_18299,N_17233,N_17943);
nand U18300 (N_18300,N_17787,N_17276);
xnor U18301 (N_18301,N_16831,N_16380);
nor U18302 (N_18302,N_16062,N_16054);
or U18303 (N_18303,N_16611,N_17790);
nand U18304 (N_18304,N_17287,N_16619);
or U18305 (N_18305,N_16626,N_17340);
xor U18306 (N_18306,N_16676,N_16566);
nand U18307 (N_18307,N_17020,N_17297);
nor U18308 (N_18308,N_17064,N_16300);
nor U18309 (N_18309,N_17409,N_16021);
and U18310 (N_18310,N_17939,N_16009);
nand U18311 (N_18311,N_17324,N_17742);
or U18312 (N_18312,N_17545,N_17981);
xor U18313 (N_18313,N_17226,N_17234);
xnor U18314 (N_18314,N_16373,N_17556);
or U18315 (N_18315,N_16103,N_16560);
or U18316 (N_18316,N_16415,N_17851);
nand U18317 (N_18317,N_17135,N_17367);
and U18318 (N_18318,N_16333,N_17942);
or U18319 (N_18319,N_16079,N_17793);
or U18320 (N_18320,N_17532,N_17497);
nor U18321 (N_18321,N_17850,N_17378);
and U18322 (N_18322,N_16149,N_17482);
and U18323 (N_18323,N_17256,N_17330);
nor U18324 (N_18324,N_17792,N_16158);
and U18325 (N_18325,N_17190,N_16383);
and U18326 (N_18326,N_17938,N_17839);
xnor U18327 (N_18327,N_16065,N_17633);
nand U18328 (N_18328,N_16472,N_17637);
and U18329 (N_18329,N_17275,N_16997);
nor U18330 (N_18330,N_17095,N_17085);
nor U18331 (N_18331,N_16684,N_16153);
xor U18332 (N_18332,N_16860,N_16862);
nor U18333 (N_18333,N_16425,N_17816);
and U18334 (N_18334,N_17620,N_17640);
xnor U18335 (N_18335,N_16407,N_17557);
or U18336 (N_18336,N_16283,N_17014);
nand U18337 (N_18337,N_17071,N_16655);
nor U18338 (N_18338,N_17982,N_16324);
or U18339 (N_18339,N_16665,N_16568);
or U18340 (N_18340,N_16050,N_17045);
and U18341 (N_18341,N_16187,N_16063);
and U18342 (N_18342,N_17120,N_17741);
and U18343 (N_18343,N_17246,N_17390);
or U18344 (N_18344,N_16590,N_17336);
xor U18345 (N_18345,N_16049,N_16530);
xnor U18346 (N_18346,N_17274,N_16427);
xnor U18347 (N_18347,N_16320,N_16730);
or U18348 (N_18348,N_16962,N_16714);
and U18349 (N_18349,N_16803,N_16791);
or U18350 (N_18350,N_16154,N_17507);
and U18351 (N_18351,N_17115,N_17100);
nand U18352 (N_18352,N_16873,N_17407);
xor U18353 (N_18353,N_16114,N_17888);
and U18354 (N_18354,N_16402,N_16341);
or U18355 (N_18355,N_16822,N_16215);
or U18356 (N_18356,N_17959,N_16168);
nor U18357 (N_18357,N_16823,N_16581);
nand U18358 (N_18358,N_16926,N_17990);
nor U18359 (N_18359,N_17450,N_16056);
and U18360 (N_18360,N_17832,N_16139);
nand U18361 (N_18361,N_17021,N_17581);
or U18362 (N_18362,N_17541,N_17963);
nand U18363 (N_18363,N_17026,N_16667);
nor U18364 (N_18364,N_16234,N_17863);
or U18365 (N_18365,N_16202,N_17719);
and U18366 (N_18366,N_16570,N_16358);
xor U18367 (N_18367,N_17894,N_17041);
xnor U18368 (N_18368,N_17774,N_17817);
and U18369 (N_18369,N_17972,N_16491);
xor U18370 (N_18370,N_17524,N_16104);
nand U18371 (N_18371,N_16393,N_16711);
and U18372 (N_18372,N_16798,N_16640);
nor U18373 (N_18373,N_17721,N_16898);
xnor U18374 (N_18374,N_17284,N_17315);
or U18375 (N_18375,N_17493,N_16145);
or U18376 (N_18376,N_16946,N_16755);
or U18377 (N_18377,N_16194,N_16875);
and U18378 (N_18378,N_16731,N_16230);
or U18379 (N_18379,N_16242,N_16169);
nand U18380 (N_18380,N_16712,N_16932);
nand U18381 (N_18381,N_16939,N_17651);
nor U18382 (N_18382,N_16817,N_17869);
nand U18383 (N_18383,N_16704,N_16291);
or U18384 (N_18384,N_16273,N_17567);
nand U18385 (N_18385,N_17862,N_16896);
or U18386 (N_18386,N_16520,N_16091);
xor U18387 (N_18387,N_16071,N_16376);
and U18388 (N_18388,N_16764,N_17919);
xnor U18389 (N_18389,N_17961,N_16717);
and U18390 (N_18390,N_17740,N_17936);
nand U18391 (N_18391,N_17443,N_16435);
and U18392 (N_18392,N_17389,N_17003);
or U18393 (N_18393,N_16867,N_16411);
and U18394 (N_18394,N_16371,N_17076);
and U18395 (N_18395,N_17149,N_17870);
nor U18396 (N_18396,N_16550,N_17013);
or U18397 (N_18397,N_17671,N_16591);
xnor U18398 (N_18398,N_16564,N_16699);
and U18399 (N_18399,N_17940,N_17141);
or U18400 (N_18400,N_17762,N_17145);
xnor U18401 (N_18401,N_17150,N_16836);
or U18402 (N_18402,N_16972,N_17768);
nor U18403 (N_18403,N_17924,N_17964);
or U18404 (N_18404,N_17857,N_16227);
nand U18405 (N_18405,N_17313,N_17188);
xor U18406 (N_18406,N_17168,N_17544);
xnor U18407 (N_18407,N_17500,N_17528);
nor U18408 (N_18408,N_17077,N_16742);
or U18409 (N_18409,N_16744,N_17323);
xnor U18410 (N_18410,N_17322,N_16018);
or U18411 (N_18411,N_16703,N_16461);
or U18412 (N_18412,N_16547,N_16330);
and U18413 (N_18413,N_17999,N_16430);
nor U18414 (N_18414,N_17465,N_16813);
nand U18415 (N_18415,N_17722,N_17570);
nor U18416 (N_18416,N_17286,N_16623);
nor U18417 (N_18417,N_16645,N_17395);
nor U18418 (N_18418,N_17868,N_17070);
and U18419 (N_18419,N_16588,N_16432);
nand U18420 (N_18420,N_17022,N_17417);
or U18421 (N_18421,N_16391,N_17241);
or U18422 (N_18422,N_16409,N_16639);
xnor U18423 (N_18423,N_16127,N_16531);
nand U18424 (N_18424,N_17778,N_16185);
or U18425 (N_18425,N_17550,N_17321);
or U18426 (N_18426,N_17192,N_17116);
or U18427 (N_18427,N_16282,N_16258);
and U18428 (N_18428,N_17734,N_17212);
nand U18429 (N_18429,N_16431,N_17459);
nor U18430 (N_18430,N_16398,N_16495);
and U18431 (N_18431,N_17352,N_17148);
and U18432 (N_18432,N_17309,N_16739);
or U18433 (N_18433,N_16775,N_16894);
xnor U18434 (N_18434,N_16356,N_17347);
nor U18435 (N_18435,N_16673,N_17517);
nand U18436 (N_18436,N_16366,N_17089);
and U18437 (N_18437,N_16524,N_16252);
xnor U18438 (N_18438,N_16672,N_17406);
xor U18439 (N_18439,N_16824,N_17215);
xor U18440 (N_18440,N_17210,N_17431);
and U18441 (N_18441,N_16038,N_16893);
or U18442 (N_18442,N_16297,N_16688);
xor U18443 (N_18443,N_17361,N_17411);
xnor U18444 (N_18444,N_17156,N_17944);
xnor U18445 (N_18445,N_17531,N_16503);
nand U18446 (N_18446,N_17703,N_16589);
or U18447 (N_18447,N_17396,N_16426);
or U18448 (N_18448,N_16609,N_16992);
or U18449 (N_18449,N_16934,N_16925);
xnor U18450 (N_18450,N_17032,N_17035);
xnor U18451 (N_18451,N_17572,N_17113);
and U18452 (N_18452,N_16417,N_17509);
nor U18453 (N_18453,N_17900,N_16785);
nand U18454 (N_18454,N_16976,N_17929);
or U18455 (N_18455,N_17059,N_16020);
nor U18456 (N_18456,N_16783,N_17828);
nand U18457 (N_18457,N_16444,N_17265);
nor U18458 (N_18458,N_17698,N_16998);
and U18459 (N_18459,N_17750,N_16064);
xnor U18460 (N_18460,N_17199,N_16882);
or U18461 (N_18461,N_17005,N_17993);
xnor U18462 (N_18462,N_17609,N_17921);
and U18463 (N_18463,N_17838,N_16734);
and U18464 (N_18464,N_16884,N_17880);
and U18465 (N_18465,N_17724,N_17400);
nor U18466 (N_18466,N_16710,N_16085);
and U18467 (N_18467,N_16059,N_16276);
and U18468 (N_18468,N_16835,N_16914);
nor U18469 (N_18469,N_16599,N_16193);
and U18470 (N_18470,N_17588,N_16770);
nor U18471 (N_18471,N_16799,N_16191);
xnor U18472 (N_18472,N_16535,N_16107);
nand U18473 (N_18473,N_16134,N_16612);
or U18474 (N_18474,N_16186,N_16845);
nand U18475 (N_18475,N_16544,N_16109);
xnor U18476 (N_18476,N_16346,N_17582);
xor U18477 (N_18477,N_16840,N_17434);
xnor U18478 (N_18478,N_17914,N_17298);
nand U18479 (N_18479,N_17080,N_16771);
nor U18480 (N_18480,N_17802,N_17757);
xor U18481 (N_18481,N_16332,N_16131);
nand U18482 (N_18482,N_16035,N_17826);
xnor U18483 (N_18483,N_16317,N_16920);
nor U18484 (N_18484,N_17288,N_17393);
xor U18485 (N_18485,N_16299,N_17043);
or U18486 (N_18486,N_17680,N_16561);
and U18487 (N_18487,N_17890,N_17560);
nand U18488 (N_18488,N_17422,N_17283);
nand U18489 (N_18489,N_16959,N_17253);
nor U18490 (N_18490,N_17538,N_16678);
xor U18491 (N_18491,N_17490,N_16111);
nor U18492 (N_18492,N_17946,N_16856);
xnor U18493 (N_18493,N_16099,N_17752);
nand U18494 (N_18494,N_16800,N_16486);
or U18495 (N_18495,N_17137,N_17649);
nor U18496 (N_18496,N_16211,N_16465);
nand U18497 (N_18497,N_16789,N_17291);
xnor U18498 (N_18498,N_17844,N_16033);
and U18499 (N_18499,N_17791,N_17780);
nand U18500 (N_18500,N_17920,N_16540);
xor U18501 (N_18501,N_16833,N_16508);
and U18502 (N_18502,N_16370,N_17454);
or U18503 (N_18503,N_16713,N_17603);
and U18504 (N_18504,N_16923,N_16449);
and U18505 (N_18505,N_16361,N_17473);
or U18506 (N_18506,N_16607,N_17858);
nor U18507 (N_18507,N_16423,N_16790);
nor U18508 (N_18508,N_17915,N_17437);
or U18509 (N_18509,N_16903,N_16631);
and U18510 (N_18510,N_17591,N_17332);
xor U18511 (N_18511,N_16752,N_16097);
nand U18512 (N_18512,N_17174,N_16219);
nor U18513 (N_18513,N_17510,N_17872);
nand U18514 (N_18514,N_16788,N_17303);
nor U18515 (N_18515,N_17764,N_17983);
nor U18516 (N_18516,N_17012,N_17800);
nor U18517 (N_18517,N_17133,N_17412);
or U18518 (N_18518,N_17318,N_16047);
and U18519 (N_18519,N_17403,N_17325);
or U18520 (N_18520,N_17720,N_17363);
or U18521 (N_18521,N_17658,N_16225);
nor U18522 (N_18522,N_17010,N_16349);
nand U18523 (N_18523,N_16510,N_16314);
or U18524 (N_18524,N_16516,N_16404);
xor U18525 (N_18525,N_17227,N_16628);
nand U18526 (N_18526,N_17598,N_16102);
and U18527 (N_18527,N_16326,N_17893);
xor U18528 (N_18528,N_17948,N_17112);
and U18529 (N_18529,N_16256,N_17966);
and U18530 (N_18530,N_17975,N_16074);
and U18531 (N_18531,N_16007,N_16944);
nand U18532 (N_18532,N_17052,N_16514);
nand U18533 (N_18533,N_17655,N_17111);
nor U18534 (N_18534,N_16166,N_17534);
nand U18535 (N_18535,N_16541,N_17480);
and U18536 (N_18536,N_17910,N_16132);
xnor U18537 (N_18537,N_17478,N_16863);
nor U18538 (N_18538,N_16724,N_16293);
nor U18539 (N_18539,N_16700,N_16577);
nor U18540 (N_18540,N_17610,N_16532);
nor U18541 (N_18541,N_17086,N_16776);
and U18542 (N_18542,N_17621,N_17926);
or U18543 (N_18543,N_16906,N_17049);
nand U18544 (N_18544,N_16130,N_16582);
xnor U18545 (N_18545,N_17672,N_16999);
and U18546 (N_18546,N_16369,N_17249);
xnor U18547 (N_18547,N_16807,N_16308);
nor U18548 (N_18548,N_17601,N_17154);
nor U18549 (N_18549,N_16192,N_17445);
and U18550 (N_18550,N_17302,N_17840);
and U18551 (N_18551,N_16077,N_17653);
xor U18552 (N_18552,N_17195,N_17605);
xor U18553 (N_18553,N_17460,N_17522);
nand U18554 (N_18554,N_17613,N_16379);
and U18555 (N_18555,N_16880,N_17383);
and U18556 (N_18556,N_17536,N_17128);
nand U18557 (N_18557,N_16253,N_16142);
and U18558 (N_18558,N_16214,N_16027);
xnor U18559 (N_18559,N_16900,N_17710);
or U18560 (N_18560,N_17729,N_17564);
nand U18561 (N_18561,N_17248,N_17813);
or U18562 (N_18562,N_17104,N_17261);
and U18563 (N_18563,N_16610,N_17264);
nor U18564 (N_18564,N_16218,N_17164);
nor U18565 (N_18565,N_17642,N_16414);
or U18566 (N_18566,N_16347,N_16952);
nand U18567 (N_18567,N_16274,N_17952);
and U18568 (N_18568,N_17980,N_16837);
xor U18569 (N_18569,N_17686,N_17065);
xor U18570 (N_18570,N_17617,N_16853);
nand U18571 (N_18571,N_16464,N_17326);
nand U18572 (N_18572,N_17555,N_16725);
nor U18573 (N_18573,N_16313,N_16922);
xor U18574 (N_18574,N_16888,N_17749);
xnor U18575 (N_18575,N_17136,N_16909);
nand U18576 (N_18576,N_17618,N_17804);
and U18577 (N_18577,N_16762,N_16196);
nand U18578 (N_18578,N_17196,N_16362);
or U18579 (N_18579,N_16285,N_17424);
xor U18580 (N_18580,N_16989,N_16759);
and U18581 (N_18581,N_16679,N_17425);
nor U18582 (N_18582,N_17576,N_17530);
nor U18583 (N_18583,N_16224,N_16808);
xnor U18584 (N_18584,N_17553,N_16298);
and U18585 (N_18585,N_17405,N_17594);
and U18586 (N_18586,N_17801,N_16696);
xor U18587 (N_18587,N_16377,N_17369);
nor U18588 (N_18588,N_16682,N_17695);
nor U18589 (N_18589,N_17803,N_16965);
and U18590 (N_18590,N_17384,N_16322);
nand U18591 (N_18591,N_16592,N_17516);
nand U18592 (N_18592,N_16182,N_16500);
xor U18593 (N_18593,N_17271,N_17379);
nand U18594 (N_18594,N_16968,N_17231);
nand U18595 (N_18595,N_16179,N_16443);
nand U18596 (N_18596,N_17194,N_17047);
nor U18597 (N_18597,N_16538,N_17169);
xor U18598 (N_18598,N_17897,N_16559);
xor U18599 (N_18599,N_16669,N_17255);
nand U18600 (N_18600,N_16636,N_17580);
nor U18601 (N_18601,N_16045,N_17206);
or U18602 (N_18602,N_16315,N_16546);
nor U18603 (N_18603,N_17751,N_17486);
or U18604 (N_18604,N_16133,N_17129);
and U18605 (N_18605,N_17786,N_16161);
nand U18606 (N_18606,N_16325,N_17270);
and U18607 (N_18607,N_17985,N_16342);
or U18608 (N_18608,N_17991,N_16010);
nand U18609 (N_18609,N_17808,N_16878);
and U18610 (N_18610,N_17927,N_17756);
nand U18611 (N_18611,N_16539,N_17181);
nand U18612 (N_18612,N_17697,N_16116);
or U18613 (N_18613,N_16498,N_17054);
nand U18614 (N_18614,N_17988,N_17171);
and U18615 (N_18615,N_17091,N_16200);
nor U18616 (N_18616,N_16526,N_16255);
nand U18617 (N_18617,N_16606,N_17540);
nand U18618 (N_18618,N_17979,N_16877);
nand U18619 (N_18619,N_17628,N_17483);
nand U18620 (N_18620,N_17351,N_16986);
xnor U18621 (N_18621,N_17166,N_17042);
and U18622 (N_18622,N_17017,N_16935);
nand U18623 (N_18623,N_16794,N_17614);
and U18624 (N_18624,N_17110,N_16094);
and U18625 (N_18625,N_17848,N_16164);
or U18626 (N_18626,N_17415,N_17362);
and U18627 (N_18627,N_17469,N_16663);
and U18628 (N_18628,N_17551,N_16784);
nor U18629 (N_18629,N_17905,N_17476);
nand U18630 (N_18630,N_16950,N_16827);
nand U18631 (N_18631,N_16633,N_17207);
xor U18632 (N_18632,N_17527,N_17596);
xnor U18633 (N_18633,N_16151,N_16720);
or U18634 (N_18634,N_17744,N_17354);
xnor U18635 (N_18635,N_17892,N_17951);
and U18636 (N_18636,N_16716,N_17027);
nor U18637 (N_18637,N_16892,N_17258);
and U18638 (N_18638,N_17777,N_17600);
nor U18639 (N_18639,N_17311,N_17590);
nand U18640 (N_18640,N_17917,N_17444);
nor U18641 (N_18641,N_17726,N_17158);
or U18642 (N_18642,N_17345,N_17702);
and U18643 (N_18643,N_16221,N_17338);
nand U18644 (N_18644,N_17986,N_17266);
nor U18645 (N_18645,N_17670,N_17167);
nor U18646 (N_18646,N_17663,N_17811);
xor U18647 (N_18647,N_17512,N_16745);
and U18648 (N_18648,N_17667,N_16485);
xnor U18649 (N_18649,N_16046,N_17094);
and U18650 (N_18650,N_17506,N_16987);
and U18651 (N_18651,N_17736,N_17358);
or U18652 (N_18652,N_17066,N_16143);
nand U18653 (N_18653,N_16263,N_17039);
nor U18654 (N_18654,N_16483,N_16973);
xnor U18655 (N_18655,N_16019,N_17903);
or U18656 (N_18656,N_17202,N_17004);
or U18657 (N_18657,N_16816,N_17487);
or U18658 (N_18658,N_17050,N_16729);
nor U18659 (N_18659,N_16406,N_16470);
xnor U18660 (N_18660,N_17498,N_16247);
xor U18661 (N_18661,N_17521,N_16337);
or U18662 (N_18662,N_17745,N_16195);
and U18663 (N_18663,N_16229,N_17696);
and U18664 (N_18664,N_16413,N_16652);
or U18665 (N_18665,N_17664,N_17707);
or U18666 (N_18666,N_17688,N_16879);
and U18667 (N_18667,N_17794,N_17489);
nand U18668 (N_18668,N_16121,N_17225);
nand U18669 (N_18669,N_16490,N_17179);
or U18670 (N_18670,N_16098,N_17627);
xnor U18671 (N_18671,N_17548,N_17307);
nor U18672 (N_18672,N_16769,N_17883);
and U18673 (N_18673,N_17151,N_16204);
or U18674 (N_18674,N_16661,N_17239);
xor U18675 (N_18675,N_17082,N_17398);
xnor U18676 (N_18676,N_16272,N_17282);
nand U18677 (N_18677,N_16162,N_16476);
nor U18678 (N_18678,N_16157,N_16677);
xor U18679 (N_18679,N_17055,N_16323);
xnor U18680 (N_18680,N_16554,N_17511);
xnor U18681 (N_18681,N_16419,N_16666);
or U18682 (N_18682,N_16635,N_17546);
or U18683 (N_18683,N_16810,N_17765);
or U18684 (N_18684,N_17681,N_17446);
nor U18685 (N_18685,N_17123,N_17947);
and U18686 (N_18686,N_17496,N_17589);
nor U18687 (N_18687,N_16504,N_17448);
nor U18688 (N_18688,N_16156,N_17428);
and U18689 (N_18689,N_17163,N_17048);
nand U18690 (N_18690,N_17998,N_16687);
and U18691 (N_18691,N_17051,N_16311);
or U18692 (N_18692,N_16148,N_17088);
nor U18693 (N_18693,N_16052,N_17037);
or U18694 (N_18694,N_17606,N_17481);
nand U18695 (N_18695,N_16181,N_16686);
xor U18696 (N_18696,N_17175,N_16284);
nor U18697 (N_18697,N_16319,N_17824);
nand U18698 (N_18698,N_16265,N_16022);
and U18699 (N_18699,N_17725,N_16165);
and U18700 (N_18700,N_16303,N_16207);
nand U18701 (N_18701,N_17693,N_17543);
nand U18702 (N_18702,N_16948,N_16838);
nand U18703 (N_18703,N_17798,N_16041);
and U18704 (N_18704,N_17312,N_16613);
xor U18705 (N_18705,N_17230,N_16685);
xor U18706 (N_18706,N_17267,N_16851);
or U18707 (N_18707,N_16534,N_16397);
and U18708 (N_18708,N_16367,N_16228);
or U18709 (N_18709,N_16437,N_17314);
nand U18710 (N_18710,N_16552,N_17854);
nand U18711 (N_18711,N_17717,N_16178);
or U18712 (N_18712,N_17038,N_16136);
and U18713 (N_18713,N_17213,N_16343);
and U18714 (N_18714,N_16767,N_17704);
xor U18715 (N_18715,N_16305,N_17016);
xnor U18716 (N_18716,N_17299,N_17399);
xnor U18717 (N_18717,N_17820,N_17391);
nand U18718 (N_18718,N_16579,N_16980);
nand U18719 (N_18719,N_17278,N_16354);
nand U18720 (N_18720,N_16081,N_16938);
and U18721 (N_18721,N_17956,N_17629);
nor U18722 (N_18722,N_16594,N_17853);
and U18723 (N_18723,N_17796,N_17477);
nor U18724 (N_18724,N_17659,N_16348);
nand U18725 (N_18725,N_17638,N_17674);
or U18726 (N_18726,N_16576,N_17107);
nand U18727 (N_18727,N_17700,N_16693);
or U18728 (N_18728,N_17730,N_17449);
xor U18729 (N_18729,N_16055,N_17355);
or U18730 (N_18730,N_17346,N_17184);
xor U18731 (N_18731,N_17146,N_17783);
nand U18732 (N_18732,N_17769,N_17272);
or U18733 (N_18733,N_16453,N_16176);
and U18734 (N_18734,N_16459,N_16820);
nor U18735 (N_18735,N_17922,N_16070);
nor U18736 (N_18736,N_17743,N_16583);
or U18737 (N_18737,N_16392,N_16213);
nor U18738 (N_18738,N_17760,N_16761);
nand U18739 (N_18739,N_16509,N_16479);
xnor U18740 (N_18740,N_16954,N_16302);
nor U18741 (N_18741,N_17401,N_17878);
and U18742 (N_18742,N_16316,N_17849);
nor U18743 (N_18743,N_16177,N_16039);
nor U18744 (N_18744,N_16586,N_17935);
nand U18745 (N_18745,N_17413,N_17715);
xnor U18746 (N_18746,N_17967,N_17418);
or U18747 (N_18747,N_16281,N_16001);
and U18748 (N_18748,N_17197,N_16659);
nand U18749 (N_18749,N_17011,N_16488);
nand U18750 (N_18750,N_17771,N_16792);
or U18751 (N_18751,N_16410,N_16585);
and U18752 (N_18752,N_17484,N_17335);
and U18753 (N_18753,N_17739,N_16804);
xor U18754 (N_18754,N_16197,N_17882);
or U18755 (N_18755,N_17087,N_16173);
xnor U18756 (N_18756,N_16174,N_17748);
nand U18757 (N_18757,N_17579,N_17814);
and U18758 (N_18758,N_17186,N_16235);
or U18759 (N_18759,N_17300,N_17223);
xnor U18760 (N_18760,N_16100,N_17974);
or U18761 (N_18761,N_16053,N_17263);
and U18762 (N_18762,N_17030,N_17861);
and U18763 (N_18763,N_16897,N_16964);
xnor U18764 (N_18764,N_17607,N_16401);
nor U18765 (N_18765,N_17685,N_17714);
nor U18766 (N_18766,N_17977,N_16331);
nand U18767 (N_18767,N_17639,N_17439);
and U18768 (N_18768,N_16985,N_16025);
or U18769 (N_18769,N_17779,N_17971);
and U18770 (N_18770,N_17679,N_17365);
nor U18771 (N_18771,N_17881,N_17386);
or U18772 (N_18772,N_16674,N_16241);
and U18773 (N_18773,N_16641,N_16467);
nor U18774 (N_18774,N_17057,N_16854);
or U18775 (N_18775,N_16614,N_17466);
nand U18776 (N_18776,N_17887,N_17250);
and U18777 (N_18777,N_17860,N_17973);
or U18778 (N_18778,N_16345,N_16825);
nor U18779 (N_18779,N_16953,N_16357);
nor U18780 (N_18780,N_16569,N_16118);
nor U18781 (N_18781,N_17867,N_16654);
or U18782 (N_18782,N_17063,N_16294);
nor U18783 (N_18783,N_16469,N_17577);
and U18784 (N_18784,N_16029,N_16350);
xnor U18785 (N_18785,N_17099,N_16680);
or U18786 (N_18786,N_17841,N_16549);
xor U18787 (N_18787,N_16885,N_17310);
or U18788 (N_18788,N_17456,N_16093);
nor U18789 (N_18789,N_16841,N_17103);
xor U18790 (N_18790,N_17008,N_16709);
or U18791 (N_18791,N_17216,N_17795);
nand U18792 (N_18792,N_17513,N_17073);
or U18793 (N_18793,N_17221,N_16754);
or U18794 (N_18794,N_17251,N_17623);
nand U18795 (N_18795,N_17441,N_17847);
xor U18796 (N_18796,N_16637,N_16057);
nand U18797 (N_18797,N_16557,N_16598);
nor U18798 (N_18798,N_17029,N_16690);
nor U18799 (N_18799,N_17992,N_16280);
and U18800 (N_18800,N_16365,N_16507);
nand U18801 (N_18801,N_17408,N_16726);
nor U18802 (N_18802,N_17575,N_17932);
or U18803 (N_18803,N_16874,N_16974);
nor U18804 (N_18804,N_16375,N_17337);
and U18805 (N_18805,N_16866,N_16681);
nor U18806 (N_18806,N_16996,N_16650);
xor U18807 (N_18807,N_17772,N_17109);
xnor U18808 (N_18808,N_16796,N_16883);
and U18809 (N_18809,N_16257,N_17941);
or U18810 (N_18810,N_17344,N_17602);
xnor U18811 (N_18811,N_17117,N_17040);
nand U18812 (N_18812,N_17502,N_16236);
nand U18813 (N_18813,N_17228,N_16124);
xnor U18814 (N_18814,N_17269,N_17001);
and U18815 (N_18815,N_16849,N_16658);
nor U18816 (N_18816,N_16573,N_16084);
xor U18817 (N_18817,N_16621,N_17877);
nand U18818 (N_18818,N_17433,N_17036);
or U18819 (N_18819,N_16457,N_17289);
xnor U18820 (N_18820,N_16955,N_17131);
nor U18821 (N_18821,N_16595,N_16140);
nand U18822 (N_18822,N_16801,N_16334);
nor U18823 (N_18823,N_17201,N_17836);
nor U18824 (N_18824,N_16604,N_16527);
nor U18825 (N_18825,N_17842,N_16551);
or U18826 (N_18826,N_17873,N_17247);
and U18827 (N_18827,N_16240,N_16889);
nor U18828 (N_18828,N_16848,N_16086);
or U18829 (N_18829,N_16916,N_17969);
nor U18830 (N_18830,N_16384,N_17193);
xnor U18831 (N_18831,N_17366,N_16513);
nand U18832 (N_18832,N_17436,N_16222);
xor U18833 (N_18833,N_16565,N_16596);
xor U18834 (N_18834,N_17805,N_17180);
nor U18835 (N_18835,N_17152,N_16543);
nor U18836 (N_18836,N_16740,N_17788);
and U18837 (N_18837,N_16876,N_17957);
or U18838 (N_18838,N_16340,N_16478);
nand U18839 (N_18839,N_16117,N_16865);
or U18840 (N_18840,N_17388,N_16756);
nand U18841 (N_18841,N_17799,N_16205);
or U18842 (N_18842,N_16578,N_17689);
or U18843 (N_18843,N_17317,N_16309);
or U18844 (N_18844,N_16243,N_16664);
xnor U18845 (N_18845,N_16120,N_17397);
or U18846 (N_18846,N_16015,N_16927);
or U18847 (N_18847,N_16858,N_17290);
and U18848 (N_18848,N_17997,N_16269);
xor U18849 (N_18849,N_17262,N_16736);
xor U18850 (N_18850,N_16378,N_17766);
nand U18851 (N_18851,N_16270,N_17090);
nor U18852 (N_18852,N_16268,N_16902);
or U18853 (N_18853,N_17471,N_17711);
or U18854 (N_18854,N_16786,N_17464);
xor U18855 (N_18855,N_17360,N_16774);
xnor U18856 (N_18856,N_17864,N_16296);
nor U18857 (N_18857,N_17024,N_17822);
or U18858 (N_18858,N_17235,N_17067);
or U18859 (N_18859,N_16921,N_17394);
xnor U18860 (N_18860,N_17837,N_16424);
and U18861 (N_18861,N_17121,N_16937);
xor U18862 (N_18862,N_16587,N_17767);
and U18863 (N_18863,N_16574,N_17033);
and U18864 (N_18864,N_16249,N_17568);
xnor U18865 (N_18865,N_16452,N_17359);
and U18866 (N_18866,N_17421,N_16949);
nor U18867 (N_18867,N_16518,N_17334);
or U18868 (N_18868,N_16480,N_16522);
nand U18869 (N_18869,N_16542,N_16830);
or U18870 (N_18870,N_17189,N_17453);
xor U18871 (N_18871,N_16758,N_16886);
or U18872 (N_18872,N_16757,N_16492);
nand U18873 (N_18873,N_16159,N_17242);
xnor U18874 (N_18874,N_17968,N_16941);
xnor U18875 (N_18875,N_17244,N_17619);
or U18876 (N_18876,N_17034,N_16850);
or U18877 (N_18877,N_16246,N_17789);
nor U18878 (N_18878,N_16870,N_17209);
and U18879 (N_18879,N_17333,N_17479);
nand U18880 (N_18880,N_17475,N_16183);
nand U18881 (N_18881,N_16943,N_16629);
xor U18882 (N_18882,N_17807,N_17416);
or U18883 (N_18883,N_17319,N_17604);
or U18884 (N_18884,N_17994,N_17746);
or U18885 (N_18885,N_17348,N_16780);
nand U18886 (N_18886,N_17132,N_17648);
and U18887 (N_18887,N_16066,N_17996);
xnor U18888 (N_18888,N_16436,N_17106);
or U18889 (N_18889,N_17833,N_16805);
or U18890 (N_18890,N_17176,N_16447);
or U18891 (N_18891,N_16988,N_17574);
nand U18892 (N_18892,N_16536,N_17173);
xnor U18893 (N_18893,N_17081,N_16030);
xor U18894 (N_18894,N_16735,N_16983);
nand U18895 (N_18895,N_17061,N_16843);
xnor U18896 (N_18896,N_17183,N_16915);
xnor U18897 (N_18897,N_16861,N_16753);
xor U18898 (N_18898,N_16254,N_16087);
nor U18899 (N_18899,N_16580,N_16175);
or U18900 (N_18900,N_17198,N_16288);
nor U18901 (N_18901,N_16445,N_17162);
and U18902 (N_18902,N_16523,N_17118);
nand U18903 (N_18903,N_17537,N_17031);
nor U18904 (N_18904,N_17668,N_16671);
and U18905 (N_18905,N_16418,N_17240);
xnor U18906 (N_18906,N_16750,N_16515);
or U18907 (N_18907,N_17586,N_17387);
nor U18908 (N_18908,N_17611,N_17122);
nand U18909 (N_18909,N_16743,N_16141);
xor U18910 (N_18910,N_16632,N_16171);
xor U18911 (N_18911,N_17683,N_17909);
xnor U18912 (N_18912,N_17753,N_17701);
or U18913 (N_18913,N_17316,N_16073);
nor U18914 (N_18914,N_16647,N_16126);
xnor U18915 (N_18915,N_17731,N_17584);
nor U18916 (N_18916,N_17023,N_17843);
or U18917 (N_18917,N_17217,N_16627);
nand U18918 (N_18918,N_17268,N_16344);
and U18919 (N_18919,N_16749,N_17368);
or U18920 (N_18920,N_17243,N_16622);
xnor U18921 (N_18921,N_16013,N_17357);
xor U18922 (N_18922,N_16147,N_16112);
nand U18923 (N_18923,N_17204,N_16484);
nand U18924 (N_18924,N_16096,N_17320);
xnor U18925 (N_18925,N_16006,N_16450);
nor U18926 (N_18926,N_16721,N_16390);
and U18927 (N_18927,N_16004,N_17342);
or U18928 (N_18928,N_17747,N_16593);
or U18929 (N_18929,N_17676,N_16387);
or U18930 (N_18930,N_17549,N_16766);
and U18931 (N_18931,N_16694,N_16408);
nand U18932 (N_18932,N_16615,N_17211);
xor U18933 (N_18933,N_16727,N_16312);
or U18934 (N_18934,N_17157,N_16608);
and U18935 (N_18935,N_17178,N_17002);
xor U18936 (N_18936,N_16600,N_17705);
or U18937 (N_18937,N_17381,N_16003);
or U18938 (N_18938,N_17254,N_16517);
nand U18939 (N_18939,N_16940,N_17827);
xor U18940 (N_18940,N_17219,N_17678);
and U18941 (N_18941,N_17904,N_16016);
xor U18942 (N_18942,N_16890,N_16990);
and U18943 (N_18943,N_16388,N_16355);
xor U18944 (N_18944,N_16493,N_17508);
or U18945 (N_18945,N_17918,N_17056);
or U18946 (N_18946,N_17727,N_17410);
and U18947 (N_18947,N_17492,N_17630);
and U18948 (N_18948,N_17806,N_16511);
or U18949 (N_18949,N_16738,N_16372);
xnor U18950 (N_18950,N_17078,N_16501);
nand U18951 (N_18951,N_16977,N_16429);
and U18952 (N_18952,N_17542,N_16722);
xnor U18953 (N_18953,N_16852,N_16567);
or U18954 (N_18954,N_16857,N_17970);
nand U18955 (N_18955,N_16321,N_16101);
and U18956 (N_18956,N_17503,N_17520);
or U18957 (N_18957,N_17208,N_16040);
xor U18958 (N_18958,N_17093,N_17224);
nor U18959 (N_18959,N_17472,N_17423);
nor U18960 (N_18960,N_16146,N_17643);
xnor U18961 (N_18961,N_17718,N_16382);
nand U18962 (N_18962,N_16905,N_16911);
nand U18963 (N_18963,N_17891,N_16092);
nor U18964 (N_18964,N_16250,N_16751);
nand U18965 (N_18965,N_17375,N_16220);
or U18966 (N_18966,N_16519,N_16806);
xor U18967 (N_18967,N_17435,N_16011);
nand U18968 (N_18968,N_16144,N_16005);
nand U18969 (N_18969,N_16113,N_17461);
nand U18970 (N_18970,N_17236,N_17652);
and U18971 (N_18971,N_16936,N_16819);
nor U18972 (N_18972,N_16651,N_16083);
nor U18973 (N_18973,N_16529,N_16634);
or U18974 (N_18974,N_17125,N_16555);
nor U18975 (N_18975,N_16339,N_17273);
and U18976 (N_18976,N_17203,N_17153);
xnor U18977 (N_18977,N_17785,N_17561);
nand U18978 (N_18978,N_17501,N_17912);
xnor U18979 (N_18979,N_16163,N_17885);
nand U18980 (N_18980,N_16000,N_17279);
xnor U18981 (N_18981,N_17819,N_16368);
nand U18982 (N_18982,N_16947,N_17587);
nor U18983 (N_18983,N_16887,N_16979);
or U18984 (N_18984,N_16496,N_17140);
xnor U18985 (N_18985,N_17634,N_16208);
xnor U18986 (N_18986,N_17429,N_16137);
nor U18987 (N_18987,N_16278,N_16649);
and U18988 (N_18988,N_17308,N_16364);
and U18989 (N_18989,N_16080,N_16812);
nor U18990 (N_18990,N_17776,N_16910);
and U18991 (N_18991,N_16942,N_17953);
or U18992 (N_18992,N_17866,N_17447);
or U18993 (N_18993,N_17733,N_16359);
and U18994 (N_18994,N_16135,N_16525);
nor U18995 (N_18995,N_16855,N_17641);
or U18996 (N_18996,N_16966,N_16123);
nand U18997 (N_18997,N_17797,N_16396);
and U18998 (N_18998,N_17728,N_17485);
nor U18999 (N_18999,N_16434,N_16975);
xnor U19000 (N_19000,N_17273,N_16771);
xor U19001 (N_19001,N_17316,N_16218);
xnor U19002 (N_19002,N_17601,N_17776);
nand U19003 (N_19003,N_16750,N_17065);
and U19004 (N_19004,N_17543,N_17807);
or U19005 (N_19005,N_16116,N_17259);
xor U19006 (N_19006,N_17258,N_17055);
nor U19007 (N_19007,N_17508,N_17671);
nor U19008 (N_19008,N_16180,N_17695);
nor U19009 (N_19009,N_17213,N_17918);
nor U19010 (N_19010,N_16030,N_16667);
nor U19011 (N_19011,N_17848,N_17017);
and U19012 (N_19012,N_16925,N_17467);
xnor U19013 (N_19013,N_16056,N_17581);
nand U19014 (N_19014,N_17078,N_17717);
nor U19015 (N_19015,N_17849,N_17187);
or U19016 (N_19016,N_16300,N_16910);
nor U19017 (N_19017,N_16526,N_17625);
and U19018 (N_19018,N_17063,N_16146);
and U19019 (N_19019,N_16199,N_16118);
or U19020 (N_19020,N_17887,N_16879);
and U19021 (N_19021,N_16492,N_17603);
and U19022 (N_19022,N_16399,N_16156);
or U19023 (N_19023,N_16728,N_16666);
nand U19024 (N_19024,N_17776,N_16887);
nor U19025 (N_19025,N_17855,N_17147);
nor U19026 (N_19026,N_16432,N_17366);
xor U19027 (N_19027,N_17607,N_16140);
and U19028 (N_19028,N_17507,N_17266);
or U19029 (N_19029,N_17506,N_17510);
xor U19030 (N_19030,N_17016,N_17093);
or U19031 (N_19031,N_16202,N_17131);
xor U19032 (N_19032,N_16257,N_17782);
or U19033 (N_19033,N_16171,N_17944);
and U19034 (N_19034,N_17364,N_17234);
nor U19035 (N_19035,N_17328,N_17326);
and U19036 (N_19036,N_17041,N_17531);
xor U19037 (N_19037,N_17720,N_16525);
nand U19038 (N_19038,N_16431,N_16163);
nand U19039 (N_19039,N_16055,N_17584);
xnor U19040 (N_19040,N_16892,N_17676);
and U19041 (N_19041,N_16319,N_17906);
nand U19042 (N_19042,N_16020,N_16945);
or U19043 (N_19043,N_16533,N_17093);
or U19044 (N_19044,N_17536,N_16059);
nand U19045 (N_19045,N_16225,N_17147);
xor U19046 (N_19046,N_17190,N_16744);
nand U19047 (N_19047,N_16798,N_16316);
or U19048 (N_19048,N_17066,N_16189);
nand U19049 (N_19049,N_16891,N_16463);
nor U19050 (N_19050,N_17833,N_17520);
nand U19051 (N_19051,N_16090,N_17043);
nor U19052 (N_19052,N_17354,N_16852);
and U19053 (N_19053,N_17459,N_17191);
and U19054 (N_19054,N_17025,N_16377);
nor U19055 (N_19055,N_17647,N_17612);
nor U19056 (N_19056,N_17680,N_16066);
nand U19057 (N_19057,N_16177,N_17265);
or U19058 (N_19058,N_16495,N_16910);
nand U19059 (N_19059,N_17483,N_16198);
and U19060 (N_19060,N_16639,N_16181);
nand U19061 (N_19061,N_16470,N_17550);
nor U19062 (N_19062,N_16399,N_16161);
xor U19063 (N_19063,N_17305,N_16647);
xor U19064 (N_19064,N_16209,N_16674);
and U19065 (N_19065,N_17846,N_17286);
nor U19066 (N_19066,N_17522,N_17089);
xor U19067 (N_19067,N_17586,N_17835);
xor U19068 (N_19068,N_17493,N_16590);
nand U19069 (N_19069,N_16397,N_17439);
and U19070 (N_19070,N_17973,N_16509);
or U19071 (N_19071,N_16933,N_16290);
and U19072 (N_19072,N_16332,N_16320);
nor U19073 (N_19073,N_17990,N_17202);
nand U19074 (N_19074,N_16607,N_16455);
or U19075 (N_19075,N_17979,N_17430);
nand U19076 (N_19076,N_17377,N_16276);
xor U19077 (N_19077,N_17616,N_17464);
and U19078 (N_19078,N_17444,N_17893);
nor U19079 (N_19079,N_16782,N_16023);
nor U19080 (N_19080,N_16932,N_17618);
and U19081 (N_19081,N_17832,N_17185);
nor U19082 (N_19082,N_17137,N_17342);
or U19083 (N_19083,N_16815,N_16359);
and U19084 (N_19084,N_17624,N_16218);
and U19085 (N_19085,N_17914,N_17493);
and U19086 (N_19086,N_17673,N_17512);
xnor U19087 (N_19087,N_16331,N_17359);
xnor U19088 (N_19088,N_16071,N_17564);
or U19089 (N_19089,N_17899,N_17619);
nand U19090 (N_19090,N_16354,N_16106);
nor U19091 (N_19091,N_16733,N_16950);
xor U19092 (N_19092,N_17818,N_16587);
or U19093 (N_19093,N_17918,N_17845);
xnor U19094 (N_19094,N_17108,N_17287);
or U19095 (N_19095,N_17050,N_16954);
nand U19096 (N_19096,N_17732,N_17919);
or U19097 (N_19097,N_16987,N_17821);
and U19098 (N_19098,N_17214,N_17525);
xor U19099 (N_19099,N_16314,N_17428);
nor U19100 (N_19100,N_16687,N_16443);
xnor U19101 (N_19101,N_16308,N_17166);
or U19102 (N_19102,N_17857,N_16520);
xnor U19103 (N_19103,N_17705,N_17880);
nor U19104 (N_19104,N_17676,N_16651);
or U19105 (N_19105,N_16705,N_17973);
nor U19106 (N_19106,N_17640,N_17449);
and U19107 (N_19107,N_16221,N_16667);
or U19108 (N_19108,N_17868,N_16974);
or U19109 (N_19109,N_16777,N_16686);
or U19110 (N_19110,N_16808,N_16465);
and U19111 (N_19111,N_16618,N_16085);
nand U19112 (N_19112,N_16405,N_16394);
or U19113 (N_19113,N_16389,N_16318);
nand U19114 (N_19114,N_16617,N_17879);
nand U19115 (N_19115,N_16346,N_17943);
and U19116 (N_19116,N_16712,N_16125);
nor U19117 (N_19117,N_17982,N_16459);
nand U19118 (N_19118,N_17735,N_17668);
or U19119 (N_19119,N_16317,N_16130);
nor U19120 (N_19120,N_16433,N_17963);
or U19121 (N_19121,N_17053,N_17371);
and U19122 (N_19122,N_16456,N_16606);
and U19123 (N_19123,N_16830,N_16510);
nor U19124 (N_19124,N_17462,N_16629);
and U19125 (N_19125,N_16016,N_16454);
or U19126 (N_19126,N_17569,N_16072);
nand U19127 (N_19127,N_16309,N_16063);
nor U19128 (N_19128,N_17311,N_16521);
xor U19129 (N_19129,N_17940,N_16691);
xor U19130 (N_19130,N_17453,N_16426);
or U19131 (N_19131,N_17333,N_17457);
xnor U19132 (N_19132,N_16085,N_17778);
xnor U19133 (N_19133,N_17859,N_17122);
nor U19134 (N_19134,N_16249,N_17400);
and U19135 (N_19135,N_16099,N_16357);
xnor U19136 (N_19136,N_16518,N_17171);
nand U19137 (N_19137,N_17596,N_16404);
nand U19138 (N_19138,N_17482,N_16685);
nand U19139 (N_19139,N_16764,N_17484);
xnor U19140 (N_19140,N_17290,N_16825);
or U19141 (N_19141,N_17220,N_17814);
nand U19142 (N_19142,N_17240,N_16625);
nor U19143 (N_19143,N_16378,N_16737);
nand U19144 (N_19144,N_16496,N_17130);
nor U19145 (N_19145,N_17261,N_16150);
xnor U19146 (N_19146,N_16725,N_16741);
nor U19147 (N_19147,N_16702,N_16573);
or U19148 (N_19148,N_16577,N_16520);
nand U19149 (N_19149,N_16706,N_17772);
nor U19150 (N_19150,N_16108,N_16230);
and U19151 (N_19151,N_17956,N_17013);
nand U19152 (N_19152,N_17094,N_16134);
nor U19153 (N_19153,N_16081,N_16955);
and U19154 (N_19154,N_16314,N_17865);
or U19155 (N_19155,N_17973,N_16806);
xor U19156 (N_19156,N_17792,N_17662);
nor U19157 (N_19157,N_16591,N_17698);
nand U19158 (N_19158,N_16708,N_16095);
nand U19159 (N_19159,N_17849,N_17998);
xor U19160 (N_19160,N_16162,N_17736);
nand U19161 (N_19161,N_16423,N_16364);
xnor U19162 (N_19162,N_16682,N_17396);
xor U19163 (N_19163,N_17529,N_16988);
xnor U19164 (N_19164,N_17966,N_16308);
nand U19165 (N_19165,N_17747,N_16055);
and U19166 (N_19166,N_17350,N_16234);
xnor U19167 (N_19167,N_17509,N_16303);
and U19168 (N_19168,N_17016,N_16545);
nand U19169 (N_19169,N_17841,N_17040);
nor U19170 (N_19170,N_17488,N_16885);
and U19171 (N_19171,N_17667,N_16988);
nor U19172 (N_19172,N_16474,N_17956);
nand U19173 (N_19173,N_16793,N_16143);
or U19174 (N_19174,N_16157,N_16890);
and U19175 (N_19175,N_17205,N_16979);
or U19176 (N_19176,N_16253,N_16085);
nand U19177 (N_19177,N_17682,N_17913);
xnor U19178 (N_19178,N_17220,N_17586);
xor U19179 (N_19179,N_16901,N_16927);
nand U19180 (N_19180,N_17393,N_16301);
xnor U19181 (N_19181,N_16018,N_17668);
or U19182 (N_19182,N_16076,N_17071);
nor U19183 (N_19183,N_16490,N_16381);
nand U19184 (N_19184,N_16858,N_17442);
or U19185 (N_19185,N_17875,N_16135);
and U19186 (N_19186,N_17509,N_17553);
nor U19187 (N_19187,N_16513,N_16369);
and U19188 (N_19188,N_17349,N_17276);
nor U19189 (N_19189,N_16763,N_17772);
nor U19190 (N_19190,N_16220,N_17656);
and U19191 (N_19191,N_16504,N_16340);
or U19192 (N_19192,N_16208,N_16015);
nand U19193 (N_19193,N_16017,N_17890);
and U19194 (N_19194,N_16310,N_17175);
nor U19195 (N_19195,N_17501,N_16699);
and U19196 (N_19196,N_17904,N_16576);
nand U19197 (N_19197,N_16439,N_16766);
nor U19198 (N_19198,N_17256,N_16884);
or U19199 (N_19199,N_17156,N_16000);
xnor U19200 (N_19200,N_16431,N_16782);
nand U19201 (N_19201,N_16409,N_16175);
or U19202 (N_19202,N_17405,N_16964);
nor U19203 (N_19203,N_16061,N_16545);
nand U19204 (N_19204,N_16336,N_17189);
and U19205 (N_19205,N_17565,N_17671);
and U19206 (N_19206,N_16761,N_17773);
or U19207 (N_19207,N_16387,N_16492);
nor U19208 (N_19208,N_17002,N_17691);
nor U19209 (N_19209,N_17774,N_17760);
nor U19210 (N_19210,N_17941,N_17223);
and U19211 (N_19211,N_16566,N_17914);
nor U19212 (N_19212,N_16764,N_17718);
nor U19213 (N_19213,N_16122,N_16009);
and U19214 (N_19214,N_17802,N_17267);
and U19215 (N_19215,N_17497,N_17735);
nand U19216 (N_19216,N_17666,N_17908);
and U19217 (N_19217,N_16607,N_16877);
or U19218 (N_19218,N_16426,N_17171);
or U19219 (N_19219,N_17936,N_17482);
xor U19220 (N_19220,N_17849,N_17055);
xnor U19221 (N_19221,N_17655,N_16521);
xor U19222 (N_19222,N_17747,N_16084);
nand U19223 (N_19223,N_16938,N_16027);
and U19224 (N_19224,N_17105,N_16430);
and U19225 (N_19225,N_17321,N_17075);
and U19226 (N_19226,N_17573,N_17139);
nand U19227 (N_19227,N_16694,N_16218);
nor U19228 (N_19228,N_17604,N_16962);
nand U19229 (N_19229,N_17951,N_17847);
nand U19230 (N_19230,N_17286,N_16914);
and U19231 (N_19231,N_16657,N_17066);
xor U19232 (N_19232,N_17664,N_16645);
nand U19233 (N_19233,N_16539,N_17928);
xnor U19234 (N_19234,N_17649,N_17958);
xnor U19235 (N_19235,N_16949,N_17847);
nor U19236 (N_19236,N_16601,N_17483);
or U19237 (N_19237,N_17041,N_16841);
or U19238 (N_19238,N_17720,N_16557);
and U19239 (N_19239,N_17614,N_16967);
or U19240 (N_19240,N_16564,N_16241);
xor U19241 (N_19241,N_17923,N_16159);
xnor U19242 (N_19242,N_16479,N_17719);
xnor U19243 (N_19243,N_17356,N_17521);
and U19244 (N_19244,N_16397,N_16684);
or U19245 (N_19245,N_16193,N_17445);
nand U19246 (N_19246,N_16436,N_16386);
or U19247 (N_19247,N_16189,N_17109);
nand U19248 (N_19248,N_17688,N_16946);
nand U19249 (N_19249,N_16466,N_16886);
nor U19250 (N_19250,N_17976,N_17713);
nor U19251 (N_19251,N_16187,N_17329);
or U19252 (N_19252,N_16563,N_16941);
nor U19253 (N_19253,N_16855,N_17014);
or U19254 (N_19254,N_17740,N_16736);
nand U19255 (N_19255,N_17254,N_17336);
nand U19256 (N_19256,N_16104,N_16281);
and U19257 (N_19257,N_17431,N_16771);
and U19258 (N_19258,N_16963,N_16717);
nor U19259 (N_19259,N_16108,N_16373);
nand U19260 (N_19260,N_16903,N_17041);
nand U19261 (N_19261,N_16934,N_17326);
and U19262 (N_19262,N_17815,N_16807);
xnor U19263 (N_19263,N_16014,N_17175);
or U19264 (N_19264,N_17240,N_16423);
nor U19265 (N_19265,N_17259,N_17834);
nor U19266 (N_19266,N_17475,N_16582);
nor U19267 (N_19267,N_16683,N_16128);
nor U19268 (N_19268,N_17525,N_17724);
and U19269 (N_19269,N_16571,N_17552);
xor U19270 (N_19270,N_16675,N_17946);
nand U19271 (N_19271,N_16370,N_16426);
or U19272 (N_19272,N_16246,N_16719);
and U19273 (N_19273,N_16482,N_16782);
nand U19274 (N_19274,N_16476,N_16319);
xor U19275 (N_19275,N_16149,N_16968);
or U19276 (N_19276,N_16374,N_16429);
and U19277 (N_19277,N_17712,N_16075);
and U19278 (N_19278,N_16458,N_17815);
nor U19279 (N_19279,N_16354,N_17723);
nand U19280 (N_19280,N_16782,N_16942);
or U19281 (N_19281,N_17958,N_17886);
or U19282 (N_19282,N_16948,N_16680);
nor U19283 (N_19283,N_16434,N_17426);
or U19284 (N_19284,N_17224,N_17692);
nand U19285 (N_19285,N_17131,N_16932);
xnor U19286 (N_19286,N_17548,N_16167);
nand U19287 (N_19287,N_16418,N_16043);
or U19288 (N_19288,N_16868,N_16285);
or U19289 (N_19289,N_17652,N_17455);
and U19290 (N_19290,N_17218,N_17633);
xnor U19291 (N_19291,N_17333,N_16181);
nand U19292 (N_19292,N_17790,N_17845);
xnor U19293 (N_19293,N_17591,N_17385);
nand U19294 (N_19294,N_17888,N_16674);
or U19295 (N_19295,N_16309,N_16845);
xor U19296 (N_19296,N_16853,N_17811);
nor U19297 (N_19297,N_17549,N_16291);
nor U19298 (N_19298,N_16393,N_16818);
nor U19299 (N_19299,N_16777,N_17480);
or U19300 (N_19300,N_17709,N_17023);
nand U19301 (N_19301,N_16935,N_17451);
nand U19302 (N_19302,N_17492,N_17245);
nand U19303 (N_19303,N_16842,N_16560);
xnor U19304 (N_19304,N_16798,N_17177);
nand U19305 (N_19305,N_16269,N_17329);
or U19306 (N_19306,N_17886,N_16625);
and U19307 (N_19307,N_16427,N_17602);
or U19308 (N_19308,N_17670,N_17990);
nor U19309 (N_19309,N_17424,N_17119);
nor U19310 (N_19310,N_16136,N_17225);
nand U19311 (N_19311,N_16741,N_17918);
or U19312 (N_19312,N_17953,N_17870);
or U19313 (N_19313,N_17128,N_17597);
and U19314 (N_19314,N_17348,N_16509);
and U19315 (N_19315,N_16028,N_17090);
xor U19316 (N_19316,N_16461,N_17128);
xnor U19317 (N_19317,N_16895,N_17809);
and U19318 (N_19318,N_17790,N_16202);
xnor U19319 (N_19319,N_17821,N_17443);
nand U19320 (N_19320,N_16863,N_16710);
or U19321 (N_19321,N_16609,N_16982);
and U19322 (N_19322,N_17496,N_17875);
xor U19323 (N_19323,N_16961,N_17953);
and U19324 (N_19324,N_17807,N_17112);
nand U19325 (N_19325,N_16749,N_17946);
or U19326 (N_19326,N_16355,N_17901);
and U19327 (N_19327,N_17233,N_17167);
or U19328 (N_19328,N_17532,N_16528);
nor U19329 (N_19329,N_17337,N_16012);
xnor U19330 (N_19330,N_17809,N_16966);
nor U19331 (N_19331,N_17768,N_17807);
or U19332 (N_19332,N_17121,N_17215);
xnor U19333 (N_19333,N_16829,N_17598);
or U19334 (N_19334,N_16460,N_17189);
or U19335 (N_19335,N_16558,N_17260);
nand U19336 (N_19336,N_17695,N_17206);
xor U19337 (N_19337,N_17116,N_16789);
or U19338 (N_19338,N_16062,N_17115);
or U19339 (N_19339,N_16306,N_17068);
nand U19340 (N_19340,N_16369,N_16942);
or U19341 (N_19341,N_17813,N_16310);
nand U19342 (N_19342,N_16544,N_16767);
nor U19343 (N_19343,N_17685,N_17065);
nand U19344 (N_19344,N_16427,N_17927);
or U19345 (N_19345,N_16134,N_16679);
xor U19346 (N_19346,N_16191,N_17872);
or U19347 (N_19347,N_17055,N_16648);
nor U19348 (N_19348,N_16732,N_17833);
nor U19349 (N_19349,N_16112,N_17084);
nor U19350 (N_19350,N_16605,N_16746);
nand U19351 (N_19351,N_16223,N_16816);
or U19352 (N_19352,N_17184,N_16198);
or U19353 (N_19353,N_17756,N_17134);
or U19354 (N_19354,N_17274,N_17242);
xor U19355 (N_19355,N_17153,N_16466);
or U19356 (N_19356,N_17378,N_17463);
nand U19357 (N_19357,N_17034,N_16125);
nor U19358 (N_19358,N_16662,N_17180);
nand U19359 (N_19359,N_16828,N_16815);
nand U19360 (N_19360,N_16683,N_16359);
or U19361 (N_19361,N_16778,N_17389);
nor U19362 (N_19362,N_17547,N_17286);
nor U19363 (N_19363,N_17782,N_16854);
nand U19364 (N_19364,N_17318,N_16697);
xor U19365 (N_19365,N_17614,N_17092);
and U19366 (N_19366,N_16626,N_16773);
and U19367 (N_19367,N_16300,N_17298);
and U19368 (N_19368,N_17041,N_16551);
nand U19369 (N_19369,N_17214,N_16033);
or U19370 (N_19370,N_16486,N_17568);
nor U19371 (N_19371,N_16573,N_16050);
nand U19372 (N_19372,N_16983,N_16941);
xnor U19373 (N_19373,N_17474,N_17592);
xnor U19374 (N_19374,N_16940,N_16058);
nand U19375 (N_19375,N_16988,N_16238);
xnor U19376 (N_19376,N_17207,N_16259);
nand U19377 (N_19377,N_16795,N_16314);
xnor U19378 (N_19378,N_16153,N_17564);
or U19379 (N_19379,N_16195,N_17020);
or U19380 (N_19380,N_17506,N_17207);
or U19381 (N_19381,N_16980,N_16698);
nand U19382 (N_19382,N_16021,N_17024);
or U19383 (N_19383,N_17816,N_17272);
and U19384 (N_19384,N_16769,N_16443);
xnor U19385 (N_19385,N_17016,N_17368);
or U19386 (N_19386,N_17731,N_16599);
xor U19387 (N_19387,N_16574,N_17369);
and U19388 (N_19388,N_16924,N_16288);
nand U19389 (N_19389,N_16596,N_16991);
and U19390 (N_19390,N_16934,N_16399);
xnor U19391 (N_19391,N_17077,N_17013);
or U19392 (N_19392,N_16163,N_16268);
nand U19393 (N_19393,N_16984,N_16613);
xor U19394 (N_19394,N_16778,N_17365);
or U19395 (N_19395,N_16562,N_16627);
xnor U19396 (N_19396,N_16727,N_17465);
and U19397 (N_19397,N_17639,N_16987);
and U19398 (N_19398,N_17708,N_17606);
xor U19399 (N_19399,N_17583,N_17412);
and U19400 (N_19400,N_16289,N_16565);
nand U19401 (N_19401,N_17433,N_16720);
or U19402 (N_19402,N_17627,N_16185);
nor U19403 (N_19403,N_16002,N_17729);
or U19404 (N_19404,N_17493,N_16012);
nand U19405 (N_19405,N_16517,N_16862);
nor U19406 (N_19406,N_17618,N_16478);
xnor U19407 (N_19407,N_17430,N_16241);
or U19408 (N_19408,N_17891,N_16827);
nor U19409 (N_19409,N_17275,N_17014);
and U19410 (N_19410,N_17789,N_16251);
and U19411 (N_19411,N_17456,N_16915);
xor U19412 (N_19412,N_16047,N_16156);
nor U19413 (N_19413,N_16347,N_17399);
nand U19414 (N_19414,N_16796,N_17237);
nor U19415 (N_19415,N_17626,N_17374);
nor U19416 (N_19416,N_16985,N_17868);
nor U19417 (N_19417,N_16124,N_16882);
or U19418 (N_19418,N_16960,N_17476);
xnor U19419 (N_19419,N_17787,N_17670);
or U19420 (N_19420,N_16909,N_16207);
xnor U19421 (N_19421,N_17077,N_17224);
xnor U19422 (N_19422,N_17811,N_16045);
or U19423 (N_19423,N_17358,N_16324);
nor U19424 (N_19424,N_17962,N_17838);
or U19425 (N_19425,N_16358,N_16644);
or U19426 (N_19426,N_17376,N_16022);
nand U19427 (N_19427,N_16981,N_16992);
nand U19428 (N_19428,N_16321,N_16603);
and U19429 (N_19429,N_16574,N_16950);
nand U19430 (N_19430,N_17735,N_16490);
xor U19431 (N_19431,N_16767,N_16052);
nand U19432 (N_19432,N_16441,N_16188);
nor U19433 (N_19433,N_17438,N_17412);
xor U19434 (N_19434,N_17453,N_17582);
nand U19435 (N_19435,N_17721,N_17442);
and U19436 (N_19436,N_17582,N_16827);
or U19437 (N_19437,N_16941,N_17319);
and U19438 (N_19438,N_16587,N_16704);
nor U19439 (N_19439,N_17374,N_17556);
nor U19440 (N_19440,N_17250,N_16016);
nand U19441 (N_19441,N_17417,N_17051);
nand U19442 (N_19442,N_16474,N_16603);
xnor U19443 (N_19443,N_17393,N_17631);
nand U19444 (N_19444,N_16151,N_16692);
nor U19445 (N_19445,N_17652,N_17358);
nor U19446 (N_19446,N_17148,N_16898);
and U19447 (N_19447,N_16108,N_16936);
nand U19448 (N_19448,N_17027,N_16824);
nand U19449 (N_19449,N_17009,N_17998);
nor U19450 (N_19450,N_16709,N_16270);
nand U19451 (N_19451,N_17160,N_16329);
xnor U19452 (N_19452,N_16870,N_17898);
nor U19453 (N_19453,N_16122,N_16722);
nand U19454 (N_19454,N_17635,N_16476);
or U19455 (N_19455,N_16246,N_16924);
or U19456 (N_19456,N_16756,N_16129);
nor U19457 (N_19457,N_16909,N_17465);
nand U19458 (N_19458,N_16485,N_17119);
nand U19459 (N_19459,N_16455,N_17325);
or U19460 (N_19460,N_16528,N_17572);
xor U19461 (N_19461,N_17603,N_16293);
nand U19462 (N_19462,N_17608,N_16696);
nor U19463 (N_19463,N_17087,N_17682);
nor U19464 (N_19464,N_17721,N_16629);
nor U19465 (N_19465,N_17098,N_17993);
and U19466 (N_19466,N_16967,N_17918);
or U19467 (N_19467,N_16929,N_16060);
xnor U19468 (N_19468,N_16122,N_17167);
and U19469 (N_19469,N_16702,N_17952);
and U19470 (N_19470,N_16868,N_17471);
xnor U19471 (N_19471,N_17136,N_16015);
xor U19472 (N_19472,N_17626,N_16200);
or U19473 (N_19473,N_17148,N_17851);
nand U19474 (N_19474,N_17441,N_17538);
nor U19475 (N_19475,N_17353,N_17701);
nor U19476 (N_19476,N_16405,N_17292);
and U19477 (N_19477,N_17263,N_17501);
or U19478 (N_19478,N_17781,N_16060);
nand U19479 (N_19479,N_17670,N_17032);
nand U19480 (N_19480,N_17268,N_17136);
nand U19481 (N_19481,N_17898,N_17026);
xnor U19482 (N_19482,N_16283,N_17167);
and U19483 (N_19483,N_16598,N_17836);
nor U19484 (N_19484,N_16587,N_16996);
nand U19485 (N_19485,N_16528,N_17983);
or U19486 (N_19486,N_16793,N_16888);
or U19487 (N_19487,N_16411,N_16020);
nand U19488 (N_19488,N_16092,N_16665);
and U19489 (N_19489,N_16560,N_17431);
or U19490 (N_19490,N_16552,N_17848);
and U19491 (N_19491,N_16385,N_17849);
or U19492 (N_19492,N_16898,N_17487);
xnor U19493 (N_19493,N_17590,N_17338);
nand U19494 (N_19494,N_16522,N_16742);
xor U19495 (N_19495,N_17389,N_17883);
and U19496 (N_19496,N_17110,N_17807);
or U19497 (N_19497,N_17748,N_17466);
or U19498 (N_19498,N_17776,N_17938);
or U19499 (N_19499,N_17453,N_16451);
xnor U19500 (N_19500,N_17718,N_17097);
nor U19501 (N_19501,N_16255,N_16767);
xor U19502 (N_19502,N_17934,N_16741);
and U19503 (N_19503,N_17527,N_16537);
xor U19504 (N_19504,N_17475,N_17191);
and U19505 (N_19505,N_16261,N_17445);
xnor U19506 (N_19506,N_17050,N_17837);
nand U19507 (N_19507,N_16887,N_16572);
or U19508 (N_19508,N_16636,N_17792);
xnor U19509 (N_19509,N_17261,N_16052);
nand U19510 (N_19510,N_16075,N_16091);
nand U19511 (N_19511,N_16870,N_16110);
nor U19512 (N_19512,N_17915,N_17369);
nor U19513 (N_19513,N_16231,N_17209);
nand U19514 (N_19514,N_17822,N_17002);
and U19515 (N_19515,N_16783,N_17523);
xnor U19516 (N_19516,N_16127,N_17200);
and U19517 (N_19517,N_16701,N_17511);
or U19518 (N_19518,N_17941,N_17836);
nand U19519 (N_19519,N_17763,N_16266);
or U19520 (N_19520,N_16122,N_16260);
and U19521 (N_19521,N_16288,N_17238);
nand U19522 (N_19522,N_17281,N_16622);
and U19523 (N_19523,N_17705,N_17817);
or U19524 (N_19524,N_17563,N_16647);
nand U19525 (N_19525,N_16469,N_17223);
and U19526 (N_19526,N_17185,N_16169);
nand U19527 (N_19527,N_16091,N_17798);
nor U19528 (N_19528,N_16881,N_16600);
or U19529 (N_19529,N_17347,N_17005);
nor U19530 (N_19530,N_16118,N_17269);
and U19531 (N_19531,N_17386,N_16586);
nor U19532 (N_19532,N_17582,N_16808);
or U19533 (N_19533,N_16029,N_17768);
or U19534 (N_19534,N_17405,N_16889);
and U19535 (N_19535,N_16795,N_16300);
or U19536 (N_19536,N_16575,N_16586);
and U19537 (N_19537,N_16608,N_17643);
xnor U19538 (N_19538,N_17373,N_17479);
or U19539 (N_19539,N_16620,N_16664);
nor U19540 (N_19540,N_17830,N_17283);
nand U19541 (N_19541,N_16281,N_16058);
nor U19542 (N_19542,N_16273,N_17364);
xnor U19543 (N_19543,N_16780,N_16974);
xnor U19544 (N_19544,N_17435,N_16773);
nand U19545 (N_19545,N_16861,N_17633);
and U19546 (N_19546,N_16375,N_16598);
or U19547 (N_19547,N_16284,N_17860);
nand U19548 (N_19548,N_16526,N_17629);
xor U19549 (N_19549,N_17253,N_17538);
nand U19550 (N_19550,N_16271,N_16043);
nor U19551 (N_19551,N_17626,N_16789);
and U19552 (N_19552,N_17374,N_17642);
nand U19553 (N_19553,N_16518,N_17492);
and U19554 (N_19554,N_16286,N_16234);
nor U19555 (N_19555,N_17526,N_17647);
nor U19556 (N_19556,N_16169,N_16087);
and U19557 (N_19557,N_17850,N_17008);
nand U19558 (N_19558,N_16834,N_16238);
or U19559 (N_19559,N_16225,N_17718);
nand U19560 (N_19560,N_17253,N_17727);
and U19561 (N_19561,N_16600,N_17104);
or U19562 (N_19562,N_16911,N_17604);
or U19563 (N_19563,N_17637,N_17846);
and U19564 (N_19564,N_17321,N_17349);
nor U19565 (N_19565,N_16152,N_16537);
xnor U19566 (N_19566,N_17839,N_17210);
xnor U19567 (N_19567,N_16635,N_17258);
nor U19568 (N_19568,N_17495,N_16264);
xor U19569 (N_19569,N_17650,N_16779);
xnor U19570 (N_19570,N_17555,N_17459);
or U19571 (N_19571,N_17009,N_16869);
xnor U19572 (N_19572,N_17106,N_17843);
nor U19573 (N_19573,N_17727,N_16665);
xor U19574 (N_19574,N_16339,N_17171);
and U19575 (N_19575,N_16338,N_17911);
nor U19576 (N_19576,N_17029,N_17398);
xor U19577 (N_19577,N_17514,N_16415);
or U19578 (N_19578,N_17909,N_16945);
nand U19579 (N_19579,N_17133,N_17359);
nand U19580 (N_19580,N_16637,N_16729);
and U19581 (N_19581,N_16626,N_17639);
or U19582 (N_19582,N_16242,N_17143);
nand U19583 (N_19583,N_16359,N_16518);
xnor U19584 (N_19584,N_16114,N_16590);
nand U19585 (N_19585,N_16810,N_16979);
xnor U19586 (N_19586,N_16478,N_16967);
xnor U19587 (N_19587,N_16275,N_16840);
xor U19588 (N_19588,N_16298,N_16255);
xnor U19589 (N_19589,N_16696,N_17525);
and U19590 (N_19590,N_16093,N_16424);
nor U19591 (N_19591,N_16798,N_16731);
and U19592 (N_19592,N_16573,N_16521);
nor U19593 (N_19593,N_17830,N_16480);
and U19594 (N_19594,N_16239,N_17373);
or U19595 (N_19595,N_17944,N_17513);
and U19596 (N_19596,N_16733,N_17927);
and U19597 (N_19597,N_16279,N_17435);
nor U19598 (N_19598,N_17909,N_17919);
xor U19599 (N_19599,N_16526,N_17089);
xor U19600 (N_19600,N_17016,N_17554);
or U19601 (N_19601,N_16136,N_17403);
or U19602 (N_19602,N_17209,N_17816);
and U19603 (N_19603,N_16920,N_16367);
or U19604 (N_19604,N_17641,N_17030);
and U19605 (N_19605,N_17678,N_17728);
nor U19606 (N_19606,N_17595,N_16699);
xnor U19607 (N_19607,N_16315,N_16443);
xor U19608 (N_19608,N_16729,N_16576);
nor U19609 (N_19609,N_16168,N_17840);
nand U19610 (N_19610,N_16659,N_16653);
or U19611 (N_19611,N_16758,N_16451);
and U19612 (N_19612,N_16933,N_17181);
or U19613 (N_19613,N_17799,N_16814);
nor U19614 (N_19614,N_17135,N_16574);
or U19615 (N_19615,N_16073,N_17930);
nor U19616 (N_19616,N_16799,N_16060);
and U19617 (N_19617,N_16621,N_16940);
and U19618 (N_19618,N_16869,N_16909);
and U19619 (N_19619,N_17297,N_16819);
and U19620 (N_19620,N_17656,N_17048);
and U19621 (N_19621,N_16057,N_17383);
nor U19622 (N_19622,N_17954,N_17860);
nand U19623 (N_19623,N_17979,N_16258);
and U19624 (N_19624,N_17799,N_17123);
or U19625 (N_19625,N_17021,N_16184);
xnor U19626 (N_19626,N_16804,N_16760);
or U19627 (N_19627,N_17680,N_16655);
nand U19628 (N_19628,N_17614,N_16127);
nand U19629 (N_19629,N_17090,N_17395);
nor U19630 (N_19630,N_16489,N_16989);
nor U19631 (N_19631,N_17645,N_17633);
and U19632 (N_19632,N_17119,N_17944);
or U19633 (N_19633,N_17567,N_16302);
or U19634 (N_19634,N_16384,N_17075);
nor U19635 (N_19635,N_16941,N_17016);
xnor U19636 (N_19636,N_17962,N_16022);
and U19637 (N_19637,N_17177,N_17512);
or U19638 (N_19638,N_16025,N_16824);
nor U19639 (N_19639,N_17758,N_17407);
and U19640 (N_19640,N_16095,N_17142);
or U19641 (N_19641,N_17417,N_16009);
xnor U19642 (N_19642,N_17562,N_17399);
nor U19643 (N_19643,N_16692,N_17155);
xor U19644 (N_19644,N_16338,N_16189);
nand U19645 (N_19645,N_16804,N_17671);
nand U19646 (N_19646,N_17947,N_17909);
xor U19647 (N_19647,N_17289,N_17171);
or U19648 (N_19648,N_17090,N_16121);
and U19649 (N_19649,N_16262,N_16636);
and U19650 (N_19650,N_16409,N_16359);
xnor U19651 (N_19651,N_16492,N_17963);
nand U19652 (N_19652,N_17516,N_16429);
and U19653 (N_19653,N_16923,N_16191);
nor U19654 (N_19654,N_16470,N_17183);
xnor U19655 (N_19655,N_16387,N_17466);
nor U19656 (N_19656,N_17437,N_17096);
xor U19657 (N_19657,N_16450,N_16228);
xnor U19658 (N_19658,N_17866,N_16817);
nand U19659 (N_19659,N_17639,N_17851);
or U19660 (N_19660,N_17036,N_17855);
or U19661 (N_19661,N_17173,N_16431);
nand U19662 (N_19662,N_16040,N_16334);
nor U19663 (N_19663,N_17327,N_16028);
xnor U19664 (N_19664,N_17141,N_17159);
nor U19665 (N_19665,N_16660,N_16928);
nor U19666 (N_19666,N_16358,N_17666);
and U19667 (N_19667,N_17429,N_17327);
nor U19668 (N_19668,N_17775,N_16044);
or U19669 (N_19669,N_17957,N_16193);
or U19670 (N_19670,N_16693,N_16742);
and U19671 (N_19671,N_16061,N_16178);
nand U19672 (N_19672,N_17902,N_16840);
or U19673 (N_19673,N_17608,N_17917);
or U19674 (N_19674,N_17548,N_16820);
nand U19675 (N_19675,N_17636,N_17232);
or U19676 (N_19676,N_17986,N_16395);
nor U19677 (N_19677,N_16118,N_16325);
and U19678 (N_19678,N_17662,N_16789);
nor U19679 (N_19679,N_16115,N_17925);
xor U19680 (N_19680,N_17020,N_16414);
or U19681 (N_19681,N_16690,N_17829);
xor U19682 (N_19682,N_16645,N_16084);
and U19683 (N_19683,N_17072,N_17557);
and U19684 (N_19684,N_16999,N_16049);
or U19685 (N_19685,N_17746,N_16878);
nand U19686 (N_19686,N_17098,N_16801);
or U19687 (N_19687,N_16111,N_17584);
nor U19688 (N_19688,N_17791,N_17563);
nand U19689 (N_19689,N_17069,N_16466);
nand U19690 (N_19690,N_16368,N_17512);
and U19691 (N_19691,N_16477,N_16599);
or U19692 (N_19692,N_17592,N_16833);
or U19693 (N_19693,N_17985,N_16969);
nor U19694 (N_19694,N_16248,N_17644);
nand U19695 (N_19695,N_16001,N_17399);
or U19696 (N_19696,N_17770,N_16204);
nand U19697 (N_19697,N_16456,N_17804);
nor U19698 (N_19698,N_17558,N_16331);
or U19699 (N_19699,N_17308,N_17515);
nand U19700 (N_19700,N_16651,N_16077);
and U19701 (N_19701,N_16258,N_17045);
or U19702 (N_19702,N_17434,N_16107);
nor U19703 (N_19703,N_16519,N_16419);
xor U19704 (N_19704,N_17548,N_16098);
and U19705 (N_19705,N_16362,N_16219);
and U19706 (N_19706,N_17106,N_16988);
nand U19707 (N_19707,N_17193,N_16761);
or U19708 (N_19708,N_17349,N_16318);
and U19709 (N_19709,N_16518,N_16347);
or U19710 (N_19710,N_16359,N_17310);
xnor U19711 (N_19711,N_17683,N_16209);
and U19712 (N_19712,N_17684,N_16091);
nand U19713 (N_19713,N_16874,N_17875);
nand U19714 (N_19714,N_17831,N_17776);
and U19715 (N_19715,N_17009,N_17700);
and U19716 (N_19716,N_16145,N_17500);
or U19717 (N_19717,N_17948,N_16100);
and U19718 (N_19718,N_16299,N_16890);
and U19719 (N_19719,N_17166,N_17975);
xor U19720 (N_19720,N_16707,N_17808);
nand U19721 (N_19721,N_16032,N_16571);
or U19722 (N_19722,N_17717,N_16995);
nor U19723 (N_19723,N_17013,N_17456);
nand U19724 (N_19724,N_17574,N_16508);
nor U19725 (N_19725,N_17333,N_16335);
nor U19726 (N_19726,N_16083,N_16344);
and U19727 (N_19727,N_16400,N_16523);
nand U19728 (N_19728,N_16418,N_17202);
or U19729 (N_19729,N_17495,N_16005);
and U19730 (N_19730,N_16424,N_16443);
and U19731 (N_19731,N_17912,N_17449);
or U19732 (N_19732,N_16310,N_17397);
nor U19733 (N_19733,N_16570,N_16773);
nor U19734 (N_19734,N_16028,N_17509);
or U19735 (N_19735,N_16169,N_17040);
nor U19736 (N_19736,N_16499,N_17862);
or U19737 (N_19737,N_16853,N_17212);
nor U19738 (N_19738,N_17080,N_16017);
nor U19739 (N_19739,N_16280,N_16835);
or U19740 (N_19740,N_16309,N_17491);
xnor U19741 (N_19741,N_17943,N_17482);
nor U19742 (N_19742,N_16132,N_17913);
nand U19743 (N_19743,N_17898,N_17421);
nand U19744 (N_19744,N_16987,N_16903);
nand U19745 (N_19745,N_16247,N_17908);
nor U19746 (N_19746,N_16083,N_17011);
nand U19747 (N_19747,N_16996,N_16174);
or U19748 (N_19748,N_16662,N_17859);
nand U19749 (N_19749,N_17343,N_16101);
nor U19750 (N_19750,N_17331,N_16296);
nand U19751 (N_19751,N_16519,N_17830);
xnor U19752 (N_19752,N_17136,N_17121);
or U19753 (N_19753,N_16702,N_17117);
nor U19754 (N_19754,N_16127,N_17243);
xor U19755 (N_19755,N_17188,N_17534);
nand U19756 (N_19756,N_16751,N_17113);
xor U19757 (N_19757,N_17974,N_16183);
or U19758 (N_19758,N_17971,N_17857);
and U19759 (N_19759,N_16487,N_16331);
xnor U19760 (N_19760,N_17964,N_16325);
or U19761 (N_19761,N_16599,N_17298);
xnor U19762 (N_19762,N_16651,N_16081);
nand U19763 (N_19763,N_16391,N_17957);
or U19764 (N_19764,N_16881,N_17517);
nand U19765 (N_19765,N_17659,N_17854);
nand U19766 (N_19766,N_17298,N_17700);
nand U19767 (N_19767,N_17398,N_16716);
nor U19768 (N_19768,N_17960,N_17035);
nor U19769 (N_19769,N_16909,N_16623);
nand U19770 (N_19770,N_16413,N_17510);
nor U19771 (N_19771,N_16510,N_17021);
nor U19772 (N_19772,N_16571,N_16587);
and U19773 (N_19773,N_16362,N_17128);
xnor U19774 (N_19774,N_17136,N_16322);
nand U19775 (N_19775,N_16109,N_16414);
or U19776 (N_19776,N_17989,N_16107);
and U19777 (N_19777,N_16618,N_17692);
xnor U19778 (N_19778,N_16348,N_17348);
xor U19779 (N_19779,N_16515,N_16566);
nand U19780 (N_19780,N_16377,N_17149);
nand U19781 (N_19781,N_17410,N_17227);
xnor U19782 (N_19782,N_17003,N_17721);
nor U19783 (N_19783,N_17310,N_16244);
xor U19784 (N_19784,N_17507,N_17076);
xor U19785 (N_19785,N_17901,N_16230);
xor U19786 (N_19786,N_16429,N_16607);
and U19787 (N_19787,N_17618,N_17632);
and U19788 (N_19788,N_16176,N_16252);
nand U19789 (N_19789,N_16322,N_16666);
or U19790 (N_19790,N_16999,N_17220);
nor U19791 (N_19791,N_17714,N_17821);
xnor U19792 (N_19792,N_17292,N_16412);
nand U19793 (N_19793,N_16679,N_16155);
xor U19794 (N_19794,N_16149,N_16175);
xnor U19795 (N_19795,N_17224,N_16163);
or U19796 (N_19796,N_16154,N_17429);
xor U19797 (N_19797,N_17740,N_17835);
nor U19798 (N_19798,N_17375,N_17393);
or U19799 (N_19799,N_17034,N_17964);
xnor U19800 (N_19800,N_16587,N_16480);
or U19801 (N_19801,N_17425,N_16004);
xor U19802 (N_19802,N_17155,N_16782);
and U19803 (N_19803,N_16103,N_17345);
xor U19804 (N_19804,N_17683,N_16007);
or U19805 (N_19805,N_17637,N_16548);
nand U19806 (N_19806,N_17963,N_17906);
xnor U19807 (N_19807,N_17645,N_17160);
and U19808 (N_19808,N_16518,N_16314);
xor U19809 (N_19809,N_16462,N_16480);
xor U19810 (N_19810,N_17677,N_17986);
nand U19811 (N_19811,N_16135,N_16817);
xnor U19812 (N_19812,N_16643,N_16438);
nand U19813 (N_19813,N_16961,N_16675);
nand U19814 (N_19814,N_16477,N_16680);
xor U19815 (N_19815,N_17035,N_17057);
nor U19816 (N_19816,N_16499,N_16913);
nand U19817 (N_19817,N_16327,N_16016);
xnor U19818 (N_19818,N_17936,N_17793);
nor U19819 (N_19819,N_16566,N_16810);
and U19820 (N_19820,N_17206,N_17338);
nor U19821 (N_19821,N_17163,N_16190);
and U19822 (N_19822,N_16685,N_17566);
nand U19823 (N_19823,N_17142,N_17022);
xor U19824 (N_19824,N_16663,N_16826);
and U19825 (N_19825,N_17540,N_17047);
and U19826 (N_19826,N_17561,N_16167);
and U19827 (N_19827,N_17708,N_17660);
and U19828 (N_19828,N_17892,N_17835);
nor U19829 (N_19829,N_16613,N_16459);
nand U19830 (N_19830,N_17401,N_16683);
or U19831 (N_19831,N_16424,N_16962);
or U19832 (N_19832,N_17798,N_17032);
nand U19833 (N_19833,N_16074,N_16878);
and U19834 (N_19834,N_17972,N_16470);
nor U19835 (N_19835,N_16757,N_17332);
and U19836 (N_19836,N_17901,N_17260);
or U19837 (N_19837,N_17455,N_16907);
and U19838 (N_19838,N_17302,N_16030);
and U19839 (N_19839,N_16899,N_17342);
or U19840 (N_19840,N_16170,N_16891);
nand U19841 (N_19841,N_16441,N_17194);
nand U19842 (N_19842,N_17906,N_17493);
and U19843 (N_19843,N_17114,N_16129);
and U19844 (N_19844,N_16876,N_16297);
and U19845 (N_19845,N_17245,N_16555);
nor U19846 (N_19846,N_16331,N_17252);
nor U19847 (N_19847,N_17289,N_17566);
nor U19848 (N_19848,N_16063,N_16032);
and U19849 (N_19849,N_16488,N_17645);
nor U19850 (N_19850,N_16673,N_17789);
nand U19851 (N_19851,N_16431,N_16758);
and U19852 (N_19852,N_17254,N_16365);
and U19853 (N_19853,N_17810,N_16205);
nor U19854 (N_19854,N_17281,N_16307);
nand U19855 (N_19855,N_16790,N_16928);
nor U19856 (N_19856,N_17631,N_16932);
and U19857 (N_19857,N_16292,N_17365);
nor U19858 (N_19858,N_16783,N_17131);
or U19859 (N_19859,N_16521,N_16741);
or U19860 (N_19860,N_17399,N_16722);
xor U19861 (N_19861,N_16386,N_17781);
or U19862 (N_19862,N_17544,N_17120);
xnor U19863 (N_19863,N_16866,N_17641);
nor U19864 (N_19864,N_16892,N_17206);
and U19865 (N_19865,N_17935,N_17888);
nor U19866 (N_19866,N_16106,N_16770);
nand U19867 (N_19867,N_17721,N_16195);
nand U19868 (N_19868,N_16665,N_17769);
nand U19869 (N_19869,N_17341,N_17855);
xor U19870 (N_19870,N_17188,N_16915);
and U19871 (N_19871,N_16854,N_17860);
and U19872 (N_19872,N_17556,N_16710);
nor U19873 (N_19873,N_16852,N_17926);
xnor U19874 (N_19874,N_17169,N_16536);
or U19875 (N_19875,N_17102,N_16893);
or U19876 (N_19876,N_17141,N_17955);
nand U19877 (N_19877,N_16207,N_16873);
nor U19878 (N_19878,N_16886,N_16665);
and U19879 (N_19879,N_17273,N_16611);
or U19880 (N_19880,N_17562,N_17012);
and U19881 (N_19881,N_17967,N_16487);
or U19882 (N_19882,N_17483,N_17016);
xor U19883 (N_19883,N_16228,N_16568);
and U19884 (N_19884,N_16790,N_17188);
or U19885 (N_19885,N_16611,N_16004);
or U19886 (N_19886,N_16942,N_16668);
nor U19887 (N_19887,N_17582,N_16277);
or U19888 (N_19888,N_16695,N_16072);
or U19889 (N_19889,N_17367,N_16759);
xor U19890 (N_19890,N_17506,N_16848);
and U19891 (N_19891,N_16640,N_16574);
nand U19892 (N_19892,N_16215,N_17000);
xor U19893 (N_19893,N_16663,N_16561);
nor U19894 (N_19894,N_17398,N_16291);
nand U19895 (N_19895,N_17654,N_17265);
and U19896 (N_19896,N_16519,N_16303);
nand U19897 (N_19897,N_17552,N_16647);
xnor U19898 (N_19898,N_16708,N_16028);
xnor U19899 (N_19899,N_16946,N_17197);
nand U19900 (N_19900,N_17227,N_17959);
or U19901 (N_19901,N_16806,N_17828);
or U19902 (N_19902,N_17378,N_17245);
and U19903 (N_19903,N_16983,N_17054);
xnor U19904 (N_19904,N_16143,N_17085);
and U19905 (N_19905,N_17521,N_16560);
nor U19906 (N_19906,N_16530,N_17469);
and U19907 (N_19907,N_17045,N_16163);
and U19908 (N_19908,N_17249,N_16286);
xor U19909 (N_19909,N_17528,N_17188);
xor U19910 (N_19910,N_17957,N_17339);
or U19911 (N_19911,N_17593,N_16962);
and U19912 (N_19912,N_16615,N_16562);
or U19913 (N_19913,N_16252,N_17864);
nor U19914 (N_19914,N_16175,N_16762);
or U19915 (N_19915,N_16045,N_17918);
or U19916 (N_19916,N_17726,N_17555);
xor U19917 (N_19917,N_16692,N_17848);
or U19918 (N_19918,N_17965,N_17048);
and U19919 (N_19919,N_17471,N_16134);
nor U19920 (N_19920,N_16630,N_16418);
or U19921 (N_19921,N_16533,N_16356);
and U19922 (N_19922,N_16349,N_16835);
or U19923 (N_19923,N_16820,N_16323);
and U19924 (N_19924,N_16513,N_16985);
nand U19925 (N_19925,N_16831,N_17266);
or U19926 (N_19926,N_17533,N_16870);
nand U19927 (N_19927,N_16088,N_17357);
nor U19928 (N_19928,N_17379,N_16958);
and U19929 (N_19929,N_17057,N_16809);
and U19930 (N_19930,N_17975,N_17990);
xor U19931 (N_19931,N_17424,N_17680);
or U19932 (N_19932,N_16232,N_17105);
nor U19933 (N_19933,N_17915,N_17473);
nand U19934 (N_19934,N_16862,N_16311);
xor U19935 (N_19935,N_16986,N_16187);
xor U19936 (N_19936,N_16576,N_16836);
xnor U19937 (N_19937,N_17468,N_17919);
nor U19938 (N_19938,N_16230,N_16933);
and U19939 (N_19939,N_17997,N_17774);
and U19940 (N_19940,N_16925,N_16429);
nor U19941 (N_19941,N_16243,N_17115);
nand U19942 (N_19942,N_17910,N_17300);
and U19943 (N_19943,N_16163,N_17268);
xnor U19944 (N_19944,N_17071,N_16379);
nand U19945 (N_19945,N_16334,N_17164);
xor U19946 (N_19946,N_16168,N_16501);
and U19947 (N_19947,N_16791,N_17601);
or U19948 (N_19948,N_16374,N_16911);
or U19949 (N_19949,N_17496,N_17306);
xnor U19950 (N_19950,N_17553,N_17524);
or U19951 (N_19951,N_17007,N_16267);
and U19952 (N_19952,N_17039,N_16669);
nor U19953 (N_19953,N_17755,N_17915);
xnor U19954 (N_19954,N_16542,N_17411);
xor U19955 (N_19955,N_17823,N_17014);
xnor U19956 (N_19956,N_17844,N_16841);
xnor U19957 (N_19957,N_17681,N_17840);
nand U19958 (N_19958,N_16125,N_17351);
xnor U19959 (N_19959,N_16839,N_16853);
and U19960 (N_19960,N_17926,N_17588);
and U19961 (N_19961,N_16415,N_17500);
or U19962 (N_19962,N_17504,N_17495);
and U19963 (N_19963,N_16670,N_16067);
or U19964 (N_19964,N_16914,N_16992);
and U19965 (N_19965,N_17745,N_16808);
xnor U19966 (N_19966,N_17668,N_16381);
or U19967 (N_19967,N_16920,N_17363);
or U19968 (N_19968,N_17056,N_16098);
nor U19969 (N_19969,N_17685,N_16609);
and U19970 (N_19970,N_16163,N_16745);
nand U19971 (N_19971,N_17230,N_17118);
nor U19972 (N_19972,N_16598,N_17414);
or U19973 (N_19973,N_16152,N_17454);
or U19974 (N_19974,N_17609,N_17641);
xnor U19975 (N_19975,N_17358,N_16714);
xnor U19976 (N_19976,N_16132,N_17802);
and U19977 (N_19977,N_17101,N_17345);
xnor U19978 (N_19978,N_16697,N_16446);
xnor U19979 (N_19979,N_16902,N_16940);
or U19980 (N_19980,N_17837,N_16903);
xnor U19981 (N_19981,N_17064,N_17737);
or U19982 (N_19982,N_17808,N_17369);
or U19983 (N_19983,N_17783,N_17132);
or U19984 (N_19984,N_16650,N_16253);
xnor U19985 (N_19985,N_16466,N_17872);
nor U19986 (N_19986,N_17810,N_16960);
nand U19987 (N_19987,N_16499,N_16276);
xnor U19988 (N_19988,N_16212,N_17178);
or U19989 (N_19989,N_16894,N_16831);
nand U19990 (N_19990,N_17053,N_17525);
nor U19991 (N_19991,N_17824,N_16776);
or U19992 (N_19992,N_16571,N_16580);
or U19993 (N_19993,N_16923,N_16414);
xor U19994 (N_19994,N_16189,N_17200);
nand U19995 (N_19995,N_16226,N_16909);
nor U19996 (N_19996,N_16643,N_17444);
and U19997 (N_19997,N_16595,N_17268);
nor U19998 (N_19998,N_17875,N_16683);
and U19999 (N_19999,N_16511,N_16117);
nand UO_0 (O_0,N_18430,N_19334);
nor UO_1 (O_1,N_19363,N_19656);
nor UO_2 (O_2,N_19103,N_19234);
nor UO_3 (O_3,N_19862,N_19383);
and UO_4 (O_4,N_19875,N_19901);
nand UO_5 (O_5,N_18402,N_19066);
xor UO_6 (O_6,N_18498,N_18306);
xnor UO_7 (O_7,N_19172,N_19518);
nor UO_8 (O_8,N_18477,N_18852);
or UO_9 (O_9,N_19540,N_19184);
or UO_10 (O_10,N_18684,N_18273);
and UO_11 (O_11,N_19799,N_19134);
nand UO_12 (O_12,N_19028,N_19398);
nor UO_13 (O_13,N_19484,N_19240);
xnor UO_14 (O_14,N_19098,N_18123);
xor UO_15 (O_15,N_19128,N_18815);
and UO_16 (O_16,N_19960,N_19824);
nor UO_17 (O_17,N_18576,N_18292);
and UO_18 (O_18,N_19507,N_19769);
nor UO_19 (O_19,N_18235,N_18893);
nand UO_20 (O_20,N_18189,N_19267);
xor UO_21 (O_21,N_18848,N_18475);
nand UO_22 (O_22,N_18332,N_19084);
nand UO_23 (O_23,N_18249,N_19569);
nand UO_24 (O_24,N_19372,N_18958);
xor UO_25 (O_25,N_19132,N_18964);
nor UO_26 (O_26,N_18146,N_19091);
nor UO_27 (O_27,N_19967,N_18379);
and UO_28 (O_28,N_18347,N_18462);
xor UO_29 (O_29,N_19150,N_19986);
xor UO_30 (O_30,N_18471,N_18868);
xnor UO_31 (O_31,N_19116,N_19972);
xnor UO_32 (O_32,N_19539,N_19852);
and UO_33 (O_33,N_18043,N_18880);
or UO_34 (O_34,N_19635,N_19042);
and UO_35 (O_35,N_19965,N_19629);
nand UO_36 (O_36,N_18951,N_19056);
xor UO_37 (O_37,N_19472,N_19532);
and UO_38 (O_38,N_18522,N_19726);
nor UO_39 (O_39,N_19316,N_18083);
nor UO_40 (O_40,N_18205,N_18225);
or UO_41 (O_41,N_18198,N_18048);
or UO_42 (O_42,N_19941,N_19191);
xnor UO_43 (O_43,N_19082,N_19711);
xnor UO_44 (O_44,N_19074,N_19996);
xor UO_45 (O_45,N_18391,N_19812);
nor UO_46 (O_46,N_19493,N_19789);
and UO_47 (O_47,N_18119,N_18765);
nand UO_48 (O_48,N_19307,N_19955);
xor UO_49 (O_49,N_18851,N_18406);
xnor UO_50 (O_50,N_18436,N_18542);
xor UO_51 (O_51,N_18137,N_18841);
xor UO_52 (O_52,N_18238,N_18375);
nand UO_53 (O_53,N_18535,N_19898);
and UO_54 (O_54,N_18905,N_18788);
xnor UO_55 (O_55,N_18835,N_18267);
and UO_56 (O_56,N_18827,N_18661);
nor UO_57 (O_57,N_19974,N_18156);
or UO_58 (O_58,N_19554,N_19110);
and UO_59 (O_59,N_19956,N_18323);
or UO_60 (O_60,N_18658,N_19089);
and UO_61 (O_61,N_18762,N_18534);
or UO_62 (O_62,N_19429,N_19130);
nor UO_63 (O_63,N_19449,N_18387);
nor UO_64 (O_64,N_18381,N_18555);
or UO_65 (O_65,N_19672,N_19969);
or UO_66 (O_66,N_18586,N_19529);
or UO_67 (O_67,N_19431,N_18473);
or UO_68 (O_68,N_19460,N_19886);
xnor UO_69 (O_69,N_18989,N_18007);
or UO_70 (O_70,N_19464,N_19676);
or UO_71 (O_71,N_19271,N_18843);
and UO_72 (O_72,N_18277,N_19229);
nand UO_73 (O_73,N_19508,N_19728);
nand UO_74 (O_74,N_18429,N_19077);
nor UO_75 (O_75,N_18701,N_19800);
xor UO_76 (O_76,N_18029,N_18897);
xnor UO_77 (O_77,N_19805,N_19818);
xnor UO_78 (O_78,N_18833,N_19264);
or UO_79 (O_79,N_18260,N_19205);
or UO_80 (O_80,N_18398,N_19669);
nor UO_81 (O_81,N_18264,N_19325);
and UO_82 (O_82,N_19285,N_18960);
and UO_83 (O_83,N_18045,N_19198);
nand UO_84 (O_84,N_19823,N_18871);
or UO_85 (O_85,N_19722,N_18840);
nand UO_86 (O_86,N_19081,N_19725);
and UO_87 (O_87,N_19147,N_18676);
xnor UO_88 (O_88,N_19262,N_18923);
nor UO_89 (O_89,N_19458,N_18806);
xor UO_90 (O_90,N_19490,N_18112);
nor UO_91 (O_91,N_19641,N_18920);
nand UO_92 (O_92,N_19739,N_19139);
or UO_93 (O_93,N_18521,N_19144);
nand UO_94 (O_94,N_18500,N_18335);
and UO_95 (O_95,N_19156,N_19872);
and UO_96 (O_96,N_19697,N_18506);
and UO_97 (O_97,N_18179,N_18180);
or UO_98 (O_98,N_19282,N_19442);
or UO_99 (O_99,N_18867,N_19837);
xor UO_100 (O_100,N_19002,N_18824);
nand UO_101 (O_101,N_18554,N_18499);
nand UO_102 (O_102,N_18305,N_19520);
nor UO_103 (O_103,N_18129,N_18977);
and UO_104 (O_104,N_19470,N_19807);
and UO_105 (O_105,N_19581,N_18731);
xnor UO_106 (O_106,N_19021,N_19806);
or UO_107 (O_107,N_18503,N_18927);
or UO_108 (O_108,N_19051,N_19162);
and UO_109 (O_109,N_19222,N_19698);
nor UO_110 (O_110,N_18875,N_18283);
nand UO_111 (O_111,N_18364,N_19369);
xnor UO_112 (O_112,N_19256,N_19375);
and UO_113 (O_113,N_18314,N_18589);
or UO_114 (O_114,N_19045,N_18693);
xor UO_115 (O_115,N_18890,N_19757);
nor UO_116 (O_116,N_18177,N_18370);
nor UO_117 (O_117,N_18312,N_18326);
or UO_118 (O_118,N_19583,N_19292);
xor UO_119 (O_119,N_18215,N_18024);
xor UO_120 (O_120,N_19311,N_19984);
xor UO_121 (O_121,N_18405,N_18208);
nand UO_122 (O_122,N_18467,N_19519);
xnor UO_123 (O_123,N_19916,N_18072);
or UO_124 (O_124,N_19025,N_19122);
or UO_125 (O_125,N_19171,N_19315);
or UO_126 (O_126,N_18207,N_18345);
nand UO_127 (O_127,N_18549,N_19489);
or UO_128 (O_128,N_18751,N_18294);
nand UO_129 (O_129,N_18466,N_18226);
nand UO_130 (O_130,N_19500,N_18584);
or UO_131 (O_131,N_18799,N_19513);
nor UO_132 (O_132,N_18154,N_19186);
xnor UO_133 (O_133,N_18708,N_19621);
xor UO_134 (O_134,N_18056,N_18607);
nor UO_135 (O_135,N_18265,N_18114);
or UO_136 (O_136,N_18758,N_19913);
nand UO_137 (O_137,N_19743,N_19269);
xnor UO_138 (O_138,N_19250,N_18970);
nor UO_139 (O_139,N_19439,N_19578);
or UO_140 (O_140,N_19868,N_19276);
nand UO_141 (O_141,N_19330,N_19355);
and UO_142 (O_142,N_19284,N_18076);
nand UO_143 (O_143,N_18856,N_19708);
nand UO_144 (O_144,N_19925,N_18930);
and UO_145 (O_145,N_19339,N_18702);
nor UO_146 (O_146,N_19000,N_19653);
nand UO_147 (O_147,N_19067,N_18057);
and UO_148 (O_148,N_19290,N_18211);
or UO_149 (O_149,N_18313,N_18626);
nand UO_150 (O_150,N_18178,N_19005);
and UO_151 (O_151,N_18540,N_18010);
or UO_152 (O_152,N_18165,N_19195);
xor UO_153 (O_153,N_18849,N_18117);
nand UO_154 (O_154,N_18531,N_18132);
or UO_155 (O_155,N_18735,N_18120);
or UO_156 (O_156,N_18094,N_19814);
xnor UO_157 (O_157,N_18968,N_19384);
xor UO_158 (O_158,N_19196,N_18403);
xor UO_159 (O_159,N_19336,N_18630);
xnor UO_160 (O_160,N_18293,N_18931);
or UO_161 (O_161,N_19504,N_19762);
or UO_162 (O_162,N_19437,N_19740);
nand UO_163 (O_163,N_18530,N_18081);
or UO_164 (O_164,N_18176,N_18459);
nor UO_165 (O_165,N_19877,N_18289);
xor UO_166 (O_166,N_18243,N_19060);
or UO_167 (O_167,N_18809,N_19933);
and UO_168 (O_168,N_18750,N_18606);
xor UO_169 (O_169,N_19286,N_18122);
and UO_170 (O_170,N_18910,N_19945);
xnor UO_171 (O_171,N_18357,N_18270);
and UO_172 (O_172,N_19623,N_18796);
nand UO_173 (O_173,N_18073,N_18533);
and UO_174 (O_174,N_19750,N_19367);
nand UO_175 (O_175,N_19395,N_18124);
or UO_176 (O_176,N_18690,N_18965);
xor UO_177 (O_177,N_19561,N_18173);
and UO_178 (O_178,N_19609,N_18934);
nand UO_179 (O_179,N_19280,N_18358);
xor UO_180 (O_180,N_18792,N_18526);
and UO_181 (O_181,N_18618,N_18109);
nor UO_182 (O_182,N_19839,N_19527);
or UO_183 (O_183,N_19380,N_18649);
or UO_184 (O_184,N_19415,N_18947);
and UO_185 (O_185,N_19982,N_18746);
and UO_186 (O_186,N_19924,N_19552);
xor UO_187 (O_187,N_19987,N_19608);
or UO_188 (O_188,N_19009,N_19037);
and UO_189 (O_189,N_18150,N_18756);
xnor UO_190 (O_190,N_19727,N_19895);
nor UO_191 (O_191,N_19085,N_19700);
xnor UO_192 (O_192,N_19246,N_19374);
xor UO_193 (O_193,N_18084,N_19188);
and UO_194 (O_194,N_19461,N_19140);
nand UO_195 (O_195,N_19345,N_18866);
nand UO_196 (O_196,N_18383,N_19633);
nor UO_197 (O_197,N_19248,N_18008);
and UO_198 (O_198,N_19602,N_18166);
nand UO_199 (O_199,N_18610,N_18494);
nor UO_200 (O_200,N_18884,N_18497);
nand UO_201 (O_201,N_18573,N_19289);
nor UO_202 (O_202,N_19764,N_19109);
xor UO_203 (O_203,N_19801,N_19036);
nand UO_204 (O_204,N_18662,N_18911);
or UO_205 (O_205,N_18537,N_19228);
and UO_206 (O_206,N_18703,N_19619);
nor UO_207 (O_207,N_18898,N_19644);
and UO_208 (O_208,N_18737,N_19971);
nand UO_209 (O_209,N_19120,N_19253);
nor UO_210 (O_210,N_18571,N_19494);
xnor UO_211 (O_211,N_18087,N_19879);
nor UO_212 (O_212,N_18206,N_18128);
or UO_213 (O_213,N_19911,N_19610);
or UO_214 (O_214,N_18134,N_19366);
and UO_215 (O_215,N_18985,N_18722);
xnor UO_216 (O_216,N_19381,N_18419);
xor UO_217 (O_217,N_19491,N_18447);
nor UO_218 (O_218,N_19255,N_19591);
xnor UO_219 (O_219,N_19317,N_19101);
nor UO_220 (O_220,N_18975,N_19358);
xnor UO_221 (O_221,N_18052,N_18183);
nand UO_222 (O_222,N_19534,N_19294);
xor UO_223 (O_223,N_19571,N_18603);
xnor UO_224 (O_224,N_18449,N_18636);
or UO_225 (O_225,N_18850,N_18304);
or UO_226 (O_226,N_19869,N_18797);
or UO_227 (O_227,N_18331,N_18940);
or UO_228 (O_228,N_19303,N_19840);
xnor UO_229 (O_229,N_19850,N_19843);
xnor UO_230 (O_230,N_18049,N_18980);
or UO_231 (O_231,N_18953,N_19048);
or UO_232 (O_232,N_19141,N_18042);
nor UO_233 (O_233,N_18480,N_19704);
nand UO_234 (O_234,N_18817,N_18291);
nor UO_235 (O_235,N_18786,N_18286);
and UO_236 (O_236,N_19992,N_19594);
nand UO_237 (O_237,N_19121,N_18779);
or UO_238 (O_238,N_18212,N_19861);
nor UO_239 (O_239,N_18365,N_18807);
xor UO_240 (O_240,N_19997,N_18111);
nor UO_241 (O_241,N_19176,N_18425);
xnor UO_242 (O_242,N_19792,N_19064);
nand UO_243 (O_243,N_18559,N_19390);
nor UO_244 (O_244,N_19846,N_19158);
xor UO_245 (O_245,N_18517,N_19018);
xor UO_246 (O_246,N_18030,N_18064);
and UO_247 (O_247,N_19313,N_19667);
and UO_248 (O_248,N_18316,N_18869);
nand UO_249 (O_249,N_19001,N_18151);
or UO_250 (O_250,N_18719,N_19133);
xor UO_251 (O_251,N_19734,N_18669);
and UO_252 (O_252,N_18632,N_18268);
nand UO_253 (O_253,N_19453,N_19268);
nand UO_254 (O_254,N_19553,N_18168);
or UO_255 (O_255,N_18925,N_18664);
or UO_256 (O_256,N_18214,N_18681);
and UO_257 (O_257,N_18857,N_18445);
nand UO_258 (O_258,N_19293,N_18752);
and UO_259 (O_259,N_19994,N_18655);
and UO_260 (O_260,N_18993,N_18432);
xnor UO_261 (O_261,N_18278,N_18638);
nor UO_262 (O_262,N_18899,N_18245);
nor UO_263 (O_263,N_18718,N_19499);
nand UO_264 (O_264,N_19220,N_19881);
or UO_265 (O_265,N_18538,N_19153);
and UO_266 (O_266,N_19265,N_19017);
or UO_267 (O_267,N_19832,N_19498);
nor UO_268 (O_268,N_18768,N_18546);
nor UO_269 (O_269,N_19679,N_18067);
and UO_270 (O_270,N_18006,N_19396);
and UO_271 (O_271,N_19995,N_19486);
nor UO_272 (O_272,N_18232,N_18290);
and UO_273 (O_273,N_18074,N_19406);
or UO_274 (O_274,N_18219,N_18650);
and UO_275 (O_275,N_19811,N_18580);
nand UO_276 (O_276,N_19346,N_19146);
or UO_277 (O_277,N_19607,N_18320);
or UO_278 (O_278,N_18324,N_19209);
nor UO_279 (O_279,N_18747,N_19076);
nand UO_280 (O_280,N_19838,N_18213);
xnor UO_281 (O_281,N_19546,N_18574);
nand UO_282 (O_282,N_18593,N_18680);
or UO_283 (O_283,N_19517,N_18368);
xnor UO_284 (O_284,N_18093,N_18928);
or UO_285 (O_285,N_18971,N_19526);
nand UO_286 (O_286,N_18981,N_18588);
and UO_287 (O_287,N_18838,N_19365);
or UO_288 (O_288,N_18879,N_18340);
xor UO_289 (O_289,N_19061,N_19598);
nor UO_290 (O_290,N_18372,N_18139);
xnor UO_291 (O_291,N_19016,N_19088);
nor UO_292 (O_292,N_19210,N_18104);
or UO_293 (O_293,N_18141,N_18915);
or UO_294 (O_294,N_19400,N_19394);
nor UO_295 (O_295,N_18793,N_19341);
xor UO_296 (O_296,N_19143,N_18862);
xor UO_297 (O_297,N_19099,N_19232);
nor UO_298 (O_298,N_18511,N_18945);
nand UO_299 (O_299,N_19634,N_18272);
and UO_300 (O_300,N_19403,N_18904);
nor UO_301 (O_301,N_18508,N_19665);
xnor UO_302 (O_302,N_18096,N_19790);
nor UO_303 (O_303,N_19378,N_19182);
xor UO_304 (O_304,N_18130,N_19897);
and UO_305 (O_305,N_19495,N_18468);
nor UO_306 (O_306,N_18998,N_19462);
and UO_307 (O_307,N_18298,N_19362);
or UO_308 (O_308,N_18696,N_19170);
nand UO_309 (O_309,N_19614,N_18539);
or UO_310 (O_310,N_18390,N_19908);
and UO_311 (O_311,N_18609,N_19509);
or UO_312 (O_312,N_19447,N_18781);
and UO_313 (O_313,N_18418,N_19957);
nand UO_314 (O_314,N_19159,N_18598);
and UO_315 (O_315,N_19417,N_18025);
nor UO_316 (O_316,N_18363,N_19864);
nor UO_317 (O_317,N_19281,N_19854);
nor UO_318 (O_318,N_18882,N_19105);
nand UO_319 (O_319,N_19759,N_18822);
and UO_320 (O_320,N_19706,N_19192);
xor UO_321 (O_321,N_18819,N_19235);
and UO_322 (O_322,N_19618,N_19966);
and UO_323 (O_323,N_19616,N_18279);
and UO_324 (O_324,N_18435,N_19709);
or UO_325 (O_325,N_18055,N_19605);
xor UO_326 (O_326,N_19558,N_18514);
xor UO_327 (O_327,N_19189,N_18821);
nor UO_328 (O_328,N_19707,N_18080);
nor UO_329 (O_329,N_19810,N_18223);
and UO_330 (O_330,N_19454,N_18501);
xnor UO_331 (O_331,N_19620,N_19151);
nor UO_332 (O_332,N_19954,N_19436);
nor UO_333 (O_333,N_18164,N_19772);
nand UO_334 (O_334,N_19819,N_18254);
nand UO_335 (O_335,N_19662,N_19632);
xor UO_336 (O_336,N_18847,N_18795);
nor UO_337 (O_337,N_19164,N_18996);
and UO_338 (O_338,N_19733,N_19003);
or UO_339 (O_339,N_19973,N_19216);
nand UO_340 (O_340,N_19218,N_18608);
or UO_341 (O_341,N_19683,N_19035);
nor UO_342 (O_342,N_18295,N_19408);
nand UO_343 (O_343,N_19181,N_18667);
xor UO_344 (O_344,N_18623,N_19108);
nand UO_345 (O_345,N_18967,N_18983);
and UO_346 (O_346,N_19044,N_18103);
nor UO_347 (O_347,N_18274,N_19568);
xnor UO_348 (O_348,N_19402,N_18182);
xnor UO_349 (O_349,N_19611,N_19079);
and UO_350 (O_350,N_18601,N_19370);
nor UO_351 (O_351,N_19659,N_19515);
xor UO_352 (O_352,N_18963,N_19226);
xor UO_353 (O_353,N_18651,N_18233);
and UO_354 (O_354,N_19677,N_19202);
nor UO_355 (O_355,N_19155,N_18617);
nand UO_356 (O_356,N_19795,N_19658);
xor UO_357 (O_357,N_18587,N_18269);
nor UO_358 (O_358,N_18763,N_18825);
nand UO_359 (O_359,N_18635,N_18186);
nor UO_360 (O_360,N_19684,N_18691);
nand UO_361 (O_361,N_19030,N_18373);
or UO_362 (O_362,N_18914,N_19421);
and UO_363 (O_363,N_18689,N_18889);
xor UO_364 (O_364,N_18836,N_19321);
and UO_365 (O_365,N_19979,N_18334);
nand UO_366 (O_366,N_18950,N_19579);
xor UO_367 (O_367,N_18948,N_18302);
and UO_368 (O_368,N_18465,N_18614);
or UO_369 (O_369,N_18870,N_18349);
nand UO_370 (O_370,N_19528,N_18369);
nand UO_371 (O_371,N_19160,N_18520);
or UO_372 (O_372,N_18749,N_19329);
nand UO_373 (O_373,N_19177,N_18644);
or UO_374 (O_374,N_19695,N_19555);
xnor UO_375 (O_375,N_19409,N_19717);
and UO_376 (O_376,N_18935,N_18878);
nand UO_377 (O_377,N_18944,N_18569);
and UO_378 (O_378,N_18367,N_18778);
or UO_379 (O_379,N_18234,N_18896);
nor UO_380 (O_380,N_19991,N_18687);
nand UO_381 (O_381,N_18297,N_18247);
and UO_382 (O_382,N_18656,N_18355);
nand UO_383 (O_383,N_18512,N_18423);
xnor UO_384 (O_384,N_18605,N_19587);
or UO_385 (O_385,N_19943,N_19425);
or UO_386 (O_386,N_19907,N_18918);
nor UO_387 (O_387,N_18683,N_19782);
nand UO_388 (O_388,N_19977,N_19919);
nor UO_389 (O_389,N_19763,N_18908);
or UO_390 (O_390,N_18757,N_18665);
nand UO_391 (O_391,N_18420,N_19465);
nand UO_392 (O_392,N_18865,N_19443);
or UO_393 (O_393,N_19320,N_18602);
nor UO_394 (O_394,N_18946,N_18054);
or UO_395 (O_395,N_19187,N_18442);
xor UO_396 (O_396,N_18634,N_19883);
and UO_397 (O_397,N_19201,N_18018);
nand UO_398 (O_398,N_19788,N_18310);
nor UO_399 (O_399,N_19012,N_18591);
and UO_400 (O_400,N_19173,N_19873);
nand UO_401 (O_401,N_18729,N_18679);
xnor UO_402 (O_402,N_18716,N_18281);
nor UO_403 (O_403,N_19719,N_19093);
xor UO_404 (O_404,N_19938,N_18811);
and UO_405 (O_405,N_18086,N_19773);
and UO_406 (O_406,N_18888,N_18738);
or UO_407 (O_407,N_18190,N_18413);
nand UO_408 (O_408,N_18009,N_18561);
nand UO_409 (O_409,N_19544,N_19716);
nor UO_410 (O_410,N_18353,N_19457);
nor UO_411 (O_411,N_19851,N_19446);
or UO_412 (O_412,N_18003,N_18395);
nand UO_413 (O_413,N_18858,N_19308);
xnor UO_414 (O_414,N_19724,N_18966);
nor UO_415 (O_415,N_18472,N_19204);
and UO_416 (O_416,N_19055,N_18396);
nand UO_417 (O_417,N_19136,N_19829);
and UO_418 (O_418,N_19175,N_18929);
nor UO_419 (O_419,N_18962,N_18239);
and UO_420 (O_420,N_19257,N_19019);
and UO_421 (O_421,N_18028,N_18912);
and UO_422 (O_422,N_18463,N_18077);
nand UO_423 (O_423,N_19312,N_19319);
nor UO_424 (O_424,N_19190,N_19249);
xnor UO_425 (O_425,N_18322,N_19351);
nand UO_426 (O_426,N_19650,N_19642);
or UO_427 (O_427,N_19224,N_18282);
xor UO_428 (O_428,N_19702,N_19137);
and UO_429 (O_429,N_19288,N_19978);
and UO_430 (O_430,N_18982,N_18155);
or UO_431 (O_431,N_18227,N_18380);
and UO_432 (O_432,N_19636,N_18577);
or UO_433 (O_433,N_18167,N_18877);
nor UO_434 (O_434,N_18633,N_19842);
xor UO_435 (O_435,N_19033,N_19350);
xor UO_436 (O_436,N_18660,N_18685);
and UO_437 (O_437,N_19344,N_18118);
xnor UO_438 (O_438,N_19444,N_19227);
nor UO_439 (O_439,N_18050,N_19287);
nand UO_440 (O_440,N_18798,N_19612);
nor UO_441 (O_441,N_19014,N_18523);
nand UO_442 (O_442,N_19456,N_18012);
nand UO_443 (O_443,N_19686,N_19793);
xor UO_444 (O_444,N_19393,N_18787);
or UO_445 (O_445,N_19223,N_18046);
xor UO_446 (O_446,N_19212,N_19451);
nand UO_447 (O_447,N_19936,N_18592);
and UO_448 (O_448,N_18484,N_18329);
and UO_449 (O_449,N_19640,N_19849);
and UO_450 (O_450,N_18366,N_19087);
xor UO_451 (O_451,N_18952,N_18377);
nand UO_452 (O_452,N_18085,N_19046);
and UO_453 (O_453,N_19723,N_18969);
nand UO_454 (O_454,N_18476,N_18416);
xor UO_455 (O_455,N_19865,N_18597);
nand UO_456 (O_456,N_18808,N_19505);
xor UO_457 (O_457,N_19391,N_19206);
xor UO_458 (O_458,N_19844,N_19673);
xor UO_459 (O_459,N_19550,N_18433);
and UO_460 (O_460,N_18613,N_19990);
and UO_461 (O_461,N_19918,N_19399);
nor UO_462 (O_462,N_19917,N_19771);
xnor UO_463 (O_463,N_18562,N_19126);
nand UO_464 (O_464,N_18051,N_19420);
nor UO_465 (O_465,N_18036,N_19435);
xor UO_466 (O_466,N_19647,N_19975);
or UO_467 (O_467,N_19735,N_18861);
and UO_468 (O_468,N_18545,N_18619);
or UO_469 (O_469,N_19423,N_18755);
nand UO_470 (O_470,N_18344,N_18611);
xor UO_471 (O_471,N_18319,N_19427);
or UO_472 (O_472,N_19300,N_18828);
nand UO_473 (O_473,N_19831,N_18612);
xor UO_474 (O_474,N_18820,N_18152);
xnor UO_475 (O_475,N_19910,N_19469);
and UO_476 (O_476,N_19856,N_18791);
and UO_477 (O_477,N_18579,N_19488);
or UO_478 (O_478,N_19915,N_18110);
or UO_479 (O_479,N_18776,N_19057);
nand UO_480 (O_480,N_19923,N_19135);
xor UO_481 (O_481,N_18263,N_19693);
and UO_482 (O_482,N_19549,N_19497);
nand UO_483 (O_483,N_18098,N_18771);
nand UO_484 (O_484,N_19951,N_19243);
xnor UO_485 (O_485,N_19455,N_19326);
nor UO_486 (O_486,N_18438,N_19687);
xnor UO_487 (O_487,N_18629,N_18259);
or UO_488 (O_488,N_19685,N_18125);
nor UO_489 (O_489,N_19360,N_19896);
nor UO_490 (O_490,N_18774,N_18678);
nor UO_491 (O_491,N_18149,N_18483);
and UO_492 (O_492,N_18456,N_18551);
or UO_493 (O_493,N_19573,N_19710);
and UO_494 (O_494,N_18519,N_19833);
and UO_495 (O_495,N_18337,N_19615);
nor UO_496 (O_496,N_19882,N_19822);
nor UO_497 (O_497,N_19627,N_18244);
nor UO_498 (O_498,N_18394,N_18102);
xnor UO_499 (O_499,N_19386,N_18622);
and UO_500 (O_500,N_19817,N_19452);
nor UO_501 (O_501,N_19606,N_19379);
nor UO_502 (O_502,N_18552,N_19349);
or UO_503 (O_503,N_19338,N_19646);
nor UO_504 (O_504,N_19247,N_18217);
nand UO_505 (O_505,N_18071,N_19930);
xor UO_506 (O_506,N_18943,N_18412);
nor UO_507 (O_507,N_19194,N_19920);
and UO_508 (O_508,N_19404,N_18895);
and UO_509 (O_509,N_18256,N_19401);
nand UO_510 (O_510,N_19145,N_18557);
nand UO_511 (O_511,N_18474,N_18011);
nor UO_512 (O_512,N_18280,N_19828);
nand UO_513 (O_513,N_19275,N_18065);
and UO_514 (O_514,N_18932,N_19768);
or UO_515 (O_515,N_18288,N_18823);
and UO_516 (O_516,N_19696,N_18327);
or UO_517 (O_517,N_18422,N_19501);
xor UO_518 (O_518,N_18812,N_18427);
nor UO_519 (O_519,N_19237,N_19661);
nor UO_520 (O_520,N_18524,N_18550);
nand UO_521 (O_521,N_19902,N_18284);
or UO_522 (O_522,N_18509,N_19547);
xor UO_523 (O_523,N_18548,N_19688);
nand UO_524 (O_524,N_18040,N_18976);
nor UO_525 (O_525,N_18978,N_19359);
nand UO_526 (O_526,N_19565,N_18830);
and UO_527 (O_527,N_18013,N_19663);
and UO_528 (O_528,N_19211,N_18753);
xnor UO_529 (O_529,N_19124,N_18770);
and UO_530 (O_530,N_19027,N_18461);
nor UO_531 (O_531,N_18328,N_18079);
nor UO_532 (O_532,N_19414,N_19600);
nor UO_533 (O_533,N_18590,N_18452);
nor UO_534 (O_534,N_18677,N_19989);
nand UO_535 (O_535,N_18299,N_18255);
nor UO_536 (O_536,N_18126,N_19584);
xnor UO_537 (O_537,N_18490,N_18454);
xor UO_538 (O_538,N_18653,N_18860);
xnor UO_539 (O_539,N_19333,N_19239);
and UO_540 (O_540,N_19068,N_18455);
or UO_541 (O_541,N_19080,N_18187);
nor UO_542 (O_542,N_19905,N_18338);
nor UO_543 (O_543,N_19241,N_19705);
or UO_544 (O_544,N_19361,N_18356);
nor UO_545 (O_545,N_19459,N_19208);
xor UO_546 (O_546,N_18495,N_18859);
nand UO_547 (O_547,N_18886,N_19075);
nor UO_548 (O_548,N_18097,N_19944);
nor UO_549 (O_549,N_19674,N_18221);
or UO_550 (O_550,N_18541,N_19556);
and UO_551 (O_551,N_19485,N_18201);
and UO_552 (O_552,N_18222,N_19523);
or UO_553 (O_553,N_18906,N_18990);
nor UO_554 (O_554,N_18321,N_18639);
xor UO_555 (O_555,N_18453,N_18318);
nand UO_556 (O_556,N_19496,N_18761);
or UO_557 (O_557,N_18956,N_19639);
or UO_558 (O_558,N_19522,N_19963);
or UO_559 (O_559,N_19117,N_19163);
nand UO_560 (O_560,N_19492,N_18641);
or UO_561 (O_561,N_18489,N_18585);
nand UO_562 (O_562,N_18019,N_19274);
nand UO_563 (O_563,N_19524,N_19049);
nor UO_564 (O_564,N_18088,N_18001);
xor UO_565 (O_565,N_18961,N_18199);
nor UO_566 (O_566,N_18262,N_18148);
nor UO_567 (O_567,N_19273,N_19730);
or UO_568 (O_568,N_18158,N_19777);
nand UO_569 (O_569,N_19655,N_19352);
nor UO_570 (O_570,N_19767,N_18804);
nor UO_571 (O_571,N_19645,N_18392);
and UO_572 (O_572,N_19948,N_19371);
and UO_573 (O_573,N_18410,N_18724);
or UO_574 (O_574,N_18894,N_19530);
or UO_575 (O_575,N_19884,N_18599);
nor UO_576 (O_576,N_18082,N_18032);
nor UO_577 (O_577,N_19595,N_18732);
nor UO_578 (O_578,N_18767,N_18491);
xor UO_579 (O_579,N_19946,N_18443);
nand UO_580 (O_580,N_18624,N_19668);
nor UO_581 (O_581,N_18625,N_18276);
nor UO_582 (O_582,N_19070,N_19157);
nand UO_583 (O_583,N_18672,N_18515);
nor UO_584 (O_584,N_18121,N_19560);
or UO_585 (O_585,N_19574,N_19535);
xor UO_586 (O_586,N_19388,N_18127);
or UO_587 (O_587,N_19567,N_19291);
or UO_588 (O_588,N_19279,N_19516);
and UO_589 (O_589,N_18901,N_19377);
and UO_590 (O_590,N_19304,N_18705);
or UO_591 (O_591,N_18136,N_19013);
xor UO_592 (O_592,N_19736,N_18038);
or UO_593 (O_593,N_19473,N_19356);
nand UO_594 (O_594,N_18553,N_19755);
nand UO_595 (O_595,N_19821,N_18106);
nor UO_596 (O_596,N_19860,N_18401);
and UO_597 (O_597,N_19154,N_19178);
nand UO_598 (O_598,N_18734,N_19738);
and UO_599 (O_599,N_19024,N_19985);
nand UO_600 (O_600,N_19357,N_18143);
nor UO_601 (O_601,N_18604,N_18138);
xor UO_602 (O_602,N_18723,N_19652);
xnor UO_603 (O_603,N_18195,N_18872);
xor UO_604 (O_604,N_18739,N_19440);
nor UO_605 (O_605,N_19214,N_18668);
xnor UO_606 (O_606,N_19900,N_19416);
or UO_607 (O_607,N_19871,N_18047);
or UO_608 (O_608,N_19701,N_19751);
or UO_609 (O_609,N_19729,N_19260);
nand UO_610 (O_610,N_18099,N_19781);
nand UO_611 (O_611,N_18090,N_18351);
xor UO_612 (O_612,N_18529,N_18855);
nand UO_613 (O_613,N_19219,N_19537);
nand UO_614 (O_614,N_19601,N_18659);
nand UO_615 (O_615,N_18285,N_19536);
and UO_616 (O_616,N_19450,N_18308);
nand UO_617 (O_617,N_18777,N_19298);
nor UO_618 (O_618,N_19432,N_19786);
and UO_619 (O_619,N_19770,N_19324);
and UO_620 (O_620,N_18754,N_19878);
xnor UO_621 (O_621,N_19775,N_18415);
xor UO_622 (O_622,N_18386,N_19760);
nor UO_623 (O_623,N_18801,N_19802);
or UO_624 (O_624,N_19467,N_18627);
xnor UO_625 (O_625,N_18730,N_19542);
or UO_626 (O_626,N_18022,N_18188);
or UO_627 (O_627,N_18873,N_18300);
or UO_628 (O_628,N_19780,N_18631);
xor UO_629 (O_629,N_18393,N_18839);
xor UO_630 (O_630,N_18984,N_18715);
or UO_631 (O_631,N_19069,N_19715);
nand UO_632 (O_632,N_18035,N_18140);
xnor UO_633 (O_633,N_19742,N_19270);
nand UO_634 (O_634,N_18959,N_19887);
xnor UO_635 (O_635,N_18014,N_18464);
and UO_636 (O_636,N_19179,N_18101);
nor UO_637 (O_637,N_18408,N_19272);
nand UO_638 (O_638,N_18907,N_18246);
nor UO_639 (O_639,N_19909,N_18439);
xor UO_640 (O_640,N_19589,N_19065);
nand UO_641 (O_641,N_19445,N_19675);
nand UO_642 (O_642,N_18039,N_18790);
and UO_643 (O_643,N_18431,N_19988);
and UO_644 (O_644,N_19323,N_19376);
nand UO_645 (O_645,N_19745,N_19422);
nor UO_646 (O_646,N_19835,N_19168);
and UO_647 (O_647,N_18926,N_19572);
or UO_648 (O_648,N_19866,N_19625);
and UO_649 (O_649,N_18949,N_18469);
nor UO_650 (O_650,N_19744,N_19090);
and UO_651 (O_651,N_18675,N_18350);
nor UO_652 (O_652,N_18287,N_19142);
nor UO_653 (O_653,N_18883,N_18002);
and UO_654 (O_654,N_18645,N_18448);
nor UO_655 (O_655,N_19949,N_18021);
nand UO_656 (O_656,N_19512,N_18502);
nand UO_657 (O_657,N_19570,N_19891);
nor UO_658 (O_658,N_18759,N_18174);
nor UO_659 (O_659,N_18686,N_18974);
xor UO_660 (O_660,N_18566,N_19327);
nor UO_661 (O_661,N_18434,N_19161);
nand UO_662 (O_662,N_19062,N_18972);
or UO_663 (O_663,N_19023,N_19820);
or UO_664 (O_664,N_18440,N_19603);
or UO_665 (O_665,N_19305,N_19511);
nand UO_666 (O_666,N_18784,N_19576);
xor UO_667 (O_667,N_19503,N_19041);
nand UO_668 (O_668,N_18348,N_18709);
or UO_669 (O_669,N_18892,N_19863);
and UO_670 (O_670,N_19754,N_19244);
or UO_671 (O_671,N_19937,N_19958);
nor UO_672 (O_672,N_18510,N_19624);
or UO_673 (O_673,N_18783,N_18023);
xor UO_674 (O_674,N_19407,N_18999);
and UO_675 (O_675,N_19976,N_18688);
or UO_676 (O_676,N_18582,N_19599);
xnor UO_677 (O_677,N_18384,N_19200);
nor UO_678 (O_678,N_18417,N_18837);
nand UO_679 (O_679,N_19731,N_18682);
nor UO_680 (O_680,N_19106,N_18070);
or UO_681 (O_681,N_18939,N_19020);
nor UO_682 (O_682,N_18089,N_19803);
xnor UO_683 (O_683,N_19113,N_19847);
or UO_684 (O_684,N_18069,N_19225);
nor UO_685 (O_685,N_19040,N_18060);
xnor UO_686 (O_686,N_19778,N_19582);
and UO_687 (O_687,N_18728,N_18075);
nor UO_688 (O_688,N_18371,N_18153);
and UO_689 (O_689,N_19588,N_18780);
nand UO_690 (O_690,N_18744,N_18424);
and UO_691 (O_691,N_18242,N_18834);
nand UO_692 (O_692,N_18171,N_19585);
or UO_693 (O_693,N_18846,N_19354);
and UO_694 (O_694,N_18437,N_18194);
or UO_695 (O_695,N_18742,N_19466);
or UO_696 (O_696,N_19566,N_19718);
and UO_697 (O_697,N_19797,N_19411);
nor UO_698 (O_698,N_18937,N_18193);
xnor UO_699 (O_699,N_18505,N_18913);
nor UO_700 (O_700,N_18095,N_19266);
or UO_701 (O_701,N_19531,N_18026);
nand UO_702 (O_702,N_18204,N_18556);
or UO_703 (O_703,N_19301,N_18210);
or UO_704 (O_704,N_18706,N_18175);
xnor UO_705 (O_705,N_19912,N_18414);
or UO_706 (O_706,N_19474,N_18250);
nor UO_707 (O_707,N_19931,N_18810);
xnor UO_708 (O_708,N_18973,N_18252);
xor UO_709 (O_709,N_19100,N_19796);
nor UO_710 (O_710,N_18400,N_18720);
or UO_711 (O_711,N_19054,N_19593);
nand UO_712 (O_712,N_18516,N_19111);
xnor UO_713 (O_713,N_18303,N_18004);
xnor UO_714 (O_714,N_19809,N_18721);
and UO_715 (O_715,N_19648,N_19434);
nand UO_716 (O_716,N_19894,N_19479);
nand UO_717 (O_717,N_19258,N_18200);
nand UO_718 (O_718,N_19318,N_19131);
nor UO_719 (O_719,N_19671,N_19699);
xor UO_720 (O_720,N_19424,N_18374);
xnor UO_721 (O_721,N_18058,N_19630);
nand UO_722 (O_722,N_19950,N_19203);
or UO_723 (O_723,N_19480,N_19929);
nand UO_724 (O_724,N_19690,N_19859);
nor UO_725 (O_725,N_18441,N_19058);
xnor UO_726 (O_726,N_19857,N_18887);
nand UO_727 (O_727,N_19322,N_19297);
xnor UO_728 (O_728,N_19410,N_18885);
nor UO_729 (O_729,N_19637,N_19193);
or UO_730 (O_730,N_19441,N_18646);
xor UO_731 (O_731,N_19029,N_18450);
nor UO_732 (O_732,N_19779,N_19123);
and UO_733 (O_733,N_18388,N_19335);
or UO_734 (O_734,N_19999,N_19245);
nor UO_735 (O_735,N_19562,N_19428);
nand UO_736 (O_736,N_18301,N_19419);
nand UO_737 (O_737,N_18652,N_19928);
xnor UO_738 (O_738,N_18710,N_18919);
or UO_739 (O_739,N_18726,N_19092);
xor UO_740 (O_740,N_19199,N_18532);
xor UO_741 (O_741,N_19808,N_18745);
nand UO_742 (O_742,N_19981,N_18241);
nor UO_743 (O_743,N_18033,N_18544);
or UO_744 (O_744,N_18640,N_18053);
xnor UO_745 (O_745,N_19332,N_18479);
or UO_746 (O_746,N_18596,N_18339);
nand UO_747 (O_747,N_18733,N_19721);
xnor UO_748 (O_748,N_18995,N_19118);
xor UO_749 (O_749,N_19899,N_18100);
xnor UO_750 (O_750,N_19302,N_18196);
xor UO_751 (O_751,N_18997,N_19694);
and UO_752 (O_752,N_18361,N_18800);
nand UO_753 (O_753,N_18078,N_19039);
nor UO_754 (O_754,N_19953,N_18564);
or UO_755 (O_755,N_19114,N_19703);
or UO_756 (O_756,N_19927,N_18900);
or UO_757 (O_757,N_18359,N_19765);
nand UO_758 (O_758,N_19283,N_19107);
nor UO_759 (O_759,N_19078,N_18113);
or UO_760 (O_760,N_18766,N_18020);
nor UO_761 (O_761,N_18954,N_18027);
nand UO_762 (O_762,N_19008,N_18876);
nor UO_763 (O_763,N_18063,N_19922);
nor UO_764 (O_764,N_18385,N_18421);
and UO_765 (O_765,N_19649,N_18657);
or UO_766 (O_766,N_19433,N_18845);
nor UO_767 (O_767,N_19236,N_18568);
and UO_768 (O_768,N_19487,N_18558);
and UO_769 (O_769,N_19478,N_19295);
and UO_770 (O_770,N_18695,N_19548);
xor UO_771 (O_771,N_18711,N_18107);
nor UO_772 (O_772,N_19221,N_18748);
nor UO_773 (O_773,N_18399,N_19010);
or UO_774 (O_774,N_19934,N_19148);
or UO_775 (O_775,N_19185,N_18988);
or UO_776 (O_776,N_18237,N_19885);
or UO_777 (O_777,N_19006,N_18428);
nand UO_778 (O_778,N_19756,N_19506);
and UO_779 (O_779,N_19774,N_19233);
nand UO_780 (O_780,N_19521,N_18628);
nor UO_781 (O_781,N_19368,N_18197);
nand UO_782 (O_782,N_19592,N_19165);
nor UO_783 (O_783,N_19026,N_19783);
nand UO_784 (O_784,N_19015,N_18874);
nor UO_785 (O_785,N_19841,N_18411);
xor UO_786 (O_786,N_19545,N_19551);
nor UO_787 (O_787,N_18378,N_19166);
nor UO_788 (O_788,N_19252,N_18513);
xor UO_789 (O_789,N_18061,N_18725);
and UO_790 (O_790,N_19510,N_19874);
xnor UO_791 (O_791,N_18570,N_19230);
xor UO_792 (O_792,N_18015,N_19418);
xnor UO_793 (O_793,N_19343,N_19557);
or UO_794 (O_794,N_18699,N_18224);
nor UO_795 (O_795,N_19127,N_18397);
nor UO_796 (O_796,N_19430,N_18409);
nand UO_797 (O_797,N_18309,N_19747);
or UO_798 (O_798,N_19766,N_19970);
nand UO_799 (O_799,N_18565,N_18987);
or UO_800 (O_800,N_18572,N_18648);
nand UO_801 (O_801,N_18330,N_18253);
nor UO_802 (O_802,N_19149,N_18647);
and UO_803 (O_803,N_18507,N_18486);
or UO_804 (O_804,N_19217,N_18666);
nand UO_805 (O_805,N_19031,N_19935);
xnor UO_806 (O_806,N_18663,N_18325);
and UO_807 (O_807,N_19306,N_19314);
and UO_808 (O_808,N_19813,N_19964);
or UO_809 (O_809,N_19848,N_18643);
nand UO_810 (O_810,N_18936,N_19053);
or UO_811 (O_811,N_18567,N_19138);
nor UO_812 (O_812,N_18903,N_19959);
nor UO_813 (O_813,N_18692,N_18775);
nand UO_814 (O_814,N_19942,N_18673);
xnor UO_815 (O_815,N_19825,N_19993);
nand UO_816 (O_816,N_18000,N_18170);
nor UO_817 (O_817,N_19468,N_18528);
nor UO_818 (O_818,N_18142,N_19961);
xnor UO_819 (O_819,N_19094,N_19152);
nand UO_820 (O_820,N_18881,N_18240);
xor UO_821 (O_821,N_19903,N_18133);
and UO_822 (O_822,N_18854,N_19613);
xor UO_823 (O_823,N_18251,N_18131);
and UO_824 (O_824,N_19836,N_19263);
nor UO_825 (O_825,N_19890,N_18059);
nand UO_826 (O_826,N_19102,N_18772);
nand UO_827 (O_827,N_19047,N_19538);
or UO_828 (O_828,N_19309,N_19340);
nor UO_829 (O_829,N_19983,N_18231);
or UO_830 (O_830,N_18578,N_19681);
nor UO_831 (O_831,N_18108,N_19277);
and UO_832 (O_832,N_19746,N_19207);
and UO_833 (O_833,N_18933,N_18518);
and UO_834 (O_834,N_18091,N_18481);
or UO_835 (O_835,N_18560,N_18220);
and UO_836 (O_836,N_19043,N_18184);
nor UO_837 (O_837,N_18760,N_19827);
and UO_838 (O_838,N_18581,N_19906);
or UO_839 (O_839,N_19853,N_18583);
nor UO_840 (O_840,N_19389,N_19296);
or UO_841 (O_841,N_18116,N_19880);
xor UO_842 (O_842,N_19980,N_18258);
xor UO_843 (O_843,N_19337,N_19405);
or UO_844 (O_844,N_18016,N_19748);
xnor UO_845 (O_845,N_18346,N_18813);
or UO_846 (O_846,N_19753,N_19784);
and UO_847 (O_847,N_18275,N_19564);
xnor UO_848 (O_848,N_19858,N_18637);
and UO_849 (O_849,N_18727,N_18621);
nand UO_850 (O_850,N_19741,N_19815);
nor UO_851 (O_851,N_18492,N_18563);
or UO_852 (O_852,N_19617,N_18909);
nand UO_853 (O_853,N_19034,N_18504);
and UO_854 (O_854,N_18891,N_19180);
nand UO_855 (O_855,N_19921,N_18740);
nand UO_856 (O_856,N_18307,N_19083);
nor UO_857 (O_857,N_18216,N_18818);
nor UO_858 (O_858,N_19834,N_18704);
xnor UO_859 (O_859,N_18209,N_19559);
and UO_860 (O_860,N_18407,N_19794);
and UO_861 (O_861,N_18485,N_18769);
nor UO_862 (O_862,N_19785,N_19940);
nand UO_863 (O_863,N_19525,N_18717);
and UO_864 (O_864,N_18712,N_19855);
nand UO_865 (O_865,N_18764,N_19119);
xnor UO_866 (O_866,N_19590,N_19626);
xor UO_867 (O_867,N_18992,N_19776);
nand UO_868 (O_868,N_18832,N_18986);
nand UO_869 (O_869,N_19475,N_19174);
or UO_870 (O_870,N_19752,N_18842);
nand UO_871 (O_871,N_18654,N_19670);
nor UO_872 (O_872,N_19643,N_19413);
or UO_873 (O_873,N_19577,N_18979);
xnor UO_874 (O_874,N_19261,N_18615);
nor UO_875 (O_875,N_19692,N_18341);
xor UO_876 (O_876,N_18230,N_18446);
nand UO_877 (O_877,N_19804,N_19364);
xnor UO_878 (O_878,N_19926,N_19628);
nor UO_879 (O_879,N_19651,N_18924);
nor UO_880 (O_880,N_19342,N_18066);
nand UO_881 (O_881,N_18714,N_18005);
and UO_882 (O_882,N_18185,N_19638);
xor UO_883 (O_883,N_19597,N_18863);
nor UO_884 (O_884,N_18041,N_18470);
nand UO_885 (O_885,N_19115,N_18487);
and UO_886 (O_886,N_19373,N_19387);
and UO_887 (O_887,N_18482,N_19032);
xnor UO_888 (O_888,N_18789,N_19050);
nand UO_889 (O_889,N_19011,N_18902);
and UO_890 (O_890,N_18343,N_18460);
or UO_891 (O_891,N_18831,N_19968);
xnor UO_892 (O_892,N_19893,N_18458);
or UO_893 (O_893,N_19476,N_19816);
xnor UO_894 (O_894,N_18311,N_18037);
or UO_895 (O_895,N_18700,N_19086);
nor UO_896 (O_896,N_19758,N_19870);
nor UO_897 (O_897,N_18814,N_18694);
nand UO_898 (O_898,N_18743,N_19382);
nor UO_899 (O_899,N_19073,N_18317);
nand UO_900 (O_900,N_19664,N_18736);
nor UO_901 (O_901,N_18352,N_18697);
xor UO_902 (O_902,N_18616,N_18955);
nor UO_903 (O_903,N_19251,N_18218);
or UO_904 (O_904,N_18938,N_18917);
and UO_905 (O_905,N_18034,N_19543);
nor UO_906 (O_906,N_19471,N_19071);
nand UO_907 (O_907,N_18266,N_18991);
nor UO_908 (O_908,N_18864,N_19392);
or UO_909 (O_909,N_18671,N_18062);
and UO_910 (O_910,N_19939,N_19348);
or UO_911 (O_911,N_18488,N_19737);
and UO_912 (O_912,N_19238,N_19952);
nor UO_913 (O_913,N_18044,N_18160);
nor UO_914 (O_914,N_18389,N_18135);
xor UO_915 (O_915,N_18698,N_18228);
and UO_916 (O_916,N_18315,N_18172);
and UO_917 (O_917,N_18805,N_18794);
or UO_918 (O_918,N_19353,N_18115);
nand UO_919 (O_919,N_18342,N_18527);
nor UO_920 (O_920,N_18741,N_19072);
and UO_921 (O_921,N_18642,N_19254);
and UO_922 (O_922,N_19038,N_19278);
and UO_923 (O_923,N_18181,N_19112);
nand UO_924 (O_924,N_18457,N_19007);
xnor UO_925 (O_925,N_19482,N_18916);
or UO_926 (O_926,N_19463,N_18547);
nor UO_927 (O_927,N_19483,N_18192);
nand UO_928 (O_928,N_19197,N_19169);
nand UO_929 (O_929,N_19845,N_19052);
and UO_930 (O_930,N_19791,N_18248);
nor UO_931 (O_931,N_18957,N_19888);
nor UO_932 (O_932,N_18941,N_19714);
nor UO_933 (O_933,N_18575,N_18942);
nand UO_934 (O_934,N_19215,N_18092);
and UO_935 (O_935,N_18144,N_19347);
xor UO_936 (O_936,N_19477,N_18360);
and UO_937 (O_937,N_19580,N_18203);
xnor UO_938 (O_938,N_18161,N_19689);
or UO_939 (O_939,N_18333,N_18229);
or UO_940 (O_940,N_18257,N_19631);
nand UO_941 (O_941,N_18163,N_19892);
xor UO_942 (O_942,N_18382,N_18816);
or UO_943 (O_943,N_19097,N_19904);
xnor UO_944 (O_944,N_19310,N_18674);
xor UO_945 (O_945,N_19259,N_19666);
and UO_946 (O_946,N_19947,N_18600);
and UO_947 (O_947,N_18191,N_19720);
or UO_948 (O_948,N_19830,N_18493);
xnor UO_949 (O_949,N_19962,N_18525);
or UO_950 (O_950,N_18782,N_18478);
or UO_951 (O_951,N_19125,N_19385);
nand UO_952 (O_952,N_19657,N_19231);
or UO_953 (O_953,N_18017,N_19914);
nand UO_954 (O_954,N_19622,N_18236);
nor UO_955 (O_955,N_18426,N_19654);
xnor UO_956 (O_956,N_18496,N_19481);
nor UO_957 (O_957,N_19213,N_19331);
or UO_958 (O_958,N_19095,N_19412);
nor UO_959 (O_959,N_19932,N_19426);
xor UO_960 (O_960,N_19541,N_19826);
xor UO_961 (O_961,N_18376,N_18922);
and UO_962 (O_962,N_18803,N_18354);
and UO_963 (O_963,N_18147,N_19732);
xnor UO_964 (O_964,N_19712,N_18773);
and UO_965 (O_965,N_19867,N_19691);
xnor UO_966 (O_966,N_18670,N_18826);
and UO_967 (O_967,N_19328,N_19299);
nor UO_968 (O_968,N_19586,N_19514);
and UO_969 (O_969,N_18536,N_18620);
nor UO_970 (O_970,N_19022,N_19397);
nand UO_971 (O_971,N_18159,N_18451);
xor UO_972 (O_972,N_19761,N_19438);
nor UO_973 (O_973,N_18594,N_18169);
and UO_974 (O_974,N_18261,N_18543);
or UO_975 (O_975,N_18362,N_18157);
nand UO_976 (O_976,N_18444,N_19183);
nand UO_977 (O_977,N_19563,N_19059);
and UO_978 (O_978,N_18336,N_18404);
nor UO_979 (O_979,N_18105,N_18162);
or UO_980 (O_980,N_19533,N_18994);
or UO_981 (O_981,N_19242,N_19680);
and UO_982 (O_982,N_19713,N_18707);
nand UO_983 (O_983,N_18145,N_19575);
or UO_984 (O_984,N_18271,N_19129);
xnor UO_985 (O_985,N_19502,N_19660);
xor UO_986 (O_986,N_19889,N_19596);
xor UO_987 (O_987,N_18921,N_18202);
and UO_988 (O_988,N_19004,N_19749);
nand UO_989 (O_989,N_18785,N_18844);
nor UO_990 (O_990,N_18031,N_18853);
and UO_991 (O_991,N_19448,N_19104);
nand UO_992 (O_992,N_18068,N_18595);
nand UO_993 (O_993,N_19063,N_19998);
or UO_994 (O_994,N_19096,N_19787);
or UO_995 (O_995,N_19876,N_18713);
or UO_996 (O_996,N_19604,N_19798);
or UO_997 (O_997,N_19167,N_18829);
and UO_998 (O_998,N_19682,N_19678);
nor UO_999 (O_999,N_18802,N_18296);
nor UO_1000 (O_1000,N_19131,N_19875);
nor UO_1001 (O_1001,N_19942,N_19241);
or UO_1002 (O_1002,N_19656,N_19214);
or UO_1003 (O_1003,N_19478,N_19026);
nor UO_1004 (O_1004,N_19862,N_18485);
nor UO_1005 (O_1005,N_18592,N_19580);
nand UO_1006 (O_1006,N_18668,N_19039);
or UO_1007 (O_1007,N_18754,N_19467);
xor UO_1008 (O_1008,N_19116,N_19104);
xor UO_1009 (O_1009,N_18464,N_19958);
nor UO_1010 (O_1010,N_18242,N_18177);
nand UO_1011 (O_1011,N_18615,N_18340);
and UO_1012 (O_1012,N_18895,N_19283);
and UO_1013 (O_1013,N_19332,N_18309);
or UO_1014 (O_1014,N_18197,N_19238);
nand UO_1015 (O_1015,N_19564,N_18620);
or UO_1016 (O_1016,N_18585,N_19857);
xnor UO_1017 (O_1017,N_18702,N_19569);
xor UO_1018 (O_1018,N_18413,N_18544);
nand UO_1019 (O_1019,N_18907,N_18696);
and UO_1020 (O_1020,N_19702,N_18468);
nand UO_1021 (O_1021,N_19734,N_18795);
nand UO_1022 (O_1022,N_18055,N_18080);
xor UO_1023 (O_1023,N_18969,N_19170);
nor UO_1024 (O_1024,N_18243,N_18762);
nor UO_1025 (O_1025,N_18723,N_19502);
or UO_1026 (O_1026,N_18609,N_18389);
xnor UO_1027 (O_1027,N_18259,N_18286);
xnor UO_1028 (O_1028,N_18547,N_19643);
or UO_1029 (O_1029,N_19427,N_18248);
or UO_1030 (O_1030,N_19637,N_18994);
xnor UO_1031 (O_1031,N_18011,N_18840);
and UO_1032 (O_1032,N_19295,N_18433);
xnor UO_1033 (O_1033,N_18967,N_19972);
nor UO_1034 (O_1034,N_19102,N_19492);
or UO_1035 (O_1035,N_18272,N_19813);
or UO_1036 (O_1036,N_18150,N_19220);
and UO_1037 (O_1037,N_19043,N_19596);
or UO_1038 (O_1038,N_19464,N_19522);
or UO_1039 (O_1039,N_19530,N_19640);
nor UO_1040 (O_1040,N_19749,N_18889);
nor UO_1041 (O_1041,N_18555,N_18487);
xor UO_1042 (O_1042,N_19346,N_19270);
xor UO_1043 (O_1043,N_19701,N_18852);
nand UO_1044 (O_1044,N_18951,N_18474);
xnor UO_1045 (O_1045,N_18944,N_19995);
and UO_1046 (O_1046,N_18265,N_19795);
xnor UO_1047 (O_1047,N_18436,N_19182);
xnor UO_1048 (O_1048,N_19678,N_19144);
nor UO_1049 (O_1049,N_18492,N_18345);
or UO_1050 (O_1050,N_19361,N_19055);
nand UO_1051 (O_1051,N_18858,N_18221);
nor UO_1052 (O_1052,N_19057,N_18480);
or UO_1053 (O_1053,N_18352,N_18369);
nand UO_1054 (O_1054,N_19158,N_19568);
xor UO_1055 (O_1055,N_18603,N_19580);
xor UO_1056 (O_1056,N_18006,N_19089);
and UO_1057 (O_1057,N_19712,N_18499);
and UO_1058 (O_1058,N_19908,N_18282);
xor UO_1059 (O_1059,N_19564,N_18630);
nand UO_1060 (O_1060,N_19517,N_18951);
nand UO_1061 (O_1061,N_19531,N_18612);
nand UO_1062 (O_1062,N_19786,N_18797);
xnor UO_1063 (O_1063,N_18222,N_19747);
or UO_1064 (O_1064,N_19247,N_19990);
and UO_1065 (O_1065,N_19735,N_19895);
nand UO_1066 (O_1066,N_18902,N_18219);
and UO_1067 (O_1067,N_19942,N_18446);
xnor UO_1068 (O_1068,N_19637,N_19735);
nand UO_1069 (O_1069,N_19271,N_19929);
nor UO_1070 (O_1070,N_19063,N_18110);
or UO_1071 (O_1071,N_18034,N_18164);
nand UO_1072 (O_1072,N_18778,N_19638);
xnor UO_1073 (O_1073,N_18560,N_19009);
nor UO_1074 (O_1074,N_19447,N_18604);
and UO_1075 (O_1075,N_18413,N_19549);
or UO_1076 (O_1076,N_19039,N_18489);
or UO_1077 (O_1077,N_19417,N_19505);
or UO_1078 (O_1078,N_18874,N_18077);
and UO_1079 (O_1079,N_18363,N_19484);
or UO_1080 (O_1080,N_19221,N_18262);
nand UO_1081 (O_1081,N_18553,N_18939);
xnor UO_1082 (O_1082,N_18960,N_19124);
xor UO_1083 (O_1083,N_18783,N_18198);
nor UO_1084 (O_1084,N_19524,N_18264);
nand UO_1085 (O_1085,N_19626,N_18187);
and UO_1086 (O_1086,N_18181,N_19170);
nand UO_1087 (O_1087,N_18480,N_19592);
or UO_1088 (O_1088,N_19654,N_18240);
or UO_1089 (O_1089,N_19514,N_18170);
xnor UO_1090 (O_1090,N_19935,N_19960);
xnor UO_1091 (O_1091,N_19595,N_19314);
or UO_1092 (O_1092,N_19433,N_19577);
nor UO_1093 (O_1093,N_19108,N_19485);
or UO_1094 (O_1094,N_19560,N_18921);
nor UO_1095 (O_1095,N_19293,N_18816);
xor UO_1096 (O_1096,N_19378,N_18821);
and UO_1097 (O_1097,N_19527,N_19554);
nor UO_1098 (O_1098,N_19793,N_18227);
nor UO_1099 (O_1099,N_18066,N_18624);
xnor UO_1100 (O_1100,N_19024,N_18669);
or UO_1101 (O_1101,N_18697,N_18795);
xnor UO_1102 (O_1102,N_19383,N_18631);
or UO_1103 (O_1103,N_18520,N_18424);
nand UO_1104 (O_1104,N_19254,N_18483);
and UO_1105 (O_1105,N_19827,N_18571);
or UO_1106 (O_1106,N_19563,N_19324);
and UO_1107 (O_1107,N_19157,N_19487);
and UO_1108 (O_1108,N_18005,N_19838);
or UO_1109 (O_1109,N_19414,N_18445);
nor UO_1110 (O_1110,N_18204,N_18003);
and UO_1111 (O_1111,N_18373,N_19079);
and UO_1112 (O_1112,N_18281,N_19797);
xor UO_1113 (O_1113,N_19012,N_18452);
nor UO_1114 (O_1114,N_18773,N_18648);
and UO_1115 (O_1115,N_19218,N_19683);
nand UO_1116 (O_1116,N_18206,N_19757);
nor UO_1117 (O_1117,N_18231,N_18142);
or UO_1118 (O_1118,N_19836,N_18515);
or UO_1119 (O_1119,N_18217,N_19970);
xnor UO_1120 (O_1120,N_19067,N_19409);
or UO_1121 (O_1121,N_19692,N_18755);
nand UO_1122 (O_1122,N_19675,N_19490);
or UO_1123 (O_1123,N_18209,N_19835);
or UO_1124 (O_1124,N_18663,N_19512);
xnor UO_1125 (O_1125,N_19843,N_19090);
and UO_1126 (O_1126,N_19871,N_19911);
and UO_1127 (O_1127,N_18765,N_18414);
and UO_1128 (O_1128,N_18329,N_18545);
nor UO_1129 (O_1129,N_19980,N_18212);
nand UO_1130 (O_1130,N_19223,N_19544);
xnor UO_1131 (O_1131,N_19781,N_19410);
or UO_1132 (O_1132,N_18824,N_19089);
nand UO_1133 (O_1133,N_18690,N_19270);
or UO_1134 (O_1134,N_19830,N_18349);
nor UO_1135 (O_1135,N_19673,N_18183);
nor UO_1136 (O_1136,N_19196,N_18528);
or UO_1137 (O_1137,N_18302,N_19150);
nand UO_1138 (O_1138,N_19987,N_19624);
nand UO_1139 (O_1139,N_18078,N_19381);
xor UO_1140 (O_1140,N_18229,N_19159);
nand UO_1141 (O_1141,N_19558,N_18131);
and UO_1142 (O_1142,N_18274,N_19513);
nor UO_1143 (O_1143,N_18733,N_19556);
and UO_1144 (O_1144,N_18457,N_19385);
nor UO_1145 (O_1145,N_18843,N_18114);
xor UO_1146 (O_1146,N_18407,N_19150);
and UO_1147 (O_1147,N_18957,N_19374);
xor UO_1148 (O_1148,N_19870,N_18719);
nor UO_1149 (O_1149,N_19182,N_18590);
nor UO_1150 (O_1150,N_18720,N_19340);
or UO_1151 (O_1151,N_18047,N_18454);
and UO_1152 (O_1152,N_19809,N_18351);
nand UO_1153 (O_1153,N_18876,N_18724);
nand UO_1154 (O_1154,N_18683,N_18995);
xnor UO_1155 (O_1155,N_18600,N_19183);
xnor UO_1156 (O_1156,N_18560,N_18059);
xor UO_1157 (O_1157,N_19059,N_18756);
xor UO_1158 (O_1158,N_18808,N_18812);
nor UO_1159 (O_1159,N_19127,N_18764);
or UO_1160 (O_1160,N_18676,N_18364);
and UO_1161 (O_1161,N_19748,N_18100);
or UO_1162 (O_1162,N_18357,N_18194);
xnor UO_1163 (O_1163,N_18563,N_19876);
nor UO_1164 (O_1164,N_19844,N_18294);
xnor UO_1165 (O_1165,N_18676,N_18841);
and UO_1166 (O_1166,N_18861,N_18092);
and UO_1167 (O_1167,N_19813,N_18532);
and UO_1168 (O_1168,N_19086,N_19293);
or UO_1169 (O_1169,N_19173,N_19438);
and UO_1170 (O_1170,N_18950,N_18834);
nor UO_1171 (O_1171,N_18715,N_19337);
xnor UO_1172 (O_1172,N_19705,N_18884);
or UO_1173 (O_1173,N_19674,N_18367);
nor UO_1174 (O_1174,N_19059,N_19013);
or UO_1175 (O_1175,N_18109,N_19554);
or UO_1176 (O_1176,N_18441,N_18877);
xnor UO_1177 (O_1177,N_18557,N_18439);
xor UO_1178 (O_1178,N_19330,N_18211);
and UO_1179 (O_1179,N_18325,N_18706);
nor UO_1180 (O_1180,N_18817,N_19136);
nor UO_1181 (O_1181,N_19990,N_18870);
xnor UO_1182 (O_1182,N_18985,N_18555);
nand UO_1183 (O_1183,N_18526,N_18128);
or UO_1184 (O_1184,N_18464,N_18227);
or UO_1185 (O_1185,N_18314,N_19793);
nor UO_1186 (O_1186,N_18330,N_19738);
nand UO_1187 (O_1187,N_19619,N_18117);
or UO_1188 (O_1188,N_18861,N_18276);
or UO_1189 (O_1189,N_19937,N_19340);
and UO_1190 (O_1190,N_18032,N_19187);
nor UO_1191 (O_1191,N_19940,N_19598);
and UO_1192 (O_1192,N_19794,N_19369);
or UO_1193 (O_1193,N_18683,N_18275);
or UO_1194 (O_1194,N_19153,N_18485);
nand UO_1195 (O_1195,N_18127,N_19253);
and UO_1196 (O_1196,N_18310,N_19495);
xor UO_1197 (O_1197,N_19763,N_18460);
or UO_1198 (O_1198,N_19701,N_18302);
nor UO_1199 (O_1199,N_19239,N_19540);
and UO_1200 (O_1200,N_18524,N_18357);
nand UO_1201 (O_1201,N_18170,N_19154);
or UO_1202 (O_1202,N_19340,N_18394);
and UO_1203 (O_1203,N_18474,N_19336);
and UO_1204 (O_1204,N_18100,N_18848);
nand UO_1205 (O_1205,N_19913,N_19199);
and UO_1206 (O_1206,N_19305,N_19253);
xnor UO_1207 (O_1207,N_19705,N_18550);
nand UO_1208 (O_1208,N_19900,N_19301);
nor UO_1209 (O_1209,N_18417,N_19876);
nor UO_1210 (O_1210,N_18221,N_19057);
and UO_1211 (O_1211,N_19223,N_19521);
nand UO_1212 (O_1212,N_19759,N_18739);
nand UO_1213 (O_1213,N_18054,N_19463);
xnor UO_1214 (O_1214,N_19748,N_18510);
and UO_1215 (O_1215,N_18865,N_18876);
and UO_1216 (O_1216,N_18649,N_19784);
xor UO_1217 (O_1217,N_19901,N_19712);
xor UO_1218 (O_1218,N_18234,N_18575);
or UO_1219 (O_1219,N_18700,N_18418);
and UO_1220 (O_1220,N_18993,N_18955);
and UO_1221 (O_1221,N_19652,N_19767);
xor UO_1222 (O_1222,N_19510,N_18550);
xor UO_1223 (O_1223,N_19099,N_18149);
xnor UO_1224 (O_1224,N_18577,N_18553);
and UO_1225 (O_1225,N_18011,N_18647);
and UO_1226 (O_1226,N_19510,N_18121);
nor UO_1227 (O_1227,N_19466,N_18591);
nor UO_1228 (O_1228,N_19665,N_19625);
and UO_1229 (O_1229,N_19936,N_19604);
or UO_1230 (O_1230,N_19124,N_18562);
nor UO_1231 (O_1231,N_19629,N_19486);
or UO_1232 (O_1232,N_18200,N_19419);
and UO_1233 (O_1233,N_18873,N_19154);
xnor UO_1234 (O_1234,N_19010,N_18450);
and UO_1235 (O_1235,N_19651,N_18138);
or UO_1236 (O_1236,N_19105,N_19270);
nand UO_1237 (O_1237,N_18288,N_19543);
xnor UO_1238 (O_1238,N_18481,N_19836);
nor UO_1239 (O_1239,N_18219,N_19485);
nand UO_1240 (O_1240,N_18395,N_18580);
nor UO_1241 (O_1241,N_18219,N_18396);
or UO_1242 (O_1242,N_18771,N_18475);
xnor UO_1243 (O_1243,N_19610,N_19353);
or UO_1244 (O_1244,N_19976,N_18690);
xor UO_1245 (O_1245,N_19140,N_18255);
nand UO_1246 (O_1246,N_19998,N_18946);
and UO_1247 (O_1247,N_18002,N_18251);
and UO_1248 (O_1248,N_19157,N_19339);
or UO_1249 (O_1249,N_19168,N_19543);
nand UO_1250 (O_1250,N_18990,N_18438);
and UO_1251 (O_1251,N_19099,N_18127);
nand UO_1252 (O_1252,N_19190,N_19855);
nand UO_1253 (O_1253,N_19858,N_18503);
xor UO_1254 (O_1254,N_19441,N_19069);
and UO_1255 (O_1255,N_19609,N_19545);
and UO_1256 (O_1256,N_18969,N_18557);
nor UO_1257 (O_1257,N_19971,N_18354);
xnor UO_1258 (O_1258,N_19239,N_19058);
nor UO_1259 (O_1259,N_19932,N_19696);
nand UO_1260 (O_1260,N_19947,N_18857);
or UO_1261 (O_1261,N_18953,N_18828);
nand UO_1262 (O_1262,N_18468,N_18690);
xnor UO_1263 (O_1263,N_18621,N_18796);
nand UO_1264 (O_1264,N_18812,N_19171);
or UO_1265 (O_1265,N_19201,N_18941);
or UO_1266 (O_1266,N_18647,N_18213);
or UO_1267 (O_1267,N_19043,N_19041);
nand UO_1268 (O_1268,N_18426,N_18694);
nor UO_1269 (O_1269,N_18869,N_19111);
xor UO_1270 (O_1270,N_18604,N_19625);
xnor UO_1271 (O_1271,N_18680,N_18145);
nor UO_1272 (O_1272,N_19084,N_19892);
xnor UO_1273 (O_1273,N_19044,N_19581);
and UO_1274 (O_1274,N_19519,N_19265);
nand UO_1275 (O_1275,N_18247,N_18023);
nand UO_1276 (O_1276,N_18444,N_18835);
nand UO_1277 (O_1277,N_18141,N_18759);
and UO_1278 (O_1278,N_18492,N_18208);
nand UO_1279 (O_1279,N_18215,N_18831);
nor UO_1280 (O_1280,N_18209,N_18084);
xnor UO_1281 (O_1281,N_19159,N_18139);
and UO_1282 (O_1282,N_19679,N_18834);
nor UO_1283 (O_1283,N_18450,N_18375);
or UO_1284 (O_1284,N_18423,N_19217);
nor UO_1285 (O_1285,N_18892,N_18844);
and UO_1286 (O_1286,N_18589,N_18745);
nand UO_1287 (O_1287,N_19997,N_18868);
nand UO_1288 (O_1288,N_18453,N_18057);
and UO_1289 (O_1289,N_18030,N_19940);
or UO_1290 (O_1290,N_18473,N_19840);
or UO_1291 (O_1291,N_19895,N_19108);
and UO_1292 (O_1292,N_18022,N_18336);
nor UO_1293 (O_1293,N_18683,N_18661);
and UO_1294 (O_1294,N_19937,N_19542);
or UO_1295 (O_1295,N_18101,N_18154);
nand UO_1296 (O_1296,N_18256,N_19888);
nand UO_1297 (O_1297,N_19981,N_19301);
or UO_1298 (O_1298,N_18524,N_18680);
xnor UO_1299 (O_1299,N_18057,N_19168);
nor UO_1300 (O_1300,N_19264,N_18162);
xnor UO_1301 (O_1301,N_19909,N_19906);
xor UO_1302 (O_1302,N_18190,N_18788);
nand UO_1303 (O_1303,N_18557,N_18564);
nand UO_1304 (O_1304,N_19516,N_18429);
xnor UO_1305 (O_1305,N_19684,N_19928);
xor UO_1306 (O_1306,N_18786,N_19864);
nand UO_1307 (O_1307,N_18361,N_18082);
nor UO_1308 (O_1308,N_18750,N_18042);
nor UO_1309 (O_1309,N_18847,N_19786);
or UO_1310 (O_1310,N_19722,N_19405);
and UO_1311 (O_1311,N_18367,N_19847);
nand UO_1312 (O_1312,N_18209,N_18046);
or UO_1313 (O_1313,N_18567,N_19000);
or UO_1314 (O_1314,N_19767,N_18325);
or UO_1315 (O_1315,N_18083,N_19766);
xnor UO_1316 (O_1316,N_18752,N_19648);
or UO_1317 (O_1317,N_18064,N_18493);
xnor UO_1318 (O_1318,N_19398,N_19618);
nor UO_1319 (O_1319,N_18942,N_18247);
or UO_1320 (O_1320,N_19684,N_18548);
or UO_1321 (O_1321,N_18674,N_19421);
xnor UO_1322 (O_1322,N_18235,N_19883);
nor UO_1323 (O_1323,N_18629,N_18698);
and UO_1324 (O_1324,N_18809,N_19474);
nor UO_1325 (O_1325,N_18234,N_18073);
nor UO_1326 (O_1326,N_19953,N_18100);
or UO_1327 (O_1327,N_19786,N_18924);
xnor UO_1328 (O_1328,N_19137,N_19653);
and UO_1329 (O_1329,N_19037,N_18092);
and UO_1330 (O_1330,N_19891,N_19127);
and UO_1331 (O_1331,N_19467,N_18924);
nand UO_1332 (O_1332,N_19647,N_19216);
nand UO_1333 (O_1333,N_19780,N_19597);
or UO_1334 (O_1334,N_18532,N_18613);
and UO_1335 (O_1335,N_19176,N_18866);
and UO_1336 (O_1336,N_18889,N_18368);
nor UO_1337 (O_1337,N_18438,N_18276);
and UO_1338 (O_1338,N_19361,N_18487);
or UO_1339 (O_1339,N_19732,N_19863);
nor UO_1340 (O_1340,N_19047,N_19111);
xor UO_1341 (O_1341,N_18473,N_18803);
nor UO_1342 (O_1342,N_18553,N_19866);
or UO_1343 (O_1343,N_19717,N_18242);
nand UO_1344 (O_1344,N_19363,N_19545);
nor UO_1345 (O_1345,N_18572,N_19537);
or UO_1346 (O_1346,N_18919,N_19928);
and UO_1347 (O_1347,N_18117,N_19372);
xor UO_1348 (O_1348,N_18432,N_19892);
nand UO_1349 (O_1349,N_18249,N_18993);
nor UO_1350 (O_1350,N_19635,N_19739);
nand UO_1351 (O_1351,N_18963,N_19711);
nand UO_1352 (O_1352,N_18799,N_19354);
nor UO_1353 (O_1353,N_18976,N_18168);
xor UO_1354 (O_1354,N_19277,N_18650);
or UO_1355 (O_1355,N_18429,N_19729);
or UO_1356 (O_1356,N_19678,N_18469);
nor UO_1357 (O_1357,N_18605,N_19092);
xnor UO_1358 (O_1358,N_18593,N_19356);
nand UO_1359 (O_1359,N_19857,N_18540);
or UO_1360 (O_1360,N_18597,N_19041);
and UO_1361 (O_1361,N_18260,N_19472);
xor UO_1362 (O_1362,N_18271,N_19225);
nand UO_1363 (O_1363,N_18147,N_19412);
or UO_1364 (O_1364,N_18271,N_19987);
or UO_1365 (O_1365,N_19813,N_19881);
nand UO_1366 (O_1366,N_18854,N_19054);
nor UO_1367 (O_1367,N_19052,N_19425);
and UO_1368 (O_1368,N_18784,N_19898);
nand UO_1369 (O_1369,N_18995,N_19857);
xor UO_1370 (O_1370,N_18857,N_19808);
and UO_1371 (O_1371,N_18248,N_19931);
nor UO_1372 (O_1372,N_18624,N_18304);
nand UO_1373 (O_1373,N_19953,N_19739);
nor UO_1374 (O_1374,N_18886,N_18507);
and UO_1375 (O_1375,N_18548,N_18235);
nand UO_1376 (O_1376,N_18267,N_19657);
and UO_1377 (O_1377,N_19332,N_18013);
nor UO_1378 (O_1378,N_18596,N_18794);
or UO_1379 (O_1379,N_18545,N_18538);
and UO_1380 (O_1380,N_19503,N_19404);
and UO_1381 (O_1381,N_19126,N_19899);
xnor UO_1382 (O_1382,N_18686,N_18423);
nor UO_1383 (O_1383,N_19600,N_19996);
and UO_1384 (O_1384,N_18351,N_19142);
nand UO_1385 (O_1385,N_19767,N_18292);
xnor UO_1386 (O_1386,N_18921,N_19598);
nand UO_1387 (O_1387,N_19264,N_19155);
nor UO_1388 (O_1388,N_19977,N_19353);
nor UO_1389 (O_1389,N_19160,N_18850);
xor UO_1390 (O_1390,N_18295,N_18178);
nor UO_1391 (O_1391,N_19216,N_18318);
xnor UO_1392 (O_1392,N_18280,N_18301);
nand UO_1393 (O_1393,N_19381,N_18247);
xor UO_1394 (O_1394,N_18504,N_18710);
and UO_1395 (O_1395,N_19832,N_18392);
and UO_1396 (O_1396,N_18576,N_18419);
or UO_1397 (O_1397,N_18233,N_19516);
nand UO_1398 (O_1398,N_18594,N_19273);
nand UO_1399 (O_1399,N_19218,N_19539);
nand UO_1400 (O_1400,N_19402,N_18160);
or UO_1401 (O_1401,N_18240,N_18461);
or UO_1402 (O_1402,N_19678,N_19439);
nor UO_1403 (O_1403,N_19712,N_18781);
and UO_1404 (O_1404,N_18385,N_19822);
and UO_1405 (O_1405,N_19965,N_19373);
nor UO_1406 (O_1406,N_18007,N_18188);
nor UO_1407 (O_1407,N_19801,N_19634);
nor UO_1408 (O_1408,N_19210,N_19574);
nand UO_1409 (O_1409,N_18118,N_18365);
and UO_1410 (O_1410,N_19593,N_18020);
nor UO_1411 (O_1411,N_19233,N_19701);
xnor UO_1412 (O_1412,N_19676,N_19551);
xor UO_1413 (O_1413,N_19244,N_18670);
nor UO_1414 (O_1414,N_19255,N_19128);
or UO_1415 (O_1415,N_19308,N_18706);
nand UO_1416 (O_1416,N_19768,N_18130);
or UO_1417 (O_1417,N_19780,N_18066);
and UO_1418 (O_1418,N_19105,N_18917);
xor UO_1419 (O_1419,N_19148,N_19157);
and UO_1420 (O_1420,N_18768,N_19439);
xnor UO_1421 (O_1421,N_18672,N_18616);
and UO_1422 (O_1422,N_18933,N_18149);
and UO_1423 (O_1423,N_19145,N_19888);
and UO_1424 (O_1424,N_18809,N_18840);
xor UO_1425 (O_1425,N_19328,N_18518);
xor UO_1426 (O_1426,N_18710,N_18514);
nand UO_1427 (O_1427,N_19896,N_18048);
and UO_1428 (O_1428,N_19878,N_18719);
nand UO_1429 (O_1429,N_18295,N_18751);
and UO_1430 (O_1430,N_19856,N_19171);
nand UO_1431 (O_1431,N_19335,N_19008);
xnor UO_1432 (O_1432,N_18873,N_18535);
and UO_1433 (O_1433,N_18252,N_19120);
xnor UO_1434 (O_1434,N_18691,N_18236);
and UO_1435 (O_1435,N_19028,N_18552);
nand UO_1436 (O_1436,N_18060,N_19165);
and UO_1437 (O_1437,N_18418,N_18954);
and UO_1438 (O_1438,N_19803,N_18946);
xnor UO_1439 (O_1439,N_19192,N_19385);
and UO_1440 (O_1440,N_19283,N_19935);
xnor UO_1441 (O_1441,N_19948,N_18118);
or UO_1442 (O_1442,N_19894,N_19238);
nand UO_1443 (O_1443,N_19841,N_18278);
and UO_1444 (O_1444,N_19932,N_18802);
nand UO_1445 (O_1445,N_19513,N_18673);
xor UO_1446 (O_1446,N_18873,N_19149);
or UO_1447 (O_1447,N_19716,N_19878);
xor UO_1448 (O_1448,N_19163,N_19929);
and UO_1449 (O_1449,N_18628,N_18658);
and UO_1450 (O_1450,N_18465,N_19177);
xor UO_1451 (O_1451,N_18937,N_18948);
or UO_1452 (O_1452,N_19554,N_19848);
and UO_1453 (O_1453,N_18383,N_19807);
or UO_1454 (O_1454,N_19859,N_19414);
or UO_1455 (O_1455,N_18548,N_19793);
nor UO_1456 (O_1456,N_18858,N_18551);
xnor UO_1457 (O_1457,N_19851,N_18880);
and UO_1458 (O_1458,N_19887,N_18570);
nor UO_1459 (O_1459,N_19764,N_19013);
nand UO_1460 (O_1460,N_18333,N_19237);
nor UO_1461 (O_1461,N_19707,N_18946);
or UO_1462 (O_1462,N_18972,N_19587);
xnor UO_1463 (O_1463,N_19297,N_19779);
nor UO_1464 (O_1464,N_19996,N_19326);
xor UO_1465 (O_1465,N_18740,N_19592);
xor UO_1466 (O_1466,N_19457,N_18393);
xnor UO_1467 (O_1467,N_18871,N_18720);
nand UO_1468 (O_1468,N_19503,N_18684);
nand UO_1469 (O_1469,N_19038,N_19528);
nor UO_1470 (O_1470,N_18747,N_18060);
nor UO_1471 (O_1471,N_18049,N_19051);
nand UO_1472 (O_1472,N_19970,N_18264);
nor UO_1473 (O_1473,N_19934,N_18609);
nor UO_1474 (O_1474,N_18016,N_18031);
or UO_1475 (O_1475,N_19172,N_19236);
nor UO_1476 (O_1476,N_18536,N_18855);
nor UO_1477 (O_1477,N_19839,N_18747);
or UO_1478 (O_1478,N_18766,N_19899);
and UO_1479 (O_1479,N_19538,N_18549);
or UO_1480 (O_1480,N_18279,N_19316);
nor UO_1481 (O_1481,N_18042,N_18348);
nor UO_1482 (O_1482,N_18549,N_18688);
nor UO_1483 (O_1483,N_18164,N_19433);
nor UO_1484 (O_1484,N_18475,N_19516);
nor UO_1485 (O_1485,N_19576,N_18751);
and UO_1486 (O_1486,N_18946,N_18343);
or UO_1487 (O_1487,N_18451,N_19641);
nand UO_1488 (O_1488,N_19305,N_19550);
xor UO_1489 (O_1489,N_18420,N_18278);
nor UO_1490 (O_1490,N_19881,N_19445);
nand UO_1491 (O_1491,N_19499,N_19955);
and UO_1492 (O_1492,N_18828,N_18211);
xor UO_1493 (O_1493,N_18380,N_19454);
nand UO_1494 (O_1494,N_19675,N_18439);
nor UO_1495 (O_1495,N_19513,N_19538);
and UO_1496 (O_1496,N_18542,N_19014);
nand UO_1497 (O_1497,N_18717,N_18837);
or UO_1498 (O_1498,N_19391,N_19896);
xor UO_1499 (O_1499,N_19222,N_19264);
nor UO_1500 (O_1500,N_19037,N_19049);
nand UO_1501 (O_1501,N_19504,N_18687);
and UO_1502 (O_1502,N_19876,N_18727);
xor UO_1503 (O_1503,N_19531,N_19053);
or UO_1504 (O_1504,N_19953,N_18977);
or UO_1505 (O_1505,N_18546,N_18582);
and UO_1506 (O_1506,N_18414,N_19097);
xnor UO_1507 (O_1507,N_19941,N_19642);
or UO_1508 (O_1508,N_18611,N_18182);
nor UO_1509 (O_1509,N_18226,N_18995);
or UO_1510 (O_1510,N_18201,N_18314);
xor UO_1511 (O_1511,N_19348,N_18736);
and UO_1512 (O_1512,N_18098,N_18187);
and UO_1513 (O_1513,N_19881,N_19429);
or UO_1514 (O_1514,N_18871,N_18249);
and UO_1515 (O_1515,N_18772,N_18265);
nand UO_1516 (O_1516,N_19428,N_19781);
xnor UO_1517 (O_1517,N_19779,N_19086);
and UO_1518 (O_1518,N_18617,N_18685);
or UO_1519 (O_1519,N_19102,N_19303);
nand UO_1520 (O_1520,N_19689,N_18421);
and UO_1521 (O_1521,N_18475,N_18339);
or UO_1522 (O_1522,N_18635,N_18864);
or UO_1523 (O_1523,N_18661,N_18656);
and UO_1524 (O_1524,N_19536,N_19598);
or UO_1525 (O_1525,N_19670,N_18380);
xnor UO_1526 (O_1526,N_18599,N_18893);
nand UO_1527 (O_1527,N_18733,N_18900);
and UO_1528 (O_1528,N_19346,N_18503);
nor UO_1529 (O_1529,N_19625,N_18928);
and UO_1530 (O_1530,N_18725,N_19372);
nor UO_1531 (O_1531,N_18365,N_18461);
nand UO_1532 (O_1532,N_18211,N_18920);
and UO_1533 (O_1533,N_18814,N_18186);
nand UO_1534 (O_1534,N_19733,N_18916);
and UO_1535 (O_1535,N_18657,N_18783);
or UO_1536 (O_1536,N_18136,N_18372);
xor UO_1537 (O_1537,N_18188,N_18818);
and UO_1538 (O_1538,N_19452,N_18890);
or UO_1539 (O_1539,N_19331,N_18218);
xnor UO_1540 (O_1540,N_19847,N_19455);
nor UO_1541 (O_1541,N_19905,N_18448);
or UO_1542 (O_1542,N_19764,N_19024);
xnor UO_1543 (O_1543,N_18984,N_19377);
nand UO_1544 (O_1544,N_19034,N_18750);
or UO_1545 (O_1545,N_19469,N_18783);
or UO_1546 (O_1546,N_18530,N_19802);
and UO_1547 (O_1547,N_18438,N_19058);
xor UO_1548 (O_1548,N_18194,N_19751);
nand UO_1549 (O_1549,N_18322,N_18009);
and UO_1550 (O_1550,N_18536,N_19117);
or UO_1551 (O_1551,N_18659,N_18430);
nand UO_1552 (O_1552,N_18218,N_19205);
xnor UO_1553 (O_1553,N_19432,N_19279);
or UO_1554 (O_1554,N_18659,N_19270);
nor UO_1555 (O_1555,N_19649,N_19526);
or UO_1556 (O_1556,N_18346,N_18484);
xnor UO_1557 (O_1557,N_19989,N_19981);
xnor UO_1558 (O_1558,N_18319,N_18313);
and UO_1559 (O_1559,N_18379,N_19025);
nor UO_1560 (O_1560,N_19628,N_18065);
or UO_1561 (O_1561,N_18126,N_19224);
xnor UO_1562 (O_1562,N_19759,N_18387);
or UO_1563 (O_1563,N_18697,N_18252);
xnor UO_1564 (O_1564,N_18049,N_19328);
or UO_1565 (O_1565,N_18858,N_19030);
xnor UO_1566 (O_1566,N_18476,N_19142);
and UO_1567 (O_1567,N_19262,N_19543);
or UO_1568 (O_1568,N_19346,N_18497);
nand UO_1569 (O_1569,N_19582,N_19336);
xnor UO_1570 (O_1570,N_18710,N_19558);
or UO_1571 (O_1571,N_18569,N_19279);
and UO_1572 (O_1572,N_19691,N_18768);
and UO_1573 (O_1573,N_19785,N_18085);
nand UO_1574 (O_1574,N_18401,N_19982);
xor UO_1575 (O_1575,N_18989,N_18710);
or UO_1576 (O_1576,N_18723,N_18412);
and UO_1577 (O_1577,N_18224,N_19660);
nand UO_1578 (O_1578,N_19172,N_19898);
and UO_1579 (O_1579,N_19037,N_18363);
nor UO_1580 (O_1580,N_19283,N_19096);
xor UO_1581 (O_1581,N_18152,N_18151);
xor UO_1582 (O_1582,N_18786,N_18388);
xor UO_1583 (O_1583,N_19757,N_18513);
or UO_1584 (O_1584,N_19202,N_19764);
or UO_1585 (O_1585,N_19629,N_19417);
or UO_1586 (O_1586,N_18222,N_19017);
or UO_1587 (O_1587,N_19318,N_18693);
nor UO_1588 (O_1588,N_19501,N_18170);
nand UO_1589 (O_1589,N_19333,N_19215);
or UO_1590 (O_1590,N_18014,N_19594);
and UO_1591 (O_1591,N_19232,N_18204);
xnor UO_1592 (O_1592,N_18556,N_18498);
and UO_1593 (O_1593,N_18886,N_18706);
nor UO_1594 (O_1594,N_18077,N_18708);
nand UO_1595 (O_1595,N_18897,N_19469);
and UO_1596 (O_1596,N_19123,N_19743);
nor UO_1597 (O_1597,N_18253,N_19175);
xnor UO_1598 (O_1598,N_18509,N_18073);
and UO_1599 (O_1599,N_19335,N_19918);
xnor UO_1600 (O_1600,N_19055,N_18964);
xor UO_1601 (O_1601,N_19016,N_19077);
or UO_1602 (O_1602,N_18845,N_18069);
or UO_1603 (O_1603,N_18543,N_19956);
nand UO_1604 (O_1604,N_19479,N_18631);
nor UO_1605 (O_1605,N_18207,N_18902);
nand UO_1606 (O_1606,N_18540,N_18183);
or UO_1607 (O_1607,N_18436,N_19138);
or UO_1608 (O_1608,N_18436,N_18475);
and UO_1609 (O_1609,N_19585,N_18454);
or UO_1610 (O_1610,N_18102,N_18192);
nand UO_1611 (O_1611,N_19435,N_18833);
xor UO_1612 (O_1612,N_18323,N_19541);
nand UO_1613 (O_1613,N_19949,N_19617);
nor UO_1614 (O_1614,N_18026,N_18594);
nand UO_1615 (O_1615,N_18084,N_19088);
and UO_1616 (O_1616,N_18751,N_18205);
nor UO_1617 (O_1617,N_19550,N_19308);
nand UO_1618 (O_1618,N_18963,N_18845);
nor UO_1619 (O_1619,N_19216,N_19331);
xor UO_1620 (O_1620,N_19444,N_19218);
nor UO_1621 (O_1621,N_19941,N_18947);
xnor UO_1622 (O_1622,N_18435,N_19972);
xor UO_1623 (O_1623,N_18374,N_18511);
nor UO_1624 (O_1624,N_18781,N_18819);
nand UO_1625 (O_1625,N_19792,N_18325);
nor UO_1626 (O_1626,N_18230,N_18781);
nand UO_1627 (O_1627,N_18739,N_19167);
and UO_1628 (O_1628,N_18056,N_19725);
and UO_1629 (O_1629,N_18255,N_18516);
nand UO_1630 (O_1630,N_19942,N_18627);
and UO_1631 (O_1631,N_19803,N_19948);
nand UO_1632 (O_1632,N_19105,N_19963);
and UO_1633 (O_1633,N_18332,N_19619);
xor UO_1634 (O_1634,N_18931,N_18202);
nand UO_1635 (O_1635,N_19830,N_19729);
nand UO_1636 (O_1636,N_19608,N_19108);
xor UO_1637 (O_1637,N_18183,N_19064);
or UO_1638 (O_1638,N_18576,N_18244);
xnor UO_1639 (O_1639,N_19059,N_18622);
or UO_1640 (O_1640,N_19410,N_19405);
or UO_1641 (O_1641,N_19037,N_19186);
nand UO_1642 (O_1642,N_18920,N_18201);
nor UO_1643 (O_1643,N_18626,N_19441);
or UO_1644 (O_1644,N_18689,N_18300);
or UO_1645 (O_1645,N_18411,N_18571);
and UO_1646 (O_1646,N_19922,N_19226);
and UO_1647 (O_1647,N_19315,N_18853);
or UO_1648 (O_1648,N_19281,N_19651);
or UO_1649 (O_1649,N_19246,N_18312);
nor UO_1650 (O_1650,N_18775,N_19805);
and UO_1651 (O_1651,N_19302,N_19205);
nand UO_1652 (O_1652,N_18362,N_19723);
and UO_1653 (O_1653,N_19387,N_19066);
xnor UO_1654 (O_1654,N_18903,N_19120);
nand UO_1655 (O_1655,N_18585,N_18968);
xor UO_1656 (O_1656,N_19002,N_18763);
and UO_1657 (O_1657,N_18402,N_18205);
nor UO_1658 (O_1658,N_18202,N_18617);
xnor UO_1659 (O_1659,N_19235,N_19938);
or UO_1660 (O_1660,N_19530,N_19531);
or UO_1661 (O_1661,N_19208,N_18673);
and UO_1662 (O_1662,N_19593,N_19185);
nor UO_1663 (O_1663,N_18814,N_19806);
nor UO_1664 (O_1664,N_19746,N_18764);
nor UO_1665 (O_1665,N_18616,N_18687);
xnor UO_1666 (O_1666,N_19393,N_19888);
or UO_1667 (O_1667,N_19161,N_19265);
xnor UO_1668 (O_1668,N_18370,N_18905);
nand UO_1669 (O_1669,N_19334,N_19055);
or UO_1670 (O_1670,N_18425,N_18373);
xor UO_1671 (O_1671,N_18610,N_19647);
or UO_1672 (O_1672,N_19917,N_18307);
nand UO_1673 (O_1673,N_19249,N_18582);
or UO_1674 (O_1674,N_18077,N_18126);
nor UO_1675 (O_1675,N_18344,N_18337);
and UO_1676 (O_1676,N_19707,N_19871);
and UO_1677 (O_1677,N_18846,N_18840);
and UO_1678 (O_1678,N_19727,N_18152);
or UO_1679 (O_1679,N_18792,N_18261);
xnor UO_1680 (O_1680,N_19648,N_18653);
xor UO_1681 (O_1681,N_18305,N_19370);
or UO_1682 (O_1682,N_19855,N_19623);
and UO_1683 (O_1683,N_19257,N_18150);
xnor UO_1684 (O_1684,N_19990,N_18924);
or UO_1685 (O_1685,N_19004,N_18118);
nor UO_1686 (O_1686,N_18984,N_19647);
xnor UO_1687 (O_1687,N_18846,N_18752);
xor UO_1688 (O_1688,N_18797,N_19274);
and UO_1689 (O_1689,N_19087,N_19727);
and UO_1690 (O_1690,N_18104,N_19471);
nor UO_1691 (O_1691,N_18494,N_18654);
or UO_1692 (O_1692,N_18505,N_19793);
or UO_1693 (O_1693,N_19344,N_18301);
and UO_1694 (O_1694,N_19818,N_18339);
and UO_1695 (O_1695,N_19640,N_18363);
or UO_1696 (O_1696,N_18523,N_18338);
or UO_1697 (O_1697,N_19991,N_18024);
and UO_1698 (O_1698,N_18486,N_18110);
or UO_1699 (O_1699,N_19528,N_19195);
and UO_1700 (O_1700,N_18315,N_18961);
xor UO_1701 (O_1701,N_18555,N_19459);
xor UO_1702 (O_1702,N_19192,N_18295);
nor UO_1703 (O_1703,N_18818,N_19572);
nand UO_1704 (O_1704,N_19930,N_18862);
or UO_1705 (O_1705,N_18741,N_18143);
xor UO_1706 (O_1706,N_19229,N_19065);
or UO_1707 (O_1707,N_18411,N_18553);
nor UO_1708 (O_1708,N_19756,N_18496);
xor UO_1709 (O_1709,N_19774,N_18546);
nand UO_1710 (O_1710,N_19204,N_19510);
nand UO_1711 (O_1711,N_19348,N_19088);
nand UO_1712 (O_1712,N_19485,N_18862);
or UO_1713 (O_1713,N_19382,N_18518);
nand UO_1714 (O_1714,N_18538,N_18486);
or UO_1715 (O_1715,N_19257,N_18691);
nand UO_1716 (O_1716,N_19180,N_19249);
nand UO_1717 (O_1717,N_19551,N_18758);
and UO_1718 (O_1718,N_19669,N_18021);
nand UO_1719 (O_1719,N_19011,N_19688);
nand UO_1720 (O_1720,N_18246,N_18171);
xnor UO_1721 (O_1721,N_19472,N_19488);
nor UO_1722 (O_1722,N_18960,N_18229);
or UO_1723 (O_1723,N_18350,N_19696);
nor UO_1724 (O_1724,N_18657,N_18789);
nor UO_1725 (O_1725,N_18686,N_19610);
nor UO_1726 (O_1726,N_18007,N_18416);
xor UO_1727 (O_1727,N_19182,N_19371);
nand UO_1728 (O_1728,N_18415,N_18783);
xnor UO_1729 (O_1729,N_19540,N_19732);
nand UO_1730 (O_1730,N_18119,N_19552);
nor UO_1731 (O_1731,N_19668,N_19441);
nor UO_1732 (O_1732,N_19797,N_19397);
or UO_1733 (O_1733,N_18532,N_19817);
nor UO_1734 (O_1734,N_19479,N_18353);
or UO_1735 (O_1735,N_18149,N_18518);
and UO_1736 (O_1736,N_19747,N_18744);
xnor UO_1737 (O_1737,N_18427,N_18489);
xnor UO_1738 (O_1738,N_18657,N_18621);
and UO_1739 (O_1739,N_19345,N_18857);
nand UO_1740 (O_1740,N_18104,N_18376);
nand UO_1741 (O_1741,N_19216,N_19253);
xnor UO_1742 (O_1742,N_19377,N_18553);
nor UO_1743 (O_1743,N_19592,N_19397);
xnor UO_1744 (O_1744,N_19749,N_18277);
or UO_1745 (O_1745,N_19794,N_18048);
and UO_1746 (O_1746,N_18835,N_18281);
and UO_1747 (O_1747,N_18237,N_19558);
or UO_1748 (O_1748,N_19442,N_18410);
nor UO_1749 (O_1749,N_18702,N_19525);
nand UO_1750 (O_1750,N_19520,N_18577);
nor UO_1751 (O_1751,N_19989,N_19455);
nand UO_1752 (O_1752,N_18291,N_18614);
or UO_1753 (O_1753,N_19408,N_19632);
nand UO_1754 (O_1754,N_18007,N_19837);
or UO_1755 (O_1755,N_18325,N_18417);
nand UO_1756 (O_1756,N_19113,N_18783);
nor UO_1757 (O_1757,N_19165,N_19935);
or UO_1758 (O_1758,N_19603,N_18102);
xnor UO_1759 (O_1759,N_18836,N_19067);
nand UO_1760 (O_1760,N_18839,N_18883);
nand UO_1761 (O_1761,N_19352,N_18398);
nor UO_1762 (O_1762,N_19757,N_18543);
nand UO_1763 (O_1763,N_18957,N_18748);
or UO_1764 (O_1764,N_18021,N_18671);
or UO_1765 (O_1765,N_19437,N_18103);
xnor UO_1766 (O_1766,N_19798,N_19078);
nand UO_1767 (O_1767,N_19434,N_19423);
xnor UO_1768 (O_1768,N_18675,N_18913);
or UO_1769 (O_1769,N_19173,N_18242);
nand UO_1770 (O_1770,N_19852,N_19328);
xor UO_1771 (O_1771,N_19900,N_18718);
nor UO_1772 (O_1772,N_19054,N_19042);
or UO_1773 (O_1773,N_18473,N_19007);
or UO_1774 (O_1774,N_19487,N_18362);
and UO_1775 (O_1775,N_18377,N_18910);
or UO_1776 (O_1776,N_19178,N_19484);
or UO_1777 (O_1777,N_19433,N_19607);
and UO_1778 (O_1778,N_19609,N_18936);
xor UO_1779 (O_1779,N_18230,N_18897);
and UO_1780 (O_1780,N_18052,N_18982);
nor UO_1781 (O_1781,N_18555,N_18592);
nand UO_1782 (O_1782,N_18121,N_18506);
and UO_1783 (O_1783,N_19937,N_19476);
xnor UO_1784 (O_1784,N_18230,N_18914);
nor UO_1785 (O_1785,N_19929,N_19382);
or UO_1786 (O_1786,N_18263,N_19273);
nor UO_1787 (O_1787,N_18200,N_18096);
nor UO_1788 (O_1788,N_18394,N_18862);
xnor UO_1789 (O_1789,N_18220,N_18710);
nand UO_1790 (O_1790,N_18406,N_19949);
nand UO_1791 (O_1791,N_19174,N_19222);
nand UO_1792 (O_1792,N_19441,N_18294);
nor UO_1793 (O_1793,N_19807,N_18020);
nand UO_1794 (O_1794,N_19510,N_19176);
nor UO_1795 (O_1795,N_19567,N_19269);
xor UO_1796 (O_1796,N_18858,N_19993);
nand UO_1797 (O_1797,N_18292,N_19790);
nand UO_1798 (O_1798,N_19067,N_18166);
or UO_1799 (O_1799,N_18481,N_18024);
nor UO_1800 (O_1800,N_19759,N_18357);
nand UO_1801 (O_1801,N_18239,N_19899);
nand UO_1802 (O_1802,N_19340,N_19346);
xor UO_1803 (O_1803,N_18384,N_18235);
nand UO_1804 (O_1804,N_19899,N_19445);
nand UO_1805 (O_1805,N_19650,N_19557);
xor UO_1806 (O_1806,N_19954,N_19096);
nor UO_1807 (O_1807,N_18010,N_19330);
xor UO_1808 (O_1808,N_18100,N_18530);
or UO_1809 (O_1809,N_18904,N_19645);
nand UO_1810 (O_1810,N_19870,N_19677);
or UO_1811 (O_1811,N_19813,N_19007);
nand UO_1812 (O_1812,N_18324,N_19558);
and UO_1813 (O_1813,N_19425,N_18920);
nor UO_1814 (O_1814,N_19068,N_18604);
xnor UO_1815 (O_1815,N_19438,N_19028);
nor UO_1816 (O_1816,N_18634,N_19602);
or UO_1817 (O_1817,N_18652,N_19310);
and UO_1818 (O_1818,N_19719,N_19170);
and UO_1819 (O_1819,N_18207,N_19738);
nor UO_1820 (O_1820,N_18308,N_19685);
xor UO_1821 (O_1821,N_18837,N_18591);
and UO_1822 (O_1822,N_18776,N_19001);
or UO_1823 (O_1823,N_19789,N_18018);
xnor UO_1824 (O_1824,N_19326,N_18777);
nand UO_1825 (O_1825,N_19548,N_18215);
nand UO_1826 (O_1826,N_18229,N_18097);
nand UO_1827 (O_1827,N_19024,N_18693);
or UO_1828 (O_1828,N_19895,N_19839);
xor UO_1829 (O_1829,N_18954,N_19533);
xnor UO_1830 (O_1830,N_19359,N_18662);
and UO_1831 (O_1831,N_19638,N_18934);
or UO_1832 (O_1832,N_19271,N_19757);
and UO_1833 (O_1833,N_19054,N_18706);
xor UO_1834 (O_1834,N_19208,N_19132);
xor UO_1835 (O_1835,N_19917,N_18100);
xor UO_1836 (O_1836,N_18000,N_19871);
and UO_1837 (O_1837,N_19735,N_18909);
nor UO_1838 (O_1838,N_18936,N_18999);
and UO_1839 (O_1839,N_19100,N_19486);
nand UO_1840 (O_1840,N_18227,N_19323);
nand UO_1841 (O_1841,N_19928,N_19758);
nor UO_1842 (O_1842,N_19504,N_18874);
nand UO_1843 (O_1843,N_18599,N_18576);
or UO_1844 (O_1844,N_18664,N_19581);
xor UO_1845 (O_1845,N_19755,N_18896);
xnor UO_1846 (O_1846,N_19264,N_19188);
nor UO_1847 (O_1847,N_19844,N_18877);
xnor UO_1848 (O_1848,N_18591,N_18390);
xnor UO_1849 (O_1849,N_18351,N_19734);
nand UO_1850 (O_1850,N_19261,N_19715);
nand UO_1851 (O_1851,N_18954,N_19309);
and UO_1852 (O_1852,N_19030,N_19294);
nor UO_1853 (O_1853,N_19480,N_19624);
nand UO_1854 (O_1854,N_18317,N_19423);
and UO_1855 (O_1855,N_19509,N_19239);
nor UO_1856 (O_1856,N_18360,N_19989);
nor UO_1857 (O_1857,N_18902,N_19496);
nand UO_1858 (O_1858,N_19434,N_19436);
or UO_1859 (O_1859,N_19118,N_18383);
and UO_1860 (O_1860,N_19448,N_18154);
or UO_1861 (O_1861,N_19229,N_18403);
xor UO_1862 (O_1862,N_19754,N_18640);
nand UO_1863 (O_1863,N_18978,N_19989);
nand UO_1864 (O_1864,N_19868,N_19592);
or UO_1865 (O_1865,N_18387,N_18628);
or UO_1866 (O_1866,N_18025,N_18413);
nand UO_1867 (O_1867,N_18409,N_18809);
or UO_1868 (O_1868,N_18990,N_18074);
nor UO_1869 (O_1869,N_19344,N_18806);
and UO_1870 (O_1870,N_19257,N_19480);
or UO_1871 (O_1871,N_18141,N_19446);
nor UO_1872 (O_1872,N_19372,N_18011);
nor UO_1873 (O_1873,N_19144,N_18868);
or UO_1874 (O_1874,N_18143,N_19423);
nor UO_1875 (O_1875,N_19259,N_19544);
xor UO_1876 (O_1876,N_19121,N_19941);
or UO_1877 (O_1877,N_18351,N_18540);
xor UO_1878 (O_1878,N_18909,N_18280);
xnor UO_1879 (O_1879,N_18778,N_18786);
nor UO_1880 (O_1880,N_19596,N_19609);
xor UO_1881 (O_1881,N_19968,N_19934);
and UO_1882 (O_1882,N_19667,N_18735);
xor UO_1883 (O_1883,N_18120,N_18437);
nor UO_1884 (O_1884,N_18716,N_18980);
or UO_1885 (O_1885,N_18790,N_19544);
or UO_1886 (O_1886,N_18466,N_19770);
nand UO_1887 (O_1887,N_19801,N_18058);
nand UO_1888 (O_1888,N_19316,N_19365);
xnor UO_1889 (O_1889,N_18352,N_19736);
nand UO_1890 (O_1890,N_19257,N_19128);
nor UO_1891 (O_1891,N_19963,N_19670);
and UO_1892 (O_1892,N_18077,N_18971);
or UO_1893 (O_1893,N_19537,N_18807);
or UO_1894 (O_1894,N_19550,N_19729);
xnor UO_1895 (O_1895,N_19413,N_19393);
or UO_1896 (O_1896,N_19741,N_19894);
or UO_1897 (O_1897,N_18221,N_18136);
xor UO_1898 (O_1898,N_19862,N_18555);
xnor UO_1899 (O_1899,N_18687,N_19020);
nand UO_1900 (O_1900,N_19757,N_18564);
nand UO_1901 (O_1901,N_19410,N_18076);
or UO_1902 (O_1902,N_19155,N_18866);
xnor UO_1903 (O_1903,N_19555,N_18484);
and UO_1904 (O_1904,N_18025,N_19746);
nand UO_1905 (O_1905,N_18218,N_18873);
or UO_1906 (O_1906,N_19976,N_19055);
nand UO_1907 (O_1907,N_18196,N_19678);
nand UO_1908 (O_1908,N_18783,N_18458);
xor UO_1909 (O_1909,N_18418,N_18116);
and UO_1910 (O_1910,N_18151,N_19407);
xor UO_1911 (O_1911,N_19445,N_19867);
xor UO_1912 (O_1912,N_18682,N_19338);
or UO_1913 (O_1913,N_19728,N_18039);
nor UO_1914 (O_1914,N_19592,N_19640);
and UO_1915 (O_1915,N_18869,N_18681);
nand UO_1916 (O_1916,N_19566,N_19960);
nor UO_1917 (O_1917,N_19251,N_18182);
nand UO_1918 (O_1918,N_18603,N_18964);
xnor UO_1919 (O_1919,N_18887,N_18745);
or UO_1920 (O_1920,N_19636,N_19524);
xor UO_1921 (O_1921,N_19429,N_19984);
xnor UO_1922 (O_1922,N_18643,N_18065);
or UO_1923 (O_1923,N_19294,N_19683);
or UO_1924 (O_1924,N_19519,N_19455);
nand UO_1925 (O_1925,N_19397,N_19879);
xnor UO_1926 (O_1926,N_19030,N_19243);
nand UO_1927 (O_1927,N_18856,N_18438);
nor UO_1928 (O_1928,N_19399,N_18562);
xor UO_1929 (O_1929,N_18942,N_19842);
and UO_1930 (O_1930,N_18702,N_18943);
or UO_1931 (O_1931,N_18589,N_19936);
nor UO_1932 (O_1932,N_19020,N_19206);
and UO_1933 (O_1933,N_18342,N_19103);
or UO_1934 (O_1934,N_18896,N_18954);
xor UO_1935 (O_1935,N_19420,N_18021);
and UO_1936 (O_1936,N_19376,N_19176);
nor UO_1937 (O_1937,N_18960,N_19367);
and UO_1938 (O_1938,N_18541,N_18061);
or UO_1939 (O_1939,N_18633,N_19696);
nand UO_1940 (O_1940,N_19465,N_19422);
xnor UO_1941 (O_1941,N_19273,N_19147);
xor UO_1942 (O_1942,N_19552,N_18594);
xnor UO_1943 (O_1943,N_19709,N_19050);
xnor UO_1944 (O_1944,N_19347,N_18596);
or UO_1945 (O_1945,N_19860,N_19394);
and UO_1946 (O_1946,N_19167,N_19220);
nand UO_1947 (O_1947,N_18117,N_18716);
and UO_1948 (O_1948,N_18172,N_19178);
and UO_1949 (O_1949,N_18012,N_18962);
and UO_1950 (O_1950,N_18907,N_18870);
and UO_1951 (O_1951,N_18080,N_18764);
nand UO_1952 (O_1952,N_18219,N_18575);
nand UO_1953 (O_1953,N_18113,N_18818);
nor UO_1954 (O_1954,N_18307,N_19462);
xor UO_1955 (O_1955,N_19272,N_19375);
and UO_1956 (O_1956,N_18175,N_18180);
nand UO_1957 (O_1957,N_18148,N_18149);
nor UO_1958 (O_1958,N_18150,N_19181);
xnor UO_1959 (O_1959,N_18135,N_18691);
nor UO_1960 (O_1960,N_18913,N_19134);
xnor UO_1961 (O_1961,N_18731,N_18033);
or UO_1962 (O_1962,N_18245,N_19613);
or UO_1963 (O_1963,N_19236,N_19281);
nand UO_1964 (O_1964,N_18872,N_18628);
xnor UO_1965 (O_1965,N_18801,N_18628);
xor UO_1966 (O_1966,N_19138,N_18179);
or UO_1967 (O_1967,N_19054,N_18232);
nor UO_1968 (O_1968,N_18305,N_19600);
and UO_1969 (O_1969,N_18172,N_18773);
or UO_1970 (O_1970,N_18088,N_18327);
nor UO_1971 (O_1971,N_19028,N_19204);
nor UO_1972 (O_1972,N_19979,N_19146);
and UO_1973 (O_1973,N_18699,N_18163);
xnor UO_1974 (O_1974,N_19966,N_19849);
xnor UO_1975 (O_1975,N_19465,N_19590);
or UO_1976 (O_1976,N_19444,N_19816);
nor UO_1977 (O_1977,N_18860,N_19660);
or UO_1978 (O_1978,N_18165,N_19456);
nor UO_1979 (O_1979,N_19233,N_18518);
or UO_1980 (O_1980,N_18149,N_18302);
nor UO_1981 (O_1981,N_19844,N_19379);
nand UO_1982 (O_1982,N_18412,N_18633);
xnor UO_1983 (O_1983,N_18326,N_19068);
xor UO_1984 (O_1984,N_19107,N_18352);
or UO_1985 (O_1985,N_18344,N_18370);
or UO_1986 (O_1986,N_18117,N_19045);
nor UO_1987 (O_1987,N_18573,N_18847);
nor UO_1988 (O_1988,N_18640,N_18762);
nand UO_1989 (O_1989,N_19652,N_19917);
and UO_1990 (O_1990,N_19877,N_19951);
xor UO_1991 (O_1991,N_19430,N_19736);
or UO_1992 (O_1992,N_19954,N_19720);
nand UO_1993 (O_1993,N_19191,N_19445);
and UO_1994 (O_1994,N_19868,N_19561);
nand UO_1995 (O_1995,N_18586,N_18892);
nor UO_1996 (O_1996,N_19981,N_18950);
and UO_1997 (O_1997,N_18016,N_18743);
and UO_1998 (O_1998,N_18123,N_19621);
nor UO_1999 (O_1999,N_18945,N_18814);
nand UO_2000 (O_2000,N_19539,N_19570);
or UO_2001 (O_2001,N_19859,N_18900);
nor UO_2002 (O_2002,N_19075,N_19650);
xnor UO_2003 (O_2003,N_18586,N_19426);
and UO_2004 (O_2004,N_18179,N_18049);
nor UO_2005 (O_2005,N_18474,N_19789);
nand UO_2006 (O_2006,N_18072,N_19158);
nand UO_2007 (O_2007,N_18952,N_19349);
nand UO_2008 (O_2008,N_19245,N_19327);
and UO_2009 (O_2009,N_18250,N_19980);
xor UO_2010 (O_2010,N_18555,N_19779);
nand UO_2011 (O_2011,N_18811,N_19042);
or UO_2012 (O_2012,N_18534,N_18389);
xnor UO_2013 (O_2013,N_18909,N_18924);
and UO_2014 (O_2014,N_18069,N_18522);
and UO_2015 (O_2015,N_19262,N_19341);
and UO_2016 (O_2016,N_18596,N_18054);
xor UO_2017 (O_2017,N_19944,N_19524);
and UO_2018 (O_2018,N_19291,N_19759);
and UO_2019 (O_2019,N_18285,N_19171);
nand UO_2020 (O_2020,N_19967,N_19531);
nand UO_2021 (O_2021,N_19560,N_19964);
and UO_2022 (O_2022,N_18121,N_18696);
nor UO_2023 (O_2023,N_19958,N_19262);
nor UO_2024 (O_2024,N_18245,N_19579);
nand UO_2025 (O_2025,N_18512,N_19941);
nor UO_2026 (O_2026,N_19015,N_19358);
nor UO_2027 (O_2027,N_19999,N_18236);
xnor UO_2028 (O_2028,N_18260,N_19925);
or UO_2029 (O_2029,N_18269,N_18558);
and UO_2030 (O_2030,N_18407,N_18542);
and UO_2031 (O_2031,N_18686,N_19166);
nand UO_2032 (O_2032,N_18582,N_18139);
and UO_2033 (O_2033,N_18750,N_19759);
nor UO_2034 (O_2034,N_19751,N_18914);
or UO_2035 (O_2035,N_19703,N_19251);
and UO_2036 (O_2036,N_19463,N_19150);
or UO_2037 (O_2037,N_18195,N_18397);
nor UO_2038 (O_2038,N_18494,N_19544);
and UO_2039 (O_2039,N_19207,N_18011);
nand UO_2040 (O_2040,N_18857,N_19358);
xnor UO_2041 (O_2041,N_18225,N_19326);
xnor UO_2042 (O_2042,N_18166,N_19412);
and UO_2043 (O_2043,N_18511,N_18789);
or UO_2044 (O_2044,N_19458,N_19404);
or UO_2045 (O_2045,N_18721,N_18930);
nand UO_2046 (O_2046,N_19718,N_19465);
nand UO_2047 (O_2047,N_18793,N_18944);
or UO_2048 (O_2048,N_18663,N_18818);
xnor UO_2049 (O_2049,N_19622,N_19090);
and UO_2050 (O_2050,N_18495,N_19198);
and UO_2051 (O_2051,N_19235,N_18890);
or UO_2052 (O_2052,N_19970,N_18131);
nor UO_2053 (O_2053,N_19310,N_19798);
nand UO_2054 (O_2054,N_19686,N_18431);
nand UO_2055 (O_2055,N_18239,N_19092);
nand UO_2056 (O_2056,N_19831,N_18901);
or UO_2057 (O_2057,N_18003,N_19634);
and UO_2058 (O_2058,N_19015,N_18362);
nor UO_2059 (O_2059,N_18484,N_19036);
xnor UO_2060 (O_2060,N_19300,N_19821);
xnor UO_2061 (O_2061,N_18825,N_18925);
nor UO_2062 (O_2062,N_19194,N_19290);
xnor UO_2063 (O_2063,N_19341,N_18071);
or UO_2064 (O_2064,N_19228,N_19733);
xor UO_2065 (O_2065,N_19823,N_18912);
or UO_2066 (O_2066,N_19428,N_18656);
and UO_2067 (O_2067,N_18999,N_19085);
and UO_2068 (O_2068,N_19318,N_19771);
and UO_2069 (O_2069,N_19557,N_19764);
nand UO_2070 (O_2070,N_18507,N_19654);
xnor UO_2071 (O_2071,N_18159,N_18171);
or UO_2072 (O_2072,N_18442,N_18237);
xor UO_2073 (O_2073,N_18088,N_18713);
xor UO_2074 (O_2074,N_18554,N_18189);
nand UO_2075 (O_2075,N_18095,N_19115);
xnor UO_2076 (O_2076,N_19108,N_18271);
xor UO_2077 (O_2077,N_19090,N_19302);
or UO_2078 (O_2078,N_18349,N_19605);
nor UO_2079 (O_2079,N_19306,N_19877);
and UO_2080 (O_2080,N_18081,N_18155);
xnor UO_2081 (O_2081,N_19624,N_19973);
nand UO_2082 (O_2082,N_18999,N_19183);
nand UO_2083 (O_2083,N_19892,N_19918);
xor UO_2084 (O_2084,N_18743,N_19095);
nand UO_2085 (O_2085,N_18764,N_18810);
nor UO_2086 (O_2086,N_18977,N_18814);
nand UO_2087 (O_2087,N_19026,N_19372);
nand UO_2088 (O_2088,N_18086,N_18950);
nor UO_2089 (O_2089,N_19357,N_18385);
nand UO_2090 (O_2090,N_19149,N_19240);
nand UO_2091 (O_2091,N_18075,N_18275);
nand UO_2092 (O_2092,N_18325,N_18035);
nor UO_2093 (O_2093,N_19582,N_18606);
and UO_2094 (O_2094,N_18714,N_18374);
or UO_2095 (O_2095,N_18858,N_18657);
nor UO_2096 (O_2096,N_19202,N_19790);
or UO_2097 (O_2097,N_19603,N_18066);
and UO_2098 (O_2098,N_19438,N_18870);
xor UO_2099 (O_2099,N_19639,N_19503);
nand UO_2100 (O_2100,N_18406,N_18649);
nor UO_2101 (O_2101,N_18149,N_18971);
nor UO_2102 (O_2102,N_19216,N_19042);
and UO_2103 (O_2103,N_18894,N_19872);
or UO_2104 (O_2104,N_18214,N_19606);
nor UO_2105 (O_2105,N_19621,N_19905);
xor UO_2106 (O_2106,N_18778,N_19465);
or UO_2107 (O_2107,N_18943,N_19015);
nand UO_2108 (O_2108,N_19444,N_18026);
or UO_2109 (O_2109,N_19156,N_18144);
nor UO_2110 (O_2110,N_18163,N_19831);
or UO_2111 (O_2111,N_18792,N_18905);
and UO_2112 (O_2112,N_18049,N_19814);
or UO_2113 (O_2113,N_19862,N_19791);
xnor UO_2114 (O_2114,N_18231,N_19678);
nor UO_2115 (O_2115,N_18113,N_18062);
xnor UO_2116 (O_2116,N_18387,N_18001);
or UO_2117 (O_2117,N_18411,N_18675);
xnor UO_2118 (O_2118,N_18331,N_18456);
nand UO_2119 (O_2119,N_19104,N_19297);
and UO_2120 (O_2120,N_18181,N_19072);
and UO_2121 (O_2121,N_19432,N_18722);
xnor UO_2122 (O_2122,N_19194,N_19386);
nor UO_2123 (O_2123,N_19903,N_18194);
nor UO_2124 (O_2124,N_19145,N_18092);
and UO_2125 (O_2125,N_19687,N_19115);
and UO_2126 (O_2126,N_19264,N_18282);
xor UO_2127 (O_2127,N_18520,N_19283);
and UO_2128 (O_2128,N_18424,N_18878);
or UO_2129 (O_2129,N_19037,N_18027);
and UO_2130 (O_2130,N_18241,N_19807);
or UO_2131 (O_2131,N_19498,N_19265);
and UO_2132 (O_2132,N_19852,N_18492);
and UO_2133 (O_2133,N_19318,N_19618);
or UO_2134 (O_2134,N_19968,N_18606);
xor UO_2135 (O_2135,N_19632,N_19009);
nand UO_2136 (O_2136,N_18099,N_19874);
nor UO_2137 (O_2137,N_18349,N_18721);
nand UO_2138 (O_2138,N_18791,N_18546);
or UO_2139 (O_2139,N_18701,N_19809);
xor UO_2140 (O_2140,N_18398,N_18219);
or UO_2141 (O_2141,N_18042,N_19150);
and UO_2142 (O_2142,N_19765,N_19550);
nand UO_2143 (O_2143,N_19060,N_18607);
or UO_2144 (O_2144,N_18562,N_19997);
xnor UO_2145 (O_2145,N_19345,N_18992);
or UO_2146 (O_2146,N_18283,N_18090);
or UO_2147 (O_2147,N_18168,N_19998);
nor UO_2148 (O_2148,N_19959,N_18692);
nor UO_2149 (O_2149,N_19977,N_18274);
nand UO_2150 (O_2150,N_19893,N_19812);
or UO_2151 (O_2151,N_18475,N_18455);
nand UO_2152 (O_2152,N_18981,N_19146);
and UO_2153 (O_2153,N_18710,N_19494);
xnor UO_2154 (O_2154,N_19803,N_19830);
nor UO_2155 (O_2155,N_18865,N_18264);
or UO_2156 (O_2156,N_18788,N_18793);
nand UO_2157 (O_2157,N_18717,N_19293);
xnor UO_2158 (O_2158,N_18652,N_19035);
xnor UO_2159 (O_2159,N_18201,N_18309);
and UO_2160 (O_2160,N_18974,N_19867);
nand UO_2161 (O_2161,N_19338,N_18983);
xnor UO_2162 (O_2162,N_19054,N_19899);
and UO_2163 (O_2163,N_19173,N_18951);
xnor UO_2164 (O_2164,N_18260,N_18910);
nor UO_2165 (O_2165,N_19794,N_19630);
and UO_2166 (O_2166,N_19992,N_18316);
nand UO_2167 (O_2167,N_19435,N_18839);
and UO_2168 (O_2168,N_19916,N_19683);
nor UO_2169 (O_2169,N_18683,N_19728);
nand UO_2170 (O_2170,N_18296,N_18327);
xnor UO_2171 (O_2171,N_19625,N_18780);
nand UO_2172 (O_2172,N_18652,N_18376);
and UO_2173 (O_2173,N_18546,N_18788);
xnor UO_2174 (O_2174,N_19685,N_19513);
and UO_2175 (O_2175,N_18358,N_19115);
and UO_2176 (O_2176,N_19585,N_19213);
nand UO_2177 (O_2177,N_19752,N_19331);
nand UO_2178 (O_2178,N_19392,N_18077);
nor UO_2179 (O_2179,N_18440,N_18043);
nand UO_2180 (O_2180,N_19194,N_19262);
or UO_2181 (O_2181,N_19041,N_19497);
nor UO_2182 (O_2182,N_18752,N_18837);
xor UO_2183 (O_2183,N_18283,N_19093);
or UO_2184 (O_2184,N_18979,N_19998);
xnor UO_2185 (O_2185,N_19512,N_19080);
nand UO_2186 (O_2186,N_19487,N_18452);
nand UO_2187 (O_2187,N_18662,N_19925);
xor UO_2188 (O_2188,N_19258,N_18124);
or UO_2189 (O_2189,N_19768,N_19003);
or UO_2190 (O_2190,N_18193,N_19827);
xor UO_2191 (O_2191,N_19919,N_18372);
and UO_2192 (O_2192,N_18311,N_19213);
xor UO_2193 (O_2193,N_19627,N_19454);
nor UO_2194 (O_2194,N_19045,N_19471);
xnor UO_2195 (O_2195,N_18885,N_18608);
and UO_2196 (O_2196,N_19007,N_18508);
xor UO_2197 (O_2197,N_18364,N_18793);
nand UO_2198 (O_2198,N_19578,N_18030);
and UO_2199 (O_2199,N_18546,N_19364);
xor UO_2200 (O_2200,N_18970,N_19039);
nor UO_2201 (O_2201,N_19901,N_19485);
nand UO_2202 (O_2202,N_18126,N_19820);
or UO_2203 (O_2203,N_18700,N_18274);
or UO_2204 (O_2204,N_19692,N_18406);
xnor UO_2205 (O_2205,N_19334,N_19022);
nand UO_2206 (O_2206,N_19833,N_19613);
or UO_2207 (O_2207,N_18455,N_19080);
xnor UO_2208 (O_2208,N_18471,N_19064);
or UO_2209 (O_2209,N_19762,N_18083);
and UO_2210 (O_2210,N_19112,N_19360);
xor UO_2211 (O_2211,N_18490,N_18255);
nor UO_2212 (O_2212,N_18896,N_19276);
or UO_2213 (O_2213,N_19394,N_19731);
nor UO_2214 (O_2214,N_19869,N_19457);
nor UO_2215 (O_2215,N_19751,N_19902);
nor UO_2216 (O_2216,N_19778,N_19863);
nand UO_2217 (O_2217,N_19030,N_18753);
and UO_2218 (O_2218,N_18358,N_18286);
xnor UO_2219 (O_2219,N_18484,N_19269);
nor UO_2220 (O_2220,N_18023,N_19123);
and UO_2221 (O_2221,N_18261,N_18062);
xnor UO_2222 (O_2222,N_19283,N_19874);
or UO_2223 (O_2223,N_18197,N_19673);
xnor UO_2224 (O_2224,N_18141,N_18530);
xor UO_2225 (O_2225,N_18952,N_19988);
xor UO_2226 (O_2226,N_19399,N_19405);
nand UO_2227 (O_2227,N_19493,N_19609);
nand UO_2228 (O_2228,N_19321,N_18486);
or UO_2229 (O_2229,N_19684,N_19710);
and UO_2230 (O_2230,N_18343,N_18061);
nor UO_2231 (O_2231,N_18861,N_18185);
nor UO_2232 (O_2232,N_18704,N_18639);
or UO_2233 (O_2233,N_18143,N_18578);
nor UO_2234 (O_2234,N_18225,N_19144);
nor UO_2235 (O_2235,N_18973,N_18257);
nand UO_2236 (O_2236,N_19788,N_18219);
and UO_2237 (O_2237,N_19219,N_19997);
nand UO_2238 (O_2238,N_18707,N_19282);
and UO_2239 (O_2239,N_19277,N_18864);
xnor UO_2240 (O_2240,N_18831,N_18643);
nor UO_2241 (O_2241,N_18531,N_19801);
or UO_2242 (O_2242,N_19779,N_18934);
xnor UO_2243 (O_2243,N_19538,N_18759);
nand UO_2244 (O_2244,N_18628,N_19277);
and UO_2245 (O_2245,N_19490,N_19905);
or UO_2246 (O_2246,N_19980,N_19467);
or UO_2247 (O_2247,N_19304,N_18123);
nand UO_2248 (O_2248,N_18898,N_18459);
nand UO_2249 (O_2249,N_18396,N_19676);
nand UO_2250 (O_2250,N_19823,N_18276);
or UO_2251 (O_2251,N_18761,N_18677);
xnor UO_2252 (O_2252,N_18505,N_18759);
nand UO_2253 (O_2253,N_18125,N_19612);
nor UO_2254 (O_2254,N_19598,N_19257);
xor UO_2255 (O_2255,N_18488,N_19445);
or UO_2256 (O_2256,N_18451,N_18807);
and UO_2257 (O_2257,N_19473,N_19299);
nor UO_2258 (O_2258,N_19361,N_19020);
or UO_2259 (O_2259,N_18464,N_19181);
or UO_2260 (O_2260,N_19361,N_18709);
nor UO_2261 (O_2261,N_18190,N_18131);
and UO_2262 (O_2262,N_18694,N_18638);
nand UO_2263 (O_2263,N_18080,N_18950);
xnor UO_2264 (O_2264,N_19847,N_18053);
nand UO_2265 (O_2265,N_18355,N_18583);
or UO_2266 (O_2266,N_19458,N_18347);
nor UO_2267 (O_2267,N_18962,N_19919);
nor UO_2268 (O_2268,N_18405,N_19246);
nand UO_2269 (O_2269,N_18045,N_19255);
and UO_2270 (O_2270,N_18362,N_19067);
nor UO_2271 (O_2271,N_18759,N_19119);
and UO_2272 (O_2272,N_18565,N_19340);
nor UO_2273 (O_2273,N_19740,N_18897);
nand UO_2274 (O_2274,N_18599,N_18608);
nor UO_2275 (O_2275,N_19877,N_18620);
nor UO_2276 (O_2276,N_18316,N_19008);
xnor UO_2277 (O_2277,N_18687,N_19377);
nand UO_2278 (O_2278,N_18883,N_19284);
or UO_2279 (O_2279,N_18550,N_18693);
and UO_2280 (O_2280,N_19830,N_19408);
and UO_2281 (O_2281,N_19711,N_19676);
xor UO_2282 (O_2282,N_19134,N_19938);
or UO_2283 (O_2283,N_19954,N_19712);
and UO_2284 (O_2284,N_19430,N_19980);
nand UO_2285 (O_2285,N_18081,N_18660);
and UO_2286 (O_2286,N_18088,N_18909);
or UO_2287 (O_2287,N_18008,N_19151);
nor UO_2288 (O_2288,N_18458,N_19537);
nand UO_2289 (O_2289,N_18467,N_19901);
and UO_2290 (O_2290,N_19051,N_19440);
and UO_2291 (O_2291,N_19186,N_19446);
nor UO_2292 (O_2292,N_19404,N_18498);
or UO_2293 (O_2293,N_19623,N_19194);
and UO_2294 (O_2294,N_18045,N_19197);
xnor UO_2295 (O_2295,N_19269,N_19137);
or UO_2296 (O_2296,N_19592,N_19641);
or UO_2297 (O_2297,N_18099,N_19373);
or UO_2298 (O_2298,N_18797,N_18199);
nand UO_2299 (O_2299,N_18921,N_19667);
and UO_2300 (O_2300,N_18184,N_18096);
nand UO_2301 (O_2301,N_19897,N_18446);
nand UO_2302 (O_2302,N_19121,N_18142);
nor UO_2303 (O_2303,N_19034,N_18785);
xor UO_2304 (O_2304,N_19470,N_19112);
nor UO_2305 (O_2305,N_19160,N_18218);
or UO_2306 (O_2306,N_18935,N_19794);
and UO_2307 (O_2307,N_19500,N_19772);
xnor UO_2308 (O_2308,N_19699,N_18588);
nor UO_2309 (O_2309,N_19456,N_19130);
xnor UO_2310 (O_2310,N_19201,N_18323);
nor UO_2311 (O_2311,N_19591,N_18961);
or UO_2312 (O_2312,N_18044,N_19258);
or UO_2313 (O_2313,N_18578,N_19098);
nor UO_2314 (O_2314,N_18487,N_18305);
and UO_2315 (O_2315,N_19045,N_19923);
nand UO_2316 (O_2316,N_18082,N_19875);
or UO_2317 (O_2317,N_19797,N_18700);
xnor UO_2318 (O_2318,N_18219,N_18813);
nand UO_2319 (O_2319,N_18940,N_18517);
xnor UO_2320 (O_2320,N_18163,N_18102);
or UO_2321 (O_2321,N_19940,N_19808);
and UO_2322 (O_2322,N_19398,N_18671);
nand UO_2323 (O_2323,N_19638,N_18244);
nand UO_2324 (O_2324,N_19422,N_18831);
nor UO_2325 (O_2325,N_19700,N_18443);
xor UO_2326 (O_2326,N_18994,N_18066);
nor UO_2327 (O_2327,N_19982,N_19827);
and UO_2328 (O_2328,N_18185,N_19345);
or UO_2329 (O_2329,N_19404,N_18675);
nor UO_2330 (O_2330,N_19605,N_18810);
nand UO_2331 (O_2331,N_18337,N_18814);
nand UO_2332 (O_2332,N_19536,N_19358);
nand UO_2333 (O_2333,N_19127,N_19988);
xnor UO_2334 (O_2334,N_19435,N_18688);
and UO_2335 (O_2335,N_18834,N_19031);
or UO_2336 (O_2336,N_19756,N_19322);
nand UO_2337 (O_2337,N_19979,N_19784);
nor UO_2338 (O_2338,N_19461,N_19761);
nand UO_2339 (O_2339,N_18086,N_19157);
nor UO_2340 (O_2340,N_19049,N_18425);
nor UO_2341 (O_2341,N_19550,N_19661);
or UO_2342 (O_2342,N_18076,N_18591);
and UO_2343 (O_2343,N_19953,N_19126);
and UO_2344 (O_2344,N_18159,N_18743);
nand UO_2345 (O_2345,N_18809,N_19775);
or UO_2346 (O_2346,N_19383,N_18683);
xnor UO_2347 (O_2347,N_18418,N_18137);
and UO_2348 (O_2348,N_19626,N_19471);
and UO_2349 (O_2349,N_19505,N_18745);
or UO_2350 (O_2350,N_18964,N_19414);
and UO_2351 (O_2351,N_18030,N_19385);
xnor UO_2352 (O_2352,N_19255,N_19958);
or UO_2353 (O_2353,N_18260,N_18173);
nor UO_2354 (O_2354,N_19853,N_19590);
or UO_2355 (O_2355,N_18051,N_18047);
and UO_2356 (O_2356,N_18281,N_19600);
nor UO_2357 (O_2357,N_18564,N_19621);
xnor UO_2358 (O_2358,N_18904,N_18246);
or UO_2359 (O_2359,N_19831,N_18552);
xor UO_2360 (O_2360,N_18498,N_18191);
and UO_2361 (O_2361,N_18382,N_19880);
and UO_2362 (O_2362,N_19660,N_19307);
or UO_2363 (O_2363,N_18972,N_19153);
xor UO_2364 (O_2364,N_18027,N_19035);
or UO_2365 (O_2365,N_18812,N_18621);
xor UO_2366 (O_2366,N_18677,N_19423);
nor UO_2367 (O_2367,N_18654,N_19127);
nor UO_2368 (O_2368,N_19408,N_18699);
and UO_2369 (O_2369,N_18889,N_18682);
xnor UO_2370 (O_2370,N_19943,N_18159);
nand UO_2371 (O_2371,N_18630,N_18644);
nand UO_2372 (O_2372,N_18062,N_18500);
and UO_2373 (O_2373,N_19134,N_19747);
nand UO_2374 (O_2374,N_19840,N_19170);
and UO_2375 (O_2375,N_18058,N_18388);
nand UO_2376 (O_2376,N_19305,N_18313);
and UO_2377 (O_2377,N_19828,N_18547);
nor UO_2378 (O_2378,N_19119,N_18149);
xnor UO_2379 (O_2379,N_18934,N_19439);
nand UO_2380 (O_2380,N_19717,N_19500);
nand UO_2381 (O_2381,N_18961,N_19823);
nor UO_2382 (O_2382,N_18084,N_19288);
or UO_2383 (O_2383,N_19044,N_18767);
nor UO_2384 (O_2384,N_18970,N_19028);
and UO_2385 (O_2385,N_18508,N_18150);
or UO_2386 (O_2386,N_18978,N_18184);
nor UO_2387 (O_2387,N_18502,N_19367);
nor UO_2388 (O_2388,N_19446,N_18117);
nor UO_2389 (O_2389,N_19438,N_19667);
xor UO_2390 (O_2390,N_19676,N_18249);
xnor UO_2391 (O_2391,N_18592,N_19233);
xnor UO_2392 (O_2392,N_18060,N_18475);
nand UO_2393 (O_2393,N_19283,N_19965);
nor UO_2394 (O_2394,N_18621,N_18872);
nand UO_2395 (O_2395,N_18222,N_19675);
nor UO_2396 (O_2396,N_18926,N_18616);
xnor UO_2397 (O_2397,N_18518,N_19455);
and UO_2398 (O_2398,N_19937,N_19922);
xor UO_2399 (O_2399,N_18941,N_18564);
nand UO_2400 (O_2400,N_18764,N_18738);
and UO_2401 (O_2401,N_18401,N_18885);
and UO_2402 (O_2402,N_18587,N_18263);
nand UO_2403 (O_2403,N_19731,N_19429);
and UO_2404 (O_2404,N_19160,N_19274);
xor UO_2405 (O_2405,N_18712,N_19573);
and UO_2406 (O_2406,N_18488,N_19900);
nor UO_2407 (O_2407,N_18049,N_18967);
or UO_2408 (O_2408,N_19789,N_18678);
nor UO_2409 (O_2409,N_19275,N_18852);
nor UO_2410 (O_2410,N_18961,N_19535);
xor UO_2411 (O_2411,N_18803,N_18059);
and UO_2412 (O_2412,N_18752,N_18882);
nand UO_2413 (O_2413,N_18769,N_18671);
xor UO_2414 (O_2414,N_19547,N_19037);
nor UO_2415 (O_2415,N_19939,N_19571);
nand UO_2416 (O_2416,N_18403,N_18480);
and UO_2417 (O_2417,N_18517,N_18351);
and UO_2418 (O_2418,N_18802,N_19799);
xnor UO_2419 (O_2419,N_18243,N_18188);
nand UO_2420 (O_2420,N_18662,N_19497);
nand UO_2421 (O_2421,N_19797,N_19072);
nand UO_2422 (O_2422,N_19825,N_18239);
or UO_2423 (O_2423,N_19871,N_18761);
or UO_2424 (O_2424,N_18177,N_18994);
nor UO_2425 (O_2425,N_18393,N_18206);
nand UO_2426 (O_2426,N_18504,N_19407);
nand UO_2427 (O_2427,N_19571,N_18273);
or UO_2428 (O_2428,N_18196,N_19210);
or UO_2429 (O_2429,N_18559,N_19532);
nor UO_2430 (O_2430,N_19788,N_19974);
xor UO_2431 (O_2431,N_19264,N_18606);
xnor UO_2432 (O_2432,N_19705,N_19691);
and UO_2433 (O_2433,N_19984,N_18680);
nand UO_2434 (O_2434,N_19476,N_19170);
and UO_2435 (O_2435,N_19020,N_19135);
xor UO_2436 (O_2436,N_19463,N_19550);
and UO_2437 (O_2437,N_19822,N_19954);
nand UO_2438 (O_2438,N_18194,N_18566);
and UO_2439 (O_2439,N_19170,N_19236);
and UO_2440 (O_2440,N_18060,N_19737);
or UO_2441 (O_2441,N_18559,N_18193);
or UO_2442 (O_2442,N_18757,N_18258);
or UO_2443 (O_2443,N_18298,N_18092);
or UO_2444 (O_2444,N_19032,N_19566);
nor UO_2445 (O_2445,N_19467,N_18525);
nand UO_2446 (O_2446,N_19343,N_19437);
nor UO_2447 (O_2447,N_19791,N_19755);
xnor UO_2448 (O_2448,N_18813,N_18649);
nand UO_2449 (O_2449,N_18321,N_19202);
and UO_2450 (O_2450,N_18582,N_19598);
nand UO_2451 (O_2451,N_19312,N_19878);
and UO_2452 (O_2452,N_18105,N_18428);
or UO_2453 (O_2453,N_18492,N_18767);
nor UO_2454 (O_2454,N_18874,N_19401);
xnor UO_2455 (O_2455,N_18519,N_18412);
nand UO_2456 (O_2456,N_19847,N_19347);
nand UO_2457 (O_2457,N_18092,N_19923);
or UO_2458 (O_2458,N_19501,N_19442);
nand UO_2459 (O_2459,N_19494,N_19367);
and UO_2460 (O_2460,N_19164,N_19818);
nand UO_2461 (O_2461,N_19764,N_18842);
xnor UO_2462 (O_2462,N_18362,N_19490);
nand UO_2463 (O_2463,N_18641,N_19549);
nor UO_2464 (O_2464,N_19955,N_19777);
xor UO_2465 (O_2465,N_18523,N_18261);
xnor UO_2466 (O_2466,N_19318,N_18779);
nor UO_2467 (O_2467,N_18127,N_19738);
xor UO_2468 (O_2468,N_18319,N_18658);
and UO_2469 (O_2469,N_18435,N_18924);
or UO_2470 (O_2470,N_19647,N_18675);
xor UO_2471 (O_2471,N_18853,N_19219);
nand UO_2472 (O_2472,N_18811,N_19923);
and UO_2473 (O_2473,N_19443,N_19349);
or UO_2474 (O_2474,N_19326,N_19056);
or UO_2475 (O_2475,N_19836,N_19060);
xnor UO_2476 (O_2476,N_18847,N_19129);
or UO_2477 (O_2477,N_19240,N_18714);
and UO_2478 (O_2478,N_19857,N_19024);
nor UO_2479 (O_2479,N_19703,N_18451);
and UO_2480 (O_2480,N_18207,N_18801);
xnor UO_2481 (O_2481,N_18088,N_19649);
nor UO_2482 (O_2482,N_18770,N_18622);
and UO_2483 (O_2483,N_19591,N_19476);
nor UO_2484 (O_2484,N_18916,N_19326);
xnor UO_2485 (O_2485,N_19295,N_19786);
and UO_2486 (O_2486,N_19098,N_19664);
nand UO_2487 (O_2487,N_19090,N_18663);
or UO_2488 (O_2488,N_19261,N_18548);
xnor UO_2489 (O_2489,N_19786,N_19757);
nand UO_2490 (O_2490,N_19987,N_18313);
nand UO_2491 (O_2491,N_18979,N_19978);
and UO_2492 (O_2492,N_19492,N_18442);
or UO_2493 (O_2493,N_19157,N_19652);
and UO_2494 (O_2494,N_18071,N_19472);
xnor UO_2495 (O_2495,N_19319,N_18658);
xnor UO_2496 (O_2496,N_19155,N_19691);
or UO_2497 (O_2497,N_18967,N_19903);
nor UO_2498 (O_2498,N_18175,N_18129);
nand UO_2499 (O_2499,N_19052,N_19796);
endmodule