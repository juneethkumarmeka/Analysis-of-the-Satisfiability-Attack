module basic_1000_10000_1500_4_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_433,In_796);
nand U1 (N_1,In_736,In_946);
nand U2 (N_2,In_636,In_704);
and U3 (N_3,In_598,In_128);
or U4 (N_4,In_981,In_2);
or U5 (N_5,In_336,In_57);
xor U6 (N_6,In_671,In_206);
nor U7 (N_7,In_640,In_919);
nor U8 (N_8,In_524,In_746);
or U9 (N_9,In_760,In_253);
or U10 (N_10,In_747,In_152);
nor U11 (N_11,In_278,In_858);
and U12 (N_12,In_205,In_562);
xnor U13 (N_13,In_609,In_254);
xnor U14 (N_14,In_276,In_975);
and U15 (N_15,In_291,In_550);
or U16 (N_16,In_395,In_717);
and U17 (N_17,In_862,In_322);
nor U18 (N_18,In_419,In_712);
xnor U19 (N_19,In_3,In_680);
nor U20 (N_20,In_134,In_413);
and U21 (N_21,In_612,In_602);
or U22 (N_22,In_860,In_664);
nand U23 (N_23,In_705,In_460);
nand U24 (N_24,In_214,In_93);
or U25 (N_25,In_149,In_71);
xor U26 (N_26,In_899,In_317);
nand U27 (N_27,In_258,In_864);
xor U28 (N_28,In_8,In_706);
and U29 (N_29,In_97,In_956);
nand U30 (N_30,In_196,In_654);
xor U31 (N_31,In_586,In_448);
nor U32 (N_32,In_262,In_283);
nor U33 (N_33,In_820,In_74);
xnor U34 (N_34,In_436,In_326);
xor U35 (N_35,In_473,In_721);
and U36 (N_36,In_937,In_776);
nor U37 (N_37,In_332,In_175);
xor U38 (N_38,In_881,In_492);
xor U39 (N_39,In_534,In_471);
nand U40 (N_40,In_571,In_288);
xor U41 (N_41,In_866,In_846);
and U42 (N_42,In_559,In_313);
or U43 (N_43,In_594,In_394);
or U44 (N_44,In_748,In_869);
nor U45 (N_45,In_201,In_236);
xnor U46 (N_46,In_857,In_979);
and U47 (N_47,In_915,In_430);
nor U48 (N_48,In_153,In_425);
xor U49 (N_49,In_268,In_588);
and U50 (N_50,In_592,In_882);
nor U51 (N_51,In_104,In_184);
nor U52 (N_52,In_303,In_852);
nand U53 (N_53,In_366,In_130);
nand U54 (N_54,In_845,In_661);
and U55 (N_55,In_749,In_652);
nor U56 (N_56,In_959,In_217);
and U57 (N_57,In_604,In_167);
xnor U58 (N_58,In_887,In_60);
xnor U59 (N_59,In_356,In_856);
nor U60 (N_60,In_733,In_825);
and U61 (N_61,In_989,In_369);
xnor U62 (N_62,In_78,In_150);
xor U63 (N_63,In_397,In_66);
and U64 (N_64,In_164,In_783);
nor U65 (N_65,In_926,In_169);
xnor U66 (N_66,In_650,In_812);
and U67 (N_67,In_391,In_916);
or U68 (N_68,In_470,In_466);
nor U69 (N_69,In_489,In_787);
or U70 (N_70,In_126,In_774);
or U71 (N_71,In_692,In_40);
or U72 (N_72,In_694,In_305);
nor U73 (N_73,In_822,In_483);
nand U74 (N_74,In_18,In_154);
nor U75 (N_75,In_73,In_280);
or U76 (N_76,In_50,In_665);
nor U77 (N_77,In_353,In_310);
and U78 (N_78,In_939,In_840);
xor U79 (N_79,In_215,In_96);
nand U80 (N_80,In_708,In_751);
or U81 (N_81,In_204,In_797);
and U82 (N_82,In_722,In_744);
nor U83 (N_83,In_940,In_584);
xnor U84 (N_84,In_848,In_182);
nor U85 (N_85,In_171,In_452);
or U86 (N_86,In_686,In_47);
nand U87 (N_87,In_597,In_298);
nor U88 (N_88,In_851,In_65);
nor U89 (N_89,In_284,In_16);
or U90 (N_90,In_231,In_372);
or U91 (N_91,In_993,In_77);
xor U92 (N_92,In_727,In_261);
and U93 (N_93,In_577,In_379);
nor U94 (N_94,In_750,In_75);
and U95 (N_95,In_859,In_933);
or U96 (N_96,In_244,In_509);
or U97 (N_97,In_403,In_438);
or U98 (N_98,In_443,In_222);
or U99 (N_99,In_341,In_789);
nor U100 (N_100,In_139,In_34);
nor U101 (N_101,In_606,In_980);
and U102 (N_102,In_177,In_872);
nor U103 (N_103,In_210,In_833);
nand U104 (N_104,In_685,In_417);
nand U105 (N_105,In_200,In_43);
and U106 (N_106,In_493,In_468);
and U107 (N_107,In_230,In_400);
nand U108 (N_108,In_663,In_761);
nand U109 (N_109,In_581,In_271);
or U110 (N_110,In_30,In_120);
nor U111 (N_111,In_319,In_823);
nand U112 (N_112,In_589,In_497);
nand U113 (N_113,In_107,In_447);
nand U114 (N_114,In_566,In_237);
or U115 (N_115,In_409,In_110);
nor U116 (N_116,In_199,In_181);
nor U117 (N_117,In_682,In_49);
nor U118 (N_118,In_243,In_905);
or U119 (N_119,In_526,In_451);
and U120 (N_120,In_131,In_977);
or U121 (N_121,In_800,In_501);
nor U122 (N_122,In_273,In_734);
nand U123 (N_123,In_963,In_404);
nand U124 (N_124,In_266,In_563);
xor U125 (N_125,In_985,In_819);
xnor U126 (N_126,In_969,In_224);
xnor U127 (N_127,In_672,In_143);
nor U128 (N_128,In_623,In_235);
or U129 (N_129,In_625,In_290);
or U130 (N_130,In_304,In_900);
xnor U131 (N_131,In_94,In_457);
or U132 (N_132,In_850,In_340);
xor U133 (N_133,In_595,In_921);
or U134 (N_134,In_945,In_407);
nor U135 (N_135,In_902,In_307);
nor U136 (N_136,In_402,In_221);
xnor U137 (N_137,In_488,In_920);
nor U138 (N_138,In_999,In_765);
or U139 (N_139,In_551,In_830);
xor U140 (N_140,In_903,In_913);
xor U141 (N_141,In_791,In_179);
and U142 (N_142,In_141,In_198);
nor U143 (N_143,In_351,In_745);
nor U144 (N_144,In_561,In_837);
xnor U145 (N_145,In_331,In_91);
nand U146 (N_146,In_620,In_114);
nor U147 (N_147,In_904,In_345);
and U148 (N_148,In_500,In_788);
xnor U149 (N_149,In_922,In_33);
xor U150 (N_150,In_737,In_659);
nor U151 (N_151,In_603,In_990);
or U152 (N_152,In_349,In_302);
nand U153 (N_153,In_378,In_113);
or U154 (N_154,In_778,In_189);
or U155 (N_155,In_677,In_1);
xor U156 (N_156,In_593,In_388);
and U157 (N_157,In_807,In_924);
nor U158 (N_158,In_260,In_781);
nand U159 (N_159,In_826,In_549);
xnor U160 (N_160,In_988,In_279);
and U161 (N_161,In_546,In_596);
nor U162 (N_162,In_365,In_14);
nor U163 (N_163,In_165,In_942);
nor U164 (N_164,In_277,In_129);
nor U165 (N_165,In_798,In_863);
or U166 (N_166,In_289,In_477);
nand U167 (N_167,In_896,In_875);
and U168 (N_168,In_622,In_491);
or U169 (N_169,In_821,In_764);
nor U170 (N_170,In_155,In_20);
and U171 (N_171,In_324,In_525);
nor U172 (N_172,In_811,In_888);
and U173 (N_173,In_907,In_478);
xnor U174 (N_174,In_930,In_576);
nor U175 (N_175,In_987,In_469);
and U176 (N_176,In_72,In_517);
and U177 (N_177,In_703,In_292);
nand U178 (N_178,In_445,In_295);
nand U179 (N_179,In_955,In_193);
nand U180 (N_180,In_118,In_618);
nor U181 (N_181,In_644,In_635);
and U182 (N_182,In_681,In_98);
and U183 (N_183,In_666,In_495);
or U184 (N_184,In_874,In_669);
nor U185 (N_185,In_886,In_670);
and U186 (N_186,In_906,In_255);
or U187 (N_187,In_232,In_754);
nor U188 (N_188,In_486,In_48);
nand U189 (N_189,In_720,In_518);
and U190 (N_190,In_505,In_371);
nand U191 (N_191,In_697,In_503);
nand U192 (N_192,In_446,In_84);
nor U193 (N_193,In_515,In_377);
and U194 (N_194,In_766,In_953);
xnor U195 (N_195,In_26,In_810);
nand U196 (N_196,In_772,In_813);
nor U197 (N_197,In_241,In_281);
and U198 (N_198,In_228,In_616);
or U199 (N_199,In_406,In_974);
nand U200 (N_200,In_743,In_502);
nor U201 (N_201,In_335,In_914);
xnor U202 (N_202,In_877,In_234);
or U203 (N_203,In_948,In_12);
nor U204 (N_204,In_27,In_983);
nor U205 (N_205,In_286,In_994);
nor U206 (N_206,In_180,In_867);
xnor U207 (N_207,In_601,In_827);
nor U208 (N_208,In_790,In_531);
nand U209 (N_209,In_490,In_358);
nor U210 (N_210,In_824,In_792);
and U211 (N_211,In_462,In_716);
and U212 (N_212,In_731,In_334);
nor U213 (N_213,In_893,In_381);
and U214 (N_214,In_192,In_111);
nor U215 (N_215,In_367,In_719);
nor U216 (N_216,In_641,In_54);
or U217 (N_217,In_634,In_116);
xor U218 (N_218,In_9,In_678);
xnor U219 (N_219,In_738,In_318);
or U220 (N_220,In_373,In_632);
nand U221 (N_221,In_984,In_769);
and U222 (N_222,In_709,In_106);
nor U223 (N_223,In_53,In_730);
nor U224 (N_224,In_39,In_7);
xnor U225 (N_225,In_784,In_207);
and U226 (N_226,In_775,In_567);
or U227 (N_227,In_572,In_718);
nand U228 (N_228,In_212,In_952);
or U229 (N_229,In_385,In_412);
and U230 (N_230,In_793,In_173);
xor U231 (N_231,In_21,In_272);
and U232 (N_232,In_465,In_961);
xor U233 (N_233,In_570,In_300);
or U234 (N_234,In_516,In_138);
nand U235 (N_235,In_814,In_533);
and U236 (N_236,In_883,In_578);
and U237 (N_237,In_575,In_558);
nor U238 (N_238,In_957,In_506);
and U239 (N_239,In_964,In_350);
and U240 (N_240,In_607,In_732);
or U241 (N_241,In_679,In_31);
nand U242 (N_242,In_947,In_756);
or U243 (N_243,In_450,In_855);
nor U244 (N_244,In_480,In_456);
or U245 (N_245,In_917,In_803);
xnor U246 (N_246,In_287,In_995);
xor U247 (N_247,In_777,In_347);
xor U248 (N_248,In_252,In_203);
and U249 (N_249,In_176,In_475);
nand U250 (N_250,In_815,In_619);
nor U251 (N_251,In_537,In_755);
or U252 (N_252,In_355,In_337);
nor U253 (N_253,In_528,In_418);
xor U254 (N_254,In_660,In_630);
and U255 (N_255,In_115,In_285);
nor U256 (N_256,In_364,In_250);
nor U257 (N_257,In_527,In_901);
nand U258 (N_258,In_529,In_521);
nand U259 (N_259,In_504,In_123);
nor U260 (N_260,In_168,In_170);
nor U261 (N_261,In_695,In_144);
xor U262 (N_262,In_376,In_297);
nor U263 (N_263,In_614,In_808);
or U264 (N_264,In_474,In_758);
xor U265 (N_265,In_380,In_631);
nand U266 (N_266,In_973,In_323);
nand U267 (N_267,In_548,In_954);
xnor U268 (N_268,In_163,In_918);
nor U269 (N_269,In_656,In_414);
xor U270 (N_270,In_218,In_794);
xnor U271 (N_271,In_348,In_458);
xor U272 (N_272,In_649,In_838);
or U273 (N_273,In_795,In_80);
nand U274 (N_274,In_997,In_628);
nand U275 (N_275,In_454,In_895);
or U276 (N_276,In_172,In_729);
or U277 (N_277,In_941,In_156);
nand U278 (N_278,In_146,In_109);
nand U279 (N_279,In_613,In_615);
nand U280 (N_280,In_352,In_481);
or U281 (N_281,In_38,In_841);
xnor U282 (N_282,In_223,In_482);
nor U283 (N_283,In_99,In_370);
nand U284 (N_284,In_740,In_725);
nor U285 (N_285,In_299,In_839);
or U286 (N_286,In_10,In_421);
or U287 (N_287,In_361,In_159);
xor U288 (N_288,In_61,In_455);
nor U289 (N_289,In_836,In_362);
nand U290 (N_290,In_148,In_157);
nand U291 (N_291,In_927,In_583);
nand U292 (N_292,In_90,In_849);
xor U293 (N_293,In_621,In_701);
nor U294 (N_294,In_105,In_690);
xor U295 (N_295,In_333,In_684);
xor U296 (N_296,In_197,In_870);
and U297 (N_297,In_962,In_103);
nor U298 (N_298,In_780,In_763);
and U299 (N_299,In_910,In_127);
nor U300 (N_300,In_158,In_805);
or U301 (N_301,In_876,In_508);
xor U302 (N_302,In_880,In_354);
xnor U303 (N_303,In_809,In_411);
xor U304 (N_304,In_11,In_687);
and U305 (N_305,In_81,In_225);
or U306 (N_306,In_965,In_715);
or U307 (N_307,In_64,In_426);
or U308 (N_308,In_368,In_676);
xnor U309 (N_309,In_294,In_599);
and U310 (N_310,In_359,In_832);
xnor U311 (N_311,In_847,In_311);
xor U312 (N_312,In_911,In_467);
nand U313 (N_313,In_321,In_142);
or U314 (N_314,In_41,In_239);
and U315 (N_315,In_100,In_536);
nor U316 (N_316,In_427,In_339);
nor U317 (N_317,In_655,In_560);
nor U318 (N_318,In_771,In_208);
or U319 (N_319,In_306,In_547);
nor U320 (N_320,In_202,In_938);
and U321 (N_321,In_651,In_137);
xor U322 (N_322,In_293,In_667);
and U323 (N_323,In_909,In_82);
and U324 (N_324,In_86,In_982);
nand U325 (N_325,In_25,In_498);
nand U326 (N_326,In_522,In_520);
nand U327 (N_327,In_88,In_42);
nor U328 (N_328,In_187,In_935);
nor U329 (N_329,In_161,In_608);
nor U330 (N_330,In_555,In_693);
or U331 (N_331,In_429,In_889);
or U332 (N_332,In_892,In_108);
nand U333 (N_333,In_390,In_532);
and U334 (N_334,In_929,In_69);
and U335 (N_335,In_868,In_986);
nand U336 (N_336,In_79,In_514);
xor U337 (N_337,In_779,In_831);
nand U338 (N_338,In_770,In_768);
nor U339 (N_339,In_101,In_136);
nand U340 (N_340,In_133,In_934);
nor U341 (N_341,In_375,In_437);
and U342 (N_342,In_219,In_316);
nor U343 (N_343,In_691,In_140);
nor U344 (N_344,In_801,In_617);
xnor U345 (N_345,In_431,In_587);
nand U346 (N_346,In_246,In_828);
or U347 (N_347,In_398,In_22);
nand U348 (N_348,In_854,In_314);
xnor U349 (N_349,In_15,In_461);
nand U350 (N_350,In_393,In_925);
xor U351 (N_351,In_541,In_55);
nand U352 (N_352,In_966,In_162);
xnor U353 (N_353,In_552,In_63);
or U354 (N_354,In_56,In_256);
xnor U355 (N_355,In_23,In_209);
nor U356 (N_356,In_229,In_569);
xor U357 (N_357,In_389,In_117);
and U358 (N_358,In_648,In_423);
xnor U359 (N_359,In_83,In_519);
or U360 (N_360,In_330,In_696);
nor U361 (N_361,In_68,In_683);
or U362 (N_362,In_259,In_211);
xor U363 (N_363,In_873,In_726);
nor U364 (N_364,In_753,In_275);
and U365 (N_365,In_978,In_36);
nand U366 (N_366,In_512,In_996);
nor U367 (N_367,In_976,In_752);
xnor U368 (N_368,In_463,In_865);
xor U369 (N_369,In_565,In_543);
xor U370 (N_370,In_713,In_51);
or U371 (N_371,In_19,In_132);
xor U372 (N_372,In_487,In_574);
and U373 (N_373,In_13,In_89);
nor U374 (N_374,In_0,In_674);
nor U375 (N_375,In_992,In_714);
nand U376 (N_376,In_439,In_220);
and U377 (N_377,In_6,In_328);
or U378 (N_378,In_639,In_600);
and U379 (N_379,In_950,In_428);
and U380 (N_380,In_401,In_943);
or U381 (N_381,In_325,In_923);
or U382 (N_382,In_611,In_52);
or U383 (N_383,In_102,In_653);
or U384 (N_384,In_309,In_449);
nand U385 (N_385,In_759,In_513);
xor U386 (N_386,In_844,In_884);
and U387 (N_387,In_556,In_44);
xor U388 (N_388,In_269,In_245);
and U389 (N_389,In_637,In_76);
nor U390 (N_390,In_786,In_879);
and U391 (N_391,In_638,In_829);
nand U392 (N_392,In_257,In_195);
nand U393 (N_393,In_312,In_32);
nand U394 (N_394,In_122,In_424);
nor U395 (N_395,In_545,In_972);
or U396 (N_396,In_186,In_124);
xnor U397 (N_397,In_960,In_530);
and U398 (N_398,In_35,In_384);
nand U399 (N_399,In_135,In_878);
or U400 (N_400,In_415,In_346);
nand U401 (N_401,In_247,In_700);
and U402 (N_402,In_580,In_668);
nand U403 (N_403,In_435,In_37);
or U404 (N_404,In_785,In_70);
nor U405 (N_405,In_591,In_213);
xnor U406 (N_406,In_951,In_5);
or U407 (N_407,In_647,In_166);
nand U408 (N_408,In_605,In_485);
nand U409 (N_409,In_510,In_185);
and U410 (N_410,In_707,In_741);
nand U411 (N_411,In_523,In_958);
and U412 (N_412,In_908,In_890);
or U413 (N_413,In_739,In_399);
nor U414 (N_414,In_762,In_564);
or U415 (N_415,In_496,In_835);
and U416 (N_416,In_912,In_773);
xnor U417 (N_417,In_579,In_440);
nor U418 (N_418,In_688,In_542);
or U419 (N_419,In_274,In_183);
or U420 (N_420,In_804,In_263);
nand U421 (N_421,In_121,In_264);
and U422 (N_422,In_344,In_675);
nor U423 (N_423,In_343,In_626);
nand U424 (N_424,In_711,In_382);
nor U425 (N_425,In_296,In_420);
or U426 (N_426,In_327,In_301);
or U427 (N_427,In_698,In_885);
xnor U428 (N_428,In_629,In_194);
and U429 (N_429,In_642,In_834);
nand U430 (N_430,In_897,In_802);
or U431 (N_431,In_816,In_444);
or U432 (N_432,In_432,In_573);
or U433 (N_433,In_405,In_342);
xor U434 (N_434,In_610,In_843);
or U435 (N_435,In_174,In_442);
nand U436 (N_436,In_932,In_112);
and U437 (N_437,In_357,In_544);
nand U438 (N_438,In_119,In_95);
or U439 (N_439,In_898,In_396);
or U440 (N_440,In_871,In_568);
nand U441 (N_441,In_476,In_125);
or U442 (N_442,In_282,In_383);
or U443 (N_443,In_817,In_87);
or U444 (N_444,In_633,In_484);
or U445 (N_445,In_338,In_28);
xor U446 (N_446,In_853,In_242);
or U447 (N_447,In_227,In_17);
xnor U448 (N_448,In_416,In_387);
or U449 (N_449,In_710,In_147);
nor U450 (N_450,In_861,In_85);
or U451 (N_451,In_360,In_818);
and U452 (N_452,In_29,In_67);
nor U453 (N_453,In_511,In_329);
nor U454 (N_454,In_645,In_58);
or U455 (N_455,In_459,In_658);
xor U456 (N_456,In_251,In_441);
and U457 (N_457,In_657,In_782);
nor U458 (N_458,In_970,In_735);
and U459 (N_459,In_553,In_554);
nor U460 (N_460,In_240,In_265);
or U461 (N_461,In_968,In_151);
nor U462 (N_462,In_190,In_410);
or U463 (N_463,In_724,In_540);
nor U464 (N_464,In_62,In_624);
nand U465 (N_465,In_538,In_160);
nor U466 (N_466,In_742,In_931);
xor U467 (N_467,In_464,In_267);
nand U468 (N_468,In_585,In_891);
nand U469 (N_469,In_24,In_757);
and U470 (N_470,In_582,In_971);
nor U471 (N_471,In_46,In_949);
and U472 (N_472,In_689,In_453);
and U473 (N_473,In_472,In_216);
and U474 (N_474,In_178,In_191);
or U475 (N_475,In_627,In_673);
xor U476 (N_476,In_842,In_45);
and U477 (N_477,In_308,In_320);
nor U478 (N_478,In_557,In_643);
nand U479 (N_479,In_392,In_894);
nand U480 (N_480,In_315,In_4);
or U481 (N_481,In_646,In_233);
xor U482 (N_482,In_507,In_238);
xor U483 (N_483,In_767,In_494);
nand U484 (N_484,In_434,In_145);
nand U485 (N_485,In_499,In_728);
and U486 (N_486,In_363,In_998);
or U487 (N_487,In_479,In_799);
or U488 (N_488,In_967,In_535);
nor U489 (N_489,In_408,In_944);
or U490 (N_490,In_806,In_699);
nor U491 (N_491,In_386,In_991);
nand U492 (N_492,In_188,In_936);
and U493 (N_493,In_59,In_723);
or U494 (N_494,In_270,In_590);
and U495 (N_495,In_248,In_702);
nor U496 (N_496,In_374,In_226);
xor U497 (N_497,In_249,In_928);
or U498 (N_498,In_662,In_422);
xor U499 (N_499,In_92,In_539);
xor U500 (N_500,In_645,In_661);
nand U501 (N_501,In_78,In_147);
nor U502 (N_502,In_447,In_682);
or U503 (N_503,In_661,In_777);
nand U504 (N_504,In_283,In_331);
nand U505 (N_505,In_694,In_890);
xor U506 (N_506,In_281,In_936);
xor U507 (N_507,In_158,In_217);
nor U508 (N_508,In_200,In_600);
nand U509 (N_509,In_230,In_333);
xnor U510 (N_510,In_386,In_402);
xor U511 (N_511,In_784,In_930);
and U512 (N_512,In_796,In_276);
or U513 (N_513,In_546,In_793);
nand U514 (N_514,In_817,In_642);
nand U515 (N_515,In_171,In_184);
nand U516 (N_516,In_37,In_319);
nor U517 (N_517,In_676,In_975);
xor U518 (N_518,In_34,In_47);
xor U519 (N_519,In_962,In_171);
nor U520 (N_520,In_322,In_549);
and U521 (N_521,In_547,In_264);
or U522 (N_522,In_442,In_969);
or U523 (N_523,In_436,In_716);
nand U524 (N_524,In_535,In_684);
nor U525 (N_525,In_792,In_694);
nand U526 (N_526,In_201,In_553);
nor U527 (N_527,In_542,In_286);
or U528 (N_528,In_917,In_28);
nor U529 (N_529,In_970,In_825);
nor U530 (N_530,In_299,In_532);
or U531 (N_531,In_266,In_782);
xnor U532 (N_532,In_469,In_422);
xor U533 (N_533,In_335,In_593);
nor U534 (N_534,In_139,In_725);
nand U535 (N_535,In_511,In_891);
or U536 (N_536,In_481,In_4);
xnor U537 (N_537,In_138,In_132);
nor U538 (N_538,In_120,In_294);
or U539 (N_539,In_616,In_930);
and U540 (N_540,In_268,In_230);
or U541 (N_541,In_894,In_887);
or U542 (N_542,In_654,In_630);
or U543 (N_543,In_94,In_86);
or U544 (N_544,In_218,In_541);
xnor U545 (N_545,In_406,In_221);
nor U546 (N_546,In_188,In_959);
and U547 (N_547,In_287,In_527);
nand U548 (N_548,In_721,In_98);
and U549 (N_549,In_755,In_234);
nor U550 (N_550,In_244,In_872);
nor U551 (N_551,In_591,In_869);
and U552 (N_552,In_579,In_244);
or U553 (N_553,In_168,In_702);
or U554 (N_554,In_151,In_872);
nor U555 (N_555,In_552,In_750);
and U556 (N_556,In_940,In_327);
nor U557 (N_557,In_841,In_44);
nand U558 (N_558,In_174,In_702);
or U559 (N_559,In_501,In_625);
nor U560 (N_560,In_757,In_290);
or U561 (N_561,In_728,In_337);
or U562 (N_562,In_90,In_135);
nor U563 (N_563,In_919,In_262);
nor U564 (N_564,In_917,In_887);
xnor U565 (N_565,In_614,In_296);
and U566 (N_566,In_973,In_991);
or U567 (N_567,In_298,In_576);
xor U568 (N_568,In_671,In_52);
or U569 (N_569,In_981,In_769);
nand U570 (N_570,In_157,In_100);
xor U571 (N_571,In_122,In_390);
or U572 (N_572,In_900,In_769);
and U573 (N_573,In_697,In_858);
xnor U574 (N_574,In_354,In_882);
xor U575 (N_575,In_839,In_550);
or U576 (N_576,In_441,In_27);
nor U577 (N_577,In_2,In_395);
nor U578 (N_578,In_474,In_13);
xnor U579 (N_579,In_920,In_837);
xnor U580 (N_580,In_476,In_691);
and U581 (N_581,In_681,In_677);
nand U582 (N_582,In_320,In_468);
or U583 (N_583,In_655,In_125);
and U584 (N_584,In_389,In_824);
nand U585 (N_585,In_581,In_526);
or U586 (N_586,In_106,In_677);
nor U587 (N_587,In_549,In_747);
and U588 (N_588,In_418,In_500);
xnor U589 (N_589,In_861,In_908);
xnor U590 (N_590,In_523,In_969);
and U591 (N_591,In_98,In_880);
and U592 (N_592,In_167,In_945);
or U593 (N_593,In_342,In_999);
and U594 (N_594,In_412,In_354);
and U595 (N_595,In_726,In_25);
nand U596 (N_596,In_98,In_727);
nand U597 (N_597,In_384,In_9);
nand U598 (N_598,In_759,In_449);
and U599 (N_599,In_660,In_184);
xnor U600 (N_600,In_863,In_618);
or U601 (N_601,In_887,In_936);
or U602 (N_602,In_558,In_827);
nand U603 (N_603,In_37,In_890);
nand U604 (N_604,In_823,In_216);
nor U605 (N_605,In_905,In_646);
xnor U606 (N_606,In_941,In_693);
xnor U607 (N_607,In_260,In_852);
or U608 (N_608,In_534,In_792);
xnor U609 (N_609,In_107,In_403);
nand U610 (N_610,In_74,In_850);
nor U611 (N_611,In_865,In_534);
or U612 (N_612,In_395,In_992);
or U613 (N_613,In_756,In_732);
nor U614 (N_614,In_518,In_243);
nand U615 (N_615,In_202,In_299);
nor U616 (N_616,In_550,In_790);
nor U617 (N_617,In_896,In_532);
or U618 (N_618,In_407,In_384);
xor U619 (N_619,In_20,In_109);
or U620 (N_620,In_919,In_141);
or U621 (N_621,In_335,In_766);
nor U622 (N_622,In_676,In_429);
nor U623 (N_623,In_145,In_429);
nand U624 (N_624,In_47,In_510);
xnor U625 (N_625,In_131,In_659);
nor U626 (N_626,In_33,In_358);
xor U627 (N_627,In_463,In_897);
and U628 (N_628,In_481,In_580);
nor U629 (N_629,In_931,In_800);
and U630 (N_630,In_737,In_53);
nor U631 (N_631,In_421,In_643);
nand U632 (N_632,In_971,In_70);
or U633 (N_633,In_171,In_881);
and U634 (N_634,In_101,In_924);
nand U635 (N_635,In_70,In_57);
nor U636 (N_636,In_134,In_660);
or U637 (N_637,In_744,In_633);
or U638 (N_638,In_943,In_1);
and U639 (N_639,In_994,In_104);
nor U640 (N_640,In_393,In_973);
nor U641 (N_641,In_464,In_146);
nand U642 (N_642,In_862,In_350);
or U643 (N_643,In_41,In_295);
nor U644 (N_644,In_840,In_332);
nand U645 (N_645,In_776,In_69);
and U646 (N_646,In_578,In_104);
xnor U647 (N_647,In_134,In_968);
and U648 (N_648,In_916,In_29);
xnor U649 (N_649,In_190,In_89);
nor U650 (N_650,In_442,In_484);
and U651 (N_651,In_843,In_836);
xor U652 (N_652,In_953,In_410);
xor U653 (N_653,In_725,In_417);
or U654 (N_654,In_793,In_554);
nand U655 (N_655,In_483,In_90);
xor U656 (N_656,In_288,In_193);
nand U657 (N_657,In_167,In_942);
nand U658 (N_658,In_996,In_818);
xnor U659 (N_659,In_179,In_275);
xor U660 (N_660,In_238,In_608);
nor U661 (N_661,In_405,In_83);
or U662 (N_662,In_98,In_904);
nand U663 (N_663,In_193,In_357);
or U664 (N_664,In_574,In_61);
nand U665 (N_665,In_874,In_390);
nor U666 (N_666,In_544,In_902);
xnor U667 (N_667,In_784,In_630);
xor U668 (N_668,In_907,In_694);
nor U669 (N_669,In_656,In_583);
nor U670 (N_670,In_720,In_366);
nor U671 (N_671,In_631,In_466);
and U672 (N_672,In_678,In_247);
nand U673 (N_673,In_560,In_553);
nor U674 (N_674,In_192,In_296);
or U675 (N_675,In_192,In_397);
or U676 (N_676,In_845,In_400);
nand U677 (N_677,In_922,In_464);
xor U678 (N_678,In_604,In_720);
nor U679 (N_679,In_574,In_519);
and U680 (N_680,In_617,In_755);
xnor U681 (N_681,In_676,In_729);
xnor U682 (N_682,In_863,In_924);
xnor U683 (N_683,In_522,In_578);
nand U684 (N_684,In_915,In_264);
and U685 (N_685,In_375,In_940);
nor U686 (N_686,In_711,In_648);
nor U687 (N_687,In_9,In_3);
or U688 (N_688,In_725,In_910);
and U689 (N_689,In_949,In_423);
xnor U690 (N_690,In_424,In_358);
nand U691 (N_691,In_557,In_998);
and U692 (N_692,In_939,In_353);
xor U693 (N_693,In_880,In_722);
nor U694 (N_694,In_426,In_998);
and U695 (N_695,In_709,In_93);
nor U696 (N_696,In_84,In_777);
nor U697 (N_697,In_403,In_991);
nand U698 (N_698,In_733,In_890);
nor U699 (N_699,In_941,In_912);
and U700 (N_700,In_520,In_789);
xor U701 (N_701,In_285,In_286);
or U702 (N_702,In_700,In_690);
nor U703 (N_703,In_325,In_629);
nor U704 (N_704,In_196,In_947);
or U705 (N_705,In_233,In_190);
and U706 (N_706,In_530,In_848);
nand U707 (N_707,In_148,In_304);
and U708 (N_708,In_40,In_712);
or U709 (N_709,In_402,In_446);
and U710 (N_710,In_305,In_954);
and U711 (N_711,In_656,In_936);
nor U712 (N_712,In_722,In_193);
nor U713 (N_713,In_942,In_80);
nand U714 (N_714,In_792,In_983);
nor U715 (N_715,In_747,In_111);
nand U716 (N_716,In_997,In_31);
nand U717 (N_717,In_908,In_610);
xnor U718 (N_718,In_923,In_608);
nor U719 (N_719,In_385,In_723);
nand U720 (N_720,In_101,In_528);
nor U721 (N_721,In_8,In_810);
and U722 (N_722,In_171,In_675);
nand U723 (N_723,In_222,In_571);
nor U724 (N_724,In_710,In_806);
or U725 (N_725,In_318,In_430);
nand U726 (N_726,In_679,In_734);
xor U727 (N_727,In_134,In_837);
and U728 (N_728,In_986,In_125);
nand U729 (N_729,In_589,In_933);
nand U730 (N_730,In_880,In_292);
nand U731 (N_731,In_71,In_804);
nor U732 (N_732,In_482,In_914);
nand U733 (N_733,In_606,In_948);
xor U734 (N_734,In_788,In_957);
xnor U735 (N_735,In_51,In_540);
or U736 (N_736,In_380,In_591);
nor U737 (N_737,In_170,In_137);
or U738 (N_738,In_736,In_565);
and U739 (N_739,In_913,In_667);
xnor U740 (N_740,In_545,In_952);
and U741 (N_741,In_240,In_332);
xor U742 (N_742,In_706,In_857);
xnor U743 (N_743,In_145,In_566);
nor U744 (N_744,In_941,In_473);
nand U745 (N_745,In_835,In_284);
or U746 (N_746,In_890,In_923);
and U747 (N_747,In_223,In_50);
xnor U748 (N_748,In_844,In_24);
or U749 (N_749,In_666,In_659);
nand U750 (N_750,In_124,In_704);
xnor U751 (N_751,In_860,In_347);
nor U752 (N_752,In_426,In_723);
nand U753 (N_753,In_645,In_600);
and U754 (N_754,In_499,In_826);
nand U755 (N_755,In_970,In_208);
xnor U756 (N_756,In_630,In_378);
or U757 (N_757,In_229,In_207);
and U758 (N_758,In_143,In_53);
and U759 (N_759,In_284,In_184);
nand U760 (N_760,In_154,In_638);
xnor U761 (N_761,In_567,In_873);
nor U762 (N_762,In_24,In_425);
or U763 (N_763,In_819,In_112);
nor U764 (N_764,In_73,In_805);
nor U765 (N_765,In_453,In_230);
nor U766 (N_766,In_993,In_336);
or U767 (N_767,In_448,In_813);
and U768 (N_768,In_619,In_408);
xnor U769 (N_769,In_676,In_339);
or U770 (N_770,In_213,In_419);
or U771 (N_771,In_282,In_292);
nand U772 (N_772,In_410,In_623);
nor U773 (N_773,In_982,In_967);
nand U774 (N_774,In_0,In_818);
or U775 (N_775,In_126,In_703);
nor U776 (N_776,In_2,In_159);
and U777 (N_777,In_826,In_725);
or U778 (N_778,In_935,In_481);
xor U779 (N_779,In_98,In_39);
xor U780 (N_780,In_582,In_383);
and U781 (N_781,In_417,In_572);
or U782 (N_782,In_166,In_285);
xor U783 (N_783,In_874,In_72);
nand U784 (N_784,In_478,In_376);
or U785 (N_785,In_288,In_940);
or U786 (N_786,In_601,In_844);
and U787 (N_787,In_452,In_640);
nor U788 (N_788,In_930,In_349);
xnor U789 (N_789,In_575,In_702);
xor U790 (N_790,In_510,In_791);
xor U791 (N_791,In_936,In_184);
xnor U792 (N_792,In_576,In_842);
xor U793 (N_793,In_438,In_949);
and U794 (N_794,In_933,In_168);
or U795 (N_795,In_571,In_335);
xor U796 (N_796,In_156,In_844);
and U797 (N_797,In_792,In_12);
nand U798 (N_798,In_479,In_705);
nor U799 (N_799,In_550,In_439);
xnor U800 (N_800,In_749,In_268);
nand U801 (N_801,In_150,In_481);
nand U802 (N_802,In_327,In_600);
or U803 (N_803,In_483,In_240);
or U804 (N_804,In_613,In_290);
and U805 (N_805,In_201,In_153);
nand U806 (N_806,In_126,In_337);
xnor U807 (N_807,In_203,In_829);
and U808 (N_808,In_449,In_957);
nand U809 (N_809,In_571,In_354);
and U810 (N_810,In_619,In_242);
xor U811 (N_811,In_440,In_797);
nand U812 (N_812,In_182,In_582);
and U813 (N_813,In_466,In_663);
nand U814 (N_814,In_563,In_180);
xor U815 (N_815,In_491,In_933);
xor U816 (N_816,In_579,In_668);
nand U817 (N_817,In_10,In_795);
nand U818 (N_818,In_17,In_313);
xor U819 (N_819,In_884,In_857);
nor U820 (N_820,In_23,In_47);
nand U821 (N_821,In_584,In_494);
nand U822 (N_822,In_725,In_845);
nor U823 (N_823,In_722,In_924);
and U824 (N_824,In_763,In_448);
nor U825 (N_825,In_991,In_181);
or U826 (N_826,In_805,In_545);
xnor U827 (N_827,In_508,In_919);
and U828 (N_828,In_177,In_991);
nor U829 (N_829,In_691,In_83);
and U830 (N_830,In_862,In_115);
or U831 (N_831,In_37,In_690);
nor U832 (N_832,In_613,In_677);
or U833 (N_833,In_735,In_942);
and U834 (N_834,In_44,In_493);
nor U835 (N_835,In_685,In_415);
nor U836 (N_836,In_60,In_701);
xor U837 (N_837,In_876,In_479);
nand U838 (N_838,In_991,In_180);
nor U839 (N_839,In_473,In_79);
nor U840 (N_840,In_137,In_127);
nand U841 (N_841,In_815,In_271);
xnor U842 (N_842,In_564,In_785);
or U843 (N_843,In_975,In_454);
nor U844 (N_844,In_129,In_502);
nand U845 (N_845,In_174,In_846);
and U846 (N_846,In_184,In_988);
nand U847 (N_847,In_14,In_478);
nand U848 (N_848,In_95,In_797);
nand U849 (N_849,In_92,In_452);
xor U850 (N_850,In_364,In_971);
and U851 (N_851,In_176,In_792);
nand U852 (N_852,In_949,In_242);
nand U853 (N_853,In_676,In_590);
xnor U854 (N_854,In_510,In_918);
or U855 (N_855,In_964,In_494);
nand U856 (N_856,In_185,In_938);
nand U857 (N_857,In_603,In_872);
or U858 (N_858,In_119,In_548);
or U859 (N_859,In_766,In_205);
nand U860 (N_860,In_138,In_39);
or U861 (N_861,In_452,In_571);
nand U862 (N_862,In_56,In_579);
xnor U863 (N_863,In_991,In_55);
nand U864 (N_864,In_802,In_54);
and U865 (N_865,In_777,In_154);
nand U866 (N_866,In_36,In_170);
nand U867 (N_867,In_541,In_324);
or U868 (N_868,In_321,In_472);
and U869 (N_869,In_373,In_272);
xor U870 (N_870,In_698,In_633);
xor U871 (N_871,In_701,In_740);
or U872 (N_872,In_39,In_510);
nand U873 (N_873,In_202,In_847);
nand U874 (N_874,In_221,In_675);
nor U875 (N_875,In_324,In_946);
or U876 (N_876,In_480,In_805);
nor U877 (N_877,In_456,In_878);
nand U878 (N_878,In_654,In_311);
xnor U879 (N_879,In_346,In_39);
nor U880 (N_880,In_647,In_985);
xnor U881 (N_881,In_345,In_50);
xnor U882 (N_882,In_240,In_364);
and U883 (N_883,In_320,In_521);
xnor U884 (N_884,In_523,In_455);
nand U885 (N_885,In_858,In_725);
or U886 (N_886,In_777,In_961);
nand U887 (N_887,In_636,In_770);
nor U888 (N_888,In_883,In_179);
or U889 (N_889,In_305,In_105);
nand U890 (N_890,In_829,In_814);
nor U891 (N_891,In_785,In_530);
nand U892 (N_892,In_298,In_672);
and U893 (N_893,In_127,In_567);
and U894 (N_894,In_307,In_54);
and U895 (N_895,In_177,In_491);
nor U896 (N_896,In_640,In_417);
nor U897 (N_897,In_232,In_912);
xnor U898 (N_898,In_463,In_689);
xor U899 (N_899,In_164,In_473);
and U900 (N_900,In_194,In_942);
or U901 (N_901,In_219,In_905);
nor U902 (N_902,In_446,In_610);
nand U903 (N_903,In_867,In_690);
xor U904 (N_904,In_749,In_404);
or U905 (N_905,In_469,In_214);
nand U906 (N_906,In_587,In_558);
nor U907 (N_907,In_413,In_853);
xnor U908 (N_908,In_457,In_932);
and U909 (N_909,In_193,In_20);
and U910 (N_910,In_986,In_739);
xor U911 (N_911,In_332,In_543);
nor U912 (N_912,In_686,In_434);
nand U913 (N_913,In_227,In_83);
xnor U914 (N_914,In_210,In_628);
and U915 (N_915,In_215,In_815);
xor U916 (N_916,In_287,In_176);
nand U917 (N_917,In_435,In_323);
or U918 (N_918,In_700,In_912);
or U919 (N_919,In_360,In_872);
xor U920 (N_920,In_615,In_429);
and U921 (N_921,In_829,In_437);
xnor U922 (N_922,In_824,In_780);
and U923 (N_923,In_246,In_336);
nor U924 (N_924,In_916,In_241);
nor U925 (N_925,In_588,In_755);
nor U926 (N_926,In_195,In_624);
or U927 (N_927,In_368,In_54);
xor U928 (N_928,In_939,In_309);
nor U929 (N_929,In_226,In_581);
xnor U930 (N_930,In_215,In_930);
nand U931 (N_931,In_679,In_795);
and U932 (N_932,In_412,In_750);
xnor U933 (N_933,In_653,In_758);
nand U934 (N_934,In_353,In_648);
and U935 (N_935,In_182,In_737);
nand U936 (N_936,In_520,In_435);
xnor U937 (N_937,In_748,In_680);
xnor U938 (N_938,In_306,In_680);
nand U939 (N_939,In_601,In_486);
nor U940 (N_940,In_348,In_431);
and U941 (N_941,In_688,In_196);
nor U942 (N_942,In_174,In_626);
nand U943 (N_943,In_170,In_660);
and U944 (N_944,In_638,In_883);
xor U945 (N_945,In_765,In_197);
nand U946 (N_946,In_29,In_876);
and U947 (N_947,In_970,In_913);
nor U948 (N_948,In_230,In_961);
or U949 (N_949,In_847,In_822);
or U950 (N_950,In_570,In_509);
nand U951 (N_951,In_351,In_936);
nand U952 (N_952,In_898,In_623);
or U953 (N_953,In_206,In_819);
nand U954 (N_954,In_21,In_409);
xor U955 (N_955,In_671,In_656);
xnor U956 (N_956,In_650,In_182);
or U957 (N_957,In_484,In_16);
or U958 (N_958,In_392,In_78);
nor U959 (N_959,In_430,In_653);
xor U960 (N_960,In_995,In_699);
and U961 (N_961,In_503,In_154);
nor U962 (N_962,In_321,In_948);
nand U963 (N_963,In_647,In_7);
xor U964 (N_964,In_404,In_488);
xor U965 (N_965,In_413,In_593);
nand U966 (N_966,In_430,In_557);
or U967 (N_967,In_567,In_387);
nor U968 (N_968,In_955,In_37);
xnor U969 (N_969,In_256,In_235);
or U970 (N_970,In_997,In_737);
nand U971 (N_971,In_828,In_3);
and U972 (N_972,In_367,In_674);
xor U973 (N_973,In_753,In_879);
nand U974 (N_974,In_199,In_540);
nand U975 (N_975,In_462,In_379);
or U976 (N_976,In_329,In_870);
xor U977 (N_977,In_634,In_862);
and U978 (N_978,In_780,In_380);
or U979 (N_979,In_365,In_977);
and U980 (N_980,In_218,In_260);
xnor U981 (N_981,In_12,In_557);
or U982 (N_982,In_235,In_570);
or U983 (N_983,In_839,In_110);
or U984 (N_984,In_127,In_546);
and U985 (N_985,In_451,In_21);
and U986 (N_986,In_664,In_286);
nor U987 (N_987,In_510,In_706);
xnor U988 (N_988,In_47,In_821);
or U989 (N_989,In_380,In_276);
and U990 (N_990,In_21,In_335);
nor U991 (N_991,In_54,In_322);
nand U992 (N_992,In_129,In_39);
or U993 (N_993,In_699,In_690);
and U994 (N_994,In_266,In_64);
and U995 (N_995,In_932,In_885);
and U996 (N_996,In_187,In_622);
xor U997 (N_997,In_189,In_208);
nand U998 (N_998,In_680,In_103);
nor U999 (N_999,In_351,In_739);
and U1000 (N_1000,In_553,In_365);
xor U1001 (N_1001,In_334,In_951);
nand U1002 (N_1002,In_251,In_931);
and U1003 (N_1003,In_561,In_426);
nor U1004 (N_1004,In_673,In_375);
nand U1005 (N_1005,In_834,In_906);
and U1006 (N_1006,In_294,In_779);
nor U1007 (N_1007,In_404,In_658);
xor U1008 (N_1008,In_878,In_157);
nand U1009 (N_1009,In_46,In_331);
nand U1010 (N_1010,In_526,In_336);
or U1011 (N_1011,In_881,In_294);
nor U1012 (N_1012,In_715,In_851);
xor U1013 (N_1013,In_715,In_329);
or U1014 (N_1014,In_988,In_839);
xnor U1015 (N_1015,In_660,In_416);
nand U1016 (N_1016,In_100,In_608);
nor U1017 (N_1017,In_354,In_565);
or U1018 (N_1018,In_368,In_857);
and U1019 (N_1019,In_58,In_594);
xnor U1020 (N_1020,In_161,In_906);
nor U1021 (N_1021,In_851,In_290);
or U1022 (N_1022,In_349,In_18);
nand U1023 (N_1023,In_625,In_842);
nand U1024 (N_1024,In_902,In_73);
xnor U1025 (N_1025,In_724,In_177);
or U1026 (N_1026,In_396,In_485);
xor U1027 (N_1027,In_297,In_916);
nand U1028 (N_1028,In_808,In_79);
or U1029 (N_1029,In_964,In_956);
xnor U1030 (N_1030,In_408,In_305);
nand U1031 (N_1031,In_798,In_551);
nor U1032 (N_1032,In_754,In_472);
nand U1033 (N_1033,In_12,In_260);
nand U1034 (N_1034,In_9,In_129);
and U1035 (N_1035,In_644,In_77);
or U1036 (N_1036,In_628,In_724);
or U1037 (N_1037,In_968,In_86);
and U1038 (N_1038,In_643,In_646);
and U1039 (N_1039,In_103,In_381);
nor U1040 (N_1040,In_857,In_120);
nor U1041 (N_1041,In_100,In_203);
nand U1042 (N_1042,In_712,In_339);
and U1043 (N_1043,In_275,In_908);
and U1044 (N_1044,In_251,In_881);
and U1045 (N_1045,In_324,In_617);
and U1046 (N_1046,In_280,In_340);
xnor U1047 (N_1047,In_22,In_835);
or U1048 (N_1048,In_858,In_495);
nor U1049 (N_1049,In_868,In_793);
and U1050 (N_1050,In_973,In_864);
nand U1051 (N_1051,In_689,In_756);
or U1052 (N_1052,In_61,In_965);
or U1053 (N_1053,In_561,In_169);
and U1054 (N_1054,In_868,In_53);
xnor U1055 (N_1055,In_721,In_929);
nor U1056 (N_1056,In_61,In_722);
nand U1057 (N_1057,In_836,In_803);
or U1058 (N_1058,In_691,In_758);
nand U1059 (N_1059,In_869,In_203);
or U1060 (N_1060,In_168,In_448);
nor U1061 (N_1061,In_551,In_129);
and U1062 (N_1062,In_581,In_298);
nand U1063 (N_1063,In_624,In_867);
or U1064 (N_1064,In_265,In_289);
nor U1065 (N_1065,In_708,In_514);
and U1066 (N_1066,In_751,In_278);
or U1067 (N_1067,In_529,In_2);
xor U1068 (N_1068,In_404,In_211);
xnor U1069 (N_1069,In_878,In_165);
nand U1070 (N_1070,In_351,In_309);
or U1071 (N_1071,In_638,In_606);
or U1072 (N_1072,In_560,In_893);
and U1073 (N_1073,In_372,In_21);
nor U1074 (N_1074,In_818,In_739);
nand U1075 (N_1075,In_638,In_1);
xnor U1076 (N_1076,In_426,In_908);
nand U1077 (N_1077,In_689,In_261);
nand U1078 (N_1078,In_648,In_188);
nor U1079 (N_1079,In_333,In_551);
nor U1080 (N_1080,In_954,In_335);
nor U1081 (N_1081,In_157,In_679);
nand U1082 (N_1082,In_856,In_804);
and U1083 (N_1083,In_648,In_257);
and U1084 (N_1084,In_452,In_522);
nor U1085 (N_1085,In_482,In_796);
or U1086 (N_1086,In_400,In_858);
or U1087 (N_1087,In_771,In_367);
nor U1088 (N_1088,In_433,In_163);
nand U1089 (N_1089,In_133,In_759);
and U1090 (N_1090,In_288,In_68);
nor U1091 (N_1091,In_114,In_207);
xnor U1092 (N_1092,In_625,In_758);
xor U1093 (N_1093,In_523,In_164);
nor U1094 (N_1094,In_544,In_92);
and U1095 (N_1095,In_71,In_800);
nand U1096 (N_1096,In_179,In_186);
and U1097 (N_1097,In_320,In_557);
xor U1098 (N_1098,In_963,In_486);
xnor U1099 (N_1099,In_15,In_416);
or U1100 (N_1100,In_372,In_934);
and U1101 (N_1101,In_845,In_621);
xnor U1102 (N_1102,In_989,In_977);
xnor U1103 (N_1103,In_923,In_876);
nand U1104 (N_1104,In_296,In_227);
and U1105 (N_1105,In_784,In_721);
nor U1106 (N_1106,In_825,In_920);
xnor U1107 (N_1107,In_854,In_660);
or U1108 (N_1108,In_963,In_676);
xor U1109 (N_1109,In_27,In_659);
or U1110 (N_1110,In_919,In_504);
nand U1111 (N_1111,In_502,In_909);
and U1112 (N_1112,In_45,In_504);
xor U1113 (N_1113,In_474,In_603);
nand U1114 (N_1114,In_221,In_266);
and U1115 (N_1115,In_153,In_388);
nand U1116 (N_1116,In_684,In_895);
xnor U1117 (N_1117,In_474,In_569);
xor U1118 (N_1118,In_150,In_504);
xor U1119 (N_1119,In_652,In_821);
nand U1120 (N_1120,In_656,In_4);
xor U1121 (N_1121,In_111,In_366);
xnor U1122 (N_1122,In_241,In_277);
or U1123 (N_1123,In_574,In_463);
nor U1124 (N_1124,In_37,In_210);
nand U1125 (N_1125,In_239,In_127);
and U1126 (N_1126,In_470,In_133);
xnor U1127 (N_1127,In_536,In_778);
or U1128 (N_1128,In_432,In_313);
or U1129 (N_1129,In_524,In_33);
and U1130 (N_1130,In_293,In_123);
and U1131 (N_1131,In_234,In_195);
nor U1132 (N_1132,In_702,In_274);
or U1133 (N_1133,In_755,In_120);
or U1134 (N_1134,In_171,In_998);
or U1135 (N_1135,In_133,In_776);
xor U1136 (N_1136,In_496,In_927);
or U1137 (N_1137,In_251,In_27);
nor U1138 (N_1138,In_241,In_227);
nor U1139 (N_1139,In_466,In_142);
and U1140 (N_1140,In_921,In_499);
and U1141 (N_1141,In_80,In_505);
xnor U1142 (N_1142,In_648,In_442);
or U1143 (N_1143,In_707,In_864);
nand U1144 (N_1144,In_841,In_90);
nand U1145 (N_1145,In_275,In_537);
nand U1146 (N_1146,In_654,In_228);
nand U1147 (N_1147,In_695,In_275);
nor U1148 (N_1148,In_468,In_852);
and U1149 (N_1149,In_43,In_169);
xor U1150 (N_1150,In_993,In_785);
and U1151 (N_1151,In_617,In_615);
and U1152 (N_1152,In_386,In_509);
nand U1153 (N_1153,In_825,In_618);
and U1154 (N_1154,In_527,In_296);
xor U1155 (N_1155,In_585,In_928);
or U1156 (N_1156,In_938,In_839);
nor U1157 (N_1157,In_725,In_581);
nand U1158 (N_1158,In_113,In_984);
and U1159 (N_1159,In_163,In_784);
nand U1160 (N_1160,In_905,In_870);
nand U1161 (N_1161,In_174,In_609);
xor U1162 (N_1162,In_875,In_780);
xor U1163 (N_1163,In_646,In_431);
and U1164 (N_1164,In_155,In_333);
xor U1165 (N_1165,In_902,In_365);
nor U1166 (N_1166,In_484,In_64);
nand U1167 (N_1167,In_271,In_973);
nor U1168 (N_1168,In_827,In_412);
xor U1169 (N_1169,In_848,In_79);
or U1170 (N_1170,In_509,In_374);
and U1171 (N_1171,In_372,In_593);
xor U1172 (N_1172,In_913,In_867);
nor U1173 (N_1173,In_818,In_468);
and U1174 (N_1174,In_766,In_200);
nor U1175 (N_1175,In_496,In_404);
and U1176 (N_1176,In_565,In_211);
nand U1177 (N_1177,In_598,In_719);
nor U1178 (N_1178,In_285,In_994);
nand U1179 (N_1179,In_165,In_360);
nand U1180 (N_1180,In_139,In_142);
nand U1181 (N_1181,In_108,In_310);
nand U1182 (N_1182,In_751,In_674);
nor U1183 (N_1183,In_116,In_94);
xnor U1184 (N_1184,In_848,In_751);
or U1185 (N_1185,In_452,In_797);
xor U1186 (N_1186,In_621,In_620);
and U1187 (N_1187,In_427,In_953);
nor U1188 (N_1188,In_537,In_25);
xnor U1189 (N_1189,In_411,In_966);
nand U1190 (N_1190,In_57,In_359);
xor U1191 (N_1191,In_373,In_318);
xnor U1192 (N_1192,In_559,In_662);
nand U1193 (N_1193,In_148,In_740);
or U1194 (N_1194,In_773,In_927);
xnor U1195 (N_1195,In_688,In_814);
xnor U1196 (N_1196,In_814,In_768);
or U1197 (N_1197,In_348,In_806);
nor U1198 (N_1198,In_394,In_175);
xor U1199 (N_1199,In_716,In_459);
xor U1200 (N_1200,In_319,In_75);
xnor U1201 (N_1201,In_98,In_374);
xnor U1202 (N_1202,In_631,In_829);
nand U1203 (N_1203,In_69,In_27);
or U1204 (N_1204,In_126,In_959);
and U1205 (N_1205,In_120,In_913);
nor U1206 (N_1206,In_545,In_352);
and U1207 (N_1207,In_677,In_792);
or U1208 (N_1208,In_1,In_43);
or U1209 (N_1209,In_955,In_647);
xnor U1210 (N_1210,In_399,In_200);
nand U1211 (N_1211,In_136,In_16);
nand U1212 (N_1212,In_109,In_577);
nor U1213 (N_1213,In_263,In_622);
xnor U1214 (N_1214,In_886,In_687);
or U1215 (N_1215,In_221,In_803);
xnor U1216 (N_1216,In_527,In_496);
nor U1217 (N_1217,In_699,In_586);
or U1218 (N_1218,In_444,In_194);
nor U1219 (N_1219,In_72,In_916);
xor U1220 (N_1220,In_214,In_249);
nand U1221 (N_1221,In_167,In_826);
or U1222 (N_1222,In_835,In_705);
nor U1223 (N_1223,In_293,In_498);
nor U1224 (N_1224,In_535,In_713);
nand U1225 (N_1225,In_558,In_333);
or U1226 (N_1226,In_365,In_761);
and U1227 (N_1227,In_715,In_257);
and U1228 (N_1228,In_521,In_574);
or U1229 (N_1229,In_40,In_485);
nand U1230 (N_1230,In_75,In_835);
nand U1231 (N_1231,In_200,In_357);
nor U1232 (N_1232,In_866,In_721);
xor U1233 (N_1233,In_32,In_795);
xor U1234 (N_1234,In_706,In_942);
or U1235 (N_1235,In_588,In_98);
xnor U1236 (N_1236,In_942,In_803);
or U1237 (N_1237,In_995,In_968);
nand U1238 (N_1238,In_835,In_776);
nand U1239 (N_1239,In_30,In_596);
nor U1240 (N_1240,In_335,In_90);
or U1241 (N_1241,In_27,In_933);
nor U1242 (N_1242,In_288,In_616);
nand U1243 (N_1243,In_751,In_99);
nor U1244 (N_1244,In_598,In_948);
nor U1245 (N_1245,In_716,In_698);
xor U1246 (N_1246,In_243,In_339);
and U1247 (N_1247,In_78,In_99);
xor U1248 (N_1248,In_162,In_473);
or U1249 (N_1249,In_618,In_886);
nand U1250 (N_1250,In_438,In_544);
nand U1251 (N_1251,In_791,In_236);
or U1252 (N_1252,In_489,In_891);
xnor U1253 (N_1253,In_199,In_529);
nand U1254 (N_1254,In_377,In_221);
and U1255 (N_1255,In_290,In_481);
xor U1256 (N_1256,In_923,In_549);
xor U1257 (N_1257,In_36,In_969);
and U1258 (N_1258,In_932,In_182);
xor U1259 (N_1259,In_7,In_171);
nor U1260 (N_1260,In_54,In_252);
nand U1261 (N_1261,In_394,In_700);
and U1262 (N_1262,In_70,In_871);
or U1263 (N_1263,In_600,In_324);
or U1264 (N_1264,In_287,In_278);
nand U1265 (N_1265,In_612,In_689);
nand U1266 (N_1266,In_991,In_296);
nor U1267 (N_1267,In_539,In_241);
nor U1268 (N_1268,In_500,In_445);
xnor U1269 (N_1269,In_219,In_904);
or U1270 (N_1270,In_212,In_504);
and U1271 (N_1271,In_871,In_516);
nand U1272 (N_1272,In_709,In_770);
nor U1273 (N_1273,In_100,In_493);
or U1274 (N_1274,In_540,In_114);
or U1275 (N_1275,In_792,In_33);
nand U1276 (N_1276,In_519,In_186);
xor U1277 (N_1277,In_352,In_89);
and U1278 (N_1278,In_194,In_322);
xor U1279 (N_1279,In_28,In_549);
or U1280 (N_1280,In_415,In_340);
nor U1281 (N_1281,In_860,In_157);
nor U1282 (N_1282,In_249,In_51);
and U1283 (N_1283,In_387,In_492);
and U1284 (N_1284,In_209,In_238);
or U1285 (N_1285,In_270,In_901);
nand U1286 (N_1286,In_891,In_361);
nand U1287 (N_1287,In_267,In_33);
or U1288 (N_1288,In_841,In_400);
xnor U1289 (N_1289,In_104,In_126);
and U1290 (N_1290,In_548,In_388);
or U1291 (N_1291,In_808,In_48);
or U1292 (N_1292,In_97,In_29);
or U1293 (N_1293,In_227,In_476);
nor U1294 (N_1294,In_992,In_962);
or U1295 (N_1295,In_607,In_233);
xnor U1296 (N_1296,In_875,In_895);
nand U1297 (N_1297,In_172,In_609);
nor U1298 (N_1298,In_144,In_810);
xnor U1299 (N_1299,In_352,In_109);
nand U1300 (N_1300,In_806,In_322);
and U1301 (N_1301,In_181,In_501);
nor U1302 (N_1302,In_86,In_275);
nor U1303 (N_1303,In_485,In_641);
xor U1304 (N_1304,In_964,In_994);
nand U1305 (N_1305,In_370,In_991);
or U1306 (N_1306,In_50,In_333);
nor U1307 (N_1307,In_511,In_715);
xnor U1308 (N_1308,In_871,In_881);
nand U1309 (N_1309,In_37,In_42);
and U1310 (N_1310,In_128,In_776);
or U1311 (N_1311,In_863,In_353);
nand U1312 (N_1312,In_246,In_651);
xnor U1313 (N_1313,In_541,In_72);
nand U1314 (N_1314,In_44,In_615);
xor U1315 (N_1315,In_626,In_524);
nand U1316 (N_1316,In_272,In_574);
and U1317 (N_1317,In_779,In_681);
or U1318 (N_1318,In_271,In_440);
xor U1319 (N_1319,In_946,In_74);
nand U1320 (N_1320,In_343,In_413);
nand U1321 (N_1321,In_175,In_874);
and U1322 (N_1322,In_661,In_535);
or U1323 (N_1323,In_842,In_943);
nor U1324 (N_1324,In_374,In_403);
and U1325 (N_1325,In_546,In_494);
nand U1326 (N_1326,In_204,In_469);
xor U1327 (N_1327,In_260,In_555);
xnor U1328 (N_1328,In_655,In_758);
or U1329 (N_1329,In_875,In_585);
xor U1330 (N_1330,In_798,In_648);
nand U1331 (N_1331,In_244,In_51);
or U1332 (N_1332,In_886,In_412);
xnor U1333 (N_1333,In_139,In_809);
and U1334 (N_1334,In_244,In_844);
nand U1335 (N_1335,In_98,In_398);
nand U1336 (N_1336,In_841,In_977);
and U1337 (N_1337,In_352,In_27);
or U1338 (N_1338,In_613,In_787);
nand U1339 (N_1339,In_811,In_577);
or U1340 (N_1340,In_884,In_229);
or U1341 (N_1341,In_133,In_531);
and U1342 (N_1342,In_963,In_859);
nor U1343 (N_1343,In_473,In_423);
and U1344 (N_1344,In_469,In_12);
or U1345 (N_1345,In_509,In_153);
or U1346 (N_1346,In_598,In_964);
and U1347 (N_1347,In_967,In_255);
xnor U1348 (N_1348,In_859,In_540);
xor U1349 (N_1349,In_689,In_698);
nor U1350 (N_1350,In_250,In_737);
and U1351 (N_1351,In_383,In_227);
or U1352 (N_1352,In_6,In_141);
or U1353 (N_1353,In_827,In_879);
and U1354 (N_1354,In_917,In_659);
or U1355 (N_1355,In_387,In_533);
or U1356 (N_1356,In_702,In_501);
nor U1357 (N_1357,In_593,In_338);
xnor U1358 (N_1358,In_219,In_797);
and U1359 (N_1359,In_40,In_555);
and U1360 (N_1360,In_962,In_855);
or U1361 (N_1361,In_618,In_616);
nor U1362 (N_1362,In_830,In_676);
nand U1363 (N_1363,In_645,In_762);
nor U1364 (N_1364,In_618,In_148);
xor U1365 (N_1365,In_515,In_113);
xor U1366 (N_1366,In_852,In_862);
xor U1367 (N_1367,In_358,In_386);
nand U1368 (N_1368,In_14,In_420);
nand U1369 (N_1369,In_41,In_277);
xor U1370 (N_1370,In_800,In_349);
xor U1371 (N_1371,In_160,In_468);
nor U1372 (N_1372,In_836,In_238);
and U1373 (N_1373,In_13,In_230);
xor U1374 (N_1374,In_549,In_869);
xor U1375 (N_1375,In_683,In_593);
nor U1376 (N_1376,In_807,In_295);
or U1377 (N_1377,In_871,In_807);
nor U1378 (N_1378,In_941,In_245);
and U1379 (N_1379,In_147,In_291);
or U1380 (N_1380,In_322,In_448);
or U1381 (N_1381,In_449,In_920);
or U1382 (N_1382,In_806,In_873);
and U1383 (N_1383,In_860,In_472);
nand U1384 (N_1384,In_406,In_702);
nor U1385 (N_1385,In_762,In_94);
nor U1386 (N_1386,In_840,In_648);
nand U1387 (N_1387,In_421,In_885);
nand U1388 (N_1388,In_297,In_483);
xor U1389 (N_1389,In_747,In_164);
nand U1390 (N_1390,In_630,In_79);
nand U1391 (N_1391,In_777,In_783);
nor U1392 (N_1392,In_639,In_657);
xnor U1393 (N_1393,In_815,In_939);
nand U1394 (N_1394,In_373,In_933);
nand U1395 (N_1395,In_706,In_703);
and U1396 (N_1396,In_547,In_626);
nand U1397 (N_1397,In_487,In_930);
nand U1398 (N_1398,In_680,In_694);
nand U1399 (N_1399,In_743,In_885);
or U1400 (N_1400,In_759,In_998);
nor U1401 (N_1401,In_281,In_185);
and U1402 (N_1402,In_25,In_769);
nand U1403 (N_1403,In_935,In_870);
and U1404 (N_1404,In_83,In_475);
nand U1405 (N_1405,In_793,In_944);
or U1406 (N_1406,In_144,In_550);
nand U1407 (N_1407,In_148,In_862);
or U1408 (N_1408,In_867,In_734);
and U1409 (N_1409,In_578,In_232);
nor U1410 (N_1410,In_58,In_322);
nor U1411 (N_1411,In_962,In_469);
nand U1412 (N_1412,In_90,In_514);
or U1413 (N_1413,In_759,In_552);
nand U1414 (N_1414,In_56,In_236);
nor U1415 (N_1415,In_991,In_245);
nand U1416 (N_1416,In_549,In_338);
nor U1417 (N_1417,In_380,In_408);
nor U1418 (N_1418,In_825,In_963);
xnor U1419 (N_1419,In_779,In_775);
nand U1420 (N_1420,In_418,In_982);
nand U1421 (N_1421,In_517,In_271);
or U1422 (N_1422,In_644,In_456);
or U1423 (N_1423,In_751,In_477);
and U1424 (N_1424,In_620,In_587);
and U1425 (N_1425,In_140,In_911);
nor U1426 (N_1426,In_786,In_151);
and U1427 (N_1427,In_885,In_618);
nand U1428 (N_1428,In_547,In_660);
or U1429 (N_1429,In_750,In_515);
nand U1430 (N_1430,In_735,In_201);
and U1431 (N_1431,In_952,In_632);
nand U1432 (N_1432,In_736,In_329);
or U1433 (N_1433,In_531,In_285);
nor U1434 (N_1434,In_555,In_188);
or U1435 (N_1435,In_813,In_999);
or U1436 (N_1436,In_195,In_877);
and U1437 (N_1437,In_17,In_104);
and U1438 (N_1438,In_611,In_62);
or U1439 (N_1439,In_853,In_723);
nor U1440 (N_1440,In_70,In_818);
nor U1441 (N_1441,In_793,In_263);
or U1442 (N_1442,In_478,In_848);
xnor U1443 (N_1443,In_873,In_96);
xor U1444 (N_1444,In_880,In_703);
and U1445 (N_1445,In_507,In_209);
and U1446 (N_1446,In_682,In_891);
xnor U1447 (N_1447,In_567,In_390);
nor U1448 (N_1448,In_755,In_35);
and U1449 (N_1449,In_77,In_984);
or U1450 (N_1450,In_643,In_422);
nand U1451 (N_1451,In_909,In_203);
nand U1452 (N_1452,In_795,In_429);
or U1453 (N_1453,In_379,In_875);
nor U1454 (N_1454,In_310,In_432);
xor U1455 (N_1455,In_733,In_6);
xor U1456 (N_1456,In_993,In_812);
nor U1457 (N_1457,In_708,In_845);
xnor U1458 (N_1458,In_422,In_613);
and U1459 (N_1459,In_348,In_905);
nor U1460 (N_1460,In_773,In_371);
xor U1461 (N_1461,In_672,In_708);
and U1462 (N_1462,In_865,In_538);
nor U1463 (N_1463,In_13,In_138);
nand U1464 (N_1464,In_943,In_193);
xnor U1465 (N_1465,In_748,In_150);
and U1466 (N_1466,In_586,In_60);
nand U1467 (N_1467,In_258,In_633);
nor U1468 (N_1468,In_713,In_353);
nor U1469 (N_1469,In_405,In_367);
nor U1470 (N_1470,In_246,In_187);
nand U1471 (N_1471,In_655,In_319);
nand U1472 (N_1472,In_874,In_783);
and U1473 (N_1473,In_887,In_822);
or U1474 (N_1474,In_591,In_568);
or U1475 (N_1475,In_200,In_944);
nand U1476 (N_1476,In_525,In_640);
nor U1477 (N_1477,In_706,In_994);
nor U1478 (N_1478,In_182,In_545);
or U1479 (N_1479,In_186,In_163);
xor U1480 (N_1480,In_255,In_248);
xnor U1481 (N_1481,In_38,In_149);
nand U1482 (N_1482,In_958,In_342);
xor U1483 (N_1483,In_834,In_556);
xnor U1484 (N_1484,In_97,In_836);
nand U1485 (N_1485,In_853,In_860);
and U1486 (N_1486,In_777,In_584);
nand U1487 (N_1487,In_431,In_949);
and U1488 (N_1488,In_772,In_402);
nand U1489 (N_1489,In_847,In_879);
or U1490 (N_1490,In_64,In_602);
nand U1491 (N_1491,In_987,In_780);
xnor U1492 (N_1492,In_297,In_254);
nor U1493 (N_1493,In_568,In_527);
nor U1494 (N_1494,In_931,In_516);
nand U1495 (N_1495,In_188,In_224);
and U1496 (N_1496,In_140,In_320);
xnor U1497 (N_1497,In_757,In_277);
xor U1498 (N_1498,In_941,In_649);
and U1499 (N_1499,In_217,In_319);
nor U1500 (N_1500,In_207,In_171);
nand U1501 (N_1501,In_463,In_290);
nor U1502 (N_1502,In_562,In_803);
nand U1503 (N_1503,In_353,In_650);
or U1504 (N_1504,In_792,In_43);
xnor U1505 (N_1505,In_617,In_718);
xnor U1506 (N_1506,In_605,In_217);
xnor U1507 (N_1507,In_582,In_571);
nand U1508 (N_1508,In_711,In_54);
xnor U1509 (N_1509,In_588,In_362);
nand U1510 (N_1510,In_667,In_127);
nor U1511 (N_1511,In_163,In_192);
xor U1512 (N_1512,In_877,In_942);
xor U1513 (N_1513,In_948,In_593);
nand U1514 (N_1514,In_315,In_956);
and U1515 (N_1515,In_801,In_613);
xor U1516 (N_1516,In_152,In_912);
xnor U1517 (N_1517,In_278,In_142);
nand U1518 (N_1518,In_519,In_624);
and U1519 (N_1519,In_891,In_140);
or U1520 (N_1520,In_783,In_564);
nor U1521 (N_1521,In_602,In_309);
nand U1522 (N_1522,In_408,In_908);
and U1523 (N_1523,In_925,In_744);
or U1524 (N_1524,In_828,In_853);
and U1525 (N_1525,In_391,In_973);
or U1526 (N_1526,In_883,In_592);
or U1527 (N_1527,In_91,In_177);
nand U1528 (N_1528,In_134,In_35);
or U1529 (N_1529,In_6,In_770);
nand U1530 (N_1530,In_799,In_562);
nand U1531 (N_1531,In_51,In_468);
nand U1532 (N_1532,In_326,In_77);
and U1533 (N_1533,In_349,In_88);
nor U1534 (N_1534,In_35,In_988);
xnor U1535 (N_1535,In_503,In_644);
or U1536 (N_1536,In_709,In_84);
nand U1537 (N_1537,In_282,In_612);
or U1538 (N_1538,In_129,In_829);
nor U1539 (N_1539,In_894,In_270);
or U1540 (N_1540,In_15,In_420);
and U1541 (N_1541,In_431,In_250);
or U1542 (N_1542,In_459,In_642);
or U1543 (N_1543,In_660,In_424);
or U1544 (N_1544,In_577,In_364);
nor U1545 (N_1545,In_805,In_329);
or U1546 (N_1546,In_996,In_988);
xnor U1547 (N_1547,In_574,In_285);
and U1548 (N_1548,In_620,In_904);
and U1549 (N_1549,In_757,In_560);
nand U1550 (N_1550,In_228,In_946);
nor U1551 (N_1551,In_871,In_727);
xnor U1552 (N_1552,In_85,In_822);
and U1553 (N_1553,In_924,In_329);
xnor U1554 (N_1554,In_152,In_103);
nand U1555 (N_1555,In_185,In_740);
xnor U1556 (N_1556,In_239,In_334);
nor U1557 (N_1557,In_624,In_793);
nand U1558 (N_1558,In_91,In_610);
nand U1559 (N_1559,In_136,In_425);
xor U1560 (N_1560,In_877,In_109);
nand U1561 (N_1561,In_416,In_555);
xor U1562 (N_1562,In_207,In_337);
or U1563 (N_1563,In_823,In_124);
nand U1564 (N_1564,In_719,In_901);
nor U1565 (N_1565,In_513,In_848);
nor U1566 (N_1566,In_664,In_743);
xor U1567 (N_1567,In_46,In_906);
xnor U1568 (N_1568,In_133,In_59);
nor U1569 (N_1569,In_188,In_890);
xnor U1570 (N_1570,In_898,In_661);
nand U1571 (N_1571,In_464,In_598);
and U1572 (N_1572,In_718,In_720);
and U1573 (N_1573,In_88,In_395);
nor U1574 (N_1574,In_657,In_783);
nor U1575 (N_1575,In_305,In_287);
or U1576 (N_1576,In_303,In_378);
or U1577 (N_1577,In_194,In_632);
and U1578 (N_1578,In_58,In_564);
and U1579 (N_1579,In_46,In_236);
and U1580 (N_1580,In_393,In_484);
nor U1581 (N_1581,In_653,In_742);
nor U1582 (N_1582,In_342,In_297);
nor U1583 (N_1583,In_174,In_568);
nor U1584 (N_1584,In_780,In_503);
or U1585 (N_1585,In_399,In_878);
xnor U1586 (N_1586,In_795,In_848);
or U1587 (N_1587,In_424,In_810);
and U1588 (N_1588,In_913,In_632);
and U1589 (N_1589,In_109,In_528);
xnor U1590 (N_1590,In_692,In_246);
and U1591 (N_1591,In_178,In_348);
and U1592 (N_1592,In_538,In_623);
xnor U1593 (N_1593,In_584,In_179);
xor U1594 (N_1594,In_448,In_467);
and U1595 (N_1595,In_649,In_161);
nor U1596 (N_1596,In_896,In_223);
and U1597 (N_1597,In_970,In_817);
or U1598 (N_1598,In_751,In_303);
and U1599 (N_1599,In_792,In_55);
nor U1600 (N_1600,In_204,In_190);
nand U1601 (N_1601,In_107,In_412);
or U1602 (N_1602,In_865,In_550);
nand U1603 (N_1603,In_889,In_166);
and U1604 (N_1604,In_978,In_766);
nand U1605 (N_1605,In_113,In_34);
or U1606 (N_1606,In_354,In_57);
nor U1607 (N_1607,In_133,In_109);
nand U1608 (N_1608,In_409,In_600);
or U1609 (N_1609,In_79,In_538);
nor U1610 (N_1610,In_246,In_727);
nand U1611 (N_1611,In_523,In_916);
and U1612 (N_1612,In_666,In_13);
nor U1613 (N_1613,In_472,In_294);
or U1614 (N_1614,In_846,In_353);
and U1615 (N_1615,In_62,In_44);
nand U1616 (N_1616,In_541,In_424);
and U1617 (N_1617,In_577,In_487);
xor U1618 (N_1618,In_485,In_626);
and U1619 (N_1619,In_449,In_497);
nor U1620 (N_1620,In_981,In_55);
and U1621 (N_1621,In_699,In_241);
and U1622 (N_1622,In_200,In_4);
nor U1623 (N_1623,In_924,In_343);
and U1624 (N_1624,In_955,In_208);
nand U1625 (N_1625,In_0,In_434);
xor U1626 (N_1626,In_944,In_383);
nand U1627 (N_1627,In_325,In_885);
or U1628 (N_1628,In_213,In_431);
or U1629 (N_1629,In_103,In_954);
nand U1630 (N_1630,In_611,In_138);
and U1631 (N_1631,In_544,In_94);
and U1632 (N_1632,In_729,In_314);
and U1633 (N_1633,In_164,In_123);
nand U1634 (N_1634,In_129,In_657);
or U1635 (N_1635,In_524,In_726);
nand U1636 (N_1636,In_292,In_727);
or U1637 (N_1637,In_89,In_808);
nor U1638 (N_1638,In_775,In_276);
xnor U1639 (N_1639,In_691,In_394);
xnor U1640 (N_1640,In_596,In_573);
nand U1641 (N_1641,In_344,In_577);
xor U1642 (N_1642,In_43,In_902);
nand U1643 (N_1643,In_80,In_578);
xnor U1644 (N_1644,In_301,In_788);
or U1645 (N_1645,In_555,In_360);
nand U1646 (N_1646,In_753,In_495);
nand U1647 (N_1647,In_779,In_778);
nand U1648 (N_1648,In_551,In_449);
and U1649 (N_1649,In_471,In_854);
nand U1650 (N_1650,In_974,In_453);
and U1651 (N_1651,In_753,In_507);
xnor U1652 (N_1652,In_590,In_93);
and U1653 (N_1653,In_207,In_605);
and U1654 (N_1654,In_997,In_427);
or U1655 (N_1655,In_980,In_329);
nand U1656 (N_1656,In_72,In_99);
nand U1657 (N_1657,In_829,In_862);
or U1658 (N_1658,In_734,In_31);
nand U1659 (N_1659,In_490,In_888);
nor U1660 (N_1660,In_542,In_33);
or U1661 (N_1661,In_86,In_468);
or U1662 (N_1662,In_32,In_239);
nand U1663 (N_1663,In_140,In_838);
xnor U1664 (N_1664,In_277,In_225);
nor U1665 (N_1665,In_473,In_821);
nand U1666 (N_1666,In_914,In_953);
nor U1667 (N_1667,In_187,In_886);
nand U1668 (N_1668,In_208,In_78);
xor U1669 (N_1669,In_12,In_265);
nor U1670 (N_1670,In_647,In_841);
or U1671 (N_1671,In_101,In_549);
nand U1672 (N_1672,In_283,In_352);
nor U1673 (N_1673,In_267,In_887);
xor U1674 (N_1674,In_58,In_944);
nand U1675 (N_1675,In_524,In_639);
or U1676 (N_1676,In_766,In_575);
nand U1677 (N_1677,In_379,In_753);
xor U1678 (N_1678,In_40,In_387);
nor U1679 (N_1679,In_548,In_664);
or U1680 (N_1680,In_258,In_393);
xor U1681 (N_1681,In_499,In_675);
xnor U1682 (N_1682,In_876,In_992);
nor U1683 (N_1683,In_551,In_166);
or U1684 (N_1684,In_487,In_452);
nor U1685 (N_1685,In_72,In_586);
nor U1686 (N_1686,In_220,In_246);
and U1687 (N_1687,In_443,In_260);
nor U1688 (N_1688,In_857,In_143);
nand U1689 (N_1689,In_501,In_582);
nand U1690 (N_1690,In_748,In_204);
nand U1691 (N_1691,In_499,In_843);
xnor U1692 (N_1692,In_785,In_958);
nor U1693 (N_1693,In_364,In_500);
and U1694 (N_1694,In_918,In_164);
or U1695 (N_1695,In_816,In_458);
xor U1696 (N_1696,In_407,In_712);
and U1697 (N_1697,In_513,In_553);
nor U1698 (N_1698,In_159,In_438);
nor U1699 (N_1699,In_229,In_282);
nor U1700 (N_1700,In_718,In_901);
nor U1701 (N_1701,In_65,In_974);
or U1702 (N_1702,In_174,In_213);
xor U1703 (N_1703,In_4,In_794);
or U1704 (N_1704,In_505,In_498);
and U1705 (N_1705,In_233,In_37);
or U1706 (N_1706,In_527,In_920);
xor U1707 (N_1707,In_366,In_92);
or U1708 (N_1708,In_75,In_291);
nor U1709 (N_1709,In_479,In_111);
or U1710 (N_1710,In_401,In_300);
nor U1711 (N_1711,In_378,In_22);
xor U1712 (N_1712,In_63,In_846);
or U1713 (N_1713,In_508,In_447);
nand U1714 (N_1714,In_910,In_243);
nand U1715 (N_1715,In_792,In_147);
nand U1716 (N_1716,In_43,In_494);
or U1717 (N_1717,In_504,In_720);
nor U1718 (N_1718,In_764,In_166);
or U1719 (N_1719,In_775,In_509);
or U1720 (N_1720,In_595,In_997);
xor U1721 (N_1721,In_643,In_513);
and U1722 (N_1722,In_133,In_959);
xnor U1723 (N_1723,In_924,In_821);
or U1724 (N_1724,In_923,In_962);
xnor U1725 (N_1725,In_197,In_831);
or U1726 (N_1726,In_741,In_17);
and U1727 (N_1727,In_878,In_938);
xor U1728 (N_1728,In_426,In_356);
or U1729 (N_1729,In_493,In_212);
nand U1730 (N_1730,In_302,In_907);
or U1731 (N_1731,In_615,In_568);
and U1732 (N_1732,In_808,In_297);
nor U1733 (N_1733,In_278,In_613);
nand U1734 (N_1734,In_950,In_504);
nand U1735 (N_1735,In_781,In_999);
or U1736 (N_1736,In_768,In_906);
nor U1737 (N_1737,In_734,In_997);
xor U1738 (N_1738,In_296,In_322);
or U1739 (N_1739,In_889,In_663);
nand U1740 (N_1740,In_594,In_978);
xor U1741 (N_1741,In_673,In_315);
xnor U1742 (N_1742,In_885,In_181);
xnor U1743 (N_1743,In_212,In_668);
and U1744 (N_1744,In_793,In_713);
or U1745 (N_1745,In_564,In_652);
xor U1746 (N_1746,In_360,In_425);
nand U1747 (N_1747,In_653,In_320);
and U1748 (N_1748,In_224,In_587);
nand U1749 (N_1749,In_998,In_26);
or U1750 (N_1750,In_367,In_829);
xnor U1751 (N_1751,In_574,In_189);
and U1752 (N_1752,In_260,In_33);
or U1753 (N_1753,In_105,In_91);
xor U1754 (N_1754,In_608,In_744);
and U1755 (N_1755,In_921,In_825);
nand U1756 (N_1756,In_336,In_157);
nand U1757 (N_1757,In_581,In_311);
nor U1758 (N_1758,In_489,In_611);
xnor U1759 (N_1759,In_388,In_716);
nor U1760 (N_1760,In_972,In_394);
and U1761 (N_1761,In_702,In_545);
and U1762 (N_1762,In_842,In_705);
or U1763 (N_1763,In_945,In_653);
xor U1764 (N_1764,In_12,In_55);
nand U1765 (N_1765,In_647,In_312);
xor U1766 (N_1766,In_94,In_289);
nor U1767 (N_1767,In_583,In_357);
nand U1768 (N_1768,In_834,In_895);
or U1769 (N_1769,In_791,In_559);
nand U1770 (N_1770,In_767,In_421);
nand U1771 (N_1771,In_439,In_424);
xor U1772 (N_1772,In_782,In_722);
or U1773 (N_1773,In_678,In_589);
and U1774 (N_1774,In_927,In_801);
xnor U1775 (N_1775,In_745,In_421);
and U1776 (N_1776,In_671,In_932);
and U1777 (N_1777,In_844,In_854);
xnor U1778 (N_1778,In_792,In_887);
or U1779 (N_1779,In_62,In_372);
nor U1780 (N_1780,In_60,In_103);
xor U1781 (N_1781,In_964,In_540);
or U1782 (N_1782,In_752,In_325);
xor U1783 (N_1783,In_547,In_307);
and U1784 (N_1784,In_731,In_699);
xor U1785 (N_1785,In_641,In_184);
or U1786 (N_1786,In_983,In_193);
xnor U1787 (N_1787,In_618,In_288);
nand U1788 (N_1788,In_849,In_860);
xnor U1789 (N_1789,In_516,In_379);
and U1790 (N_1790,In_162,In_45);
xor U1791 (N_1791,In_696,In_900);
nand U1792 (N_1792,In_153,In_369);
or U1793 (N_1793,In_430,In_85);
and U1794 (N_1794,In_424,In_557);
or U1795 (N_1795,In_715,In_27);
nor U1796 (N_1796,In_23,In_616);
xnor U1797 (N_1797,In_860,In_672);
nor U1798 (N_1798,In_39,In_180);
nand U1799 (N_1799,In_229,In_972);
and U1800 (N_1800,In_134,In_953);
and U1801 (N_1801,In_317,In_261);
xnor U1802 (N_1802,In_481,In_85);
or U1803 (N_1803,In_106,In_551);
or U1804 (N_1804,In_16,In_989);
or U1805 (N_1805,In_497,In_457);
and U1806 (N_1806,In_469,In_346);
nand U1807 (N_1807,In_694,In_302);
nor U1808 (N_1808,In_920,In_305);
nor U1809 (N_1809,In_892,In_763);
nand U1810 (N_1810,In_647,In_856);
nor U1811 (N_1811,In_260,In_276);
xor U1812 (N_1812,In_891,In_135);
nor U1813 (N_1813,In_224,In_586);
and U1814 (N_1814,In_142,In_158);
and U1815 (N_1815,In_76,In_575);
or U1816 (N_1816,In_498,In_943);
nor U1817 (N_1817,In_734,In_837);
or U1818 (N_1818,In_616,In_160);
or U1819 (N_1819,In_233,In_556);
or U1820 (N_1820,In_497,In_388);
and U1821 (N_1821,In_188,In_760);
nand U1822 (N_1822,In_874,In_682);
nor U1823 (N_1823,In_60,In_349);
nor U1824 (N_1824,In_553,In_883);
xnor U1825 (N_1825,In_43,In_979);
or U1826 (N_1826,In_13,In_396);
or U1827 (N_1827,In_734,In_130);
xor U1828 (N_1828,In_680,In_243);
nor U1829 (N_1829,In_997,In_586);
nor U1830 (N_1830,In_813,In_993);
and U1831 (N_1831,In_904,In_673);
nor U1832 (N_1832,In_99,In_136);
nor U1833 (N_1833,In_37,In_285);
nor U1834 (N_1834,In_624,In_973);
nand U1835 (N_1835,In_676,In_736);
nand U1836 (N_1836,In_540,In_828);
or U1837 (N_1837,In_514,In_192);
nor U1838 (N_1838,In_721,In_620);
nor U1839 (N_1839,In_805,In_783);
nand U1840 (N_1840,In_470,In_796);
or U1841 (N_1841,In_978,In_565);
or U1842 (N_1842,In_842,In_633);
or U1843 (N_1843,In_686,In_173);
or U1844 (N_1844,In_645,In_862);
nand U1845 (N_1845,In_537,In_692);
or U1846 (N_1846,In_439,In_514);
nand U1847 (N_1847,In_692,In_989);
nor U1848 (N_1848,In_522,In_934);
nand U1849 (N_1849,In_707,In_364);
or U1850 (N_1850,In_376,In_943);
and U1851 (N_1851,In_531,In_640);
and U1852 (N_1852,In_770,In_300);
nor U1853 (N_1853,In_764,In_118);
xnor U1854 (N_1854,In_80,In_748);
and U1855 (N_1855,In_80,In_218);
nor U1856 (N_1856,In_355,In_108);
nand U1857 (N_1857,In_458,In_463);
and U1858 (N_1858,In_807,In_329);
nand U1859 (N_1859,In_802,In_599);
or U1860 (N_1860,In_664,In_991);
or U1861 (N_1861,In_391,In_932);
and U1862 (N_1862,In_624,In_869);
nand U1863 (N_1863,In_885,In_362);
and U1864 (N_1864,In_900,In_534);
or U1865 (N_1865,In_288,In_705);
nand U1866 (N_1866,In_726,In_690);
and U1867 (N_1867,In_548,In_399);
nor U1868 (N_1868,In_142,In_131);
and U1869 (N_1869,In_15,In_9);
nor U1870 (N_1870,In_824,In_555);
nand U1871 (N_1871,In_931,In_838);
or U1872 (N_1872,In_387,In_69);
or U1873 (N_1873,In_423,In_974);
and U1874 (N_1874,In_662,In_446);
or U1875 (N_1875,In_289,In_208);
nand U1876 (N_1876,In_777,In_198);
nor U1877 (N_1877,In_685,In_353);
and U1878 (N_1878,In_225,In_197);
and U1879 (N_1879,In_414,In_766);
xor U1880 (N_1880,In_991,In_127);
or U1881 (N_1881,In_946,In_512);
and U1882 (N_1882,In_938,In_672);
nand U1883 (N_1883,In_15,In_52);
nand U1884 (N_1884,In_896,In_77);
and U1885 (N_1885,In_404,In_569);
nor U1886 (N_1886,In_135,In_502);
or U1887 (N_1887,In_279,In_714);
xor U1888 (N_1888,In_881,In_962);
or U1889 (N_1889,In_50,In_285);
nor U1890 (N_1890,In_349,In_431);
xor U1891 (N_1891,In_774,In_969);
xnor U1892 (N_1892,In_604,In_169);
or U1893 (N_1893,In_46,In_229);
nand U1894 (N_1894,In_314,In_957);
or U1895 (N_1895,In_741,In_415);
or U1896 (N_1896,In_911,In_143);
or U1897 (N_1897,In_988,In_602);
xor U1898 (N_1898,In_604,In_764);
nand U1899 (N_1899,In_650,In_634);
xor U1900 (N_1900,In_94,In_569);
or U1901 (N_1901,In_944,In_327);
and U1902 (N_1902,In_410,In_223);
and U1903 (N_1903,In_833,In_258);
and U1904 (N_1904,In_68,In_432);
nand U1905 (N_1905,In_596,In_595);
and U1906 (N_1906,In_168,In_846);
and U1907 (N_1907,In_975,In_83);
nor U1908 (N_1908,In_422,In_549);
or U1909 (N_1909,In_233,In_156);
nor U1910 (N_1910,In_743,In_943);
and U1911 (N_1911,In_443,In_303);
and U1912 (N_1912,In_705,In_228);
xnor U1913 (N_1913,In_856,In_585);
or U1914 (N_1914,In_953,In_282);
or U1915 (N_1915,In_581,In_474);
nand U1916 (N_1916,In_762,In_754);
and U1917 (N_1917,In_328,In_748);
nand U1918 (N_1918,In_343,In_605);
and U1919 (N_1919,In_126,In_649);
and U1920 (N_1920,In_261,In_323);
xor U1921 (N_1921,In_822,In_394);
and U1922 (N_1922,In_852,In_746);
nand U1923 (N_1923,In_743,In_247);
or U1924 (N_1924,In_186,In_444);
nand U1925 (N_1925,In_947,In_131);
xor U1926 (N_1926,In_927,In_839);
xor U1927 (N_1927,In_253,In_831);
or U1928 (N_1928,In_394,In_991);
nand U1929 (N_1929,In_312,In_465);
and U1930 (N_1930,In_137,In_939);
and U1931 (N_1931,In_189,In_171);
or U1932 (N_1932,In_287,In_624);
nand U1933 (N_1933,In_50,In_759);
and U1934 (N_1934,In_336,In_570);
xnor U1935 (N_1935,In_357,In_727);
and U1936 (N_1936,In_903,In_374);
nand U1937 (N_1937,In_180,In_50);
xnor U1938 (N_1938,In_632,In_839);
and U1939 (N_1939,In_747,In_755);
and U1940 (N_1940,In_57,In_490);
nor U1941 (N_1941,In_801,In_90);
and U1942 (N_1942,In_921,In_540);
and U1943 (N_1943,In_664,In_604);
and U1944 (N_1944,In_228,In_324);
or U1945 (N_1945,In_399,In_657);
and U1946 (N_1946,In_653,In_581);
and U1947 (N_1947,In_7,In_80);
xor U1948 (N_1948,In_4,In_161);
and U1949 (N_1949,In_987,In_501);
xnor U1950 (N_1950,In_456,In_678);
xnor U1951 (N_1951,In_115,In_284);
and U1952 (N_1952,In_632,In_388);
and U1953 (N_1953,In_908,In_240);
or U1954 (N_1954,In_466,In_457);
xor U1955 (N_1955,In_866,In_496);
nand U1956 (N_1956,In_545,In_964);
nand U1957 (N_1957,In_196,In_332);
nand U1958 (N_1958,In_868,In_993);
or U1959 (N_1959,In_261,In_510);
nand U1960 (N_1960,In_65,In_929);
and U1961 (N_1961,In_990,In_142);
nand U1962 (N_1962,In_214,In_62);
or U1963 (N_1963,In_995,In_885);
nor U1964 (N_1964,In_517,In_590);
nand U1965 (N_1965,In_595,In_932);
nor U1966 (N_1966,In_323,In_195);
and U1967 (N_1967,In_267,In_391);
and U1968 (N_1968,In_973,In_15);
or U1969 (N_1969,In_97,In_431);
nor U1970 (N_1970,In_331,In_829);
nand U1971 (N_1971,In_962,In_368);
or U1972 (N_1972,In_904,In_14);
and U1973 (N_1973,In_368,In_649);
or U1974 (N_1974,In_805,In_76);
nor U1975 (N_1975,In_102,In_305);
or U1976 (N_1976,In_395,In_581);
xor U1977 (N_1977,In_390,In_444);
or U1978 (N_1978,In_446,In_645);
or U1979 (N_1979,In_24,In_214);
nand U1980 (N_1980,In_866,In_324);
nor U1981 (N_1981,In_537,In_466);
nand U1982 (N_1982,In_587,In_64);
xnor U1983 (N_1983,In_263,In_900);
nand U1984 (N_1984,In_591,In_787);
xnor U1985 (N_1985,In_815,In_318);
nor U1986 (N_1986,In_8,In_258);
and U1987 (N_1987,In_43,In_600);
or U1988 (N_1988,In_93,In_163);
xor U1989 (N_1989,In_505,In_569);
nor U1990 (N_1990,In_269,In_672);
nor U1991 (N_1991,In_125,In_704);
or U1992 (N_1992,In_665,In_975);
and U1993 (N_1993,In_7,In_345);
xor U1994 (N_1994,In_892,In_110);
nor U1995 (N_1995,In_829,In_91);
and U1996 (N_1996,In_476,In_62);
and U1997 (N_1997,In_139,In_516);
nand U1998 (N_1998,In_628,In_702);
xnor U1999 (N_1999,In_161,In_48);
or U2000 (N_2000,In_57,In_349);
nor U2001 (N_2001,In_186,In_333);
xor U2002 (N_2002,In_526,In_280);
and U2003 (N_2003,In_105,In_677);
xor U2004 (N_2004,In_814,In_846);
nand U2005 (N_2005,In_934,In_505);
nand U2006 (N_2006,In_703,In_666);
nor U2007 (N_2007,In_96,In_268);
nand U2008 (N_2008,In_437,In_661);
nand U2009 (N_2009,In_759,In_838);
and U2010 (N_2010,In_887,In_102);
xor U2011 (N_2011,In_883,In_850);
xnor U2012 (N_2012,In_76,In_207);
or U2013 (N_2013,In_424,In_203);
and U2014 (N_2014,In_188,In_723);
and U2015 (N_2015,In_562,In_996);
xor U2016 (N_2016,In_666,In_486);
nand U2017 (N_2017,In_147,In_791);
nand U2018 (N_2018,In_693,In_573);
nor U2019 (N_2019,In_694,In_502);
or U2020 (N_2020,In_115,In_761);
nor U2021 (N_2021,In_8,In_51);
or U2022 (N_2022,In_288,In_625);
xnor U2023 (N_2023,In_89,In_223);
or U2024 (N_2024,In_676,In_182);
nand U2025 (N_2025,In_223,In_361);
nand U2026 (N_2026,In_844,In_555);
nand U2027 (N_2027,In_775,In_526);
nor U2028 (N_2028,In_460,In_888);
nor U2029 (N_2029,In_880,In_617);
and U2030 (N_2030,In_399,In_46);
xnor U2031 (N_2031,In_317,In_936);
or U2032 (N_2032,In_796,In_942);
nor U2033 (N_2033,In_304,In_718);
nand U2034 (N_2034,In_897,In_10);
nand U2035 (N_2035,In_930,In_551);
nor U2036 (N_2036,In_524,In_885);
and U2037 (N_2037,In_180,In_857);
and U2038 (N_2038,In_373,In_299);
and U2039 (N_2039,In_400,In_737);
or U2040 (N_2040,In_701,In_291);
nand U2041 (N_2041,In_93,In_605);
nor U2042 (N_2042,In_333,In_157);
nor U2043 (N_2043,In_293,In_460);
or U2044 (N_2044,In_834,In_342);
xnor U2045 (N_2045,In_405,In_78);
xnor U2046 (N_2046,In_330,In_124);
nor U2047 (N_2047,In_260,In_183);
xnor U2048 (N_2048,In_195,In_841);
xnor U2049 (N_2049,In_757,In_173);
nand U2050 (N_2050,In_224,In_195);
xnor U2051 (N_2051,In_785,In_863);
or U2052 (N_2052,In_624,In_207);
xnor U2053 (N_2053,In_76,In_406);
or U2054 (N_2054,In_189,In_788);
nand U2055 (N_2055,In_596,In_97);
xnor U2056 (N_2056,In_722,In_403);
xnor U2057 (N_2057,In_821,In_363);
or U2058 (N_2058,In_451,In_770);
and U2059 (N_2059,In_965,In_884);
or U2060 (N_2060,In_761,In_857);
xor U2061 (N_2061,In_579,In_216);
xnor U2062 (N_2062,In_938,In_201);
nand U2063 (N_2063,In_65,In_889);
nor U2064 (N_2064,In_125,In_92);
nor U2065 (N_2065,In_807,In_206);
nor U2066 (N_2066,In_873,In_660);
xnor U2067 (N_2067,In_925,In_259);
xnor U2068 (N_2068,In_443,In_7);
and U2069 (N_2069,In_211,In_363);
and U2070 (N_2070,In_72,In_682);
and U2071 (N_2071,In_57,In_202);
nor U2072 (N_2072,In_531,In_340);
and U2073 (N_2073,In_645,In_961);
and U2074 (N_2074,In_643,In_804);
and U2075 (N_2075,In_189,In_149);
nor U2076 (N_2076,In_685,In_317);
nor U2077 (N_2077,In_122,In_20);
xnor U2078 (N_2078,In_827,In_30);
nand U2079 (N_2079,In_874,In_780);
xnor U2080 (N_2080,In_75,In_17);
nor U2081 (N_2081,In_403,In_109);
nor U2082 (N_2082,In_155,In_41);
nor U2083 (N_2083,In_429,In_146);
and U2084 (N_2084,In_750,In_827);
or U2085 (N_2085,In_213,In_0);
nand U2086 (N_2086,In_859,In_659);
nand U2087 (N_2087,In_921,In_797);
and U2088 (N_2088,In_130,In_51);
nand U2089 (N_2089,In_565,In_668);
nand U2090 (N_2090,In_874,In_521);
nor U2091 (N_2091,In_814,In_821);
xor U2092 (N_2092,In_605,In_593);
and U2093 (N_2093,In_178,In_864);
or U2094 (N_2094,In_575,In_414);
nor U2095 (N_2095,In_812,In_427);
nor U2096 (N_2096,In_402,In_810);
nor U2097 (N_2097,In_210,In_679);
or U2098 (N_2098,In_550,In_975);
nor U2099 (N_2099,In_534,In_136);
xor U2100 (N_2100,In_999,In_166);
and U2101 (N_2101,In_423,In_315);
xor U2102 (N_2102,In_268,In_698);
and U2103 (N_2103,In_814,In_321);
and U2104 (N_2104,In_851,In_994);
and U2105 (N_2105,In_716,In_906);
or U2106 (N_2106,In_228,In_687);
and U2107 (N_2107,In_65,In_488);
nor U2108 (N_2108,In_149,In_816);
nand U2109 (N_2109,In_341,In_726);
xor U2110 (N_2110,In_952,In_24);
nor U2111 (N_2111,In_346,In_998);
nor U2112 (N_2112,In_107,In_25);
xor U2113 (N_2113,In_436,In_140);
nand U2114 (N_2114,In_311,In_599);
and U2115 (N_2115,In_427,In_96);
nor U2116 (N_2116,In_365,In_711);
nor U2117 (N_2117,In_358,In_882);
xnor U2118 (N_2118,In_653,In_78);
and U2119 (N_2119,In_56,In_633);
xnor U2120 (N_2120,In_196,In_112);
nand U2121 (N_2121,In_275,In_800);
or U2122 (N_2122,In_633,In_629);
xnor U2123 (N_2123,In_634,In_416);
nand U2124 (N_2124,In_117,In_302);
or U2125 (N_2125,In_266,In_476);
nor U2126 (N_2126,In_775,In_746);
nor U2127 (N_2127,In_153,In_432);
nor U2128 (N_2128,In_516,In_70);
or U2129 (N_2129,In_925,In_875);
nor U2130 (N_2130,In_594,In_127);
or U2131 (N_2131,In_722,In_412);
and U2132 (N_2132,In_529,In_203);
xor U2133 (N_2133,In_169,In_479);
nor U2134 (N_2134,In_58,In_782);
xnor U2135 (N_2135,In_812,In_320);
nor U2136 (N_2136,In_979,In_911);
nand U2137 (N_2137,In_586,In_519);
xnor U2138 (N_2138,In_262,In_831);
nor U2139 (N_2139,In_870,In_411);
xor U2140 (N_2140,In_638,In_454);
and U2141 (N_2141,In_21,In_239);
and U2142 (N_2142,In_569,In_822);
and U2143 (N_2143,In_54,In_268);
or U2144 (N_2144,In_677,In_656);
nand U2145 (N_2145,In_294,In_855);
or U2146 (N_2146,In_964,In_272);
and U2147 (N_2147,In_436,In_371);
nand U2148 (N_2148,In_73,In_309);
and U2149 (N_2149,In_567,In_565);
nor U2150 (N_2150,In_414,In_923);
and U2151 (N_2151,In_84,In_253);
and U2152 (N_2152,In_996,In_791);
nor U2153 (N_2153,In_688,In_444);
or U2154 (N_2154,In_457,In_714);
or U2155 (N_2155,In_949,In_41);
nor U2156 (N_2156,In_956,In_621);
or U2157 (N_2157,In_732,In_897);
nor U2158 (N_2158,In_692,In_679);
or U2159 (N_2159,In_437,In_390);
xnor U2160 (N_2160,In_77,In_999);
and U2161 (N_2161,In_688,In_358);
nor U2162 (N_2162,In_788,In_204);
nor U2163 (N_2163,In_196,In_365);
or U2164 (N_2164,In_929,In_138);
nand U2165 (N_2165,In_648,In_606);
nor U2166 (N_2166,In_658,In_265);
nor U2167 (N_2167,In_668,In_421);
nor U2168 (N_2168,In_162,In_527);
or U2169 (N_2169,In_646,In_359);
or U2170 (N_2170,In_106,In_952);
nor U2171 (N_2171,In_72,In_301);
xor U2172 (N_2172,In_481,In_97);
or U2173 (N_2173,In_95,In_841);
and U2174 (N_2174,In_194,In_760);
nor U2175 (N_2175,In_36,In_926);
nand U2176 (N_2176,In_787,In_231);
nand U2177 (N_2177,In_17,In_671);
nor U2178 (N_2178,In_347,In_189);
xnor U2179 (N_2179,In_119,In_871);
nand U2180 (N_2180,In_763,In_678);
xor U2181 (N_2181,In_125,In_668);
and U2182 (N_2182,In_315,In_191);
or U2183 (N_2183,In_381,In_71);
and U2184 (N_2184,In_137,In_627);
nand U2185 (N_2185,In_795,In_40);
nand U2186 (N_2186,In_450,In_708);
or U2187 (N_2187,In_453,In_601);
nand U2188 (N_2188,In_524,In_817);
and U2189 (N_2189,In_393,In_629);
or U2190 (N_2190,In_241,In_236);
nand U2191 (N_2191,In_104,In_73);
and U2192 (N_2192,In_126,In_5);
or U2193 (N_2193,In_669,In_703);
or U2194 (N_2194,In_576,In_94);
or U2195 (N_2195,In_28,In_41);
nand U2196 (N_2196,In_120,In_586);
xor U2197 (N_2197,In_646,In_568);
or U2198 (N_2198,In_574,In_205);
xor U2199 (N_2199,In_987,In_509);
nand U2200 (N_2200,In_818,In_958);
or U2201 (N_2201,In_83,In_851);
nand U2202 (N_2202,In_699,In_609);
xnor U2203 (N_2203,In_34,In_814);
or U2204 (N_2204,In_808,In_180);
nor U2205 (N_2205,In_329,In_222);
xnor U2206 (N_2206,In_313,In_443);
and U2207 (N_2207,In_394,In_542);
or U2208 (N_2208,In_507,In_436);
xnor U2209 (N_2209,In_73,In_138);
nor U2210 (N_2210,In_424,In_157);
or U2211 (N_2211,In_187,In_300);
or U2212 (N_2212,In_609,In_69);
or U2213 (N_2213,In_917,In_15);
xor U2214 (N_2214,In_925,In_994);
xor U2215 (N_2215,In_222,In_673);
or U2216 (N_2216,In_416,In_185);
nor U2217 (N_2217,In_636,In_957);
and U2218 (N_2218,In_181,In_121);
xor U2219 (N_2219,In_366,In_454);
nand U2220 (N_2220,In_312,In_837);
or U2221 (N_2221,In_658,In_771);
and U2222 (N_2222,In_759,In_945);
and U2223 (N_2223,In_816,In_879);
or U2224 (N_2224,In_24,In_129);
and U2225 (N_2225,In_287,In_591);
nor U2226 (N_2226,In_24,In_146);
nor U2227 (N_2227,In_333,In_110);
nand U2228 (N_2228,In_982,In_455);
or U2229 (N_2229,In_263,In_592);
xnor U2230 (N_2230,In_60,In_767);
and U2231 (N_2231,In_313,In_693);
xnor U2232 (N_2232,In_298,In_998);
and U2233 (N_2233,In_933,In_993);
nor U2234 (N_2234,In_762,In_918);
or U2235 (N_2235,In_578,In_603);
xor U2236 (N_2236,In_991,In_786);
and U2237 (N_2237,In_870,In_787);
or U2238 (N_2238,In_710,In_169);
xnor U2239 (N_2239,In_754,In_147);
xnor U2240 (N_2240,In_756,In_763);
and U2241 (N_2241,In_275,In_57);
xnor U2242 (N_2242,In_284,In_475);
or U2243 (N_2243,In_62,In_747);
nor U2244 (N_2244,In_713,In_680);
nor U2245 (N_2245,In_481,In_634);
or U2246 (N_2246,In_372,In_295);
nor U2247 (N_2247,In_604,In_535);
and U2248 (N_2248,In_814,In_35);
xnor U2249 (N_2249,In_999,In_716);
xnor U2250 (N_2250,In_469,In_364);
nand U2251 (N_2251,In_877,In_245);
nor U2252 (N_2252,In_607,In_774);
nand U2253 (N_2253,In_685,In_281);
nor U2254 (N_2254,In_717,In_943);
nor U2255 (N_2255,In_118,In_350);
and U2256 (N_2256,In_944,In_974);
nor U2257 (N_2257,In_941,In_930);
nor U2258 (N_2258,In_825,In_541);
and U2259 (N_2259,In_809,In_736);
xor U2260 (N_2260,In_995,In_643);
xnor U2261 (N_2261,In_308,In_625);
nor U2262 (N_2262,In_386,In_385);
xnor U2263 (N_2263,In_562,In_66);
nand U2264 (N_2264,In_287,In_270);
xnor U2265 (N_2265,In_694,In_28);
and U2266 (N_2266,In_534,In_814);
and U2267 (N_2267,In_822,In_347);
and U2268 (N_2268,In_497,In_41);
nand U2269 (N_2269,In_701,In_159);
nand U2270 (N_2270,In_299,In_598);
nand U2271 (N_2271,In_152,In_809);
nand U2272 (N_2272,In_763,In_800);
nand U2273 (N_2273,In_931,In_65);
or U2274 (N_2274,In_567,In_249);
nor U2275 (N_2275,In_834,In_961);
xor U2276 (N_2276,In_709,In_117);
or U2277 (N_2277,In_616,In_736);
xor U2278 (N_2278,In_338,In_504);
or U2279 (N_2279,In_481,In_536);
and U2280 (N_2280,In_229,In_725);
and U2281 (N_2281,In_795,In_768);
or U2282 (N_2282,In_511,In_690);
or U2283 (N_2283,In_149,In_488);
nand U2284 (N_2284,In_892,In_295);
nor U2285 (N_2285,In_528,In_416);
or U2286 (N_2286,In_177,In_426);
nor U2287 (N_2287,In_996,In_441);
and U2288 (N_2288,In_767,In_67);
xnor U2289 (N_2289,In_42,In_654);
nor U2290 (N_2290,In_669,In_698);
nand U2291 (N_2291,In_408,In_684);
and U2292 (N_2292,In_485,In_477);
and U2293 (N_2293,In_387,In_804);
or U2294 (N_2294,In_859,In_179);
nand U2295 (N_2295,In_4,In_658);
and U2296 (N_2296,In_476,In_375);
nand U2297 (N_2297,In_14,In_120);
nor U2298 (N_2298,In_500,In_550);
and U2299 (N_2299,In_481,In_679);
and U2300 (N_2300,In_879,In_717);
and U2301 (N_2301,In_581,In_713);
nand U2302 (N_2302,In_42,In_21);
and U2303 (N_2303,In_306,In_497);
nand U2304 (N_2304,In_667,In_572);
nand U2305 (N_2305,In_95,In_378);
nand U2306 (N_2306,In_524,In_866);
xor U2307 (N_2307,In_619,In_330);
and U2308 (N_2308,In_696,In_586);
xor U2309 (N_2309,In_726,In_789);
nor U2310 (N_2310,In_564,In_988);
xnor U2311 (N_2311,In_990,In_361);
and U2312 (N_2312,In_641,In_241);
nand U2313 (N_2313,In_25,In_86);
or U2314 (N_2314,In_277,In_901);
nand U2315 (N_2315,In_348,In_936);
nor U2316 (N_2316,In_552,In_744);
or U2317 (N_2317,In_736,In_845);
nor U2318 (N_2318,In_732,In_739);
or U2319 (N_2319,In_678,In_53);
xnor U2320 (N_2320,In_395,In_512);
and U2321 (N_2321,In_649,In_388);
and U2322 (N_2322,In_15,In_373);
and U2323 (N_2323,In_768,In_375);
or U2324 (N_2324,In_587,In_622);
nand U2325 (N_2325,In_489,In_846);
nand U2326 (N_2326,In_11,In_991);
xor U2327 (N_2327,In_499,In_439);
or U2328 (N_2328,In_446,In_420);
or U2329 (N_2329,In_959,In_892);
nand U2330 (N_2330,In_774,In_586);
nor U2331 (N_2331,In_663,In_565);
nor U2332 (N_2332,In_738,In_863);
and U2333 (N_2333,In_869,In_343);
or U2334 (N_2334,In_786,In_798);
and U2335 (N_2335,In_990,In_287);
nand U2336 (N_2336,In_185,In_61);
nor U2337 (N_2337,In_96,In_871);
xnor U2338 (N_2338,In_936,In_603);
xor U2339 (N_2339,In_505,In_720);
and U2340 (N_2340,In_101,In_757);
xor U2341 (N_2341,In_385,In_161);
xnor U2342 (N_2342,In_302,In_914);
xnor U2343 (N_2343,In_996,In_488);
xor U2344 (N_2344,In_81,In_301);
and U2345 (N_2345,In_24,In_5);
and U2346 (N_2346,In_981,In_158);
xnor U2347 (N_2347,In_698,In_399);
xnor U2348 (N_2348,In_883,In_297);
or U2349 (N_2349,In_797,In_677);
nand U2350 (N_2350,In_749,In_626);
xor U2351 (N_2351,In_245,In_579);
nor U2352 (N_2352,In_369,In_371);
nand U2353 (N_2353,In_384,In_983);
nand U2354 (N_2354,In_144,In_931);
or U2355 (N_2355,In_485,In_725);
nor U2356 (N_2356,In_925,In_121);
xor U2357 (N_2357,In_998,In_62);
and U2358 (N_2358,In_27,In_578);
nor U2359 (N_2359,In_118,In_101);
nand U2360 (N_2360,In_652,In_330);
and U2361 (N_2361,In_570,In_467);
or U2362 (N_2362,In_555,In_45);
and U2363 (N_2363,In_812,In_197);
nor U2364 (N_2364,In_910,In_786);
or U2365 (N_2365,In_800,In_496);
and U2366 (N_2366,In_448,In_882);
and U2367 (N_2367,In_109,In_91);
nand U2368 (N_2368,In_551,In_564);
nor U2369 (N_2369,In_919,In_89);
or U2370 (N_2370,In_697,In_682);
or U2371 (N_2371,In_804,In_100);
and U2372 (N_2372,In_836,In_859);
or U2373 (N_2373,In_312,In_226);
or U2374 (N_2374,In_665,In_541);
nand U2375 (N_2375,In_449,In_501);
xor U2376 (N_2376,In_168,In_900);
nand U2377 (N_2377,In_428,In_514);
or U2378 (N_2378,In_793,In_331);
xnor U2379 (N_2379,In_621,In_48);
nor U2380 (N_2380,In_427,In_83);
nor U2381 (N_2381,In_325,In_156);
and U2382 (N_2382,In_527,In_587);
and U2383 (N_2383,In_53,In_757);
nand U2384 (N_2384,In_783,In_71);
nor U2385 (N_2385,In_969,In_116);
nand U2386 (N_2386,In_395,In_150);
nand U2387 (N_2387,In_410,In_290);
nor U2388 (N_2388,In_673,In_69);
nand U2389 (N_2389,In_867,In_36);
or U2390 (N_2390,In_174,In_813);
xnor U2391 (N_2391,In_199,In_40);
and U2392 (N_2392,In_576,In_420);
nand U2393 (N_2393,In_750,In_639);
xor U2394 (N_2394,In_352,In_840);
nand U2395 (N_2395,In_448,In_221);
or U2396 (N_2396,In_312,In_760);
or U2397 (N_2397,In_322,In_386);
xor U2398 (N_2398,In_642,In_65);
xnor U2399 (N_2399,In_949,In_455);
or U2400 (N_2400,In_894,In_178);
nor U2401 (N_2401,In_831,In_477);
nand U2402 (N_2402,In_812,In_916);
or U2403 (N_2403,In_635,In_66);
nor U2404 (N_2404,In_225,In_363);
xor U2405 (N_2405,In_96,In_891);
nor U2406 (N_2406,In_283,In_952);
xnor U2407 (N_2407,In_700,In_732);
nor U2408 (N_2408,In_219,In_719);
or U2409 (N_2409,In_177,In_137);
nand U2410 (N_2410,In_869,In_668);
and U2411 (N_2411,In_3,In_10);
nor U2412 (N_2412,In_611,In_782);
nor U2413 (N_2413,In_836,In_566);
and U2414 (N_2414,In_852,In_18);
or U2415 (N_2415,In_872,In_179);
and U2416 (N_2416,In_92,In_70);
nand U2417 (N_2417,In_196,In_381);
nand U2418 (N_2418,In_702,In_660);
xor U2419 (N_2419,In_510,In_554);
nand U2420 (N_2420,In_531,In_582);
nand U2421 (N_2421,In_313,In_523);
xnor U2422 (N_2422,In_708,In_103);
and U2423 (N_2423,In_88,In_346);
nand U2424 (N_2424,In_847,In_723);
nand U2425 (N_2425,In_396,In_437);
xnor U2426 (N_2426,In_485,In_50);
nand U2427 (N_2427,In_856,In_441);
and U2428 (N_2428,In_547,In_340);
and U2429 (N_2429,In_976,In_819);
xnor U2430 (N_2430,In_102,In_912);
xor U2431 (N_2431,In_975,In_67);
nand U2432 (N_2432,In_832,In_651);
or U2433 (N_2433,In_897,In_56);
xnor U2434 (N_2434,In_250,In_577);
or U2435 (N_2435,In_748,In_195);
xnor U2436 (N_2436,In_791,In_313);
nand U2437 (N_2437,In_537,In_843);
xnor U2438 (N_2438,In_408,In_552);
xnor U2439 (N_2439,In_818,In_15);
and U2440 (N_2440,In_379,In_779);
xnor U2441 (N_2441,In_414,In_368);
nand U2442 (N_2442,In_501,In_335);
and U2443 (N_2443,In_840,In_983);
xnor U2444 (N_2444,In_597,In_513);
xor U2445 (N_2445,In_690,In_69);
or U2446 (N_2446,In_603,In_467);
nor U2447 (N_2447,In_870,In_651);
and U2448 (N_2448,In_815,In_701);
xnor U2449 (N_2449,In_269,In_759);
nor U2450 (N_2450,In_527,In_489);
and U2451 (N_2451,In_112,In_650);
nor U2452 (N_2452,In_155,In_839);
and U2453 (N_2453,In_448,In_265);
or U2454 (N_2454,In_416,In_74);
xor U2455 (N_2455,In_891,In_939);
nand U2456 (N_2456,In_847,In_619);
xnor U2457 (N_2457,In_472,In_617);
nor U2458 (N_2458,In_91,In_703);
nor U2459 (N_2459,In_185,In_872);
or U2460 (N_2460,In_408,In_285);
nand U2461 (N_2461,In_586,In_550);
nor U2462 (N_2462,In_616,In_394);
or U2463 (N_2463,In_612,In_331);
or U2464 (N_2464,In_346,In_996);
nor U2465 (N_2465,In_470,In_396);
and U2466 (N_2466,In_240,In_396);
or U2467 (N_2467,In_228,In_581);
nand U2468 (N_2468,In_931,In_254);
nor U2469 (N_2469,In_48,In_373);
nor U2470 (N_2470,In_113,In_431);
or U2471 (N_2471,In_644,In_906);
nand U2472 (N_2472,In_644,In_563);
and U2473 (N_2473,In_253,In_336);
and U2474 (N_2474,In_720,In_341);
or U2475 (N_2475,In_702,In_440);
nand U2476 (N_2476,In_735,In_369);
nand U2477 (N_2477,In_230,In_542);
nor U2478 (N_2478,In_128,In_312);
nor U2479 (N_2479,In_68,In_706);
nor U2480 (N_2480,In_69,In_821);
and U2481 (N_2481,In_817,In_485);
or U2482 (N_2482,In_342,In_750);
nand U2483 (N_2483,In_249,In_170);
nor U2484 (N_2484,In_443,In_482);
and U2485 (N_2485,In_948,In_723);
nor U2486 (N_2486,In_869,In_250);
nand U2487 (N_2487,In_769,In_29);
xor U2488 (N_2488,In_781,In_342);
nor U2489 (N_2489,In_511,In_785);
nand U2490 (N_2490,In_509,In_776);
xor U2491 (N_2491,In_105,In_851);
and U2492 (N_2492,In_946,In_189);
xnor U2493 (N_2493,In_435,In_866);
or U2494 (N_2494,In_993,In_574);
xnor U2495 (N_2495,In_6,In_372);
xnor U2496 (N_2496,In_382,In_716);
xor U2497 (N_2497,In_421,In_461);
nor U2498 (N_2498,In_416,In_789);
nor U2499 (N_2499,In_524,In_95);
and U2500 (N_2500,N_982,N_973);
nor U2501 (N_2501,N_1719,N_670);
and U2502 (N_2502,N_2224,N_923);
and U2503 (N_2503,N_846,N_854);
and U2504 (N_2504,N_819,N_924);
or U2505 (N_2505,N_68,N_293);
nor U2506 (N_2506,N_2348,N_2210);
or U2507 (N_2507,N_288,N_2225);
and U2508 (N_2508,N_768,N_2311);
and U2509 (N_2509,N_1302,N_1487);
nand U2510 (N_2510,N_1139,N_1718);
or U2511 (N_2511,N_1284,N_1547);
or U2512 (N_2512,N_2250,N_2393);
or U2513 (N_2513,N_2255,N_2291);
nor U2514 (N_2514,N_860,N_180);
nor U2515 (N_2515,N_378,N_993);
or U2516 (N_2516,N_1278,N_2156);
nor U2517 (N_2517,N_1150,N_1168);
nor U2518 (N_2518,N_704,N_2340);
nand U2519 (N_2519,N_1829,N_1409);
nand U2520 (N_2520,N_2419,N_876);
and U2521 (N_2521,N_1592,N_1845);
xnor U2522 (N_2522,N_1596,N_125);
or U2523 (N_2523,N_302,N_2219);
and U2524 (N_2524,N_803,N_1173);
or U2525 (N_2525,N_832,N_2367);
nor U2526 (N_2526,N_1686,N_1821);
nand U2527 (N_2527,N_2397,N_1064);
and U2528 (N_2528,N_201,N_1439);
nor U2529 (N_2529,N_1419,N_216);
and U2530 (N_2530,N_1362,N_2489);
xor U2531 (N_2531,N_1820,N_1051);
and U2532 (N_2532,N_1584,N_1887);
nand U2533 (N_2533,N_1210,N_476);
and U2534 (N_2534,N_245,N_958);
and U2535 (N_2535,N_2478,N_1878);
or U2536 (N_2536,N_667,N_162);
nand U2537 (N_2537,N_1026,N_1776);
xor U2538 (N_2538,N_1262,N_1342);
nor U2539 (N_2539,N_344,N_1532);
nor U2540 (N_2540,N_1629,N_1874);
nand U2541 (N_2541,N_1739,N_2009);
nor U2542 (N_2542,N_2346,N_1812);
and U2543 (N_2543,N_405,N_530);
or U2544 (N_2544,N_1666,N_711);
and U2545 (N_2545,N_959,N_1452);
and U2546 (N_2546,N_985,N_2206);
xnor U2547 (N_2547,N_424,N_601);
or U2548 (N_2548,N_1404,N_2363);
and U2549 (N_2549,N_1918,N_1883);
nand U2550 (N_2550,N_285,N_842);
and U2551 (N_2551,N_273,N_64);
or U2552 (N_2552,N_1661,N_1499);
nand U2553 (N_2553,N_955,N_1091);
or U2554 (N_2554,N_2004,N_2422);
nand U2555 (N_2555,N_886,N_557);
or U2556 (N_2556,N_2099,N_422);
or U2557 (N_2557,N_1917,N_1814);
and U2558 (N_2558,N_412,N_213);
xnor U2559 (N_2559,N_2108,N_1222);
and U2560 (N_2560,N_1065,N_2302);
and U2561 (N_2561,N_487,N_1399);
nor U2562 (N_2562,N_1044,N_2001);
nand U2563 (N_2563,N_631,N_57);
or U2564 (N_2564,N_408,N_1077);
xnor U2565 (N_2565,N_1481,N_231);
and U2566 (N_2566,N_1194,N_2492);
xnor U2567 (N_2567,N_1197,N_239);
and U2568 (N_2568,N_1340,N_2046);
nor U2569 (N_2569,N_2216,N_2034);
nand U2570 (N_2570,N_1742,N_1901);
nand U2571 (N_2571,N_814,N_658);
or U2572 (N_2572,N_1466,N_1250);
xnor U2573 (N_2573,N_222,N_1941);
and U2574 (N_2574,N_544,N_2023);
xor U2575 (N_2575,N_2223,N_1708);
nand U2576 (N_2576,N_1552,N_1743);
and U2577 (N_2577,N_910,N_1273);
nor U2578 (N_2578,N_1684,N_1563);
xnor U2579 (N_2579,N_80,N_18);
or U2580 (N_2580,N_1645,N_2270);
and U2581 (N_2581,N_1354,N_103);
xnor U2582 (N_2582,N_2173,N_2214);
and U2583 (N_2583,N_547,N_1279);
nor U2584 (N_2584,N_1848,N_2349);
xor U2585 (N_2585,N_279,N_1036);
and U2586 (N_2586,N_46,N_1798);
nor U2587 (N_2587,N_1834,N_779);
nand U2588 (N_2588,N_2030,N_1028);
nor U2589 (N_2589,N_1549,N_2081);
nand U2590 (N_2590,N_2027,N_1581);
nand U2591 (N_2591,N_1382,N_514);
nand U2592 (N_2592,N_1530,N_1724);
and U2593 (N_2593,N_582,N_2433);
nor U2594 (N_2594,N_710,N_1327);
nand U2595 (N_2595,N_1430,N_808);
and U2596 (N_2596,N_553,N_2356);
nand U2597 (N_2597,N_2403,N_2065);
and U2598 (N_2598,N_2036,N_903);
nor U2599 (N_2599,N_1653,N_988);
xor U2600 (N_2600,N_2385,N_87);
nor U2601 (N_2601,N_1866,N_787);
or U2602 (N_2602,N_468,N_1121);
nand U2603 (N_2603,N_1215,N_1349);
and U2604 (N_2604,N_828,N_581);
xor U2605 (N_2605,N_995,N_1253);
and U2606 (N_2606,N_869,N_2067);
nand U2607 (N_2607,N_1759,N_1948);
nand U2608 (N_2608,N_98,N_856);
or U2609 (N_2609,N_1945,N_1132);
xnor U2610 (N_2610,N_1185,N_2059);
nand U2611 (N_2611,N_2080,N_1620);
nand U2612 (N_2612,N_2435,N_1939);
or U2613 (N_2613,N_1375,N_1523);
nor U2614 (N_2614,N_2186,N_1300);
xor U2615 (N_2615,N_2353,N_1040);
or U2616 (N_2616,N_2342,N_2215);
nor U2617 (N_2617,N_259,N_784);
nor U2618 (N_2618,N_1078,N_1839);
nor U2619 (N_2619,N_2290,N_480);
nor U2620 (N_2620,N_1591,N_2303);
nor U2621 (N_2621,N_1492,N_1063);
nor U2622 (N_2622,N_1745,N_618);
and U2623 (N_2623,N_587,N_1736);
and U2624 (N_2624,N_861,N_1444);
nor U2625 (N_2625,N_2241,N_884);
nand U2626 (N_2626,N_1183,N_423);
nand U2627 (N_2627,N_983,N_1735);
nor U2628 (N_2628,N_2171,N_1694);
nand U2629 (N_2629,N_574,N_358);
nand U2630 (N_2630,N_392,N_181);
nor U2631 (N_2631,N_502,N_1485);
and U2632 (N_2632,N_2273,N_2107);
nand U2633 (N_2633,N_1593,N_830);
and U2634 (N_2634,N_641,N_1695);
or U2635 (N_2635,N_1384,N_1338);
or U2636 (N_2636,N_615,N_911);
nand U2637 (N_2637,N_622,N_2324);
nand U2638 (N_2638,N_10,N_2076);
nor U2639 (N_2639,N_1956,N_1234);
or U2640 (N_2640,N_1585,N_1154);
nand U2641 (N_2641,N_610,N_25);
nand U2642 (N_2642,N_2304,N_1270);
or U2643 (N_2643,N_2077,N_486);
or U2644 (N_2644,N_383,N_1947);
or U2645 (N_2645,N_588,N_2196);
xnor U2646 (N_2646,N_1934,N_396);
nor U2647 (N_2647,N_338,N_1491);
nor U2648 (N_2648,N_798,N_1892);
or U2649 (N_2649,N_1120,N_2305);
xor U2650 (N_2650,N_345,N_1931);
or U2651 (N_2651,N_2084,N_1321);
or U2652 (N_2652,N_2198,N_60);
nor U2653 (N_2653,N_1606,N_218);
nand U2654 (N_2654,N_1468,N_987);
nor U2655 (N_2655,N_592,N_347);
or U2656 (N_2656,N_159,N_2058);
xor U2657 (N_2657,N_1847,N_74);
xor U2658 (N_2658,N_2280,N_1192);
and U2659 (N_2659,N_141,N_124);
nor U2660 (N_2660,N_1095,N_1923);
nor U2661 (N_2661,N_2070,N_744);
and U2662 (N_2662,N_1318,N_2142);
xnor U2663 (N_2663,N_2380,N_1649);
nand U2664 (N_2664,N_1449,N_1004);
xor U2665 (N_2665,N_752,N_1993);
nand U2666 (N_2666,N_1025,N_470);
and U2667 (N_2667,N_1520,N_1152);
and U2668 (N_2668,N_168,N_908);
xor U2669 (N_2669,N_745,N_805);
nor U2670 (N_2670,N_2037,N_2319);
or U2671 (N_2671,N_1307,N_1978);
nand U2672 (N_2672,N_1637,N_2078);
or U2673 (N_2673,N_106,N_1136);
or U2674 (N_2674,N_1348,N_1752);
nor U2675 (N_2675,N_2443,N_1269);
xnor U2676 (N_2676,N_1674,N_128);
xnor U2677 (N_2677,N_1431,N_2330);
or U2678 (N_2678,N_1971,N_2329);
nand U2679 (N_2679,N_2149,N_278);
and U2680 (N_2680,N_1778,N_1761);
or U2681 (N_2681,N_1018,N_2405);
and U2682 (N_2682,N_203,N_1359);
xor U2683 (N_2683,N_975,N_2098);
or U2684 (N_2684,N_2121,N_1385);
nor U2685 (N_2685,N_1692,N_1545);
or U2686 (N_2686,N_1147,N_611);
nand U2687 (N_2687,N_1495,N_1981);
nand U2688 (N_2688,N_935,N_529);
nand U2689 (N_2689,N_12,N_1073);
and U2690 (N_2690,N_1097,N_685);
nand U2691 (N_2691,N_1083,N_1935);
nand U2692 (N_2692,N_533,N_1779);
or U2693 (N_2693,N_503,N_35);
nor U2694 (N_2694,N_1976,N_393);
nor U2695 (N_2695,N_1140,N_312);
and U2696 (N_2696,N_1067,N_1980);
or U2697 (N_2697,N_1339,N_85);
nor U2698 (N_2698,N_849,N_2274);
xor U2699 (N_2699,N_100,N_1703);
and U2700 (N_2700,N_1762,N_1462);
xor U2701 (N_2701,N_2378,N_1247);
nand U2702 (N_2702,N_646,N_1497);
nor U2703 (N_2703,N_913,N_1212);
or U2704 (N_2704,N_2082,N_2165);
nand U2705 (N_2705,N_1589,N_1391);
nand U2706 (N_2706,N_1070,N_786);
and U2707 (N_2707,N_292,N_1201);
xnor U2708 (N_2708,N_889,N_878);
nor U2709 (N_2709,N_2394,N_402);
and U2710 (N_2710,N_1451,N_840);
and U2711 (N_2711,N_1282,N_621);
or U2712 (N_2712,N_1794,N_1780);
xor U2713 (N_2713,N_991,N_2477);
and U2714 (N_2714,N_1425,N_943);
and U2715 (N_2715,N_1149,N_683);
or U2716 (N_2716,N_1526,N_1472);
and U2717 (N_2717,N_1930,N_1470);
nor U2718 (N_2718,N_1647,N_2170);
and U2719 (N_2719,N_382,N_2155);
and U2720 (N_2720,N_1870,N_2406);
xnor U2721 (N_2721,N_1254,N_2145);
xor U2722 (N_2722,N_1207,N_1218);
nor U2723 (N_2723,N_2494,N_947);
or U2724 (N_2724,N_1330,N_1769);
and U2725 (N_2725,N_1505,N_2334);
or U2726 (N_2726,N_1211,N_1341);
or U2727 (N_2727,N_2337,N_482);
and U2728 (N_2728,N_174,N_1689);
or U2729 (N_2729,N_137,N_1288);
and U2730 (N_2730,N_1543,N_1411);
nor U2731 (N_2731,N_1236,N_2229);
xor U2732 (N_2732,N_864,N_1746);
nor U2733 (N_2733,N_2177,N_770);
xor U2734 (N_2734,N_275,N_1872);
nor U2735 (N_2735,N_411,N_1099);
or U2736 (N_2736,N_1295,N_504);
nor U2737 (N_2737,N_2021,N_1754);
or U2738 (N_2738,N_2128,N_1271);
nor U2739 (N_2739,N_1611,N_780);
or U2740 (N_2740,N_2057,N_569);
nor U2741 (N_2741,N_435,N_1831);
xor U2742 (N_2742,N_283,N_1500);
or U2743 (N_2743,N_2462,N_820);
nand U2744 (N_2744,N_1668,N_1909);
nor U2745 (N_2745,N_909,N_2153);
xnor U2746 (N_2746,N_1888,N_2429);
xor U2747 (N_2747,N_62,N_2201);
xor U2748 (N_2748,N_1021,N_414);
or U2749 (N_2749,N_1628,N_138);
or U2750 (N_2750,N_1170,N_1166);
nor U2751 (N_2751,N_1416,N_308);
or U2752 (N_2752,N_32,N_438);
xor U2753 (N_2753,N_1214,N_1165);
nand U2754 (N_2754,N_1199,N_576);
nand U2755 (N_2755,N_2253,N_1267);
nand U2756 (N_2756,N_2402,N_1962);
nand U2757 (N_2757,N_371,N_1502);
and U2758 (N_2758,N_1846,N_2481);
and U2759 (N_2759,N_1400,N_2460);
nand U2760 (N_2760,N_977,N_2438);
xnor U2761 (N_2761,N_296,N_591);
nor U2762 (N_2762,N_251,N_1937);
xor U2763 (N_2763,N_1347,N_49);
or U2764 (N_2764,N_2442,N_1541);
xnor U2765 (N_2765,N_1929,N_2260);
or U2766 (N_2766,N_204,N_1710);
or U2767 (N_2767,N_206,N_2176);
nor U2768 (N_2768,N_1108,N_782);
and U2769 (N_2769,N_1678,N_894);
and U2770 (N_2770,N_2127,N_2445);
or U2771 (N_2771,N_173,N_1727);
nor U2772 (N_2772,N_1806,N_1960);
nor U2773 (N_2773,N_2482,N_1670);
xor U2774 (N_2774,N_531,N_1730);
nor U2775 (N_2775,N_150,N_627);
and U2776 (N_2776,N_1102,N_2191);
or U2777 (N_2777,N_523,N_580);
nor U2778 (N_2778,N_1413,N_2420);
xor U2779 (N_2779,N_682,N_1777);
xnor U2780 (N_2780,N_449,N_101);
or U2781 (N_2781,N_2415,N_2190);
nand U2782 (N_2782,N_1792,N_342);
nand U2783 (N_2783,N_28,N_2427);
xnor U2784 (N_2784,N_1967,N_243);
and U2785 (N_2785,N_2103,N_295);
or U2786 (N_2786,N_1904,N_1319);
nand U2787 (N_2787,N_1554,N_681);
nand U2788 (N_2788,N_1423,N_326);
nor U2789 (N_2789,N_1702,N_2079);
xnor U2790 (N_2790,N_1949,N_1486);
nand U2791 (N_2791,N_1179,N_1442);
nand U2792 (N_2792,N_1986,N_997);
nand U2793 (N_2793,N_316,N_2400);
or U2794 (N_2794,N_735,N_859);
or U2795 (N_2795,N_756,N_2134);
and U2796 (N_2796,N_1094,N_208);
and U2797 (N_2797,N_30,N_925);
nand U2798 (N_2798,N_2172,N_1357);
or U2799 (N_2799,N_817,N_834);
or U2800 (N_2800,N_2424,N_1117);
or U2801 (N_2801,N_1496,N_1617);
and U2802 (N_2802,N_1813,N_1894);
nor U2803 (N_2803,N_234,N_1196);
nor U2804 (N_2804,N_269,N_823);
and U2805 (N_2805,N_1501,N_1047);
and U2806 (N_2806,N_2275,N_693);
and U2807 (N_2807,N_1298,N_1368);
or U2808 (N_2808,N_471,N_1195);
nand U2809 (N_2809,N_2091,N_540);
and U2810 (N_2810,N_1490,N_1334);
and U2811 (N_2811,N_198,N_792);
nor U2812 (N_2812,N_390,N_1571);
xor U2813 (N_2813,N_2207,N_113);
nand U2814 (N_2814,N_1907,N_1609);
or U2815 (N_2815,N_1729,N_264);
or U2816 (N_2816,N_309,N_2106);
nand U2817 (N_2817,N_2020,N_1310);
nor U2818 (N_2818,N_984,N_282);
nand U2819 (N_2819,N_188,N_75);
and U2820 (N_2820,N_1602,N_45);
xor U2821 (N_2821,N_1809,N_2317);
nand U2822 (N_2822,N_43,N_2094);
or U2823 (N_2823,N_1358,N_1405);
nand U2824 (N_2824,N_539,N_696);
and U2825 (N_2825,N_19,N_205);
or U2826 (N_2826,N_2088,N_1473);
xnor U2827 (N_2827,N_2484,N_2452);
xor U2828 (N_2828,N_289,N_2351);
nand U2829 (N_2829,N_266,N_455);
xor U2830 (N_2830,N_2,N_1054);
nor U2831 (N_2831,N_81,N_845);
xor U2832 (N_2832,N_324,N_2209);
nor U2833 (N_2833,N_1407,N_1240);
or U2834 (N_2834,N_2022,N_72);
and U2835 (N_2835,N_1263,N_1005);
nor U2836 (N_2836,N_2417,N_1660);
xnor U2837 (N_2837,N_1824,N_2265);
nor U2838 (N_2838,N_1910,N_1885);
xnor U2839 (N_2839,N_2310,N_1968);
or U2840 (N_2840,N_1424,N_701);
nand U2841 (N_2841,N_1876,N_1420);
nand U2842 (N_2842,N_1445,N_1011);
nand U2843 (N_2843,N_769,N_837);
nor U2844 (N_2844,N_1182,N_1950);
or U2845 (N_2845,N_413,N_636);
and U2846 (N_2846,N_2217,N_1903);
xnor U2847 (N_2847,N_2294,N_1112);
nand U2848 (N_2848,N_1533,N_738);
xor U2849 (N_2849,N_2343,N_1280);
nor U2850 (N_2850,N_1050,N_156);
or U2851 (N_2851,N_1386,N_2289);
nand U2852 (N_2852,N_1027,N_1482);
nor U2853 (N_2853,N_1257,N_1364);
or U2854 (N_2854,N_310,N_560);
and U2855 (N_2855,N_931,N_1772);
and U2856 (N_2856,N_1817,N_1721);
or U2857 (N_2857,N_2408,N_2257);
xor U2858 (N_2858,N_1638,N_1744);
or U2859 (N_2859,N_432,N_1972);
or U2860 (N_2860,N_488,N_2109);
xnor U2861 (N_2861,N_672,N_479);
xor U2862 (N_2862,N_585,N_418);
or U2863 (N_2863,N_1291,N_2008);
nand U2864 (N_2864,N_885,N_771);
nor U2865 (N_2865,N_1896,N_518);
or U2866 (N_2866,N_1305,N_599);
or U2867 (N_2867,N_370,N_1356);
nand U2868 (N_2868,N_1900,N_96);
and U2869 (N_2869,N_2017,N_299);
nand U2870 (N_2870,N_1914,N_1110);
or U2871 (N_2871,N_1880,N_2032);
xor U2872 (N_2872,N_905,N_73);
nand U2873 (N_2873,N_2398,N_620);
and U2874 (N_2874,N_1636,N_1317);
nand U2875 (N_2875,N_195,N_2062);
and U2876 (N_2876,N_2167,N_104);
or U2877 (N_2877,N_388,N_721);
nor U2878 (N_2878,N_2071,N_831);
xnor U2879 (N_2879,N_1161,N_298);
nand U2880 (N_2880,N_240,N_2249);
or U2881 (N_2881,N_202,N_1374);
nor U2882 (N_2882,N_20,N_565);
nor U2883 (N_2883,N_743,N_1000);
and U2884 (N_2884,N_110,N_2464);
or U2885 (N_2885,N_1863,N_841);
xnor U2886 (N_2886,N_536,N_1861);
nor U2887 (N_2887,N_1088,N_178);
or U2888 (N_2888,N_1174,N_1773);
nor U2889 (N_2889,N_1494,N_1457);
and U2890 (N_2890,N_873,N_349);
or U2891 (N_2891,N_1017,N_879);
xnor U2892 (N_2892,N_1961,N_687);
or U2893 (N_2893,N_791,N_1177);
nor U2894 (N_2894,N_848,N_598);
nor U2895 (N_2895,N_2471,N_1134);
xor U2896 (N_2896,N_556,N_495);
nand U2897 (N_2897,N_1373,N_2479);
nor U2898 (N_2898,N_1432,N_1020);
or U2899 (N_2899,N_1558,N_739);
nand U2900 (N_2900,N_1474,N_2000);
xor U2901 (N_2901,N_1749,N_2193);
or U2902 (N_2902,N_507,N_2288);
nor U2903 (N_2903,N_1332,N_1285);
or U2904 (N_2904,N_2212,N_2320);
nor U2905 (N_2905,N_510,N_2323);
nor U2906 (N_2906,N_447,N_1632);
or U2907 (N_2907,N_2028,N_800);
nor U2908 (N_2908,N_1815,N_545);
and U2909 (N_2909,N_380,N_1768);
xnor U2910 (N_2910,N_996,N_1066);
nand U2911 (N_2911,N_1408,N_1869);
xor U2912 (N_2912,N_790,N_90);
nor U2913 (N_2913,N_774,N_2095);
nand U2914 (N_2914,N_331,N_1517);
xor U2915 (N_2915,N_2025,N_132);
nor U2916 (N_2916,N_2432,N_2235);
or U2917 (N_2917,N_2497,N_645);
nand U2918 (N_2918,N_753,N_961);
xnor U2919 (N_2919,N_1631,N_538);
or U2920 (N_2920,N_1458,N_1042);
nand U2921 (N_2921,N_1297,N_136);
xnor U2922 (N_2922,N_709,N_1920);
nor U2923 (N_2923,N_1426,N_2299);
nand U2924 (N_2924,N_1220,N_1979);
xor U2925 (N_2925,N_1700,N_1855);
nand U2926 (N_2926,N_1213,N_2019);
xnor U2927 (N_2927,N_850,N_1277);
nor U2928 (N_2928,N_664,N_77);
xor U2929 (N_2929,N_515,N_1884);
xnor U2930 (N_2930,N_29,N_82);
nand U2931 (N_2931,N_2033,N_1440);
or U2932 (N_2932,N_1072,N_163);
and U2933 (N_2933,N_472,N_1613);
and U2934 (N_2934,N_1033,N_656);
xnor U2935 (N_2935,N_433,N_732);
or U2936 (N_2936,N_967,N_2383);
and U2937 (N_2937,N_2463,N_2117);
nor U2938 (N_2938,N_1394,N_1323);
xor U2939 (N_2939,N_2388,N_1512);
and U2940 (N_2940,N_2096,N_1728);
or U2941 (N_2941,N_362,N_1463);
or U2942 (N_2942,N_403,N_1441);
xor U2943 (N_2943,N_1844,N_917);
xor U2944 (N_2944,N_969,N_51);
xor U2945 (N_2945,N_1264,N_2024);
nor U2946 (N_2946,N_2203,N_384);
nor U2947 (N_2947,N_2202,N_66);
or U2948 (N_2948,N_1239,N_1219);
and U2949 (N_2949,N_1864,N_86);
or U2950 (N_2950,N_1524,N_2087);
or U2951 (N_2951,N_1315,N_1178);
xor U2952 (N_2952,N_1757,N_577);
nor U2953 (N_2953,N_17,N_920);
nor U2954 (N_2954,N_1306,N_149);
and U2955 (N_2955,N_437,N_1790);
nand U2956 (N_2956,N_15,N_1938);
or U2957 (N_2957,N_61,N_2188);
and U2958 (N_2958,N_1796,N_2011);
and U2959 (N_2959,N_968,N_1115);
nor U2960 (N_2960,N_1521,N_58);
or U2961 (N_2961,N_123,N_356);
nand U2962 (N_2962,N_327,N_963);
xor U2963 (N_2963,N_2245,N_166);
nand U2964 (N_2964,N_1974,N_2016);
nor U2965 (N_2965,N_2184,N_169);
or U2966 (N_2966,N_1651,N_56);
and U2967 (N_2967,N_214,N_254);
xnor U2968 (N_2968,N_579,N_1260);
or U2969 (N_2969,N_1576,N_1557);
xor U2970 (N_2970,N_706,N_2258);
nor U2971 (N_2971,N_2179,N_1417);
nand U2972 (N_2972,N_1807,N_1553);
or U2973 (N_2973,N_941,N_1418);
xor U2974 (N_2974,N_1387,N_1311);
and U2975 (N_2975,N_882,N_895);
nand U2976 (N_2976,N_720,N_33);
or U2977 (N_2977,N_2136,N_2227);
xor U2978 (N_2978,N_140,N_2355);
xnor U2979 (N_2979,N_586,N_614);
xor U2980 (N_2980,N_1741,N_1770);
and U2981 (N_2981,N_1325,N_130);
nand U2982 (N_2982,N_41,N_2230);
nand U2983 (N_2983,N_1610,N_767);
xnor U2984 (N_2984,N_1249,N_899);
or U2985 (N_2985,N_2376,N_478);
or U2986 (N_2986,N_318,N_50);
nand U2987 (N_2987,N_2072,N_1231);
xor U2988 (N_2988,N_2371,N_443);
xnor U2989 (N_2989,N_1126,N_1588);
xnor U2990 (N_2990,N_1160,N_8);
nand U2991 (N_2991,N_303,N_276);
xor U2992 (N_2992,N_2174,N_1826);
nor U2993 (N_2993,N_1598,N_1226);
nand U2994 (N_2994,N_1453,N_1975);
or U2995 (N_2995,N_1955,N_2013);
or U2996 (N_2996,N_1621,N_1525);
nor U2997 (N_2997,N_212,N_762);
and U2998 (N_2998,N_1990,N_2461);
nor U2999 (N_2999,N_1329,N_2105);
nor U3000 (N_3000,N_1723,N_1352);
or U3001 (N_3001,N_1819,N_1756);
and U3002 (N_3002,N_684,N_2097);
nor U3003 (N_3003,N_1052,N_1936);
nor U3004 (N_3004,N_604,N_1331);
or U3005 (N_3005,N_1654,N_1566);
nand U3006 (N_3006,N_2104,N_2358);
nand U3007 (N_3007,N_332,N_1912);
or U3008 (N_3008,N_906,N_902);
xor U3009 (N_3009,N_2469,N_48);
nand U3010 (N_3010,N_1682,N_1345);
and U3011 (N_3011,N_2029,N_660);
or U3012 (N_3012,N_623,N_2456);
or U3013 (N_3013,N_1528,N_2026);
nor U3014 (N_3014,N_97,N_2401);
and U3015 (N_3015,N_1590,N_272);
and U3016 (N_3016,N_458,N_1751);
or U3017 (N_3017,N_2467,N_232);
nor U3018 (N_3018,N_1053,N_228);
nand U3019 (N_3019,N_524,N_1268);
nand U3020 (N_3020,N_1802,N_2437);
nor U3021 (N_3021,N_603,N_1350);
and U3022 (N_3022,N_705,N_2159);
and U3023 (N_3023,N_255,N_764);
xor U3024 (N_3024,N_367,N_1252);
nand U3025 (N_3025,N_2440,N_427);
nand U3026 (N_3026,N_1858,N_1607);
or U3027 (N_3027,N_253,N_1248);
and U3028 (N_3028,N_2352,N_929);
nor U3029 (N_3029,N_1952,N_669);
or U3030 (N_3030,N_152,N_446);
xnor U3031 (N_3031,N_334,N_1080);
nor U3032 (N_3032,N_750,N_1146);
or U3033 (N_3033,N_2269,N_1414);
nor U3034 (N_3034,N_2493,N_401);
and U3035 (N_3035,N_813,N_2093);
nor U3036 (N_3036,N_2446,N_2333);
nand U3037 (N_3037,N_1141,N_2436);
nor U3038 (N_3038,N_1232,N_690);
xor U3039 (N_3039,N_2266,N_835);
xnor U3040 (N_3040,N_1003,N_1478);
xor U3041 (N_3041,N_450,N_1580);
xor U3042 (N_3042,N_67,N_1618);
and U3043 (N_3043,N_933,N_1477);
nand U3044 (N_3044,N_2354,N_111);
nor U3045 (N_3045,N_191,N_862);
nor U3046 (N_3046,N_724,N_1604);
nor U3047 (N_3047,N_2189,N_160);
and U3048 (N_3048,N_1789,N_2277);
and U3049 (N_3049,N_2130,N_385);
or U3050 (N_3050,N_102,N_1369);
nor U3051 (N_3051,N_439,N_1856);
xnor U3052 (N_3052,N_506,N_237);
and U3053 (N_3053,N_1039,N_336);
xnor U3054 (N_3054,N_807,N_1434);
and U3055 (N_3055,N_1410,N_1225);
nand U3056 (N_3056,N_824,N_1206);
and U3057 (N_3057,N_148,N_1626);
and U3058 (N_3058,N_668,N_1919);
xor U3059 (N_3059,N_516,N_1828);
nor U3060 (N_3060,N_265,N_333);
nor U3061 (N_3061,N_2180,N_2232);
xor U3062 (N_3062,N_1514,N_1717);
and U3063 (N_3063,N_1469,N_2138);
or U3064 (N_3064,N_794,N_689);
and U3065 (N_3065,N_1246,N_1337);
nand U3066 (N_3066,N_270,N_896);
nand U3067 (N_3067,N_1940,N_1476);
nand U3068 (N_3068,N_1172,N_281);
nand U3069 (N_3069,N_1098,N_2123);
nor U3070 (N_3070,N_1467,N_2090);
nand U3071 (N_3071,N_880,N_1679);
and U3072 (N_3072,N_1111,N_2444);
nand U3073 (N_3073,N_733,N_575);
and U3074 (N_3074,N_1933,N_1062);
xnor U3075 (N_3075,N_360,N_2339);
nand U3076 (N_3076,N_654,N_227);
nand U3077 (N_3077,N_1289,N_1958);
xor U3078 (N_3078,N_425,N_772);
nor U3079 (N_3079,N_236,N_2267);
and U3080 (N_3080,N_1133,N_94);
xnor U3081 (N_3081,N_165,N_319);
nand U3082 (N_3082,N_186,N_2459);
xor U3083 (N_3083,N_6,N_230);
nand U3084 (N_3084,N_1748,N_99);
nand U3085 (N_3085,N_1301,N_277);
and U3086 (N_3086,N_26,N_2296);
nor U3087 (N_3087,N_286,N_1326);
nor U3088 (N_3088,N_2491,N_2005);
and U3089 (N_3089,N_1393,N_1797);
and U3090 (N_3090,N_2499,N_589);
xnor U3091 (N_3091,N_346,N_948);
nand U3092 (N_3092,N_1565,N_426);
or U3093 (N_3093,N_389,N_2345);
nand U3094 (N_3094,N_2178,N_2231);
and U3095 (N_3095,N_1634,N_2146);
xor U3096 (N_3096,N_1276,N_725);
or U3097 (N_3097,N_1084,N_1119);
nor U3098 (N_3098,N_1693,N_1163);
and U3099 (N_3099,N_1957,N_1635);
nand U3100 (N_3100,N_2238,N_262);
and U3101 (N_3101,N_673,N_1022);
and U3102 (N_3102,N_1493,N_1652);
xnor U3103 (N_3103,N_1100,N_688);
xor U3104 (N_3104,N_562,N_167);
nand U3105 (N_3105,N_2018,N_1989);
and U3106 (N_3106,N_554,N_335);
xnor U3107 (N_3107,N_2006,N_1437);
xnor U3108 (N_3108,N_747,N_1737);
xor U3109 (N_3109,N_409,N_2047);
or U3110 (N_3110,N_215,N_107);
nor U3111 (N_3111,N_1535,N_2426);
or U3112 (N_3112,N_2069,N_494);
or U3113 (N_3113,N_1805,N_1573);
nor U3114 (N_3114,N_322,N_1456);
nand U3115 (N_3115,N_261,N_1488);
or U3116 (N_3116,N_1529,N_2295);
and U3117 (N_3117,N_1304,N_1622);
xnor U3118 (N_3118,N_887,N_444);
nor U3119 (N_3119,N_1616,N_2472);
nor U3120 (N_3120,N_535,N_1908);
and U3121 (N_3121,N_1037,N_157);
xor U3122 (N_3122,N_2066,N_484);
and U3123 (N_3123,N_1964,N_1765);
or U3124 (N_3124,N_2244,N_2074);
and U3125 (N_3125,N_1842,N_1605);
nor U3126 (N_3126,N_337,N_2423);
nand U3127 (N_3127,N_2197,N_1363);
xnor U3128 (N_3128,N_135,N_1687);
xor U3129 (N_3129,N_2053,N_1461);
and U3130 (N_3130,N_2132,N_2369);
xnor U3131 (N_3131,N_1074,N_224);
xnor U3132 (N_3132,N_1123,N_1881);
or U3133 (N_3133,N_1895,N_399);
and U3134 (N_3134,N_1379,N_1024);
and U3135 (N_3135,N_763,N_69);
nor U3136 (N_3136,N_2042,N_93);
and U3137 (N_3137,N_2218,N_115);
xor U3138 (N_3138,N_1542,N_1564);
xnor U3139 (N_3139,N_1446,N_2344);
and U3140 (N_3140,N_919,N_519);
nand U3141 (N_3141,N_257,N_1186);
or U3142 (N_3142,N_785,N_799);
or U3143 (N_3143,N_1658,N_146);
nor U3144 (N_3144,N_1447,N_2116);
and U3145 (N_3145,N_456,N_2125);
or U3146 (N_3146,N_1312,N_1244);
and U3147 (N_3147,N_1046,N_1720);
xor U3148 (N_3148,N_914,N_1791);
xor U3149 (N_3149,N_2364,N_1832);
nand U3150 (N_3150,N_252,N_1010);
xor U3151 (N_3151,N_1992,N_1175);
xor U3152 (N_3152,N_1109,N_893);
or U3153 (N_3153,N_176,N_981);
nor U3154 (N_3154,N_1125,N_827);
xor U3155 (N_3155,N_315,N_729);
nor U3156 (N_3156,N_694,N_713);
and U3157 (N_3157,N_294,N_1650);
and U3158 (N_3158,N_1559,N_777);
nor U3159 (N_3159,N_91,N_407);
xnor U3160 (N_3160,N_2236,N_1403);
nand U3161 (N_3161,N_1714,N_2439);
nor U3162 (N_3162,N_1680,N_14);
and U3163 (N_3163,N_2297,N_1838);
or U3164 (N_3164,N_1551,N_151);
or U3165 (N_3165,N_1657,N_2455);
nand U3166 (N_3166,N_398,N_1711);
nand U3167 (N_3167,N_436,N_945);
or U3168 (N_3168,N_1675,N_2233);
or U3169 (N_3169,N_1619,N_825);
or U3170 (N_3170,N_1167,N_1999);
or U3171 (N_3171,N_2396,N_716);
xor U3172 (N_3172,N_1672,N_1854);
nand U3173 (N_3173,N_730,N_1498);
or U3174 (N_3174,N_1019,N_121);
nor U3175 (N_3175,N_70,N_182);
xor U3176 (N_3176,N_223,N_609);
and U3177 (N_3177,N_868,N_1454);
nand U3178 (N_3178,N_874,N_534);
and U3179 (N_3179,N_1664,N_1709);
nor U3180 (N_3180,N_1138,N_194);
nor U3181 (N_3181,N_1561,N_129);
or U3182 (N_3182,N_1816,N_2453);
or U3183 (N_3183,N_915,N_740);
nor U3184 (N_3184,N_1238,N_932);
nor U3185 (N_3185,N_189,N_2040);
nand U3186 (N_3186,N_2060,N_2390);
nand U3187 (N_3187,N_2157,N_665);
nand U3188 (N_3188,N_1153,N_1055);
and U3189 (N_3189,N_2281,N_2391);
and U3190 (N_3190,N_248,N_2411);
nor U3191 (N_3191,N_498,N_133);
nand U3192 (N_3192,N_726,N_1243);
xor U3193 (N_3193,N_1471,N_1292);
nor U3194 (N_3194,N_2089,N_1731);
nor U3195 (N_3195,N_473,N_1370);
nor U3196 (N_3196,N_590,N_2122);
or U3197 (N_3197,N_271,N_1366);
nor U3198 (N_3198,N_467,N_306);
nor U3199 (N_3199,N_2002,N_2200);
xnor U3200 (N_3200,N_934,N_907);
or U3201 (N_3201,N_1642,N_235);
xor U3202 (N_3202,N_2341,N_260);
xnor U3203 (N_3203,N_1023,N_2237);
nor U3204 (N_3204,N_1582,N_815);
xnor U3205 (N_3205,N_1436,N_1915);
nand U3206 (N_3206,N_1706,N_79);
and U3207 (N_3207,N_1313,N_2470);
nor U3208 (N_3208,N_1090,N_2316);
or U3209 (N_3209,N_2395,N_1516);
and U3210 (N_3210,N_1823,N_2362);
or U3211 (N_3211,N_2049,N_1793);
xor U3212 (N_3212,N_1732,N_1314);
nand U3213 (N_3213,N_2496,N_1515);
and U3214 (N_3214,N_1480,N_541);
and U3215 (N_3215,N_937,N_1145);
nor U3216 (N_3216,N_1261,N_2007);
and U3217 (N_3217,N_2286,N_225);
nor U3218 (N_3218,N_354,N_5);
and U3219 (N_3219,N_826,N_812);
nand U3220 (N_3220,N_966,N_699);
or U3221 (N_3221,N_2300,N_863);
nor U3222 (N_3222,N_329,N_1716);
and U3223 (N_3223,N_131,N_2414);
and U3224 (N_3224,N_1274,N_47);
and U3225 (N_3225,N_290,N_2366);
xor U3226 (N_3226,N_1045,N_2050);
nor U3227 (N_3227,N_1612,N_1928);
nor U3228 (N_3228,N_715,N_89);
or U3229 (N_3229,N_666,N_978);
nor U3230 (N_3230,N_1506,N_606);
or U3231 (N_3231,N_1540,N_2264);
nor U3232 (N_3232,N_663,N_972);
and U3233 (N_3233,N_1587,N_629);
nor U3234 (N_3234,N_1873,N_571);
nand U3235 (N_3235,N_851,N_1600);
or U3236 (N_3236,N_1963,N_1891);
or U3237 (N_3237,N_220,N_561);
nor U3238 (N_3238,N_638,N_707);
nand U3239 (N_3239,N_1283,N_1367);
nand U3240 (N_3240,N_2465,N_1371);
xor U3241 (N_3241,N_1324,N_1184);
nor U3242 (N_3242,N_1550,N_691);
nand U3243 (N_3243,N_2483,N_676);
nand U3244 (N_3244,N_776,N_1868);
and U3245 (N_3245,N_2137,N_221);
or U3246 (N_3246,N_1667,N_513);
and U3247 (N_3247,N_2321,N_1129);
nand U3248 (N_3248,N_2382,N_2309);
xor U3249 (N_3249,N_1851,N_1401);
or U3250 (N_3250,N_451,N_280);
xnor U3251 (N_3251,N_1849,N_1061);
xnor U3252 (N_3252,N_1171,N_2262);
and U3253 (N_3253,N_83,N_2327);
and U3254 (N_3254,N_2228,N_965);
nand U3255 (N_3255,N_686,N_718);
and U3256 (N_3256,N_1007,N_695);
nor U3257 (N_3257,N_430,N_793);
xnor U3258 (N_3258,N_644,N_1322);
xnor U3259 (N_3259,N_1775,N_737);
nand U3260 (N_3260,N_496,N_1412);
nor U3261 (N_3261,N_179,N_567);
nor U3262 (N_3262,N_1548,N_760);
nand U3263 (N_3263,N_875,N_918);
nor U3264 (N_3264,N_844,N_52);
xnor U3265 (N_3265,N_505,N_512);
nand U3266 (N_3266,N_734,N_651);
xnor U3267 (N_3267,N_1015,N_613);
nor U3268 (N_3268,N_352,N_1227);
nor U3269 (N_3269,N_2211,N_247);
xnor U3270 (N_3270,N_778,N_199);
nor U3271 (N_3271,N_2487,N_1715);
nor U3272 (N_3272,N_145,N_1504);
xor U3273 (N_3273,N_1784,N_192);
and U3274 (N_3274,N_1395,N_2115);
or U3275 (N_3275,N_2268,N_1713);
xnor U3276 (N_3276,N_2256,N_364);
nor U3277 (N_3277,N_2221,N_381);
nor U3278 (N_3278,N_2162,N_804);
nand U3279 (N_3279,N_2075,N_674);
xor U3280 (N_3280,N_1767,N_2185);
nor U3281 (N_3281,N_2263,N_1987);
nor U3282 (N_3282,N_796,N_1641);
nand U3283 (N_3283,N_2441,N_0);
xor U3284 (N_3284,N_1118,N_183);
nor U3285 (N_3285,N_1503,N_766);
xor U3286 (N_3286,N_1537,N_749);
nor U3287 (N_3287,N_2301,N_2466);
or U3288 (N_3288,N_369,N_2490);
nor U3289 (N_3289,N_209,N_1006);
xnor U3290 (N_3290,N_477,N_1640);
nand U3291 (N_3291,N_986,N_2039);
and U3292 (N_3292,N_499,N_1902);
or U3293 (N_3293,N_2251,N_1205);
nand U3294 (N_3294,N_1169,N_1190);
xor U3295 (N_3295,N_619,N_1843);
or U3296 (N_3296,N_1,N_1082);
nor U3297 (N_3297,N_2335,N_1209);
or U3298 (N_3298,N_2118,N_1187);
nor U3299 (N_3299,N_942,N_926);
nor U3300 (N_3300,N_142,N_1673);
nor U3301 (N_3301,N_980,N_184);
nand U3302 (N_3302,N_1351,N_2350);
and U3303 (N_3303,N_550,N_1508);
nand U3304 (N_3304,N_2293,N_821);
nand U3305 (N_3305,N_1995,N_1105);
or U3306 (N_3306,N_419,N_960);
and U3307 (N_3307,N_2163,N_1202);
or U3308 (N_3308,N_1361,N_2252);
and U3309 (N_3309,N_491,N_1833);
and U3310 (N_3310,N_490,N_1519);
and U3311 (N_3311,N_1421,N_434);
nand U3312 (N_3312,N_361,N_1959);
and U3313 (N_3313,N_2292,N_2166);
and U3314 (N_3314,N_114,N_1122);
nand U3315 (N_3315,N_1886,N_117);
or U3316 (N_3316,N_2447,N_1705);
xnor U3317 (N_3317,N_1290,N_440);
and U3318 (N_3318,N_2486,N_679);
or U3319 (N_3319,N_1586,N_653);
xnor U3320 (N_3320,N_1624,N_1882);
nand U3321 (N_3321,N_1556,N_1683);
nand U3322 (N_3322,N_1946,N_1627);
and U3323 (N_3323,N_998,N_1085);
xnor U3324 (N_3324,N_2377,N_1343);
or U3325 (N_3325,N_1799,N_1155);
nor U3326 (N_3326,N_1124,N_649);
nor U3327 (N_3327,N_1603,N_2404);
nand U3328 (N_3328,N_1795,N_754);
nor U3329 (N_3329,N_936,N_809);
xnor U3330 (N_3330,N_2152,N_320);
xor U3331 (N_3331,N_2208,N_602);
nor U3332 (N_3332,N_532,N_2416);
or U3333 (N_3333,N_2322,N_703);
and U3334 (N_3334,N_1460,N_27);
nor U3335 (N_3335,N_1544,N_1860);
xor U3336 (N_3336,N_421,N_2370);
or U3337 (N_3337,N_748,N_1942);
nor U3338 (N_3338,N_552,N_24);
xnor U3339 (N_3339,N_1726,N_2083);
nand U3340 (N_3340,N_1002,N_775);
or U3341 (N_3341,N_872,N_200);
nor U3342 (N_3342,N_2048,N_368);
nand U3343 (N_3343,N_1639,N_357);
nand U3344 (N_3344,N_454,N_1804);
or U3345 (N_3345,N_2012,N_373);
and U3346 (N_3346,N_2234,N_2325);
or U3347 (N_3347,N_1738,N_989);
nor U3348 (N_3348,N_1659,N_1841);
and U3349 (N_3349,N_1998,N_1048);
xnor U3350 (N_3350,N_1309,N_143);
nand U3351 (N_3351,N_921,N_938);
or U3352 (N_3352,N_1595,N_979);
xor U3353 (N_3353,N_109,N_727);
xor U3354 (N_3354,N_1608,N_2110);
or U3355 (N_3355,N_642,N_1648);
nand U3356 (N_3356,N_2410,N_417);
xor U3357 (N_3357,N_2328,N_992);
or U3358 (N_3358,N_2141,N_1058);
xnor U3359 (N_3359,N_1701,N_2164);
and U3360 (N_3360,N_951,N_953);
and U3361 (N_3361,N_464,N_1181);
or U3362 (N_3362,N_1835,N_1272);
and U3363 (N_3363,N_1725,N_343);
and U3364 (N_3364,N_2374,N_1293);
nand U3365 (N_3365,N_1377,N_153);
or U3366 (N_3366,N_1286,N_452);
xnor U3367 (N_3367,N_526,N_2051);
xnor U3368 (N_3368,N_2379,N_677);
and U3369 (N_3369,N_1255,N_172);
or U3370 (N_3370,N_258,N_1996);
or U3371 (N_3371,N_806,N_1867);
and U3372 (N_3372,N_463,N_2331);
xor U3373 (N_3373,N_1857,N_154);
nor U3374 (N_3374,N_836,N_1381);
xor U3375 (N_3375,N_2120,N_922);
or U3376 (N_3376,N_287,N_1256);
nand U3377 (N_3377,N_2458,N_1579);
and U3378 (N_3378,N_1951,N_1555);
nor U3379 (N_3379,N_866,N_1113);
and U3380 (N_3380,N_829,N_1875);
nand U3381 (N_3381,N_1335,N_839);
xnor U3382 (N_3382,N_1685,N_2112);
and U3383 (N_3383,N_1266,N_3);
xnor U3384 (N_3384,N_789,N_1148);
and U3385 (N_3385,N_1489,N_2148);
nand U3386 (N_3386,N_1583,N_2154);
nand U3387 (N_3387,N_1696,N_2041);
nand U3388 (N_3388,N_643,N_2035);
xor U3389 (N_3389,N_1699,N_1840);
nor U3390 (N_3390,N_95,N_1057);
nand U3391 (N_3391,N_892,N_1223);
or U3392 (N_3392,N_1698,N_323);
and U3393 (N_3393,N_460,N_1800);
xor U3394 (N_3394,N_1994,N_1188);
and U3395 (N_3395,N_612,N_1750);
nand U3396 (N_3396,N_40,N_219);
and U3397 (N_3397,N_1060,N_1911);
or U3398 (N_3398,N_406,N_1013);
and U3399 (N_3399,N_898,N_1983);
nand U3400 (N_3400,N_1104,N_2407);
or U3401 (N_3401,N_1056,N_375);
nor U3402 (N_3402,N_1862,N_2308);
nand U3403 (N_3403,N_1422,N_1825);
xor U3404 (N_3404,N_650,N_1151);
nand U3405 (N_3405,N_2204,N_416);
nand U3406 (N_3406,N_1221,N_2449);
nor U3407 (N_3407,N_1303,N_122);
nor U3408 (N_3408,N_1296,N_267);
and U3409 (N_3409,N_2054,N_697);
or U3410 (N_3410,N_492,N_2044);
and U3411 (N_3411,N_2287,N_481);
xor U3412 (N_3412,N_410,N_2038);
or U3413 (N_3413,N_1671,N_2399);
xnor U3414 (N_3414,N_1574,N_1159);
or U3415 (N_3415,N_2213,N_147);
xnor U3416 (N_3416,N_572,N_1803);
and U3417 (N_3417,N_1527,N_317);
nor U3418 (N_3418,N_1890,N_597);
or U3419 (N_3419,N_1755,N_2114);
nand U3420 (N_3420,N_648,N_1443);
or U3421 (N_3421,N_465,N_1320);
xnor U3422 (N_3422,N_1038,N_1546);
and U3423 (N_3423,N_640,N_1143);
nor U3424 (N_3424,N_1235,N_2064);
and U3425 (N_3425,N_340,N_36);
or U3426 (N_3426,N_781,N_217);
nand U3427 (N_3427,N_1899,N_177);
nand U3428 (N_3428,N_702,N_1130);
and U3429 (N_3429,N_2135,N_962);
nand U3430 (N_3430,N_1509,N_717);
xor U3431 (N_3431,N_657,N_2158);
nor U3432 (N_3432,N_256,N_628);
or U3433 (N_3433,N_1953,N_448);
nand U3434 (N_3434,N_1785,N_626);
nand U3435 (N_3435,N_2387,N_78);
nor U3436 (N_3436,N_2318,N_185);
or U3437 (N_3437,N_250,N_2315);
or U3438 (N_3438,N_1984,N_119);
nand U3439 (N_3439,N_474,N_2312);
nor U3440 (N_3440,N_2085,N_1032);
or U3441 (N_3441,N_847,N_927);
xor U3442 (N_3442,N_1753,N_1200);
xnor U3443 (N_3443,N_1747,N_1216);
and U3444 (N_3444,N_2119,N_2347);
xnor U3445 (N_3445,N_542,N_1435);
nand U3446 (N_3446,N_916,N_2052);
and U3447 (N_3447,N_2043,N_551);
or U3448 (N_3448,N_1853,N_700);
xor U3449 (N_3449,N_990,N_853);
and U3450 (N_3450,N_2475,N_2063);
xor U3451 (N_3451,N_956,N_431);
nor U3452 (N_3452,N_1224,N_9);
xor U3453 (N_3453,N_1764,N_394);
nor U3454 (N_3454,N_374,N_1808);
and U3455 (N_3455,N_843,N_783);
nor U3456 (N_3456,N_1889,N_522);
and U3457 (N_3457,N_578,N_1801);
and U3458 (N_3458,N_795,N_2151);
xnor U3459 (N_3459,N_2307,N_1360);
or U3460 (N_3460,N_118,N_822);
nor U3461 (N_3461,N_1575,N_1597);
or U3462 (N_3462,N_2314,N_459);
xor U3463 (N_3463,N_838,N_1093);
or U3464 (N_3464,N_946,N_1811);
or U3465 (N_3465,N_788,N_2498);
nand U3466 (N_3466,N_2428,N_1766);
and U3467 (N_3467,N_126,N_634);
xor U3468 (N_3468,N_1396,N_1014);
nor U3469 (N_3469,N_2239,N_616);
nand U3470 (N_3470,N_1771,N_719);
xor U3471 (N_3471,N_1049,N_197);
nor U3472 (N_3472,N_1397,N_2056);
or U3473 (N_3473,N_2181,N_2143);
nor U3474 (N_3474,N_350,N_244);
nor U3475 (N_3475,N_1081,N_2413);
nor U3476 (N_3476,N_675,N_387);
nand U3477 (N_3477,N_1897,N_714);
nand U3478 (N_3478,N_1572,N_1086);
nand U3479 (N_3479,N_400,N_2272);
or U3480 (N_3480,N_1001,N_1092);
or U3481 (N_3481,N_722,N_84);
and U3482 (N_3482,N_751,N_1191);
and U3483 (N_3483,N_2248,N_1836);
or U3484 (N_3484,N_1538,N_7);
xnor U3485 (N_3485,N_2384,N_944);
or U3486 (N_3486,N_1599,N_1103);
nand U3487 (N_3487,N_2276,N_120);
and U3488 (N_3488,N_954,N_1164);
or U3489 (N_3489,N_1560,N_2480);
nor U3490 (N_3490,N_637,N_1913);
xor U3491 (N_3491,N_330,N_351);
and U3492 (N_3492,N_2100,N_211);
and U3493 (N_3493,N_521,N_2450);
nor U3494 (N_3494,N_2140,N_698);
or U3495 (N_3495,N_797,N_1997);
nand U3496 (N_3496,N_1041,N_897);
nand U3497 (N_3497,N_583,N_2361);
nand U3498 (N_3498,N_2144,N_1344);
and U3499 (N_3499,N_1783,N_23);
nand U3500 (N_3500,N_595,N_1237);
nand U3501 (N_3501,N_746,N_680);
or U3502 (N_3502,N_1906,N_1398);
and U3503 (N_3503,N_2102,N_196);
nor U3504 (N_3504,N_741,N_558);
xnor U3505 (N_3505,N_1534,N_207);
or U3506 (N_3506,N_1570,N_2381);
or U3507 (N_3507,N_600,N_1850);
or U3508 (N_3508,N_1459,N_1144);
nand U3509 (N_3509,N_311,N_355);
nor U3510 (N_3510,N_1615,N_1646);
or U3511 (N_3511,N_1353,N_1877);
nand U3512 (N_3512,N_31,N_971);
nand U3513 (N_3513,N_928,N_39);
xnor U3514 (N_3514,N_2222,N_300);
and U3515 (N_3515,N_453,N_2454);
or U3516 (N_3516,N_801,N_736);
nand U3517 (N_3517,N_1656,N_1204);
nor U3518 (N_3518,N_1380,N_659);
xnor U3519 (N_3519,N_1569,N_584);
nand U3520 (N_3520,N_1507,N_1176);
nor U3521 (N_3521,N_1415,N_1287);
or U3522 (N_3522,N_16,N_692);
nor U3523 (N_3523,N_2015,N_605);
or U3524 (N_3524,N_2372,N_55);
xor U3525 (N_3525,N_1135,N_939);
or U3526 (N_3526,N_1096,N_475);
nor U3527 (N_3527,N_2147,N_2357);
nand U3528 (N_3528,N_742,N_870);
nand U3529 (N_3529,N_139,N_964);
or U3530 (N_3530,N_1106,N_2278);
and U3531 (N_3531,N_632,N_1071);
nand U3532 (N_3532,N_1734,N_1536);
xnor U3533 (N_3533,N_1712,N_625);
xnor U3534 (N_3534,N_957,N_37);
or U3535 (N_3535,N_457,N_2192);
and U3536 (N_3536,N_53,N_363);
xnor U3537 (N_3537,N_164,N_566);
xnor U3538 (N_3538,N_1688,N_65);
nand U3539 (N_3539,N_155,N_268);
or U3540 (N_3540,N_1944,N_1924);
xor U3541 (N_3541,N_904,N_528);
and U3542 (N_3542,N_1786,N_1774);
nor U3543 (N_3543,N_1677,N_2003);
nand U3544 (N_3544,N_2246,N_1193);
nor U3545 (N_3545,N_1365,N_1275);
nor U3546 (N_3546,N_1614,N_1241);
nand U3547 (N_3547,N_1827,N_249);
xnor U3548 (N_3548,N_1782,N_1128);
nor U3549 (N_3549,N_161,N_549);
nor U3550 (N_3550,N_1787,N_2282);
xor U3551 (N_3551,N_307,N_2365);
or U3552 (N_3552,N_1328,N_2086);
xor U3553 (N_3553,N_1016,N_112);
xnor U3554 (N_3554,N_1669,N_755);
nand U3555 (N_3555,N_1916,N_428);
nand U3556 (N_3556,N_1601,N_246);
and U3557 (N_3557,N_2113,N_2359);
xor U3558 (N_3558,N_881,N_1229);
or U3559 (N_3559,N_2392,N_379);
xor U3560 (N_3560,N_2474,N_563);
nor U3561 (N_3561,N_1905,N_2055);
and U3562 (N_3562,N_2313,N_857);
xor U3563 (N_3563,N_802,N_301);
or U3564 (N_3564,N_1763,N_1079);
xor U3565 (N_3565,N_2010,N_508);
or U3566 (N_3566,N_1127,N_1389);
nor U3567 (N_3567,N_1921,N_2368);
xor U3568 (N_3568,N_1740,N_190);
nand U3569 (N_3569,N_994,N_593);
xnor U3570 (N_3570,N_2205,N_314);
nand U3571 (N_3571,N_377,N_13);
nand U3572 (N_3572,N_1879,N_1142);
nor U3573 (N_3573,N_2254,N_757);
xnor U3574 (N_3574,N_1372,N_647);
nand U3575 (N_3575,N_1623,N_548);
or U3576 (N_3576,N_1562,N_127);
and U3577 (N_3577,N_855,N_1251);
nand U3578 (N_3578,N_365,N_420);
nand U3579 (N_3579,N_1510,N_509);
nand U3580 (N_3580,N_1378,N_1059);
or U3581 (N_3581,N_573,N_500);
and U3582 (N_3582,N_1390,N_1518);
nand U3583 (N_3583,N_639,N_1158);
nor U3584 (N_3584,N_366,N_1531);
xnor U3585 (N_3585,N_624,N_2279);
xnor U3586 (N_3586,N_1676,N_1406);
nand U3587 (N_3587,N_2261,N_339);
nor U3588 (N_3588,N_1852,N_833);
nand U3589 (N_3589,N_1388,N_527);
and U3590 (N_3590,N_226,N_1198);
nand U3591 (N_3591,N_2126,N_171);
nor U3592 (N_3592,N_901,N_2160);
and U3593 (N_3593,N_607,N_2183);
nor U3594 (N_3594,N_2045,N_397);
and U3595 (N_3595,N_810,N_1076);
or U3596 (N_3596,N_88,N_2194);
nor U3597 (N_3597,N_1943,N_1733);
or U3598 (N_3598,N_712,N_1131);
or U3599 (N_3599,N_22,N_2412);
nor U3600 (N_3600,N_1475,N_671);
nor U3601 (N_3601,N_1567,N_2195);
nor U3602 (N_3602,N_2495,N_2240);
xor U3603 (N_3603,N_1114,N_229);
or U3604 (N_3604,N_2386,N_655);
or U3605 (N_3605,N_242,N_1346);
or U3606 (N_3606,N_391,N_1483);
nor U3607 (N_3607,N_1336,N_1758);
xnor U3608 (N_3608,N_1043,N_359);
nor U3609 (N_3609,N_883,N_1788);
xor U3610 (N_3610,N_1012,N_1871);
and U3611 (N_3611,N_2199,N_596);
nand U3612 (N_3612,N_1427,N_761);
or U3613 (N_3613,N_1455,N_341);
nand U3614 (N_3614,N_708,N_1316);
xnor U3615 (N_3615,N_297,N_2068);
and U3616 (N_3616,N_1954,N_2175);
nand U3617 (N_3617,N_891,N_635);
xor U3618 (N_3618,N_193,N_678);
nand U3619 (N_3619,N_1203,N_867);
and U3620 (N_3620,N_1030,N_21);
or U3621 (N_3621,N_1208,N_1704);
nor U3622 (N_3622,N_34,N_305);
xor U3623 (N_3623,N_2133,N_999);
nor U3624 (N_3624,N_2031,N_1402);
nand U3625 (N_3625,N_348,N_594);
nand U3626 (N_3626,N_1830,N_2457);
and U3627 (N_3627,N_376,N_758);
or U3628 (N_3628,N_1781,N_1438);
xnor U3629 (N_3629,N_2431,N_517);
and U3630 (N_3630,N_2488,N_1927);
and U3631 (N_3631,N_11,N_2259);
and U3632 (N_3632,N_1760,N_662);
nor U3633 (N_3633,N_1087,N_1089);
xor U3634 (N_3634,N_559,N_1697);
or U3635 (N_3635,N_1392,N_2061);
and U3636 (N_3636,N_2336,N_442);
and U3637 (N_3637,N_2129,N_321);
nor U3638 (N_3638,N_2468,N_608);
nand U3639 (N_3639,N_1630,N_483);
or U3640 (N_3640,N_1116,N_2150);
or U3641 (N_3641,N_372,N_1722);
and U3642 (N_3642,N_4,N_1008);
and U3643 (N_3643,N_2485,N_858);
nand U3644 (N_3644,N_1157,N_2169);
nand U3645 (N_3645,N_2338,N_1355);
and U3646 (N_3646,N_462,N_1031);
xnor U3647 (N_3647,N_108,N_888);
nor U3648 (N_3648,N_1837,N_497);
and U3649 (N_3649,N_2243,N_1822);
xnor U3650 (N_3650,N_2421,N_865);
nand U3651 (N_3651,N_1859,N_76);
or U3652 (N_3652,N_1982,N_395);
and U3653 (N_3653,N_2448,N_2306);
and U3654 (N_3654,N_493,N_1988);
or U3655 (N_3655,N_1810,N_441);
xnor U3656 (N_3656,N_2182,N_501);
and U3657 (N_3657,N_1228,N_328);
and U3658 (N_3658,N_274,N_1299);
xor U3659 (N_3659,N_890,N_1969);
or U3660 (N_3660,N_633,N_2389);
nor U3661 (N_3661,N_2360,N_728);
nand U3662 (N_3662,N_1258,N_900);
xnor U3663 (N_3663,N_1662,N_2168);
or U3664 (N_3664,N_2373,N_2425);
nor U3665 (N_3665,N_116,N_59);
nor U3666 (N_3666,N_1308,N_1242);
nor U3667 (N_3667,N_353,N_2298);
or U3668 (N_3668,N_2073,N_568);
nor U3669 (N_3669,N_1594,N_1991);
nand U3670 (N_3670,N_1230,N_263);
and U3671 (N_3671,N_1655,N_1691);
nor U3672 (N_3672,N_92,N_520);
nand U3673 (N_3673,N_2139,N_1925);
nand U3674 (N_3674,N_940,N_912);
and U3675 (N_3675,N_304,N_54);
nand U3676 (N_3676,N_2418,N_2131);
xor U3677 (N_3677,N_2375,N_2451);
and U3678 (N_3678,N_949,N_2187);
xor U3679 (N_3679,N_2434,N_877);
xor U3680 (N_3680,N_1428,N_1429);
and U3681 (N_3681,N_1484,N_210);
xnor U3682 (N_3682,N_2220,N_511);
and U3683 (N_3683,N_546,N_1479);
xnor U3684 (N_3684,N_1977,N_970);
xor U3685 (N_3685,N_445,N_1265);
nor U3686 (N_3686,N_1376,N_652);
or U3687 (N_3687,N_1511,N_2014);
or U3688 (N_3688,N_1539,N_1162);
nand U3689 (N_3689,N_2247,N_284);
nand U3690 (N_3690,N_241,N_63);
or U3691 (N_3691,N_1294,N_976);
xor U3692 (N_3692,N_1707,N_1464);
and U3693 (N_3693,N_187,N_543);
and U3694 (N_3694,N_1932,N_2285);
and U3695 (N_3695,N_1578,N_44);
xnor U3696 (N_3696,N_950,N_811);
xnor U3697 (N_3697,N_2430,N_461);
or U3698 (N_3698,N_1101,N_71);
or U3699 (N_3699,N_871,N_537);
and U3700 (N_3700,N_2332,N_773);
nand U3701 (N_3701,N_2124,N_555);
nand U3702 (N_3702,N_1156,N_1568);
nor U3703 (N_3703,N_974,N_158);
nand U3704 (N_3704,N_1029,N_2161);
or U3705 (N_3705,N_1625,N_759);
xor U3706 (N_3706,N_485,N_525);
xnor U3707 (N_3707,N_1034,N_1450);
or U3708 (N_3708,N_661,N_564);
and U3709 (N_3709,N_1926,N_1448);
xnor U3710 (N_3710,N_313,N_1966);
nand U3711 (N_3711,N_1665,N_175);
nor U3712 (N_3712,N_38,N_404);
nor U3713 (N_3713,N_1690,N_1522);
nand U3714 (N_3714,N_170,N_1681);
and U3715 (N_3715,N_1259,N_1865);
xor U3716 (N_3716,N_630,N_1985);
or U3717 (N_3717,N_469,N_386);
xnor U3718 (N_3718,N_2473,N_1633);
nor U3719 (N_3719,N_2476,N_42);
or U3720 (N_3720,N_1245,N_1281);
nor U3721 (N_3721,N_1973,N_429);
xor U3722 (N_3722,N_2326,N_2101);
and U3723 (N_3723,N_2092,N_233);
nand U3724 (N_3724,N_930,N_1035);
xnor U3725 (N_3725,N_489,N_1217);
nor U3726 (N_3726,N_105,N_291);
xor U3727 (N_3727,N_852,N_1644);
nand U3728 (N_3728,N_1189,N_1465);
nand U3729 (N_3729,N_723,N_765);
nand U3730 (N_3730,N_818,N_1069);
or U3731 (N_3731,N_816,N_952);
xor U3732 (N_3732,N_238,N_617);
nand U3733 (N_3733,N_1107,N_1970);
nor U3734 (N_3734,N_1137,N_1898);
and U3735 (N_3735,N_1965,N_1009);
xnor U3736 (N_3736,N_466,N_134);
xor U3737 (N_3737,N_1818,N_1893);
and U3738 (N_3738,N_2271,N_1383);
nand U3739 (N_3739,N_1922,N_1233);
xnor U3740 (N_3740,N_570,N_2283);
or U3741 (N_3741,N_1663,N_1180);
or U3742 (N_3742,N_2284,N_325);
xor U3743 (N_3743,N_144,N_1068);
nand U3744 (N_3744,N_2409,N_1333);
xnor U3745 (N_3745,N_1513,N_1577);
and U3746 (N_3746,N_2226,N_1643);
and U3747 (N_3747,N_2242,N_731);
xnor U3748 (N_3748,N_2111,N_1075);
nor U3749 (N_3749,N_415,N_1433);
nor U3750 (N_3750,N_1988,N_1339);
nor U3751 (N_3751,N_215,N_829);
and U3752 (N_3752,N_1218,N_791);
or U3753 (N_3753,N_1348,N_2090);
and U3754 (N_3754,N_100,N_2094);
nand U3755 (N_3755,N_888,N_2093);
xnor U3756 (N_3756,N_2368,N_1343);
nor U3757 (N_3757,N_676,N_1738);
and U3758 (N_3758,N_1737,N_342);
nor U3759 (N_3759,N_2228,N_1883);
nand U3760 (N_3760,N_1335,N_472);
or U3761 (N_3761,N_403,N_1117);
nor U3762 (N_3762,N_676,N_2252);
nor U3763 (N_3763,N_2286,N_1753);
and U3764 (N_3764,N_168,N_925);
nor U3765 (N_3765,N_1981,N_1061);
xor U3766 (N_3766,N_1683,N_358);
or U3767 (N_3767,N_1503,N_1669);
nand U3768 (N_3768,N_1457,N_1346);
or U3769 (N_3769,N_1110,N_1330);
nor U3770 (N_3770,N_1746,N_2031);
nand U3771 (N_3771,N_2417,N_1836);
or U3772 (N_3772,N_2099,N_1807);
and U3773 (N_3773,N_200,N_705);
xnor U3774 (N_3774,N_1385,N_1134);
nor U3775 (N_3775,N_520,N_1042);
and U3776 (N_3776,N_1377,N_416);
nor U3777 (N_3777,N_1164,N_1634);
nor U3778 (N_3778,N_1459,N_508);
xor U3779 (N_3779,N_2008,N_395);
xor U3780 (N_3780,N_1351,N_1252);
nor U3781 (N_3781,N_1318,N_691);
nor U3782 (N_3782,N_1654,N_1138);
nor U3783 (N_3783,N_1948,N_2152);
xnor U3784 (N_3784,N_2407,N_1149);
or U3785 (N_3785,N_2495,N_2092);
nand U3786 (N_3786,N_552,N_2448);
nand U3787 (N_3787,N_1218,N_337);
xnor U3788 (N_3788,N_566,N_396);
or U3789 (N_3789,N_339,N_2309);
nor U3790 (N_3790,N_2258,N_2016);
nand U3791 (N_3791,N_240,N_2161);
or U3792 (N_3792,N_2483,N_454);
nand U3793 (N_3793,N_1760,N_1354);
nor U3794 (N_3794,N_1257,N_755);
nor U3795 (N_3795,N_925,N_947);
or U3796 (N_3796,N_1775,N_461);
nand U3797 (N_3797,N_1483,N_604);
xnor U3798 (N_3798,N_2216,N_1641);
xor U3799 (N_3799,N_1339,N_1567);
xor U3800 (N_3800,N_1174,N_380);
nand U3801 (N_3801,N_2048,N_1850);
or U3802 (N_3802,N_2324,N_347);
and U3803 (N_3803,N_2169,N_1833);
and U3804 (N_3804,N_1841,N_336);
or U3805 (N_3805,N_603,N_218);
xor U3806 (N_3806,N_638,N_2116);
nand U3807 (N_3807,N_943,N_1294);
and U3808 (N_3808,N_710,N_1527);
xnor U3809 (N_3809,N_1572,N_145);
xnor U3810 (N_3810,N_1287,N_859);
nand U3811 (N_3811,N_260,N_376);
xor U3812 (N_3812,N_1406,N_1305);
xnor U3813 (N_3813,N_298,N_739);
or U3814 (N_3814,N_848,N_766);
or U3815 (N_3815,N_1918,N_1402);
and U3816 (N_3816,N_171,N_704);
xnor U3817 (N_3817,N_1700,N_86);
and U3818 (N_3818,N_489,N_777);
and U3819 (N_3819,N_2259,N_433);
or U3820 (N_3820,N_1688,N_631);
or U3821 (N_3821,N_651,N_193);
or U3822 (N_3822,N_480,N_1177);
and U3823 (N_3823,N_1614,N_1008);
or U3824 (N_3824,N_2404,N_1627);
nor U3825 (N_3825,N_1015,N_2222);
nand U3826 (N_3826,N_2377,N_1830);
or U3827 (N_3827,N_1056,N_742);
or U3828 (N_3828,N_1723,N_1008);
xnor U3829 (N_3829,N_624,N_389);
nand U3830 (N_3830,N_495,N_1001);
or U3831 (N_3831,N_2322,N_2452);
nand U3832 (N_3832,N_1210,N_2323);
and U3833 (N_3833,N_1638,N_2266);
nand U3834 (N_3834,N_79,N_2144);
nor U3835 (N_3835,N_1265,N_2434);
xor U3836 (N_3836,N_1490,N_1020);
and U3837 (N_3837,N_171,N_602);
and U3838 (N_3838,N_329,N_1575);
and U3839 (N_3839,N_180,N_1658);
nor U3840 (N_3840,N_1143,N_1599);
and U3841 (N_3841,N_30,N_724);
nor U3842 (N_3842,N_353,N_1012);
or U3843 (N_3843,N_121,N_165);
or U3844 (N_3844,N_306,N_526);
or U3845 (N_3845,N_1378,N_1645);
and U3846 (N_3846,N_1451,N_1474);
nand U3847 (N_3847,N_1493,N_753);
or U3848 (N_3848,N_928,N_1489);
nand U3849 (N_3849,N_1040,N_239);
nor U3850 (N_3850,N_404,N_1218);
or U3851 (N_3851,N_1516,N_578);
xnor U3852 (N_3852,N_790,N_865);
xor U3853 (N_3853,N_698,N_844);
or U3854 (N_3854,N_2390,N_1648);
nand U3855 (N_3855,N_231,N_2263);
or U3856 (N_3856,N_44,N_833);
and U3857 (N_3857,N_1967,N_1086);
nand U3858 (N_3858,N_2000,N_1926);
and U3859 (N_3859,N_2131,N_2074);
xor U3860 (N_3860,N_2460,N_2096);
xnor U3861 (N_3861,N_314,N_20);
xnor U3862 (N_3862,N_2214,N_746);
and U3863 (N_3863,N_1168,N_1558);
xor U3864 (N_3864,N_1012,N_2432);
nand U3865 (N_3865,N_2456,N_2472);
nand U3866 (N_3866,N_1512,N_1649);
nand U3867 (N_3867,N_1035,N_1037);
and U3868 (N_3868,N_2100,N_1908);
nor U3869 (N_3869,N_227,N_1063);
xnor U3870 (N_3870,N_70,N_175);
nand U3871 (N_3871,N_1305,N_354);
or U3872 (N_3872,N_2239,N_1097);
and U3873 (N_3873,N_110,N_1107);
nor U3874 (N_3874,N_1529,N_1030);
xnor U3875 (N_3875,N_1870,N_923);
xnor U3876 (N_3876,N_839,N_379);
or U3877 (N_3877,N_43,N_1817);
or U3878 (N_3878,N_724,N_88);
nand U3879 (N_3879,N_1908,N_1798);
or U3880 (N_3880,N_2408,N_95);
nor U3881 (N_3881,N_2284,N_1777);
or U3882 (N_3882,N_627,N_581);
or U3883 (N_3883,N_1334,N_2053);
nor U3884 (N_3884,N_2095,N_1486);
and U3885 (N_3885,N_34,N_281);
nor U3886 (N_3886,N_1447,N_1900);
or U3887 (N_3887,N_2045,N_1126);
and U3888 (N_3888,N_313,N_2491);
or U3889 (N_3889,N_1753,N_182);
or U3890 (N_3890,N_1228,N_985);
nor U3891 (N_3891,N_1369,N_945);
and U3892 (N_3892,N_1263,N_1187);
xnor U3893 (N_3893,N_1152,N_272);
or U3894 (N_3894,N_1158,N_1891);
or U3895 (N_3895,N_1211,N_740);
or U3896 (N_3896,N_87,N_2455);
or U3897 (N_3897,N_2305,N_1019);
nor U3898 (N_3898,N_171,N_2401);
or U3899 (N_3899,N_1854,N_935);
and U3900 (N_3900,N_294,N_457);
nand U3901 (N_3901,N_241,N_2399);
or U3902 (N_3902,N_2054,N_10);
xor U3903 (N_3903,N_613,N_1733);
and U3904 (N_3904,N_636,N_1529);
nor U3905 (N_3905,N_2298,N_1695);
and U3906 (N_3906,N_80,N_2347);
or U3907 (N_3907,N_1640,N_2478);
nor U3908 (N_3908,N_592,N_1709);
xnor U3909 (N_3909,N_1820,N_1061);
or U3910 (N_3910,N_790,N_2167);
and U3911 (N_3911,N_1657,N_1629);
nor U3912 (N_3912,N_1772,N_109);
nor U3913 (N_3913,N_1053,N_1650);
xnor U3914 (N_3914,N_1529,N_2277);
or U3915 (N_3915,N_1317,N_2466);
and U3916 (N_3916,N_524,N_1075);
nor U3917 (N_3917,N_1858,N_2028);
xor U3918 (N_3918,N_1755,N_1364);
nand U3919 (N_3919,N_2189,N_917);
and U3920 (N_3920,N_10,N_2325);
nor U3921 (N_3921,N_890,N_2231);
nand U3922 (N_3922,N_1036,N_1216);
or U3923 (N_3923,N_734,N_1926);
and U3924 (N_3924,N_1393,N_1024);
or U3925 (N_3925,N_965,N_2234);
and U3926 (N_3926,N_2148,N_1734);
xor U3927 (N_3927,N_2153,N_1464);
xor U3928 (N_3928,N_676,N_303);
and U3929 (N_3929,N_578,N_1197);
xor U3930 (N_3930,N_812,N_365);
or U3931 (N_3931,N_1023,N_1118);
nand U3932 (N_3932,N_559,N_586);
or U3933 (N_3933,N_1846,N_2049);
nand U3934 (N_3934,N_530,N_69);
and U3935 (N_3935,N_862,N_428);
nand U3936 (N_3936,N_551,N_350);
or U3937 (N_3937,N_2373,N_763);
and U3938 (N_3938,N_1927,N_2031);
nor U3939 (N_3939,N_2283,N_59);
nor U3940 (N_3940,N_1685,N_2481);
xor U3941 (N_3941,N_1985,N_2211);
xnor U3942 (N_3942,N_847,N_1615);
nand U3943 (N_3943,N_735,N_2343);
nor U3944 (N_3944,N_725,N_104);
or U3945 (N_3945,N_535,N_144);
nor U3946 (N_3946,N_2130,N_1674);
or U3947 (N_3947,N_1344,N_94);
xor U3948 (N_3948,N_1516,N_666);
xor U3949 (N_3949,N_553,N_899);
xor U3950 (N_3950,N_2153,N_259);
and U3951 (N_3951,N_978,N_243);
nand U3952 (N_3952,N_2230,N_1597);
nor U3953 (N_3953,N_1576,N_2475);
xor U3954 (N_3954,N_1926,N_1626);
or U3955 (N_3955,N_124,N_159);
nor U3956 (N_3956,N_2468,N_30);
xnor U3957 (N_3957,N_1451,N_429);
nor U3958 (N_3958,N_1995,N_831);
nor U3959 (N_3959,N_1025,N_1890);
xnor U3960 (N_3960,N_1564,N_320);
xor U3961 (N_3961,N_1137,N_2449);
and U3962 (N_3962,N_979,N_736);
or U3963 (N_3963,N_2254,N_1043);
and U3964 (N_3964,N_184,N_32);
and U3965 (N_3965,N_1523,N_2453);
or U3966 (N_3966,N_506,N_300);
or U3967 (N_3967,N_2110,N_991);
or U3968 (N_3968,N_840,N_330);
nand U3969 (N_3969,N_829,N_784);
nand U3970 (N_3970,N_1011,N_1148);
or U3971 (N_3971,N_337,N_2303);
xnor U3972 (N_3972,N_867,N_1350);
or U3973 (N_3973,N_2062,N_1536);
and U3974 (N_3974,N_1144,N_187);
and U3975 (N_3975,N_700,N_122);
nand U3976 (N_3976,N_2190,N_1058);
xnor U3977 (N_3977,N_1076,N_1246);
and U3978 (N_3978,N_2230,N_1754);
and U3979 (N_3979,N_875,N_1597);
or U3980 (N_3980,N_869,N_1061);
and U3981 (N_3981,N_1776,N_681);
nand U3982 (N_3982,N_1296,N_1971);
or U3983 (N_3983,N_541,N_553);
and U3984 (N_3984,N_790,N_2339);
nor U3985 (N_3985,N_394,N_1461);
and U3986 (N_3986,N_101,N_1299);
nor U3987 (N_3987,N_895,N_2459);
and U3988 (N_3988,N_227,N_2472);
nand U3989 (N_3989,N_2266,N_281);
nand U3990 (N_3990,N_887,N_1423);
nor U3991 (N_3991,N_2303,N_2195);
and U3992 (N_3992,N_374,N_185);
and U3993 (N_3993,N_393,N_1788);
or U3994 (N_3994,N_599,N_2121);
nand U3995 (N_3995,N_1587,N_1450);
xnor U3996 (N_3996,N_1227,N_108);
and U3997 (N_3997,N_845,N_765);
nand U3998 (N_3998,N_1902,N_52);
nand U3999 (N_3999,N_1448,N_1590);
or U4000 (N_4000,N_1135,N_2443);
or U4001 (N_4001,N_1502,N_977);
nor U4002 (N_4002,N_36,N_322);
xnor U4003 (N_4003,N_311,N_2358);
nor U4004 (N_4004,N_2117,N_929);
xnor U4005 (N_4005,N_2217,N_1685);
nand U4006 (N_4006,N_1012,N_1701);
and U4007 (N_4007,N_721,N_1865);
nor U4008 (N_4008,N_2303,N_629);
or U4009 (N_4009,N_1160,N_2432);
and U4010 (N_4010,N_842,N_580);
or U4011 (N_4011,N_2388,N_1492);
xor U4012 (N_4012,N_1979,N_1377);
nor U4013 (N_4013,N_978,N_212);
xor U4014 (N_4014,N_1973,N_880);
and U4015 (N_4015,N_456,N_315);
xor U4016 (N_4016,N_1227,N_766);
or U4017 (N_4017,N_1542,N_758);
xnor U4018 (N_4018,N_1147,N_113);
nand U4019 (N_4019,N_2281,N_113);
and U4020 (N_4020,N_439,N_2329);
nand U4021 (N_4021,N_386,N_1736);
or U4022 (N_4022,N_20,N_1626);
or U4023 (N_4023,N_194,N_2065);
nand U4024 (N_4024,N_88,N_2214);
and U4025 (N_4025,N_1037,N_1161);
and U4026 (N_4026,N_2230,N_1264);
nand U4027 (N_4027,N_1692,N_1183);
xnor U4028 (N_4028,N_1907,N_2111);
and U4029 (N_4029,N_2270,N_2244);
nor U4030 (N_4030,N_559,N_2300);
or U4031 (N_4031,N_825,N_1209);
xor U4032 (N_4032,N_1645,N_2497);
xnor U4033 (N_4033,N_1702,N_435);
and U4034 (N_4034,N_776,N_851);
xnor U4035 (N_4035,N_1496,N_604);
xnor U4036 (N_4036,N_2456,N_1586);
or U4037 (N_4037,N_2145,N_796);
and U4038 (N_4038,N_1823,N_313);
xnor U4039 (N_4039,N_2241,N_2351);
nor U4040 (N_4040,N_474,N_359);
and U4041 (N_4041,N_2209,N_343);
nor U4042 (N_4042,N_970,N_2304);
and U4043 (N_4043,N_2043,N_1696);
and U4044 (N_4044,N_447,N_558);
xnor U4045 (N_4045,N_1090,N_967);
nor U4046 (N_4046,N_2350,N_560);
nor U4047 (N_4047,N_1142,N_2182);
nor U4048 (N_4048,N_2215,N_1377);
and U4049 (N_4049,N_1812,N_476);
and U4050 (N_4050,N_1443,N_1816);
and U4051 (N_4051,N_1354,N_2360);
and U4052 (N_4052,N_1763,N_1965);
and U4053 (N_4053,N_243,N_509);
nand U4054 (N_4054,N_1700,N_2357);
xor U4055 (N_4055,N_2223,N_558);
or U4056 (N_4056,N_1536,N_19);
or U4057 (N_4057,N_299,N_1917);
xnor U4058 (N_4058,N_782,N_672);
nand U4059 (N_4059,N_1289,N_811);
or U4060 (N_4060,N_497,N_1644);
xnor U4061 (N_4061,N_1902,N_1981);
or U4062 (N_4062,N_2079,N_1942);
xor U4063 (N_4063,N_1587,N_1378);
nor U4064 (N_4064,N_143,N_542);
xnor U4065 (N_4065,N_948,N_239);
nor U4066 (N_4066,N_1438,N_510);
nand U4067 (N_4067,N_261,N_903);
nor U4068 (N_4068,N_139,N_170);
xnor U4069 (N_4069,N_1744,N_1604);
xnor U4070 (N_4070,N_1881,N_1150);
and U4071 (N_4071,N_1419,N_2115);
nand U4072 (N_4072,N_48,N_1298);
nand U4073 (N_4073,N_699,N_1537);
and U4074 (N_4074,N_2453,N_1416);
xor U4075 (N_4075,N_1870,N_1032);
nand U4076 (N_4076,N_776,N_1197);
or U4077 (N_4077,N_566,N_1290);
or U4078 (N_4078,N_651,N_1361);
nor U4079 (N_4079,N_1763,N_1583);
nor U4080 (N_4080,N_407,N_2027);
nor U4081 (N_4081,N_649,N_291);
xor U4082 (N_4082,N_17,N_1723);
or U4083 (N_4083,N_1534,N_2035);
xnor U4084 (N_4084,N_948,N_713);
nand U4085 (N_4085,N_528,N_2028);
and U4086 (N_4086,N_49,N_620);
nor U4087 (N_4087,N_2369,N_2013);
xnor U4088 (N_4088,N_1497,N_1199);
and U4089 (N_4089,N_2406,N_213);
and U4090 (N_4090,N_2185,N_1262);
xor U4091 (N_4091,N_90,N_611);
nand U4092 (N_4092,N_276,N_1449);
or U4093 (N_4093,N_1061,N_1451);
or U4094 (N_4094,N_767,N_628);
nor U4095 (N_4095,N_794,N_2117);
nand U4096 (N_4096,N_1288,N_197);
xnor U4097 (N_4097,N_890,N_630);
and U4098 (N_4098,N_1068,N_1727);
xor U4099 (N_4099,N_962,N_115);
or U4100 (N_4100,N_1572,N_429);
nand U4101 (N_4101,N_1398,N_1458);
nand U4102 (N_4102,N_439,N_212);
xor U4103 (N_4103,N_92,N_2328);
xor U4104 (N_4104,N_889,N_1490);
or U4105 (N_4105,N_4,N_1571);
and U4106 (N_4106,N_1068,N_1488);
nor U4107 (N_4107,N_2046,N_1612);
and U4108 (N_4108,N_101,N_2085);
nor U4109 (N_4109,N_14,N_2421);
xor U4110 (N_4110,N_374,N_1061);
nand U4111 (N_4111,N_893,N_1448);
nand U4112 (N_4112,N_1763,N_1860);
nor U4113 (N_4113,N_1742,N_2204);
and U4114 (N_4114,N_2107,N_1732);
nand U4115 (N_4115,N_458,N_1189);
xor U4116 (N_4116,N_105,N_18);
and U4117 (N_4117,N_820,N_1301);
or U4118 (N_4118,N_1801,N_1575);
xnor U4119 (N_4119,N_1404,N_1753);
nand U4120 (N_4120,N_700,N_2331);
nand U4121 (N_4121,N_1420,N_915);
nor U4122 (N_4122,N_1398,N_955);
nand U4123 (N_4123,N_462,N_1837);
nor U4124 (N_4124,N_2291,N_1272);
nand U4125 (N_4125,N_241,N_2267);
or U4126 (N_4126,N_2281,N_396);
xor U4127 (N_4127,N_397,N_41);
nor U4128 (N_4128,N_598,N_1134);
or U4129 (N_4129,N_921,N_2166);
nand U4130 (N_4130,N_1797,N_1854);
nor U4131 (N_4131,N_1729,N_361);
or U4132 (N_4132,N_211,N_527);
nor U4133 (N_4133,N_699,N_1624);
nor U4134 (N_4134,N_260,N_1708);
and U4135 (N_4135,N_1321,N_1841);
and U4136 (N_4136,N_354,N_118);
xor U4137 (N_4137,N_677,N_2473);
or U4138 (N_4138,N_1021,N_1965);
or U4139 (N_4139,N_28,N_168);
or U4140 (N_4140,N_66,N_603);
and U4141 (N_4141,N_1086,N_929);
nand U4142 (N_4142,N_2231,N_2012);
nor U4143 (N_4143,N_1524,N_1827);
nand U4144 (N_4144,N_2210,N_1951);
nand U4145 (N_4145,N_1902,N_866);
and U4146 (N_4146,N_1502,N_1954);
and U4147 (N_4147,N_113,N_1883);
or U4148 (N_4148,N_185,N_917);
nor U4149 (N_4149,N_1754,N_508);
and U4150 (N_4150,N_866,N_552);
or U4151 (N_4151,N_315,N_1726);
or U4152 (N_4152,N_1479,N_681);
or U4153 (N_4153,N_1881,N_1948);
nand U4154 (N_4154,N_2495,N_665);
and U4155 (N_4155,N_2312,N_1859);
or U4156 (N_4156,N_191,N_36);
nand U4157 (N_4157,N_997,N_1443);
xor U4158 (N_4158,N_779,N_1713);
nor U4159 (N_4159,N_2466,N_1474);
xor U4160 (N_4160,N_2447,N_503);
or U4161 (N_4161,N_819,N_882);
xor U4162 (N_4162,N_561,N_2159);
and U4163 (N_4163,N_1696,N_269);
or U4164 (N_4164,N_1006,N_1116);
xnor U4165 (N_4165,N_1600,N_2194);
or U4166 (N_4166,N_1757,N_1721);
and U4167 (N_4167,N_538,N_2386);
nor U4168 (N_4168,N_1270,N_614);
nand U4169 (N_4169,N_1234,N_805);
nor U4170 (N_4170,N_505,N_1758);
and U4171 (N_4171,N_493,N_1081);
and U4172 (N_4172,N_1739,N_614);
and U4173 (N_4173,N_1238,N_1371);
xor U4174 (N_4174,N_325,N_889);
nor U4175 (N_4175,N_1059,N_55);
nand U4176 (N_4176,N_156,N_733);
nor U4177 (N_4177,N_784,N_838);
or U4178 (N_4178,N_1281,N_1335);
nor U4179 (N_4179,N_1798,N_1549);
nor U4180 (N_4180,N_939,N_560);
nand U4181 (N_4181,N_1860,N_1434);
xor U4182 (N_4182,N_1561,N_618);
nor U4183 (N_4183,N_587,N_1415);
nand U4184 (N_4184,N_2147,N_53);
nor U4185 (N_4185,N_799,N_696);
or U4186 (N_4186,N_425,N_2319);
nand U4187 (N_4187,N_743,N_2185);
or U4188 (N_4188,N_1275,N_2193);
nand U4189 (N_4189,N_1696,N_1456);
xnor U4190 (N_4190,N_1073,N_629);
or U4191 (N_4191,N_2372,N_1639);
or U4192 (N_4192,N_2396,N_1225);
xor U4193 (N_4193,N_693,N_1091);
and U4194 (N_4194,N_143,N_1080);
or U4195 (N_4195,N_1088,N_2114);
nand U4196 (N_4196,N_2101,N_1864);
xor U4197 (N_4197,N_84,N_222);
nor U4198 (N_4198,N_1316,N_1635);
nor U4199 (N_4199,N_1387,N_1868);
and U4200 (N_4200,N_712,N_252);
nand U4201 (N_4201,N_1677,N_1157);
nand U4202 (N_4202,N_2457,N_251);
xor U4203 (N_4203,N_2141,N_2435);
and U4204 (N_4204,N_1182,N_1520);
or U4205 (N_4205,N_1932,N_1145);
or U4206 (N_4206,N_861,N_1943);
xnor U4207 (N_4207,N_1920,N_2284);
or U4208 (N_4208,N_929,N_2157);
and U4209 (N_4209,N_9,N_1860);
nand U4210 (N_4210,N_174,N_1956);
nor U4211 (N_4211,N_2021,N_1835);
and U4212 (N_4212,N_2159,N_1006);
and U4213 (N_4213,N_2097,N_767);
xor U4214 (N_4214,N_192,N_315);
nand U4215 (N_4215,N_2308,N_786);
xor U4216 (N_4216,N_914,N_1543);
xnor U4217 (N_4217,N_1562,N_303);
nand U4218 (N_4218,N_1137,N_917);
or U4219 (N_4219,N_2359,N_74);
and U4220 (N_4220,N_250,N_169);
nor U4221 (N_4221,N_245,N_964);
nor U4222 (N_4222,N_1670,N_294);
nor U4223 (N_4223,N_183,N_1778);
nand U4224 (N_4224,N_1314,N_821);
or U4225 (N_4225,N_456,N_737);
xor U4226 (N_4226,N_969,N_1027);
and U4227 (N_4227,N_982,N_1551);
and U4228 (N_4228,N_1941,N_420);
nand U4229 (N_4229,N_2033,N_1140);
and U4230 (N_4230,N_2380,N_1354);
or U4231 (N_4231,N_815,N_1396);
xor U4232 (N_4232,N_946,N_2418);
nor U4233 (N_4233,N_2056,N_1659);
and U4234 (N_4234,N_1968,N_1541);
xnor U4235 (N_4235,N_260,N_1161);
and U4236 (N_4236,N_1118,N_250);
xnor U4237 (N_4237,N_764,N_1721);
nor U4238 (N_4238,N_2457,N_792);
and U4239 (N_4239,N_885,N_927);
xor U4240 (N_4240,N_250,N_923);
nand U4241 (N_4241,N_1744,N_608);
or U4242 (N_4242,N_1668,N_2045);
or U4243 (N_4243,N_1487,N_2446);
and U4244 (N_4244,N_666,N_1844);
xnor U4245 (N_4245,N_817,N_1360);
nand U4246 (N_4246,N_366,N_1764);
xor U4247 (N_4247,N_390,N_966);
or U4248 (N_4248,N_1457,N_640);
xor U4249 (N_4249,N_704,N_2171);
nor U4250 (N_4250,N_285,N_1797);
nand U4251 (N_4251,N_1540,N_128);
or U4252 (N_4252,N_2039,N_707);
or U4253 (N_4253,N_1360,N_290);
or U4254 (N_4254,N_525,N_410);
nor U4255 (N_4255,N_1941,N_2010);
and U4256 (N_4256,N_578,N_1906);
or U4257 (N_4257,N_1919,N_2402);
nor U4258 (N_4258,N_2216,N_995);
and U4259 (N_4259,N_2252,N_496);
nor U4260 (N_4260,N_540,N_1076);
and U4261 (N_4261,N_2285,N_1107);
nand U4262 (N_4262,N_1405,N_2320);
and U4263 (N_4263,N_2109,N_1938);
or U4264 (N_4264,N_1880,N_393);
xor U4265 (N_4265,N_66,N_1243);
or U4266 (N_4266,N_1736,N_1014);
nor U4267 (N_4267,N_287,N_2252);
nand U4268 (N_4268,N_1812,N_1856);
nand U4269 (N_4269,N_2152,N_2079);
nand U4270 (N_4270,N_958,N_1986);
xnor U4271 (N_4271,N_574,N_195);
nor U4272 (N_4272,N_967,N_895);
or U4273 (N_4273,N_41,N_1272);
nand U4274 (N_4274,N_2208,N_1383);
xor U4275 (N_4275,N_448,N_1966);
xor U4276 (N_4276,N_1393,N_681);
and U4277 (N_4277,N_563,N_1986);
nor U4278 (N_4278,N_2266,N_283);
nor U4279 (N_4279,N_1206,N_2480);
nor U4280 (N_4280,N_1463,N_1879);
nor U4281 (N_4281,N_992,N_2238);
nor U4282 (N_4282,N_350,N_2165);
and U4283 (N_4283,N_2033,N_2284);
or U4284 (N_4284,N_1797,N_1593);
and U4285 (N_4285,N_1770,N_1701);
nand U4286 (N_4286,N_517,N_1944);
xnor U4287 (N_4287,N_1920,N_673);
xor U4288 (N_4288,N_1063,N_1594);
or U4289 (N_4289,N_2260,N_24);
xor U4290 (N_4290,N_1544,N_2383);
and U4291 (N_4291,N_1911,N_1257);
or U4292 (N_4292,N_326,N_1183);
or U4293 (N_4293,N_2098,N_2191);
nor U4294 (N_4294,N_216,N_466);
or U4295 (N_4295,N_1930,N_396);
or U4296 (N_4296,N_1556,N_1835);
or U4297 (N_4297,N_342,N_2059);
nor U4298 (N_4298,N_1451,N_2204);
xnor U4299 (N_4299,N_1998,N_1086);
nand U4300 (N_4300,N_1705,N_2163);
and U4301 (N_4301,N_464,N_2046);
and U4302 (N_4302,N_2174,N_212);
nor U4303 (N_4303,N_1784,N_320);
xnor U4304 (N_4304,N_2387,N_1863);
nor U4305 (N_4305,N_976,N_855);
and U4306 (N_4306,N_623,N_1806);
and U4307 (N_4307,N_1526,N_644);
and U4308 (N_4308,N_699,N_1759);
or U4309 (N_4309,N_489,N_440);
xnor U4310 (N_4310,N_1561,N_1039);
nor U4311 (N_4311,N_1440,N_583);
xnor U4312 (N_4312,N_1074,N_1856);
xnor U4313 (N_4313,N_943,N_2433);
or U4314 (N_4314,N_94,N_907);
and U4315 (N_4315,N_695,N_1327);
nand U4316 (N_4316,N_1374,N_941);
or U4317 (N_4317,N_849,N_60);
xnor U4318 (N_4318,N_1584,N_2078);
and U4319 (N_4319,N_1711,N_1038);
nor U4320 (N_4320,N_1772,N_966);
nand U4321 (N_4321,N_824,N_12);
xor U4322 (N_4322,N_2191,N_1485);
or U4323 (N_4323,N_2192,N_1871);
and U4324 (N_4324,N_30,N_60);
nand U4325 (N_4325,N_465,N_570);
nand U4326 (N_4326,N_388,N_1039);
nand U4327 (N_4327,N_2382,N_1260);
and U4328 (N_4328,N_1813,N_1239);
nor U4329 (N_4329,N_1176,N_2434);
nand U4330 (N_4330,N_1784,N_783);
xor U4331 (N_4331,N_1435,N_1955);
and U4332 (N_4332,N_2183,N_1598);
and U4333 (N_4333,N_1793,N_251);
nand U4334 (N_4334,N_1225,N_1862);
or U4335 (N_4335,N_485,N_1200);
nand U4336 (N_4336,N_1067,N_158);
nand U4337 (N_4337,N_2479,N_115);
and U4338 (N_4338,N_1943,N_223);
and U4339 (N_4339,N_666,N_1520);
xnor U4340 (N_4340,N_1044,N_1823);
nor U4341 (N_4341,N_2312,N_1874);
nand U4342 (N_4342,N_238,N_1419);
and U4343 (N_4343,N_1721,N_1502);
or U4344 (N_4344,N_754,N_783);
or U4345 (N_4345,N_2125,N_117);
xor U4346 (N_4346,N_929,N_1157);
nand U4347 (N_4347,N_1798,N_1429);
nor U4348 (N_4348,N_1043,N_726);
nand U4349 (N_4349,N_241,N_153);
and U4350 (N_4350,N_1375,N_1685);
nand U4351 (N_4351,N_2227,N_22);
nor U4352 (N_4352,N_783,N_1466);
nor U4353 (N_4353,N_1286,N_1085);
or U4354 (N_4354,N_867,N_71);
nor U4355 (N_4355,N_271,N_1510);
or U4356 (N_4356,N_2255,N_767);
nor U4357 (N_4357,N_1249,N_966);
nor U4358 (N_4358,N_1551,N_1988);
nand U4359 (N_4359,N_2191,N_661);
nor U4360 (N_4360,N_1211,N_819);
or U4361 (N_4361,N_376,N_210);
nand U4362 (N_4362,N_737,N_381);
nor U4363 (N_4363,N_2330,N_2169);
xor U4364 (N_4364,N_359,N_1127);
and U4365 (N_4365,N_1855,N_318);
nand U4366 (N_4366,N_2357,N_2456);
and U4367 (N_4367,N_2388,N_66);
nor U4368 (N_4368,N_1009,N_766);
and U4369 (N_4369,N_15,N_2485);
xor U4370 (N_4370,N_630,N_1251);
xnor U4371 (N_4371,N_1537,N_524);
xor U4372 (N_4372,N_2294,N_2252);
nand U4373 (N_4373,N_2481,N_317);
nand U4374 (N_4374,N_885,N_1900);
xor U4375 (N_4375,N_1192,N_2145);
xnor U4376 (N_4376,N_1069,N_1696);
or U4377 (N_4377,N_2267,N_175);
or U4378 (N_4378,N_2470,N_2419);
xor U4379 (N_4379,N_312,N_280);
xor U4380 (N_4380,N_2426,N_1833);
nor U4381 (N_4381,N_2347,N_1776);
xor U4382 (N_4382,N_1152,N_274);
xor U4383 (N_4383,N_1893,N_1348);
xnor U4384 (N_4384,N_1032,N_1552);
or U4385 (N_4385,N_2429,N_1946);
xnor U4386 (N_4386,N_2335,N_1073);
and U4387 (N_4387,N_1409,N_2387);
or U4388 (N_4388,N_894,N_250);
nor U4389 (N_4389,N_2270,N_1852);
and U4390 (N_4390,N_1857,N_1350);
nand U4391 (N_4391,N_1214,N_6);
and U4392 (N_4392,N_2035,N_792);
and U4393 (N_4393,N_736,N_2436);
and U4394 (N_4394,N_1535,N_1138);
xnor U4395 (N_4395,N_1755,N_923);
xnor U4396 (N_4396,N_1866,N_746);
nand U4397 (N_4397,N_2480,N_2161);
nand U4398 (N_4398,N_1706,N_1848);
or U4399 (N_4399,N_1236,N_64);
and U4400 (N_4400,N_385,N_967);
or U4401 (N_4401,N_2206,N_983);
or U4402 (N_4402,N_2088,N_326);
and U4403 (N_4403,N_940,N_233);
xnor U4404 (N_4404,N_1723,N_2153);
nor U4405 (N_4405,N_2223,N_1728);
xor U4406 (N_4406,N_697,N_1336);
or U4407 (N_4407,N_1833,N_1291);
nor U4408 (N_4408,N_890,N_1134);
or U4409 (N_4409,N_2285,N_1094);
xnor U4410 (N_4410,N_2140,N_1136);
or U4411 (N_4411,N_2404,N_2292);
nand U4412 (N_4412,N_658,N_1033);
nor U4413 (N_4413,N_142,N_1456);
xnor U4414 (N_4414,N_951,N_1123);
and U4415 (N_4415,N_1426,N_2428);
nor U4416 (N_4416,N_339,N_74);
nand U4417 (N_4417,N_57,N_1964);
xnor U4418 (N_4418,N_1832,N_509);
nand U4419 (N_4419,N_2046,N_132);
xor U4420 (N_4420,N_1906,N_2008);
nor U4421 (N_4421,N_51,N_1830);
or U4422 (N_4422,N_1392,N_534);
nor U4423 (N_4423,N_520,N_1894);
xor U4424 (N_4424,N_2339,N_222);
xnor U4425 (N_4425,N_1442,N_1476);
xor U4426 (N_4426,N_1746,N_132);
nor U4427 (N_4427,N_776,N_1924);
or U4428 (N_4428,N_1378,N_489);
nor U4429 (N_4429,N_1085,N_875);
xnor U4430 (N_4430,N_866,N_1610);
nor U4431 (N_4431,N_2047,N_687);
or U4432 (N_4432,N_884,N_2495);
nand U4433 (N_4433,N_1501,N_2290);
or U4434 (N_4434,N_572,N_997);
xnor U4435 (N_4435,N_1345,N_930);
nor U4436 (N_4436,N_1914,N_612);
nand U4437 (N_4437,N_1919,N_2081);
xor U4438 (N_4438,N_112,N_817);
nand U4439 (N_4439,N_1500,N_1213);
or U4440 (N_4440,N_1725,N_2175);
xor U4441 (N_4441,N_539,N_1765);
nor U4442 (N_4442,N_342,N_1628);
nor U4443 (N_4443,N_1300,N_1191);
nor U4444 (N_4444,N_1204,N_230);
or U4445 (N_4445,N_1667,N_2156);
nor U4446 (N_4446,N_1960,N_1645);
nand U4447 (N_4447,N_480,N_1106);
and U4448 (N_4448,N_1517,N_1146);
xor U4449 (N_4449,N_2433,N_2430);
and U4450 (N_4450,N_2303,N_852);
nand U4451 (N_4451,N_483,N_789);
nand U4452 (N_4452,N_763,N_2177);
xnor U4453 (N_4453,N_1371,N_2112);
xor U4454 (N_4454,N_2132,N_1528);
and U4455 (N_4455,N_443,N_2059);
xor U4456 (N_4456,N_635,N_18);
and U4457 (N_4457,N_925,N_1468);
xnor U4458 (N_4458,N_1490,N_704);
nand U4459 (N_4459,N_2412,N_406);
nand U4460 (N_4460,N_1537,N_2109);
or U4461 (N_4461,N_2488,N_504);
and U4462 (N_4462,N_2216,N_1019);
nor U4463 (N_4463,N_645,N_2491);
nand U4464 (N_4464,N_2062,N_2014);
nand U4465 (N_4465,N_1871,N_652);
nor U4466 (N_4466,N_768,N_1716);
nand U4467 (N_4467,N_1201,N_2470);
xnor U4468 (N_4468,N_2384,N_500);
or U4469 (N_4469,N_2173,N_2406);
nand U4470 (N_4470,N_392,N_1856);
nor U4471 (N_4471,N_551,N_455);
or U4472 (N_4472,N_1768,N_1793);
nand U4473 (N_4473,N_890,N_1697);
nor U4474 (N_4474,N_2237,N_644);
and U4475 (N_4475,N_2113,N_1088);
xor U4476 (N_4476,N_1524,N_496);
nor U4477 (N_4477,N_911,N_1071);
nand U4478 (N_4478,N_151,N_801);
xnor U4479 (N_4479,N_1885,N_1090);
or U4480 (N_4480,N_2309,N_2257);
and U4481 (N_4481,N_1308,N_15);
and U4482 (N_4482,N_2363,N_1991);
nand U4483 (N_4483,N_2145,N_2255);
and U4484 (N_4484,N_2258,N_2169);
nand U4485 (N_4485,N_1300,N_942);
nor U4486 (N_4486,N_569,N_714);
nand U4487 (N_4487,N_2449,N_1186);
and U4488 (N_4488,N_54,N_133);
nor U4489 (N_4489,N_400,N_2184);
nor U4490 (N_4490,N_2099,N_350);
and U4491 (N_4491,N_1656,N_2352);
nor U4492 (N_4492,N_2119,N_212);
and U4493 (N_4493,N_1092,N_571);
xor U4494 (N_4494,N_686,N_1757);
nand U4495 (N_4495,N_2442,N_2384);
or U4496 (N_4496,N_1646,N_1504);
or U4497 (N_4497,N_1824,N_78);
nand U4498 (N_4498,N_1633,N_2098);
nand U4499 (N_4499,N_124,N_901);
nand U4500 (N_4500,N_2128,N_1131);
nand U4501 (N_4501,N_1382,N_2387);
and U4502 (N_4502,N_1501,N_1395);
and U4503 (N_4503,N_1238,N_778);
xor U4504 (N_4504,N_595,N_2092);
nor U4505 (N_4505,N_2150,N_594);
and U4506 (N_4506,N_106,N_1145);
nand U4507 (N_4507,N_2156,N_1874);
nand U4508 (N_4508,N_926,N_1039);
or U4509 (N_4509,N_2190,N_2142);
xor U4510 (N_4510,N_1404,N_2094);
or U4511 (N_4511,N_157,N_2045);
and U4512 (N_4512,N_34,N_2343);
xor U4513 (N_4513,N_391,N_2163);
and U4514 (N_4514,N_1063,N_1821);
nand U4515 (N_4515,N_2148,N_1939);
or U4516 (N_4516,N_1977,N_1305);
and U4517 (N_4517,N_1315,N_1598);
xor U4518 (N_4518,N_711,N_1037);
and U4519 (N_4519,N_1167,N_1298);
or U4520 (N_4520,N_22,N_1508);
xor U4521 (N_4521,N_2319,N_2484);
nand U4522 (N_4522,N_2034,N_24);
or U4523 (N_4523,N_1268,N_2483);
xor U4524 (N_4524,N_375,N_257);
xnor U4525 (N_4525,N_2085,N_2325);
or U4526 (N_4526,N_815,N_818);
nor U4527 (N_4527,N_183,N_502);
and U4528 (N_4528,N_1492,N_1383);
or U4529 (N_4529,N_2361,N_499);
or U4530 (N_4530,N_880,N_105);
xor U4531 (N_4531,N_340,N_1137);
xor U4532 (N_4532,N_1812,N_2029);
nor U4533 (N_4533,N_1035,N_1863);
nand U4534 (N_4534,N_1467,N_1981);
and U4535 (N_4535,N_1616,N_741);
and U4536 (N_4536,N_746,N_2329);
nand U4537 (N_4537,N_558,N_777);
nor U4538 (N_4538,N_757,N_1837);
xor U4539 (N_4539,N_360,N_1609);
or U4540 (N_4540,N_1497,N_1139);
nand U4541 (N_4541,N_984,N_525);
nor U4542 (N_4542,N_222,N_1542);
nor U4543 (N_4543,N_1936,N_1102);
and U4544 (N_4544,N_2329,N_109);
xnor U4545 (N_4545,N_1293,N_2433);
xor U4546 (N_4546,N_2166,N_1469);
or U4547 (N_4547,N_527,N_1498);
nor U4548 (N_4548,N_2023,N_1307);
nand U4549 (N_4549,N_1861,N_2342);
and U4550 (N_4550,N_422,N_1530);
and U4551 (N_4551,N_2084,N_372);
nand U4552 (N_4552,N_1722,N_460);
xor U4553 (N_4553,N_424,N_2188);
nor U4554 (N_4554,N_317,N_393);
xor U4555 (N_4555,N_338,N_170);
xnor U4556 (N_4556,N_502,N_712);
and U4557 (N_4557,N_1146,N_1003);
and U4558 (N_4558,N_2258,N_1295);
nand U4559 (N_4559,N_955,N_1545);
xnor U4560 (N_4560,N_2044,N_2060);
or U4561 (N_4561,N_895,N_1484);
nor U4562 (N_4562,N_1924,N_2098);
and U4563 (N_4563,N_940,N_1436);
and U4564 (N_4564,N_1702,N_2047);
or U4565 (N_4565,N_477,N_1189);
and U4566 (N_4566,N_1905,N_679);
nand U4567 (N_4567,N_114,N_780);
and U4568 (N_4568,N_1175,N_1012);
nand U4569 (N_4569,N_1527,N_2041);
nand U4570 (N_4570,N_843,N_13);
and U4571 (N_4571,N_567,N_473);
nand U4572 (N_4572,N_1353,N_1450);
xnor U4573 (N_4573,N_2339,N_1427);
nand U4574 (N_4574,N_494,N_93);
xnor U4575 (N_4575,N_1566,N_601);
nand U4576 (N_4576,N_1971,N_767);
nor U4577 (N_4577,N_1988,N_940);
and U4578 (N_4578,N_2129,N_270);
and U4579 (N_4579,N_1764,N_2194);
and U4580 (N_4580,N_1981,N_1805);
xnor U4581 (N_4581,N_2041,N_42);
xor U4582 (N_4582,N_1203,N_93);
nor U4583 (N_4583,N_419,N_1453);
nor U4584 (N_4584,N_943,N_1301);
or U4585 (N_4585,N_1056,N_1761);
or U4586 (N_4586,N_559,N_2099);
nand U4587 (N_4587,N_318,N_109);
nand U4588 (N_4588,N_1431,N_71);
and U4589 (N_4589,N_1215,N_1526);
xor U4590 (N_4590,N_48,N_618);
xor U4591 (N_4591,N_887,N_1145);
nand U4592 (N_4592,N_823,N_246);
nand U4593 (N_4593,N_1270,N_1989);
and U4594 (N_4594,N_2019,N_1374);
nand U4595 (N_4595,N_1839,N_1916);
or U4596 (N_4596,N_1712,N_735);
and U4597 (N_4597,N_2087,N_64);
nand U4598 (N_4598,N_2499,N_1412);
nand U4599 (N_4599,N_445,N_2340);
nor U4600 (N_4600,N_754,N_631);
nor U4601 (N_4601,N_876,N_558);
nand U4602 (N_4602,N_559,N_2257);
xnor U4603 (N_4603,N_2142,N_1689);
nand U4604 (N_4604,N_650,N_145);
xnor U4605 (N_4605,N_1184,N_1719);
nand U4606 (N_4606,N_1868,N_1057);
and U4607 (N_4607,N_2252,N_877);
or U4608 (N_4608,N_1504,N_72);
xnor U4609 (N_4609,N_1035,N_486);
and U4610 (N_4610,N_2274,N_184);
and U4611 (N_4611,N_128,N_2056);
xor U4612 (N_4612,N_1384,N_694);
nand U4613 (N_4613,N_2176,N_678);
xnor U4614 (N_4614,N_2046,N_37);
and U4615 (N_4615,N_2301,N_1589);
nor U4616 (N_4616,N_1736,N_2477);
or U4617 (N_4617,N_40,N_1228);
nor U4618 (N_4618,N_265,N_2177);
xor U4619 (N_4619,N_2012,N_1247);
nor U4620 (N_4620,N_1186,N_1388);
or U4621 (N_4621,N_1143,N_2137);
nand U4622 (N_4622,N_241,N_257);
and U4623 (N_4623,N_1021,N_692);
nand U4624 (N_4624,N_768,N_2202);
nor U4625 (N_4625,N_1333,N_1602);
xor U4626 (N_4626,N_431,N_1362);
and U4627 (N_4627,N_918,N_440);
nor U4628 (N_4628,N_1946,N_1250);
or U4629 (N_4629,N_905,N_677);
xor U4630 (N_4630,N_1861,N_1697);
nor U4631 (N_4631,N_1660,N_1253);
or U4632 (N_4632,N_455,N_2012);
nor U4633 (N_4633,N_1079,N_1757);
nor U4634 (N_4634,N_1346,N_1200);
or U4635 (N_4635,N_873,N_649);
nor U4636 (N_4636,N_2373,N_1254);
or U4637 (N_4637,N_2105,N_606);
and U4638 (N_4638,N_790,N_1230);
nor U4639 (N_4639,N_1436,N_1644);
nor U4640 (N_4640,N_1628,N_1437);
nand U4641 (N_4641,N_2479,N_1067);
nand U4642 (N_4642,N_2174,N_609);
and U4643 (N_4643,N_2468,N_2216);
nand U4644 (N_4644,N_126,N_1057);
nand U4645 (N_4645,N_2139,N_588);
and U4646 (N_4646,N_549,N_515);
or U4647 (N_4647,N_91,N_799);
or U4648 (N_4648,N_1783,N_441);
or U4649 (N_4649,N_66,N_1281);
and U4650 (N_4650,N_1573,N_1617);
or U4651 (N_4651,N_1910,N_611);
and U4652 (N_4652,N_1593,N_1139);
and U4653 (N_4653,N_512,N_2050);
or U4654 (N_4654,N_642,N_648);
nand U4655 (N_4655,N_1515,N_396);
or U4656 (N_4656,N_823,N_1226);
nor U4657 (N_4657,N_792,N_1196);
nor U4658 (N_4658,N_2462,N_401);
and U4659 (N_4659,N_1372,N_1388);
xor U4660 (N_4660,N_1229,N_892);
xor U4661 (N_4661,N_221,N_983);
xnor U4662 (N_4662,N_1881,N_980);
xnor U4663 (N_4663,N_1343,N_2349);
nand U4664 (N_4664,N_238,N_1457);
nor U4665 (N_4665,N_1521,N_420);
or U4666 (N_4666,N_215,N_471);
or U4667 (N_4667,N_880,N_2);
nand U4668 (N_4668,N_1076,N_2217);
nand U4669 (N_4669,N_1601,N_1373);
nand U4670 (N_4670,N_1690,N_2478);
nor U4671 (N_4671,N_1346,N_1639);
nand U4672 (N_4672,N_674,N_1215);
xnor U4673 (N_4673,N_435,N_851);
nor U4674 (N_4674,N_698,N_152);
xor U4675 (N_4675,N_1151,N_173);
nor U4676 (N_4676,N_2062,N_2006);
and U4677 (N_4677,N_1238,N_945);
and U4678 (N_4678,N_376,N_1769);
and U4679 (N_4679,N_1385,N_2251);
and U4680 (N_4680,N_553,N_1075);
and U4681 (N_4681,N_2272,N_600);
and U4682 (N_4682,N_1339,N_971);
or U4683 (N_4683,N_1597,N_1785);
and U4684 (N_4684,N_716,N_7);
or U4685 (N_4685,N_1445,N_149);
nor U4686 (N_4686,N_1664,N_63);
nor U4687 (N_4687,N_2132,N_957);
xor U4688 (N_4688,N_1286,N_1366);
or U4689 (N_4689,N_843,N_185);
nor U4690 (N_4690,N_491,N_113);
or U4691 (N_4691,N_259,N_1343);
nand U4692 (N_4692,N_1683,N_1605);
xor U4693 (N_4693,N_1073,N_610);
and U4694 (N_4694,N_1840,N_2392);
xor U4695 (N_4695,N_2102,N_1461);
nor U4696 (N_4696,N_416,N_1703);
nand U4697 (N_4697,N_1735,N_1844);
and U4698 (N_4698,N_1324,N_2305);
nand U4699 (N_4699,N_1147,N_675);
xnor U4700 (N_4700,N_2231,N_647);
nand U4701 (N_4701,N_1764,N_1016);
or U4702 (N_4702,N_2440,N_1345);
nand U4703 (N_4703,N_211,N_76);
nor U4704 (N_4704,N_1559,N_2049);
xor U4705 (N_4705,N_2166,N_647);
and U4706 (N_4706,N_2395,N_2298);
nand U4707 (N_4707,N_1604,N_1540);
nand U4708 (N_4708,N_1428,N_2214);
xor U4709 (N_4709,N_1831,N_2242);
nand U4710 (N_4710,N_620,N_471);
and U4711 (N_4711,N_1819,N_803);
and U4712 (N_4712,N_2470,N_807);
or U4713 (N_4713,N_1135,N_747);
nand U4714 (N_4714,N_2270,N_1767);
or U4715 (N_4715,N_2082,N_1061);
or U4716 (N_4716,N_1127,N_1738);
nor U4717 (N_4717,N_2228,N_594);
xnor U4718 (N_4718,N_1599,N_511);
xnor U4719 (N_4719,N_1155,N_917);
and U4720 (N_4720,N_287,N_541);
and U4721 (N_4721,N_2044,N_1407);
nor U4722 (N_4722,N_892,N_595);
nand U4723 (N_4723,N_804,N_1784);
nand U4724 (N_4724,N_2226,N_986);
xor U4725 (N_4725,N_2287,N_1940);
and U4726 (N_4726,N_444,N_2140);
xor U4727 (N_4727,N_1001,N_453);
xor U4728 (N_4728,N_107,N_84);
or U4729 (N_4729,N_859,N_1555);
and U4730 (N_4730,N_957,N_601);
nor U4731 (N_4731,N_1617,N_1937);
or U4732 (N_4732,N_901,N_1173);
and U4733 (N_4733,N_800,N_1908);
xnor U4734 (N_4734,N_798,N_1336);
nand U4735 (N_4735,N_1671,N_2031);
nand U4736 (N_4736,N_1078,N_2328);
xnor U4737 (N_4737,N_1360,N_1861);
and U4738 (N_4738,N_1863,N_2338);
or U4739 (N_4739,N_767,N_1608);
nand U4740 (N_4740,N_2179,N_2475);
and U4741 (N_4741,N_798,N_55);
and U4742 (N_4742,N_1235,N_1646);
nor U4743 (N_4743,N_2314,N_1595);
nor U4744 (N_4744,N_443,N_1562);
nand U4745 (N_4745,N_299,N_1015);
nor U4746 (N_4746,N_928,N_941);
and U4747 (N_4747,N_1094,N_1276);
xor U4748 (N_4748,N_1481,N_2304);
and U4749 (N_4749,N_1151,N_2378);
or U4750 (N_4750,N_2271,N_784);
nor U4751 (N_4751,N_1381,N_1546);
or U4752 (N_4752,N_282,N_963);
or U4753 (N_4753,N_1141,N_564);
xnor U4754 (N_4754,N_26,N_675);
or U4755 (N_4755,N_1870,N_1376);
nand U4756 (N_4756,N_1604,N_529);
or U4757 (N_4757,N_1995,N_471);
xor U4758 (N_4758,N_1554,N_539);
nand U4759 (N_4759,N_610,N_982);
xnor U4760 (N_4760,N_295,N_441);
and U4761 (N_4761,N_1465,N_1846);
xnor U4762 (N_4762,N_446,N_1040);
and U4763 (N_4763,N_2165,N_2299);
xnor U4764 (N_4764,N_151,N_570);
nor U4765 (N_4765,N_1892,N_1475);
xnor U4766 (N_4766,N_1882,N_473);
nand U4767 (N_4767,N_2486,N_628);
nand U4768 (N_4768,N_1390,N_1688);
nor U4769 (N_4769,N_2165,N_897);
nor U4770 (N_4770,N_1456,N_383);
or U4771 (N_4771,N_1912,N_1420);
and U4772 (N_4772,N_1232,N_894);
xnor U4773 (N_4773,N_100,N_604);
and U4774 (N_4774,N_187,N_2427);
and U4775 (N_4775,N_842,N_252);
nor U4776 (N_4776,N_1499,N_1629);
xnor U4777 (N_4777,N_828,N_1907);
xnor U4778 (N_4778,N_2332,N_223);
or U4779 (N_4779,N_2025,N_674);
xor U4780 (N_4780,N_746,N_1567);
or U4781 (N_4781,N_114,N_1717);
nor U4782 (N_4782,N_343,N_1163);
and U4783 (N_4783,N_593,N_2446);
xor U4784 (N_4784,N_1602,N_2109);
and U4785 (N_4785,N_245,N_222);
and U4786 (N_4786,N_1810,N_1725);
nor U4787 (N_4787,N_1277,N_2136);
and U4788 (N_4788,N_2072,N_2066);
or U4789 (N_4789,N_1040,N_582);
nand U4790 (N_4790,N_2081,N_226);
xor U4791 (N_4791,N_241,N_619);
nand U4792 (N_4792,N_923,N_1743);
and U4793 (N_4793,N_2295,N_1254);
and U4794 (N_4794,N_994,N_1666);
or U4795 (N_4795,N_2253,N_2293);
or U4796 (N_4796,N_804,N_687);
nor U4797 (N_4797,N_556,N_721);
and U4798 (N_4798,N_1764,N_1200);
xnor U4799 (N_4799,N_140,N_1480);
nor U4800 (N_4800,N_601,N_127);
xnor U4801 (N_4801,N_1679,N_787);
nand U4802 (N_4802,N_974,N_1405);
nor U4803 (N_4803,N_114,N_1547);
nor U4804 (N_4804,N_579,N_508);
nand U4805 (N_4805,N_2019,N_1517);
and U4806 (N_4806,N_466,N_1818);
xnor U4807 (N_4807,N_166,N_1109);
or U4808 (N_4808,N_371,N_2080);
and U4809 (N_4809,N_611,N_1616);
and U4810 (N_4810,N_2269,N_1250);
and U4811 (N_4811,N_1995,N_2489);
and U4812 (N_4812,N_1937,N_1037);
nand U4813 (N_4813,N_693,N_825);
xor U4814 (N_4814,N_85,N_1491);
xor U4815 (N_4815,N_1965,N_1590);
or U4816 (N_4816,N_935,N_1551);
nand U4817 (N_4817,N_1751,N_2255);
xor U4818 (N_4818,N_152,N_1069);
nor U4819 (N_4819,N_603,N_2013);
nand U4820 (N_4820,N_1191,N_34);
or U4821 (N_4821,N_629,N_987);
and U4822 (N_4822,N_403,N_2367);
nand U4823 (N_4823,N_1175,N_1174);
and U4824 (N_4824,N_1033,N_496);
or U4825 (N_4825,N_459,N_583);
and U4826 (N_4826,N_458,N_398);
nand U4827 (N_4827,N_1322,N_419);
nor U4828 (N_4828,N_137,N_2317);
nor U4829 (N_4829,N_2077,N_2091);
and U4830 (N_4830,N_173,N_2160);
or U4831 (N_4831,N_2147,N_1899);
nor U4832 (N_4832,N_1544,N_369);
nand U4833 (N_4833,N_28,N_1703);
nor U4834 (N_4834,N_2064,N_2273);
and U4835 (N_4835,N_1237,N_2465);
and U4836 (N_4836,N_1231,N_2085);
nor U4837 (N_4837,N_214,N_967);
or U4838 (N_4838,N_1996,N_2394);
and U4839 (N_4839,N_334,N_2377);
nand U4840 (N_4840,N_122,N_1320);
and U4841 (N_4841,N_1355,N_1758);
xnor U4842 (N_4842,N_1659,N_274);
nand U4843 (N_4843,N_1700,N_2084);
nor U4844 (N_4844,N_1500,N_2150);
or U4845 (N_4845,N_1820,N_1647);
and U4846 (N_4846,N_1126,N_1554);
and U4847 (N_4847,N_1813,N_186);
nor U4848 (N_4848,N_454,N_1674);
and U4849 (N_4849,N_341,N_834);
nor U4850 (N_4850,N_840,N_346);
nor U4851 (N_4851,N_806,N_256);
xor U4852 (N_4852,N_1558,N_2439);
nor U4853 (N_4853,N_246,N_2013);
nor U4854 (N_4854,N_1417,N_2099);
nand U4855 (N_4855,N_2165,N_979);
xnor U4856 (N_4856,N_569,N_1365);
nor U4857 (N_4857,N_130,N_2458);
xnor U4858 (N_4858,N_442,N_899);
nand U4859 (N_4859,N_817,N_1013);
or U4860 (N_4860,N_1661,N_35);
and U4861 (N_4861,N_2017,N_1392);
nor U4862 (N_4862,N_1544,N_49);
or U4863 (N_4863,N_2082,N_2229);
nand U4864 (N_4864,N_1182,N_2310);
nand U4865 (N_4865,N_195,N_657);
nand U4866 (N_4866,N_1851,N_156);
xor U4867 (N_4867,N_276,N_669);
and U4868 (N_4868,N_1344,N_1793);
and U4869 (N_4869,N_1301,N_2163);
or U4870 (N_4870,N_166,N_2005);
xor U4871 (N_4871,N_651,N_1418);
xnor U4872 (N_4872,N_1000,N_1065);
and U4873 (N_4873,N_1399,N_578);
and U4874 (N_4874,N_870,N_1946);
or U4875 (N_4875,N_2284,N_1085);
nor U4876 (N_4876,N_120,N_878);
nand U4877 (N_4877,N_377,N_64);
or U4878 (N_4878,N_2214,N_1842);
nand U4879 (N_4879,N_1596,N_1714);
nand U4880 (N_4880,N_1392,N_2076);
or U4881 (N_4881,N_2301,N_1182);
xor U4882 (N_4882,N_171,N_1964);
and U4883 (N_4883,N_1791,N_133);
and U4884 (N_4884,N_446,N_310);
nand U4885 (N_4885,N_87,N_531);
nand U4886 (N_4886,N_2052,N_1948);
xnor U4887 (N_4887,N_245,N_1190);
xnor U4888 (N_4888,N_110,N_940);
nor U4889 (N_4889,N_10,N_788);
and U4890 (N_4890,N_2289,N_1322);
and U4891 (N_4891,N_88,N_413);
xor U4892 (N_4892,N_1101,N_152);
nand U4893 (N_4893,N_1815,N_724);
nand U4894 (N_4894,N_2212,N_1845);
or U4895 (N_4895,N_46,N_1982);
or U4896 (N_4896,N_664,N_2423);
nor U4897 (N_4897,N_1844,N_932);
nand U4898 (N_4898,N_1240,N_1398);
nand U4899 (N_4899,N_157,N_1402);
nand U4900 (N_4900,N_1450,N_2288);
or U4901 (N_4901,N_506,N_269);
or U4902 (N_4902,N_195,N_1082);
xor U4903 (N_4903,N_2218,N_408);
and U4904 (N_4904,N_1235,N_2227);
and U4905 (N_4905,N_1005,N_804);
nor U4906 (N_4906,N_360,N_1054);
nor U4907 (N_4907,N_423,N_429);
nor U4908 (N_4908,N_1610,N_873);
xor U4909 (N_4909,N_58,N_1358);
nor U4910 (N_4910,N_945,N_1708);
nor U4911 (N_4911,N_1518,N_1043);
xor U4912 (N_4912,N_1118,N_748);
nor U4913 (N_4913,N_810,N_614);
xor U4914 (N_4914,N_1003,N_1694);
nor U4915 (N_4915,N_2428,N_1693);
or U4916 (N_4916,N_12,N_2057);
nor U4917 (N_4917,N_80,N_96);
nor U4918 (N_4918,N_231,N_909);
or U4919 (N_4919,N_2217,N_54);
nor U4920 (N_4920,N_402,N_269);
xnor U4921 (N_4921,N_633,N_992);
and U4922 (N_4922,N_2473,N_1553);
and U4923 (N_4923,N_802,N_1051);
or U4924 (N_4924,N_492,N_1291);
nand U4925 (N_4925,N_644,N_1594);
or U4926 (N_4926,N_503,N_1919);
xor U4927 (N_4927,N_53,N_1603);
or U4928 (N_4928,N_1844,N_243);
and U4929 (N_4929,N_1970,N_693);
and U4930 (N_4930,N_2303,N_180);
nor U4931 (N_4931,N_2145,N_1017);
and U4932 (N_4932,N_229,N_1725);
or U4933 (N_4933,N_938,N_2155);
nor U4934 (N_4934,N_1409,N_343);
nand U4935 (N_4935,N_1,N_2170);
nand U4936 (N_4936,N_265,N_2217);
and U4937 (N_4937,N_333,N_1530);
xnor U4938 (N_4938,N_118,N_78);
and U4939 (N_4939,N_1976,N_936);
nand U4940 (N_4940,N_1811,N_2198);
nor U4941 (N_4941,N_1780,N_144);
nor U4942 (N_4942,N_1055,N_836);
nor U4943 (N_4943,N_244,N_1251);
xnor U4944 (N_4944,N_822,N_2253);
xnor U4945 (N_4945,N_835,N_1209);
and U4946 (N_4946,N_2085,N_92);
or U4947 (N_4947,N_1775,N_45);
nand U4948 (N_4948,N_1199,N_1460);
nand U4949 (N_4949,N_1928,N_2494);
nor U4950 (N_4950,N_419,N_237);
nand U4951 (N_4951,N_1869,N_2491);
nand U4952 (N_4952,N_1286,N_1620);
nand U4953 (N_4953,N_1958,N_789);
nor U4954 (N_4954,N_567,N_1265);
nand U4955 (N_4955,N_921,N_2153);
and U4956 (N_4956,N_688,N_2189);
nand U4957 (N_4957,N_1268,N_905);
or U4958 (N_4958,N_1035,N_910);
nand U4959 (N_4959,N_386,N_1783);
and U4960 (N_4960,N_2499,N_666);
and U4961 (N_4961,N_2084,N_1554);
or U4962 (N_4962,N_1562,N_1463);
and U4963 (N_4963,N_920,N_1289);
xor U4964 (N_4964,N_643,N_2114);
nand U4965 (N_4965,N_1691,N_2499);
nand U4966 (N_4966,N_608,N_2323);
nor U4967 (N_4967,N_387,N_2304);
and U4968 (N_4968,N_355,N_2251);
and U4969 (N_4969,N_490,N_1182);
nand U4970 (N_4970,N_671,N_2035);
nor U4971 (N_4971,N_1296,N_1151);
and U4972 (N_4972,N_1985,N_1667);
and U4973 (N_4973,N_1620,N_288);
xnor U4974 (N_4974,N_172,N_2012);
xor U4975 (N_4975,N_999,N_1902);
nor U4976 (N_4976,N_1681,N_2073);
nand U4977 (N_4977,N_645,N_1235);
xnor U4978 (N_4978,N_2099,N_2045);
nor U4979 (N_4979,N_941,N_214);
nand U4980 (N_4980,N_1871,N_753);
or U4981 (N_4981,N_309,N_1839);
nand U4982 (N_4982,N_2192,N_240);
nand U4983 (N_4983,N_644,N_384);
nand U4984 (N_4984,N_2116,N_1548);
xor U4985 (N_4985,N_1121,N_1423);
and U4986 (N_4986,N_1070,N_1632);
nor U4987 (N_4987,N_1268,N_227);
nor U4988 (N_4988,N_2129,N_2434);
nor U4989 (N_4989,N_254,N_884);
nand U4990 (N_4990,N_581,N_1353);
xor U4991 (N_4991,N_1063,N_930);
and U4992 (N_4992,N_654,N_1442);
and U4993 (N_4993,N_2212,N_2419);
or U4994 (N_4994,N_1747,N_2007);
nor U4995 (N_4995,N_701,N_265);
xnor U4996 (N_4996,N_501,N_255);
xor U4997 (N_4997,N_2117,N_2233);
and U4998 (N_4998,N_1722,N_1437);
nor U4999 (N_4999,N_2203,N_445);
xnor U5000 (N_5000,N_3956,N_2741);
nand U5001 (N_5001,N_3145,N_2671);
or U5002 (N_5002,N_4479,N_4434);
and U5003 (N_5003,N_4999,N_4315);
or U5004 (N_5004,N_3204,N_3497);
and U5005 (N_5005,N_3042,N_3149);
or U5006 (N_5006,N_4218,N_4612);
or U5007 (N_5007,N_4905,N_2724);
and U5008 (N_5008,N_4445,N_2949);
or U5009 (N_5009,N_3669,N_4217);
nand U5010 (N_5010,N_2532,N_3107);
xor U5011 (N_5011,N_3033,N_2934);
and U5012 (N_5012,N_4356,N_3783);
nor U5013 (N_5013,N_4990,N_4478);
and U5014 (N_5014,N_4875,N_3993);
or U5015 (N_5015,N_4524,N_2789);
or U5016 (N_5016,N_3231,N_3096);
nor U5017 (N_5017,N_2810,N_4673);
or U5018 (N_5018,N_4930,N_2831);
xnor U5019 (N_5019,N_2749,N_4614);
or U5020 (N_5020,N_3892,N_2933);
nor U5021 (N_5021,N_3934,N_3561);
xnor U5022 (N_5022,N_3282,N_4362);
and U5023 (N_5023,N_4343,N_3525);
and U5024 (N_5024,N_3379,N_4628);
nor U5025 (N_5025,N_4283,N_4661);
nand U5026 (N_5026,N_4163,N_3472);
nand U5027 (N_5027,N_4937,N_4371);
xor U5028 (N_5028,N_4507,N_2552);
or U5029 (N_5029,N_2726,N_3110);
xor U5030 (N_5030,N_4592,N_2969);
nand U5031 (N_5031,N_3015,N_2911);
nand U5032 (N_5032,N_4108,N_2594);
and U5033 (N_5033,N_2694,N_3404);
and U5034 (N_5034,N_4641,N_2672);
nand U5035 (N_5035,N_2589,N_2889);
nand U5036 (N_5036,N_3461,N_3513);
xor U5037 (N_5037,N_4494,N_4794);
nor U5038 (N_5038,N_4901,N_2835);
xor U5039 (N_5039,N_4327,N_3467);
nor U5040 (N_5040,N_4448,N_3400);
and U5041 (N_5041,N_2982,N_3364);
nand U5042 (N_5042,N_4307,N_2579);
nand U5043 (N_5043,N_4765,N_3428);
nor U5044 (N_5044,N_2992,N_2971);
nor U5045 (N_5045,N_2972,N_3061);
nand U5046 (N_5046,N_2799,N_3920);
or U5047 (N_5047,N_4138,N_2998);
xor U5048 (N_5048,N_3703,N_4897);
xor U5049 (N_5049,N_2800,N_4469);
xnor U5050 (N_5050,N_2605,N_4426);
and U5051 (N_5051,N_4211,N_2941);
or U5052 (N_5052,N_4646,N_2687);
and U5053 (N_5053,N_3658,N_4586);
or U5054 (N_5054,N_3209,N_3849);
and U5055 (N_5055,N_4702,N_4121);
nand U5056 (N_5056,N_4926,N_4314);
or U5057 (N_5057,N_2868,N_3770);
nor U5058 (N_5058,N_4397,N_3190);
or U5059 (N_5059,N_3049,N_2565);
and U5060 (N_5060,N_4459,N_2660);
and U5061 (N_5061,N_4944,N_3531);
or U5062 (N_5062,N_3242,N_4969);
nor U5063 (N_5063,N_3548,N_4219);
xnor U5064 (N_5064,N_4373,N_4255);
xor U5065 (N_5065,N_4609,N_2519);
or U5066 (N_5066,N_4210,N_2878);
nor U5067 (N_5067,N_3429,N_3225);
nand U5068 (N_5068,N_3763,N_4579);
nor U5069 (N_5069,N_4348,N_3581);
nor U5070 (N_5070,N_2797,N_3396);
and U5071 (N_5071,N_2711,N_2961);
and U5072 (N_5072,N_4027,N_4569);
and U5073 (N_5073,N_4635,N_4573);
nand U5074 (N_5074,N_2830,N_2935);
nor U5075 (N_5075,N_2955,N_3069);
xnor U5076 (N_5076,N_3269,N_4645);
or U5077 (N_5077,N_3728,N_4410);
or U5078 (N_5078,N_4537,N_2920);
nor U5079 (N_5079,N_4886,N_4328);
and U5080 (N_5080,N_4072,N_4557);
nor U5081 (N_5081,N_3991,N_4487);
and U5082 (N_5082,N_4078,N_4923);
xnor U5083 (N_5083,N_3918,N_4510);
or U5084 (N_5084,N_3504,N_4962);
xnor U5085 (N_5085,N_2960,N_3906);
and U5086 (N_5086,N_4268,N_2567);
nand U5087 (N_5087,N_3311,N_4009);
and U5088 (N_5088,N_4960,N_3682);
or U5089 (N_5089,N_4739,N_2625);
nand U5090 (N_5090,N_4711,N_2836);
nand U5091 (N_5091,N_2699,N_3059);
nand U5092 (N_5092,N_4772,N_3321);
nand U5093 (N_5093,N_2895,N_3651);
or U5094 (N_5094,N_3283,N_3649);
and U5095 (N_5095,N_4617,N_2866);
nand U5096 (N_5096,N_4808,N_2500);
or U5097 (N_5097,N_3772,N_4764);
nand U5098 (N_5098,N_3474,N_3455);
and U5099 (N_5099,N_3541,N_4180);
xnor U5100 (N_5100,N_4892,N_4919);
nand U5101 (N_5101,N_3449,N_4023);
and U5102 (N_5102,N_4848,N_4101);
or U5103 (N_5103,N_4073,N_4413);
xor U5104 (N_5104,N_4908,N_3383);
and U5105 (N_5105,N_3919,N_3961);
xor U5106 (N_5106,N_4452,N_2632);
or U5107 (N_5107,N_3385,N_4753);
nor U5108 (N_5108,N_4607,N_4812);
or U5109 (N_5109,N_3362,N_2582);
and U5110 (N_5110,N_3478,N_2824);
nand U5111 (N_5111,N_3515,N_2675);
nor U5112 (N_5112,N_3071,N_4568);
and U5113 (N_5113,N_4780,N_3861);
nand U5114 (N_5114,N_2839,N_3024);
or U5115 (N_5115,N_4201,N_2502);
and U5116 (N_5116,N_3271,N_3280);
nor U5117 (N_5117,N_4380,N_2544);
and U5118 (N_5118,N_4683,N_3030);
or U5119 (N_5119,N_2788,N_4778);
nor U5120 (N_5120,N_2524,N_4828);
xnor U5121 (N_5121,N_3766,N_4054);
and U5122 (N_5122,N_4040,N_3473);
and U5123 (N_5123,N_4734,N_2898);
nand U5124 (N_5124,N_3664,N_2790);
nand U5125 (N_5125,N_3366,N_3996);
or U5126 (N_5126,N_3980,N_3814);
or U5127 (N_5127,N_2572,N_3045);
nor U5128 (N_5128,N_2883,N_2630);
nor U5129 (N_5129,N_2855,N_4948);
nand U5130 (N_5130,N_2650,N_4925);
nor U5131 (N_5131,N_2867,N_4735);
nand U5132 (N_5132,N_4161,N_3369);
nand U5133 (N_5133,N_4632,N_4625);
nor U5134 (N_5134,N_3141,N_3494);
or U5135 (N_5135,N_2943,N_3538);
and U5136 (N_5136,N_4500,N_4252);
or U5137 (N_5137,N_4706,N_4953);
xnor U5138 (N_5138,N_2617,N_3318);
and U5139 (N_5139,N_4300,N_2522);
or U5140 (N_5140,N_4987,N_4316);
or U5141 (N_5141,N_2718,N_4758);
and U5142 (N_5142,N_3896,N_4643);
nand U5143 (N_5143,N_2608,N_2956);
and U5144 (N_5144,N_3930,N_4081);
nand U5145 (N_5145,N_4552,N_3866);
nor U5146 (N_5146,N_3706,N_2802);
nand U5147 (N_5147,N_3232,N_3983);
and U5148 (N_5148,N_2980,N_4564);
nand U5149 (N_5149,N_4233,N_4025);
nor U5150 (N_5150,N_3674,N_3464);
and U5151 (N_5151,N_2588,N_2514);
and U5152 (N_5152,N_4146,N_4486);
nor U5153 (N_5153,N_2592,N_2919);
nor U5154 (N_5154,N_4319,N_4277);
or U5155 (N_5155,N_4680,N_3129);
xor U5156 (N_5156,N_2816,N_3398);
xor U5157 (N_5157,N_3941,N_3089);
nor U5158 (N_5158,N_3559,N_3433);
or U5159 (N_5159,N_3818,N_2740);
or U5160 (N_5160,N_3990,N_4104);
xnor U5161 (N_5161,N_4384,N_4869);
nor U5162 (N_5162,N_3493,N_4427);
xnor U5163 (N_5163,N_4057,N_3079);
nor U5164 (N_5164,N_2783,N_3431);
or U5165 (N_5165,N_2606,N_2778);
or U5166 (N_5166,N_3477,N_3981);
nor U5167 (N_5167,N_3660,N_4446);
and U5168 (N_5168,N_4387,N_4237);
nand U5169 (N_5169,N_4118,N_3838);
or U5170 (N_5170,N_4823,N_3935);
nor U5171 (N_5171,N_4689,N_4119);
xnor U5172 (N_5172,N_3698,N_3900);
or U5173 (N_5173,N_2910,N_4931);
xor U5174 (N_5174,N_4241,N_4405);
and U5175 (N_5175,N_4274,N_4723);
and U5176 (N_5176,N_4276,N_2758);
nand U5177 (N_5177,N_4726,N_3953);
nor U5178 (N_5178,N_3816,N_4326);
or U5179 (N_5179,N_3829,N_4621);
nand U5180 (N_5180,N_2786,N_4800);
nor U5181 (N_5181,N_2593,N_4199);
nor U5182 (N_5182,N_4587,N_3987);
nand U5183 (N_5183,N_3685,N_4705);
nor U5184 (N_5184,N_4728,N_3593);
or U5185 (N_5185,N_3267,N_3960);
xnor U5186 (N_5186,N_2604,N_4456);
xor U5187 (N_5187,N_4333,N_4016);
or U5188 (N_5188,N_3744,N_4257);
nor U5189 (N_5189,N_2653,N_3874);
or U5190 (N_5190,N_3249,N_4109);
xnor U5191 (N_5191,N_3457,N_4549);
nor U5192 (N_5192,N_2813,N_4667);
nor U5193 (N_5193,N_3454,N_3540);
nor U5194 (N_5194,N_3533,N_4350);
nor U5195 (N_5195,N_3147,N_3725);
xnor U5196 (N_5196,N_4790,N_4022);
or U5197 (N_5197,N_4822,N_2622);
xnor U5198 (N_5198,N_2663,N_3647);
nand U5199 (N_5199,N_2882,N_3140);
xnor U5200 (N_5200,N_2781,N_4291);
nand U5201 (N_5201,N_3786,N_3088);
xor U5202 (N_5202,N_4499,N_4653);
nand U5203 (N_5203,N_3543,N_3572);
xnor U5204 (N_5204,N_4001,N_4911);
or U5205 (N_5205,N_4658,N_4660);
nand U5206 (N_5206,N_3388,N_4866);
xnor U5207 (N_5207,N_2766,N_3169);
nor U5208 (N_5208,N_4857,N_4142);
nor U5209 (N_5209,N_3914,N_3436);
nand U5210 (N_5210,N_4697,N_4256);
xnor U5211 (N_5211,N_3797,N_3005);
nand U5212 (N_5212,N_3729,N_3508);
and U5213 (N_5213,N_2569,N_4884);
or U5214 (N_5214,N_4872,N_3211);
nand U5215 (N_5215,N_4150,N_3569);
nor U5216 (N_5216,N_2837,N_2966);
nand U5217 (N_5217,N_4228,N_2975);
and U5218 (N_5218,N_4634,N_4484);
nor U5219 (N_5219,N_3985,N_3095);
xnor U5220 (N_5220,N_2794,N_3004);
xnor U5221 (N_5221,N_3189,N_4074);
nand U5222 (N_5222,N_3272,N_4388);
nor U5223 (N_5223,N_4249,N_3387);
nand U5224 (N_5224,N_2570,N_4442);
and U5225 (N_5225,N_4289,N_4732);
and U5226 (N_5226,N_3078,N_4815);
or U5227 (N_5227,N_3812,N_3805);
xor U5228 (N_5228,N_4725,N_2750);
nor U5229 (N_5229,N_2994,N_3998);
xnor U5230 (N_5230,N_4224,N_4605);
nand U5231 (N_5231,N_2731,N_4584);
nand U5232 (N_5232,N_4311,N_4203);
or U5233 (N_5233,N_4803,N_2964);
xor U5234 (N_5234,N_3828,N_3687);
nand U5235 (N_5235,N_3984,N_3306);
xor U5236 (N_5236,N_2550,N_3488);
xor U5237 (N_5237,N_3394,N_4465);
nand U5238 (N_5238,N_4436,N_3689);
nor U5239 (N_5239,N_2525,N_2619);
xor U5240 (N_5240,N_4582,N_3865);
xor U5241 (N_5241,N_4096,N_3066);
or U5242 (N_5242,N_4120,N_2643);
and U5243 (N_5243,N_3928,N_2917);
nand U5244 (N_5244,N_3416,N_2627);
nor U5245 (N_5245,N_3475,N_4796);
nor U5246 (N_5246,N_4451,N_3320);
and U5247 (N_5247,N_3266,N_3135);
xnor U5248 (N_5248,N_2838,N_4981);
or U5249 (N_5249,N_3758,N_2674);
nor U5250 (N_5250,N_4756,N_2859);
and U5251 (N_5251,N_3261,N_2996);
xnor U5252 (N_5252,N_4378,N_4048);
xor U5253 (N_5253,N_3880,N_2747);
and U5254 (N_5254,N_2506,N_2944);
nand U5255 (N_5255,N_3926,N_3380);
nand U5256 (N_5256,N_3695,N_3646);
xor U5257 (N_5257,N_4175,N_4988);
nand U5258 (N_5258,N_2691,N_4793);
nand U5259 (N_5259,N_4966,N_4100);
or U5260 (N_5260,N_3236,N_4135);
and U5261 (N_5261,N_4058,N_4932);
nor U5262 (N_5262,N_2976,N_3372);
nor U5263 (N_5263,N_4019,N_3636);
nor U5264 (N_5264,N_4774,N_3375);
nor U5265 (N_5265,N_4453,N_3281);
nand U5266 (N_5266,N_3331,N_2776);
nor U5267 (N_5267,N_4066,N_4983);
and U5268 (N_5268,N_3679,N_3127);
nand U5269 (N_5269,N_4795,N_4585);
xnor U5270 (N_5270,N_3847,N_4460);
and U5271 (N_5271,N_4916,N_4782);
or U5272 (N_5272,N_4320,N_4128);
or U5273 (N_5273,N_4766,N_4712);
nand U5274 (N_5274,N_4084,N_4090);
and U5275 (N_5275,N_4671,N_3684);
or U5276 (N_5276,N_4659,N_3344);
nor U5277 (N_5277,N_4532,N_2530);
and U5278 (N_5278,N_3518,N_3507);
and U5279 (N_5279,N_4438,N_2730);
or U5280 (N_5280,N_4391,N_3046);
or U5281 (N_5281,N_3670,N_3026);
nand U5282 (N_5282,N_2598,N_3512);
xnor U5283 (N_5283,N_4489,N_3622);
nor U5284 (N_5284,N_3313,N_4724);
and U5285 (N_5285,N_4721,N_3459);
xor U5286 (N_5286,N_3090,N_4535);
or U5287 (N_5287,N_3598,N_3999);
or U5288 (N_5288,N_4745,N_3997);
xnor U5289 (N_5289,N_3378,N_3184);
xnor U5290 (N_5290,N_4703,N_4352);
or U5291 (N_5291,N_3040,N_3133);
or U5292 (N_5292,N_3963,N_3479);
xor U5293 (N_5293,N_2862,N_2990);
nand U5294 (N_5294,N_2967,N_4555);
and U5295 (N_5295,N_2702,N_3946);
and U5296 (N_5296,N_2833,N_4996);
or U5297 (N_5297,N_4622,N_2549);
nand U5298 (N_5298,N_2775,N_4473);
and U5299 (N_5299,N_4949,N_2692);
nand U5300 (N_5300,N_2652,N_3086);
xnor U5301 (N_5301,N_2561,N_2720);
and U5302 (N_5302,N_4106,N_4225);
xor U5303 (N_5303,N_3910,N_2693);
nand U5304 (N_5304,N_2773,N_4443);
nand U5305 (N_5305,N_3823,N_4136);
nand U5306 (N_5306,N_2997,N_3354);
nand U5307 (N_5307,N_4518,N_3099);
nor U5308 (N_5308,N_4692,N_4768);
xnor U5309 (N_5309,N_4825,N_4687);
or U5310 (N_5310,N_2707,N_3709);
nand U5311 (N_5311,N_2849,N_2932);
or U5312 (N_5312,N_3254,N_3315);
nor U5313 (N_5313,N_4860,N_4189);
and U5314 (N_5314,N_4088,N_3060);
nor U5315 (N_5315,N_4519,N_3970);
xor U5316 (N_5316,N_4110,N_4554);
and U5317 (N_5317,N_3864,N_4686);
nor U5318 (N_5318,N_4207,N_3583);
nor U5319 (N_5319,N_3294,N_3530);
and U5320 (N_5320,N_4160,N_3337);
xor U5321 (N_5321,N_3973,N_3314);
or U5322 (N_5322,N_2686,N_2542);
or U5323 (N_5323,N_4964,N_3064);
or U5324 (N_5324,N_3075,N_2658);
or U5325 (N_5325,N_3549,N_4430);
and U5326 (N_5326,N_3050,N_2858);
and U5327 (N_5327,N_3992,N_3460);
nor U5328 (N_5328,N_3959,N_2962);
nor U5329 (N_5329,N_4067,N_4527);
nand U5330 (N_5330,N_3006,N_3853);
and U5331 (N_5331,N_4655,N_2583);
and U5332 (N_5332,N_3811,N_3936);
nor U5333 (N_5333,N_3913,N_4947);
xor U5334 (N_5334,N_4992,N_2755);
nor U5335 (N_5335,N_3542,N_4903);
and U5336 (N_5336,N_4475,N_3869);
xnor U5337 (N_5337,N_3951,N_4046);
nor U5338 (N_5338,N_4385,N_4334);
nor U5339 (N_5339,N_4439,N_2843);
nand U5340 (N_5340,N_2973,N_4701);
or U5341 (N_5341,N_4536,N_2950);
and U5342 (N_5342,N_3343,N_4841);
nor U5343 (N_5343,N_3470,N_2688);
nand U5344 (N_5344,N_3719,N_4624);
nand U5345 (N_5345,N_4381,N_4998);
or U5346 (N_5346,N_2508,N_4253);
xnor U5347 (N_5347,N_2513,N_4239);
xor U5348 (N_5348,N_3017,N_4989);
and U5349 (N_5349,N_4243,N_4458);
and U5350 (N_5350,N_2769,N_4312);
and U5351 (N_5351,N_4457,N_2983);
nor U5352 (N_5352,N_3944,N_3787);
xor U5353 (N_5353,N_3327,N_4377);
xnor U5354 (N_5354,N_4137,N_3007);
nand U5355 (N_5355,N_4595,N_4240);
nand U5356 (N_5356,N_4164,N_4546);
xor U5357 (N_5357,N_3053,N_2556);
or U5358 (N_5358,N_4056,N_4041);
nand U5359 (N_5359,N_3789,N_4797);
xor U5360 (N_5360,N_3820,N_4193);
or U5361 (N_5361,N_3577,N_2659);
nand U5362 (N_5362,N_4275,N_4230);
nor U5363 (N_5363,N_3265,N_3018);
nand U5364 (N_5364,N_2716,N_4008);
nand U5365 (N_5365,N_3368,N_4153);
nor U5366 (N_5366,N_4491,N_4303);
or U5367 (N_5367,N_2979,N_4918);
and U5368 (N_5368,N_3250,N_4294);
xor U5369 (N_5369,N_4053,N_3545);
nand U5370 (N_5370,N_4805,N_4332);
xor U5371 (N_5371,N_3120,N_4205);
or U5372 (N_5372,N_4154,N_3534);
xor U5373 (N_5373,N_3877,N_3841);
and U5374 (N_5374,N_4783,N_4954);
and U5375 (N_5375,N_3589,N_3037);
or U5376 (N_5376,N_3529,N_4995);
and U5377 (N_5377,N_4092,N_4868);
or U5378 (N_5378,N_4375,N_3241);
and U5379 (N_5379,N_2743,N_3203);
xor U5380 (N_5380,N_4238,N_2585);
xnor U5381 (N_5381,N_3904,N_4912);
or U5382 (N_5382,N_3642,N_2640);
and U5383 (N_5383,N_3503,N_4831);
xor U5384 (N_5384,N_2517,N_4824);
or U5385 (N_5385,N_4955,N_2504);
and U5386 (N_5386,N_3384,N_3794);
xnor U5387 (N_5387,N_3633,N_3735);
or U5388 (N_5388,N_2861,N_2842);
and U5389 (N_5389,N_3224,N_4492);
nand U5390 (N_5390,N_4729,N_4047);
nand U5391 (N_5391,N_2577,N_2545);
nand U5392 (N_5392,N_3159,N_4416);
nand U5393 (N_5393,N_2587,N_4619);
nand U5394 (N_5394,N_4364,N_3312);
nand U5395 (N_5395,N_3562,N_4178);
and U5396 (N_5396,N_4418,N_3625);
nand U5397 (N_5397,N_3616,N_3523);
or U5398 (N_5398,N_4222,N_4784);
and U5399 (N_5399,N_2916,N_3898);
and U5400 (N_5400,N_2888,N_3976);
and U5401 (N_5401,N_3938,N_3825);
nand U5402 (N_5402,N_3350,N_4340);
nor U5403 (N_5403,N_4927,N_4907);
and U5404 (N_5404,N_3964,N_3626);
nand U5405 (N_5405,N_2623,N_2558);
and U5406 (N_5406,N_2963,N_3336);
and U5407 (N_5407,N_4490,N_4921);
and U5408 (N_5408,N_4666,N_3764);
and U5409 (N_5409,N_3038,N_4887);
or U5410 (N_5410,N_3044,N_4123);
nor U5411 (N_5411,N_3273,N_3889);
nor U5412 (N_5412,N_4227,N_3937);
xnor U5413 (N_5413,N_3551,N_3391);
nor U5414 (N_5414,N_3422,N_4260);
or U5415 (N_5415,N_4112,N_3346);
nor U5416 (N_5416,N_4080,N_4898);
or U5417 (N_5417,N_3573,N_4130);
nor U5418 (N_5418,N_2828,N_4829);
nor U5419 (N_5419,N_4093,N_2951);
and U5420 (N_5420,N_4415,N_4117);
nor U5421 (N_5421,N_3329,N_4280);
xor U5422 (N_5422,N_3897,N_3335);
nand U5423 (N_5423,N_3305,N_4042);
or U5424 (N_5424,N_4144,N_4681);
and U5425 (N_5425,N_4893,N_4360);
nor U5426 (N_5426,N_3355,N_3844);
or U5427 (N_5427,N_3003,N_4107);
and U5428 (N_5428,N_2526,N_4105);
and U5429 (N_5429,N_4122,N_3367);
or U5430 (N_5430,N_3717,N_3068);
and U5431 (N_5431,N_4447,N_2885);
or U5432 (N_5432,N_4335,N_4917);
nor U5433 (N_5433,N_2708,N_2779);
nand U5434 (N_5434,N_3251,N_4976);
or U5435 (N_5435,N_2746,N_4113);
xor U5436 (N_5436,N_3702,N_3942);
nor U5437 (N_5437,N_2586,N_3048);
nor U5438 (N_5438,N_4615,N_4533);
and U5439 (N_5439,N_3381,N_4888);
and U5440 (N_5440,N_3975,N_2921);
xnor U5441 (N_5441,N_3021,N_3894);
or U5442 (N_5442,N_2760,N_3667);
and U5443 (N_5443,N_3578,N_4836);
or U5444 (N_5444,N_3732,N_3229);
nand U5445 (N_5445,N_3840,N_3317);
xor U5446 (N_5446,N_3087,N_3255);
or U5447 (N_5447,N_3954,N_3776);
or U5448 (N_5448,N_4349,N_2689);
nand U5449 (N_5449,N_4134,N_4678);
and U5450 (N_5450,N_4077,N_4206);
nor U5451 (N_5451,N_2903,N_2841);
xor U5452 (N_5452,N_4337,N_2596);
nor U5453 (N_5453,N_3268,N_3832);
xnor U5454 (N_5454,N_3230,N_3067);
nand U5455 (N_5455,N_4091,N_3704);
nor U5456 (N_5456,N_3219,N_4910);
nand U5457 (N_5457,N_2578,N_2697);
or U5458 (N_5458,N_2808,N_2827);
nor U5459 (N_5459,N_3753,N_4853);
or U5460 (N_5460,N_3167,N_3444);
xnor U5461 (N_5461,N_3752,N_4936);
or U5462 (N_5462,N_3179,N_3610);
and U5463 (N_5463,N_3425,N_4596);
nand U5464 (N_5464,N_4620,N_4834);
or U5465 (N_5465,N_4993,N_4155);
xnor U5466 (N_5466,N_4561,N_2668);
nor U5467 (N_5467,N_4980,N_4742);
xnor U5468 (N_5468,N_3187,N_4299);
xor U5469 (N_5469,N_3966,N_3174);
xor U5470 (N_5470,N_3803,N_3575);
nand U5471 (N_5471,N_4075,N_4059);
xor U5472 (N_5472,N_2677,N_3916);
xnor U5473 (N_5473,N_2854,N_2928);
and U5474 (N_5474,N_3831,N_2533);
and U5475 (N_5475,N_3597,N_2722);
nand U5476 (N_5476,N_3675,N_3256);
and U5477 (N_5477,N_4578,N_4082);
and U5478 (N_5478,N_4179,N_3855);
nand U5479 (N_5479,N_2822,N_3165);
nand U5480 (N_5480,N_3836,N_3032);
nor U5481 (N_5481,N_2865,N_4633);
nor U5482 (N_5482,N_4613,N_3923);
or U5483 (N_5483,N_3223,N_4324);
xnor U5484 (N_5484,N_4608,N_4220);
or U5485 (N_5485,N_4979,N_4719);
or U5486 (N_5486,N_3592,N_2853);
and U5487 (N_5487,N_3138,N_4407);
nand U5488 (N_5488,N_3083,N_3215);
xnor U5489 (N_5489,N_4272,N_2661);
nor U5490 (N_5490,N_4269,N_4344);
xor U5491 (N_5491,N_3481,N_4165);
and U5492 (N_5492,N_3492,N_3392);
nand U5493 (N_5493,N_4736,N_2678);
nand U5494 (N_5494,N_3487,N_3723);
nand U5495 (N_5495,N_4688,N_4971);
and U5496 (N_5496,N_2757,N_4662);
xor U5497 (N_5497,N_4474,N_4235);
nor U5498 (N_5498,N_2712,N_3058);
or U5499 (N_5499,N_4039,N_3274);
or U5500 (N_5500,N_4743,N_2795);
nand U5501 (N_5501,N_4099,N_2629);
xor U5502 (N_5502,N_3289,N_3390);
nand U5503 (N_5503,N_4221,N_4062);
nor U5504 (N_5504,N_4354,N_4773);
nand U5505 (N_5505,N_3057,N_3308);
nor U5506 (N_5506,N_3415,N_2864);
nor U5507 (N_5507,N_3842,N_2559);
or U5508 (N_5508,N_4762,N_4177);
nor U5509 (N_5509,N_2573,N_4977);
or U5510 (N_5510,N_3438,N_2890);
or U5511 (N_5511,N_3476,N_3582);
xnor U5512 (N_5512,N_3374,N_3365);
nor U5513 (N_5513,N_3092,N_2557);
nand U5514 (N_5514,N_3322,N_3419);
or U5515 (N_5515,N_2832,N_4330);
xor U5516 (N_5516,N_3621,N_4367);
nand U5517 (N_5517,N_4351,N_2646);
nand U5518 (N_5518,N_3663,N_3188);
nand U5519 (N_5519,N_3349,N_4064);
or U5520 (N_5520,N_3292,N_3371);
or U5521 (N_5521,N_3253,N_3002);
nand U5522 (N_5522,N_4506,N_2914);
xnor U5523 (N_5523,N_4567,N_3264);
nand U5524 (N_5524,N_2732,N_3631);
nand U5525 (N_5525,N_3287,N_3641);
nor U5526 (N_5526,N_3566,N_4470);
xor U5527 (N_5527,N_2698,N_4583);
nor U5528 (N_5528,N_4406,N_3074);
and U5529 (N_5529,N_4368,N_4158);
and U5530 (N_5530,N_3688,N_4421);
nor U5531 (N_5531,N_4419,N_4631);
nand U5532 (N_5532,N_2682,N_2829);
and U5533 (N_5533,N_2931,N_4279);
xor U5534 (N_5534,N_4755,N_3962);
xnor U5535 (N_5535,N_3862,N_3565);
xnor U5536 (N_5536,N_3686,N_4847);
xnor U5537 (N_5537,N_3259,N_3712);
nor U5538 (N_5538,N_3857,N_3200);
nand U5539 (N_5539,N_3699,N_4696);
and U5540 (N_5540,N_3270,N_4116);
and U5541 (N_5541,N_4139,N_3012);
or U5542 (N_5542,N_4727,N_3263);
and U5543 (N_5543,N_2958,N_4810);
and U5544 (N_5544,N_4412,N_3750);
or U5545 (N_5545,N_2984,N_4896);
and U5546 (N_5546,N_4885,N_4844);
nor U5547 (N_5547,N_4145,N_4601);
or U5548 (N_5548,N_2897,N_4234);
and U5549 (N_5549,N_4485,N_3940);
xor U5550 (N_5550,N_3500,N_4864);
nand U5551 (N_5551,N_3871,N_3304);
nor U5552 (N_5552,N_2551,N_3432);
and U5553 (N_5553,N_2803,N_3197);
nand U5554 (N_5554,N_3103,N_3496);
nor U5555 (N_5555,N_3205,N_3708);
xnor U5556 (N_5556,N_3100,N_2762);
or U5557 (N_5557,N_3157,N_3228);
or U5558 (N_5558,N_3791,N_3466);
or U5559 (N_5559,N_3295,N_3608);
and U5560 (N_5560,N_3891,N_4730);
nand U5561 (N_5561,N_4909,N_4821);
xor U5562 (N_5562,N_3553,N_4775);
nor U5563 (N_5563,N_4306,N_3939);
or U5564 (N_5564,N_4192,N_4867);
nand U5565 (N_5565,N_3690,N_3222);
or U5566 (N_5566,N_3377,N_4604);
nor U5567 (N_5567,N_3325,N_4390);
nor U5568 (N_5568,N_4403,N_3340);
nand U5569 (N_5569,N_3353,N_4920);
xnor U5570 (N_5570,N_4209,N_3453);
or U5571 (N_5571,N_4437,N_2631);
nand U5572 (N_5572,N_2507,N_2834);
and U5573 (N_5573,N_4749,N_4664);
and U5574 (N_5574,N_3645,N_3810);
or U5575 (N_5575,N_3279,N_4176);
or U5576 (N_5576,N_4037,N_3278);
xnor U5577 (N_5577,N_2884,N_3697);
or U5578 (N_5578,N_3155,N_4162);
or U5579 (N_5579,N_4709,N_3546);
and U5580 (N_5580,N_3168,N_4792);
nor U5581 (N_5581,N_3243,N_2723);
xor U5582 (N_5582,N_4677,N_2957);
nor U5583 (N_5583,N_2667,N_2751);
nand U5584 (N_5584,N_2748,N_4036);
and U5585 (N_5585,N_3514,N_3677);
xor U5586 (N_5586,N_3132,N_2923);
nand U5587 (N_5587,N_3440,N_3809);
and U5588 (N_5588,N_4694,N_2767);
and U5589 (N_5589,N_4392,N_4684);
xnor U5590 (N_5590,N_4346,N_4747);
xor U5591 (N_5591,N_2742,N_2785);
and U5592 (N_5592,N_3550,N_3134);
nor U5593 (N_5593,N_3054,N_2793);
and U5594 (N_5594,N_3175,N_2706);
and U5595 (N_5595,N_2942,N_3673);
and U5596 (N_5596,N_2534,N_4400);
nor U5597 (N_5597,N_3678,N_2818);
xor U5598 (N_5598,N_3301,N_2597);
xnor U5599 (N_5599,N_4505,N_4833);
or U5600 (N_5600,N_3574,N_3151);
xor U5601 (N_5601,N_2715,N_3019);
and U5602 (N_5602,N_3290,N_3217);
xor U5603 (N_5603,N_3376,N_3055);
xor U5604 (N_5604,N_2709,N_3348);
nor U5605 (N_5605,N_3931,N_3560);
or U5606 (N_5606,N_3846,N_3212);
and U5607 (N_5607,N_3947,N_3220);
nand U5608 (N_5608,N_4642,N_3208);
or U5609 (N_5609,N_3815,N_4353);
and U5610 (N_5610,N_4501,N_3863);
xor U5611 (N_5611,N_3927,N_4156);
nor U5612 (N_5612,N_3310,N_2805);
xnor U5613 (N_5613,N_2913,N_4504);
or U5614 (N_5614,N_4250,N_4508);
and U5615 (N_5615,N_3620,N_3720);
nor U5616 (N_5616,N_2871,N_4889);
or U5617 (N_5617,N_3591,N_4838);
xnor U5618 (N_5618,N_4763,N_3480);
and U5619 (N_5619,N_4700,N_2621);
nand U5620 (N_5620,N_3644,N_3716);
xor U5621 (N_5621,N_4355,N_4126);
xor U5622 (N_5622,N_4562,N_3393);
or U5623 (N_5623,N_2780,N_4097);
and U5624 (N_5624,N_4710,N_4804);
nand U5625 (N_5625,N_3244,N_4835);
or U5626 (N_5626,N_4802,N_3106);
or U5627 (N_5627,N_3835,N_3520);
nand U5628 (N_5628,N_3813,N_2806);
and U5629 (N_5629,N_3902,N_4603);
or U5630 (N_5630,N_2905,N_3933);
nand U5631 (N_5631,N_2940,N_3734);
and U5632 (N_5632,N_4191,N_2807);
xnor U5633 (N_5633,N_3554,N_2618);
xor U5634 (N_5634,N_3754,N_3957);
nor U5635 (N_5635,N_3326,N_3619);
or U5636 (N_5636,N_2628,N_3924);
xor U5637 (N_5637,N_4934,N_4004);
nand U5638 (N_5638,N_3884,N_2759);
nor U5639 (N_5639,N_4590,N_4089);
xor U5640 (N_5640,N_3323,N_4467);
xnor U5641 (N_5641,N_4454,N_2616);
xnor U5642 (N_5642,N_2512,N_3439);
nand U5643 (N_5643,N_4513,N_4006);
or U5644 (N_5644,N_2700,N_3749);
xor U5645 (N_5645,N_2739,N_4304);
xnor U5646 (N_5646,N_4157,N_3207);
and U5647 (N_5647,N_3402,N_2937);
or U5648 (N_5648,N_3907,N_3276);
nor U5649 (N_5649,N_3181,N_3130);
or U5650 (N_5650,N_4420,N_3537);
nor U5651 (N_5651,N_3564,N_3826);
or U5652 (N_5652,N_4807,N_3128);
nor U5653 (N_5653,N_4849,N_4215);
nor U5654 (N_5654,N_3922,N_4281);
nand U5655 (N_5655,N_2986,N_3822);
xnor U5656 (N_5656,N_4197,N_3299);
and U5657 (N_5657,N_3652,N_3361);
nor U5658 (N_5658,N_2679,N_4786);
and U5659 (N_5659,N_3839,N_3206);
or U5660 (N_5660,N_4102,N_2575);
nand U5661 (N_5661,N_4026,N_2717);
nand U5662 (N_5662,N_4650,N_3210);
nand U5663 (N_5663,N_4941,N_3700);
nand U5664 (N_5664,N_2753,N_3463);
or U5665 (N_5665,N_2648,N_3201);
and U5666 (N_5666,N_3760,N_3657);
xor U5667 (N_5667,N_3628,N_4411);
nand U5668 (N_5668,N_4094,N_2515);
or U5669 (N_5669,N_4288,N_3683);
and U5670 (N_5670,N_4011,N_3781);
nand U5671 (N_5671,N_2863,N_3406);
nor U5672 (N_5672,N_3397,N_4565);
xnor U5673 (N_5673,N_3882,N_3780);
or U5674 (N_5674,N_3629,N_4214);
xor U5675 (N_5675,N_3691,N_2856);
and U5676 (N_5676,N_4184,N_3234);
or U5677 (N_5677,N_3114,N_3437);
or U5678 (N_5678,N_3676,N_3701);
or U5679 (N_5679,N_4817,N_2684);
and U5680 (N_5680,N_4539,N_4129);
or U5681 (N_5681,N_4152,N_2814);
nand U5682 (N_5682,N_3421,N_4168);
nand U5683 (N_5683,N_4593,N_3257);
nand U5684 (N_5684,N_2527,N_3302);
or U5685 (N_5685,N_4408,N_2591);
and U5686 (N_5686,N_4174,N_4127);
nor U5687 (N_5687,N_3634,N_3972);
nand U5688 (N_5688,N_2909,N_2611);
nor U5689 (N_5689,N_4173,N_4693);
nor U5690 (N_5690,N_3909,N_4744);
and U5691 (N_5691,N_3858,N_4051);
nand U5692 (N_5692,N_3486,N_3091);
and U5693 (N_5693,N_4482,N_3604);
and U5694 (N_5694,N_4297,N_3659);
nand U5695 (N_5695,N_3782,N_4750);
nor U5696 (N_5696,N_4423,N_4757);
nor U5697 (N_5697,N_4965,N_2595);
xor U5698 (N_5698,N_4985,N_4842);
and U5699 (N_5699,N_3407,N_3202);
or U5700 (N_5700,N_2662,N_3804);
nor U5701 (N_5701,N_4323,N_4318);
or U5702 (N_5702,N_2511,N_2509);
nand U5703 (N_5703,N_3465,N_2791);
nand U5704 (N_5704,N_2782,N_2615);
or U5705 (N_5705,N_4715,N_3423);
nand U5706 (N_5706,N_3097,N_4978);
xor U5707 (N_5707,N_3859,N_4440);
or U5708 (N_5708,N_3875,N_4309);
and U5709 (N_5709,N_3563,N_4781);
nor U5710 (N_5710,N_4785,N_3426);
nand U5711 (N_5711,N_4629,N_2945);
and U5712 (N_5712,N_4183,N_4050);
nand U5713 (N_5713,N_3029,N_4531);
nand U5714 (N_5714,N_3733,N_3784);
nor U5715 (N_5715,N_3655,N_3411);
or U5716 (N_5716,N_4424,N_3656);
or U5717 (N_5717,N_2685,N_2874);
nand U5718 (N_5718,N_3968,N_4959);
nor U5719 (N_5719,N_3605,N_4534);
nor U5720 (N_5720,N_2891,N_3352);
or U5721 (N_5721,N_4287,N_3532);
and U5722 (N_5722,N_3932,N_3170);
nor U5723 (N_5723,N_4248,N_2737);
or U5724 (N_5724,N_3298,N_3417);
nand U5725 (N_5725,N_4246,N_4878);
and U5726 (N_5726,N_3408,N_2614);
nor U5727 (N_5727,N_3558,N_4347);
nand U5728 (N_5728,N_3020,N_3765);
nand U5729 (N_5729,N_4811,N_4746);
and U5730 (N_5730,N_4929,N_3731);
xor U5731 (N_5731,N_3176,N_4021);
or U5732 (N_5732,N_2804,N_2815);
nand U5733 (N_5733,N_4331,N_4704);
nand U5734 (N_5734,N_2851,N_4891);
nor U5735 (N_5735,N_3609,N_3216);
nor U5736 (N_5736,N_3405,N_4832);
xnor U5737 (N_5737,N_2879,N_3711);
xnor U5738 (N_5738,N_3412,N_4141);
nor U5739 (N_5739,N_4414,N_3166);
xnor U5740 (N_5740,N_3817,N_3041);
xor U5741 (N_5741,N_2654,N_3757);
and U5742 (N_5742,N_3307,N_3915);
nor U5743 (N_5743,N_4379,N_3485);
nand U5744 (N_5744,N_2645,N_4862);
or U5745 (N_5745,N_3180,N_3579);
or U5746 (N_5746,N_2505,N_3653);
or U5747 (N_5747,N_3977,N_2680);
nand U5748 (N_5748,N_4986,N_2696);
nand U5749 (N_5749,N_3434,N_3777);
nor U5750 (N_5750,N_3602,N_2965);
nor U5751 (N_5751,N_2535,N_2812);
nor U5752 (N_5752,N_3011,N_3116);
xnor U5753 (N_5753,N_4263,N_3967);
or U5754 (N_5754,N_2995,N_3108);
nand U5755 (N_5755,N_3627,N_4972);
and U5756 (N_5756,N_3821,N_4882);
nand U5757 (N_5757,N_4871,N_2539);
or U5758 (N_5758,N_2705,N_4321);
xnor U5759 (N_5759,N_3885,N_4883);
and U5760 (N_5760,N_3662,N_4575);
and U5761 (N_5761,N_4267,N_2735);
nand U5762 (N_5762,N_3123,N_4663);
xnor U5763 (N_5763,N_3028,N_4402);
xor U5764 (N_5764,N_3905,N_2554);
nand U5765 (N_5765,N_4963,N_3277);
xor U5766 (N_5766,N_3043,N_3389);
nor U5767 (N_5767,N_3363,N_4143);
nor U5768 (N_5768,N_2947,N_3447);
nor U5769 (N_5769,N_3001,N_4169);
and U5770 (N_5770,N_4468,N_3430);
nand U5771 (N_5771,N_4591,N_2736);
nand U5772 (N_5772,N_3601,N_3136);
or U5773 (N_5773,N_3737,N_4874);
nand U5774 (N_5774,N_3401,N_4713);
and U5775 (N_5775,N_4751,N_3759);
or U5776 (N_5776,N_4266,N_2666);
xor U5777 (N_5777,N_4361,N_3286);
and U5778 (N_5778,N_3878,N_4545);
nand U5779 (N_5779,N_2719,N_4293);
or U5780 (N_5780,N_3639,N_3945);
nor U5781 (N_5781,N_3718,N_3876);
xnor U5782 (N_5782,N_4791,N_4095);
or U5783 (N_5783,N_4043,N_4851);
nand U5784 (N_5784,N_4873,N_2690);
or U5785 (N_5785,N_4695,N_4572);
nor U5786 (N_5786,N_4086,N_4284);
xnor U5787 (N_5787,N_4760,N_4651);
and U5788 (N_5788,N_4471,N_2752);
and U5789 (N_5789,N_3198,N_3668);
nand U5790 (N_5790,N_4902,N_3798);
nand U5791 (N_5791,N_4776,N_2501);
nor U5792 (N_5792,N_3879,N_2738);
and U5793 (N_5793,N_3988,N_3595);
or U5794 (N_5794,N_3117,N_3519);
or U5795 (N_5795,N_3192,N_4386);
and U5796 (N_5796,N_3288,N_2787);
nand U5797 (N_5797,N_3952,N_3539);
nand U5798 (N_5798,N_4970,N_2852);
and U5799 (N_5799,N_3025,N_2902);
and U5800 (N_5800,N_3873,N_3693);
or U5801 (N_5801,N_3386,N_2528);
and U5802 (N_5802,N_4517,N_3482);
or U5803 (N_5803,N_4190,N_3445);
nand U5804 (N_5804,N_4213,N_2580);
or U5805 (N_5805,N_4188,N_4806);
or U5806 (N_5806,N_4496,N_3881);
xnor U5807 (N_5807,N_3774,N_3359);
or U5808 (N_5808,N_4525,N_4425);
or U5809 (N_5809,N_3587,N_3252);
xor U5810 (N_5810,N_3351,N_3741);
and U5811 (N_5811,N_4556,N_2704);
and U5812 (N_5812,N_2906,N_4589);
nor U5813 (N_5813,N_3239,N_2912);
or U5814 (N_5814,N_3483,N_3556);
xor U5815 (N_5815,N_4541,N_4159);
nand U5816 (N_5816,N_4242,N_4290);
nor U5817 (N_5817,N_3214,N_2873);
nor U5818 (N_5818,N_4623,N_3247);
nand U5819 (N_5819,N_3218,N_4033);
nand U5820 (N_5820,N_4961,N_3146);
xor U5821 (N_5821,N_3908,N_3333);
and U5822 (N_5822,N_3316,N_2574);
nand U5823 (N_5823,N_4639,N_3801);
and U5824 (N_5824,N_3607,N_4087);
xor U5825 (N_5825,N_3016,N_3319);
nand U5826 (N_5826,N_2681,N_2846);
or U5827 (N_5827,N_2987,N_3779);
nand U5828 (N_5828,N_2763,N_2538);
nand U5829 (N_5829,N_3285,N_3755);
and U5830 (N_5830,N_3854,N_3661);
or U5831 (N_5831,N_4370,N_2899);
xnor U5832 (N_5832,N_4818,N_2634);
and U5833 (N_5833,N_3194,N_4055);
nand U5834 (N_5834,N_2811,N_4495);
nor U5835 (N_5835,N_3009,N_3768);
and U5836 (N_5836,N_2930,N_4699);
and U5837 (N_5837,N_2518,N_3469);
nor U5838 (N_5838,N_3413,N_3338);
xnor U5839 (N_5839,N_2721,N_3612);
nor U5840 (N_5840,N_3245,N_2857);
and U5841 (N_5841,N_3921,N_2584);
xnor U5842 (N_5842,N_3738,N_2655);
or U5843 (N_5843,N_3890,N_4759);
and U5844 (N_5844,N_2503,N_4265);
xor U5845 (N_5845,N_4770,N_4881);
and U5846 (N_5846,N_4707,N_3000);
xnor U5847 (N_5847,N_4598,N_3022);
and U5848 (N_5848,N_4310,N_3056);
xor U5849 (N_5849,N_3895,N_4668);
xnor U5850 (N_5850,N_4131,N_4974);
and U5851 (N_5851,N_3137,N_3788);
or U5852 (N_5852,N_3995,N_4717);
nand U5853 (N_5853,N_4060,N_2860);
xor U5854 (N_5854,N_3509,N_4147);
and U5855 (N_5855,N_3111,N_2985);
nor U5856 (N_5856,N_3051,N_4401);
nand U5857 (N_5857,N_3585,N_2881);
and U5858 (N_5858,N_2918,N_2988);
nand U5859 (N_5859,N_4529,N_3736);
nand U5860 (N_5860,N_2880,N_4738);
and U5861 (N_5861,N_4298,N_3036);
nand U5862 (N_5862,N_3101,N_4685);
and U5863 (N_5863,N_4644,N_4991);
nand U5864 (N_5864,N_4843,N_4208);
and U5865 (N_5865,N_4422,N_2734);
and U5866 (N_5866,N_3521,N_3570);
nand U5867 (N_5867,N_4543,N_3442);
nor U5868 (N_5868,N_3424,N_2657);
nor U5869 (N_5869,N_4212,N_3484);
and U5870 (N_5870,N_3240,N_3911);
xor U5871 (N_5871,N_3112,N_4928);
xnor U5872 (N_5872,N_4200,N_2970);
and U5873 (N_5873,N_4956,N_4398);
xnor U5874 (N_5874,N_4846,N_4914);
or U5875 (N_5875,N_3451,N_3221);
and U5876 (N_5876,N_2978,N_4031);
xnor U5877 (N_5877,N_4943,N_2547);
or U5878 (N_5878,N_3152,N_3692);
xor U5879 (N_5879,N_3450,N_3063);
nand U5880 (N_5880,N_3544,N_2981);
xnor U5881 (N_5881,N_4394,N_2770);
nor U5882 (N_5882,N_3303,N_3606);
nand U5883 (N_5883,N_4005,N_2840);
nor U5884 (N_5884,N_3796,N_4665);
xnor U5885 (N_5885,N_3526,N_4827);
and U5886 (N_5886,N_2516,N_3747);
and U5887 (N_5887,N_4994,N_4748);
and U5888 (N_5888,N_4935,N_4720);
xor U5889 (N_5889,N_2948,N_3435);
nand U5890 (N_5890,N_3727,N_2590);
or U5891 (N_5891,N_4924,N_4895);
xor U5892 (N_5892,N_3756,N_3742);
or U5893 (N_5893,N_4570,N_2887);
and U5894 (N_5894,N_4389,N_3258);
or U5895 (N_5895,N_3767,N_2703);
or U5896 (N_5896,N_2581,N_3516);
xnor U5897 (N_5897,N_4566,N_4271);
nor U5898 (N_5898,N_4185,N_4444);
nor U5899 (N_5899,N_3062,N_3183);
xor U5900 (N_5900,N_3568,N_2817);
and U5901 (N_5901,N_3226,N_3989);
or U5902 (N_5902,N_3773,N_4863);
and U5903 (N_5903,N_3227,N_3722);
or U5904 (N_5904,N_4450,N_3883);
nor U5905 (N_5905,N_4950,N_3119);
or U5906 (N_5906,N_3164,N_4463);
or U5907 (N_5907,N_3081,N_2626);
xor U5908 (N_5908,N_2922,N_3085);
xnor U5909 (N_5909,N_4296,N_3547);
nand U5910 (N_5910,N_4481,N_2639);
xnor U5911 (N_5911,N_2896,N_3499);
xnor U5912 (N_5912,N_3511,N_4877);
nand U5913 (N_5913,N_2974,N_3125);
and U5914 (N_5914,N_3173,N_4839);
nand U5915 (N_5915,N_3860,N_4383);
and U5916 (N_5916,N_2929,N_4626);
nor U5917 (N_5917,N_2541,N_2641);
or U5918 (N_5918,N_4476,N_2847);
or U5919 (N_5919,N_3193,N_4588);
xnor U5920 (N_5920,N_2892,N_4079);
and U5921 (N_5921,N_2607,N_4530);
xor U5922 (N_5922,N_3360,N_3807);
xor U5923 (N_5923,N_3034,N_4859);
nor U5924 (N_5924,N_3148,N_4559);
xor U5925 (N_5925,N_3347,N_3917);
and U5926 (N_5926,N_3925,N_4366);
nand U5927 (N_5927,N_4069,N_3505);
nand U5928 (N_5928,N_4798,N_2875);
or U5929 (N_5929,N_4325,N_4488);
xnor U5930 (N_5930,N_4035,N_4837);
xor U5931 (N_5931,N_2901,N_4581);
xor U5932 (N_5932,N_4455,N_3502);
nand U5933 (N_5933,N_4861,N_3399);
or U5934 (N_5934,N_2714,N_4065);
nand U5935 (N_5935,N_2600,N_3600);
nor U5936 (N_5936,N_4070,N_4550);
nand U5937 (N_5937,N_4111,N_4657);
and U5938 (N_5938,N_4984,N_4083);
xnor U5939 (N_5939,N_4216,N_3834);
xnor U5940 (N_5940,N_2764,N_2612);
xnor U5941 (N_5941,N_2908,N_3899);
nand U5942 (N_5942,N_4852,N_4018);
or U5943 (N_5943,N_3233,N_4906);
nor U5944 (N_5944,N_4571,N_3833);
and U5945 (N_5945,N_4483,N_4733);
nand U5946 (N_5946,N_3456,N_3109);
or U5947 (N_5947,N_4722,N_4826);
or U5948 (N_5948,N_3238,N_3495);
xor U5949 (N_5949,N_2894,N_4514);
or U5950 (N_5950,N_2809,N_3491);
or U5951 (N_5951,N_4103,N_4945);
and U5952 (N_5952,N_3342,N_4396);
nor U5953 (N_5953,N_4814,N_4967);
nor U5954 (N_5954,N_4076,N_4431);
nor U5955 (N_5955,N_4597,N_2744);
or U5956 (N_5956,N_4542,N_3872);
nand U5957 (N_5957,N_4151,N_3681);
or U5958 (N_5958,N_4433,N_3739);
nor U5959 (N_5959,N_3624,N_2877);
and U5960 (N_5960,N_3775,N_4754);
and U5961 (N_5961,N_4957,N_4880);
xor U5962 (N_5962,N_4820,N_4198);
nor U5963 (N_5963,N_2553,N_3949);
and U5964 (N_5964,N_4627,N_2959);
xnor U5965 (N_5965,N_4187,N_4345);
nand U5966 (N_5966,N_4997,N_3070);
nor U5967 (N_5967,N_4771,N_4594);
nand U5968 (N_5968,N_4195,N_3131);
xnor U5969 (N_5969,N_2821,N_3971);
nand U5970 (N_5970,N_4204,N_3013);
or U5971 (N_5971,N_3617,N_4858);
and U5972 (N_5972,N_4286,N_4462);
xor U5973 (N_5973,N_4435,N_4801);
xnor U5974 (N_5974,N_4939,N_4301);
nand U5975 (N_5975,N_4672,N_4675);
and U5976 (N_5976,N_2904,N_2993);
or U5977 (N_5977,N_4295,N_4952);
or U5978 (N_5978,N_3552,N_2826);
xor U5979 (N_5979,N_2564,N_4395);
nor U5980 (N_5980,N_4512,N_4558);
nor U5981 (N_5981,N_3745,N_4840);
nor U5982 (N_5982,N_4922,N_3666);
nand U5983 (N_5983,N_4777,N_4171);
nor U5984 (N_5984,N_3824,N_3665);
and U5985 (N_5985,N_3751,N_4466);
and U5986 (N_5986,N_3158,N_2665);
nor U5987 (N_5987,N_4876,N_4879);
and U5988 (N_5988,N_2798,N_4509);
nand U5989 (N_5989,N_4548,N_3856);
xnor U5990 (N_5990,N_4357,N_2673);
nand U5991 (N_5991,N_4731,N_2644);
nor U5992 (N_5992,N_3640,N_2927);
nor U5993 (N_5993,N_3635,N_4809);
or U5994 (N_5994,N_3851,N_3746);
xor U5995 (N_5995,N_2774,N_3008);
or U5996 (N_5996,N_3172,N_4052);
and U5997 (N_5997,N_3297,N_4503);
nand U5998 (N_5998,N_3613,N_4982);
nor U5999 (N_5999,N_2601,N_3958);
or U6000 (N_6000,N_4098,N_3162);
nand U6001 (N_6001,N_2936,N_4679);
nand U6002 (N_6002,N_4372,N_4850);
and U6003 (N_6003,N_3291,N_3443);
nor U6004 (N_6004,N_4020,N_3357);
xor U6005 (N_6005,N_3650,N_3150);
or U6006 (N_6006,N_3458,N_4226);
or U6007 (N_6007,N_4779,N_2870);
xor U6008 (N_6008,N_2546,N_4329);
or U6009 (N_6009,N_4149,N_3848);
or U6010 (N_6010,N_2801,N_3196);
and U6011 (N_6011,N_3031,N_4520);
nor U6012 (N_6012,N_3707,N_4652);
nand U6013 (N_6013,N_3035,N_2642);
nand U6014 (N_6014,N_3144,N_4856);
xor U6015 (N_6015,N_4030,N_4015);
nor U6016 (N_6016,N_3073,N_3576);
and U6017 (N_6017,N_3827,N_3596);
and U6018 (N_6018,N_3237,N_4973);
nand U6019 (N_6019,N_4477,N_4611);
nor U6020 (N_6020,N_3052,N_4322);
and U6021 (N_6021,N_2729,N_3118);
nand U6022 (N_6022,N_2568,N_4038);
nor U6023 (N_6023,N_2939,N_3262);
xnor U6024 (N_6024,N_2676,N_3948);
xnor U6025 (N_6025,N_4262,N_4085);
nor U6026 (N_6026,N_2991,N_2761);
and U6027 (N_6027,N_3182,N_4515);
and U6028 (N_6028,N_4528,N_3837);
and U6029 (N_6029,N_3724,N_4968);
xnor U6030 (N_6030,N_4637,N_4502);
nor U6031 (N_6031,N_4049,N_3867);
and U6032 (N_6032,N_3740,N_2756);
and U6033 (N_6033,N_4428,N_2777);
or U6034 (N_6034,N_3328,N_3588);
nor U6035 (N_6035,N_4270,N_4132);
nor U6036 (N_6036,N_4045,N_4247);
xnor U6037 (N_6037,N_4061,N_3014);
or U6038 (N_6038,N_3195,N_4610);
nand U6039 (N_6039,N_3330,N_3671);
nor U6040 (N_6040,N_4480,N_2820);
nor U6041 (N_6041,N_3771,N_4409);
and U6042 (N_6042,N_3721,N_3446);
nor U6043 (N_6043,N_3082,N_3714);
xnor U6044 (N_6044,N_3886,N_3468);
nor U6045 (N_6045,N_4449,N_3395);
xnor U6046 (N_6046,N_2695,N_2953);
and U6047 (N_6047,N_3614,N_4654);
and U6048 (N_6048,N_2670,N_2637);
nor U6049 (N_6049,N_3710,N_3793);
xor U6050 (N_6050,N_4472,N_4133);
nor U6051 (N_6051,N_4894,N_3339);
or U6052 (N_6052,N_2999,N_3010);
or U6053 (N_6053,N_3567,N_2599);
nand U6054 (N_6054,N_4273,N_3555);
or U6055 (N_6055,N_3943,N_3527);
and U6056 (N_6056,N_4417,N_3160);
and U6057 (N_6057,N_2647,N_3743);
nor U6058 (N_6058,N_2543,N_4245);
nor U6059 (N_6059,N_4251,N_3638);
or U6060 (N_6060,N_2656,N_3694);
xor U6061 (N_6061,N_4202,N_4140);
nor U6062 (N_6062,N_4574,N_2768);
xnor U6063 (N_6063,N_2529,N_4071);
nand U6064 (N_6064,N_3888,N_4148);
nand U6065 (N_6065,N_3868,N_3161);
or U6066 (N_6066,N_3808,N_4359);
or U6067 (N_6067,N_3065,N_4313);
xor U6068 (N_6068,N_2523,N_3618);
xnor U6069 (N_6069,N_4034,N_3615);
and U6070 (N_6070,N_3969,N_4167);
or U6071 (N_6071,N_3802,N_3039);
or U6072 (N_6072,N_2792,N_2872);
and U6073 (N_6073,N_3528,N_4547);
or U6074 (N_6074,N_3084,N_3580);
nor U6075 (N_6075,N_2907,N_4232);
and U6076 (N_6076,N_2844,N_2989);
and U6077 (N_6077,N_4830,N_3901);
or U6078 (N_6078,N_3420,N_4551);
nor U6079 (N_6079,N_2540,N_4014);
or U6080 (N_6080,N_3643,N_3696);
nand U6081 (N_6081,N_2536,N_2745);
nor U6082 (N_6082,N_3522,N_3382);
xnor U6083 (N_6083,N_4649,N_2765);
xor U6084 (N_6084,N_4317,N_2823);
nand U6085 (N_6085,N_4676,N_4170);
and U6086 (N_6086,N_4068,N_2728);
xnor U6087 (N_6087,N_3785,N_4799);
xnor U6088 (N_6088,N_3630,N_4236);
nand U6089 (N_6089,N_4813,N_2520);
and U6090 (N_6090,N_3489,N_4958);
or U6091 (N_6091,N_3748,N_4669);
xor U6092 (N_6092,N_4264,N_4338);
or U6093 (N_6093,N_2571,N_4526);
nor U6094 (N_6094,N_4017,N_4461);
xnor U6095 (N_6095,N_3762,N_3623);
nand U6096 (N_6096,N_3163,N_3296);
nor U6097 (N_6097,N_4308,N_2727);
xor U6098 (N_6098,N_2548,N_4716);
nand U6099 (N_6099,N_4942,N_4441);
xnor U6100 (N_6100,N_2633,N_3462);
nor U6101 (N_6101,N_4698,N_3284);
nor U6102 (N_6102,N_2954,N_4181);
and U6103 (N_6103,N_4616,N_3955);
and U6104 (N_6104,N_4032,N_3590);
nand U6105 (N_6105,N_3047,N_3490);
xor U6106 (N_6106,N_4708,N_4464);
xor U6107 (N_6107,N_4599,N_2562);
and U6108 (N_6108,N_4259,N_4404);
or U6109 (N_6109,N_2664,N_4865);
xor U6110 (N_6110,N_4010,N_2819);
xnor U6111 (N_6111,N_3715,N_2701);
or U6112 (N_6112,N_3177,N_3524);
xor U6113 (N_6113,N_3994,N_3414);
or U6114 (N_6114,N_3121,N_4114);
nor U6115 (N_6115,N_4282,N_2713);
or U6116 (N_6116,N_2733,N_3654);
nor U6117 (N_6117,N_3156,N_3403);
nand U6118 (N_6118,N_4115,N_2845);
xor U6119 (N_6119,N_4341,N_2869);
and U6120 (N_6120,N_4761,N_3769);
and U6121 (N_6121,N_2772,N_3260);
xor U6122 (N_6122,N_2636,N_3191);
or U6123 (N_6123,N_3113,N_4261);
xor U6124 (N_6124,N_4670,N_3792);
nand U6125 (N_6125,N_4374,N_2669);
or U6126 (N_6126,N_4024,N_3246);
nand U6127 (N_6127,N_3632,N_4498);
nor U6128 (N_6128,N_4376,N_3098);
nand U6129 (N_6129,N_3199,N_4691);
nand U6130 (N_6130,N_3023,N_3594);
nor U6131 (N_6131,N_4196,N_4182);
and U6132 (N_6132,N_3334,N_4740);
or U6133 (N_6133,N_2900,N_3845);
or U6134 (N_6134,N_3843,N_4855);
or U6135 (N_6135,N_3235,N_3730);
nor U6136 (N_6136,N_2771,N_4540);
and U6137 (N_6137,N_2635,N_3713);
nand U6138 (N_6138,N_4602,N_4690);
nand U6139 (N_6139,N_4339,N_4305);
xnor U6140 (N_6140,N_3122,N_4522);
nor U6141 (N_6141,N_4124,N_3309);
nand U6142 (N_6142,N_3887,N_4029);
and U6143 (N_6143,N_3300,N_3441);
nor U6144 (N_6144,N_3076,N_2537);
and U6145 (N_6145,N_4125,N_3409);
or U6146 (N_6146,N_4648,N_2977);
nor U6147 (N_6147,N_3830,N_4012);
and U6148 (N_6148,N_3819,N_3586);
and U6149 (N_6149,N_2620,N_2925);
xnor U6150 (N_6150,N_4258,N_4769);
or U6151 (N_6151,N_3571,N_4640);
nor U6152 (N_6152,N_3672,N_4845);
nand U6153 (N_6153,N_4789,N_2510);
nor U6154 (N_6154,N_3341,N_2651);
or U6155 (N_6155,N_3452,N_3517);
nor U6156 (N_6156,N_4028,N_2563);
xnor U6157 (N_6157,N_3726,N_4002);
nand U6158 (N_6158,N_4899,N_3903);
nor U6159 (N_6159,N_3536,N_4342);
or U6160 (N_6160,N_3986,N_3324);
xnor U6161 (N_6161,N_4741,N_2968);
or U6162 (N_6162,N_3680,N_2848);
or U6163 (N_6163,N_4951,N_2796);
or U6164 (N_6164,N_3448,N_4560);
nand U6165 (N_6165,N_3080,N_3275);
or U6166 (N_6166,N_4493,N_4553);
xor U6167 (N_6167,N_4600,N_2915);
nand U6168 (N_6168,N_4576,N_2825);
and U6169 (N_6169,N_4563,N_3761);
nor U6170 (N_6170,N_4938,N_4302);
nand U6171 (N_6171,N_3124,N_2638);
nor U6172 (N_6172,N_4606,N_4521);
or U6173 (N_6173,N_4618,N_4636);
or U6174 (N_6174,N_4656,N_3185);
or U6175 (N_6175,N_3893,N_4358);
or U6176 (N_6176,N_3077,N_4630);
xnor U6177 (N_6177,N_3105,N_3102);
nand U6178 (N_6178,N_2566,N_3603);
nand U6179 (N_6179,N_3950,N_3799);
or U6180 (N_6180,N_3982,N_3332);
and U6181 (N_6181,N_4674,N_3535);
nand U6182 (N_6182,N_2603,N_3072);
xnor U6183 (N_6183,N_4369,N_3599);
nor U6184 (N_6184,N_2784,N_4577);
xor U6185 (N_6185,N_3790,N_2924);
xor U6186 (N_6186,N_3370,N_2613);
and U6187 (N_6187,N_4363,N_3611);
nor U6188 (N_6188,N_2609,N_4382);
nand U6189 (N_6189,N_3510,N_4933);
nand U6190 (N_6190,N_3126,N_4647);
and U6191 (N_6191,N_3115,N_3965);
or U6192 (N_6192,N_4229,N_3705);
and U6193 (N_6193,N_4254,N_4900);
nor U6194 (N_6194,N_4432,N_4854);
or U6195 (N_6195,N_3501,N_4223);
and U6196 (N_6196,N_4516,N_4285);
nor U6197 (N_6197,N_3186,N_3418);
and U6198 (N_6198,N_4682,N_4523);
and U6199 (N_6199,N_4752,N_4365);
xnor U6200 (N_6200,N_4166,N_3978);
xor U6201 (N_6201,N_3795,N_2725);
xnor U6202 (N_6202,N_2610,N_4393);
nor U6203 (N_6203,N_2876,N_4003);
and U6204 (N_6204,N_4497,N_3093);
nor U6205 (N_6205,N_4231,N_4870);
nor U6206 (N_6206,N_4915,N_3974);
nor U6207 (N_6207,N_3806,N_2560);
xor U6208 (N_6208,N_3648,N_4186);
and U6209 (N_6209,N_4714,N_4787);
nand U6210 (N_6210,N_4913,N_3356);
nand U6211 (N_6211,N_2649,N_4278);
and U6212 (N_6212,N_3345,N_4975);
or U6213 (N_6213,N_2754,N_4904);
xnor U6214 (N_6214,N_3143,N_4429);
nor U6215 (N_6215,N_3471,N_3027);
nor U6216 (N_6216,N_3979,N_4336);
nor U6217 (N_6217,N_2602,N_4292);
or U6218 (N_6218,N_4816,N_4013);
nand U6219 (N_6219,N_4044,N_4399);
nand U6220 (N_6220,N_4194,N_4767);
or U6221 (N_6221,N_3142,N_3800);
xor U6222 (N_6222,N_3358,N_3178);
or U6223 (N_6223,N_2683,N_4000);
nor U6224 (N_6224,N_2521,N_4819);
nand U6225 (N_6225,N_3293,N_3154);
xnor U6226 (N_6226,N_4638,N_2952);
xor U6227 (N_6227,N_4007,N_2624);
nor U6228 (N_6228,N_4511,N_4172);
or U6229 (N_6229,N_3870,N_2531);
nor U6230 (N_6230,N_2555,N_3929);
or U6231 (N_6231,N_3584,N_3373);
nand U6232 (N_6232,N_3094,N_4940);
nand U6233 (N_6233,N_3852,N_3506);
nor U6234 (N_6234,N_3139,N_2926);
xnor U6235 (N_6235,N_3153,N_3248);
or U6236 (N_6236,N_3912,N_2850);
nor U6237 (N_6237,N_3498,N_3557);
nand U6238 (N_6238,N_3427,N_4788);
nand U6239 (N_6239,N_4580,N_2576);
xnor U6240 (N_6240,N_3171,N_3213);
or U6241 (N_6241,N_4063,N_4718);
xor U6242 (N_6242,N_3637,N_4946);
xor U6243 (N_6243,N_4737,N_4538);
nor U6244 (N_6244,N_4544,N_2938);
and U6245 (N_6245,N_3104,N_2886);
xnor U6246 (N_6246,N_2946,N_3850);
nor U6247 (N_6247,N_3410,N_4890);
or U6248 (N_6248,N_2710,N_4244);
xor U6249 (N_6249,N_2893,N_3778);
xor U6250 (N_6250,N_2647,N_2904);
and U6251 (N_6251,N_2760,N_4097);
nor U6252 (N_6252,N_4561,N_3133);
nand U6253 (N_6253,N_3011,N_4564);
nor U6254 (N_6254,N_4191,N_3559);
nand U6255 (N_6255,N_4202,N_4895);
nor U6256 (N_6256,N_3174,N_3085);
nor U6257 (N_6257,N_4395,N_3830);
nand U6258 (N_6258,N_3816,N_4065);
and U6259 (N_6259,N_4864,N_3836);
nor U6260 (N_6260,N_4271,N_4763);
xor U6261 (N_6261,N_3204,N_3266);
xor U6262 (N_6262,N_4898,N_4021);
nor U6263 (N_6263,N_4046,N_3241);
nand U6264 (N_6264,N_2740,N_3280);
and U6265 (N_6265,N_4680,N_4652);
or U6266 (N_6266,N_2531,N_3159);
nor U6267 (N_6267,N_3790,N_3981);
xor U6268 (N_6268,N_4854,N_4925);
and U6269 (N_6269,N_4660,N_4890);
and U6270 (N_6270,N_2839,N_4930);
nor U6271 (N_6271,N_3546,N_2860);
and U6272 (N_6272,N_3007,N_2529);
or U6273 (N_6273,N_2960,N_4160);
or U6274 (N_6274,N_3174,N_4882);
nand U6275 (N_6275,N_2518,N_3870);
xnor U6276 (N_6276,N_3372,N_4202);
and U6277 (N_6277,N_4977,N_2990);
xnor U6278 (N_6278,N_3362,N_4684);
or U6279 (N_6279,N_4551,N_4266);
and U6280 (N_6280,N_2544,N_3859);
nand U6281 (N_6281,N_3050,N_3323);
nor U6282 (N_6282,N_3129,N_2640);
or U6283 (N_6283,N_4817,N_4189);
xnor U6284 (N_6284,N_2703,N_3741);
nor U6285 (N_6285,N_3231,N_3655);
nand U6286 (N_6286,N_3420,N_3925);
nand U6287 (N_6287,N_3422,N_4854);
xor U6288 (N_6288,N_4705,N_3289);
nor U6289 (N_6289,N_2931,N_3706);
and U6290 (N_6290,N_4172,N_4731);
nor U6291 (N_6291,N_3716,N_4107);
or U6292 (N_6292,N_3803,N_4929);
nor U6293 (N_6293,N_3588,N_3367);
xnor U6294 (N_6294,N_3337,N_3753);
or U6295 (N_6295,N_3914,N_4475);
and U6296 (N_6296,N_3510,N_3109);
nor U6297 (N_6297,N_4995,N_3017);
and U6298 (N_6298,N_3647,N_4120);
nand U6299 (N_6299,N_4558,N_3409);
or U6300 (N_6300,N_4525,N_3627);
nor U6301 (N_6301,N_3656,N_4119);
or U6302 (N_6302,N_4262,N_3528);
or U6303 (N_6303,N_4121,N_4592);
nand U6304 (N_6304,N_4248,N_3052);
xor U6305 (N_6305,N_4199,N_3289);
or U6306 (N_6306,N_4270,N_3877);
or U6307 (N_6307,N_3246,N_4456);
xnor U6308 (N_6308,N_3379,N_3143);
and U6309 (N_6309,N_4955,N_3499);
nand U6310 (N_6310,N_4677,N_3167);
nand U6311 (N_6311,N_3419,N_3686);
xnor U6312 (N_6312,N_2969,N_3094);
or U6313 (N_6313,N_4620,N_3788);
or U6314 (N_6314,N_4652,N_4018);
or U6315 (N_6315,N_2971,N_3961);
nor U6316 (N_6316,N_4630,N_2798);
nor U6317 (N_6317,N_2940,N_3037);
and U6318 (N_6318,N_4542,N_2955);
nand U6319 (N_6319,N_4972,N_3562);
xor U6320 (N_6320,N_4618,N_3623);
or U6321 (N_6321,N_4659,N_3293);
xnor U6322 (N_6322,N_4733,N_4397);
nor U6323 (N_6323,N_4041,N_3758);
nand U6324 (N_6324,N_4431,N_3273);
nor U6325 (N_6325,N_3016,N_3141);
nor U6326 (N_6326,N_2853,N_2740);
nor U6327 (N_6327,N_4684,N_3398);
xor U6328 (N_6328,N_4121,N_4404);
xor U6329 (N_6329,N_3783,N_3800);
nand U6330 (N_6330,N_4003,N_3097);
and U6331 (N_6331,N_4397,N_2963);
xnor U6332 (N_6332,N_3366,N_2866);
xor U6333 (N_6333,N_3074,N_4302);
nand U6334 (N_6334,N_3130,N_2895);
nor U6335 (N_6335,N_3741,N_3248);
nand U6336 (N_6336,N_4323,N_2616);
nand U6337 (N_6337,N_4200,N_4769);
and U6338 (N_6338,N_3210,N_4428);
nor U6339 (N_6339,N_3117,N_3492);
and U6340 (N_6340,N_4049,N_4839);
nand U6341 (N_6341,N_3716,N_4392);
and U6342 (N_6342,N_4085,N_3415);
xor U6343 (N_6343,N_3658,N_4956);
and U6344 (N_6344,N_4064,N_3714);
nand U6345 (N_6345,N_4178,N_4913);
nand U6346 (N_6346,N_3267,N_4227);
nand U6347 (N_6347,N_3263,N_3671);
and U6348 (N_6348,N_4002,N_3555);
nor U6349 (N_6349,N_4667,N_3750);
or U6350 (N_6350,N_4031,N_4521);
and U6351 (N_6351,N_3574,N_3452);
and U6352 (N_6352,N_3957,N_2667);
xnor U6353 (N_6353,N_2949,N_3553);
xor U6354 (N_6354,N_4590,N_4625);
xnor U6355 (N_6355,N_4042,N_3818);
or U6356 (N_6356,N_4367,N_3231);
nand U6357 (N_6357,N_4588,N_2988);
nor U6358 (N_6358,N_4711,N_3035);
nor U6359 (N_6359,N_4984,N_2721);
xnor U6360 (N_6360,N_3290,N_3275);
xor U6361 (N_6361,N_2927,N_2913);
nand U6362 (N_6362,N_4383,N_3934);
xnor U6363 (N_6363,N_3166,N_4607);
or U6364 (N_6364,N_4858,N_4871);
nand U6365 (N_6365,N_4495,N_4316);
or U6366 (N_6366,N_3664,N_4703);
or U6367 (N_6367,N_4356,N_2799);
or U6368 (N_6368,N_3565,N_3779);
and U6369 (N_6369,N_2570,N_2935);
or U6370 (N_6370,N_4202,N_4022);
nor U6371 (N_6371,N_3226,N_4084);
and U6372 (N_6372,N_3376,N_2968);
and U6373 (N_6373,N_4317,N_3571);
nor U6374 (N_6374,N_4723,N_4669);
nor U6375 (N_6375,N_4522,N_4096);
nand U6376 (N_6376,N_3418,N_4073);
xor U6377 (N_6377,N_4679,N_4077);
nand U6378 (N_6378,N_4450,N_3174);
xnor U6379 (N_6379,N_4458,N_3798);
and U6380 (N_6380,N_2964,N_4149);
xnor U6381 (N_6381,N_3598,N_4942);
nor U6382 (N_6382,N_2738,N_4899);
xor U6383 (N_6383,N_3178,N_4170);
and U6384 (N_6384,N_2840,N_3217);
or U6385 (N_6385,N_3766,N_2511);
nand U6386 (N_6386,N_2583,N_2724);
xor U6387 (N_6387,N_3246,N_3850);
and U6388 (N_6388,N_4645,N_4133);
nand U6389 (N_6389,N_2567,N_3600);
xor U6390 (N_6390,N_4146,N_2698);
xnor U6391 (N_6391,N_3028,N_2886);
nor U6392 (N_6392,N_4455,N_2591);
nand U6393 (N_6393,N_3727,N_3185);
nor U6394 (N_6394,N_3305,N_3521);
nand U6395 (N_6395,N_4927,N_3327);
xor U6396 (N_6396,N_2622,N_3180);
nand U6397 (N_6397,N_4558,N_3074);
xnor U6398 (N_6398,N_4244,N_3661);
nor U6399 (N_6399,N_3197,N_2946);
and U6400 (N_6400,N_3971,N_4827);
or U6401 (N_6401,N_4658,N_2662);
nor U6402 (N_6402,N_3999,N_2619);
nand U6403 (N_6403,N_3283,N_3915);
and U6404 (N_6404,N_3185,N_3757);
nand U6405 (N_6405,N_4940,N_4014);
and U6406 (N_6406,N_4459,N_4118);
or U6407 (N_6407,N_4508,N_3434);
and U6408 (N_6408,N_3046,N_4934);
or U6409 (N_6409,N_2829,N_2697);
xor U6410 (N_6410,N_3568,N_4780);
xor U6411 (N_6411,N_4256,N_2712);
or U6412 (N_6412,N_2561,N_3863);
xnor U6413 (N_6413,N_2541,N_4727);
or U6414 (N_6414,N_3989,N_3937);
nor U6415 (N_6415,N_4780,N_2609);
or U6416 (N_6416,N_4512,N_3327);
nand U6417 (N_6417,N_3657,N_2693);
xor U6418 (N_6418,N_4316,N_3602);
or U6419 (N_6419,N_3133,N_3317);
xor U6420 (N_6420,N_2855,N_4608);
or U6421 (N_6421,N_3875,N_3179);
and U6422 (N_6422,N_2820,N_3010);
xnor U6423 (N_6423,N_2678,N_2561);
and U6424 (N_6424,N_2652,N_4420);
nand U6425 (N_6425,N_4347,N_3555);
and U6426 (N_6426,N_3957,N_3716);
xor U6427 (N_6427,N_3240,N_3625);
xor U6428 (N_6428,N_4534,N_3073);
or U6429 (N_6429,N_3193,N_3963);
nor U6430 (N_6430,N_2732,N_2561);
nand U6431 (N_6431,N_3352,N_3239);
and U6432 (N_6432,N_2668,N_4778);
and U6433 (N_6433,N_4116,N_4004);
nand U6434 (N_6434,N_4152,N_4554);
xnor U6435 (N_6435,N_3025,N_4786);
and U6436 (N_6436,N_4502,N_3446);
and U6437 (N_6437,N_3101,N_3129);
or U6438 (N_6438,N_4675,N_2912);
and U6439 (N_6439,N_3416,N_3995);
and U6440 (N_6440,N_2945,N_3148);
nand U6441 (N_6441,N_3633,N_3680);
xor U6442 (N_6442,N_2579,N_3795);
nor U6443 (N_6443,N_3636,N_2863);
nor U6444 (N_6444,N_4829,N_3129);
and U6445 (N_6445,N_3930,N_3064);
nand U6446 (N_6446,N_2831,N_3312);
nor U6447 (N_6447,N_4380,N_3436);
xor U6448 (N_6448,N_3406,N_2767);
xor U6449 (N_6449,N_4634,N_4415);
or U6450 (N_6450,N_4495,N_2557);
or U6451 (N_6451,N_3769,N_3330);
xor U6452 (N_6452,N_3869,N_4047);
xnor U6453 (N_6453,N_2719,N_4616);
or U6454 (N_6454,N_4146,N_3967);
and U6455 (N_6455,N_3176,N_2974);
xnor U6456 (N_6456,N_3981,N_4751);
or U6457 (N_6457,N_4014,N_2775);
nand U6458 (N_6458,N_3254,N_3364);
xnor U6459 (N_6459,N_2897,N_4687);
and U6460 (N_6460,N_3865,N_3150);
nor U6461 (N_6461,N_3183,N_2528);
nor U6462 (N_6462,N_3702,N_4036);
nor U6463 (N_6463,N_4404,N_4762);
and U6464 (N_6464,N_4584,N_3714);
and U6465 (N_6465,N_4196,N_4437);
nand U6466 (N_6466,N_3856,N_3433);
or U6467 (N_6467,N_3230,N_4223);
nor U6468 (N_6468,N_4129,N_4604);
nor U6469 (N_6469,N_2936,N_3472);
and U6470 (N_6470,N_3356,N_3143);
or U6471 (N_6471,N_4173,N_4902);
or U6472 (N_6472,N_2977,N_3719);
or U6473 (N_6473,N_4724,N_4305);
xnor U6474 (N_6474,N_2926,N_4730);
or U6475 (N_6475,N_2975,N_3289);
nor U6476 (N_6476,N_2791,N_2590);
nand U6477 (N_6477,N_3221,N_4917);
or U6478 (N_6478,N_4739,N_4956);
nand U6479 (N_6479,N_4006,N_2822);
nand U6480 (N_6480,N_4193,N_3116);
and U6481 (N_6481,N_3585,N_3228);
xnor U6482 (N_6482,N_3015,N_3616);
xor U6483 (N_6483,N_4458,N_3214);
or U6484 (N_6484,N_2932,N_3279);
nand U6485 (N_6485,N_3216,N_2923);
xor U6486 (N_6486,N_2532,N_3916);
xor U6487 (N_6487,N_2562,N_3943);
nand U6488 (N_6488,N_3287,N_4686);
xnor U6489 (N_6489,N_4356,N_3055);
or U6490 (N_6490,N_3556,N_4841);
and U6491 (N_6491,N_4187,N_3546);
and U6492 (N_6492,N_3703,N_4505);
xnor U6493 (N_6493,N_3461,N_2629);
nand U6494 (N_6494,N_2505,N_4193);
and U6495 (N_6495,N_4449,N_3157);
nor U6496 (N_6496,N_2557,N_2895);
or U6497 (N_6497,N_4229,N_2646);
xnor U6498 (N_6498,N_3020,N_2776);
nand U6499 (N_6499,N_3950,N_3620);
and U6500 (N_6500,N_2917,N_2860);
or U6501 (N_6501,N_3416,N_3510);
and U6502 (N_6502,N_3357,N_3454);
nand U6503 (N_6503,N_3829,N_4903);
nor U6504 (N_6504,N_2836,N_2888);
nor U6505 (N_6505,N_2705,N_4275);
and U6506 (N_6506,N_4583,N_4758);
or U6507 (N_6507,N_4890,N_4260);
nand U6508 (N_6508,N_2882,N_3277);
or U6509 (N_6509,N_4201,N_2936);
xor U6510 (N_6510,N_2989,N_4560);
nor U6511 (N_6511,N_4853,N_3662);
xnor U6512 (N_6512,N_3794,N_3338);
nor U6513 (N_6513,N_3418,N_3696);
nand U6514 (N_6514,N_4434,N_2924);
and U6515 (N_6515,N_3989,N_2644);
nand U6516 (N_6516,N_4755,N_4121);
or U6517 (N_6517,N_3825,N_3820);
nand U6518 (N_6518,N_4783,N_3714);
nor U6519 (N_6519,N_3791,N_3169);
nand U6520 (N_6520,N_4012,N_4775);
and U6521 (N_6521,N_3270,N_3608);
nor U6522 (N_6522,N_4925,N_4799);
or U6523 (N_6523,N_4584,N_3626);
nor U6524 (N_6524,N_4511,N_2641);
or U6525 (N_6525,N_4852,N_3956);
nand U6526 (N_6526,N_2882,N_3334);
or U6527 (N_6527,N_3600,N_3808);
and U6528 (N_6528,N_3607,N_2853);
xnor U6529 (N_6529,N_4933,N_2611);
or U6530 (N_6530,N_4635,N_2861);
nand U6531 (N_6531,N_3226,N_4202);
or U6532 (N_6532,N_4100,N_4206);
nand U6533 (N_6533,N_4464,N_4968);
and U6534 (N_6534,N_2538,N_4709);
and U6535 (N_6535,N_4345,N_4887);
and U6536 (N_6536,N_3615,N_3855);
and U6537 (N_6537,N_2950,N_3361);
nor U6538 (N_6538,N_3420,N_4077);
or U6539 (N_6539,N_3131,N_2921);
or U6540 (N_6540,N_3583,N_3154);
nor U6541 (N_6541,N_4461,N_2575);
or U6542 (N_6542,N_3114,N_3895);
nor U6543 (N_6543,N_3360,N_3815);
xnor U6544 (N_6544,N_3716,N_4262);
nor U6545 (N_6545,N_4407,N_3441);
nand U6546 (N_6546,N_4594,N_2911);
nand U6547 (N_6547,N_4067,N_3187);
or U6548 (N_6548,N_3722,N_4193);
nand U6549 (N_6549,N_3728,N_3961);
nor U6550 (N_6550,N_4519,N_4504);
and U6551 (N_6551,N_3749,N_3552);
xor U6552 (N_6552,N_4708,N_3247);
and U6553 (N_6553,N_3858,N_3474);
and U6554 (N_6554,N_4241,N_2582);
xor U6555 (N_6555,N_2839,N_2944);
nor U6556 (N_6556,N_2532,N_3469);
xnor U6557 (N_6557,N_3273,N_3270);
nand U6558 (N_6558,N_4389,N_4619);
nor U6559 (N_6559,N_3440,N_3896);
and U6560 (N_6560,N_4811,N_4932);
nand U6561 (N_6561,N_3297,N_2930);
and U6562 (N_6562,N_3973,N_4970);
or U6563 (N_6563,N_3020,N_4866);
xnor U6564 (N_6564,N_4202,N_4518);
or U6565 (N_6565,N_4559,N_3229);
nand U6566 (N_6566,N_4018,N_3528);
xnor U6567 (N_6567,N_3825,N_2693);
nand U6568 (N_6568,N_3502,N_3424);
and U6569 (N_6569,N_3985,N_2809);
xor U6570 (N_6570,N_3776,N_4442);
nand U6571 (N_6571,N_4476,N_4091);
and U6572 (N_6572,N_4231,N_4874);
nor U6573 (N_6573,N_3243,N_3319);
xor U6574 (N_6574,N_3599,N_4903);
nor U6575 (N_6575,N_2944,N_4844);
nand U6576 (N_6576,N_3011,N_3814);
nand U6577 (N_6577,N_2593,N_3753);
and U6578 (N_6578,N_3040,N_3572);
nor U6579 (N_6579,N_4923,N_3483);
nand U6580 (N_6580,N_3574,N_4278);
xor U6581 (N_6581,N_2808,N_2997);
nor U6582 (N_6582,N_2905,N_4812);
xor U6583 (N_6583,N_3573,N_2609);
nand U6584 (N_6584,N_3324,N_3571);
or U6585 (N_6585,N_3468,N_3184);
xnor U6586 (N_6586,N_3937,N_2737);
or U6587 (N_6587,N_2617,N_2993);
and U6588 (N_6588,N_3219,N_4214);
nor U6589 (N_6589,N_4536,N_3411);
nand U6590 (N_6590,N_3422,N_3377);
and U6591 (N_6591,N_3473,N_4165);
nand U6592 (N_6592,N_3895,N_3364);
or U6593 (N_6593,N_3088,N_4138);
nand U6594 (N_6594,N_3225,N_3302);
nor U6595 (N_6595,N_3308,N_4994);
and U6596 (N_6596,N_3700,N_3141);
and U6597 (N_6597,N_4888,N_3110);
nor U6598 (N_6598,N_4560,N_3962);
or U6599 (N_6599,N_4640,N_4431);
and U6600 (N_6600,N_4652,N_3709);
xnor U6601 (N_6601,N_3451,N_3405);
or U6602 (N_6602,N_2942,N_3989);
nor U6603 (N_6603,N_3836,N_3970);
xnor U6604 (N_6604,N_3672,N_4771);
and U6605 (N_6605,N_3046,N_3224);
and U6606 (N_6606,N_3400,N_3596);
xor U6607 (N_6607,N_3688,N_4543);
xor U6608 (N_6608,N_2541,N_4792);
and U6609 (N_6609,N_3633,N_4591);
nor U6610 (N_6610,N_3871,N_3146);
or U6611 (N_6611,N_2943,N_3892);
or U6612 (N_6612,N_3961,N_2855);
nor U6613 (N_6613,N_3376,N_2615);
nor U6614 (N_6614,N_4820,N_4858);
nand U6615 (N_6615,N_4199,N_4728);
xnor U6616 (N_6616,N_4570,N_3092);
xnor U6617 (N_6617,N_3963,N_4561);
xor U6618 (N_6618,N_4470,N_3656);
or U6619 (N_6619,N_4415,N_2636);
xnor U6620 (N_6620,N_3641,N_4445);
xnor U6621 (N_6621,N_3430,N_4215);
xor U6622 (N_6622,N_4270,N_3902);
nor U6623 (N_6623,N_4775,N_3111);
or U6624 (N_6624,N_4644,N_2888);
and U6625 (N_6625,N_4061,N_3920);
nand U6626 (N_6626,N_4741,N_3976);
nand U6627 (N_6627,N_4575,N_4468);
and U6628 (N_6628,N_3248,N_3958);
and U6629 (N_6629,N_3069,N_3822);
nor U6630 (N_6630,N_4154,N_3366);
nand U6631 (N_6631,N_3597,N_3247);
nand U6632 (N_6632,N_2769,N_4720);
and U6633 (N_6633,N_3522,N_4255);
nor U6634 (N_6634,N_4534,N_3910);
xnor U6635 (N_6635,N_4191,N_4619);
nor U6636 (N_6636,N_4116,N_4863);
xnor U6637 (N_6637,N_4534,N_3484);
nor U6638 (N_6638,N_3870,N_4541);
or U6639 (N_6639,N_4327,N_3143);
xnor U6640 (N_6640,N_4469,N_4407);
and U6641 (N_6641,N_4794,N_3422);
and U6642 (N_6642,N_4078,N_3800);
nand U6643 (N_6643,N_3467,N_3876);
or U6644 (N_6644,N_2955,N_2601);
nand U6645 (N_6645,N_4402,N_3740);
nand U6646 (N_6646,N_3522,N_3294);
nor U6647 (N_6647,N_3137,N_3271);
xor U6648 (N_6648,N_2961,N_4783);
and U6649 (N_6649,N_3008,N_3817);
or U6650 (N_6650,N_4502,N_3774);
nand U6651 (N_6651,N_3389,N_3748);
xnor U6652 (N_6652,N_2760,N_4999);
and U6653 (N_6653,N_3843,N_4412);
or U6654 (N_6654,N_3073,N_3247);
and U6655 (N_6655,N_4461,N_2566);
nand U6656 (N_6656,N_3703,N_4198);
and U6657 (N_6657,N_4633,N_3688);
or U6658 (N_6658,N_3122,N_3102);
nand U6659 (N_6659,N_3785,N_3791);
and U6660 (N_6660,N_4836,N_4384);
and U6661 (N_6661,N_3511,N_4925);
nand U6662 (N_6662,N_4331,N_3855);
or U6663 (N_6663,N_3952,N_2536);
or U6664 (N_6664,N_4786,N_3981);
or U6665 (N_6665,N_3661,N_3348);
or U6666 (N_6666,N_4415,N_4109);
or U6667 (N_6667,N_4880,N_2937);
or U6668 (N_6668,N_4459,N_3384);
nor U6669 (N_6669,N_4494,N_3565);
nor U6670 (N_6670,N_3761,N_3049);
nand U6671 (N_6671,N_3172,N_3025);
and U6672 (N_6672,N_4023,N_4695);
and U6673 (N_6673,N_2634,N_2746);
and U6674 (N_6674,N_3819,N_4779);
nand U6675 (N_6675,N_3881,N_4503);
nor U6676 (N_6676,N_4666,N_4617);
and U6677 (N_6677,N_2699,N_2588);
or U6678 (N_6678,N_2765,N_4489);
or U6679 (N_6679,N_3864,N_3945);
xor U6680 (N_6680,N_3606,N_4472);
and U6681 (N_6681,N_4594,N_3179);
xor U6682 (N_6682,N_3061,N_3173);
nor U6683 (N_6683,N_2777,N_4667);
nand U6684 (N_6684,N_3753,N_4554);
or U6685 (N_6685,N_3394,N_4317);
xor U6686 (N_6686,N_4363,N_3920);
or U6687 (N_6687,N_4420,N_3856);
or U6688 (N_6688,N_3866,N_2688);
and U6689 (N_6689,N_2590,N_3466);
and U6690 (N_6690,N_3412,N_3504);
or U6691 (N_6691,N_3361,N_4803);
nand U6692 (N_6692,N_4942,N_3926);
nand U6693 (N_6693,N_3946,N_2729);
and U6694 (N_6694,N_2610,N_3186);
xnor U6695 (N_6695,N_2804,N_2642);
nor U6696 (N_6696,N_3584,N_2512);
and U6697 (N_6697,N_4590,N_4375);
nand U6698 (N_6698,N_3479,N_4789);
xnor U6699 (N_6699,N_4127,N_3020);
xor U6700 (N_6700,N_3176,N_4202);
nand U6701 (N_6701,N_3932,N_3251);
xnor U6702 (N_6702,N_4024,N_4953);
nand U6703 (N_6703,N_4346,N_4687);
and U6704 (N_6704,N_4964,N_4403);
xnor U6705 (N_6705,N_4427,N_2956);
nor U6706 (N_6706,N_4374,N_4237);
nand U6707 (N_6707,N_4855,N_2531);
or U6708 (N_6708,N_4857,N_4315);
nor U6709 (N_6709,N_4830,N_3690);
nand U6710 (N_6710,N_4607,N_3958);
nand U6711 (N_6711,N_2820,N_3748);
or U6712 (N_6712,N_4545,N_4155);
or U6713 (N_6713,N_3885,N_4784);
nor U6714 (N_6714,N_4441,N_3817);
and U6715 (N_6715,N_3143,N_2562);
xor U6716 (N_6716,N_3691,N_4520);
or U6717 (N_6717,N_3577,N_4387);
nand U6718 (N_6718,N_4464,N_4995);
and U6719 (N_6719,N_4669,N_4811);
or U6720 (N_6720,N_3120,N_3856);
or U6721 (N_6721,N_4048,N_4568);
nand U6722 (N_6722,N_3105,N_4533);
and U6723 (N_6723,N_3135,N_2654);
or U6724 (N_6724,N_4424,N_2981);
xor U6725 (N_6725,N_2516,N_4634);
and U6726 (N_6726,N_3076,N_4221);
and U6727 (N_6727,N_4883,N_4503);
or U6728 (N_6728,N_4515,N_2889);
nor U6729 (N_6729,N_2921,N_3380);
xor U6730 (N_6730,N_4816,N_3106);
nand U6731 (N_6731,N_2568,N_2774);
nand U6732 (N_6732,N_4216,N_4395);
and U6733 (N_6733,N_3607,N_4748);
and U6734 (N_6734,N_3114,N_3892);
or U6735 (N_6735,N_4374,N_3360);
nand U6736 (N_6736,N_2733,N_3598);
nand U6737 (N_6737,N_3854,N_3417);
nor U6738 (N_6738,N_4149,N_3412);
nor U6739 (N_6739,N_4449,N_2975);
nor U6740 (N_6740,N_2971,N_3475);
or U6741 (N_6741,N_4277,N_2617);
nor U6742 (N_6742,N_3493,N_4738);
nor U6743 (N_6743,N_4551,N_3843);
nor U6744 (N_6744,N_2670,N_3784);
nor U6745 (N_6745,N_2866,N_3027);
xor U6746 (N_6746,N_3865,N_4286);
xor U6747 (N_6747,N_4346,N_3658);
nor U6748 (N_6748,N_4369,N_4372);
nand U6749 (N_6749,N_3883,N_4904);
nand U6750 (N_6750,N_4019,N_3003);
nand U6751 (N_6751,N_3150,N_3790);
or U6752 (N_6752,N_2620,N_4690);
nor U6753 (N_6753,N_2965,N_4330);
or U6754 (N_6754,N_3144,N_3077);
nor U6755 (N_6755,N_4371,N_4723);
nor U6756 (N_6756,N_3441,N_3763);
or U6757 (N_6757,N_4320,N_4232);
xor U6758 (N_6758,N_2795,N_4722);
nor U6759 (N_6759,N_3411,N_4481);
and U6760 (N_6760,N_4756,N_3988);
xnor U6761 (N_6761,N_2701,N_3857);
nor U6762 (N_6762,N_3480,N_4823);
xor U6763 (N_6763,N_4076,N_4366);
or U6764 (N_6764,N_2765,N_4341);
nor U6765 (N_6765,N_3094,N_4474);
or U6766 (N_6766,N_4173,N_2664);
or U6767 (N_6767,N_4480,N_4666);
nor U6768 (N_6768,N_2714,N_2950);
and U6769 (N_6769,N_2573,N_3721);
nand U6770 (N_6770,N_3814,N_3530);
nor U6771 (N_6771,N_2690,N_3669);
xnor U6772 (N_6772,N_4535,N_3100);
xnor U6773 (N_6773,N_4162,N_4011);
nor U6774 (N_6774,N_2988,N_3675);
and U6775 (N_6775,N_2764,N_3805);
or U6776 (N_6776,N_3802,N_2961);
or U6777 (N_6777,N_3649,N_3188);
and U6778 (N_6778,N_4008,N_3972);
and U6779 (N_6779,N_4436,N_4806);
nand U6780 (N_6780,N_2691,N_2898);
or U6781 (N_6781,N_4085,N_2662);
nand U6782 (N_6782,N_4994,N_4815);
xor U6783 (N_6783,N_2968,N_3840);
and U6784 (N_6784,N_4605,N_4821);
nand U6785 (N_6785,N_3935,N_3146);
and U6786 (N_6786,N_3303,N_2863);
and U6787 (N_6787,N_4989,N_4691);
nor U6788 (N_6788,N_2569,N_3395);
or U6789 (N_6789,N_3043,N_2637);
xnor U6790 (N_6790,N_4786,N_4677);
nor U6791 (N_6791,N_3259,N_2859);
nor U6792 (N_6792,N_4800,N_4113);
or U6793 (N_6793,N_4778,N_3900);
xnor U6794 (N_6794,N_3843,N_3874);
nand U6795 (N_6795,N_3228,N_4863);
xor U6796 (N_6796,N_3406,N_3374);
and U6797 (N_6797,N_4899,N_4451);
xor U6798 (N_6798,N_2750,N_3420);
or U6799 (N_6799,N_3935,N_3753);
nor U6800 (N_6800,N_3675,N_2733);
nand U6801 (N_6801,N_3722,N_4829);
nor U6802 (N_6802,N_3567,N_4064);
nor U6803 (N_6803,N_4942,N_4791);
nand U6804 (N_6804,N_2719,N_3498);
and U6805 (N_6805,N_3410,N_3068);
or U6806 (N_6806,N_3370,N_4363);
or U6807 (N_6807,N_4547,N_3095);
nor U6808 (N_6808,N_3507,N_4506);
nor U6809 (N_6809,N_3512,N_2524);
and U6810 (N_6810,N_3493,N_4985);
and U6811 (N_6811,N_4593,N_3690);
and U6812 (N_6812,N_2730,N_3909);
or U6813 (N_6813,N_2688,N_4028);
nor U6814 (N_6814,N_3286,N_2556);
or U6815 (N_6815,N_3844,N_3390);
or U6816 (N_6816,N_4408,N_3357);
nand U6817 (N_6817,N_3576,N_2507);
nand U6818 (N_6818,N_2606,N_4990);
and U6819 (N_6819,N_4644,N_3276);
or U6820 (N_6820,N_2613,N_2946);
xnor U6821 (N_6821,N_4826,N_3340);
or U6822 (N_6822,N_3117,N_2920);
or U6823 (N_6823,N_4236,N_4972);
and U6824 (N_6824,N_4112,N_2975);
nand U6825 (N_6825,N_2930,N_4050);
and U6826 (N_6826,N_2849,N_4047);
xor U6827 (N_6827,N_4449,N_2655);
or U6828 (N_6828,N_4262,N_3312);
nor U6829 (N_6829,N_3596,N_3998);
or U6830 (N_6830,N_3477,N_4639);
nor U6831 (N_6831,N_4837,N_3696);
nand U6832 (N_6832,N_3752,N_3522);
or U6833 (N_6833,N_4899,N_3552);
nand U6834 (N_6834,N_4230,N_4635);
or U6835 (N_6835,N_3375,N_4299);
nand U6836 (N_6836,N_4544,N_3030);
and U6837 (N_6837,N_3576,N_3274);
or U6838 (N_6838,N_3473,N_2923);
and U6839 (N_6839,N_2880,N_4391);
or U6840 (N_6840,N_4620,N_3605);
xnor U6841 (N_6841,N_4031,N_4206);
nand U6842 (N_6842,N_2978,N_3907);
or U6843 (N_6843,N_4264,N_2932);
or U6844 (N_6844,N_2740,N_3870);
nor U6845 (N_6845,N_2776,N_4684);
nor U6846 (N_6846,N_4237,N_4595);
and U6847 (N_6847,N_3371,N_3038);
and U6848 (N_6848,N_4834,N_3118);
xor U6849 (N_6849,N_2616,N_3434);
and U6850 (N_6850,N_3343,N_4025);
xor U6851 (N_6851,N_4528,N_3940);
and U6852 (N_6852,N_3835,N_4007);
nor U6853 (N_6853,N_3087,N_3962);
nand U6854 (N_6854,N_2787,N_2947);
or U6855 (N_6855,N_4402,N_3139);
nor U6856 (N_6856,N_2737,N_4262);
nand U6857 (N_6857,N_3048,N_2629);
and U6858 (N_6858,N_2656,N_4336);
or U6859 (N_6859,N_4257,N_3977);
nor U6860 (N_6860,N_3766,N_2651);
nor U6861 (N_6861,N_2833,N_2948);
nor U6862 (N_6862,N_3493,N_4499);
or U6863 (N_6863,N_3555,N_4418);
and U6864 (N_6864,N_4689,N_3115);
nor U6865 (N_6865,N_4822,N_4635);
or U6866 (N_6866,N_3553,N_4184);
nor U6867 (N_6867,N_4461,N_3084);
nand U6868 (N_6868,N_3963,N_2992);
xor U6869 (N_6869,N_2551,N_3389);
xor U6870 (N_6870,N_3433,N_3034);
or U6871 (N_6871,N_4204,N_2568);
nand U6872 (N_6872,N_4020,N_3703);
xor U6873 (N_6873,N_4463,N_3063);
nor U6874 (N_6874,N_3724,N_4609);
nor U6875 (N_6875,N_4340,N_4903);
nand U6876 (N_6876,N_3981,N_4760);
xor U6877 (N_6877,N_4704,N_3612);
nor U6878 (N_6878,N_3631,N_3145);
xor U6879 (N_6879,N_4997,N_4193);
nand U6880 (N_6880,N_4828,N_4124);
or U6881 (N_6881,N_4778,N_3194);
xor U6882 (N_6882,N_4221,N_3421);
xnor U6883 (N_6883,N_3286,N_4966);
and U6884 (N_6884,N_4904,N_3774);
nand U6885 (N_6885,N_3361,N_2917);
or U6886 (N_6886,N_2803,N_2619);
and U6887 (N_6887,N_3227,N_3136);
xor U6888 (N_6888,N_2553,N_4880);
and U6889 (N_6889,N_4951,N_3531);
nor U6890 (N_6890,N_3701,N_3028);
and U6891 (N_6891,N_3594,N_3953);
xnor U6892 (N_6892,N_3022,N_3799);
or U6893 (N_6893,N_2967,N_3213);
nor U6894 (N_6894,N_4480,N_2839);
nor U6895 (N_6895,N_4816,N_4518);
and U6896 (N_6896,N_3885,N_4703);
xor U6897 (N_6897,N_3691,N_2576);
nor U6898 (N_6898,N_4633,N_3825);
nor U6899 (N_6899,N_4893,N_3226);
nand U6900 (N_6900,N_3885,N_2647);
nand U6901 (N_6901,N_3405,N_4715);
nand U6902 (N_6902,N_4590,N_3620);
nor U6903 (N_6903,N_3660,N_2929);
or U6904 (N_6904,N_2889,N_3486);
or U6905 (N_6905,N_4160,N_3369);
nand U6906 (N_6906,N_4199,N_2572);
xnor U6907 (N_6907,N_4548,N_4425);
xor U6908 (N_6908,N_3018,N_3795);
and U6909 (N_6909,N_3317,N_2505);
nand U6910 (N_6910,N_3409,N_4890);
nand U6911 (N_6911,N_3392,N_3811);
and U6912 (N_6912,N_4235,N_4188);
or U6913 (N_6913,N_4258,N_4430);
nor U6914 (N_6914,N_4290,N_4756);
or U6915 (N_6915,N_3641,N_2518);
nand U6916 (N_6916,N_3648,N_4984);
and U6917 (N_6917,N_3649,N_3216);
nand U6918 (N_6918,N_3952,N_3646);
nand U6919 (N_6919,N_3190,N_4395);
nand U6920 (N_6920,N_4961,N_3209);
nand U6921 (N_6921,N_2554,N_3967);
and U6922 (N_6922,N_4754,N_3934);
xnor U6923 (N_6923,N_4308,N_3651);
and U6924 (N_6924,N_4975,N_3139);
and U6925 (N_6925,N_3762,N_4297);
or U6926 (N_6926,N_2558,N_3004);
xor U6927 (N_6927,N_3003,N_3160);
nor U6928 (N_6928,N_3780,N_2895);
nand U6929 (N_6929,N_2809,N_2541);
and U6930 (N_6930,N_4652,N_2714);
xor U6931 (N_6931,N_2935,N_2927);
and U6932 (N_6932,N_4490,N_3072);
or U6933 (N_6933,N_2511,N_2783);
or U6934 (N_6934,N_3986,N_3443);
or U6935 (N_6935,N_3732,N_2860);
xnor U6936 (N_6936,N_4126,N_2763);
xnor U6937 (N_6937,N_2826,N_3415);
nor U6938 (N_6938,N_3823,N_4652);
xor U6939 (N_6939,N_2984,N_2500);
xnor U6940 (N_6940,N_3437,N_4368);
and U6941 (N_6941,N_3438,N_4558);
xnor U6942 (N_6942,N_4500,N_3695);
and U6943 (N_6943,N_2682,N_3994);
xor U6944 (N_6944,N_3163,N_3390);
and U6945 (N_6945,N_3698,N_4557);
and U6946 (N_6946,N_3008,N_4764);
nor U6947 (N_6947,N_2713,N_4048);
or U6948 (N_6948,N_4601,N_4657);
nand U6949 (N_6949,N_4377,N_4525);
nand U6950 (N_6950,N_2614,N_2585);
nand U6951 (N_6951,N_4144,N_3322);
and U6952 (N_6952,N_3304,N_4757);
nor U6953 (N_6953,N_4591,N_3102);
and U6954 (N_6954,N_4188,N_4549);
nor U6955 (N_6955,N_3751,N_4801);
or U6956 (N_6956,N_3421,N_2759);
and U6957 (N_6957,N_4763,N_3548);
and U6958 (N_6958,N_3515,N_3010);
or U6959 (N_6959,N_4633,N_2740);
and U6960 (N_6960,N_4921,N_4180);
xnor U6961 (N_6961,N_4958,N_3512);
and U6962 (N_6962,N_2811,N_4551);
nor U6963 (N_6963,N_3964,N_3115);
and U6964 (N_6964,N_2894,N_3060);
nor U6965 (N_6965,N_3360,N_3752);
nor U6966 (N_6966,N_4500,N_4572);
nand U6967 (N_6967,N_2968,N_2790);
xnor U6968 (N_6968,N_2626,N_4337);
xor U6969 (N_6969,N_4353,N_4452);
xnor U6970 (N_6970,N_3225,N_3508);
nor U6971 (N_6971,N_4184,N_4853);
xor U6972 (N_6972,N_2578,N_3993);
and U6973 (N_6973,N_3789,N_4698);
nor U6974 (N_6974,N_3985,N_3922);
xor U6975 (N_6975,N_3620,N_4917);
nand U6976 (N_6976,N_3880,N_2854);
xor U6977 (N_6977,N_3796,N_3021);
and U6978 (N_6978,N_4833,N_4925);
or U6979 (N_6979,N_4788,N_3720);
and U6980 (N_6980,N_4643,N_3892);
nor U6981 (N_6981,N_3320,N_4827);
nor U6982 (N_6982,N_4252,N_4250);
nand U6983 (N_6983,N_4611,N_3404);
and U6984 (N_6984,N_4365,N_4782);
and U6985 (N_6985,N_4400,N_4730);
and U6986 (N_6986,N_2882,N_4388);
or U6987 (N_6987,N_4089,N_3066);
and U6988 (N_6988,N_2515,N_4548);
or U6989 (N_6989,N_3780,N_3980);
or U6990 (N_6990,N_3632,N_4362);
nor U6991 (N_6991,N_3377,N_3281);
and U6992 (N_6992,N_2726,N_3692);
nor U6993 (N_6993,N_2523,N_3797);
or U6994 (N_6994,N_3290,N_3315);
or U6995 (N_6995,N_3918,N_2847);
and U6996 (N_6996,N_3790,N_4909);
nor U6997 (N_6997,N_3550,N_2851);
and U6998 (N_6998,N_3226,N_3836);
nand U6999 (N_6999,N_3617,N_2934);
nand U7000 (N_7000,N_2917,N_2794);
xnor U7001 (N_7001,N_3826,N_3050);
xnor U7002 (N_7002,N_2940,N_3993);
nand U7003 (N_7003,N_3572,N_4681);
nor U7004 (N_7004,N_2588,N_4089);
nand U7005 (N_7005,N_2657,N_4486);
nand U7006 (N_7006,N_2903,N_3246);
or U7007 (N_7007,N_3433,N_4710);
or U7008 (N_7008,N_4529,N_2780);
and U7009 (N_7009,N_4097,N_2692);
nand U7010 (N_7010,N_2708,N_3279);
or U7011 (N_7011,N_3358,N_4837);
xnor U7012 (N_7012,N_4890,N_3916);
or U7013 (N_7013,N_4139,N_3204);
xnor U7014 (N_7014,N_3072,N_2889);
nand U7015 (N_7015,N_2540,N_4699);
nand U7016 (N_7016,N_3120,N_3312);
or U7017 (N_7017,N_3024,N_2986);
and U7018 (N_7018,N_3361,N_2562);
nor U7019 (N_7019,N_3221,N_4919);
nand U7020 (N_7020,N_4262,N_4225);
nand U7021 (N_7021,N_3433,N_3348);
and U7022 (N_7022,N_2618,N_4592);
nand U7023 (N_7023,N_4157,N_4951);
xnor U7024 (N_7024,N_4460,N_4836);
or U7025 (N_7025,N_4772,N_3471);
nand U7026 (N_7026,N_4236,N_4046);
xnor U7027 (N_7027,N_4755,N_4715);
nor U7028 (N_7028,N_3138,N_3957);
and U7029 (N_7029,N_4102,N_4220);
nand U7030 (N_7030,N_4525,N_3651);
or U7031 (N_7031,N_3585,N_3574);
and U7032 (N_7032,N_3091,N_4482);
nor U7033 (N_7033,N_4687,N_2806);
nor U7034 (N_7034,N_4838,N_2558);
xor U7035 (N_7035,N_4877,N_4467);
xor U7036 (N_7036,N_4849,N_4710);
nand U7037 (N_7037,N_4708,N_2999);
or U7038 (N_7038,N_2701,N_4315);
xnor U7039 (N_7039,N_3606,N_3239);
xor U7040 (N_7040,N_3893,N_4407);
nand U7041 (N_7041,N_3665,N_3515);
xor U7042 (N_7042,N_4163,N_4939);
xor U7043 (N_7043,N_2979,N_4366);
nor U7044 (N_7044,N_3190,N_3162);
nor U7045 (N_7045,N_3135,N_4655);
xnor U7046 (N_7046,N_4949,N_4919);
and U7047 (N_7047,N_4076,N_3243);
and U7048 (N_7048,N_4781,N_3325);
nand U7049 (N_7049,N_4790,N_4344);
or U7050 (N_7050,N_4195,N_3962);
xnor U7051 (N_7051,N_2593,N_4982);
or U7052 (N_7052,N_4479,N_3504);
nand U7053 (N_7053,N_4536,N_4070);
or U7054 (N_7054,N_4738,N_3102);
nor U7055 (N_7055,N_3554,N_4076);
xor U7056 (N_7056,N_4110,N_2791);
xnor U7057 (N_7057,N_3422,N_4019);
xor U7058 (N_7058,N_4394,N_4646);
or U7059 (N_7059,N_3405,N_4888);
or U7060 (N_7060,N_4539,N_3101);
nor U7061 (N_7061,N_4849,N_3011);
nand U7062 (N_7062,N_4147,N_4460);
xnor U7063 (N_7063,N_4412,N_4868);
nand U7064 (N_7064,N_4467,N_3920);
nand U7065 (N_7065,N_2898,N_4095);
and U7066 (N_7066,N_4064,N_2585);
or U7067 (N_7067,N_2830,N_4109);
or U7068 (N_7068,N_2568,N_3653);
or U7069 (N_7069,N_3956,N_4213);
nor U7070 (N_7070,N_2873,N_4495);
xnor U7071 (N_7071,N_4158,N_4219);
xnor U7072 (N_7072,N_4452,N_3586);
nand U7073 (N_7073,N_4192,N_3215);
nand U7074 (N_7074,N_4606,N_3758);
or U7075 (N_7075,N_3976,N_4002);
xnor U7076 (N_7076,N_4467,N_4306);
xnor U7077 (N_7077,N_4440,N_4635);
or U7078 (N_7078,N_2994,N_2507);
and U7079 (N_7079,N_3693,N_4522);
or U7080 (N_7080,N_3521,N_2996);
nand U7081 (N_7081,N_3435,N_4385);
xor U7082 (N_7082,N_4778,N_4966);
and U7083 (N_7083,N_3191,N_3446);
nand U7084 (N_7084,N_4153,N_3695);
xor U7085 (N_7085,N_4775,N_4037);
and U7086 (N_7086,N_3769,N_4141);
nand U7087 (N_7087,N_3572,N_4043);
nand U7088 (N_7088,N_3094,N_2569);
nor U7089 (N_7089,N_4212,N_3912);
nor U7090 (N_7090,N_2766,N_4170);
and U7091 (N_7091,N_4590,N_4897);
or U7092 (N_7092,N_4524,N_4268);
nor U7093 (N_7093,N_4911,N_2933);
nor U7094 (N_7094,N_2824,N_3753);
nand U7095 (N_7095,N_4948,N_3272);
or U7096 (N_7096,N_3108,N_2575);
xor U7097 (N_7097,N_3262,N_3132);
nor U7098 (N_7098,N_3866,N_3380);
nand U7099 (N_7099,N_3928,N_2857);
or U7100 (N_7100,N_4118,N_3256);
and U7101 (N_7101,N_4326,N_3971);
nor U7102 (N_7102,N_2638,N_3018);
nand U7103 (N_7103,N_4391,N_4800);
nand U7104 (N_7104,N_3397,N_4686);
nor U7105 (N_7105,N_3987,N_3472);
xnor U7106 (N_7106,N_2789,N_3540);
and U7107 (N_7107,N_2613,N_3363);
xnor U7108 (N_7108,N_3842,N_4791);
xor U7109 (N_7109,N_4174,N_3560);
nor U7110 (N_7110,N_4577,N_3412);
or U7111 (N_7111,N_4763,N_3298);
nor U7112 (N_7112,N_3397,N_4349);
and U7113 (N_7113,N_2858,N_3075);
xor U7114 (N_7114,N_3543,N_4826);
nand U7115 (N_7115,N_2764,N_2958);
nand U7116 (N_7116,N_4197,N_4718);
and U7117 (N_7117,N_3222,N_4685);
nor U7118 (N_7118,N_3392,N_2761);
nand U7119 (N_7119,N_4936,N_4385);
or U7120 (N_7120,N_3668,N_2994);
nand U7121 (N_7121,N_3475,N_4861);
nand U7122 (N_7122,N_4128,N_4352);
nand U7123 (N_7123,N_3388,N_2959);
nor U7124 (N_7124,N_4094,N_4146);
nor U7125 (N_7125,N_4508,N_4271);
nand U7126 (N_7126,N_2536,N_3594);
xnor U7127 (N_7127,N_3623,N_4468);
or U7128 (N_7128,N_2904,N_3058);
or U7129 (N_7129,N_4889,N_2999);
xnor U7130 (N_7130,N_3934,N_4830);
and U7131 (N_7131,N_3664,N_4137);
or U7132 (N_7132,N_3145,N_4385);
and U7133 (N_7133,N_2823,N_3478);
or U7134 (N_7134,N_4737,N_3014);
and U7135 (N_7135,N_2953,N_2529);
nor U7136 (N_7136,N_2762,N_3232);
xnor U7137 (N_7137,N_2700,N_4706);
nor U7138 (N_7138,N_2745,N_4133);
nand U7139 (N_7139,N_3860,N_4527);
nor U7140 (N_7140,N_2573,N_4164);
xnor U7141 (N_7141,N_4343,N_4945);
xnor U7142 (N_7142,N_3513,N_2998);
nor U7143 (N_7143,N_3896,N_3172);
nand U7144 (N_7144,N_3829,N_4596);
and U7145 (N_7145,N_2769,N_2722);
nor U7146 (N_7146,N_2599,N_4249);
nor U7147 (N_7147,N_3904,N_4299);
xnor U7148 (N_7148,N_4329,N_2995);
nor U7149 (N_7149,N_3552,N_4369);
nor U7150 (N_7150,N_4507,N_4942);
xor U7151 (N_7151,N_3337,N_4782);
xor U7152 (N_7152,N_3515,N_3046);
nand U7153 (N_7153,N_3748,N_2823);
nor U7154 (N_7154,N_2719,N_4157);
nand U7155 (N_7155,N_2621,N_4652);
nor U7156 (N_7156,N_2506,N_4956);
and U7157 (N_7157,N_4080,N_4747);
nor U7158 (N_7158,N_3958,N_2880);
xnor U7159 (N_7159,N_3994,N_3524);
xnor U7160 (N_7160,N_4413,N_4471);
xor U7161 (N_7161,N_3052,N_4818);
or U7162 (N_7162,N_4980,N_2811);
nand U7163 (N_7163,N_2531,N_4830);
nor U7164 (N_7164,N_3559,N_2885);
or U7165 (N_7165,N_4262,N_3499);
xnor U7166 (N_7166,N_4600,N_3539);
and U7167 (N_7167,N_2536,N_4074);
xnor U7168 (N_7168,N_2864,N_3731);
and U7169 (N_7169,N_2637,N_3890);
and U7170 (N_7170,N_2978,N_3089);
or U7171 (N_7171,N_2969,N_4059);
nor U7172 (N_7172,N_2719,N_3041);
nand U7173 (N_7173,N_4623,N_3671);
nand U7174 (N_7174,N_3081,N_2507);
nand U7175 (N_7175,N_4973,N_3155);
nor U7176 (N_7176,N_3686,N_2945);
xnor U7177 (N_7177,N_4743,N_3660);
nor U7178 (N_7178,N_3850,N_3701);
nand U7179 (N_7179,N_2944,N_2523);
and U7180 (N_7180,N_3388,N_3804);
nor U7181 (N_7181,N_3177,N_4707);
and U7182 (N_7182,N_4460,N_3157);
nand U7183 (N_7183,N_3442,N_3948);
xor U7184 (N_7184,N_3304,N_4302);
or U7185 (N_7185,N_4342,N_4612);
nor U7186 (N_7186,N_4224,N_3844);
nor U7187 (N_7187,N_4939,N_4472);
and U7188 (N_7188,N_3926,N_4056);
xnor U7189 (N_7189,N_4680,N_3477);
nand U7190 (N_7190,N_3798,N_4702);
nor U7191 (N_7191,N_4304,N_3533);
nor U7192 (N_7192,N_3508,N_3883);
and U7193 (N_7193,N_4935,N_2904);
nand U7194 (N_7194,N_3412,N_3975);
and U7195 (N_7195,N_4028,N_4782);
xnor U7196 (N_7196,N_2702,N_2619);
xnor U7197 (N_7197,N_4474,N_4993);
and U7198 (N_7198,N_4185,N_4826);
nor U7199 (N_7199,N_4536,N_3875);
or U7200 (N_7200,N_2826,N_4931);
and U7201 (N_7201,N_4563,N_2838);
nand U7202 (N_7202,N_3953,N_3008);
or U7203 (N_7203,N_4902,N_2560);
or U7204 (N_7204,N_2875,N_2693);
nor U7205 (N_7205,N_2611,N_3973);
and U7206 (N_7206,N_3801,N_2869);
nor U7207 (N_7207,N_2925,N_4946);
xnor U7208 (N_7208,N_4923,N_2698);
nor U7209 (N_7209,N_2892,N_4907);
or U7210 (N_7210,N_3571,N_3433);
nand U7211 (N_7211,N_3118,N_3614);
or U7212 (N_7212,N_3722,N_4683);
nand U7213 (N_7213,N_3333,N_2614);
nand U7214 (N_7214,N_4522,N_3318);
xor U7215 (N_7215,N_4504,N_4179);
or U7216 (N_7216,N_4357,N_4545);
nor U7217 (N_7217,N_3235,N_2880);
or U7218 (N_7218,N_4894,N_3057);
nor U7219 (N_7219,N_4925,N_3165);
nand U7220 (N_7220,N_2668,N_4085);
xnor U7221 (N_7221,N_3562,N_4918);
nand U7222 (N_7222,N_3967,N_4691);
nand U7223 (N_7223,N_3005,N_3724);
nand U7224 (N_7224,N_4199,N_3310);
and U7225 (N_7225,N_2523,N_3462);
and U7226 (N_7226,N_4305,N_3272);
nand U7227 (N_7227,N_4972,N_3795);
or U7228 (N_7228,N_3520,N_3900);
xnor U7229 (N_7229,N_4290,N_3258);
or U7230 (N_7230,N_4168,N_2501);
or U7231 (N_7231,N_3181,N_2825);
nor U7232 (N_7232,N_4520,N_4447);
and U7233 (N_7233,N_2586,N_3762);
xor U7234 (N_7234,N_4082,N_3903);
nand U7235 (N_7235,N_3029,N_4353);
and U7236 (N_7236,N_3322,N_4297);
or U7237 (N_7237,N_3633,N_2811);
and U7238 (N_7238,N_2520,N_2638);
nor U7239 (N_7239,N_4965,N_3113);
nor U7240 (N_7240,N_3502,N_4537);
nand U7241 (N_7241,N_4259,N_4134);
or U7242 (N_7242,N_4101,N_3555);
or U7243 (N_7243,N_4536,N_4992);
nand U7244 (N_7244,N_3798,N_3590);
nor U7245 (N_7245,N_2661,N_3710);
or U7246 (N_7246,N_2728,N_3641);
and U7247 (N_7247,N_3806,N_3627);
xnor U7248 (N_7248,N_4211,N_2803);
nand U7249 (N_7249,N_3406,N_4573);
nor U7250 (N_7250,N_3092,N_3320);
or U7251 (N_7251,N_2671,N_4786);
and U7252 (N_7252,N_4879,N_3822);
xnor U7253 (N_7253,N_3194,N_3925);
nor U7254 (N_7254,N_2565,N_2864);
nor U7255 (N_7255,N_2778,N_3395);
nand U7256 (N_7256,N_4628,N_3246);
nor U7257 (N_7257,N_4406,N_4184);
nor U7258 (N_7258,N_4310,N_4910);
xnor U7259 (N_7259,N_3255,N_3098);
and U7260 (N_7260,N_2965,N_4993);
or U7261 (N_7261,N_3800,N_3570);
xnor U7262 (N_7262,N_4723,N_2948);
nand U7263 (N_7263,N_3233,N_2729);
nor U7264 (N_7264,N_3344,N_4030);
nor U7265 (N_7265,N_3397,N_2739);
and U7266 (N_7266,N_3758,N_4091);
nor U7267 (N_7267,N_4473,N_2593);
nor U7268 (N_7268,N_4494,N_4695);
nand U7269 (N_7269,N_3636,N_4463);
nand U7270 (N_7270,N_4938,N_4043);
nand U7271 (N_7271,N_2784,N_4042);
and U7272 (N_7272,N_4510,N_2912);
and U7273 (N_7273,N_4959,N_2806);
nand U7274 (N_7274,N_4160,N_4580);
or U7275 (N_7275,N_3112,N_4202);
nand U7276 (N_7276,N_4458,N_2877);
or U7277 (N_7277,N_4906,N_3330);
nand U7278 (N_7278,N_3745,N_2561);
xnor U7279 (N_7279,N_2631,N_3626);
nor U7280 (N_7280,N_4234,N_3756);
nor U7281 (N_7281,N_4504,N_3922);
nor U7282 (N_7282,N_3264,N_2521);
and U7283 (N_7283,N_3696,N_4127);
xnor U7284 (N_7284,N_2715,N_3451);
nand U7285 (N_7285,N_4633,N_4161);
nor U7286 (N_7286,N_4843,N_4572);
and U7287 (N_7287,N_2721,N_3070);
or U7288 (N_7288,N_4992,N_3392);
and U7289 (N_7289,N_4196,N_3381);
nand U7290 (N_7290,N_4558,N_2647);
or U7291 (N_7291,N_3236,N_3708);
and U7292 (N_7292,N_2876,N_3403);
xor U7293 (N_7293,N_2502,N_4344);
and U7294 (N_7294,N_4347,N_4173);
and U7295 (N_7295,N_3477,N_3474);
or U7296 (N_7296,N_3052,N_3037);
nand U7297 (N_7297,N_2652,N_4501);
xnor U7298 (N_7298,N_3013,N_3716);
and U7299 (N_7299,N_2617,N_4398);
nand U7300 (N_7300,N_3074,N_4517);
xor U7301 (N_7301,N_4031,N_4721);
and U7302 (N_7302,N_4524,N_2753);
nor U7303 (N_7303,N_2976,N_3215);
nand U7304 (N_7304,N_3969,N_3237);
nor U7305 (N_7305,N_3578,N_3545);
and U7306 (N_7306,N_3647,N_3585);
or U7307 (N_7307,N_2950,N_4301);
and U7308 (N_7308,N_2944,N_4413);
xor U7309 (N_7309,N_3723,N_3826);
xnor U7310 (N_7310,N_4338,N_2738);
nor U7311 (N_7311,N_3849,N_3032);
and U7312 (N_7312,N_3592,N_3199);
and U7313 (N_7313,N_3670,N_3918);
nor U7314 (N_7314,N_2556,N_3384);
xor U7315 (N_7315,N_2524,N_4675);
and U7316 (N_7316,N_4106,N_4381);
nand U7317 (N_7317,N_2859,N_3230);
and U7318 (N_7318,N_3494,N_3202);
xnor U7319 (N_7319,N_2983,N_4111);
xnor U7320 (N_7320,N_4908,N_2524);
or U7321 (N_7321,N_3943,N_3305);
xnor U7322 (N_7322,N_2693,N_2626);
or U7323 (N_7323,N_2500,N_3330);
nand U7324 (N_7324,N_3326,N_4822);
or U7325 (N_7325,N_3332,N_3249);
or U7326 (N_7326,N_4432,N_4797);
nand U7327 (N_7327,N_4069,N_4849);
or U7328 (N_7328,N_2501,N_3292);
or U7329 (N_7329,N_2547,N_2784);
or U7330 (N_7330,N_4740,N_4671);
xnor U7331 (N_7331,N_2539,N_4637);
nor U7332 (N_7332,N_4850,N_4513);
nand U7333 (N_7333,N_4574,N_2662);
nor U7334 (N_7334,N_4229,N_2678);
nor U7335 (N_7335,N_2968,N_3198);
or U7336 (N_7336,N_3023,N_3376);
or U7337 (N_7337,N_2508,N_3566);
and U7338 (N_7338,N_2968,N_4351);
nor U7339 (N_7339,N_3637,N_4925);
xor U7340 (N_7340,N_4652,N_2810);
nand U7341 (N_7341,N_4652,N_4933);
xnor U7342 (N_7342,N_4443,N_4745);
nor U7343 (N_7343,N_3078,N_4284);
and U7344 (N_7344,N_3926,N_4574);
and U7345 (N_7345,N_3105,N_3932);
and U7346 (N_7346,N_4504,N_3325);
nor U7347 (N_7347,N_3748,N_4371);
xnor U7348 (N_7348,N_4156,N_3352);
and U7349 (N_7349,N_3919,N_2885);
nor U7350 (N_7350,N_3357,N_4041);
xor U7351 (N_7351,N_3220,N_4139);
xor U7352 (N_7352,N_4662,N_2587);
nand U7353 (N_7353,N_2563,N_3658);
nand U7354 (N_7354,N_3648,N_2915);
nand U7355 (N_7355,N_3861,N_3690);
nand U7356 (N_7356,N_3891,N_2997);
or U7357 (N_7357,N_2870,N_4395);
nor U7358 (N_7358,N_4574,N_2891);
xnor U7359 (N_7359,N_3292,N_3402);
nor U7360 (N_7360,N_4531,N_2513);
and U7361 (N_7361,N_3770,N_4023);
or U7362 (N_7362,N_2736,N_4914);
and U7363 (N_7363,N_2657,N_3966);
or U7364 (N_7364,N_3913,N_4019);
xor U7365 (N_7365,N_3482,N_4088);
xor U7366 (N_7366,N_4545,N_2525);
nand U7367 (N_7367,N_3310,N_4032);
nor U7368 (N_7368,N_4727,N_2569);
or U7369 (N_7369,N_3329,N_4352);
and U7370 (N_7370,N_3112,N_4325);
or U7371 (N_7371,N_4501,N_4304);
and U7372 (N_7372,N_3543,N_4999);
and U7373 (N_7373,N_4793,N_3025);
nor U7374 (N_7374,N_3402,N_2524);
and U7375 (N_7375,N_2684,N_3729);
or U7376 (N_7376,N_4388,N_4124);
or U7377 (N_7377,N_3611,N_4088);
nor U7378 (N_7378,N_2724,N_4524);
nand U7379 (N_7379,N_3221,N_4795);
nor U7380 (N_7380,N_3093,N_4329);
nor U7381 (N_7381,N_4103,N_3914);
xor U7382 (N_7382,N_4140,N_2522);
nor U7383 (N_7383,N_3044,N_2920);
or U7384 (N_7384,N_2773,N_4087);
nor U7385 (N_7385,N_2856,N_3239);
nand U7386 (N_7386,N_3663,N_2743);
nor U7387 (N_7387,N_4854,N_3524);
or U7388 (N_7388,N_4939,N_4272);
nor U7389 (N_7389,N_2943,N_3596);
xor U7390 (N_7390,N_4322,N_3480);
nor U7391 (N_7391,N_4422,N_2803);
or U7392 (N_7392,N_4721,N_3383);
xor U7393 (N_7393,N_4694,N_4070);
nor U7394 (N_7394,N_3358,N_3048);
or U7395 (N_7395,N_4491,N_2853);
and U7396 (N_7396,N_3587,N_3323);
nand U7397 (N_7397,N_4249,N_4030);
nor U7398 (N_7398,N_3634,N_4517);
nand U7399 (N_7399,N_4886,N_4017);
xor U7400 (N_7400,N_4867,N_3537);
or U7401 (N_7401,N_4281,N_4260);
or U7402 (N_7402,N_3754,N_3586);
and U7403 (N_7403,N_2826,N_4057);
or U7404 (N_7404,N_3029,N_3870);
and U7405 (N_7405,N_3019,N_3932);
and U7406 (N_7406,N_4555,N_4639);
or U7407 (N_7407,N_2663,N_4662);
and U7408 (N_7408,N_2807,N_4527);
nand U7409 (N_7409,N_4403,N_4752);
and U7410 (N_7410,N_3309,N_3865);
nand U7411 (N_7411,N_2565,N_3733);
xnor U7412 (N_7412,N_3606,N_4987);
and U7413 (N_7413,N_3071,N_2869);
and U7414 (N_7414,N_2520,N_4849);
or U7415 (N_7415,N_2643,N_3963);
nor U7416 (N_7416,N_4206,N_4065);
or U7417 (N_7417,N_2960,N_3530);
nor U7418 (N_7418,N_4054,N_3996);
or U7419 (N_7419,N_2769,N_3259);
and U7420 (N_7420,N_2804,N_2896);
and U7421 (N_7421,N_2699,N_3527);
xnor U7422 (N_7422,N_3547,N_4265);
or U7423 (N_7423,N_4511,N_4435);
nand U7424 (N_7424,N_2734,N_4133);
xnor U7425 (N_7425,N_3762,N_2615);
nand U7426 (N_7426,N_4645,N_4194);
xnor U7427 (N_7427,N_3169,N_3128);
nor U7428 (N_7428,N_3723,N_2525);
or U7429 (N_7429,N_3453,N_3099);
and U7430 (N_7430,N_4301,N_4409);
nor U7431 (N_7431,N_3090,N_3135);
xor U7432 (N_7432,N_2808,N_3257);
nor U7433 (N_7433,N_4726,N_3752);
nor U7434 (N_7434,N_3268,N_4496);
nor U7435 (N_7435,N_3042,N_4753);
xor U7436 (N_7436,N_4307,N_4073);
nand U7437 (N_7437,N_4466,N_4592);
and U7438 (N_7438,N_4603,N_3864);
nor U7439 (N_7439,N_2508,N_3833);
xor U7440 (N_7440,N_3456,N_2723);
xor U7441 (N_7441,N_4659,N_4770);
nand U7442 (N_7442,N_3423,N_3649);
nand U7443 (N_7443,N_3599,N_2874);
xnor U7444 (N_7444,N_2529,N_4208);
nor U7445 (N_7445,N_4385,N_4139);
and U7446 (N_7446,N_2954,N_3850);
or U7447 (N_7447,N_4009,N_4317);
xor U7448 (N_7448,N_3985,N_3681);
and U7449 (N_7449,N_3524,N_3819);
or U7450 (N_7450,N_3583,N_3626);
xor U7451 (N_7451,N_2913,N_4383);
or U7452 (N_7452,N_4895,N_4341);
xnor U7453 (N_7453,N_4299,N_4412);
xor U7454 (N_7454,N_4520,N_3601);
nor U7455 (N_7455,N_3364,N_4713);
or U7456 (N_7456,N_4115,N_3404);
or U7457 (N_7457,N_3523,N_4916);
nor U7458 (N_7458,N_3119,N_2865);
and U7459 (N_7459,N_4139,N_3240);
or U7460 (N_7460,N_3789,N_4395);
and U7461 (N_7461,N_4684,N_3669);
and U7462 (N_7462,N_3298,N_2657);
and U7463 (N_7463,N_3610,N_4792);
or U7464 (N_7464,N_2843,N_3964);
and U7465 (N_7465,N_2601,N_4759);
nor U7466 (N_7466,N_4315,N_4916);
or U7467 (N_7467,N_3668,N_4290);
and U7468 (N_7468,N_3296,N_4912);
and U7469 (N_7469,N_4803,N_4748);
or U7470 (N_7470,N_3674,N_2682);
and U7471 (N_7471,N_2726,N_4014);
xnor U7472 (N_7472,N_3173,N_4242);
or U7473 (N_7473,N_4435,N_4718);
or U7474 (N_7474,N_2768,N_4277);
xnor U7475 (N_7475,N_4506,N_3116);
or U7476 (N_7476,N_3669,N_3440);
and U7477 (N_7477,N_3029,N_3768);
and U7478 (N_7478,N_4058,N_3444);
or U7479 (N_7479,N_3889,N_3667);
or U7480 (N_7480,N_4493,N_4735);
or U7481 (N_7481,N_4635,N_2752);
nor U7482 (N_7482,N_4983,N_4988);
xor U7483 (N_7483,N_3678,N_3117);
xor U7484 (N_7484,N_3066,N_2702);
xnor U7485 (N_7485,N_4811,N_3511);
nor U7486 (N_7486,N_3962,N_4138);
and U7487 (N_7487,N_3049,N_2593);
or U7488 (N_7488,N_4289,N_3304);
nand U7489 (N_7489,N_4740,N_2994);
or U7490 (N_7490,N_2886,N_2796);
nand U7491 (N_7491,N_2508,N_2636);
nor U7492 (N_7492,N_3905,N_4574);
nor U7493 (N_7493,N_4635,N_2692);
xnor U7494 (N_7494,N_4218,N_3574);
nand U7495 (N_7495,N_4229,N_3468);
or U7496 (N_7496,N_3540,N_3493);
nor U7497 (N_7497,N_3377,N_4773);
nor U7498 (N_7498,N_3418,N_3893);
nor U7499 (N_7499,N_3928,N_3850);
xnor U7500 (N_7500,N_5123,N_7096);
nor U7501 (N_7501,N_6199,N_6283);
or U7502 (N_7502,N_6439,N_5351);
xnor U7503 (N_7503,N_7064,N_6751);
or U7504 (N_7504,N_5155,N_6104);
xor U7505 (N_7505,N_6264,N_7146);
or U7506 (N_7506,N_5931,N_7321);
nor U7507 (N_7507,N_7311,N_5977);
and U7508 (N_7508,N_7115,N_5450);
xnor U7509 (N_7509,N_5554,N_5688);
nor U7510 (N_7510,N_7305,N_5367);
and U7511 (N_7511,N_6643,N_7280);
xnor U7512 (N_7512,N_7150,N_5836);
xor U7513 (N_7513,N_6685,N_6630);
nand U7514 (N_7514,N_5006,N_5508);
and U7515 (N_7515,N_6143,N_7273);
and U7516 (N_7516,N_5192,N_5734);
nor U7517 (N_7517,N_6815,N_5899);
nor U7518 (N_7518,N_7034,N_5762);
nand U7519 (N_7519,N_7399,N_5505);
nor U7520 (N_7520,N_5622,N_6581);
and U7521 (N_7521,N_5736,N_5510);
nor U7522 (N_7522,N_5991,N_5541);
or U7523 (N_7523,N_5781,N_6835);
xor U7524 (N_7524,N_5612,N_5267);
nand U7525 (N_7525,N_5535,N_5002);
or U7526 (N_7526,N_5520,N_5865);
or U7527 (N_7527,N_5513,N_5840);
and U7528 (N_7528,N_5237,N_6267);
xnor U7529 (N_7529,N_5335,N_6065);
xor U7530 (N_7530,N_5570,N_5858);
nor U7531 (N_7531,N_5043,N_6524);
nor U7532 (N_7532,N_6902,N_5708);
nor U7533 (N_7533,N_5031,N_6301);
xnor U7534 (N_7534,N_6183,N_5700);
xnor U7535 (N_7535,N_6971,N_5608);
nor U7536 (N_7536,N_5221,N_6704);
nand U7537 (N_7537,N_5739,N_6466);
nand U7538 (N_7538,N_6378,N_5414);
and U7539 (N_7539,N_5423,N_7038);
nand U7540 (N_7540,N_6872,N_6450);
nor U7541 (N_7541,N_6540,N_5299);
xor U7542 (N_7542,N_5584,N_6443);
xnor U7543 (N_7543,N_5086,N_6913);
xor U7544 (N_7544,N_6693,N_7429);
or U7545 (N_7545,N_7239,N_5907);
nor U7546 (N_7546,N_7075,N_6401);
or U7547 (N_7547,N_6613,N_5302);
xor U7548 (N_7548,N_7380,N_5326);
xnor U7549 (N_7549,N_6232,N_5764);
xnor U7550 (N_7550,N_5240,N_7136);
or U7551 (N_7551,N_5293,N_6603);
nor U7552 (N_7552,N_5112,N_5916);
nand U7553 (N_7553,N_7308,N_5782);
or U7554 (N_7554,N_5814,N_7194);
nor U7555 (N_7555,N_5507,N_7293);
xnor U7556 (N_7556,N_5895,N_7095);
and U7557 (N_7557,N_5312,N_7379);
xor U7558 (N_7558,N_7411,N_5184);
xnor U7559 (N_7559,N_5376,N_5362);
and U7560 (N_7560,N_5677,N_5021);
xnor U7561 (N_7561,N_5853,N_6438);
nand U7562 (N_7562,N_5429,N_7483);
nand U7563 (N_7563,N_5494,N_5911);
nor U7564 (N_7564,N_6492,N_6873);
or U7565 (N_7565,N_6729,N_6719);
xnor U7566 (N_7566,N_6277,N_6561);
and U7567 (N_7567,N_6817,N_6593);
xor U7568 (N_7568,N_5170,N_7487);
or U7569 (N_7569,N_6149,N_7430);
or U7570 (N_7570,N_5973,N_6521);
and U7571 (N_7571,N_7418,N_6255);
xnor U7572 (N_7572,N_5971,N_5649);
nor U7573 (N_7573,N_7477,N_6698);
or U7574 (N_7574,N_5648,N_6186);
or U7575 (N_7575,N_5859,N_6976);
nand U7576 (N_7576,N_6319,N_7207);
nor U7577 (N_7577,N_5551,N_5458);
nor U7578 (N_7578,N_6753,N_6477);
nand U7579 (N_7579,N_5871,N_6457);
nand U7580 (N_7580,N_7147,N_5442);
and U7581 (N_7581,N_6615,N_5877);
nor U7582 (N_7582,N_6080,N_5862);
nand U7583 (N_7583,N_6249,N_5193);
and U7584 (N_7584,N_7154,N_7347);
nand U7585 (N_7585,N_6800,N_7404);
xnor U7586 (N_7586,N_6054,N_6335);
xnor U7587 (N_7587,N_5477,N_5214);
and U7588 (N_7588,N_6625,N_5425);
nand U7589 (N_7589,N_7359,N_6519);
nor U7590 (N_7590,N_6985,N_5091);
or U7591 (N_7591,N_5107,N_5157);
xnor U7592 (N_7592,N_7310,N_5845);
or U7593 (N_7593,N_7468,N_6629);
or U7594 (N_7594,N_6922,N_6589);
nand U7595 (N_7595,N_5744,N_6906);
or U7596 (N_7596,N_6274,N_6946);
nand U7597 (N_7597,N_5875,N_5227);
nand U7598 (N_7598,N_7386,N_6898);
nor U7599 (N_7599,N_5276,N_6127);
nand U7600 (N_7600,N_6454,N_6317);
nor U7601 (N_7601,N_5571,N_6330);
nor U7602 (N_7602,N_6992,N_6395);
nor U7603 (N_7603,N_5891,N_6265);
or U7604 (N_7604,N_5111,N_6484);
xnor U7605 (N_7605,N_5523,N_5357);
or U7606 (N_7606,N_5934,N_5947);
nand U7607 (N_7607,N_5495,N_5786);
xnor U7608 (N_7608,N_6494,N_5345);
nor U7609 (N_7609,N_5999,N_6754);
and U7610 (N_7610,N_7345,N_6056);
or U7611 (N_7611,N_7159,N_6688);
nor U7612 (N_7612,N_5469,N_5933);
or U7613 (N_7613,N_5745,N_5359);
xor U7614 (N_7614,N_5272,N_5851);
or U7615 (N_7615,N_6787,N_5893);
nand U7616 (N_7616,N_6113,N_6293);
and U7617 (N_7617,N_6522,N_5939);
and U7618 (N_7618,N_5219,N_7098);
or U7619 (N_7619,N_7161,N_7103);
or U7620 (N_7620,N_5210,N_6597);
nor U7621 (N_7621,N_5472,N_6322);
nor U7622 (N_7622,N_7303,N_6558);
or U7623 (N_7623,N_5471,N_6649);
nand U7624 (N_7624,N_5905,N_5779);
and U7625 (N_7625,N_5595,N_7447);
and U7626 (N_7626,N_5106,N_6196);
and U7627 (N_7627,N_7274,N_5810);
and U7628 (N_7628,N_7340,N_5743);
or U7629 (N_7629,N_6633,N_6708);
xnor U7630 (N_7630,N_6563,N_7058);
or U7631 (N_7631,N_7223,N_6642);
and U7632 (N_7632,N_6099,N_5169);
or U7633 (N_7633,N_7383,N_7391);
nand U7634 (N_7634,N_6346,N_6987);
nor U7635 (N_7635,N_6115,N_7489);
nand U7636 (N_7636,N_5678,N_7290);
nand U7637 (N_7637,N_7461,N_7426);
and U7638 (N_7638,N_7334,N_5249);
and U7639 (N_7639,N_7382,N_5640);
xnor U7640 (N_7640,N_7494,N_5398);
xnor U7641 (N_7641,N_5147,N_6570);
nand U7642 (N_7642,N_5830,N_6647);
xnor U7643 (N_7643,N_5569,N_5572);
nor U7644 (N_7644,N_6308,N_5360);
xnor U7645 (N_7645,N_5912,N_6388);
and U7646 (N_7646,N_5672,N_7476);
xor U7647 (N_7647,N_6098,N_6179);
or U7648 (N_7648,N_5248,N_5509);
xor U7649 (N_7649,N_6961,N_7165);
nand U7650 (N_7650,N_7116,N_6081);
and U7651 (N_7651,N_6152,N_7271);
nor U7652 (N_7652,N_6877,N_6211);
nor U7653 (N_7653,N_5839,N_6072);
nor U7654 (N_7654,N_6057,N_5396);
and U7655 (N_7655,N_5431,N_7142);
xnor U7656 (N_7656,N_6997,N_7080);
xnor U7657 (N_7657,N_7145,N_7229);
and U7658 (N_7658,N_6654,N_5987);
xnor U7659 (N_7659,N_6447,N_6053);
nor U7660 (N_7660,N_5778,N_7173);
nand U7661 (N_7661,N_7330,N_5769);
and U7662 (N_7662,N_6448,N_6444);
or U7663 (N_7663,N_5946,N_5522);
or U7664 (N_7664,N_5497,N_7104);
xnor U7665 (N_7665,N_5110,N_6914);
nand U7666 (N_7666,N_5481,N_5553);
nand U7667 (N_7667,N_5149,N_5646);
and U7668 (N_7668,N_6016,N_5488);
nand U7669 (N_7669,N_5186,N_6910);
and U7670 (N_7670,N_7414,N_5888);
nand U7671 (N_7671,N_7451,N_6969);
nand U7672 (N_7672,N_5255,N_5320);
or U7673 (N_7673,N_7130,N_6320);
nor U7674 (N_7674,N_6943,N_5329);
nor U7675 (N_7675,N_7008,N_5462);
and U7676 (N_7676,N_6370,N_6890);
xor U7677 (N_7677,N_5651,N_5856);
xor U7678 (N_7678,N_7067,N_6187);
nor U7679 (N_7679,N_7059,N_5883);
and U7680 (N_7680,N_6495,N_6701);
nor U7681 (N_7681,N_6758,N_6036);
xnor U7682 (N_7682,N_6281,N_5078);
nor U7683 (N_7683,N_6528,N_5115);
nor U7684 (N_7684,N_6634,N_5041);
nor U7685 (N_7685,N_7247,N_5948);
xor U7686 (N_7686,N_6402,N_5670);
xnor U7687 (N_7687,N_7295,N_6584);
xor U7688 (N_7688,N_7433,N_5722);
nand U7689 (N_7689,N_5775,N_7195);
xor U7690 (N_7690,N_6692,N_6614);
and U7691 (N_7691,N_7302,N_5172);
or U7692 (N_7692,N_6657,N_5981);
or U7693 (N_7693,N_6555,N_6476);
or U7694 (N_7694,N_6923,N_6793);
or U7695 (N_7695,N_7301,N_5354);
nor U7696 (N_7696,N_6208,N_6653);
and U7697 (N_7697,N_6605,N_5323);
nor U7698 (N_7698,N_6210,N_7373);
and U7699 (N_7699,N_6203,N_6215);
xnor U7700 (N_7700,N_5310,N_6844);
xor U7701 (N_7701,N_6911,N_6327);
nor U7702 (N_7702,N_6357,N_6938);
nor U7703 (N_7703,N_7360,N_5198);
nand U7704 (N_7704,N_6690,N_5464);
nand U7705 (N_7705,N_5604,N_7389);
and U7706 (N_7706,N_6188,N_7422);
nor U7707 (N_7707,N_5521,N_7263);
nor U7708 (N_7708,N_6518,N_6193);
nand U7709 (N_7709,N_6512,N_6046);
nand U7710 (N_7710,N_6422,N_6921);
and U7711 (N_7711,N_5783,N_6001);
nor U7712 (N_7712,N_6811,N_6172);
xor U7713 (N_7713,N_6768,N_5927);
or U7714 (N_7714,N_6766,N_5873);
or U7715 (N_7715,N_6334,N_7306);
and U7716 (N_7716,N_7498,N_5724);
xnor U7717 (N_7717,N_6393,N_5166);
or U7718 (N_7718,N_5846,N_5005);
or U7719 (N_7719,N_6156,N_5190);
nor U7720 (N_7720,N_6373,N_5487);
nor U7721 (N_7721,N_6082,N_7106);
or U7722 (N_7722,N_5140,N_5995);
nand U7723 (N_7723,N_6431,N_6602);
nor U7724 (N_7724,N_6529,N_7000);
nor U7725 (N_7725,N_6288,N_5832);
nand U7726 (N_7726,N_5099,N_5093);
nand U7727 (N_7727,N_7465,N_6383);
nor U7728 (N_7728,N_7090,N_6060);
and U7729 (N_7729,N_7289,N_5165);
nor U7730 (N_7730,N_6120,N_5673);
or U7731 (N_7731,N_6740,N_7358);
nor U7732 (N_7732,N_6869,N_5909);
xnor U7733 (N_7733,N_7419,N_7296);
xor U7734 (N_7734,N_5544,N_5686);
and U7735 (N_7735,N_7336,N_5038);
and U7736 (N_7736,N_6639,N_6441);
or U7737 (N_7737,N_6485,N_6066);
nor U7738 (N_7738,N_5387,N_5715);
nand U7739 (N_7739,N_5275,N_5558);
nand U7740 (N_7740,N_7457,N_6285);
xnor U7741 (N_7741,N_7438,N_5656);
or U7742 (N_7742,N_7252,N_7172);
nand U7743 (N_7743,N_7456,N_5930);
nand U7744 (N_7744,N_5784,N_7291);
nor U7745 (N_7745,N_6076,N_5375);
nor U7746 (N_7746,N_6313,N_5628);
or U7747 (N_7747,N_6445,N_6576);
xnor U7748 (N_7748,N_7108,N_6207);
nor U7749 (N_7749,N_6064,N_6631);
xnor U7750 (N_7750,N_5799,N_7472);
nand U7751 (N_7751,N_6842,N_6075);
xnor U7752 (N_7752,N_5056,N_6339);
nor U7753 (N_7753,N_7285,N_6089);
or U7754 (N_7754,N_7228,N_5615);
nor U7755 (N_7755,N_5108,N_5328);
and U7756 (N_7756,N_5459,N_6783);
nand U7757 (N_7757,N_7351,N_5261);
nor U7758 (N_7758,N_7026,N_7353);
xor U7759 (N_7759,N_6079,N_5908);
and U7760 (N_7760,N_5153,N_6325);
nand U7761 (N_7761,N_6471,N_6717);
or U7762 (N_7762,N_5607,N_5687);
nand U7763 (N_7763,N_5330,N_5511);
and U7764 (N_7764,N_5215,N_6045);
nor U7765 (N_7765,N_5904,N_5380);
nand U7766 (N_7766,N_6947,N_5674);
and U7767 (N_7767,N_5089,N_6318);
xnor U7768 (N_7768,N_6165,N_7240);
xnor U7769 (N_7769,N_6122,N_6509);
nand U7770 (N_7770,N_7315,N_6336);
xor U7771 (N_7771,N_6580,N_6718);
xnor U7772 (N_7772,N_5561,N_7188);
and U7773 (N_7773,N_5760,N_5366);
or U7774 (N_7774,N_5139,N_7220);
or U7775 (N_7775,N_6579,N_6983);
nor U7776 (N_7776,N_7467,N_6741);
nand U7777 (N_7777,N_6469,N_6233);
nor U7778 (N_7778,N_5207,N_6041);
nor U7779 (N_7779,N_6533,N_7237);
nor U7780 (N_7780,N_7078,N_6575);
nand U7781 (N_7781,N_6669,N_7062);
xnor U7782 (N_7782,N_5759,N_6531);
nand U7783 (N_7783,N_6350,N_7403);
xor U7784 (N_7784,N_5774,N_5493);
xnor U7785 (N_7785,N_5885,N_6909);
and U7786 (N_7786,N_5046,N_7342);
nand U7787 (N_7787,N_5447,N_7168);
nor U7788 (N_7788,N_7283,N_6564);
nor U7789 (N_7789,N_6356,N_6475);
nor U7790 (N_7790,N_5436,N_7163);
and U7791 (N_7791,N_6456,N_7299);
nand U7792 (N_7792,N_6377,N_7268);
nor U7793 (N_7793,N_6899,N_6414);
nand U7794 (N_7794,N_6884,N_7453);
or U7795 (N_7795,N_6731,N_7160);
and U7796 (N_7796,N_6147,N_6772);
or U7797 (N_7797,N_6744,N_6945);
xor U7798 (N_7798,N_6261,N_7431);
or U7799 (N_7799,N_7335,N_6604);
or U7800 (N_7800,N_5457,N_6358);
xnor U7801 (N_7801,N_5325,N_7029);
nand U7802 (N_7802,N_7117,N_6182);
and U7803 (N_7803,N_7152,N_5286);
nor U7804 (N_7804,N_6197,N_6962);
nand U7805 (N_7805,N_7089,N_6086);
nor U7806 (N_7806,N_6990,N_6472);
xnor U7807 (N_7807,N_5303,N_6506);
and U7808 (N_7808,N_5121,N_5684);
nor U7809 (N_7809,N_6146,N_5158);
and U7810 (N_7810,N_5298,N_7212);
nor U7811 (N_7811,N_5199,N_5151);
or U7812 (N_7812,N_5979,N_7475);
or U7813 (N_7813,N_6620,N_5805);
nand U7814 (N_7814,N_5412,N_6425);
nand U7815 (N_7815,N_6430,N_7164);
xnor U7816 (N_7816,N_5294,N_5009);
or U7817 (N_7817,N_5707,N_6617);
or U7818 (N_7818,N_6982,N_5564);
or U7819 (N_7819,N_6209,N_5653);
or U7820 (N_7820,N_6672,N_6903);
nor U7821 (N_7821,N_5938,N_6025);
and U7822 (N_7822,N_5590,N_6746);
or U7823 (N_7823,N_6515,N_6141);
xnor U7824 (N_7824,N_5800,N_5498);
and U7825 (N_7825,N_6090,N_6473);
xor U7826 (N_7826,N_6608,N_5034);
or U7827 (N_7827,N_5704,N_6360);
xor U7828 (N_7828,N_6889,N_6859);
nor U7829 (N_7829,N_5040,N_6040);
nor U7830 (N_7830,N_6458,N_6635);
xor U7831 (N_7831,N_6453,N_6668);
nand U7832 (N_7832,N_5780,N_6234);
and U7833 (N_7833,N_5465,N_5542);
nand U7834 (N_7834,N_6102,N_5940);
nand U7835 (N_7835,N_6520,N_6153);
nor U7836 (N_7836,N_6488,N_5892);
nand U7837 (N_7837,N_5660,N_6816);
nand U7838 (N_7838,N_5758,N_5452);
nand U7839 (N_7839,N_6640,N_6479);
or U7840 (N_7840,N_6765,N_5007);
nor U7841 (N_7841,N_6478,N_6256);
or U7842 (N_7842,N_5476,N_7462);
nor U7843 (N_7843,N_5338,N_6042);
or U7844 (N_7844,N_6100,N_5277);
and U7845 (N_7845,N_6932,N_5440);
nor U7846 (N_7846,N_5059,N_5378);
and U7847 (N_7847,N_6230,N_5141);
or U7848 (N_7848,N_5812,N_6324);
xor U7849 (N_7849,N_6435,N_5070);
nor U7850 (N_7850,N_6808,N_7409);
xor U7851 (N_7851,N_5787,N_7131);
or U7852 (N_7852,N_5563,N_7407);
and U7853 (N_7853,N_6006,N_6201);
or U7854 (N_7854,N_6023,N_6567);
nand U7855 (N_7855,N_5902,N_5596);
xor U7856 (N_7856,N_6830,N_5101);
nand U7857 (N_7857,N_6134,N_5388);
or U7858 (N_7858,N_5691,N_5071);
nand U7859 (N_7859,N_5096,N_5461);
and U7860 (N_7860,N_6737,N_5868);
and U7861 (N_7861,N_5116,N_5725);
xnor U7862 (N_7862,N_5284,N_5698);
and U7863 (N_7863,N_5755,N_5103);
or U7864 (N_7864,N_6725,N_6694);
nor U7865 (N_7865,N_6964,N_6467);
nand U7866 (N_7866,N_6862,N_7233);
xnor U7867 (N_7867,N_5234,N_6845);
or U7868 (N_7868,N_5316,N_5581);
or U7869 (N_7869,N_7074,N_6278);
xnor U7870 (N_7870,N_5950,N_5647);
and U7871 (N_7871,N_5582,N_6535);
nand U7872 (N_7872,N_7392,N_5247);
and U7873 (N_7873,N_5964,N_6761);
nor U7874 (N_7874,N_5454,N_7366);
nor U7875 (N_7875,N_5918,N_5777);
and U7876 (N_7876,N_6508,N_6497);
or U7877 (N_7877,N_5919,N_6131);
xor U7878 (N_7878,N_5641,N_5797);
and U7879 (N_7879,N_7191,N_5179);
xor U7880 (N_7880,N_7390,N_6756);
and U7881 (N_7881,N_5706,N_5194);
nand U7882 (N_7882,N_5057,N_6666);
nand U7883 (N_7883,N_5680,N_6005);
and U7884 (N_7884,N_6097,N_5183);
or U7885 (N_7885,N_6794,N_5424);
nand U7886 (N_7886,N_6534,N_6658);
or U7887 (N_7887,N_7063,N_5518);
and U7888 (N_7888,N_6651,N_6352);
xnor U7889 (N_7889,N_5568,N_6687);
and U7890 (N_7890,N_5420,N_5419);
and U7891 (N_7891,N_5529,N_5597);
xor U7892 (N_7892,N_5264,N_5125);
nand U7893 (N_7893,N_5746,N_7322);
xnor U7894 (N_7894,N_6219,N_5491);
and U7895 (N_7895,N_6245,N_5382);
xnor U7896 (N_7896,N_6895,N_5445);
and U7897 (N_7897,N_6118,N_6721);
xor U7898 (N_7898,N_5932,N_6771);
and U7899 (N_7899,N_6674,N_7046);
xor U7900 (N_7900,N_7143,N_6926);
nor U7901 (N_7901,N_7225,N_7129);
or U7902 (N_7902,N_5010,N_7425);
nand U7903 (N_7903,N_5716,N_6483);
nand U7904 (N_7904,N_6828,N_5478);
or U7905 (N_7905,N_5289,N_5747);
nand U7906 (N_7906,N_5854,N_6091);
and U7907 (N_7907,N_6979,N_5233);
nand U7908 (N_7908,N_5355,N_5557);
nand U7909 (N_7909,N_5976,N_5609);
nor U7910 (N_7910,N_6349,N_6601);
and U7911 (N_7911,N_7023,N_7434);
xor U7912 (N_7912,N_5980,N_6646);
or U7913 (N_7913,N_5404,N_5941);
xnor U7914 (N_7914,N_7236,N_6364);
or U7915 (N_7915,N_5258,N_7332);
xnor U7916 (N_7916,N_5524,N_7053);
or U7917 (N_7917,N_7428,N_7230);
xor U7918 (N_7918,N_5954,N_6585);
nor U7919 (N_7919,N_5681,N_5957);
xnor U7920 (N_7920,N_5291,N_5336);
or U7921 (N_7921,N_5882,N_6752);
xor U7922 (N_7922,N_5666,N_6019);
xor U7923 (N_7923,N_6367,N_7479);
and U7924 (N_7924,N_5339,N_6956);
and U7925 (N_7925,N_5699,N_5826);
xnor U7926 (N_7926,N_5663,N_5765);
nor U7927 (N_7927,N_7288,N_6764);
nand U7928 (N_7928,N_7370,N_5131);
or U7929 (N_7929,N_6386,N_5062);
xor U7930 (N_7930,N_5923,N_5257);
nand U7931 (N_7931,N_6517,N_5438);
or U7932 (N_7932,N_5978,N_5824);
xnor U7933 (N_7933,N_5128,N_6774);
xnor U7934 (N_7934,N_7348,N_7112);
nor U7935 (N_7935,N_6696,N_5566);
xnor U7936 (N_7936,N_7197,N_5280);
or U7937 (N_7937,N_6341,N_6437);
nor U7938 (N_7938,N_7329,N_5313);
xnor U7939 (N_7939,N_7208,N_5792);
xnor U7940 (N_7940,N_6482,N_7134);
nor U7941 (N_7941,N_7304,N_5421);
or U7942 (N_7942,N_6587,N_7174);
nor U7943 (N_7943,N_5771,N_6821);
or U7944 (N_7944,N_6825,N_5206);
or U7945 (N_7945,N_5889,N_5178);
xnor U7946 (N_7946,N_7454,N_6032);
and U7947 (N_7947,N_6121,N_7210);
or U7948 (N_7948,N_7258,N_5113);
or U7949 (N_7949,N_7242,N_7193);
nand U7950 (N_7950,N_6361,N_7056);
and U7951 (N_7951,N_5614,N_7003);
and U7952 (N_7952,N_6228,N_5334);
and U7953 (N_7953,N_6214,N_5573);
xnor U7954 (N_7954,N_5422,N_5547);
nor U7955 (N_7955,N_5742,N_5872);
and U7956 (N_7956,N_6148,N_6499);
xor U7957 (N_7957,N_7234,N_6018);
nor U7958 (N_7958,N_7372,N_6927);
or U7959 (N_7959,N_5230,N_5047);
nor U7960 (N_7960,N_5342,N_5504);
nand U7961 (N_7961,N_6296,N_6843);
and U7962 (N_7962,N_5023,N_5994);
xnor U7963 (N_7963,N_7109,N_5637);
or U7964 (N_7964,N_5966,N_7265);
and U7965 (N_7965,N_6407,N_5201);
or U7966 (N_7966,N_6807,N_6298);
xnor U7967 (N_7967,N_7297,N_7149);
or U7968 (N_7968,N_7044,N_7338);
nand U7969 (N_7969,N_6790,N_6770);
or U7970 (N_7970,N_5019,N_6415);
nor U7971 (N_7971,N_5229,N_6136);
and U7972 (N_7972,N_5801,N_6857);
and U7973 (N_7973,N_6596,N_6954);
or U7974 (N_7974,N_6837,N_6714);
nand U7975 (N_7975,N_7460,N_7097);
or U7976 (N_7976,N_7226,N_5446);
nor U7977 (N_7977,N_5097,N_5848);
xor U7978 (N_7978,N_5444,N_5161);
nor U7979 (N_7979,N_5245,N_5593);
and U7980 (N_7980,N_7073,N_6546);
nand U7981 (N_7981,N_7474,N_5060);
or U7982 (N_7982,N_7125,N_6695);
or U7983 (N_7983,N_6510,N_7402);
nand U7984 (N_7984,N_5552,N_5730);
nand U7985 (N_7985,N_6159,N_5528);
and U7986 (N_7986,N_5135,N_5661);
and U7987 (N_7987,N_5349,N_7211);
and U7988 (N_7988,N_7140,N_6096);
or U7989 (N_7989,N_6051,N_5386);
xnor U7990 (N_7990,N_5390,N_6144);
nor U7991 (N_7991,N_5654,N_6542);
nand U7992 (N_7992,N_7014,N_6022);
nor U7993 (N_7993,N_6491,N_7202);
nor U7994 (N_7994,N_5353,N_6167);
and U7995 (N_7995,N_5667,N_6034);
nand U7996 (N_7996,N_6242,N_5600);
nor U7997 (N_7997,N_5304,N_5945);
nand U7998 (N_7998,N_6446,N_5986);
nor U7999 (N_7999,N_6059,N_6282);
nand U8000 (N_8000,N_5935,N_6015);
or U8001 (N_8001,N_6128,N_5583);
nor U8002 (N_8002,N_6111,N_5441);
or U8003 (N_8003,N_5344,N_6470);
xnor U8004 (N_8004,N_5560,N_7279);
nor U8005 (N_8005,N_5844,N_6739);
nand U8006 (N_8006,N_5181,N_5537);
xnor U8007 (N_8007,N_5499,N_6610);
or U8008 (N_8008,N_6254,N_5928);
or U8009 (N_8009,N_6958,N_5900);
nand U8010 (N_8010,N_5049,N_7488);
and U8011 (N_8011,N_5623,N_7272);
or U8012 (N_8012,N_6489,N_5997);
or U8013 (N_8013,N_6526,N_6310);
or U8014 (N_8014,N_5861,N_5831);
nor U8015 (N_8015,N_7024,N_6673);
nand U8016 (N_8016,N_6568,N_7385);
or U8017 (N_8017,N_7033,N_6951);
nor U8018 (N_8018,N_5118,N_5352);
xor U8019 (N_8019,N_7365,N_7035);
xor U8020 (N_8020,N_5290,N_5263);
nor U8021 (N_8021,N_6260,N_5625);
nand U8022 (N_8022,N_6027,N_7138);
nor U8023 (N_8023,N_5100,N_6290);
nor U8024 (N_8024,N_6138,N_7085);
xnor U8025 (N_8025,N_6942,N_5629);
nand U8026 (N_8026,N_7388,N_5119);
nand U8027 (N_8027,N_5350,N_5061);
or U8028 (N_8028,N_5105,N_5087);
and U8029 (N_8029,N_6554,N_6607);
xor U8030 (N_8030,N_5400,N_6061);
xnor U8031 (N_8031,N_6924,N_6164);
or U8032 (N_8032,N_5642,N_7256);
nor U8033 (N_8033,N_5223,N_7170);
xor U8034 (N_8034,N_6730,N_7042);
nand U8035 (N_8035,N_5188,N_6331);
nand U8036 (N_8036,N_6953,N_5260);
xor U8037 (N_8037,N_7400,N_6728);
xnor U8038 (N_8038,N_5189,N_5205);
xor U8039 (N_8039,N_5798,N_6052);
xnor U8040 (N_8040,N_6952,N_5515);
or U8041 (N_8041,N_6720,N_6659);
nor U8042 (N_8042,N_5114,N_5225);
or U8043 (N_8043,N_6565,N_5033);
xor U8044 (N_8044,N_6315,N_6680);
and U8045 (N_8045,N_7206,N_6621);
nor U8046 (N_8046,N_5703,N_5137);
nand U8047 (N_8047,N_6660,N_6050);
and U8048 (N_8048,N_5012,N_7017);
nor U8049 (N_8049,N_5657,N_5837);
or U8050 (N_8050,N_5852,N_5624);
nand U8051 (N_8051,N_5791,N_5901);
or U8052 (N_8052,N_6819,N_5228);
nand U8053 (N_8053,N_5381,N_6973);
nor U8054 (N_8054,N_7442,N_7496);
or U8055 (N_8055,N_6462,N_5167);
and U8056 (N_8056,N_5058,N_6917);
xor U8057 (N_8057,N_6636,N_6748);
xnor U8058 (N_8058,N_6440,N_5702);
and U8059 (N_8059,N_5500,N_5617);
nor U8060 (N_8060,N_6609,N_6455);
and U8061 (N_8061,N_6792,N_5035);
nor U8062 (N_8062,N_6896,N_6875);
or U8063 (N_8063,N_5811,N_6525);
nand U8064 (N_8064,N_7482,N_6216);
nor U8065 (N_8065,N_6665,N_6780);
or U8066 (N_8066,N_6411,N_6433);
or U8067 (N_8067,N_6362,N_5341);
and U8068 (N_8068,N_5463,N_5603);
xnor U8069 (N_8069,N_6221,N_5449);
or U8070 (N_8070,N_5083,N_5253);
xnor U8071 (N_8071,N_6847,N_6724);
nor U8072 (N_8072,N_6691,N_5146);
and U8073 (N_8073,N_5003,N_5202);
and U8074 (N_8074,N_5154,N_6246);
and U8075 (N_8075,N_5072,N_7405);
and U8076 (N_8076,N_6206,N_7436);
xor U8077 (N_8077,N_5453,N_7377);
or U8078 (N_8078,N_5363,N_6312);
and U8079 (N_8079,N_5017,N_7314);
nor U8080 (N_8080,N_5894,N_6426);
and U8081 (N_8081,N_6957,N_5567);
nand U8082 (N_8082,N_6933,N_5970);
nor U8083 (N_8083,N_6271,N_6169);
nor U8084 (N_8084,N_6105,N_7213);
xnor U8085 (N_8085,N_6493,N_5881);
or U8086 (N_8086,N_5098,N_5559);
or U8087 (N_8087,N_6174,N_7259);
xor U8088 (N_8088,N_6231,N_6885);
or U8089 (N_8089,N_6574,N_6849);
nand U8090 (N_8090,N_6897,N_5308);
or U8091 (N_8091,N_5630,N_6963);
nand U8092 (N_8092,N_5655,N_5589);
and U8093 (N_8093,N_5711,N_7452);
nor U8094 (N_8094,N_5196,N_6781);
nor U8095 (N_8095,N_7371,N_5937);
nor U8096 (N_8096,N_5693,N_7316);
and U8097 (N_8097,N_5432,N_6502);
nor U8098 (N_8098,N_5530,N_6432);
nand U8099 (N_8099,N_6805,N_5870);
and U8100 (N_8100,N_6755,N_5555);
nand U8101 (N_8101,N_6262,N_6275);
nand U8102 (N_8102,N_5988,N_6126);
nor U8103 (N_8103,N_6888,N_5803);
xnor U8104 (N_8104,N_6676,N_5216);
nand U8105 (N_8105,N_5361,N_5850);
xor U8106 (N_8106,N_5371,N_7368);
and U8107 (N_8107,N_6294,N_5823);
xnor U8108 (N_8108,N_5252,N_5906);
nand U8109 (N_8109,N_7463,N_6707);
nand U8110 (N_8110,N_5018,N_6514);
or U8111 (N_8111,N_5054,N_6038);
nor U8112 (N_8112,N_6195,N_5752);
nand U8113 (N_8113,N_5773,N_5827);
nor U8114 (N_8114,N_5200,N_6263);
or U8115 (N_8115,N_7217,N_5849);
and U8116 (N_8116,N_6396,N_5406);
or U8117 (N_8117,N_7126,N_6516);
and U8118 (N_8118,N_5879,N_6176);
xor U8119 (N_8119,N_5632,N_5546);
nor U8120 (N_8120,N_5726,N_6628);
nor U8121 (N_8121,N_6276,N_6129);
or U8122 (N_8122,N_7241,N_5953);
and U8123 (N_8123,N_6348,N_6011);
or U8124 (N_8124,N_5480,N_6881);
and U8125 (N_8125,N_5203,N_5282);
nand U8126 (N_8126,N_5321,N_7459);
and U8127 (N_8127,N_5996,N_6305);
and U8128 (N_8128,N_6966,N_5250);
xnor U8129 (N_8129,N_5145,N_7048);
nor U8130 (N_8130,N_5269,N_5794);
xnor U8131 (N_8131,N_7439,N_6536);
and U8132 (N_8132,N_5993,N_5143);
and U8133 (N_8133,N_7019,N_5770);
and U8134 (N_8134,N_6977,N_6400);
or U8135 (N_8135,N_5768,N_6763);
nor U8136 (N_8136,N_5394,N_7093);
nand U8137 (N_8137,N_6851,N_6392);
nor U8138 (N_8138,N_7284,N_5032);
or U8139 (N_8139,N_5506,N_7031);
and U8140 (N_8140,N_6908,N_6049);
or U8141 (N_8141,N_7069,N_7327);
nand U8142 (N_8142,N_5377,N_7437);
or U8143 (N_8143,N_6405,N_7473);
nor U8144 (N_8144,N_7423,N_6008);
and U8145 (N_8145,N_7278,N_5683);
or U8146 (N_8146,N_7015,N_5696);
and U8147 (N_8147,N_5370,N_5731);
xor U8148 (N_8148,N_5397,N_5177);
nand U8149 (N_8149,N_6907,N_6648);
xnor U8150 (N_8150,N_6641,N_6829);
nor U8151 (N_8151,N_5473,N_6996);
or U8152 (N_8152,N_5833,N_7443);
xnor U8153 (N_8153,N_6480,N_6871);
nor U8154 (N_8154,N_5079,N_7186);
and U8155 (N_8155,N_5695,N_6381);
xor U8156 (N_8156,N_7374,N_6675);
nand U8157 (N_8157,N_6451,N_5929);
xor U8158 (N_8158,N_5820,N_7415);
nand U8159 (N_8159,N_6304,N_5287);
nor U8160 (N_8160,N_5268,N_5825);
xor U8161 (N_8161,N_6836,N_5712);
or U8162 (N_8162,N_5358,N_6010);
nor U8163 (N_8163,N_6767,N_6637);
nor U8164 (N_8164,N_6026,N_6747);
or U8165 (N_8165,N_7216,N_6865);
nand U8166 (N_8166,N_6021,N_5922);
nor U8167 (N_8167,N_7413,N_6814);
nand U8168 (N_8168,N_5485,N_5343);
xor U8169 (N_8169,N_5949,N_7339);
or U8170 (N_8170,N_5897,N_5331);
xnor U8171 (N_8171,N_7282,N_6709);
nor U8172 (N_8172,N_6178,N_5761);
xor U8173 (N_8173,N_7333,N_7445);
xor U8174 (N_8174,N_6959,N_7354);
nand U8175 (N_8175,N_7416,N_5750);
nand U8176 (N_8176,N_7187,N_5163);
or U8177 (N_8177,N_6539,N_7018);
or U8178 (N_8178,N_6645,N_5887);
nand U8179 (N_8179,N_6980,N_7045);
and U8180 (N_8180,N_6723,N_6618);
nand U8181 (N_8181,N_5244,N_6240);
nor U8182 (N_8182,N_6595,N_5664);
nand U8183 (N_8183,N_6173,N_7153);
and U8184 (N_8184,N_7004,N_6928);
xnor U8185 (N_8185,N_5014,N_7037);
and U8186 (N_8186,N_5468,N_6839);
nor U8187 (N_8187,N_6627,N_6202);
xor U8188 (N_8188,N_6846,N_5127);
nor U8189 (N_8189,N_7262,N_6861);
xor U8190 (N_8190,N_7199,N_5278);
or U8191 (N_8191,N_6496,N_6226);
and U8192 (N_8192,N_6158,N_6340);
xnor U8193 (N_8193,N_6850,N_6578);
and U8194 (N_8194,N_5633,N_6684);
and U8195 (N_8195,N_5317,N_6092);
and U8196 (N_8196,N_6530,N_5254);
nand U8197 (N_8197,N_6656,N_5435);
nand U8198 (N_8198,N_5484,N_5975);
and U8199 (N_8199,N_6190,N_6112);
nand U8200 (N_8200,N_7255,N_6583);
xor U8201 (N_8201,N_6670,N_6244);
or U8202 (N_8202,N_7367,N_7013);
or U8203 (N_8203,N_7012,N_6915);
nand U8204 (N_8204,N_5585,N_5346);
or U8205 (N_8205,N_7406,N_5502);
xor U8206 (N_8206,N_5273,N_6474);
or U8207 (N_8207,N_5598,N_6775);
xnor U8208 (N_8208,N_6797,N_7209);
and U8209 (N_8209,N_6505,N_5389);
nand U8210 (N_8210,N_5374,N_6853);
or U8211 (N_8211,N_6991,N_5989);
xnor U8212 (N_8212,N_6960,N_6043);
or U8213 (N_8213,N_6429,N_7065);
and U8214 (N_8214,N_5327,N_5857);
nand U8215 (N_8215,N_5483,N_5514);
xor U8216 (N_8216,N_6920,N_6420);
nor U8217 (N_8217,N_7054,N_6044);
and U8218 (N_8218,N_6886,N_6399);
nor U8219 (N_8219,N_5393,N_6095);
xnor U8220 (N_8220,N_5486,N_6257);
and U8221 (N_8221,N_5090,N_7070);
or U8222 (N_8222,N_6380,N_6268);
and U8223 (N_8223,N_6247,N_5044);
and U8224 (N_8224,N_6088,N_6093);
or U8225 (N_8225,N_6711,N_7312);
nor U8226 (N_8226,N_5246,N_6541);
nor U8227 (N_8227,N_6697,N_6342);
nand U8228 (N_8228,N_6880,N_6918);
xnor U8229 (N_8229,N_5265,N_5016);
and U8230 (N_8230,N_5448,N_5133);
nand U8231 (N_8231,N_5878,N_7183);
nor U8232 (N_8232,N_7319,N_5088);
and U8233 (N_8233,N_5218,N_7051);
nand U8234 (N_8234,N_5643,N_5160);
or U8235 (N_8235,N_5843,N_5659);
nor U8236 (N_8236,N_5064,N_5466);
xor U8237 (N_8237,N_5309,N_6727);
nand U8238 (N_8238,N_7355,N_7123);
nand U8239 (N_8239,N_7200,N_6108);
or U8240 (N_8240,N_7076,N_5094);
xor U8241 (N_8241,N_6874,N_5295);
or U8242 (N_8242,N_6087,N_6409);
and U8243 (N_8243,N_7100,N_5682);
nor U8244 (N_8244,N_6504,N_7432);
and U8245 (N_8245,N_5052,N_7260);
or U8246 (N_8246,N_6418,N_7277);
or U8247 (N_8247,N_6882,N_6988);
xnor U8248 (N_8248,N_7251,N_7410);
xnor U8249 (N_8249,N_5130,N_6366);
and U8250 (N_8250,N_7323,N_5379);
and U8251 (N_8251,N_5685,N_6838);
xor U8252 (N_8252,N_7395,N_5226);
nand U8253 (N_8253,N_6700,N_5733);
nor U8254 (N_8254,N_5776,N_5150);
nor U8255 (N_8255,N_6316,N_6738);
xor U8256 (N_8256,N_6236,N_6981);
or U8257 (N_8257,N_6802,N_6559);
xnor U8258 (N_8258,N_6218,N_7270);
and U8259 (N_8259,N_5972,N_7009);
or U8260 (N_8260,N_5301,N_6363);
and U8261 (N_8261,N_7077,N_5588);
or U8262 (N_8262,N_5479,N_5605);
and U8263 (N_8263,N_6778,N_5576);
xnor U8264 (N_8264,N_6020,N_7326);
nand U8265 (N_8265,N_6856,N_5208);
and U8266 (N_8266,N_5174,N_7384);
nor U8267 (N_8267,N_6253,N_5220);
or U8268 (N_8268,N_6181,N_5817);
xor U8269 (N_8269,N_6735,N_5408);
and U8270 (N_8270,N_5645,N_6795);
nor U8271 (N_8271,N_5512,N_6679);
nand U8272 (N_8272,N_6130,N_6822);
or U8273 (N_8273,N_5525,N_5965);
and U8274 (N_8274,N_6481,N_6867);
and U8275 (N_8275,N_6513,N_6171);
xnor U8276 (N_8276,N_7253,N_6408);
nor U8277 (N_8277,N_6599,N_6769);
xor U8278 (N_8278,N_6904,N_6860);
xor U8279 (N_8279,N_6826,N_6905);
or U8280 (N_8280,N_6039,N_5124);
nor U8281 (N_8281,N_6343,N_5884);
or U8282 (N_8282,N_5960,N_5719);
nand U8283 (N_8283,N_7091,N_6419);
nor U8284 (N_8284,N_5292,N_5077);
and U8285 (N_8285,N_7440,N_7151);
nand U8286 (N_8286,N_5209,N_6101);
xor U8287 (N_8287,N_5333,N_6252);
nor U8288 (N_8288,N_6062,N_6619);
xor U8289 (N_8289,N_6177,N_5754);
nor U8290 (N_8290,N_6998,N_7158);
xnor U8291 (N_8291,N_5136,N_5262);
nand U8292 (N_8292,N_5575,N_6355);
xnor U8293 (N_8293,N_5142,N_6289);
and U8294 (N_8294,N_7309,N_6894);
nor U8295 (N_8295,N_7114,N_6354);
and U8296 (N_8296,N_6213,N_6083);
or U8297 (N_8297,N_7396,N_6681);
or U8298 (N_8298,N_6259,N_6624);
or U8299 (N_8299,N_7027,N_6511);
and U8300 (N_8300,N_5772,N_6110);
and U8301 (N_8301,N_5045,N_5156);
and U8302 (N_8302,N_6750,N_6328);
and U8303 (N_8303,N_7398,N_7470);
or U8304 (N_8304,N_7124,N_5159);
nand U8305 (N_8305,N_6047,N_5531);
or U8306 (N_8306,N_5626,N_6248);
nor U8307 (N_8307,N_6133,N_5241);
and U8308 (N_8308,N_6855,N_6663);
xor U8309 (N_8309,N_6107,N_5539);
nand U8310 (N_8310,N_6229,N_5385);
nor U8311 (N_8311,N_6017,N_6333);
and U8312 (N_8312,N_6594,N_7491);
or U8313 (N_8313,N_6337,N_7362);
and U8314 (N_8314,N_5439,N_5917);
nor U8315 (N_8315,N_6742,N_6776);
nand U8316 (N_8316,N_6180,N_5834);
nor U8317 (N_8317,N_7055,N_7184);
nand U8318 (N_8318,N_7375,N_5679);
or U8319 (N_8319,N_5281,N_5815);
or U8320 (N_8320,N_5855,N_7011);
nor U8321 (N_8321,N_6031,N_7072);
or U8322 (N_8322,N_6103,N_6759);
or U8323 (N_8323,N_5984,N_6200);
nand U8324 (N_8324,N_5259,N_5802);
nor U8325 (N_8325,N_5869,N_7376);
or U8326 (N_8326,N_6194,N_5224);
or U8327 (N_8327,N_5222,N_6500);
nand U8328 (N_8328,N_7417,N_5270);
and U8329 (N_8329,N_5735,N_6912);
xnor U8330 (N_8330,N_5104,N_6548);
and U8331 (N_8331,N_5428,N_5565);
xnor U8332 (N_8332,N_5134,N_6870);
and U8333 (N_8333,N_7249,N_5211);
xor U8334 (N_8334,N_6858,N_7171);
nor U8335 (N_8335,N_5652,N_7478);
or U8336 (N_8336,N_5689,N_7235);
and U8337 (N_8337,N_6823,N_6225);
and U8338 (N_8338,N_6820,N_6854);
or U8339 (N_8339,N_6662,N_6063);
or U8340 (N_8340,N_5721,N_6667);
nor U8341 (N_8341,N_6323,N_7485);
or U8342 (N_8342,N_6273,N_5838);
nor U8343 (N_8343,N_6372,N_7245);
xor U8344 (N_8344,N_7205,N_5740);
nor U8345 (N_8345,N_7250,N_5671);
xnor U8346 (N_8346,N_5517,N_6217);
xnor U8347 (N_8347,N_5821,N_6132);
xor U8348 (N_8348,N_5662,N_5443);
or U8349 (N_8349,N_5409,N_7088);
or U8350 (N_8350,N_6163,N_5451);
or U8351 (N_8351,N_6577,N_6067);
or U8352 (N_8352,N_7198,N_7137);
and U8353 (N_8353,N_5713,N_5243);
nor U8354 (N_8354,N_5332,N_5709);
nor U8355 (N_8355,N_6002,N_5718);
and U8356 (N_8356,N_7120,N_6029);
or U8357 (N_8357,N_5180,N_6978);
nand U8358 (N_8358,N_5430,N_6804);
xor U8359 (N_8359,N_6238,N_5732);
nor U8360 (N_8360,N_6677,N_5545);
or U8361 (N_8361,N_7182,N_5050);
or U8362 (N_8362,N_7328,N_6591);
nor U8363 (N_8363,N_6123,N_6785);
and U8364 (N_8364,N_6192,N_6227);
nand U8365 (N_8365,N_7110,N_5000);
nor U8366 (N_8366,N_7084,N_6833);
nor U8367 (N_8367,N_6726,N_7175);
and U8368 (N_8368,N_5026,N_7361);
xnor U8369 (N_8369,N_5069,N_5053);
and U8370 (N_8370,N_5470,N_5591);
nand U8371 (N_8371,N_5516,N_6948);
nor U8372 (N_8372,N_5788,N_5129);
nor U8373 (N_8373,N_7068,N_7381);
nor U8374 (N_8374,N_6427,N_7156);
and U8375 (N_8375,N_5990,N_5785);
or U8376 (N_8376,N_6465,N_5437);
nand U8377 (N_8377,N_6999,N_7421);
nand U8378 (N_8378,N_5011,N_7081);
and U8379 (N_8379,N_5126,N_5300);
xor U8380 (N_8380,N_5627,N_5191);
xor U8381 (N_8381,N_6773,N_7082);
and U8382 (N_8382,N_7458,N_6376);
nand U8383 (N_8383,N_6713,N_7119);
xnor U8384 (N_8384,N_6368,N_6705);
nor U8385 (N_8385,N_5004,N_7397);
and U8386 (N_8386,N_5022,N_7050);
and U8387 (N_8387,N_5025,N_6224);
nor U8388 (N_8388,N_7052,N_5757);
xor U8389 (N_8389,N_5492,N_7061);
and U8390 (N_8390,N_6950,N_5921);
nor U8391 (N_8391,N_7356,N_6459);
or U8392 (N_8392,N_6678,N_6543);
and U8393 (N_8393,N_6616,N_6280);
or U8394 (N_8394,N_7364,N_6406);
nand U8395 (N_8395,N_6840,N_7313);
nor U8396 (N_8396,N_5055,N_6832);
nor U8397 (N_8397,N_5863,N_5401);
nand U8398 (N_8398,N_5538,N_7441);
and U8399 (N_8399,N_5968,N_5434);
and U8400 (N_8400,N_5503,N_7435);
xnor U8401 (N_8401,N_5416,N_6387);
nand U8402 (N_8402,N_6250,N_5587);
xor U8403 (N_8403,N_5318,N_6403);
and U8404 (N_8404,N_5081,N_6307);
nor U8405 (N_8405,N_5138,N_6004);
or U8406 (N_8406,N_6930,N_6611);
nand U8407 (N_8407,N_7480,N_5251);
nor U8408 (N_8408,N_6109,N_5232);
nor U8409 (N_8409,N_7148,N_5102);
and U8410 (N_8410,N_6955,N_6119);
and U8411 (N_8411,N_6371,N_6085);
nor U8412 (N_8412,N_6410,N_6161);
xnor U8413 (N_8413,N_6314,N_7185);
nand U8414 (N_8414,N_6142,N_6498);
or U8415 (N_8415,N_6757,N_5319);
nor U8416 (N_8416,N_7261,N_5807);
nand U8417 (N_8417,N_5082,N_5204);
and U8418 (N_8418,N_6916,N_7060);
and U8419 (N_8419,N_7101,N_7446);
nand U8420 (N_8420,N_6235,N_7246);
xnor U8421 (N_8421,N_6799,N_5037);
nand U8422 (N_8422,N_7144,N_7083);
xor U8423 (N_8423,N_7218,N_6784);
and U8424 (N_8424,N_5534,N_5373);
xor U8425 (N_8425,N_5296,N_5148);
and U8426 (N_8426,N_5231,N_5383);
nand U8427 (N_8427,N_5117,N_6683);
or U8428 (N_8428,N_7203,N_6827);
or U8429 (N_8429,N_5306,N_7320);
and U8430 (N_8430,N_5274,N_7341);
and U8431 (N_8431,N_5829,N_7464);
nand U8432 (N_8432,N_7307,N_7243);
nand U8433 (N_8433,N_5618,N_7025);
and U8434 (N_8434,N_5675,N_5242);
nor U8435 (N_8435,N_6189,N_5967);
nand U8436 (N_8436,N_6806,N_5796);
xnor U8437 (N_8437,N_6818,N_7427);
nand U8438 (N_8438,N_6623,N_5867);
and U8439 (N_8439,N_6501,N_6949);
or U8440 (N_8440,N_5490,N_5084);
xnor U8441 (N_8441,N_6241,N_7275);
nor U8442 (N_8442,N_7020,N_6421);
and U8443 (N_8443,N_6592,N_5407);
and U8444 (N_8444,N_7344,N_6879);
xor U8445 (N_8445,N_7286,N_6931);
or U8446 (N_8446,N_5533,N_5369);
nand U8447 (N_8447,N_5063,N_5594);
or U8448 (N_8448,N_5795,N_5616);
nor U8449 (N_8449,N_5433,N_5818);
nor U8450 (N_8450,N_6716,N_6791);
xnor U8451 (N_8451,N_6024,N_6299);
xor U8452 (N_8452,N_6606,N_7047);
xnor U8453 (N_8453,N_6801,N_6993);
xnor U8454 (N_8454,N_6303,N_5956);
or U8455 (N_8455,N_5961,N_6940);
nor U8456 (N_8456,N_6237,N_5197);
nand U8457 (N_8457,N_5903,N_7214);
nor U8458 (N_8458,N_6139,N_6632);
xor U8459 (N_8459,N_6655,N_7484);
nor U8460 (N_8460,N_7162,N_6212);
nor U8461 (N_8461,N_7139,N_6048);
nor U8462 (N_8462,N_6550,N_5074);
and U8463 (N_8463,N_7267,N_6798);
or U8464 (N_8464,N_5816,N_6106);
xnor U8465 (N_8465,N_6598,N_7281);
xnor U8466 (N_8466,N_7040,N_7181);
nor U8467 (N_8467,N_6891,N_6967);
or U8468 (N_8468,N_7132,N_6864);
xor U8469 (N_8469,N_6413,N_5550);
nand U8470 (N_8470,N_6557,N_6664);
xnor U8471 (N_8471,N_7420,N_5285);
xor U8472 (N_8472,N_6151,N_5283);
or U8473 (N_8473,N_6786,N_5579);
xnor U8474 (N_8474,N_7448,N_6590);
nor U8475 (N_8475,N_6428,N_6135);
nand U8476 (N_8476,N_5985,N_6291);
and U8477 (N_8477,N_6184,N_5368);
nor U8478 (N_8478,N_5926,N_5898);
nand U8479 (N_8479,N_5162,N_6321);
and U8480 (N_8480,N_6682,N_7486);
or U8481 (N_8481,N_7300,N_5789);
or U8482 (N_8482,N_7254,N_6652);
and U8483 (N_8483,N_7121,N_5024);
or U8484 (N_8484,N_6077,N_6586);
and U8485 (N_8485,N_7133,N_6311);
nand U8486 (N_8486,N_6671,N_6689);
nor U8487 (N_8487,N_7169,N_5475);
nor U8488 (N_8488,N_5650,N_5212);
nor U8489 (N_8489,N_6394,N_6813);
nand U8490 (N_8490,N_5890,N_5413);
nand U8491 (N_8491,N_5297,N_5235);
nor U8492 (N_8492,N_6416,N_7128);
or U8493 (N_8493,N_7079,N_7028);
and U8494 (N_8494,N_7412,N_5910);
or U8495 (N_8495,N_6168,N_5668);
and U8496 (N_8496,N_5015,N_6556);
or U8497 (N_8497,N_5426,N_5697);
xnor U8498 (N_8498,N_7127,N_5766);
or U8499 (N_8499,N_7378,N_6258);
nor U8500 (N_8500,N_5415,N_5418);
xor U8501 (N_8501,N_5164,N_5720);
xnor U8502 (N_8502,N_7298,N_5028);
or U8503 (N_8503,N_6078,N_5701);
or U8504 (N_8504,N_5455,N_6390);
or U8505 (N_8505,N_5029,N_6270);
xor U8506 (N_8506,N_5866,N_5809);
nand U8507 (N_8507,N_5543,N_7107);
nand U8508 (N_8508,N_7001,N_5864);
and U8509 (N_8509,N_6644,N_5171);
xnor U8510 (N_8510,N_5364,N_6243);
nand U8511 (N_8511,N_6941,N_6359);
or U8512 (N_8512,N_6760,N_7022);
or U8513 (N_8513,N_7481,N_6436);
nand U8514 (N_8514,N_6000,N_5601);
or U8515 (N_8515,N_6013,N_5068);
nand U8516 (N_8516,N_5548,N_5738);
or U8517 (N_8517,N_6033,N_6703);
nor U8518 (N_8518,N_5239,N_5638);
or U8519 (N_8519,N_5658,N_5384);
xnor U8520 (N_8520,N_6841,N_7357);
and U8521 (N_8521,N_6222,N_6154);
nand U8522 (N_8522,N_6338,N_7492);
nor U8523 (N_8523,N_5348,N_6734);
and U8524 (N_8524,N_6789,N_5813);
nand U8525 (N_8525,N_5144,N_5606);
nor U8526 (N_8526,N_7238,N_6191);
nand U8527 (N_8527,N_6369,N_5727);
and U8528 (N_8528,N_6175,N_7244);
or U8529 (N_8529,N_5936,N_6553);
or U8530 (N_8530,N_5372,N_5279);
and U8531 (N_8531,N_7094,N_5763);
xor U8532 (N_8532,N_5556,N_5992);
nor U8533 (N_8533,N_6058,N_6397);
or U8534 (N_8534,N_6162,N_7192);
nand U8535 (N_8535,N_5639,N_6464);
nor U8536 (N_8536,N_6434,N_5613);
and U8537 (N_8537,N_6944,N_6347);
nor U8538 (N_8538,N_6365,N_6710);
xnor U8539 (N_8539,N_7257,N_5185);
xnor U8540 (N_8540,N_6204,N_6573);
xor U8541 (N_8541,N_6600,N_7294);
and U8542 (N_8542,N_7266,N_5036);
nor U8543 (N_8543,N_5636,N_7352);
or U8544 (N_8544,N_6030,N_7167);
nor U8545 (N_8545,N_6686,N_5073);
or U8546 (N_8546,N_5578,N_6145);
and U8547 (N_8547,N_5152,N_7039);
and U8548 (N_8548,N_7227,N_7043);
and U8549 (N_8549,N_6834,N_6824);
nand U8550 (N_8550,N_6094,N_6155);
or U8551 (N_8551,N_7221,N_7215);
nand U8552 (N_8552,N_5602,N_6572);
or U8553 (N_8553,N_6661,N_6185);
and U8554 (N_8554,N_5705,N_5847);
xor U8555 (N_8555,N_6706,N_6385);
nor U8556 (N_8556,N_6626,N_6702);
nand U8557 (N_8557,N_6284,N_6545);
nor U8558 (N_8558,N_6287,N_6452);
or U8559 (N_8559,N_6345,N_7346);
xor U8560 (N_8560,N_7324,N_5963);
and U8561 (N_8561,N_5195,N_5013);
and U8562 (N_8562,N_5405,N_7049);
and U8563 (N_8563,N_5737,N_5008);
and U8564 (N_8564,N_6986,N_6035);
nand U8565 (N_8565,N_6582,N_5001);
nand U8566 (N_8566,N_5266,N_6544);
xnor U8567 (N_8567,N_6012,N_5886);
nor U8568 (N_8568,N_6295,N_5305);
or U8569 (N_8569,N_5876,N_5496);
or U8570 (N_8570,N_6935,N_5519);
or U8571 (N_8571,N_5925,N_6461);
nor U8572 (N_8572,N_6353,N_5467);
nand U8573 (N_8573,N_6069,N_5690);
and U8574 (N_8574,N_5790,N_5621);
nand U8575 (N_8575,N_7495,N_5536);
xor U8576 (N_8576,N_7102,N_5669);
nor U8577 (N_8577,N_5175,N_6975);
xor U8578 (N_8578,N_5048,N_6551);
nor U8579 (N_8579,N_7016,N_6170);
or U8580 (N_8580,N_6125,N_7092);
and U8581 (N_8581,N_5756,N_5042);
xnor U8582 (N_8582,N_6507,N_6070);
xor U8583 (N_8583,N_6743,N_5611);
nor U8584 (N_8584,N_7086,N_7444);
nor U8585 (N_8585,N_6302,N_5365);
xor U8586 (N_8586,N_5109,N_6382);
and U8587 (N_8587,N_6537,N_5474);
or U8588 (N_8588,N_5080,N_5694);
nor U8589 (N_8589,N_7066,N_5692);
or U8590 (N_8590,N_5767,N_6934);
xor U8591 (N_8591,N_7394,N_5095);
nor U8592 (N_8592,N_7113,N_6486);
xor U8593 (N_8593,N_5549,N_7224);
or U8594 (N_8594,N_6549,N_5051);
xor U8595 (N_8595,N_6003,N_6749);
or U8596 (N_8596,N_6566,N_5027);
and U8597 (N_8597,N_7189,N_6965);
xor U8598 (N_8598,N_5634,N_5644);
or U8599 (N_8599,N_5714,N_6852);
xor U8600 (N_8600,N_5896,N_5914);
and U8601 (N_8601,N_7325,N_5340);
nor U8602 (N_8602,N_6084,N_5122);
nand U8603 (N_8603,N_7343,N_7449);
nand U8604 (N_8604,N_5314,N_6028);
or U8605 (N_8605,N_6715,N_5599);
and U8606 (N_8606,N_6166,N_5974);
and U8607 (N_8607,N_6925,N_5793);
nor U8608 (N_8608,N_5808,N_6269);
nor U8609 (N_8609,N_6994,N_6562);
and U8610 (N_8610,N_5676,N_6984);
nand U8611 (N_8611,N_6468,N_7455);
and U8612 (N_8612,N_7331,N_6523);
nand U8613 (N_8613,N_7196,N_7497);
or U8614 (N_8614,N_6292,N_5066);
and U8615 (N_8615,N_5959,N_5913);
and U8616 (N_8616,N_6391,N_5874);
or U8617 (N_8617,N_5085,N_6007);
nand U8618 (N_8618,N_6071,N_6995);
nand U8619 (N_8619,N_5238,N_7248);
or U8620 (N_8620,N_6398,N_6286);
nor U8621 (N_8621,N_6848,N_6300);
and U8622 (N_8622,N_5943,N_5819);
nor U8623 (N_8623,N_5391,N_5806);
nand U8624 (N_8624,N_5322,N_6074);
nor U8625 (N_8625,N_5958,N_5417);
nor U8626 (N_8626,N_5527,N_7493);
nand U8627 (N_8627,N_6638,N_6160);
nand U8628 (N_8628,N_5577,N_6442);
nor U8629 (N_8629,N_5456,N_6114);
xor U8630 (N_8630,N_6968,N_5962);
nor U8631 (N_8631,N_5176,N_5482);
nor U8632 (N_8632,N_6198,N_7118);
and U8633 (N_8633,N_6712,N_7006);
or U8634 (N_8634,N_6157,N_5460);
or U8635 (N_8635,N_7041,N_5665);
xor U8636 (N_8636,N_5951,N_6812);
nor U8637 (N_8637,N_6332,N_5307);
nand U8638 (N_8638,N_5860,N_7471);
and U8639 (N_8639,N_6887,N_7490);
and U8640 (N_8640,N_6863,N_6389);
or U8641 (N_8641,N_6762,N_6929);
nor U8642 (N_8642,N_6037,N_6073);
xor U8643 (N_8643,N_6463,N_5574);
and U8644 (N_8644,N_6375,N_6239);
and U8645 (N_8645,N_5631,N_5236);
nand U8646 (N_8646,N_6733,N_7450);
or U8647 (N_8647,N_7499,N_5915);
nor U8648 (N_8648,N_5347,N_5065);
and U8649 (N_8649,N_5710,N_7276);
and U8650 (N_8650,N_6868,N_7337);
or U8651 (N_8651,N_7387,N_5120);
nand U8652 (N_8652,N_6272,N_6972);
nor U8653 (N_8653,N_7105,N_7349);
nand U8654 (N_8654,N_6055,N_5828);
and U8655 (N_8655,N_5213,N_5256);
nor U8656 (N_8656,N_6788,N_5998);
nor U8657 (N_8657,N_6412,N_6279);
nor U8658 (N_8658,N_6384,N_7292);
nand U8659 (N_8659,N_5804,N_6892);
xor U8660 (N_8660,N_6974,N_6068);
nor U8661 (N_8661,N_6329,N_7030);
nor U8662 (N_8662,N_5841,N_5092);
xor U8663 (N_8663,N_6503,N_6901);
nand U8664 (N_8664,N_6936,N_7219);
nand U8665 (N_8665,N_6650,N_5075);
or U8666 (N_8666,N_5132,N_6223);
and U8667 (N_8667,N_5395,N_5729);
nand U8668 (N_8668,N_7111,N_7264);
xnor U8669 (N_8669,N_7036,N_5842);
nand U8670 (N_8670,N_6779,N_6612);
xnor U8671 (N_8671,N_5182,N_5822);
nand U8672 (N_8672,N_6532,N_6527);
or U8673 (N_8673,N_7190,N_5982);
xor U8674 (N_8674,N_5489,N_7005);
or U8675 (N_8675,N_6351,N_7010);
or U8676 (N_8676,N_6777,N_6919);
or U8677 (N_8677,N_6803,N_6449);
and U8678 (N_8678,N_5427,N_6014);
or U8679 (N_8679,N_5983,N_5030);
and U8680 (N_8680,N_6404,N_7177);
xor U8681 (N_8681,N_6939,N_5717);
or U8682 (N_8682,N_6344,N_5532);
nor U8683 (N_8683,N_7469,N_7021);
nor U8684 (N_8684,N_6722,N_5337);
nand U8685 (N_8685,N_7122,N_5271);
xor U8686 (N_8686,N_5411,N_6205);
or U8687 (N_8687,N_7155,N_5592);
nand U8688 (N_8688,N_6306,N_7222);
and U8689 (N_8689,N_6490,N_5610);
nand U8690 (N_8690,N_5168,N_7317);
nor U8691 (N_8691,N_5635,N_6893);
nand U8692 (N_8692,N_7166,N_6266);
nand U8693 (N_8693,N_6009,N_5067);
xnor U8694 (N_8694,N_7180,N_5356);
or U8695 (N_8695,N_5217,N_6878);
nand U8696 (N_8696,N_5020,N_5723);
nor U8697 (N_8697,N_5324,N_7087);
nor U8698 (N_8698,N_6116,N_6989);
and U8699 (N_8699,N_6732,N_5402);
or U8700 (N_8700,N_5835,N_7032);
nor U8701 (N_8701,N_5751,N_7466);
and U8702 (N_8702,N_5748,N_6117);
nor U8703 (N_8703,N_7424,N_7231);
xnor U8704 (N_8704,N_5410,N_6588);
nor U8705 (N_8705,N_5392,N_5749);
xnor U8706 (N_8706,N_5187,N_7176);
or U8707 (N_8707,N_6876,N_6417);
xnor U8708 (N_8708,N_6124,N_6251);
xnor U8709 (N_8709,N_5619,N_6970);
nor U8710 (N_8710,N_6937,N_5540);
or U8711 (N_8711,N_5399,N_7135);
nand U8712 (N_8712,N_7007,N_5920);
nand U8713 (N_8713,N_6552,N_6796);
and U8714 (N_8714,N_6831,N_5880);
or U8715 (N_8715,N_5562,N_6309);
xnor U8716 (N_8716,N_6423,N_6866);
or U8717 (N_8717,N_5969,N_5526);
or U8718 (N_8718,N_7201,N_5753);
xor U8719 (N_8719,N_6571,N_6220);
nor U8720 (N_8720,N_5076,N_6424);
and U8721 (N_8721,N_6137,N_5952);
nor U8722 (N_8722,N_5924,N_5944);
or U8723 (N_8723,N_7350,N_7157);
and U8724 (N_8724,N_6326,N_5955);
nand U8725 (N_8725,N_7287,N_5942);
xor U8726 (N_8726,N_6140,N_7408);
xor U8727 (N_8727,N_5580,N_7369);
xor U8728 (N_8728,N_7057,N_6374);
or U8729 (N_8729,N_5741,N_5403);
nand U8730 (N_8730,N_5501,N_5728);
and U8731 (N_8731,N_7269,N_6547);
nor U8732 (N_8732,N_6900,N_6560);
xor U8733 (N_8733,N_7204,N_6809);
xor U8734 (N_8734,N_5173,N_5315);
nand U8735 (N_8735,N_6297,N_6460);
nor U8736 (N_8736,N_5620,N_7179);
or U8737 (N_8737,N_6699,N_6569);
and U8738 (N_8738,N_5039,N_6736);
or U8739 (N_8739,N_6745,N_7141);
nor U8740 (N_8740,N_5586,N_5311);
and U8741 (N_8741,N_6538,N_7071);
or U8742 (N_8742,N_7232,N_7178);
nor U8743 (N_8743,N_6883,N_6810);
nand U8744 (N_8744,N_7318,N_7002);
nand U8745 (N_8745,N_6622,N_6487);
xor U8746 (N_8746,N_7393,N_5288);
nor U8747 (N_8747,N_6782,N_6150);
or U8748 (N_8748,N_6379,N_7099);
and U8749 (N_8749,N_7401,N_7363);
nand U8750 (N_8750,N_5609,N_5768);
nor U8751 (N_8751,N_6502,N_6463);
nor U8752 (N_8752,N_6728,N_5000);
or U8753 (N_8753,N_6095,N_6980);
and U8754 (N_8754,N_7408,N_6284);
nand U8755 (N_8755,N_5415,N_6137);
nor U8756 (N_8756,N_6482,N_6476);
xor U8757 (N_8757,N_5597,N_7355);
nor U8758 (N_8758,N_6306,N_5433);
nand U8759 (N_8759,N_7292,N_6126);
nand U8760 (N_8760,N_6749,N_6089);
and U8761 (N_8761,N_5301,N_5876);
nor U8762 (N_8762,N_6680,N_5202);
nor U8763 (N_8763,N_6392,N_5822);
nand U8764 (N_8764,N_6422,N_5693);
or U8765 (N_8765,N_7093,N_5010);
nor U8766 (N_8766,N_6755,N_6193);
xnor U8767 (N_8767,N_6587,N_5168);
nor U8768 (N_8768,N_6241,N_6079);
nand U8769 (N_8769,N_5231,N_5861);
and U8770 (N_8770,N_6888,N_6322);
or U8771 (N_8771,N_6319,N_6757);
or U8772 (N_8772,N_7225,N_5263);
nor U8773 (N_8773,N_6668,N_5901);
or U8774 (N_8774,N_5320,N_5215);
nor U8775 (N_8775,N_5743,N_7445);
xor U8776 (N_8776,N_6353,N_7112);
nand U8777 (N_8777,N_7005,N_6058);
and U8778 (N_8778,N_6453,N_6375);
and U8779 (N_8779,N_5512,N_5611);
nand U8780 (N_8780,N_5044,N_5349);
xor U8781 (N_8781,N_5044,N_6309);
nand U8782 (N_8782,N_7113,N_6885);
and U8783 (N_8783,N_6835,N_7190);
xnor U8784 (N_8784,N_7288,N_5433);
and U8785 (N_8785,N_6195,N_5537);
or U8786 (N_8786,N_5516,N_7411);
or U8787 (N_8787,N_5739,N_6944);
or U8788 (N_8788,N_6923,N_6251);
nand U8789 (N_8789,N_5383,N_7276);
or U8790 (N_8790,N_5152,N_6723);
xor U8791 (N_8791,N_7016,N_5626);
or U8792 (N_8792,N_7352,N_6199);
or U8793 (N_8793,N_5209,N_6691);
xor U8794 (N_8794,N_7035,N_7180);
nand U8795 (N_8795,N_6812,N_6427);
xnor U8796 (N_8796,N_6674,N_6080);
or U8797 (N_8797,N_6274,N_5217);
nand U8798 (N_8798,N_6154,N_7100);
and U8799 (N_8799,N_6108,N_7315);
nor U8800 (N_8800,N_5147,N_5217);
and U8801 (N_8801,N_5934,N_5716);
xor U8802 (N_8802,N_7347,N_5292);
nand U8803 (N_8803,N_5782,N_6392);
xor U8804 (N_8804,N_6187,N_5188);
xor U8805 (N_8805,N_5341,N_5250);
nor U8806 (N_8806,N_5165,N_6509);
or U8807 (N_8807,N_6419,N_5442);
nand U8808 (N_8808,N_6089,N_6372);
xnor U8809 (N_8809,N_5567,N_5563);
xor U8810 (N_8810,N_5399,N_5139);
and U8811 (N_8811,N_5807,N_6730);
and U8812 (N_8812,N_7279,N_6956);
nor U8813 (N_8813,N_5002,N_5806);
nand U8814 (N_8814,N_6700,N_6650);
nor U8815 (N_8815,N_6191,N_5689);
xnor U8816 (N_8816,N_6812,N_6093);
xor U8817 (N_8817,N_7338,N_7446);
nand U8818 (N_8818,N_5671,N_6429);
and U8819 (N_8819,N_5732,N_6601);
and U8820 (N_8820,N_5662,N_6744);
nand U8821 (N_8821,N_7363,N_6369);
and U8822 (N_8822,N_5920,N_7203);
xnor U8823 (N_8823,N_5685,N_7170);
nor U8824 (N_8824,N_6456,N_6999);
nand U8825 (N_8825,N_5466,N_6586);
xor U8826 (N_8826,N_7467,N_5158);
xnor U8827 (N_8827,N_6397,N_6685);
nand U8828 (N_8828,N_5242,N_5678);
nand U8829 (N_8829,N_5574,N_6362);
and U8830 (N_8830,N_6810,N_7107);
xor U8831 (N_8831,N_5314,N_7477);
and U8832 (N_8832,N_5452,N_5825);
nand U8833 (N_8833,N_5911,N_5749);
or U8834 (N_8834,N_6107,N_6960);
nor U8835 (N_8835,N_7271,N_6378);
xnor U8836 (N_8836,N_6228,N_5534);
xnor U8837 (N_8837,N_6522,N_5729);
xor U8838 (N_8838,N_6952,N_5866);
or U8839 (N_8839,N_6142,N_7178);
xor U8840 (N_8840,N_5829,N_5808);
xor U8841 (N_8841,N_6940,N_7283);
and U8842 (N_8842,N_7034,N_5619);
and U8843 (N_8843,N_6156,N_6802);
nand U8844 (N_8844,N_5460,N_6553);
and U8845 (N_8845,N_5671,N_6131);
nand U8846 (N_8846,N_6910,N_6329);
xor U8847 (N_8847,N_7042,N_5791);
and U8848 (N_8848,N_7106,N_6566);
nor U8849 (N_8849,N_5849,N_5113);
nand U8850 (N_8850,N_7463,N_7148);
or U8851 (N_8851,N_6523,N_5775);
and U8852 (N_8852,N_7476,N_5451);
and U8853 (N_8853,N_7456,N_5682);
and U8854 (N_8854,N_6706,N_7118);
nor U8855 (N_8855,N_7491,N_6656);
or U8856 (N_8856,N_5649,N_5825);
nand U8857 (N_8857,N_7343,N_7358);
xor U8858 (N_8858,N_6193,N_5470);
and U8859 (N_8859,N_5998,N_5750);
and U8860 (N_8860,N_5354,N_5638);
nor U8861 (N_8861,N_6721,N_7454);
or U8862 (N_8862,N_6155,N_7469);
or U8863 (N_8863,N_5829,N_6568);
or U8864 (N_8864,N_6555,N_5027);
nor U8865 (N_8865,N_6246,N_6690);
or U8866 (N_8866,N_6793,N_5682);
nor U8867 (N_8867,N_7009,N_6770);
and U8868 (N_8868,N_7246,N_6333);
or U8869 (N_8869,N_7138,N_6266);
and U8870 (N_8870,N_5778,N_5104);
nor U8871 (N_8871,N_6470,N_7388);
nand U8872 (N_8872,N_7100,N_5132);
xor U8873 (N_8873,N_5285,N_7042);
and U8874 (N_8874,N_7344,N_7392);
nor U8875 (N_8875,N_5567,N_6183);
or U8876 (N_8876,N_6083,N_5523);
or U8877 (N_8877,N_5476,N_6974);
and U8878 (N_8878,N_6204,N_5731);
nor U8879 (N_8879,N_6132,N_5179);
xor U8880 (N_8880,N_7313,N_5157);
nand U8881 (N_8881,N_5282,N_6059);
or U8882 (N_8882,N_6361,N_5601);
nand U8883 (N_8883,N_6667,N_5439);
or U8884 (N_8884,N_5956,N_5855);
and U8885 (N_8885,N_5089,N_7467);
nand U8886 (N_8886,N_5771,N_6933);
xor U8887 (N_8887,N_6005,N_5742);
nor U8888 (N_8888,N_7272,N_5111);
or U8889 (N_8889,N_5068,N_6969);
nand U8890 (N_8890,N_5668,N_7217);
xnor U8891 (N_8891,N_6982,N_7013);
or U8892 (N_8892,N_7116,N_5208);
or U8893 (N_8893,N_5169,N_5060);
nand U8894 (N_8894,N_5079,N_5647);
and U8895 (N_8895,N_6890,N_6820);
xnor U8896 (N_8896,N_6176,N_5034);
xnor U8897 (N_8897,N_5545,N_6181);
or U8898 (N_8898,N_6005,N_6343);
nor U8899 (N_8899,N_6955,N_6498);
xnor U8900 (N_8900,N_5119,N_6771);
xor U8901 (N_8901,N_7329,N_5094);
nor U8902 (N_8902,N_5377,N_6327);
nand U8903 (N_8903,N_7035,N_5450);
nor U8904 (N_8904,N_5264,N_5136);
and U8905 (N_8905,N_6085,N_6315);
nor U8906 (N_8906,N_5997,N_5812);
and U8907 (N_8907,N_7197,N_6575);
xnor U8908 (N_8908,N_5360,N_6275);
and U8909 (N_8909,N_6339,N_6513);
nor U8910 (N_8910,N_6837,N_5320);
nor U8911 (N_8911,N_6913,N_6066);
or U8912 (N_8912,N_6694,N_6519);
xnor U8913 (N_8913,N_5010,N_6682);
and U8914 (N_8914,N_5620,N_6257);
or U8915 (N_8915,N_7178,N_6775);
nor U8916 (N_8916,N_7288,N_5910);
and U8917 (N_8917,N_6048,N_7122);
or U8918 (N_8918,N_6615,N_5717);
nor U8919 (N_8919,N_6398,N_7323);
xor U8920 (N_8920,N_5069,N_5566);
xnor U8921 (N_8921,N_7116,N_5216);
or U8922 (N_8922,N_6289,N_5980);
or U8923 (N_8923,N_5324,N_6387);
or U8924 (N_8924,N_6876,N_6577);
nor U8925 (N_8925,N_6615,N_5362);
nor U8926 (N_8926,N_5326,N_5943);
nor U8927 (N_8927,N_6204,N_6650);
nor U8928 (N_8928,N_5375,N_7160);
nand U8929 (N_8929,N_7322,N_5527);
nand U8930 (N_8930,N_7081,N_5295);
or U8931 (N_8931,N_6824,N_6204);
nand U8932 (N_8932,N_5935,N_7422);
xnor U8933 (N_8933,N_6684,N_6038);
nand U8934 (N_8934,N_6314,N_6319);
xor U8935 (N_8935,N_7075,N_5668);
or U8936 (N_8936,N_7259,N_6476);
xor U8937 (N_8937,N_6855,N_6566);
or U8938 (N_8938,N_7042,N_6468);
xor U8939 (N_8939,N_5163,N_5524);
nand U8940 (N_8940,N_5341,N_6764);
and U8941 (N_8941,N_7434,N_6699);
nand U8942 (N_8942,N_5076,N_5462);
nand U8943 (N_8943,N_6947,N_6629);
nor U8944 (N_8944,N_6422,N_7317);
nor U8945 (N_8945,N_6307,N_5284);
and U8946 (N_8946,N_5900,N_6775);
or U8947 (N_8947,N_5480,N_5890);
nor U8948 (N_8948,N_5492,N_7051);
nand U8949 (N_8949,N_6060,N_7184);
or U8950 (N_8950,N_7469,N_6327);
nor U8951 (N_8951,N_6845,N_7254);
and U8952 (N_8952,N_7484,N_7257);
or U8953 (N_8953,N_7209,N_5841);
xnor U8954 (N_8954,N_5242,N_7186);
and U8955 (N_8955,N_6990,N_5725);
nand U8956 (N_8956,N_6668,N_7002);
xor U8957 (N_8957,N_6318,N_6236);
or U8958 (N_8958,N_5903,N_5691);
xor U8959 (N_8959,N_6719,N_5655);
nand U8960 (N_8960,N_6817,N_7217);
and U8961 (N_8961,N_5203,N_5024);
nor U8962 (N_8962,N_7282,N_7246);
and U8963 (N_8963,N_6094,N_5296);
xor U8964 (N_8964,N_5475,N_6578);
and U8965 (N_8965,N_6169,N_5643);
xnor U8966 (N_8966,N_6217,N_6560);
and U8967 (N_8967,N_6320,N_6215);
xnor U8968 (N_8968,N_6921,N_6508);
nor U8969 (N_8969,N_5067,N_7371);
nor U8970 (N_8970,N_5473,N_7044);
nand U8971 (N_8971,N_5651,N_7248);
xor U8972 (N_8972,N_6890,N_6252);
and U8973 (N_8973,N_6869,N_7469);
and U8974 (N_8974,N_5536,N_5584);
nand U8975 (N_8975,N_5337,N_5458);
xnor U8976 (N_8976,N_5111,N_7163);
nand U8977 (N_8977,N_5358,N_6264);
and U8978 (N_8978,N_5791,N_5233);
nand U8979 (N_8979,N_5240,N_5888);
nor U8980 (N_8980,N_5754,N_5233);
and U8981 (N_8981,N_7183,N_6391);
nor U8982 (N_8982,N_7105,N_6872);
nor U8983 (N_8983,N_6935,N_5979);
or U8984 (N_8984,N_6787,N_5344);
and U8985 (N_8985,N_6893,N_7053);
xnor U8986 (N_8986,N_5637,N_5492);
nor U8987 (N_8987,N_6528,N_6954);
xor U8988 (N_8988,N_7286,N_6937);
xnor U8989 (N_8989,N_5118,N_6342);
nand U8990 (N_8990,N_6578,N_6788);
or U8991 (N_8991,N_5117,N_5016);
or U8992 (N_8992,N_5844,N_7098);
nand U8993 (N_8993,N_6910,N_6447);
and U8994 (N_8994,N_5272,N_6550);
nor U8995 (N_8995,N_6577,N_6031);
nor U8996 (N_8996,N_5319,N_6589);
or U8997 (N_8997,N_6485,N_5322);
xnor U8998 (N_8998,N_6010,N_5527);
and U8999 (N_8999,N_6087,N_6626);
nand U9000 (N_9000,N_5105,N_6829);
and U9001 (N_9001,N_6374,N_6384);
or U9002 (N_9002,N_7469,N_7065);
and U9003 (N_9003,N_6987,N_5224);
nor U9004 (N_9004,N_7241,N_7024);
nor U9005 (N_9005,N_6668,N_6388);
and U9006 (N_9006,N_6954,N_6779);
xor U9007 (N_9007,N_5672,N_5493);
or U9008 (N_9008,N_5605,N_7317);
and U9009 (N_9009,N_6905,N_5115);
or U9010 (N_9010,N_7138,N_6035);
and U9011 (N_9011,N_6739,N_5084);
nor U9012 (N_9012,N_7258,N_5958);
xnor U9013 (N_9013,N_7348,N_6747);
xor U9014 (N_9014,N_6709,N_5657);
xor U9015 (N_9015,N_5946,N_7304);
nor U9016 (N_9016,N_6922,N_5227);
nand U9017 (N_9017,N_5112,N_6917);
xnor U9018 (N_9018,N_6336,N_5150);
nor U9019 (N_9019,N_6629,N_7491);
nor U9020 (N_9020,N_6994,N_5616);
nor U9021 (N_9021,N_5605,N_5073);
xor U9022 (N_9022,N_5577,N_6006);
and U9023 (N_9023,N_6619,N_7045);
nand U9024 (N_9024,N_6821,N_7336);
and U9025 (N_9025,N_7099,N_6951);
nand U9026 (N_9026,N_5816,N_6602);
nand U9027 (N_9027,N_5888,N_5830);
nand U9028 (N_9028,N_7247,N_5319);
xnor U9029 (N_9029,N_6629,N_5732);
nor U9030 (N_9030,N_7308,N_5634);
and U9031 (N_9031,N_6900,N_6451);
nor U9032 (N_9032,N_6626,N_5863);
nand U9033 (N_9033,N_6179,N_5089);
and U9034 (N_9034,N_6672,N_6847);
nand U9035 (N_9035,N_5408,N_5836);
nor U9036 (N_9036,N_5193,N_6813);
nor U9037 (N_9037,N_5913,N_5902);
and U9038 (N_9038,N_5527,N_6905);
or U9039 (N_9039,N_6785,N_5896);
nand U9040 (N_9040,N_5063,N_7280);
xnor U9041 (N_9041,N_5778,N_5668);
and U9042 (N_9042,N_5131,N_6010);
xnor U9043 (N_9043,N_6188,N_5656);
nor U9044 (N_9044,N_6282,N_6030);
or U9045 (N_9045,N_6715,N_5049);
nand U9046 (N_9046,N_7221,N_6017);
or U9047 (N_9047,N_6565,N_6792);
nor U9048 (N_9048,N_7156,N_5252);
nor U9049 (N_9049,N_7044,N_6589);
and U9050 (N_9050,N_7453,N_6597);
xnor U9051 (N_9051,N_6809,N_6067);
or U9052 (N_9052,N_6244,N_5256);
xor U9053 (N_9053,N_6975,N_7297);
and U9054 (N_9054,N_5288,N_6990);
or U9055 (N_9055,N_5352,N_5786);
nand U9056 (N_9056,N_5519,N_6323);
and U9057 (N_9057,N_6222,N_6403);
and U9058 (N_9058,N_5399,N_6045);
nor U9059 (N_9059,N_6559,N_6036);
xnor U9060 (N_9060,N_5511,N_5892);
or U9061 (N_9061,N_5190,N_5564);
xnor U9062 (N_9062,N_5021,N_6219);
xor U9063 (N_9063,N_6991,N_7294);
and U9064 (N_9064,N_5613,N_6686);
nor U9065 (N_9065,N_7300,N_6807);
or U9066 (N_9066,N_6290,N_5820);
and U9067 (N_9067,N_5845,N_6932);
or U9068 (N_9068,N_5427,N_6336);
or U9069 (N_9069,N_5748,N_6282);
and U9070 (N_9070,N_7213,N_7457);
nand U9071 (N_9071,N_6234,N_5186);
xor U9072 (N_9072,N_6674,N_6894);
or U9073 (N_9073,N_5590,N_6958);
nand U9074 (N_9074,N_6524,N_7032);
nand U9075 (N_9075,N_5479,N_6327);
or U9076 (N_9076,N_5851,N_6059);
xor U9077 (N_9077,N_7194,N_7172);
or U9078 (N_9078,N_5582,N_7426);
xnor U9079 (N_9079,N_6087,N_6133);
or U9080 (N_9080,N_6121,N_5688);
and U9081 (N_9081,N_6276,N_6858);
and U9082 (N_9082,N_7181,N_6186);
nor U9083 (N_9083,N_6402,N_6272);
nor U9084 (N_9084,N_6658,N_5717);
nand U9085 (N_9085,N_5145,N_7408);
or U9086 (N_9086,N_7060,N_7253);
xnor U9087 (N_9087,N_7270,N_6079);
and U9088 (N_9088,N_6590,N_5641);
or U9089 (N_9089,N_6417,N_7412);
xor U9090 (N_9090,N_7406,N_7342);
nor U9091 (N_9091,N_5017,N_6100);
nand U9092 (N_9092,N_7183,N_5469);
xnor U9093 (N_9093,N_6463,N_6190);
nand U9094 (N_9094,N_6290,N_5667);
and U9095 (N_9095,N_7478,N_7365);
nor U9096 (N_9096,N_6961,N_7381);
and U9097 (N_9097,N_7257,N_6523);
xnor U9098 (N_9098,N_6670,N_5263);
xor U9099 (N_9099,N_6016,N_6055);
xnor U9100 (N_9100,N_5622,N_7041);
or U9101 (N_9101,N_7079,N_5207);
or U9102 (N_9102,N_6264,N_7287);
or U9103 (N_9103,N_6480,N_5870);
xnor U9104 (N_9104,N_6520,N_7036);
nand U9105 (N_9105,N_6735,N_5443);
or U9106 (N_9106,N_7152,N_5499);
nand U9107 (N_9107,N_7302,N_6959);
nor U9108 (N_9108,N_7059,N_6564);
xor U9109 (N_9109,N_7330,N_6511);
xnor U9110 (N_9110,N_5899,N_7460);
xor U9111 (N_9111,N_5022,N_5259);
xor U9112 (N_9112,N_7460,N_6937);
or U9113 (N_9113,N_6554,N_5847);
and U9114 (N_9114,N_6562,N_6186);
or U9115 (N_9115,N_6308,N_6064);
and U9116 (N_9116,N_6622,N_5733);
nand U9117 (N_9117,N_5577,N_6397);
nor U9118 (N_9118,N_5639,N_6603);
nor U9119 (N_9119,N_6223,N_5859);
xnor U9120 (N_9120,N_6032,N_5998);
or U9121 (N_9121,N_6323,N_5096);
or U9122 (N_9122,N_6869,N_5984);
and U9123 (N_9123,N_6542,N_6791);
nand U9124 (N_9124,N_7063,N_6411);
or U9125 (N_9125,N_6670,N_6260);
and U9126 (N_9126,N_6786,N_6192);
nor U9127 (N_9127,N_5241,N_5431);
xnor U9128 (N_9128,N_6839,N_6364);
and U9129 (N_9129,N_5410,N_5990);
xor U9130 (N_9130,N_5097,N_6824);
nand U9131 (N_9131,N_5488,N_5475);
or U9132 (N_9132,N_6180,N_6807);
or U9133 (N_9133,N_6384,N_6354);
xnor U9134 (N_9134,N_5912,N_6412);
nor U9135 (N_9135,N_6044,N_5992);
or U9136 (N_9136,N_7499,N_6868);
xor U9137 (N_9137,N_5758,N_6698);
or U9138 (N_9138,N_5827,N_5706);
xnor U9139 (N_9139,N_5023,N_6442);
nor U9140 (N_9140,N_7063,N_5501);
xor U9141 (N_9141,N_5082,N_6561);
xnor U9142 (N_9142,N_7165,N_5457);
xnor U9143 (N_9143,N_5929,N_5905);
nand U9144 (N_9144,N_5822,N_6274);
or U9145 (N_9145,N_6486,N_5797);
xor U9146 (N_9146,N_7254,N_6834);
nand U9147 (N_9147,N_7426,N_5817);
nand U9148 (N_9148,N_5142,N_5183);
or U9149 (N_9149,N_5646,N_6089);
or U9150 (N_9150,N_5953,N_6720);
xnor U9151 (N_9151,N_5120,N_5891);
and U9152 (N_9152,N_5366,N_5609);
and U9153 (N_9153,N_5454,N_7011);
nand U9154 (N_9154,N_5546,N_6465);
nor U9155 (N_9155,N_6641,N_5959);
nand U9156 (N_9156,N_5699,N_5213);
nand U9157 (N_9157,N_5561,N_7270);
nand U9158 (N_9158,N_7450,N_6756);
nor U9159 (N_9159,N_5597,N_5177);
or U9160 (N_9160,N_7351,N_5968);
xnor U9161 (N_9161,N_7281,N_7196);
and U9162 (N_9162,N_5772,N_7126);
or U9163 (N_9163,N_6561,N_5159);
or U9164 (N_9164,N_6082,N_5024);
nor U9165 (N_9165,N_5351,N_6843);
or U9166 (N_9166,N_6403,N_6458);
xor U9167 (N_9167,N_7388,N_5470);
nand U9168 (N_9168,N_5847,N_6171);
and U9169 (N_9169,N_5290,N_7034);
or U9170 (N_9170,N_5709,N_5333);
nand U9171 (N_9171,N_5662,N_7250);
nand U9172 (N_9172,N_5970,N_7209);
or U9173 (N_9173,N_7121,N_6953);
or U9174 (N_9174,N_6035,N_5221);
or U9175 (N_9175,N_5212,N_6514);
xnor U9176 (N_9176,N_6379,N_7354);
and U9177 (N_9177,N_6049,N_5640);
xnor U9178 (N_9178,N_6091,N_5847);
or U9179 (N_9179,N_5673,N_5485);
or U9180 (N_9180,N_7291,N_5247);
nor U9181 (N_9181,N_6170,N_5853);
or U9182 (N_9182,N_6711,N_5298);
and U9183 (N_9183,N_7233,N_6978);
xor U9184 (N_9184,N_5965,N_5943);
and U9185 (N_9185,N_6080,N_5696);
nand U9186 (N_9186,N_7055,N_7442);
nor U9187 (N_9187,N_6640,N_5377);
and U9188 (N_9188,N_6271,N_7248);
or U9189 (N_9189,N_6994,N_6239);
nor U9190 (N_9190,N_6740,N_5071);
or U9191 (N_9191,N_5715,N_5490);
and U9192 (N_9192,N_5695,N_6038);
and U9193 (N_9193,N_5514,N_7259);
nor U9194 (N_9194,N_6141,N_5518);
or U9195 (N_9195,N_6337,N_6118);
or U9196 (N_9196,N_7039,N_5689);
or U9197 (N_9197,N_5164,N_5887);
nor U9198 (N_9198,N_5429,N_5994);
and U9199 (N_9199,N_6106,N_5137);
xnor U9200 (N_9200,N_5909,N_5136);
nor U9201 (N_9201,N_5959,N_6600);
xnor U9202 (N_9202,N_6874,N_6349);
or U9203 (N_9203,N_6501,N_5506);
xnor U9204 (N_9204,N_7383,N_5123);
nand U9205 (N_9205,N_5046,N_5271);
or U9206 (N_9206,N_6742,N_5799);
and U9207 (N_9207,N_5164,N_7070);
nor U9208 (N_9208,N_6818,N_7391);
or U9209 (N_9209,N_6884,N_6721);
and U9210 (N_9210,N_6862,N_5187);
xnor U9211 (N_9211,N_6409,N_6305);
and U9212 (N_9212,N_5406,N_7266);
xor U9213 (N_9213,N_5366,N_6418);
nor U9214 (N_9214,N_5427,N_5370);
xor U9215 (N_9215,N_5840,N_6134);
xnor U9216 (N_9216,N_5158,N_6292);
xnor U9217 (N_9217,N_7227,N_5737);
and U9218 (N_9218,N_5125,N_5717);
xnor U9219 (N_9219,N_6219,N_7262);
nand U9220 (N_9220,N_6603,N_5929);
nor U9221 (N_9221,N_5320,N_6065);
or U9222 (N_9222,N_7040,N_5171);
nor U9223 (N_9223,N_6962,N_6076);
xnor U9224 (N_9224,N_6568,N_6049);
nand U9225 (N_9225,N_5356,N_5648);
xor U9226 (N_9226,N_7350,N_5568);
and U9227 (N_9227,N_5261,N_6549);
nand U9228 (N_9228,N_5153,N_7228);
and U9229 (N_9229,N_5439,N_6177);
or U9230 (N_9230,N_5862,N_5610);
nor U9231 (N_9231,N_5764,N_5494);
xor U9232 (N_9232,N_6331,N_5524);
nor U9233 (N_9233,N_6188,N_5378);
or U9234 (N_9234,N_7275,N_5639);
or U9235 (N_9235,N_6924,N_6746);
and U9236 (N_9236,N_7492,N_6367);
nand U9237 (N_9237,N_5589,N_7225);
nand U9238 (N_9238,N_7009,N_7280);
nand U9239 (N_9239,N_7037,N_7025);
or U9240 (N_9240,N_5093,N_6682);
nor U9241 (N_9241,N_6520,N_5785);
and U9242 (N_9242,N_6065,N_6682);
nor U9243 (N_9243,N_7003,N_5313);
and U9244 (N_9244,N_6716,N_7322);
nor U9245 (N_9245,N_5134,N_6818);
or U9246 (N_9246,N_7316,N_6695);
xnor U9247 (N_9247,N_5468,N_5480);
nand U9248 (N_9248,N_6151,N_5400);
xnor U9249 (N_9249,N_6228,N_6015);
nand U9250 (N_9250,N_5558,N_6615);
nor U9251 (N_9251,N_7076,N_6745);
nand U9252 (N_9252,N_6121,N_5823);
or U9253 (N_9253,N_6343,N_5783);
and U9254 (N_9254,N_5616,N_6751);
nor U9255 (N_9255,N_6064,N_5083);
and U9256 (N_9256,N_7101,N_7225);
nand U9257 (N_9257,N_5463,N_7051);
nand U9258 (N_9258,N_6317,N_5464);
nor U9259 (N_9259,N_6702,N_5271);
nand U9260 (N_9260,N_6324,N_6515);
xor U9261 (N_9261,N_6074,N_5775);
or U9262 (N_9262,N_5655,N_5268);
and U9263 (N_9263,N_5650,N_5259);
or U9264 (N_9264,N_7345,N_5522);
or U9265 (N_9265,N_5328,N_5437);
xnor U9266 (N_9266,N_7221,N_5076);
nand U9267 (N_9267,N_7022,N_6720);
and U9268 (N_9268,N_7417,N_6610);
nand U9269 (N_9269,N_5899,N_6781);
and U9270 (N_9270,N_5282,N_5997);
xnor U9271 (N_9271,N_5744,N_6116);
nand U9272 (N_9272,N_7046,N_6033);
and U9273 (N_9273,N_7118,N_6015);
nand U9274 (N_9274,N_5804,N_5559);
or U9275 (N_9275,N_6088,N_7255);
nor U9276 (N_9276,N_6941,N_5098);
nand U9277 (N_9277,N_7404,N_7450);
or U9278 (N_9278,N_6290,N_6802);
nor U9279 (N_9279,N_6864,N_6214);
xor U9280 (N_9280,N_5730,N_5499);
nor U9281 (N_9281,N_5875,N_5224);
nand U9282 (N_9282,N_6790,N_6705);
xnor U9283 (N_9283,N_7044,N_6827);
xnor U9284 (N_9284,N_6443,N_5018);
nand U9285 (N_9285,N_7495,N_5820);
nand U9286 (N_9286,N_5431,N_7086);
nand U9287 (N_9287,N_5353,N_6015);
and U9288 (N_9288,N_5840,N_5446);
nor U9289 (N_9289,N_5482,N_6183);
nor U9290 (N_9290,N_5431,N_7357);
or U9291 (N_9291,N_5439,N_6236);
nor U9292 (N_9292,N_7065,N_5057);
nor U9293 (N_9293,N_5264,N_5005);
nor U9294 (N_9294,N_6083,N_6818);
xor U9295 (N_9295,N_7472,N_5550);
nand U9296 (N_9296,N_5785,N_6313);
or U9297 (N_9297,N_7188,N_5090);
xnor U9298 (N_9298,N_6861,N_5615);
or U9299 (N_9299,N_6955,N_6055);
nand U9300 (N_9300,N_5210,N_6697);
and U9301 (N_9301,N_5149,N_7392);
nor U9302 (N_9302,N_5181,N_5165);
nand U9303 (N_9303,N_6373,N_6598);
nand U9304 (N_9304,N_5929,N_5148);
or U9305 (N_9305,N_6870,N_6484);
xnor U9306 (N_9306,N_6872,N_6727);
nor U9307 (N_9307,N_6833,N_5135);
and U9308 (N_9308,N_7408,N_6706);
and U9309 (N_9309,N_6667,N_6301);
nor U9310 (N_9310,N_6706,N_6246);
nor U9311 (N_9311,N_6020,N_6239);
nor U9312 (N_9312,N_7325,N_6425);
nor U9313 (N_9313,N_5769,N_5538);
nor U9314 (N_9314,N_6798,N_6254);
nor U9315 (N_9315,N_5747,N_5769);
xnor U9316 (N_9316,N_6181,N_5682);
xnor U9317 (N_9317,N_6212,N_5237);
nor U9318 (N_9318,N_6067,N_6759);
and U9319 (N_9319,N_7397,N_5982);
nor U9320 (N_9320,N_6674,N_6135);
xor U9321 (N_9321,N_6058,N_6721);
nor U9322 (N_9322,N_6091,N_6609);
nand U9323 (N_9323,N_5253,N_7159);
xnor U9324 (N_9324,N_6393,N_5316);
and U9325 (N_9325,N_7405,N_6390);
xor U9326 (N_9326,N_6702,N_6839);
or U9327 (N_9327,N_6452,N_6792);
nor U9328 (N_9328,N_6452,N_6423);
nand U9329 (N_9329,N_6444,N_6270);
and U9330 (N_9330,N_5028,N_6073);
nor U9331 (N_9331,N_5426,N_6092);
and U9332 (N_9332,N_5519,N_6859);
nor U9333 (N_9333,N_7179,N_7142);
or U9334 (N_9334,N_6292,N_6909);
nand U9335 (N_9335,N_6164,N_5538);
nor U9336 (N_9336,N_6344,N_6614);
and U9337 (N_9337,N_6841,N_6235);
nor U9338 (N_9338,N_5736,N_7272);
nand U9339 (N_9339,N_7402,N_5788);
nor U9340 (N_9340,N_5557,N_6641);
xnor U9341 (N_9341,N_5134,N_5081);
xnor U9342 (N_9342,N_6465,N_6326);
xor U9343 (N_9343,N_7170,N_7141);
nor U9344 (N_9344,N_6960,N_6835);
and U9345 (N_9345,N_5308,N_6178);
or U9346 (N_9346,N_6930,N_7446);
or U9347 (N_9347,N_5407,N_5744);
nor U9348 (N_9348,N_5431,N_6318);
nor U9349 (N_9349,N_6730,N_5598);
nand U9350 (N_9350,N_6101,N_6115);
nand U9351 (N_9351,N_5759,N_6184);
or U9352 (N_9352,N_6457,N_6987);
nor U9353 (N_9353,N_6281,N_5337);
or U9354 (N_9354,N_5821,N_5498);
or U9355 (N_9355,N_7236,N_5944);
nand U9356 (N_9356,N_6048,N_6441);
xor U9357 (N_9357,N_6328,N_5661);
and U9358 (N_9358,N_5648,N_5286);
nand U9359 (N_9359,N_6746,N_6386);
nor U9360 (N_9360,N_6490,N_6397);
or U9361 (N_9361,N_7397,N_5620);
and U9362 (N_9362,N_5547,N_5793);
xnor U9363 (N_9363,N_6940,N_5598);
nand U9364 (N_9364,N_5256,N_7454);
xnor U9365 (N_9365,N_5408,N_6893);
nand U9366 (N_9366,N_7335,N_5869);
xnor U9367 (N_9367,N_7374,N_6631);
and U9368 (N_9368,N_5005,N_5382);
nand U9369 (N_9369,N_7262,N_5623);
and U9370 (N_9370,N_6619,N_7285);
xnor U9371 (N_9371,N_7070,N_7431);
nand U9372 (N_9372,N_6042,N_7098);
nor U9373 (N_9373,N_6839,N_7427);
xor U9374 (N_9374,N_6490,N_5762);
and U9375 (N_9375,N_5478,N_6794);
xor U9376 (N_9376,N_5238,N_5025);
nand U9377 (N_9377,N_7369,N_5620);
and U9378 (N_9378,N_5778,N_6552);
xnor U9379 (N_9379,N_5623,N_6385);
xor U9380 (N_9380,N_7172,N_6529);
nand U9381 (N_9381,N_7137,N_6738);
or U9382 (N_9382,N_6364,N_5942);
xnor U9383 (N_9383,N_6361,N_5061);
or U9384 (N_9384,N_5452,N_7156);
nand U9385 (N_9385,N_6719,N_6636);
and U9386 (N_9386,N_5810,N_6446);
or U9387 (N_9387,N_6743,N_7124);
xor U9388 (N_9388,N_6055,N_7058);
nand U9389 (N_9389,N_6662,N_7164);
nor U9390 (N_9390,N_6919,N_6017);
or U9391 (N_9391,N_6666,N_6053);
and U9392 (N_9392,N_5636,N_5352);
or U9393 (N_9393,N_5947,N_6412);
and U9394 (N_9394,N_5930,N_5666);
or U9395 (N_9395,N_6871,N_6464);
nor U9396 (N_9396,N_7194,N_5140);
nand U9397 (N_9397,N_7449,N_6580);
nand U9398 (N_9398,N_5566,N_5052);
nand U9399 (N_9399,N_6106,N_6152);
xnor U9400 (N_9400,N_5965,N_5736);
xor U9401 (N_9401,N_6487,N_6823);
nor U9402 (N_9402,N_5355,N_7198);
xor U9403 (N_9403,N_5844,N_6959);
nor U9404 (N_9404,N_6238,N_5811);
nand U9405 (N_9405,N_6656,N_5425);
xnor U9406 (N_9406,N_6392,N_5937);
and U9407 (N_9407,N_5457,N_7119);
and U9408 (N_9408,N_6284,N_6420);
nor U9409 (N_9409,N_5595,N_6710);
nand U9410 (N_9410,N_5799,N_5255);
nand U9411 (N_9411,N_5669,N_5544);
or U9412 (N_9412,N_5854,N_7272);
and U9413 (N_9413,N_5384,N_6684);
xnor U9414 (N_9414,N_6291,N_7483);
nor U9415 (N_9415,N_6953,N_6352);
and U9416 (N_9416,N_6234,N_5615);
and U9417 (N_9417,N_5437,N_6024);
nor U9418 (N_9418,N_5669,N_7166);
nor U9419 (N_9419,N_5312,N_6676);
nand U9420 (N_9420,N_6548,N_6598);
and U9421 (N_9421,N_6540,N_5694);
xnor U9422 (N_9422,N_5332,N_5743);
and U9423 (N_9423,N_5766,N_5981);
nor U9424 (N_9424,N_6161,N_6229);
and U9425 (N_9425,N_5811,N_6917);
nand U9426 (N_9426,N_6091,N_6499);
nor U9427 (N_9427,N_5733,N_5761);
xnor U9428 (N_9428,N_5835,N_6497);
nor U9429 (N_9429,N_6175,N_5419);
nor U9430 (N_9430,N_5453,N_7247);
xor U9431 (N_9431,N_5249,N_6701);
nand U9432 (N_9432,N_6065,N_6149);
xor U9433 (N_9433,N_6372,N_5444);
or U9434 (N_9434,N_5350,N_5101);
nor U9435 (N_9435,N_6044,N_6560);
or U9436 (N_9436,N_6683,N_6303);
xnor U9437 (N_9437,N_5883,N_6997);
or U9438 (N_9438,N_6262,N_6194);
nor U9439 (N_9439,N_5429,N_5360);
nand U9440 (N_9440,N_5375,N_5250);
xor U9441 (N_9441,N_6627,N_6906);
nand U9442 (N_9442,N_5672,N_5135);
nand U9443 (N_9443,N_7435,N_5284);
nor U9444 (N_9444,N_7203,N_5393);
or U9445 (N_9445,N_5849,N_6287);
and U9446 (N_9446,N_6820,N_5438);
nand U9447 (N_9447,N_5293,N_5765);
nor U9448 (N_9448,N_5257,N_6121);
nor U9449 (N_9449,N_6762,N_5761);
nor U9450 (N_9450,N_6031,N_6275);
and U9451 (N_9451,N_5933,N_5268);
xor U9452 (N_9452,N_6640,N_6894);
nand U9453 (N_9453,N_7124,N_5588);
or U9454 (N_9454,N_5587,N_6907);
nand U9455 (N_9455,N_5080,N_5253);
nand U9456 (N_9456,N_5942,N_5893);
and U9457 (N_9457,N_5794,N_6955);
xnor U9458 (N_9458,N_6618,N_6296);
or U9459 (N_9459,N_5706,N_7199);
nor U9460 (N_9460,N_6342,N_5034);
or U9461 (N_9461,N_7135,N_6150);
nor U9462 (N_9462,N_5001,N_5022);
nor U9463 (N_9463,N_5380,N_5238);
nor U9464 (N_9464,N_5053,N_7195);
nand U9465 (N_9465,N_5175,N_5262);
nand U9466 (N_9466,N_6493,N_7337);
xor U9467 (N_9467,N_5431,N_6222);
or U9468 (N_9468,N_6016,N_6548);
nand U9469 (N_9469,N_7118,N_6872);
xnor U9470 (N_9470,N_5201,N_5867);
nor U9471 (N_9471,N_7262,N_6000);
xnor U9472 (N_9472,N_6296,N_6074);
or U9473 (N_9473,N_5800,N_7331);
or U9474 (N_9474,N_7190,N_5295);
and U9475 (N_9475,N_6106,N_5678);
and U9476 (N_9476,N_7297,N_5844);
xor U9477 (N_9477,N_7224,N_6520);
xor U9478 (N_9478,N_6947,N_7348);
and U9479 (N_9479,N_6898,N_6447);
nand U9480 (N_9480,N_7013,N_6686);
and U9481 (N_9481,N_7028,N_7082);
and U9482 (N_9482,N_5027,N_5792);
nor U9483 (N_9483,N_5358,N_5084);
or U9484 (N_9484,N_5463,N_7480);
nand U9485 (N_9485,N_5495,N_6647);
and U9486 (N_9486,N_6451,N_6887);
nor U9487 (N_9487,N_6010,N_6710);
nor U9488 (N_9488,N_7263,N_6127);
and U9489 (N_9489,N_7181,N_5016);
and U9490 (N_9490,N_6639,N_5921);
nand U9491 (N_9491,N_5320,N_5703);
nor U9492 (N_9492,N_5329,N_5732);
nand U9493 (N_9493,N_5247,N_5189);
and U9494 (N_9494,N_7201,N_5033);
nor U9495 (N_9495,N_6456,N_5951);
or U9496 (N_9496,N_6547,N_5537);
nor U9497 (N_9497,N_5548,N_7365);
xnor U9498 (N_9498,N_5411,N_6308);
and U9499 (N_9499,N_5572,N_5065);
nor U9500 (N_9500,N_7163,N_5689);
nor U9501 (N_9501,N_6123,N_7402);
nand U9502 (N_9502,N_6396,N_7313);
xor U9503 (N_9503,N_7309,N_5094);
xnor U9504 (N_9504,N_6290,N_5676);
and U9505 (N_9505,N_7104,N_7356);
xor U9506 (N_9506,N_5230,N_7233);
nor U9507 (N_9507,N_7016,N_6767);
and U9508 (N_9508,N_5164,N_6270);
and U9509 (N_9509,N_6988,N_7237);
and U9510 (N_9510,N_6161,N_6573);
nand U9511 (N_9511,N_5706,N_7387);
nand U9512 (N_9512,N_7164,N_5543);
and U9513 (N_9513,N_5348,N_5835);
xor U9514 (N_9514,N_6440,N_6817);
or U9515 (N_9515,N_6161,N_5259);
nand U9516 (N_9516,N_5616,N_5555);
xor U9517 (N_9517,N_6161,N_7176);
nand U9518 (N_9518,N_6414,N_6036);
xnor U9519 (N_9519,N_5549,N_6674);
xnor U9520 (N_9520,N_6040,N_5130);
or U9521 (N_9521,N_5692,N_5538);
and U9522 (N_9522,N_6379,N_6698);
nor U9523 (N_9523,N_6453,N_5965);
nor U9524 (N_9524,N_6054,N_6314);
xnor U9525 (N_9525,N_6964,N_6271);
xnor U9526 (N_9526,N_6445,N_5746);
and U9527 (N_9527,N_5583,N_6424);
or U9528 (N_9528,N_5843,N_7131);
and U9529 (N_9529,N_5700,N_7214);
xor U9530 (N_9530,N_5264,N_7221);
xor U9531 (N_9531,N_6553,N_7461);
and U9532 (N_9532,N_5858,N_6982);
nand U9533 (N_9533,N_7063,N_5080);
nor U9534 (N_9534,N_7204,N_6546);
nand U9535 (N_9535,N_6929,N_5532);
nand U9536 (N_9536,N_7258,N_5637);
nor U9537 (N_9537,N_5688,N_6824);
and U9538 (N_9538,N_6837,N_6759);
nand U9539 (N_9539,N_5551,N_5115);
nand U9540 (N_9540,N_6319,N_5632);
nand U9541 (N_9541,N_5887,N_6348);
or U9542 (N_9542,N_5206,N_5887);
and U9543 (N_9543,N_5600,N_6462);
nand U9544 (N_9544,N_6170,N_7106);
and U9545 (N_9545,N_7312,N_6612);
xor U9546 (N_9546,N_6989,N_5955);
and U9547 (N_9547,N_5050,N_6103);
nor U9548 (N_9548,N_6963,N_5003);
and U9549 (N_9549,N_5491,N_5334);
nor U9550 (N_9550,N_5958,N_6762);
or U9551 (N_9551,N_5955,N_5060);
or U9552 (N_9552,N_5407,N_5255);
xor U9553 (N_9553,N_5772,N_6069);
xnor U9554 (N_9554,N_5822,N_5320);
and U9555 (N_9555,N_7252,N_7228);
and U9556 (N_9556,N_5312,N_5695);
and U9557 (N_9557,N_7061,N_7135);
nor U9558 (N_9558,N_6130,N_5416);
or U9559 (N_9559,N_6262,N_5261);
or U9560 (N_9560,N_7380,N_6915);
nand U9561 (N_9561,N_6905,N_6466);
and U9562 (N_9562,N_6672,N_5536);
or U9563 (N_9563,N_5366,N_5349);
and U9564 (N_9564,N_5084,N_6329);
nand U9565 (N_9565,N_6251,N_7298);
or U9566 (N_9566,N_5063,N_6739);
xnor U9567 (N_9567,N_7085,N_6822);
and U9568 (N_9568,N_6440,N_5291);
nand U9569 (N_9569,N_7311,N_6725);
xor U9570 (N_9570,N_7310,N_5305);
nand U9571 (N_9571,N_6991,N_7251);
xor U9572 (N_9572,N_7067,N_6141);
or U9573 (N_9573,N_6557,N_5853);
or U9574 (N_9574,N_6312,N_5432);
or U9575 (N_9575,N_6376,N_6413);
or U9576 (N_9576,N_7355,N_5715);
and U9577 (N_9577,N_6317,N_6353);
nor U9578 (N_9578,N_5757,N_7421);
and U9579 (N_9579,N_7354,N_6878);
and U9580 (N_9580,N_5004,N_5150);
or U9581 (N_9581,N_7379,N_7086);
nand U9582 (N_9582,N_6941,N_5745);
or U9583 (N_9583,N_5418,N_5061);
xnor U9584 (N_9584,N_6858,N_6215);
and U9585 (N_9585,N_5612,N_6048);
or U9586 (N_9586,N_5866,N_5920);
or U9587 (N_9587,N_5208,N_5431);
or U9588 (N_9588,N_7398,N_7481);
xor U9589 (N_9589,N_6579,N_7488);
nor U9590 (N_9590,N_7097,N_6174);
and U9591 (N_9591,N_7208,N_5352);
nor U9592 (N_9592,N_6170,N_7377);
nand U9593 (N_9593,N_6796,N_6185);
or U9594 (N_9594,N_7173,N_6005);
and U9595 (N_9595,N_7428,N_7383);
or U9596 (N_9596,N_6047,N_6369);
nand U9597 (N_9597,N_7120,N_5234);
or U9598 (N_9598,N_5705,N_6515);
nand U9599 (N_9599,N_6230,N_5526);
nand U9600 (N_9600,N_7360,N_6801);
nor U9601 (N_9601,N_6768,N_5832);
nand U9602 (N_9602,N_6793,N_5875);
and U9603 (N_9603,N_6879,N_7039);
or U9604 (N_9604,N_5345,N_5952);
or U9605 (N_9605,N_5895,N_6483);
xor U9606 (N_9606,N_6856,N_6717);
and U9607 (N_9607,N_7272,N_5825);
nor U9608 (N_9608,N_5101,N_5523);
and U9609 (N_9609,N_6159,N_5443);
or U9610 (N_9610,N_6132,N_5039);
xor U9611 (N_9611,N_6883,N_6131);
xor U9612 (N_9612,N_5224,N_5133);
or U9613 (N_9613,N_6045,N_7063);
xor U9614 (N_9614,N_6291,N_5431);
nor U9615 (N_9615,N_7372,N_6225);
nand U9616 (N_9616,N_5887,N_7412);
nand U9617 (N_9617,N_6156,N_6046);
nor U9618 (N_9618,N_5572,N_5664);
xnor U9619 (N_9619,N_7307,N_5802);
xnor U9620 (N_9620,N_5507,N_5096);
nor U9621 (N_9621,N_6319,N_5818);
and U9622 (N_9622,N_5174,N_5120);
xnor U9623 (N_9623,N_7003,N_6977);
nand U9624 (N_9624,N_6672,N_7368);
xor U9625 (N_9625,N_6939,N_7279);
or U9626 (N_9626,N_6793,N_5329);
nor U9627 (N_9627,N_5021,N_7275);
nand U9628 (N_9628,N_6113,N_6650);
or U9629 (N_9629,N_5669,N_7193);
nor U9630 (N_9630,N_6864,N_7215);
nor U9631 (N_9631,N_7316,N_6251);
nand U9632 (N_9632,N_5416,N_5916);
and U9633 (N_9633,N_5379,N_5492);
nand U9634 (N_9634,N_7158,N_6714);
nand U9635 (N_9635,N_5013,N_5177);
and U9636 (N_9636,N_6833,N_6559);
nor U9637 (N_9637,N_6951,N_5324);
xor U9638 (N_9638,N_5751,N_5655);
nor U9639 (N_9639,N_5490,N_5690);
and U9640 (N_9640,N_5852,N_6292);
xnor U9641 (N_9641,N_6496,N_7358);
nor U9642 (N_9642,N_5543,N_5332);
and U9643 (N_9643,N_5485,N_6783);
nor U9644 (N_9644,N_7079,N_5188);
nand U9645 (N_9645,N_5471,N_5586);
nor U9646 (N_9646,N_7045,N_5312);
xor U9647 (N_9647,N_5990,N_6099);
nand U9648 (N_9648,N_6318,N_7310);
and U9649 (N_9649,N_6662,N_7489);
and U9650 (N_9650,N_5373,N_6554);
or U9651 (N_9651,N_6329,N_5940);
or U9652 (N_9652,N_7028,N_6505);
and U9653 (N_9653,N_5891,N_5690);
nor U9654 (N_9654,N_5886,N_6516);
xnor U9655 (N_9655,N_5220,N_6115);
or U9656 (N_9656,N_7086,N_6082);
nor U9657 (N_9657,N_5199,N_5314);
nand U9658 (N_9658,N_7009,N_5598);
nand U9659 (N_9659,N_6626,N_5600);
and U9660 (N_9660,N_5456,N_6449);
xor U9661 (N_9661,N_5666,N_6053);
nand U9662 (N_9662,N_5648,N_7332);
or U9663 (N_9663,N_7451,N_5180);
xnor U9664 (N_9664,N_7424,N_5603);
or U9665 (N_9665,N_6841,N_6588);
or U9666 (N_9666,N_7152,N_6781);
xor U9667 (N_9667,N_7367,N_6522);
nand U9668 (N_9668,N_7250,N_5888);
or U9669 (N_9669,N_6178,N_5044);
nand U9670 (N_9670,N_6480,N_5337);
nor U9671 (N_9671,N_6122,N_6829);
or U9672 (N_9672,N_5803,N_6366);
nor U9673 (N_9673,N_5431,N_6553);
and U9674 (N_9674,N_6541,N_5550);
or U9675 (N_9675,N_7047,N_6442);
nand U9676 (N_9676,N_5459,N_5302);
or U9677 (N_9677,N_6566,N_7419);
or U9678 (N_9678,N_6671,N_6438);
nand U9679 (N_9679,N_5763,N_7360);
or U9680 (N_9680,N_5776,N_7089);
and U9681 (N_9681,N_5788,N_5411);
and U9682 (N_9682,N_6899,N_6292);
nor U9683 (N_9683,N_6043,N_5905);
and U9684 (N_9684,N_5289,N_5493);
nor U9685 (N_9685,N_6211,N_5006);
nand U9686 (N_9686,N_5723,N_5946);
and U9687 (N_9687,N_6202,N_6951);
or U9688 (N_9688,N_5316,N_7081);
nor U9689 (N_9689,N_6487,N_5962);
xnor U9690 (N_9690,N_7108,N_5964);
and U9691 (N_9691,N_5660,N_5751);
or U9692 (N_9692,N_7441,N_5492);
xnor U9693 (N_9693,N_6206,N_5565);
and U9694 (N_9694,N_5764,N_6591);
nor U9695 (N_9695,N_6748,N_7009);
nor U9696 (N_9696,N_6978,N_6558);
or U9697 (N_9697,N_5879,N_7420);
nor U9698 (N_9698,N_5600,N_6019);
and U9699 (N_9699,N_7473,N_6217);
nand U9700 (N_9700,N_5289,N_6385);
xor U9701 (N_9701,N_5699,N_5996);
nand U9702 (N_9702,N_7392,N_7404);
nor U9703 (N_9703,N_5361,N_7012);
and U9704 (N_9704,N_5034,N_7035);
xnor U9705 (N_9705,N_6473,N_5659);
and U9706 (N_9706,N_5756,N_5183);
and U9707 (N_9707,N_6153,N_7149);
nand U9708 (N_9708,N_5425,N_7280);
nand U9709 (N_9709,N_5609,N_6155);
and U9710 (N_9710,N_6442,N_5690);
or U9711 (N_9711,N_5780,N_6578);
nand U9712 (N_9712,N_5400,N_5965);
nor U9713 (N_9713,N_6777,N_7125);
xor U9714 (N_9714,N_6694,N_7026);
nand U9715 (N_9715,N_7297,N_6493);
nor U9716 (N_9716,N_7102,N_5345);
or U9717 (N_9717,N_7049,N_5410);
xor U9718 (N_9718,N_5787,N_5402);
nor U9719 (N_9719,N_5320,N_5612);
nand U9720 (N_9720,N_5656,N_7218);
and U9721 (N_9721,N_5753,N_6995);
nor U9722 (N_9722,N_6848,N_6952);
nor U9723 (N_9723,N_5368,N_6463);
and U9724 (N_9724,N_7050,N_5413);
xnor U9725 (N_9725,N_6885,N_6585);
nand U9726 (N_9726,N_6002,N_6473);
and U9727 (N_9727,N_7213,N_6491);
and U9728 (N_9728,N_5088,N_5796);
nand U9729 (N_9729,N_6457,N_7159);
nor U9730 (N_9730,N_6647,N_6725);
or U9731 (N_9731,N_6862,N_7208);
nor U9732 (N_9732,N_6937,N_6139);
nor U9733 (N_9733,N_5791,N_6685);
nor U9734 (N_9734,N_7369,N_6162);
nand U9735 (N_9735,N_7419,N_6086);
or U9736 (N_9736,N_6653,N_6500);
nor U9737 (N_9737,N_5279,N_6284);
xnor U9738 (N_9738,N_6490,N_5012);
xor U9739 (N_9739,N_6092,N_7315);
xor U9740 (N_9740,N_5567,N_6707);
xnor U9741 (N_9741,N_6152,N_5810);
and U9742 (N_9742,N_7360,N_5622);
and U9743 (N_9743,N_5674,N_6866);
and U9744 (N_9744,N_6045,N_5535);
nor U9745 (N_9745,N_5135,N_6915);
and U9746 (N_9746,N_7477,N_5181);
or U9747 (N_9747,N_6468,N_5850);
or U9748 (N_9748,N_5190,N_5821);
nand U9749 (N_9749,N_6851,N_6378);
nor U9750 (N_9750,N_5913,N_6454);
and U9751 (N_9751,N_6387,N_6262);
nand U9752 (N_9752,N_5075,N_5093);
nor U9753 (N_9753,N_7480,N_5082);
or U9754 (N_9754,N_7069,N_6961);
xor U9755 (N_9755,N_5952,N_5279);
xor U9756 (N_9756,N_6363,N_5621);
nor U9757 (N_9757,N_5572,N_5517);
xor U9758 (N_9758,N_5796,N_6776);
nand U9759 (N_9759,N_7485,N_7461);
or U9760 (N_9760,N_6704,N_5705);
xnor U9761 (N_9761,N_6829,N_5766);
xnor U9762 (N_9762,N_6688,N_5590);
nand U9763 (N_9763,N_5371,N_7089);
or U9764 (N_9764,N_6255,N_5856);
xor U9765 (N_9765,N_5708,N_5897);
nand U9766 (N_9766,N_5374,N_5075);
and U9767 (N_9767,N_7111,N_6331);
or U9768 (N_9768,N_7153,N_5477);
and U9769 (N_9769,N_5264,N_6614);
xor U9770 (N_9770,N_6427,N_5462);
nand U9771 (N_9771,N_7288,N_5208);
nor U9772 (N_9772,N_5775,N_6911);
nor U9773 (N_9773,N_5957,N_5686);
nand U9774 (N_9774,N_6155,N_5399);
or U9775 (N_9775,N_6395,N_6998);
xor U9776 (N_9776,N_6666,N_5493);
and U9777 (N_9777,N_6185,N_6830);
or U9778 (N_9778,N_7471,N_6087);
xor U9779 (N_9779,N_5937,N_6923);
nand U9780 (N_9780,N_7301,N_5247);
nand U9781 (N_9781,N_6236,N_6056);
or U9782 (N_9782,N_6538,N_6511);
or U9783 (N_9783,N_5191,N_5333);
nor U9784 (N_9784,N_5151,N_5101);
nand U9785 (N_9785,N_6806,N_5936);
nand U9786 (N_9786,N_7259,N_5853);
and U9787 (N_9787,N_5930,N_7236);
or U9788 (N_9788,N_6727,N_6656);
nor U9789 (N_9789,N_5578,N_6681);
and U9790 (N_9790,N_5716,N_5578);
and U9791 (N_9791,N_5943,N_5822);
nand U9792 (N_9792,N_5806,N_5663);
and U9793 (N_9793,N_5896,N_6398);
or U9794 (N_9794,N_7062,N_7163);
or U9795 (N_9795,N_5223,N_5618);
nand U9796 (N_9796,N_5298,N_5134);
xor U9797 (N_9797,N_5872,N_6053);
or U9798 (N_9798,N_7056,N_6358);
or U9799 (N_9799,N_5061,N_5722);
xor U9800 (N_9800,N_7425,N_5315);
nand U9801 (N_9801,N_5285,N_5083);
nand U9802 (N_9802,N_5496,N_5646);
nor U9803 (N_9803,N_7140,N_5541);
nor U9804 (N_9804,N_7342,N_6004);
nor U9805 (N_9805,N_5813,N_5275);
nor U9806 (N_9806,N_5274,N_6954);
nand U9807 (N_9807,N_6869,N_7427);
or U9808 (N_9808,N_7275,N_5819);
or U9809 (N_9809,N_6631,N_5376);
xor U9810 (N_9810,N_6924,N_5888);
nand U9811 (N_9811,N_7380,N_5727);
xnor U9812 (N_9812,N_5279,N_6276);
and U9813 (N_9813,N_5383,N_5593);
and U9814 (N_9814,N_6882,N_5167);
or U9815 (N_9815,N_5714,N_7017);
xor U9816 (N_9816,N_7287,N_7272);
nand U9817 (N_9817,N_6189,N_6717);
and U9818 (N_9818,N_6871,N_5059);
xor U9819 (N_9819,N_5124,N_6576);
xnor U9820 (N_9820,N_5509,N_6771);
nand U9821 (N_9821,N_7382,N_5588);
nand U9822 (N_9822,N_6100,N_7424);
and U9823 (N_9823,N_5435,N_7105);
nor U9824 (N_9824,N_5827,N_5154);
xor U9825 (N_9825,N_6523,N_7463);
or U9826 (N_9826,N_6255,N_5364);
xor U9827 (N_9827,N_7266,N_5717);
nor U9828 (N_9828,N_6026,N_6031);
xnor U9829 (N_9829,N_6573,N_5836);
and U9830 (N_9830,N_6447,N_6099);
nor U9831 (N_9831,N_6470,N_5385);
or U9832 (N_9832,N_6684,N_5646);
or U9833 (N_9833,N_5504,N_5884);
nand U9834 (N_9834,N_6530,N_5920);
nand U9835 (N_9835,N_6635,N_6863);
and U9836 (N_9836,N_7141,N_6664);
xnor U9837 (N_9837,N_6374,N_5454);
and U9838 (N_9838,N_7212,N_6741);
nand U9839 (N_9839,N_7496,N_6376);
xor U9840 (N_9840,N_6787,N_7326);
xnor U9841 (N_9841,N_6612,N_6551);
nand U9842 (N_9842,N_6870,N_6313);
nand U9843 (N_9843,N_7368,N_5404);
or U9844 (N_9844,N_5156,N_6855);
and U9845 (N_9845,N_5449,N_6448);
xnor U9846 (N_9846,N_5179,N_5566);
or U9847 (N_9847,N_6517,N_6609);
nand U9848 (N_9848,N_6919,N_7381);
nor U9849 (N_9849,N_7491,N_6434);
xor U9850 (N_9850,N_5486,N_5243);
xnor U9851 (N_9851,N_6685,N_6503);
and U9852 (N_9852,N_5327,N_5471);
and U9853 (N_9853,N_6808,N_6691);
nand U9854 (N_9854,N_6116,N_6020);
or U9855 (N_9855,N_7388,N_5544);
nand U9856 (N_9856,N_7193,N_5634);
nor U9857 (N_9857,N_5738,N_5487);
xnor U9858 (N_9858,N_6739,N_5524);
nor U9859 (N_9859,N_5299,N_7305);
xnor U9860 (N_9860,N_5899,N_6099);
nor U9861 (N_9861,N_6213,N_6040);
xnor U9862 (N_9862,N_6218,N_6064);
xnor U9863 (N_9863,N_6492,N_5392);
or U9864 (N_9864,N_5159,N_6781);
xnor U9865 (N_9865,N_6856,N_6183);
nor U9866 (N_9866,N_6642,N_5690);
or U9867 (N_9867,N_7371,N_5493);
and U9868 (N_9868,N_6136,N_5622);
xor U9869 (N_9869,N_6972,N_6192);
and U9870 (N_9870,N_6638,N_5196);
xnor U9871 (N_9871,N_6846,N_6743);
xnor U9872 (N_9872,N_6315,N_7259);
nor U9873 (N_9873,N_5880,N_6771);
nand U9874 (N_9874,N_6702,N_7170);
xnor U9875 (N_9875,N_5082,N_6142);
and U9876 (N_9876,N_6815,N_7104);
nor U9877 (N_9877,N_5837,N_7396);
nor U9878 (N_9878,N_6676,N_6040);
nor U9879 (N_9879,N_5885,N_5455);
xor U9880 (N_9880,N_6895,N_5619);
nand U9881 (N_9881,N_6855,N_7438);
xor U9882 (N_9882,N_5975,N_6738);
and U9883 (N_9883,N_5246,N_5728);
nor U9884 (N_9884,N_5040,N_6909);
nand U9885 (N_9885,N_6977,N_6986);
nand U9886 (N_9886,N_5434,N_6312);
and U9887 (N_9887,N_6237,N_5532);
or U9888 (N_9888,N_6952,N_6143);
and U9889 (N_9889,N_7271,N_6537);
xor U9890 (N_9890,N_6007,N_5320);
nand U9891 (N_9891,N_5962,N_5792);
nor U9892 (N_9892,N_6924,N_7028);
nand U9893 (N_9893,N_7249,N_6785);
nor U9894 (N_9894,N_5375,N_6450);
xor U9895 (N_9895,N_5946,N_5259);
and U9896 (N_9896,N_6731,N_5631);
nor U9897 (N_9897,N_7264,N_5091);
nor U9898 (N_9898,N_6857,N_6483);
and U9899 (N_9899,N_5401,N_5443);
or U9900 (N_9900,N_6700,N_5028);
and U9901 (N_9901,N_5258,N_7256);
and U9902 (N_9902,N_5897,N_6655);
nand U9903 (N_9903,N_5836,N_5193);
nand U9904 (N_9904,N_6770,N_6486);
nand U9905 (N_9905,N_6265,N_5874);
xor U9906 (N_9906,N_6166,N_7014);
or U9907 (N_9907,N_7127,N_5085);
and U9908 (N_9908,N_7254,N_6794);
xnor U9909 (N_9909,N_6930,N_5304);
nand U9910 (N_9910,N_5594,N_5298);
nor U9911 (N_9911,N_5384,N_6960);
nand U9912 (N_9912,N_6795,N_5796);
xnor U9913 (N_9913,N_6406,N_6569);
nand U9914 (N_9914,N_6375,N_7239);
nor U9915 (N_9915,N_5522,N_5061);
nor U9916 (N_9916,N_6934,N_6191);
and U9917 (N_9917,N_6101,N_5905);
xor U9918 (N_9918,N_7286,N_6614);
xor U9919 (N_9919,N_6115,N_6512);
xnor U9920 (N_9920,N_6489,N_7471);
or U9921 (N_9921,N_7018,N_5038);
xnor U9922 (N_9922,N_5619,N_6934);
and U9923 (N_9923,N_5393,N_7477);
xor U9924 (N_9924,N_5382,N_6506);
and U9925 (N_9925,N_6379,N_7483);
and U9926 (N_9926,N_5028,N_6749);
or U9927 (N_9927,N_6418,N_6821);
nand U9928 (N_9928,N_7126,N_5816);
nor U9929 (N_9929,N_6454,N_5666);
xor U9930 (N_9930,N_7339,N_5699);
nand U9931 (N_9931,N_5570,N_5680);
or U9932 (N_9932,N_5860,N_5020);
and U9933 (N_9933,N_5125,N_6229);
xor U9934 (N_9934,N_5532,N_5183);
and U9935 (N_9935,N_6884,N_5487);
xnor U9936 (N_9936,N_6375,N_7342);
or U9937 (N_9937,N_6002,N_6947);
nand U9938 (N_9938,N_7179,N_6323);
and U9939 (N_9939,N_6645,N_6504);
nand U9940 (N_9940,N_5184,N_7220);
xnor U9941 (N_9941,N_6914,N_5588);
or U9942 (N_9942,N_6350,N_5188);
xnor U9943 (N_9943,N_6106,N_5431);
or U9944 (N_9944,N_5905,N_5001);
and U9945 (N_9945,N_6464,N_6118);
and U9946 (N_9946,N_5442,N_6772);
or U9947 (N_9947,N_7062,N_6391);
or U9948 (N_9948,N_6220,N_5838);
nand U9949 (N_9949,N_6241,N_5205);
nor U9950 (N_9950,N_5223,N_5815);
nand U9951 (N_9951,N_6734,N_6662);
and U9952 (N_9952,N_6690,N_6368);
and U9953 (N_9953,N_6976,N_6136);
nand U9954 (N_9954,N_5697,N_6428);
nand U9955 (N_9955,N_5501,N_7408);
and U9956 (N_9956,N_5373,N_5650);
and U9957 (N_9957,N_7223,N_5349);
nor U9958 (N_9958,N_6516,N_6323);
nand U9959 (N_9959,N_5044,N_6898);
or U9960 (N_9960,N_5635,N_5160);
or U9961 (N_9961,N_5401,N_5184);
nor U9962 (N_9962,N_5250,N_5912);
or U9963 (N_9963,N_5788,N_6523);
nand U9964 (N_9964,N_7243,N_6132);
and U9965 (N_9965,N_6658,N_7258);
and U9966 (N_9966,N_5562,N_5908);
nand U9967 (N_9967,N_6693,N_6530);
nand U9968 (N_9968,N_6591,N_5078);
nand U9969 (N_9969,N_7250,N_6823);
or U9970 (N_9970,N_5716,N_6405);
nor U9971 (N_9971,N_6091,N_7463);
or U9972 (N_9972,N_5124,N_7433);
or U9973 (N_9973,N_5689,N_7060);
xnor U9974 (N_9974,N_5133,N_5629);
and U9975 (N_9975,N_5288,N_5749);
and U9976 (N_9976,N_6231,N_5301);
or U9977 (N_9977,N_6299,N_6628);
nor U9978 (N_9978,N_5891,N_5595);
nand U9979 (N_9979,N_7376,N_5019);
or U9980 (N_9980,N_5104,N_6369);
xor U9981 (N_9981,N_6790,N_6409);
xor U9982 (N_9982,N_5481,N_7350);
nand U9983 (N_9983,N_6606,N_5652);
xnor U9984 (N_9984,N_6721,N_5023);
nand U9985 (N_9985,N_6774,N_5052);
nand U9986 (N_9986,N_5266,N_5714);
nand U9987 (N_9987,N_6000,N_5167);
nor U9988 (N_9988,N_7136,N_7469);
or U9989 (N_9989,N_5396,N_7439);
or U9990 (N_9990,N_5372,N_7260);
or U9991 (N_9991,N_6703,N_5059);
or U9992 (N_9992,N_5233,N_6696);
or U9993 (N_9993,N_7103,N_7227);
nor U9994 (N_9994,N_6607,N_6958);
xnor U9995 (N_9995,N_6633,N_5493);
xnor U9996 (N_9996,N_5926,N_6183);
nor U9997 (N_9997,N_5651,N_5091);
nor U9998 (N_9998,N_6033,N_5174);
or U9999 (N_9999,N_5906,N_5578);
nand UO_0 (O_0,N_8261,N_9788);
and UO_1 (O_1,N_9297,N_9374);
nor UO_2 (O_2,N_9579,N_9695);
nor UO_3 (O_3,N_9764,N_9000);
nor UO_4 (O_4,N_8691,N_8075);
nand UO_5 (O_5,N_9068,N_8052);
nor UO_6 (O_6,N_9699,N_9077);
xor UO_7 (O_7,N_8316,N_7665);
nor UO_8 (O_8,N_8095,N_7649);
xor UO_9 (O_9,N_9108,N_9658);
xnor UO_10 (O_10,N_8839,N_8670);
and UO_11 (O_11,N_8562,N_7854);
nor UO_12 (O_12,N_8388,N_7982);
nor UO_13 (O_13,N_9516,N_9005);
xnor UO_14 (O_14,N_8641,N_7821);
nor UO_15 (O_15,N_9765,N_8235);
nand UO_16 (O_16,N_8448,N_9295);
nand UO_17 (O_17,N_8460,N_7595);
or UO_18 (O_18,N_8440,N_9274);
nand UO_19 (O_19,N_9489,N_7747);
xnor UO_20 (O_20,N_8006,N_9288);
and UO_21 (O_21,N_8592,N_7704);
xnor UO_22 (O_22,N_9736,N_8512);
or UO_23 (O_23,N_9359,N_8395);
or UO_24 (O_24,N_7577,N_9133);
or UO_25 (O_25,N_7550,N_8738);
xor UO_26 (O_26,N_9460,N_7823);
nor UO_27 (O_27,N_8702,N_8265);
nand UO_28 (O_28,N_8736,N_8497);
nor UO_29 (O_29,N_9299,N_9267);
nor UO_30 (O_30,N_9845,N_9852);
nand UO_31 (O_31,N_8200,N_9661);
or UO_32 (O_32,N_8508,N_8994);
or UO_33 (O_33,N_9006,N_8314);
or UO_34 (O_34,N_9698,N_8864);
nor UO_35 (O_35,N_8809,N_8877);
and UO_36 (O_36,N_7906,N_9724);
nor UO_37 (O_37,N_7565,N_8124);
nor UO_38 (O_38,N_9450,N_7913);
nand UO_39 (O_39,N_8403,N_8014);
xnor UO_40 (O_40,N_9825,N_7500);
and UO_41 (O_41,N_9449,N_9200);
and UO_42 (O_42,N_8062,N_9749);
nand UO_43 (O_43,N_8746,N_8713);
nor UO_44 (O_44,N_7518,N_9697);
nor UO_45 (O_45,N_8367,N_8925);
nand UO_46 (O_46,N_9562,N_9790);
nor UO_47 (O_47,N_8791,N_8456);
and UO_48 (O_48,N_9254,N_9167);
and UO_49 (O_49,N_8682,N_8649);
xor UO_50 (O_50,N_8948,N_7922);
or UO_51 (O_51,N_9421,N_8930);
or UO_52 (O_52,N_7775,N_7613);
and UO_53 (O_53,N_9193,N_8607);
nor UO_54 (O_54,N_8897,N_8125);
or UO_55 (O_55,N_8960,N_9856);
or UO_56 (O_56,N_8179,N_7576);
and UO_57 (O_57,N_9387,N_8916);
nand UO_58 (O_58,N_7621,N_8459);
nor UO_59 (O_59,N_8424,N_9255);
and UO_60 (O_60,N_9090,N_9438);
or UO_61 (O_61,N_8548,N_8787);
or UO_62 (O_62,N_7637,N_8084);
nand UO_63 (O_63,N_7698,N_8374);
or UO_64 (O_64,N_8264,N_9269);
nor UO_65 (O_65,N_9596,N_7584);
and UO_66 (O_66,N_9178,N_9205);
xor UO_67 (O_67,N_9853,N_8131);
nor UO_68 (O_68,N_8701,N_7663);
or UO_69 (O_69,N_8222,N_9055);
xor UO_70 (O_70,N_8003,N_9545);
nor UO_71 (O_71,N_8704,N_9715);
and UO_72 (O_72,N_8248,N_8656);
nor UO_73 (O_73,N_7763,N_8441);
or UO_74 (O_74,N_8804,N_9160);
nor UO_75 (O_75,N_9147,N_9637);
or UO_76 (O_76,N_9215,N_8784);
xnor UO_77 (O_77,N_8438,N_7749);
xnor UO_78 (O_78,N_9426,N_9718);
or UO_79 (O_79,N_8573,N_8342);
nor UO_80 (O_80,N_8046,N_8636);
nand UO_81 (O_81,N_7623,N_9956);
nor UO_82 (O_82,N_7762,N_8333);
and UO_83 (O_83,N_9286,N_8490);
and UO_84 (O_84,N_8532,N_7596);
xnor UO_85 (O_85,N_8243,N_7607);
or UO_86 (O_86,N_8935,N_9702);
nor UO_87 (O_87,N_9456,N_8149);
and UO_88 (O_88,N_8580,N_9747);
or UO_89 (O_89,N_8435,N_7620);
or UO_90 (O_90,N_9007,N_8683);
nor UO_91 (O_91,N_9692,N_7758);
nor UO_92 (O_92,N_9879,N_9099);
nor UO_93 (O_93,N_8090,N_7836);
xnor UO_94 (O_94,N_8760,N_7547);
or UO_95 (O_95,N_7664,N_9491);
xor UO_96 (O_96,N_7598,N_7632);
or UO_97 (O_97,N_7514,N_7809);
nor UO_98 (O_98,N_9248,N_9835);
nor UO_99 (O_99,N_7880,N_9244);
nand UO_100 (O_100,N_8277,N_7626);
xor UO_101 (O_101,N_9534,N_9246);
or UO_102 (O_102,N_8345,N_7734);
nand UO_103 (O_103,N_7895,N_9739);
nand UO_104 (O_104,N_7805,N_9733);
nor UO_105 (O_105,N_9612,N_7509);
xnor UO_106 (O_106,N_8303,N_7594);
and UO_107 (O_107,N_7801,N_9549);
and UO_108 (O_108,N_8574,N_8962);
and UO_109 (O_109,N_8487,N_9506);
nor UO_110 (O_110,N_8624,N_7811);
nor UO_111 (O_111,N_8387,N_8069);
nor UO_112 (O_112,N_9618,N_7606);
xnor UO_113 (O_113,N_8833,N_8423);
or UO_114 (O_114,N_8537,N_8085);
xor UO_115 (O_115,N_7830,N_7671);
xor UO_116 (O_116,N_7817,N_7877);
xor UO_117 (O_117,N_7773,N_9798);
nor UO_118 (O_118,N_8807,N_8462);
nor UO_119 (O_119,N_9293,N_8304);
or UO_120 (O_120,N_9891,N_9253);
nand UO_121 (O_121,N_8461,N_8359);
nor UO_122 (O_122,N_7701,N_8128);
nand UO_123 (O_123,N_8584,N_9496);
or UO_124 (O_124,N_8789,N_9303);
or UO_125 (O_125,N_7683,N_8778);
or UO_126 (O_126,N_7693,N_7807);
and UO_127 (O_127,N_9581,N_8376);
nor UO_128 (O_128,N_7639,N_8365);
and UO_129 (O_129,N_9616,N_9560);
or UO_130 (O_130,N_8305,N_8059);
nor UO_131 (O_131,N_8337,N_9672);
or UO_132 (O_132,N_8381,N_9398);
xnor UO_133 (O_133,N_7988,N_7881);
or UO_134 (O_134,N_9732,N_9084);
or UO_135 (O_135,N_9706,N_8735);
or UO_136 (O_136,N_8765,N_8004);
nand UO_137 (O_137,N_8801,N_8141);
or UO_138 (O_138,N_9757,N_9360);
nor UO_139 (O_139,N_8500,N_9775);
and UO_140 (O_140,N_8744,N_9608);
or UO_141 (O_141,N_8126,N_9985);
xor UO_142 (O_142,N_8712,N_8457);
or UO_143 (O_143,N_9745,N_8266);
nor UO_144 (O_144,N_8215,N_7666);
nand UO_145 (O_145,N_7964,N_9582);
nand UO_146 (O_146,N_8521,N_9174);
nor UO_147 (O_147,N_8174,N_9002);
xnor UO_148 (O_148,N_8687,N_9164);
or UO_149 (O_149,N_9901,N_9479);
xnor UO_150 (O_150,N_8080,N_7923);
xor UO_151 (O_151,N_8282,N_8905);
nor UO_152 (O_152,N_8398,N_7902);
nor UO_153 (O_153,N_9268,N_8386);
and UO_154 (O_154,N_9277,N_7806);
and UO_155 (O_155,N_9216,N_9371);
and UO_156 (O_156,N_9323,N_8703);
nor UO_157 (O_157,N_9641,N_9141);
xor UO_158 (O_158,N_9633,N_9016);
nor UO_159 (O_159,N_9234,N_9703);
or UO_160 (O_160,N_9709,N_9568);
xnor UO_161 (O_161,N_9273,N_9003);
or UO_162 (O_162,N_8055,N_8137);
or UO_163 (O_163,N_9792,N_8957);
nand UO_164 (O_164,N_9784,N_9224);
xor UO_165 (O_165,N_7772,N_7670);
xor UO_166 (O_166,N_8254,N_8100);
or UO_167 (O_167,N_9721,N_8696);
nand UO_168 (O_168,N_9292,N_7861);
nand UO_169 (O_169,N_7888,N_9567);
nor UO_170 (O_170,N_7711,N_8298);
nor UO_171 (O_171,N_7825,N_8952);
xor UO_172 (O_172,N_8155,N_9806);
xor UO_173 (O_173,N_8477,N_7644);
nand UO_174 (O_174,N_9123,N_8534);
or UO_175 (O_175,N_7757,N_9822);
and UO_176 (O_176,N_7692,N_9649);
nand UO_177 (O_177,N_8788,N_9380);
and UO_178 (O_178,N_9899,N_7927);
and UO_179 (O_179,N_9827,N_9731);
nor UO_180 (O_180,N_9409,N_9113);
or UO_181 (O_181,N_8945,N_8627);
nand UO_182 (O_182,N_9465,N_8446);
nand UO_183 (O_183,N_8191,N_9168);
nor UO_184 (O_184,N_8991,N_8544);
xnor UO_185 (O_185,N_9689,N_8325);
xnor UO_186 (O_186,N_9848,N_9635);
and UO_187 (O_187,N_8979,N_9281);
and UO_188 (O_188,N_8582,N_8831);
and UO_189 (O_189,N_8944,N_9861);
nand UO_190 (O_190,N_9786,N_8120);
or UO_191 (O_191,N_9128,N_8781);
xor UO_192 (O_192,N_8363,N_8357);
nor UO_193 (O_193,N_9801,N_8165);
nand UO_194 (O_194,N_7508,N_8160);
nand UO_195 (O_195,N_9038,N_8927);
and UO_196 (O_196,N_8830,N_8545);
and UO_197 (O_197,N_9197,N_9066);
or UO_198 (O_198,N_8060,N_9129);
and UO_199 (O_199,N_8465,N_8714);
nor UO_200 (O_200,N_9550,N_8541);
or UO_201 (O_201,N_9261,N_8980);
nand UO_202 (O_202,N_9134,N_9961);
nor UO_203 (O_203,N_9930,N_9483);
nor UO_204 (O_204,N_9741,N_9411);
nor UO_205 (O_205,N_8271,N_8552);
nor UO_206 (O_206,N_9119,N_8810);
nor UO_207 (O_207,N_8053,N_9225);
nor UO_208 (O_208,N_8482,N_7891);
xor UO_209 (O_209,N_7769,N_7829);
nand UO_210 (O_210,N_9235,N_9585);
xor UO_211 (O_211,N_8189,N_7789);
xnor UO_212 (O_212,N_9714,N_9774);
or UO_213 (O_213,N_7737,N_9796);
nor UO_214 (O_214,N_9748,N_8523);
nand UO_215 (O_215,N_8321,N_7616);
xor UO_216 (O_216,N_8026,N_7914);
or UO_217 (O_217,N_7656,N_8042);
xor UO_218 (O_218,N_9684,N_8132);
nor UO_219 (O_219,N_9683,N_8108);
xor UO_220 (O_220,N_9753,N_7986);
or UO_221 (O_221,N_7778,N_7999);
and UO_222 (O_222,N_9884,N_7928);
or UO_223 (O_223,N_8276,N_9535);
xnor UO_224 (O_224,N_8700,N_9112);
xnor UO_225 (O_225,N_9795,N_9911);
nor UO_226 (O_226,N_8318,N_8772);
xnor UO_227 (O_227,N_8615,N_7591);
xor UO_228 (O_228,N_9817,N_7978);
xor UO_229 (O_229,N_9812,N_9425);
nand UO_230 (O_230,N_8390,N_7736);
xor UO_231 (O_231,N_9785,N_8525);
xor UO_232 (O_232,N_7702,N_8157);
nand UO_233 (O_233,N_9626,N_8756);
or UO_234 (O_234,N_8954,N_8777);
and UO_235 (O_235,N_8098,N_9576);
nor UO_236 (O_236,N_7731,N_7535);
nor UO_237 (O_237,N_9855,N_8392);
nand UO_238 (O_238,N_8074,N_8564);
nor UO_239 (O_239,N_8589,N_9400);
nor UO_240 (O_240,N_7796,N_9650);
nand UO_241 (O_241,N_7781,N_9645);
and UO_242 (O_242,N_8814,N_9605);
and UO_243 (O_243,N_7968,N_9945);
nand UO_244 (O_244,N_9843,N_7912);
and UO_245 (O_245,N_9609,N_9898);
nor UO_246 (O_246,N_9457,N_7552);
and UO_247 (O_247,N_9892,N_8193);
xnor UO_248 (O_248,N_9484,N_8009);
and UO_249 (O_249,N_9953,N_8535);
nor UO_250 (O_250,N_8766,N_9392);
xor UO_251 (O_251,N_9181,N_9433);
or UO_252 (O_252,N_9461,N_8470);
nor UO_253 (O_253,N_9333,N_9493);
or UO_254 (O_254,N_7609,N_9969);
and UO_255 (O_255,N_8983,N_8492);
nor UO_256 (O_256,N_9651,N_9106);
xor UO_257 (O_257,N_8826,N_9452);
and UO_258 (O_258,N_7983,N_8414);
nand UO_259 (O_259,N_9245,N_9551);
or UO_260 (O_260,N_8360,N_9826);
and UO_261 (O_261,N_9663,N_8516);
and UO_262 (O_262,N_7712,N_7558);
or UO_263 (O_263,N_8031,N_8763);
nand UO_264 (O_264,N_8602,N_8058);
and UO_265 (O_265,N_7991,N_8166);
nand UO_266 (O_266,N_8597,N_8295);
xor UO_267 (O_267,N_9690,N_8102);
nor UO_268 (O_268,N_9907,N_7507);
xnor UO_269 (O_269,N_7858,N_8761);
xnor UO_270 (O_270,N_8513,N_7766);
or UO_271 (O_271,N_7973,N_9091);
or UO_272 (O_272,N_8307,N_8843);
and UO_273 (O_273,N_7889,N_8168);
nand UO_274 (O_274,N_8237,N_9617);
nand UO_275 (O_275,N_7933,N_9354);
and UO_276 (O_276,N_8474,N_9638);
and UO_277 (O_277,N_8593,N_9236);
nand UO_278 (O_278,N_7943,N_9280);
and UO_279 (O_279,N_9184,N_9981);
and UO_280 (O_280,N_8982,N_9588);
xor UO_281 (O_281,N_8167,N_9109);
nor UO_282 (O_282,N_9086,N_9972);
nand UO_283 (O_283,N_9209,N_9327);
and UO_284 (O_284,N_9126,N_8664);
or UO_285 (O_285,N_9150,N_9422);
and UO_286 (O_286,N_7629,N_8421);
xor UO_287 (O_287,N_7564,N_8451);
or UO_288 (O_288,N_8351,N_8107);
nand UO_289 (O_289,N_9487,N_9230);
nand UO_290 (O_290,N_9910,N_7708);
xnor UO_291 (O_291,N_8480,N_7602);
nor UO_292 (O_292,N_9473,N_9231);
and UO_293 (O_293,N_9631,N_8119);
or UO_294 (O_294,N_7697,N_8384);
nand UO_295 (O_295,N_8299,N_9815);
nand UO_296 (O_296,N_8139,N_7980);
and UO_297 (O_297,N_8192,N_9221);
and UO_298 (O_298,N_9922,N_8901);
nand UO_299 (O_299,N_7897,N_8017);
xor UO_300 (O_300,N_8319,N_7718);
and UO_301 (O_301,N_7568,N_9919);
or UO_302 (O_302,N_9020,N_8648);
nor UO_303 (O_303,N_8280,N_8389);
xnor UO_304 (O_304,N_9693,N_9357);
or UO_305 (O_305,N_8837,N_8908);
nor UO_306 (O_306,N_8391,N_8289);
or UO_307 (O_307,N_8063,N_9833);
xor UO_308 (O_308,N_7625,N_9475);
nand UO_309 (O_309,N_9575,N_8479);
nor UO_310 (O_310,N_9139,N_8154);
nand UO_311 (O_311,N_8731,N_7622);
xnor UO_312 (O_312,N_8841,N_9681);
nor UO_313 (O_313,N_8618,N_8002);
xor UO_314 (O_314,N_7904,N_9862);
and UO_315 (O_315,N_9031,N_9740);
nor UO_316 (O_316,N_8655,N_8922);
nand UO_317 (O_317,N_8657,N_8041);
nand UO_318 (O_318,N_7959,N_7593);
xnor UO_319 (O_319,N_8818,N_8850);
and UO_320 (O_320,N_9111,N_9060);
or UO_321 (O_321,N_8116,N_8078);
nand UO_322 (O_322,N_9530,N_8247);
nand UO_323 (O_323,N_8676,N_9694);
nand UO_324 (O_324,N_9451,N_9571);
or UO_325 (O_325,N_9305,N_7803);
and UO_326 (O_326,N_8370,N_7585);
nand UO_327 (O_327,N_8997,N_8951);
nor UO_328 (O_328,N_8163,N_9569);
nand UO_329 (O_329,N_9625,N_9517);
and UO_330 (O_330,N_7865,N_7990);
xnor UO_331 (O_331,N_8976,N_7810);
and UO_332 (O_332,N_9180,N_7946);
nor UO_333 (O_333,N_7926,N_9828);
xor UO_334 (O_334,N_9199,N_8768);
and UO_335 (O_335,N_9799,N_8396);
nor UO_336 (O_336,N_8220,N_8216);
and UO_337 (O_337,N_7727,N_8955);
nor UO_338 (O_338,N_7759,N_8311);
nor UO_339 (O_339,N_9183,N_9980);
nor UO_340 (O_340,N_9201,N_9557);
xor UO_341 (O_341,N_7791,N_9104);
or UO_342 (O_342,N_8404,N_7971);
and UO_343 (O_343,N_7843,N_9987);
nor UO_344 (O_344,N_9434,N_8038);
nand UO_345 (O_345,N_9204,N_9037);
and UO_346 (O_346,N_7551,N_9591);
or UO_347 (O_347,N_7937,N_7726);
nand UO_348 (O_348,N_7715,N_8050);
nor UO_349 (O_349,N_9275,N_8054);
or UO_350 (O_350,N_8273,N_9272);
or UO_351 (O_351,N_8229,N_7835);
nor UO_352 (O_352,N_7667,N_8458);
nor UO_353 (O_353,N_7828,N_9103);
nand UO_354 (O_354,N_8015,N_7932);
nor UO_355 (O_355,N_7753,N_9124);
or UO_356 (O_356,N_7700,N_8358);
xor UO_357 (O_357,N_9355,N_8426);
and UO_358 (O_358,N_7634,N_8348);
xor UO_359 (O_359,N_8025,N_7890);
and UO_360 (O_360,N_8817,N_9726);
and UO_361 (O_361,N_9379,N_8684);
xor UO_362 (O_362,N_9873,N_8048);
and UO_363 (O_363,N_8967,N_9377);
and UO_364 (O_364,N_8324,N_8661);
xor UO_365 (O_365,N_8596,N_8913);
and UO_366 (O_366,N_9614,N_8747);
nand UO_367 (O_367,N_9927,N_7545);
nor UO_368 (O_368,N_9797,N_7741);
xor UO_369 (O_369,N_8653,N_7570);
and UO_370 (O_370,N_8775,N_7905);
or UO_371 (O_371,N_8865,N_8730);
nor UO_372 (O_372,N_9895,N_8505);
xor UO_373 (O_373,N_8999,N_8892);
and UO_374 (O_374,N_8151,N_8043);
nand UO_375 (O_375,N_9207,N_8981);
nand UO_376 (O_376,N_7915,N_8232);
xnor UO_377 (O_377,N_8087,N_9120);
or UO_378 (O_378,N_9814,N_9722);
and UO_379 (O_379,N_8932,N_8566);
nor UO_380 (O_380,N_9250,N_8340);
xor UO_381 (O_381,N_7841,N_9561);
and UO_382 (O_382,N_7870,N_7953);
nor UO_383 (O_383,N_8104,N_7921);
or UO_384 (O_384,N_9679,N_9064);
nand UO_385 (O_385,N_9140,N_8745);
and UO_386 (O_386,N_8561,N_7739);
xnor UO_387 (O_387,N_7838,N_9877);
nand UO_388 (O_388,N_9312,N_9361);
nand UO_389 (O_389,N_7962,N_8924);
nand UO_390 (O_390,N_8503,N_8428);
nor UO_391 (O_391,N_7651,N_7722);
nand UO_392 (O_392,N_9889,N_9583);
nor UO_393 (O_393,N_8947,N_7504);
xnor UO_394 (O_394,N_8287,N_7853);
and UO_395 (O_395,N_9198,N_8175);
nand UO_396 (O_396,N_9321,N_8239);
nor UO_397 (O_397,N_8840,N_8507);
nor UO_398 (O_398,N_7575,N_9763);
nor UO_399 (O_399,N_9659,N_9830);
or UO_400 (O_400,N_8278,N_9701);
and UO_401 (O_401,N_7658,N_8708);
or UO_402 (O_402,N_8963,N_9941);
nor UO_403 (O_403,N_8728,N_9915);
nor UO_404 (O_404,N_9364,N_9508);
and UO_405 (O_405,N_9787,N_7929);
or UO_406 (O_406,N_8614,N_7976);
nand UO_407 (O_407,N_8134,N_9931);
nand UO_408 (O_408,N_9604,N_8995);
and UO_409 (O_409,N_9378,N_8045);
and UO_410 (O_410,N_9202,N_8820);
or UO_411 (O_411,N_9023,N_9428);
nand UO_412 (O_412,N_8306,N_9559);
xnor UO_413 (O_413,N_9840,N_8996);
or UO_414 (O_414,N_9166,N_7779);
nand UO_415 (O_415,N_9908,N_8432);
or UO_416 (O_416,N_9570,N_9952);
or UO_417 (O_417,N_7909,N_7761);
nor UO_418 (O_418,N_7813,N_8591);
xor UO_419 (O_419,N_7530,N_7919);
and UO_420 (O_420,N_7957,N_8493);
and UO_421 (O_421,N_8242,N_8622);
and UO_422 (O_422,N_8005,N_8628);
or UO_423 (O_423,N_9929,N_8214);
xnor UO_424 (O_424,N_9300,N_8016);
or UO_425 (O_425,N_9586,N_8612);
and UO_426 (O_426,N_9213,N_8647);
or UO_427 (O_427,N_7820,N_8118);
nand UO_428 (O_428,N_9781,N_8904);
xor UO_429 (O_429,N_7689,N_9105);
and UO_430 (O_430,N_8091,N_9917);
or UO_431 (O_431,N_9427,N_9059);
or UO_432 (O_432,N_8133,N_9011);
nor UO_433 (O_433,N_9282,N_7846);
or UO_434 (O_434,N_7636,N_9418);
and UO_435 (O_435,N_9542,N_7750);
and UO_436 (O_436,N_8724,N_9170);
nor UO_437 (O_437,N_8604,N_8184);
nand UO_438 (O_438,N_9494,N_9990);
nor UO_439 (O_439,N_8172,N_9847);
nor UO_440 (O_440,N_8297,N_9013);
xnor UO_441 (O_441,N_9511,N_9851);
nor UO_442 (O_442,N_8586,N_8339);
or UO_443 (O_443,N_9610,N_8244);
nand UO_444 (O_444,N_8848,N_8308);
and UO_445 (O_445,N_8136,N_9358);
nor UO_446 (O_446,N_7874,N_9544);
or UO_447 (O_447,N_9519,N_8634);
nor UO_448 (O_448,N_9131,N_8842);
or UO_449 (O_449,N_9498,N_7855);
xor UO_450 (O_450,N_7541,N_7647);
nand UO_451 (O_451,N_8685,N_9802);
xor UO_452 (O_452,N_8067,N_8590);
xnor UO_453 (O_453,N_7967,N_8506);
or UO_454 (O_454,N_9222,N_7615);
and UO_455 (O_455,N_8181,N_8212);
nand UO_456 (O_456,N_9803,N_9432);
or UO_457 (O_457,N_7679,N_9030);
xnor UO_458 (O_458,N_8553,N_8066);
nor UO_459 (O_459,N_9039,N_8617);
or UO_460 (O_460,N_8742,N_8950);
or UO_461 (O_461,N_9986,N_8675);
nand UO_462 (O_462,N_7794,N_9668);
xor UO_463 (O_463,N_9442,N_9622);
or UO_464 (O_464,N_7676,N_8099);
and UO_465 (O_465,N_8910,N_7903);
and UO_466 (O_466,N_8517,N_7760);
xnor UO_467 (O_467,N_9725,N_9742);
and UO_468 (O_468,N_7966,N_8186);
or UO_469 (O_469,N_8977,N_8511);
nand UO_470 (O_470,N_7643,N_7804);
xnor UO_471 (O_471,N_9029,N_9791);
nor UO_472 (O_472,N_8419,N_8729);
or UO_473 (O_473,N_8519,N_9353);
xor UO_474 (O_474,N_7723,N_9329);
nor UO_475 (O_475,N_9291,N_8883);
xnor UO_476 (O_476,N_9769,N_7951);
and UO_477 (O_477,N_9708,N_7834);
nor UO_478 (O_478,N_9439,N_8262);
and UO_479 (O_479,N_9263,N_9677);
nand UO_480 (O_480,N_9497,N_8228);
and UO_481 (O_481,N_9276,N_8620);
nor UO_482 (O_482,N_7981,N_9652);
nand UO_483 (O_483,N_8679,N_9767);
and UO_484 (O_484,N_9351,N_7856);
nor UO_485 (O_485,N_9867,N_7566);
nor UO_486 (O_486,N_9186,N_8606);
xnor UO_487 (O_487,N_8037,N_9441);
nor UO_488 (O_488,N_9088,N_9459);
nand UO_489 (O_489,N_7538,N_8431);
nor UO_490 (O_490,N_7640,N_9868);
or UO_491 (O_491,N_7876,N_9553);
xor UO_492 (O_492,N_7540,N_8434);
and UO_493 (O_493,N_8029,N_9707);
xor UO_494 (O_494,N_8281,N_7785);
or UO_495 (O_495,N_9149,N_9240);
nand UO_496 (O_496,N_8430,N_7970);
or UO_497 (O_497,N_9151,N_8260);
xnor UO_498 (O_498,N_7567,N_8613);
or UO_499 (O_499,N_8476,N_9301);
nor UO_500 (O_500,N_9334,N_8514);
xor UO_501 (O_501,N_9607,N_9455);
xnor UO_502 (O_502,N_7886,N_8007);
or UO_503 (O_503,N_8824,N_8364);
xor UO_504 (O_504,N_7502,N_7808);
or UO_505 (O_505,N_8044,N_9682);
nand UO_506 (O_506,N_9807,N_7703);
nor UO_507 (O_507,N_8130,N_9860);
or UO_508 (O_508,N_8678,N_9482);
and UO_509 (O_509,N_9532,N_9925);
and UO_510 (O_510,N_8733,N_8206);
nor UO_511 (O_511,N_9022,N_9948);
nand UO_512 (O_512,N_8393,N_9114);
nor UO_513 (O_513,N_9079,N_9713);
nand UO_514 (O_514,N_9720,N_7742);
and UO_515 (O_515,N_8484,N_9623);
nor UO_516 (O_516,N_8556,N_8699);
or UO_517 (O_517,N_9369,N_9805);
and UO_518 (O_518,N_7604,N_9127);
xor UO_519 (O_519,N_8536,N_7956);
xor UO_520 (O_520,N_9778,N_7797);
or UO_521 (O_521,N_7767,N_7544);
and UO_522 (O_522,N_8473,N_7916);
nor UO_523 (O_523,N_8998,N_7503);
nand UO_524 (O_524,N_9759,N_9846);
and UO_525 (O_525,N_7580,N_8540);
and UO_526 (O_526,N_9082,N_8605);
or UO_527 (O_527,N_9440,N_8145);
nand UO_528 (O_528,N_8326,N_8366);
and UO_529 (O_529,N_9995,N_9252);
nor UO_530 (O_530,N_9574,N_8094);
nand UO_531 (O_531,N_8176,N_9971);
nand UO_532 (O_532,N_8320,N_7728);
nand UO_533 (O_533,N_9993,N_7994);
xor UO_534 (O_534,N_9964,N_9831);
or UO_535 (O_535,N_8086,N_9716);
nand UO_536 (O_536,N_8719,N_8375);
nor UO_537 (O_537,N_9172,N_8092);
or UO_538 (O_538,N_7522,N_7673);
nand UO_539 (O_539,N_8485,N_8483);
xnor UO_540 (O_540,N_8764,N_8491);
xnor UO_541 (O_541,N_8579,N_9335);
xnor UO_542 (O_542,N_9619,N_9678);
and UO_543 (O_543,N_8631,N_8328);
or UO_544 (O_544,N_7788,N_9620);
xor UO_545 (O_545,N_9777,N_8912);
or UO_546 (O_546,N_9156,N_8792);
xor UO_547 (O_547,N_8301,N_8857);
and UO_548 (O_548,N_8774,N_8797);
and UO_549 (O_549,N_8429,N_8626);
or UO_550 (O_550,N_7935,N_9918);
or UO_551 (O_551,N_8732,N_8692);
nor UO_552 (O_552,N_7589,N_9004);
and UO_553 (O_553,N_9158,N_9988);
xnor UO_554 (O_554,N_7938,N_7710);
or UO_555 (O_555,N_9025,N_8726);
xnor UO_556 (O_556,N_7832,N_9284);
and UO_557 (O_557,N_9841,N_7755);
xor UO_558 (O_558,N_9142,N_8401);
and UO_559 (O_559,N_9932,N_8362);
nand UO_560 (O_560,N_8970,N_9546);
nand UO_561 (O_561,N_9942,N_8501);
nand UO_562 (O_562,N_7885,N_8721);
nand UO_563 (O_563,N_7678,N_7506);
and UO_564 (O_564,N_8233,N_8587);
nand UO_565 (O_565,N_9920,N_7780);
or UO_566 (O_566,N_8852,N_9524);
or UO_567 (O_567,N_7985,N_8601);
nor UO_568 (O_568,N_8868,N_8658);
nand UO_569 (O_569,N_8638,N_9959);
and UO_570 (O_570,N_9429,N_9026);
nand UO_571 (O_571,N_8853,N_8891);
nand UO_572 (O_572,N_7941,N_9674);
nor UO_573 (O_573,N_9865,N_8464);
or UO_574 (O_574,N_8936,N_9144);
nor UO_575 (O_575,N_7992,N_8915);
nand UO_576 (O_576,N_9983,N_8013);
nand UO_577 (O_577,N_7539,N_9239);
and UO_578 (O_578,N_8697,N_7572);
and UO_579 (O_579,N_8070,N_8709);
nand UO_580 (O_580,N_8077,N_9259);
or UO_581 (O_581,N_8407,N_7515);
or UO_582 (O_582,N_8861,N_9478);
or UO_583 (O_583,N_7523,N_8855);
nor UO_584 (O_584,N_9154,N_7501);
xnor UO_585 (O_585,N_7592,N_9548);
nand UO_586 (O_586,N_7652,N_9049);
or UO_587 (O_587,N_8518,N_8274);
nor UO_588 (O_588,N_8866,N_8822);
nand UO_589 (O_589,N_8032,N_9220);
xor UO_590 (O_590,N_9687,N_8563);
xor UO_591 (O_591,N_9311,N_8867);
nand UO_592 (O_592,N_9600,N_9711);
nor UO_593 (O_593,N_8650,N_9406);
or UO_594 (O_594,N_8140,N_8113);
or UO_595 (O_595,N_9271,N_9776);
nor UO_596 (O_596,N_9515,N_8047);
xor UO_597 (O_597,N_9664,N_9019);
nand UO_598 (O_598,N_8224,N_8870);
nor UO_599 (O_599,N_7955,N_9671);
nand UO_600 (O_600,N_9704,N_8219);
nor UO_601 (O_601,N_8068,N_8028);
and UO_602 (O_602,N_9045,N_9021);
nor UO_603 (O_603,N_9161,N_8309);
nor UO_604 (O_604,N_9595,N_8813);
xnor UO_605 (O_605,N_7864,N_8410);
or UO_606 (O_606,N_9010,N_9938);
and UO_607 (O_607,N_7768,N_8975);
or UO_608 (O_608,N_7685,N_8882);
nand UO_609 (O_609,N_7849,N_8173);
or UO_610 (O_610,N_8382,N_9320);
or UO_611 (O_611,N_9458,N_8489);
or UO_612 (O_612,N_7691,N_8406);
nor UO_613 (O_613,N_7560,N_9839);
or UO_614 (O_614,N_8990,N_9470);
xnor UO_615 (O_615,N_8373,N_9886);
xor UO_616 (O_616,N_8105,N_7793);
nand UO_617 (O_617,N_8832,N_9325);
or UO_618 (O_618,N_7979,N_8021);
and UO_619 (O_619,N_8494,N_9522);
nor UO_620 (O_620,N_9116,N_7960);
nor UO_621 (O_621,N_9394,N_7635);
nand UO_622 (O_622,N_9093,N_7826);
and UO_623 (O_623,N_9613,N_8802);
and UO_624 (O_624,N_8899,N_8111);
xnor UO_625 (O_625,N_8368,N_9405);
nor UO_626 (O_626,N_8437,N_9627);
xor UO_627 (O_627,N_9653,N_8103);
or UO_628 (O_628,N_9590,N_8888);
nand UO_629 (O_629,N_9445,N_9710);
nor UO_630 (O_630,N_9761,N_8812);
or UO_631 (O_631,N_9842,N_9555);
nor UO_632 (O_632,N_8667,N_9780);
and UO_633 (O_633,N_9285,N_9307);
or UO_634 (O_634,N_9115,N_8420);
nand UO_635 (O_635,N_7562,N_9556);
and UO_636 (O_636,N_9770,N_8547);
or UO_637 (O_637,N_7725,N_7827);
and UO_638 (O_638,N_9177,N_8268);
nor UO_639 (O_639,N_9243,N_7939);
or UO_640 (O_640,N_8201,N_7677);
and UO_641 (O_641,N_8569,N_9363);
and UO_642 (O_642,N_7574,N_7945);
nor UO_643 (O_643,N_9396,N_7944);
xnor UO_644 (O_644,N_8958,N_8409);
nor UO_645 (O_645,N_9366,N_7873);
xor UO_646 (O_646,N_8666,N_9008);
xnor UO_647 (O_647,N_9476,N_8992);
and UO_648 (O_648,N_9464,N_8939);
nand UO_649 (O_649,N_7543,N_8024);
nand UO_650 (O_650,N_7917,N_9505);
nand UO_651 (O_651,N_8862,N_7668);
and UO_652 (O_652,N_9381,N_9738);
nor UO_653 (O_653,N_8203,N_8397);
or UO_654 (O_654,N_9996,N_7818);
and UO_655 (O_655,N_9593,N_9502);
nand UO_656 (O_656,N_7969,N_7798);
nand UO_657 (O_657,N_7989,N_7995);
xor UO_658 (O_658,N_9880,N_7925);
or UO_659 (O_659,N_9080,N_9523);
xor UO_660 (O_660,N_9352,N_8283);
and UO_661 (O_661,N_9310,N_9431);
nand UO_662 (O_662,N_8115,N_7631);
xor UO_663 (O_663,N_8478,N_8475);
nand UO_664 (O_664,N_9318,N_8199);
xor UO_665 (O_665,N_9989,N_7896);
xor UO_666 (O_666,N_7682,N_9266);
or UO_667 (O_667,N_8369,N_9666);
nor UO_668 (O_668,N_9420,N_8941);
nor UO_669 (O_669,N_7901,N_7687);
xnor UO_670 (O_670,N_7561,N_8616);
and UO_671 (O_671,N_7614,N_8422);
xor UO_672 (O_672,N_7573,N_9818);
or UO_673 (O_673,N_8875,N_8879);
xnor UO_674 (O_674,N_7654,N_7842);
or UO_675 (O_675,N_8205,N_8471);
and UO_676 (O_676,N_9153,N_8466);
or UO_677 (O_677,N_9504,N_8705);
nor UO_678 (O_678,N_8245,N_8942);
nor UO_679 (O_679,N_7920,N_7748);
xor UO_680 (O_680,N_8858,N_8023);
and UO_681 (O_681,N_8863,N_8093);
or UO_682 (O_682,N_8633,N_8827);
or UO_683 (O_683,N_9069,N_7586);
nand UO_684 (O_684,N_8076,N_8698);
nor UO_685 (O_685,N_7765,N_8290);
nor UO_686 (O_686,N_9376,N_8639);
and UO_687 (O_687,N_8127,N_9192);
nor UO_688 (O_688,N_8135,N_9727);
nor UO_689 (O_689,N_8836,N_8680);
nand UO_690 (O_690,N_8334,N_9488);
nor UO_691 (O_691,N_8323,N_7918);
and UO_692 (O_692,N_8218,N_9756);
nand UO_693 (O_693,N_7744,N_9477);
or UO_694 (O_694,N_9249,N_8011);
nand UO_695 (O_695,N_9423,N_9913);
and UO_696 (O_696,N_7930,N_9700);
xor UO_697 (O_697,N_9223,N_9095);
and UO_698 (O_698,N_7833,N_9028);
nand UO_699 (O_699,N_8416,N_9760);
nand UO_700 (O_700,N_8896,N_9287);
and UO_701 (O_701,N_8845,N_9415);
and UO_702 (O_702,N_9081,N_9552);
and UO_703 (O_703,N_8989,N_7510);
xnor UO_704 (O_704,N_8794,N_7675);
nor UO_705 (O_705,N_7735,N_8454);
or UO_706 (O_706,N_9940,N_9165);
or UO_707 (O_707,N_9863,N_9657);
or UO_708 (O_708,N_7972,N_9467);
xnor UO_709 (O_709,N_8909,N_9175);
or UO_710 (O_710,N_7659,N_8625);
and UO_711 (O_711,N_8660,N_8344);
or UO_712 (O_712,N_9316,N_7984);
nor UO_713 (O_713,N_9135,N_8110);
xor UO_714 (O_714,N_9044,N_9132);
nor UO_715 (O_715,N_9572,N_9251);
nor UO_716 (O_716,N_8327,N_9169);
or UO_717 (O_717,N_9946,N_9966);
and UO_718 (O_718,N_8550,N_7852);
and UO_719 (O_719,N_9949,N_9217);
nand UO_720 (O_720,N_8956,N_7517);
nor UO_721 (O_721,N_9829,N_8400);
or UO_722 (O_722,N_8121,N_9370);
xnor UO_723 (O_723,N_9054,N_7894);
nand UO_724 (O_724,N_8762,N_9869);
and UO_725 (O_725,N_9844,N_7578);
or UO_726 (O_726,N_9190,N_7840);
nand UO_727 (O_727,N_9226,N_8659);
or UO_728 (O_728,N_9187,N_9974);
nor UO_729 (O_729,N_9723,N_9654);
and UO_730 (O_730,N_8717,N_9870);
or UO_731 (O_731,N_8377,N_8986);
nor UO_732 (O_732,N_9669,N_8643);
or UO_733 (O_733,N_9043,N_8436);
nor UO_734 (O_734,N_8109,N_9036);
or UO_735 (O_735,N_7642,N_9834);
nor UO_736 (O_736,N_9118,N_8722);
nand UO_737 (O_737,N_8546,N_9962);
nor UO_738 (O_738,N_8972,N_8669);
nand UO_739 (O_739,N_8162,N_9500);
or UO_740 (O_740,N_8515,N_8849);
xor UO_741 (O_741,N_7590,N_9466);
nand UO_742 (O_742,N_9955,N_9728);
nor UO_743 (O_743,N_8816,N_7581);
nand UO_744 (O_744,N_7648,N_7860);
xnor UO_745 (O_745,N_9278,N_8677);
or UO_746 (O_746,N_7940,N_9258);
and UO_747 (O_747,N_9237,N_8710);
nor UO_748 (O_748,N_8294,N_8776);
nor UO_749 (O_749,N_8748,N_8502);
or UO_750 (O_750,N_8468,N_8522);
nand UO_751 (O_751,N_9436,N_9598);
xor UO_752 (O_752,N_8240,N_9382);
and UO_753 (O_753,N_8197,N_8549);
nand UO_754 (O_754,N_9762,N_9162);
nor UO_755 (O_755,N_9977,N_9138);
nor UO_756 (O_756,N_9185,N_9024);
xnor UO_757 (O_757,N_8906,N_8292);
or UO_758 (O_758,N_9463,N_9897);
nand UO_759 (O_759,N_7819,N_8275);
or UO_760 (O_760,N_8572,N_9348);
xnor UO_761 (O_761,N_8354,N_9730);
nor UO_762 (O_762,N_9472,N_8187);
and UO_763 (O_763,N_9794,N_9324);
nor UO_764 (O_764,N_9046,N_8415);
nand UO_765 (O_765,N_7563,N_8585);
nand UO_766 (O_766,N_9058,N_8651);
nand UO_767 (O_767,N_9110,N_9577);
xor UO_768 (O_768,N_8158,N_8238);
and UO_769 (O_769,N_8751,N_9592);
and UO_770 (O_770,N_7872,N_7548);
nor UO_771 (O_771,N_9705,N_9388);
and UO_772 (O_772,N_8259,N_8079);
xor UO_773 (O_773,N_9533,N_7850);
nand UO_774 (O_774,N_9691,N_7790);
nand UO_775 (O_775,N_7542,N_9850);
nand UO_776 (O_776,N_7863,N_8695);
and UO_777 (O_777,N_9540,N_7837);
xnor UO_778 (O_778,N_8226,N_8190);
nand UO_779 (O_779,N_8114,N_8467);
and UO_780 (O_780,N_9597,N_8805);
nand UO_781 (O_781,N_8565,N_7893);
or UO_782 (O_782,N_9014,N_7709);
nand UO_783 (O_783,N_9662,N_9580);
nor UO_784 (O_784,N_9083,N_9390);
and UO_785 (O_785,N_8182,N_8061);
xnor UO_786 (O_786,N_8153,N_9978);
xor UO_787 (O_787,N_8161,N_8894);
xor UO_788 (O_788,N_9041,N_8959);
nor UO_789 (O_789,N_9034,N_9998);
or UO_790 (O_790,N_9543,N_9735);
nand UO_791 (O_791,N_9208,N_9052);
and UO_792 (O_792,N_8177,N_7745);
or UO_793 (O_793,N_7655,N_9410);
xnor UO_794 (O_794,N_9302,N_8012);
xnor UO_795 (O_795,N_9256,N_7730);
nor UO_796 (O_796,N_7546,N_8159);
nor UO_797 (O_797,N_8767,N_8893);
xnor UO_798 (O_798,N_8331,N_9893);
and UO_799 (O_799,N_9751,N_8185);
nand UO_800 (O_800,N_9934,N_7892);
and UO_801 (O_801,N_9821,N_8928);
and UO_802 (O_802,N_9474,N_8917);
nand UO_803 (O_803,N_9073,N_9085);
xnor UO_804 (O_804,N_9937,N_7936);
nand UO_805 (O_805,N_7998,N_8341);
nor UO_806 (O_806,N_9636,N_8811);
or UO_807 (O_807,N_9800,N_7724);
or UO_808 (O_808,N_8138,N_8973);
or UO_809 (O_809,N_7537,N_8251);
xnor UO_810 (O_810,N_8723,N_9290);
nor UO_811 (O_811,N_9408,N_7961);
nand UO_812 (O_812,N_7868,N_9789);
or UO_813 (O_813,N_9349,N_8610);
nor UO_814 (O_814,N_7599,N_9935);
and UO_815 (O_815,N_8444,N_9339);
and UO_816 (O_816,N_8008,N_8623);
and UO_817 (O_817,N_9009,N_8757);
nor UO_818 (O_818,N_7582,N_8707);
nand UO_819 (O_819,N_8529,N_9783);
xnor UO_820 (O_820,N_9584,N_8921);
nand UO_821 (O_821,N_8884,N_9878);
and UO_822 (O_822,N_8234,N_8258);
or UO_823 (O_823,N_7569,N_8727);
nor UO_824 (O_824,N_9196,N_7800);
nand UO_825 (O_825,N_7924,N_9182);
or UO_826 (O_826,N_9210,N_8293);
xnor UO_827 (O_827,N_8886,N_8943);
nor UO_828 (O_828,N_8144,N_7680);
nand UO_829 (O_829,N_9823,N_8640);
and UO_830 (O_830,N_8753,N_9510);
and UO_831 (O_831,N_7695,N_9729);
and UO_832 (O_832,N_9212,N_7624);
nand UO_833 (O_833,N_7645,N_9675);
nand UO_834 (O_834,N_8964,N_8447);
and UO_835 (O_835,N_8088,N_9639);
xor UO_836 (O_836,N_8889,N_8035);
or UO_837 (O_837,N_7511,N_8770);
and UO_838 (O_838,N_8347,N_9896);
nor UO_839 (O_839,N_7694,N_8241);
or UO_840 (O_840,N_9885,N_7740);
nand UO_841 (O_841,N_8030,N_8823);
nor UO_842 (O_842,N_8551,N_8689);
nand UO_843 (O_843,N_9242,N_8594);
nand UO_844 (O_844,N_9107,N_9589);
nor UO_845 (O_845,N_8630,N_9773);
and UO_846 (O_846,N_9179,N_7815);
and UO_847 (O_847,N_9991,N_8887);
xnor UO_848 (O_848,N_9900,N_9538);
nand UO_849 (O_849,N_9328,N_9832);
nor UO_850 (O_850,N_9951,N_9067);
xor UO_851 (O_851,N_8412,N_8279);
nand UO_852 (O_852,N_8040,N_9737);
nor UO_853 (O_853,N_9070,N_9298);
xnor UO_854 (O_854,N_8734,N_8350);
nor UO_855 (O_855,N_9499,N_8785);
and UO_856 (O_856,N_9536,N_8417);
xor UO_857 (O_857,N_9176,N_7662);
and UO_858 (O_858,N_7713,N_8267);
xnor UO_859 (O_859,N_8263,N_9630);
xnor UO_860 (O_860,N_8272,N_7879);
nand UO_861 (O_861,N_9241,N_8588);
xor UO_862 (O_862,N_9734,N_7954);
or UO_863 (O_863,N_8799,N_7553);
xor UO_864 (O_864,N_9501,N_7965);
nor UO_865 (O_865,N_7633,N_8195);
nand UO_866 (O_866,N_9963,N_9365);
nor UO_867 (O_867,N_8800,N_9914);
and UO_868 (O_868,N_8652,N_9894);
xor UO_869 (O_869,N_8619,N_8567);
or UO_870 (O_870,N_8496,N_8914);
or UO_871 (O_871,N_9558,N_7526);
and UO_872 (O_872,N_9837,N_7660);
or UO_873 (O_873,N_7947,N_8152);
nor UO_874 (O_874,N_8411,N_9979);
xor UO_875 (O_875,N_7696,N_9816);
xnor UO_876 (O_876,N_8743,N_8056);
or UO_877 (O_877,N_7610,N_8284);
nand UO_878 (O_878,N_8577,N_9027);
xnor UO_879 (O_879,N_8568,N_8129);
nor UO_880 (O_880,N_9820,N_9076);
or UO_881 (O_881,N_9053,N_8371);
nand UO_882 (O_882,N_9033,N_8902);
nand UO_883 (O_883,N_9015,N_9766);
and UO_884 (O_884,N_7774,N_9960);
or UO_885 (O_885,N_7549,N_8338);
and UO_886 (O_886,N_9824,N_9326);
xor UO_887 (O_887,N_9507,N_7630);
and UO_888 (O_888,N_9874,N_8739);
nor UO_889 (O_889,N_7525,N_9304);
nand UO_890 (O_890,N_8253,N_7862);
xnor UO_891 (O_891,N_7669,N_8829);
nor UO_892 (O_892,N_9512,N_9383);
nor UO_893 (O_893,N_7812,N_8524);
nand UO_894 (O_894,N_8662,N_9094);
nor UO_895 (O_895,N_8688,N_8372);
nand UO_896 (O_896,N_8644,N_8408);
and UO_897 (O_897,N_8270,N_8296);
xor UO_898 (O_898,N_7688,N_7733);
and UO_899 (O_899,N_8595,N_9599);
and UO_900 (O_900,N_9191,N_7608);
nor UO_901 (O_901,N_8033,N_9143);
nand UO_902 (O_902,N_8790,N_9446);
xnor UO_903 (O_903,N_9750,N_7646);
and UO_904 (O_904,N_7674,N_9130);
nor UO_905 (O_905,N_9744,N_7882);
nor UO_906 (O_906,N_9811,N_9531);
or UO_907 (O_907,N_9566,N_8231);
and UO_908 (O_908,N_9621,N_9624);
nand UO_909 (O_909,N_8759,N_8286);
nor UO_910 (O_910,N_9994,N_7934);
or UO_911 (O_911,N_9537,N_8538);
xor UO_912 (O_912,N_8854,N_8427);
and UO_913 (O_913,N_8057,N_9443);
nand UO_914 (O_914,N_9984,N_8204);
nor UO_915 (O_915,N_9883,N_9976);
nand UO_916 (O_916,N_8629,N_8504);
and UO_917 (O_917,N_8463,N_9965);
nand UO_918 (O_918,N_9218,N_8907);
or UO_919 (O_919,N_9074,N_7975);
nand UO_920 (O_920,N_9283,N_8122);
or UO_921 (O_921,N_9001,N_7583);
xor UO_922 (O_922,N_7963,N_9975);
nand UO_923 (O_923,N_7716,N_9447);
or UO_924 (O_924,N_8112,N_8796);
nand UO_925 (O_925,N_8143,N_9928);
nor UO_926 (O_926,N_8183,N_9492);
or UO_927 (O_927,N_8346,N_8081);
xnor UO_928 (O_928,N_8971,N_8198);
or UO_929 (O_929,N_8196,N_9152);
nor UO_930 (O_930,N_8073,N_8609);
xor UO_931 (O_931,N_7847,N_8509);
nor UO_932 (O_932,N_9453,N_8938);
xor UO_933 (O_933,N_7977,N_7958);
nand UO_934 (O_934,N_9051,N_7641);
xor UO_935 (O_935,N_8929,N_7782);
nor UO_936 (O_936,N_8872,N_9854);
nor UO_937 (O_937,N_9876,N_8352);
nor UO_938 (O_938,N_8528,N_9100);
nand UO_939 (O_939,N_7529,N_8715);
xnor UO_940 (O_940,N_7617,N_9875);
xor UO_941 (O_941,N_8209,N_9206);
and UO_942 (O_942,N_9048,N_9102);
nor UO_943 (O_943,N_8018,N_8096);
xnor UO_944 (O_944,N_9528,N_9350);
and UO_945 (O_945,N_7650,N_9999);
or UO_946 (O_946,N_8065,N_8071);
nand UO_947 (O_947,N_9262,N_9640);
nand UO_948 (O_948,N_9122,N_8673);
or UO_949 (O_949,N_8285,N_9012);
nand UO_950 (O_950,N_8900,N_9146);
nand UO_951 (O_951,N_8693,N_7884);
and UO_952 (O_952,N_7653,N_7601);
xor UO_953 (O_953,N_9057,N_8844);
nand UO_954 (O_954,N_8332,N_9970);
or UO_955 (O_955,N_8225,N_8082);
nand UO_956 (O_956,N_8808,N_8988);
nor UO_957 (O_957,N_9958,N_8300);
or UO_958 (O_958,N_8559,N_9688);
nand UO_959 (O_959,N_9188,N_7557);
nand UO_960 (O_960,N_7887,N_8828);
nor UO_961 (O_961,N_9189,N_9468);
xnor UO_962 (O_962,N_8725,N_8903);
or UO_963 (O_963,N_9634,N_8291);
and UO_964 (O_964,N_7556,N_8984);
nand UO_965 (O_965,N_9315,N_9098);
or UO_966 (O_966,N_9503,N_9173);
and UO_967 (O_967,N_8472,N_8488);
xnor UO_968 (O_968,N_8001,N_8250);
nand UO_969 (O_969,N_7579,N_9758);
xor UO_970 (O_970,N_7786,N_9890);
xor UO_971 (O_971,N_9905,N_9078);
or UO_972 (O_972,N_9346,N_8949);
nor UO_973 (O_973,N_9362,N_8890);
nand UO_974 (O_974,N_9793,N_8637);
xor UO_975 (O_975,N_9228,N_9838);
nor UO_976 (O_976,N_9643,N_9279);
xnor UO_977 (O_977,N_7814,N_8142);
nand UO_978 (O_978,N_9332,N_7520);
xnor UO_979 (O_979,N_9075,N_9909);
or UO_980 (O_980,N_7859,N_9404);
nand UO_981 (O_981,N_9849,N_8083);
nor UO_982 (O_982,N_9121,N_8211);
nand UO_983 (O_983,N_7597,N_8310);
nor UO_984 (O_984,N_9950,N_9772);
xor UO_985 (O_985,N_7952,N_9338);
xnor UO_986 (O_986,N_8330,N_8170);
xor UO_987 (O_987,N_8317,N_9211);
nand UO_988 (O_988,N_9717,N_7802);
xnor UO_989 (O_989,N_8786,N_8608);
xnor UO_990 (O_990,N_9089,N_8940);
nor UO_991 (O_991,N_9092,N_9926);
and UO_992 (O_992,N_8019,N_7721);
xnor UO_993 (O_993,N_8531,N_7512);
or UO_994 (O_994,N_9340,N_8315);
and UO_995 (O_995,N_8213,N_8453);
nand UO_996 (O_996,N_9071,N_7611);
xnor UO_997 (O_997,N_8780,N_8150);
and UO_998 (O_998,N_7777,N_8449);
xor UO_999 (O_999,N_9485,N_8499);
xor UO_1000 (O_1000,N_7875,N_9424);
or UO_1001 (O_1001,N_9903,N_9696);
nand UO_1002 (O_1002,N_8895,N_8642);
nor UO_1003 (O_1003,N_7784,N_8754);
nor UO_1004 (O_1004,N_8571,N_9628);
nor UO_1005 (O_1005,N_9399,N_9412);
and UO_1006 (O_1006,N_8539,N_7824);
xnor UO_1007 (O_1007,N_8542,N_8993);
nor UO_1008 (O_1008,N_7756,N_9344);
xor UO_1009 (O_1009,N_8322,N_9881);
and UO_1010 (O_1010,N_9345,N_7707);
nand UO_1011 (O_1011,N_8825,N_8686);
and UO_1012 (O_1012,N_9264,N_7822);
or UO_1013 (O_1013,N_9386,N_8969);
nand UO_1014 (O_1014,N_7505,N_8581);
nand UO_1015 (O_1015,N_7949,N_9247);
nor UO_1016 (O_1016,N_9403,N_8968);
nor UO_1017 (O_1017,N_9393,N_9061);
or UO_1018 (O_1018,N_8526,N_9936);
nand UO_1019 (O_1019,N_8869,N_7729);
or UO_1020 (O_1020,N_8455,N_8690);
xnor UO_1021 (O_1021,N_8399,N_9655);
xor UO_1022 (O_1022,N_9319,N_8312);
and UO_1023 (O_1023,N_9063,N_8672);
and UO_1024 (O_1024,N_7997,N_7587);
nand UO_1025 (O_1025,N_9539,N_8834);
or UO_1026 (O_1026,N_9065,N_8918);
and UO_1027 (O_1027,N_8469,N_9454);
nand UO_1028 (O_1028,N_8881,N_7738);
xor UO_1029 (O_1029,N_7974,N_8510);
nor UO_1030 (O_1030,N_9047,N_8445);
xor UO_1031 (O_1031,N_9866,N_8156);
xor UO_1032 (O_1032,N_8450,N_9097);
nor UO_1033 (O_1033,N_8878,N_7871);
xnor UO_1034 (O_1034,N_9509,N_8442);
or UO_1035 (O_1035,N_8575,N_9656);
and UO_1036 (O_1036,N_7771,N_9857);
or UO_1037 (O_1037,N_9194,N_8885);
or UO_1038 (O_1038,N_8755,N_9018);
nor UO_1039 (O_1039,N_8769,N_9331);
nor UO_1040 (O_1040,N_8741,N_8919);
nand UO_1041 (O_1041,N_7839,N_9944);
xor UO_1042 (O_1042,N_9660,N_8815);
and UO_1043 (O_1043,N_9603,N_9872);
xor UO_1044 (O_1044,N_8558,N_8926);
nand UO_1045 (O_1045,N_7743,N_9342);
nand UO_1046 (O_1046,N_9602,N_7720);
nand UO_1047 (O_1047,N_8227,N_8385);
and UO_1048 (O_1048,N_8335,N_7684);
xnor UO_1049 (O_1049,N_8355,N_9771);
nand UO_1050 (O_1050,N_9125,N_8064);
nor UO_1051 (O_1051,N_9385,N_9858);
xor UO_1052 (O_1052,N_7681,N_9486);
xnor UO_1053 (O_1053,N_9471,N_9481);
nor UO_1054 (O_1054,N_9615,N_7848);
and UO_1055 (O_1055,N_9308,N_8578);
nor UO_1056 (O_1056,N_7783,N_7686);
or UO_1057 (O_1057,N_9670,N_8188);
nor UO_1058 (O_1058,N_8795,N_8148);
xnor UO_1059 (O_1059,N_9163,N_9087);
xor UO_1060 (O_1060,N_9809,N_8933);
nand UO_1061 (O_1061,N_9968,N_8208);
and UO_1062 (O_1062,N_9673,N_9871);
nand UO_1063 (O_1063,N_9573,N_8486);
nand UO_1064 (O_1064,N_7705,N_9768);
xnor UO_1065 (O_1065,N_9227,N_7751);
and UO_1066 (O_1066,N_8750,N_9437);
or UO_1067 (O_1067,N_9313,N_9887);
nand UO_1068 (O_1068,N_8694,N_9395);
xnor UO_1069 (O_1069,N_8383,N_8527);
nand UO_1070 (O_1070,N_9565,N_8394);
nor UO_1071 (O_1071,N_8737,N_8302);
or UO_1072 (O_1072,N_9541,N_7513);
or UO_1073 (O_1073,N_8758,N_9062);
xnor UO_1074 (O_1074,N_9719,N_9265);
nor UO_1075 (O_1075,N_8570,N_8749);
or UO_1076 (O_1076,N_8873,N_9686);
nor UO_1077 (O_1077,N_8665,N_9676);
xnor UO_1078 (O_1078,N_8533,N_8543);
and UO_1079 (O_1079,N_7527,N_8560);
nor UO_1080 (O_1080,N_9755,N_9096);
nand UO_1081 (O_1081,N_9912,N_7867);
and UO_1082 (O_1082,N_8646,N_9916);
or UO_1083 (O_1083,N_8603,N_8530);
nor UO_1084 (O_1084,N_8946,N_8217);
xnor UO_1085 (O_1085,N_8378,N_9072);
nor UO_1086 (O_1086,N_7516,N_7627);
and UO_1087 (O_1087,N_8706,N_8288);
nand UO_1088 (O_1088,N_8269,N_8223);
or UO_1089 (O_1089,N_7795,N_7898);
xor UO_1090 (O_1090,N_8987,N_7787);
and UO_1091 (O_1091,N_8418,N_9665);
or UO_1092 (O_1092,N_8336,N_8978);
or UO_1093 (O_1093,N_8931,N_9982);
and UO_1094 (O_1094,N_7851,N_8847);
nand UO_1095 (O_1095,N_8106,N_9520);
xnor UO_1096 (O_1096,N_7533,N_9219);
or UO_1097 (O_1097,N_9367,N_9171);
nor UO_1098 (O_1098,N_8961,N_8674);
nand UO_1099 (O_1099,N_9973,N_9314);
and UO_1100 (O_1100,N_9294,N_9117);
nor UO_1101 (O_1101,N_9554,N_9341);
or UO_1102 (O_1102,N_7706,N_9939);
nor UO_1103 (O_1103,N_8171,N_9397);
and UO_1104 (O_1104,N_8835,N_9859);
or UO_1105 (O_1105,N_8180,N_8598);
xor UO_1106 (O_1106,N_7559,N_9924);
and UO_1107 (O_1107,N_7869,N_7519);
nand UO_1108 (O_1108,N_9148,N_7931);
and UO_1109 (O_1109,N_8876,N_8405);
nand UO_1110 (O_1110,N_9337,N_7524);
and UO_1111 (O_1111,N_8498,N_9155);
nand UO_1112 (O_1112,N_9646,N_7603);
and UO_1113 (O_1113,N_8246,N_8495);
nor UO_1114 (O_1114,N_8937,N_9752);
or UO_1115 (O_1115,N_8663,N_9810);
or UO_1116 (O_1116,N_8039,N_9435);
nor UO_1117 (O_1117,N_7605,N_7993);
or UO_1118 (O_1118,N_9384,N_9289);
nor UO_1119 (O_1119,N_9992,N_7908);
nand UO_1120 (O_1120,N_9214,N_8027);
xnor UO_1121 (O_1121,N_8554,N_9564);
nand UO_1122 (O_1122,N_7987,N_8819);
nand UO_1123 (O_1123,N_9368,N_8020);
and UO_1124 (O_1124,N_8798,N_9947);
xor UO_1125 (O_1125,N_7618,N_7752);
or UO_1126 (O_1126,N_9322,N_9270);
xnor UO_1127 (O_1127,N_7831,N_8860);
and UO_1128 (O_1128,N_9448,N_9336);
xnor UO_1129 (O_1129,N_7588,N_7878);
and UO_1130 (O_1130,N_8966,N_8147);
and UO_1131 (O_1131,N_9902,N_8803);
nand UO_1132 (O_1132,N_8036,N_8920);
nand UO_1133 (O_1133,N_8207,N_8349);
nand UO_1134 (O_1134,N_8911,N_9257);
and UO_1135 (O_1135,N_7554,N_7899);
and UO_1136 (O_1136,N_7661,N_8221);
or UO_1137 (O_1137,N_7612,N_8313);
xor UO_1138 (O_1138,N_8413,N_9606);
nor UO_1139 (O_1139,N_9375,N_9819);
or UO_1140 (O_1140,N_7555,N_8520);
nand UO_1141 (O_1141,N_9933,N_8923);
and UO_1142 (O_1142,N_9526,N_9347);
or UO_1143 (O_1143,N_8452,N_8934);
xor UO_1144 (O_1144,N_7534,N_9685);
nand UO_1145 (O_1145,N_8838,N_7628);
and UO_1146 (O_1146,N_9195,N_9882);
and UO_1147 (O_1147,N_8402,N_9419);
nor UO_1148 (O_1148,N_7719,N_9407);
and UO_1149 (O_1149,N_9527,N_8117);
or UO_1150 (O_1150,N_8718,N_8953);
nand UO_1151 (O_1151,N_9921,N_8583);
nor UO_1152 (O_1152,N_9997,N_7844);
nor UO_1153 (O_1153,N_8752,N_9563);
nand UO_1154 (O_1154,N_9356,N_8256);
and UO_1155 (O_1155,N_9040,N_8000);
or UO_1156 (O_1156,N_9480,N_8782);
or UO_1157 (O_1157,N_8178,N_9518);
nand UO_1158 (O_1158,N_9957,N_9414);
or UO_1159 (O_1159,N_9904,N_8681);
and UO_1160 (O_1160,N_7776,N_9495);
nor UO_1161 (O_1161,N_7900,N_9469);
and UO_1162 (O_1162,N_9032,N_9157);
nand UO_1163 (O_1163,N_9229,N_9746);
xnor UO_1164 (O_1164,N_7532,N_7816);
nor UO_1165 (O_1165,N_9525,N_9372);
or UO_1166 (O_1166,N_9391,N_9238);
xor UO_1167 (O_1167,N_8611,N_8806);
or UO_1168 (O_1168,N_9056,N_9648);
nand UO_1169 (O_1169,N_9782,N_9808);
xnor UO_1170 (O_1170,N_9601,N_8874);
and UO_1171 (O_1171,N_7521,N_8194);
nor UO_1172 (O_1172,N_9836,N_8600);
or UO_1173 (O_1173,N_8974,N_9042);
or UO_1174 (O_1174,N_8425,N_7699);
or UO_1175 (O_1175,N_8343,N_9514);
nor UO_1176 (O_1176,N_8051,N_8353);
and UO_1177 (O_1177,N_8379,N_8793);
xnor UO_1178 (O_1178,N_9521,N_8671);
nand UO_1179 (O_1179,N_9444,N_8783);
and UO_1180 (O_1180,N_8097,N_8236);
nor UO_1181 (O_1181,N_8871,N_9813);
or UO_1182 (O_1182,N_9203,N_9513);
xor UO_1183 (O_1183,N_7996,N_8859);
or UO_1184 (O_1184,N_9260,N_8599);
and UO_1185 (O_1185,N_9233,N_9779);
xor UO_1186 (O_1186,N_8645,N_8101);
and UO_1187 (O_1187,N_7950,N_8668);
xor UO_1188 (O_1188,N_8439,N_9389);
or UO_1189 (O_1189,N_9137,N_9712);
and UO_1190 (O_1190,N_8164,N_8356);
nand UO_1191 (O_1191,N_8846,N_8361);
or UO_1192 (O_1192,N_8773,N_7638);
nor UO_1193 (O_1193,N_7746,N_8210);
xnor UO_1194 (O_1194,N_8202,N_9462);
and UO_1195 (O_1195,N_7911,N_8034);
and UO_1196 (O_1196,N_8022,N_9667);
nand UO_1197 (O_1197,N_9629,N_9611);
and UO_1198 (O_1198,N_8779,N_8255);
nor UO_1199 (O_1199,N_9954,N_7857);
nor UO_1200 (O_1200,N_9402,N_8252);
xor UO_1201 (O_1201,N_7942,N_7528);
nand UO_1202 (O_1202,N_9888,N_7910);
nor UO_1203 (O_1203,N_9490,N_8089);
nand UO_1204 (O_1204,N_7948,N_8123);
nand UO_1205 (O_1205,N_9644,N_8146);
or UO_1206 (O_1206,N_7536,N_8880);
and UO_1207 (O_1207,N_7619,N_8481);
xor UO_1208 (O_1208,N_8898,N_9923);
and UO_1209 (O_1209,N_7792,N_8049);
or UO_1210 (O_1210,N_8654,N_8555);
or UO_1211 (O_1211,N_9145,N_8621);
or UO_1212 (O_1212,N_9101,N_7907);
nand UO_1213 (O_1213,N_9017,N_9050);
and UO_1214 (O_1214,N_8257,N_9343);
nor UO_1215 (O_1215,N_8443,N_8635);
or UO_1216 (O_1216,N_9943,N_9864);
xnor UO_1217 (O_1217,N_8965,N_9413);
and UO_1218 (O_1218,N_9159,N_9906);
nand UO_1219 (O_1219,N_9296,N_9754);
or UO_1220 (O_1220,N_7531,N_9232);
and UO_1221 (O_1221,N_9401,N_8720);
nor UO_1222 (O_1222,N_7717,N_7571);
xor UO_1223 (O_1223,N_8740,N_9547);
nand UO_1224 (O_1224,N_8380,N_9594);
and UO_1225 (O_1225,N_8557,N_7770);
and UO_1226 (O_1226,N_9430,N_8632);
nor UO_1227 (O_1227,N_8249,N_9373);
or UO_1228 (O_1228,N_7672,N_9330);
nor UO_1229 (O_1229,N_8821,N_7883);
and UO_1230 (O_1230,N_7600,N_9642);
or UO_1231 (O_1231,N_9529,N_9035);
xnor UO_1232 (O_1232,N_7845,N_9743);
and UO_1233 (O_1233,N_8851,N_8856);
xor UO_1234 (O_1234,N_8711,N_7866);
xnor UO_1235 (O_1235,N_8169,N_7799);
and UO_1236 (O_1236,N_7732,N_7754);
and UO_1237 (O_1237,N_8072,N_9647);
nor UO_1238 (O_1238,N_9587,N_7764);
and UO_1239 (O_1239,N_8985,N_9804);
nor UO_1240 (O_1240,N_9416,N_7657);
nor UO_1241 (O_1241,N_8230,N_8716);
or UO_1242 (O_1242,N_8433,N_9306);
nor UO_1243 (O_1243,N_9967,N_9680);
xnor UO_1244 (O_1244,N_8329,N_8771);
xnor UO_1245 (O_1245,N_7690,N_9136);
nand UO_1246 (O_1246,N_9309,N_8010);
nand UO_1247 (O_1247,N_9317,N_9578);
and UO_1248 (O_1248,N_7714,N_9417);
nor UO_1249 (O_1249,N_8576,N_9632);
nand UO_1250 (O_1250,N_9941,N_8586);
nor UO_1251 (O_1251,N_9073,N_7873);
nor UO_1252 (O_1252,N_9438,N_9069);
or UO_1253 (O_1253,N_8428,N_8408);
nor UO_1254 (O_1254,N_9037,N_7630);
nor UO_1255 (O_1255,N_9504,N_8294);
or UO_1256 (O_1256,N_8195,N_9776);
and UO_1257 (O_1257,N_9731,N_8480);
nand UO_1258 (O_1258,N_8655,N_7512);
xor UO_1259 (O_1259,N_8941,N_9865);
and UO_1260 (O_1260,N_9563,N_8415);
or UO_1261 (O_1261,N_7514,N_9325);
nor UO_1262 (O_1262,N_9775,N_8426);
nand UO_1263 (O_1263,N_9258,N_8740);
or UO_1264 (O_1264,N_8292,N_9347);
nand UO_1265 (O_1265,N_7779,N_9211);
and UO_1266 (O_1266,N_9901,N_7960);
or UO_1267 (O_1267,N_8103,N_7933);
or UO_1268 (O_1268,N_9219,N_7760);
nand UO_1269 (O_1269,N_8301,N_9721);
nor UO_1270 (O_1270,N_8770,N_9739);
nand UO_1271 (O_1271,N_9241,N_8132);
or UO_1272 (O_1272,N_7742,N_9739);
nor UO_1273 (O_1273,N_8502,N_8432);
nor UO_1274 (O_1274,N_8505,N_8627);
nand UO_1275 (O_1275,N_9398,N_9363);
nand UO_1276 (O_1276,N_8747,N_9025);
nand UO_1277 (O_1277,N_8266,N_9810);
or UO_1278 (O_1278,N_8251,N_7708);
or UO_1279 (O_1279,N_8245,N_9406);
xnor UO_1280 (O_1280,N_8602,N_8890);
and UO_1281 (O_1281,N_7806,N_9539);
xor UO_1282 (O_1282,N_9088,N_7634);
nor UO_1283 (O_1283,N_9154,N_7519);
nor UO_1284 (O_1284,N_9417,N_9149);
and UO_1285 (O_1285,N_9892,N_9910);
xnor UO_1286 (O_1286,N_9202,N_8338);
xor UO_1287 (O_1287,N_8137,N_8977);
nor UO_1288 (O_1288,N_9978,N_7676);
nand UO_1289 (O_1289,N_7590,N_7735);
xor UO_1290 (O_1290,N_8440,N_8346);
nor UO_1291 (O_1291,N_9207,N_8731);
or UO_1292 (O_1292,N_8450,N_8733);
and UO_1293 (O_1293,N_7814,N_7856);
nand UO_1294 (O_1294,N_8176,N_8944);
nor UO_1295 (O_1295,N_7512,N_9205);
or UO_1296 (O_1296,N_8764,N_8003);
xnor UO_1297 (O_1297,N_8487,N_8827);
and UO_1298 (O_1298,N_7516,N_7942);
xnor UO_1299 (O_1299,N_8166,N_7764);
nor UO_1300 (O_1300,N_9032,N_7584);
nor UO_1301 (O_1301,N_9463,N_8657);
or UO_1302 (O_1302,N_8970,N_7815);
xor UO_1303 (O_1303,N_9653,N_9788);
or UO_1304 (O_1304,N_8340,N_9764);
nand UO_1305 (O_1305,N_8991,N_9814);
xor UO_1306 (O_1306,N_9228,N_9769);
nand UO_1307 (O_1307,N_8992,N_9624);
xnor UO_1308 (O_1308,N_9651,N_9025);
and UO_1309 (O_1309,N_8413,N_9297);
xor UO_1310 (O_1310,N_7885,N_8062);
and UO_1311 (O_1311,N_9635,N_9250);
xnor UO_1312 (O_1312,N_8051,N_8390);
nor UO_1313 (O_1313,N_7518,N_7514);
or UO_1314 (O_1314,N_8881,N_7633);
nand UO_1315 (O_1315,N_9690,N_8409);
nand UO_1316 (O_1316,N_7906,N_7674);
nor UO_1317 (O_1317,N_9924,N_9585);
nand UO_1318 (O_1318,N_7546,N_8898);
and UO_1319 (O_1319,N_8658,N_7563);
and UO_1320 (O_1320,N_9355,N_9746);
nor UO_1321 (O_1321,N_7705,N_9673);
and UO_1322 (O_1322,N_9284,N_8540);
nand UO_1323 (O_1323,N_9334,N_9197);
nor UO_1324 (O_1324,N_8792,N_9936);
nor UO_1325 (O_1325,N_8781,N_7645);
or UO_1326 (O_1326,N_9668,N_9601);
and UO_1327 (O_1327,N_7867,N_9038);
or UO_1328 (O_1328,N_8031,N_9816);
nor UO_1329 (O_1329,N_9806,N_8341);
and UO_1330 (O_1330,N_8286,N_8243);
nand UO_1331 (O_1331,N_9717,N_9776);
nand UO_1332 (O_1332,N_9662,N_8402);
xor UO_1333 (O_1333,N_7854,N_7902);
xor UO_1334 (O_1334,N_7789,N_9494);
xnor UO_1335 (O_1335,N_7777,N_9089);
and UO_1336 (O_1336,N_8499,N_8630);
nor UO_1337 (O_1337,N_7549,N_8927);
nand UO_1338 (O_1338,N_8069,N_9507);
nand UO_1339 (O_1339,N_7777,N_7700);
and UO_1340 (O_1340,N_9075,N_8610);
or UO_1341 (O_1341,N_9562,N_7650);
or UO_1342 (O_1342,N_8912,N_9658);
or UO_1343 (O_1343,N_9301,N_7835);
xnor UO_1344 (O_1344,N_9711,N_7859);
and UO_1345 (O_1345,N_7845,N_9929);
or UO_1346 (O_1346,N_9187,N_9423);
or UO_1347 (O_1347,N_9107,N_7567);
nand UO_1348 (O_1348,N_7545,N_9859);
or UO_1349 (O_1349,N_8297,N_7726);
or UO_1350 (O_1350,N_7616,N_9305);
and UO_1351 (O_1351,N_8967,N_8464);
nand UO_1352 (O_1352,N_8474,N_7966);
nand UO_1353 (O_1353,N_9128,N_7549);
nor UO_1354 (O_1354,N_7877,N_8098);
nor UO_1355 (O_1355,N_8083,N_9264);
and UO_1356 (O_1356,N_8118,N_8259);
xor UO_1357 (O_1357,N_8848,N_8042);
nor UO_1358 (O_1358,N_9678,N_7632);
nand UO_1359 (O_1359,N_8058,N_8020);
nor UO_1360 (O_1360,N_8440,N_8301);
nand UO_1361 (O_1361,N_9845,N_9721);
and UO_1362 (O_1362,N_9728,N_9161);
nor UO_1363 (O_1363,N_7793,N_7579);
nand UO_1364 (O_1364,N_7902,N_9741);
nor UO_1365 (O_1365,N_9187,N_7566);
and UO_1366 (O_1366,N_9405,N_8518);
xnor UO_1367 (O_1367,N_9903,N_7622);
xnor UO_1368 (O_1368,N_8823,N_8059);
nor UO_1369 (O_1369,N_9792,N_8636);
nand UO_1370 (O_1370,N_9671,N_8143);
nor UO_1371 (O_1371,N_7754,N_8650);
nor UO_1372 (O_1372,N_7897,N_8802);
or UO_1373 (O_1373,N_8024,N_8639);
xor UO_1374 (O_1374,N_7870,N_8993);
nand UO_1375 (O_1375,N_8870,N_8587);
and UO_1376 (O_1376,N_9474,N_8143);
nor UO_1377 (O_1377,N_7573,N_8559);
and UO_1378 (O_1378,N_7566,N_7558);
nor UO_1379 (O_1379,N_9494,N_8128);
nor UO_1380 (O_1380,N_9344,N_9862);
nand UO_1381 (O_1381,N_9059,N_9804);
nand UO_1382 (O_1382,N_8057,N_9804);
nor UO_1383 (O_1383,N_9258,N_9472);
and UO_1384 (O_1384,N_9161,N_7755);
nand UO_1385 (O_1385,N_8764,N_8999);
nor UO_1386 (O_1386,N_9427,N_8970);
nor UO_1387 (O_1387,N_8738,N_9999);
xor UO_1388 (O_1388,N_8400,N_7856);
and UO_1389 (O_1389,N_7738,N_7899);
xor UO_1390 (O_1390,N_7645,N_8489);
and UO_1391 (O_1391,N_9494,N_9641);
nand UO_1392 (O_1392,N_8331,N_9334);
nor UO_1393 (O_1393,N_7936,N_9256);
xnor UO_1394 (O_1394,N_9193,N_7525);
and UO_1395 (O_1395,N_9096,N_7707);
nand UO_1396 (O_1396,N_8685,N_8662);
xor UO_1397 (O_1397,N_7652,N_7707);
and UO_1398 (O_1398,N_8800,N_7773);
or UO_1399 (O_1399,N_7647,N_8634);
xnor UO_1400 (O_1400,N_7883,N_9322);
or UO_1401 (O_1401,N_9214,N_7701);
xnor UO_1402 (O_1402,N_9817,N_9398);
nand UO_1403 (O_1403,N_9585,N_9199);
nor UO_1404 (O_1404,N_7988,N_8750);
nor UO_1405 (O_1405,N_8518,N_8516);
xor UO_1406 (O_1406,N_7577,N_7820);
or UO_1407 (O_1407,N_8895,N_9419);
nand UO_1408 (O_1408,N_8618,N_9962);
nor UO_1409 (O_1409,N_7559,N_8977);
xnor UO_1410 (O_1410,N_8526,N_8380);
nand UO_1411 (O_1411,N_7832,N_9176);
xor UO_1412 (O_1412,N_8233,N_9848);
nor UO_1413 (O_1413,N_9568,N_8593);
xnor UO_1414 (O_1414,N_9396,N_7839);
and UO_1415 (O_1415,N_8386,N_8706);
nand UO_1416 (O_1416,N_8927,N_7865);
and UO_1417 (O_1417,N_7518,N_8124);
nor UO_1418 (O_1418,N_9095,N_8143);
nand UO_1419 (O_1419,N_8365,N_9637);
or UO_1420 (O_1420,N_9909,N_7630);
and UO_1421 (O_1421,N_8201,N_9866);
nor UO_1422 (O_1422,N_9019,N_8318);
or UO_1423 (O_1423,N_9994,N_7576);
or UO_1424 (O_1424,N_9058,N_7826);
xnor UO_1425 (O_1425,N_8253,N_8145);
and UO_1426 (O_1426,N_8323,N_9220);
xnor UO_1427 (O_1427,N_7516,N_9350);
xnor UO_1428 (O_1428,N_9215,N_9342);
and UO_1429 (O_1429,N_8843,N_8750);
xor UO_1430 (O_1430,N_8531,N_9435);
and UO_1431 (O_1431,N_8488,N_8344);
xnor UO_1432 (O_1432,N_9224,N_9658);
nor UO_1433 (O_1433,N_8373,N_7702);
or UO_1434 (O_1434,N_9659,N_8918);
xor UO_1435 (O_1435,N_9148,N_9133);
or UO_1436 (O_1436,N_7962,N_9937);
and UO_1437 (O_1437,N_9409,N_7847);
nor UO_1438 (O_1438,N_8157,N_8266);
nor UO_1439 (O_1439,N_8200,N_9472);
nor UO_1440 (O_1440,N_8835,N_8296);
nand UO_1441 (O_1441,N_9766,N_8146);
nand UO_1442 (O_1442,N_9744,N_8973);
and UO_1443 (O_1443,N_9070,N_7544);
nand UO_1444 (O_1444,N_7740,N_8451);
and UO_1445 (O_1445,N_8053,N_8246);
xor UO_1446 (O_1446,N_9867,N_9923);
or UO_1447 (O_1447,N_7996,N_9949);
nor UO_1448 (O_1448,N_7750,N_9097);
nor UO_1449 (O_1449,N_8764,N_9434);
nor UO_1450 (O_1450,N_8132,N_7622);
nand UO_1451 (O_1451,N_9779,N_8803);
nand UO_1452 (O_1452,N_9491,N_8858);
or UO_1453 (O_1453,N_9132,N_7556);
nand UO_1454 (O_1454,N_7738,N_8188);
nor UO_1455 (O_1455,N_9690,N_8305);
and UO_1456 (O_1456,N_9766,N_8497);
or UO_1457 (O_1457,N_8304,N_8757);
xnor UO_1458 (O_1458,N_9755,N_8785);
nor UO_1459 (O_1459,N_8709,N_8780);
xor UO_1460 (O_1460,N_8899,N_9411);
and UO_1461 (O_1461,N_9172,N_8863);
nor UO_1462 (O_1462,N_8078,N_8976);
and UO_1463 (O_1463,N_8469,N_7650);
nand UO_1464 (O_1464,N_8238,N_9904);
and UO_1465 (O_1465,N_8276,N_8430);
or UO_1466 (O_1466,N_7789,N_8034);
xor UO_1467 (O_1467,N_9181,N_9629);
and UO_1468 (O_1468,N_9802,N_7534);
and UO_1469 (O_1469,N_9972,N_8592);
and UO_1470 (O_1470,N_7520,N_9183);
nand UO_1471 (O_1471,N_8184,N_9168);
or UO_1472 (O_1472,N_8396,N_8924);
xnor UO_1473 (O_1473,N_8360,N_9470);
xor UO_1474 (O_1474,N_7591,N_9076);
nand UO_1475 (O_1475,N_9874,N_9178);
and UO_1476 (O_1476,N_8181,N_7662);
xor UO_1477 (O_1477,N_8209,N_9299);
nor UO_1478 (O_1478,N_8545,N_8426);
nand UO_1479 (O_1479,N_9856,N_8763);
xnor UO_1480 (O_1480,N_9044,N_7905);
xnor UO_1481 (O_1481,N_8704,N_8685);
nor UO_1482 (O_1482,N_7757,N_9865);
and UO_1483 (O_1483,N_7721,N_8233);
xnor UO_1484 (O_1484,N_7781,N_9873);
nand UO_1485 (O_1485,N_9473,N_9342);
nor UO_1486 (O_1486,N_7727,N_8232);
nand UO_1487 (O_1487,N_8660,N_9153);
and UO_1488 (O_1488,N_7965,N_8045);
nand UO_1489 (O_1489,N_8551,N_8647);
or UO_1490 (O_1490,N_7637,N_7669);
nand UO_1491 (O_1491,N_9158,N_9617);
and UO_1492 (O_1492,N_9672,N_8858);
xnor UO_1493 (O_1493,N_8028,N_9115);
and UO_1494 (O_1494,N_9351,N_9849);
nand UO_1495 (O_1495,N_7949,N_8220);
or UO_1496 (O_1496,N_7720,N_8757);
xor UO_1497 (O_1497,N_9784,N_9200);
or UO_1498 (O_1498,N_8077,N_9685);
and UO_1499 (O_1499,N_8565,N_8654);
endmodule