module basic_5000_50000_5000_10_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nand U0 (N_0,In_25,In_1101);
nor U1 (N_1,In_2588,In_4145);
nand U2 (N_2,In_4577,In_1044);
nor U3 (N_3,In_1442,In_4879);
or U4 (N_4,In_3882,In_1857);
nand U5 (N_5,In_4380,In_2323);
nand U6 (N_6,In_33,In_1320);
and U7 (N_7,In_1169,In_1740);
nand U8 (N_8,In_565,In_3674);
and U9 (N_9,In_3770,In_1623);
xor U10 (N_10,In_2015,In_1591);
nor U11 (N_11,In_3205,In_1855);
and U12 (N_12,In_2358,In_2395);
or U13 (N_13,In_3255,In_800);
and U14 (N_14,In_2642,In_2888);
nand U15 (N_15,In_75,In_2553);
and U16 (N_16,In_4221,In_2992);
or U17 (N_17,In_3667,In_876);
xnor U18 (N_18,In_4764,In_3656);
nor U19 (N_19,In_3813,In_534);
nand U20 (N_20,In_4456,In_4773);
and U21 (N_21,In_1722,In_689);
nand U22 (N_22,In_4056,In_3727);
xor U23 (N_23,In_30,In_20);
nand U24 (N_24,In_2089,In_1231);
nor U25 (N_25,In_922,In_222);
nor U26 (N_26,In_2177,In_4003);
nor U27 (N_27,In_2394,In_974);
nand U28 (N_28,In_4935,In_697);
nor U29 (N_29,In_2523,In_2643);
and U30 (N_30,In_2105,In_2499);
nand U31 (N_31,In_4703,In_103);
and U32 (N_32,In_4360,In_446);
nor U33 (N_33,In_2220,In_3897);
or U34 (N_34,In_3764,In_3757);
or U35 (N_35,In_1967,In_1802);
and U36 (N_36,In_2117,In_4967);
nand U37 (N_37,In_1684,In_3990);
and U38 (N_38,In_2272,In_2939);
and U39 (N_39,In_1352,In_1912);
xnor U40 (N_40,In_4678,In_2620);
nor U41 (N_41,In_3288,In_2974);
and U42 (N_42,In_2330,In_4851);
nand U43 (N_43,In_4763,In_3438);
and U44 (N_44,In_2245,In_2614);
nand U45 (N_45,In_3215,In_2839);
nand U46 (N_46,In_2243,In_1055);
nor U47 (N_47,In_3901,In_4511);
or U48 (N_48,In_3352,In_588);
or U49 (N_49,In_2862,In_3407);
nor U50 (N_50,In_2900,In_246);
nor U51 (N_51,In_351,In_2185);
nand U52 (N_52,In_4154,In_3361);
or U53 (N_53,In_4979,In_293);
nor U54 (N_54,In_3156,In_1200);
xnor U55 (N_55,In_2752,In_4923);
and U56 (N_56,In_3341,In_2537);
nand U57 (N_57,In_741,In_616);
nand U58 (N_58,In_4447,In_100);
or U59 (N_59,In_587,In_2647);
xnor U60 (N_60,In_2759,In_2656);
and U61 (N_61,In_723,In_3179);
nand U62 (N_62,In_1037,In_1970);
and U63 (N_63,In_2476,In_521);
nand U64 (N_64,In_4120,In_3745);
nand U65 (N_65,In_4589,In_4059);
nor U66 (N_66,In_4322,In_952);
xnor U67 (N_67,In_1248,In_2035);
or U68 (N_68,In_2118,In_2281);
xnor U69 (N_69,In_2670,In_1581);
nor U70 (N_70,In_4884,In_3340);
nor U71 (N_71,In_2590,In_2836);
nor U72 (N_72,In_3768,In_1412);
xnor U73 (N_73,In_4585,In_2750);
nor U74 (N_74,In_1693,In_4378);
nand U75 (N_75,In_2819,In_4581);
and U76 (N_76,In_1256,In_4917);
and U77 (N_77,In_1923,In_4445);
nand U78 (N_78,In_474,In_776);
or U79 (N_79,In_4252,In_1506);
nor U80 (N_80,In_16,In_462);
nand U81 (N_81,In_992,In_1666);
xnor U82 (N_82,In_963,In_3685);
nor U83 (N_83,In_2041,In_1141);
xor U84 (N_84,In_3710,In_3636);
and U85 (N_85,In_178,In_607);
nand U86 (N_86,In_4153,In_2705);
nor U87 (N_87,In_903,In_4093);
and U88 (N_88,In_3962,In_2183);
nand U89 (N_89,In_865,In_2333);
nor U90 (N_90,In_1495,In_2026);
nand U91 (N_91,In_327,In_4098);
and U92 (N_92,In_850,In_4115);
nor U93 (N_93,In_1307,In_816);
nand U94 (N_94,In_1113,In_3647);
nor U95 (N_95,In_3848,In_1709);
nor U96 (N_96,In_4213,In_4474);
and U97 (N_97,In_2916,In_1992);
and U98 (N_98,In_3084,In_4076);
nand U99 (N_99,In_2389,In_2192);
nand U100 (N_100,In_3322,In_4468);
nor U101 (N_101,In_887,In_606);
or U102 (N_102,In_4391,In_2547);
nand U103 (N_103,In_433,In_104);
nor U104 (N_104,In_495,In_1456);
nor U105 (N_105,In_806,In_4743);
nor U106 (N_106,In_35,In_86);
nor U107 (N_107,In_1767,In_333);
or U108 (N_108,In_3476,In_3478);
or U109 (N_109,In_3890,In_2515);
nor U110 (N_110,In_2188,In_2033);
xor U111 (N_111,In_1136,In_4049);
or U112 (N_112,In_2132,In_4858);
nand U113 (N_113,In_4926,In_255);
nand U114 (N_114,In_853,In_1370);
and U115 (N_115,In_182,In_114);
nor U116 (N_116,In_1462,In_2677);
and U117 (N_117,In_4205,In_2881);
nand U118 (N_118,In_634,In_3113);
nand U119 (N_119,In_4455,In_3171);
nand U120 (N_120,In_3226,In_4625);
and U121 (N_121,In_1934,In_4035);
nor U122 (N_122,In_4290,In_2227);
or U123 (N_123,In_2686,In_3256);
xor U124 (N_124,In_3716,In_3465);
nor U125 (N_125,In_2849,In_4509);
and U126 (N_126,In_1409,In_1651);
nand U127 (N_127,In_4730,In_2594);
xnor U128 (N_128,In_4044,In_2599);
nor U129 (N_129,In_3872,In_2372);
nand U130 (N_130,In_113,In_2887);
and U131 (N_131,In_595,In_4141);
nand U132 (N_132,In_1478,In_4948);
nand U133 (N_133,In_2497,In_3860);
and U134 (N_134,In_4195,In_190);
and U135 (N_135,In_2167,In_1368);
nand U136 (N_136,In_301,In_3999);
and U137 (N_137,In_1217,In_4641);
nor U138 (N_138,In_1800,In_3431);
and U139 (N_139,In_1833,In_4092);
and U140 (N_140,In_3167,In_4578);
or U141 (N_141,In_986,In_4868);
nand U142 (N_142,In_3106,In_2271);
and U143 (N_143,In_73,In_2926);
xnor U144 (N_144,In_1510,In_1030);
or U145 (N_145,In_3974,In_413);
nand U146 (N_146,In_2469,In_4435);
or U147 (N_147,In_2287,In_3114);
nor U148 (N_148,In_4862,In_747);
and U149 (N_149,In_4083,In_620);
nor U150 (N_150,In_2332,In_1156);
or U151 (N_151,In_2601,In_4089);
nor U152 (N_152,In_3027,In_200);
or U153 (N_153,In_2247,In_356);
nor U154 (N_154,In_664,In_4551);
and U155 (N_155,In_1405,In_3212);
and U156 (N_156,In_2181,In_716);
and U157 (N_157,In_757,In_684);
and U158 (N_158,In_4159,In_3249);
and U159 (N_159,In_1790,In_2827);
nand U160 (N_160,In_4684,In_624);
xor U161 (N_161,In_4466,In_4579);
or U162 (N_162,In_3376,In_4584);
xnor U163 (N_163,In_3096,In_4876);
and U164 (N_164,In_774,In_2139);
nor U165 (N_165,In_3837,In_2291);
and U166 (N_166,In_1218,In_3581);
nor U167 (N_167,In_1836,In_2712);
or U168 (N_168,In_1877,In_2756);
and U169 (N_169,In_2847,In_694);
or U170 (N_170,In_766,In_3323);
or U171 (N_171,In_4515,In_4355);
and U172 (N_172,In_528,In_1189);
nand U173 (N_173,In_3912,In_4042);
nand U174 (N_174,In_4530,In_3511);
or U175 (N_175,In_3827,In_2918);
or U176 (N_176,In_1897,In_4898);
xor U177 (N_177,In_2725,In_2096);
nor U178 (N_178,In_1521,In_2978);
nand U179 (N_179,In_242,In_3992);
or U180 (N_180,In_4800,In_2025);
and U181 (N_181,In_1016,In_3499);
nor U182 (N_182,In_1702,In_3540);
xor U183 (N_183,In_4889,In_947);
or U184 (N_184,In_2806,In_3895);
or U185 (N_185,In_2904,In_532);
or U186 (N_186,In_3326,In_1057);
xnor U187 (N_187,In_203,In_2619);
xnor U188 (N_188,In_3842,In_3738);
xnor U189 (N_189,In_323,In_7);
or U190 (N_190,In_4314,In_4254);
xnor U191 (N_191,In_2492,In_2267);
nand U192 (N_192,In_1783,In_3053);
nor U193 (N_193,In_1332,In_1282);
nand U194 (N_194,In_3362,In_1237);
nor U195 (N_195,In_744,In_3316);
or U196 (N_196,In_4971,In_4993);
nor U197 (N_197,In_526,In_2006);
nand U198 (N_198,In_4497,In_3169);
nor U199 (N_199,In_2844,In_2010);
and U200 (N_200,In_2152,In_4528);
nand U201 (N_201,In_4552,In_463);
nand U202 (N_202,In_1007,In_4178);
and U203 (N_203,In_3535,In_171);
and U204 (N_204,In_1508,In_3480);
or U205 (N_205,In_514,In_4163);
or U206 (N_206,In_2023,In_4481);
xnor U207 (N_207,In_4111,In_2415);
or U208 (N_208,In_4257,In_4925);
and U209 (N_209,In_1979,In_3408);
nand U210 (N_210,In_4675,In_938);
and U211 (N_211,In_2316,In_556);
or U212 (N_212,In_4592,In_983);
nor U213 (N_213,In_321,In_1348);
and U214 (N_214,In_3708,In_782);
nor U215 (N_215,In_2814,In_995);
nor U216 (N_216,In_2997,In_2279);
nand U217 (N_217,In_1496,In_2748);
and U218 (N_218,In_3858,In_1664);
or U219 (N_219,In_3088,In_1536);
or U220 (N_220,In_3730,In_2283);
nor U221 (N_221,In_575,In_2371);
and U222 (N_222,In_1394,In_2954);
nor U223 (N_223,In_4021,In_2672);
xnor U224 (N_224,In_3285,In_1885);
xor U225 (N_225,In_1959,In_2445);
and U226 (N_226,In_2095,In_921);
and U227 (N_227,In_205,In_3485);
nand U228 (N_228,In_2674,In_3204);
and U229 (N_229,In_2576,In_3268);
nor U230 (N_230,In_2509,In_3449);
nor U231 (N_231,In_506,In_3909);
or U232 (N_232,In_3589,In_4693);
or U233 (N_233,In_2928,In_2561);
and U234 (N_234,In_4636,In_4704);
nand U235 (N_235,In_4335,In_3217);
nor U236 (N_236,In_2713,In_955);
nor U237 (N_237,In_2606,In_1406);
nand U238 (N_238,In_1077,In_3039);
or U239 (N_239,In_2650,In_1728);
or U240 (N_240,In_3903,In_3756);
and U241 (N_241,In_1955,In_2083);
and U242 (N_242,In_4458,In_2593);
nand U243 (N_243,In_4787,In_803);
nor U244 (N_244,In_430,In_4866);
and U245 (N_245,In_954,In_4157);
or U246 (N_246,In_303,In_4104);
and U247 (N_247,In_4751,In_2150);
or U248 (N_248,In_2193,In_1056);
nand U249 (N_249,In_1619,In_655);
nand U250 (N_250,In_1339,In_4177);
xnor U251 (N_251,In_1595,In_4526);
nand U252 (N_252,In_1918,In_623);
or U253 (N_253,In_1115,In_4038);
or U254 (N_254,In_2976,In_3759);
nand U255 (N_255,In_4150,In_1854);
nand U256 (N_256,In_4962,In_3261);
and U257 (N_257,In_1514,In_3594);
nor U258 (N_258,In_2305,In_4223);
and U259 (N_259,In_2443,In_3128);
nor U260 (N_260,In_4399,In_3926);
xnor U261 (N_261,In_1608,In_3963);
xnor U262 (N_262,In_2176,In_3307);
nor U263 (N_263,In_2482,In_4306);
or U264 (N_264,In_4087,In_3120);
nor U265 (N_265,In_263,In_2716);
nand U266 (N_266,In_4231,In_2453);
nor U267 (N_267,In_552,In_567);
nor U268 (N_268,In_789,In_346);
or U269 (N_269,In_2094,In_2514);
xnor U270 (N_270,In_4544,In_3082);
xor U271 (N_271,In_1816,In_1289);
and U272 (N_272,In_2765,In_1924);
nor U273 (N_273,In_1050,In_810);
nor U274 (N_274,In_4311,In_3512);
nand U275 (N_275,In_1299,In_4268);
or U276 (N_276,In_571,In_4521);
nand U277 (N_277,In_3464,In_594);
nand U278 (N_278,In_1054,In_2584);
nor U279 (N_279,In_4886,In_507);
nand U280 (N_280,In_4132,In_4953);
nand U281 (N_281,In_4988,In_754);
and U282 (N_282,In_2334,In_4016);
nor U283 (N_283,In_2504,In_2373);
xor U284 (N_284,In_404,In_2696);
nor U285 (N_285,In_2815,In_4700);
xnor U286 (N_286,In_3717,In_2627);
nor U287 (N_287,In_4464,In_2400);
and U288 (N_288,In_54,In_972);
and U289 (N_289,In_3871,In_1484);
and U290 (N_290,In_3467,In_2479);
nor U291 (N_291,In_1525,In_4325);
nand U292 (N_292,In_4756,In_4989);
nor U293 (N_293,In_2860,In_3771);
and U294 (N_294,In_1603,In_2161);
nand U295 (N_295,In_2983,In_1759);
nand U296 (N_296,In_2922,In_4346);
and U297 (N_297,In_1383,In_3552);
nand U298 (N_298,In_4845,In_1911);
and U299 (N_299,In_4643,In_968);
nor U300 (N_300,In_1397,In_1474);
or U301 (N_301,In_2222,In_470);
xnor U302 (N_302,In_2800,In_3908);
and U303 (N_303,In_4742,In_3705);
or U304 (N_304,In_913,In_1365);
and U305 (N_305,In_72,In_3418);
nand U306 (N_306,In_1734,In_4749);
or U307 (N_307,In_2551,In_4631);
or U308 (N_308,In_4976,In_3928);
or U309 (N_309,In_885,In_527);
or U310 (N_310,In_4187,In_3373);
nor U311 (N_311,In_3211,In_3331);
nor U312 (N_312,In_4614,In_4940);
nor U313 (N_313,In_306,In_3339);
xnor U314 (N_314,In_4672,In_603);
nor U315 (N_315,In_2409,In_408);
nand U316 (N_316,In_3392,In_1517);
nor U317 (N_317,In_1028,In_671);
nor U318 (N_318,In_183,In_1909);
or U319 (N_319,In_1308,In_258);
or U320 (N_320,In_4258,In_1275);
nor U321 (N_321,In_2496,In_317);
or U322 (N_322,In_918,In_4011);
nor U323 (N_323,In_1434,In_331);
nand U324 (N_324,In_3722,In_2592);
or U325 (N_325,In_4739,In_2254);
or U326 (N_326,In_1989,In_1481);
nor U327 (N_327,In_4379,In_2940);
nor U328 (N_328,In_329,In_287);
and U329 (N_329,In_3295,In_4433);
nand U330 (N_330,In_4333,In_4102);
nand U331 (N_331,In_718,In_1433);
xor U332 (N_332,In_4808,In_2336);
nor U333 (N_333,In_3777,In_1888);
nor U334 (N_334,In_4710,In_3593);
and U335 (N_335,In_4320,In_345);
nor U336 (N_336,In_1605,In_4899);
nor U337 (N_337,In_748,In_310);
and U338 (N_338,In_488,In_2159);
nor U339 (N_339,In_1703,In_259);
nor U340 (N_340,In_2019,In_1825);
or U341 (N_341,In_3976,In_4780);
or U342 (N_342,In_3763,In_4356);
nor U343 (N_343,In_1554,In_792);
nand U344 (N_344,In_4376,In_3134);
nand U345 (N_345,In_4431,In_1229);
nor U346 (N_346,In_3784,In_612);
nor U347 (N_347,In_3429,In_27);
or U348 (N_348,In_4279,In_2968);
nor U349 (N_349,In_4189,In_2513);
and U350 (N_350,In_557,In_3124);
or U351 (N_351,In_2345,In_4927);
and U352 (N_352,In_358,In_4226);
or U353 (N_353,In_3490,In_825);
nand U354 (N_354,In_2113,In_221);
nor U355 (N_355,In_217,In_4383);
and U356 (N_356,In_959,In_4519);
or U357 (N_357,In_1944,In_883);
nor U358 (N_358,In_896,In_1827);
and U359 (N_359,In_3216,In_2869);
or U360 (N_360,In_964,In_3917);
nand U361 (N_361,In_3208,In_3196);
nand U362 (N_362,In_1475,In_1931);
nand U363 (N_363,In_237,In_949);
nand U364 (N_364,In_906,In_2544);
and U365 (N_365,In_2003,In_1920);
or U366 (N_366,In_4538,In_4911);
nand U367 (N_367,In_1815,In_4357);
and U368 (N_368,In_2277,In_2249);
and U369 (N_369,In_3437,In_3733);
or U370 (N_370,In_1534,In_350);
nand U371 (N_371,In_2246,In_861);
nand U372 (N_372,In_3247,In_3282);
or U373 (N_373,In_3781,In_3849);
xor U374 (N_374,In_1502,In_2374);
and U375 (N_375,In_1636,In_4545);
nand U376 (N_376,In_4348,In_3422);
and U377 (N_377,In_2407,In_3083);
nand U378 (N_378,In_2299,In_3330);
nor U379 (N_379,In_4687,In_2856);
and U380 (N_380,In_551,In_4449);
or U381 (N_381,In_4135,In_4492);
nor U382 (N_382,In_988,In_236);
nand U383 (N_383,In_3371,In_119);
nor U384 (N_384,In_2726,In_984);
xnor U385 (N_385,In_1158,In_251);
or U386 (N_386,In_1874,In_4305);
xnor U387 (N_387,In_475,In_2166);
nor U388 (N_388,In_1257,In_2558);
nor U389 (N_389,In_406,In_3989);
and U390 (N_390,In_3670,In_4754);
and U391 (N_391,In_733,In_1606);
and U392 (N_392,In_2196,In_132);
nor U393 (N_393,In_3328,In_3309);
nand U394 (N_394,In_3075,In_4733);
and U395 (N_395,In_617,In_1467);
nand U396 (N_396,In_4653,In_1135);
nor U397 (N_397,In_2956,In_2131);
and U398 (N_398,In_529,In_4487);
nand U399 (N_399,In_4156,In_3633);
nand U400 (N_400,In_3740,In_2195);
nand U401 (N_401,In_1476,In_2895);
and U402 (N_402,In_480,In_1807);
or U403 (N_403,In_875,In_1696);
or U404 (N_404,In_586,In_3752);
or U405 (N_405,In_3380,In_4740);
xnor U406 (N_406,In_759,In_2424);
nor U407 (N_407,In_1327,In_4827);
and U408 (N_408,In_2425,In_543);
or U409 (N_409,In_4164,In_2431);
or U410 (N_410,In_2045,In_1260);
xor U411 (N_411,In_1335,In_767);
or U412 (N_412,In_1657,In_3704);
or U413 (N_413,In_1343,In_1376);
and U414 (N_414,In_4611,In_2802);
xnor U415 (N_415,In_3206,In_4478);
or U416 (N_416,In_3946,In_4676);
xor U417 (N_417,In_1389,In_1809);
nor U418 (N_418,In_3095,In_4280);
or U419 (N_419,In_636,In_3676);
nor U420 (N_420,In_1498,In_711);
nor U421 (N_421,In_4339,In_3673);
or U422 (N_422,In_688,In_4473);
and U423 (N_423,In_1744,In_2794);
xor U424 (N_424,In_699,In_4639);
nand U425 (N_425,In_518,In_2318);
and U426 (N_426,In_1949,In_666);
nand U427 (N_427,In_3152,In_1139);
xor U428 (N_428,In_169,In_2327);
and U429 (N_429,In_2893,In_1901);
nand U430 (N_430,In_4599,In_1147);
nor U431 (N_431,In_4591,In_1691);
nand U432 (N_432,In_38,In_715);
or U433 (N_433,In_1943,In_1259);
nor U434 (N_434,In_2224,In_2434);
or U435 (N_435,In_4313,In_1234);
xor U436 (N_436,In_1298,In_3627);
nor U437 (N_437,In_1494,In_2321);
xnor U438 (N_438,In_197,In_281);
or U439 (N_439,In_4186,In_1860);
xor U440 (N_440,In_3808,In_4843);
nand U441 (N_441,In_31,In_3462);
nand U442 (N_442,In_3719,In_2457);
nor U443 (N_443,In_3644,In_3875);
xnor U444 (N_444,In_3229,In_2353);
xor U445 (N_445,In_2823,In_418);
xor U446 (N_446,In_3679,In_564);
or U447 (N_447,In_1176,In_1133);
nor U448 (N_448,In_669,In_2259);
nor U449 (N_449,In_1617,In_3130);
nand U450 (N_450,In_597,In_1239);
nor U451 (N_451,In_2863,In_4029);
nor U452 (N_452,In_3142,In_4662);
or U453 (N_453,In_3898,In_173);
or U454 (N_454,In_878,In_3358);
and U455 (N_455,In_1680,In_1822);
and U456 (N_456,In_873,In_1798);
and U457 (N_457,In_3811,In_3273);
and U458 (N_458,In_3894,In_212);
or U459 (N_459,In_3718,In_34);
nand U460 (N_460,In_1648,In_1527);
nor U461 (N_461,In_1839,In_3393);
and U462 (N_462,In_821,In_3655);
or U463 (N_463,In_2760,In_2543);
nand U464 (N_464,In_1123,In_1326);
or U465 (N_465,In_1177,In_277);
nor U466 (N_466,In_4941,In_4727);
nor U467 (N_467,In_3172,In_1919);
or U468 (N_468,In_2528,In_2265);
nor U469 (N_469,In_3213,In_1889);
and U470 (N_470,In_1817,In_1227);
nand U471 (N_471,In_2986,In_4161);
or U472 (N_472,In_3582,In_1199);
nor U473 (N_473,In_4185,In_3961);
nor U474 (N_474,In_3631,In_3042);
and U475 (N_475,In_1639,In_1408);
nor U476 (N_476,In_4908,In_2737);
and U477 (N_477,In_3109,In_1473);
xor U478 (N_478,In_892,In_3420);
nand U479 (N_479,In_884,In_77);
nor U480 (N_480,In_308,In_1160);
or U481 (N_481,In_1029,In_4426);
nand U482 (N_482,In_3365,In_2683);
and U483 (N_483,In_2158,In_4882);
nor U484 (N_484,In_3048,In_4437);
and U485 (N_485,In_1183,In_4785);
nor U486 (N_486,In_4783,In_1220);
and U487 (N_487,In_1721,In_2142);
nor U488 (N_488,In_4615,In_3214);
and U489 (N_489,In_2987,In_2664);
nor U490 (N_490,In_3641,In_2396);
nand U491 (N_491,In_1203,In_1454);
nor U492 (N_492,In_1678,In_1196);
and U493 (N_493,In_2116,In_2600);
xor U494 (N_494,In_4351,In_3528);
or U495 (N_495,In_1228,In_36);
nor U496 (N_496,In_4462,In_3866);
or U497 (N_497,In_2153,In_547);
nand U498 (N_498,In_1466,In_2521);
and U499 (N_499,In_4789,In_1537);
or U500 (N_500,In_2949,In_720);
and U501 (N_501,In_1532,In_1472);
or U502 (N_502,In_3680,In_713);
or U503 (N_503,In_919,In_4430);
nand U504 (N_504,In_442,In_2659);
or U505 (N_505,In_2668,In_2519);
or U506 (N_506,In_460,In_783);
nor U507 (N_507,In_621,In_4373);
and U508 (N_508,In_4116,In_3436);
nor U509 (N_509,In_1813,In_2882);
and U510 (N_510,In_2439,In_2897);
nand U511 (N_511,In_1641,In_1179);
nand U512 (N_512,In_3297,In_4318);
nor U513 (N_513,In_1863,In_4007);
or U514 (N_514,In_4208,In_3078);
nor U515 (N_515,In_315,In_3906);
nor U516 (N_516,In_253,In_1533);
nand U517 (N_517,In_4230,In_1907);
nor U518 (N_518,In_3222,In_976);
and U519 (N_519,In_1006,In_3948);
or U520 (N_520,In_1302,In_2228);
xnor U521 (N_521,In_2364,In_1729);
nor U522 (N_522,In_4316,In_4147);
or U523 (N_523,In_1589,In_4819);
or U524 (N_524,In_1892,In_4304);
nand U525 (N_525,In_4243,In_1245);
and U526 (N_526,In_3915,In_2084);
and U527 (N_527,In_3703,In_3426);
and U528 (N_528,In_248,In_439);
nor U529 (N_529,In_2461,In_3313);
or U530 (N_530,In_2915,In_3584);
and U531 (N_531,In_2982,In_4802);
or U532 (N_532,In_3723,In_828);
and U533 (N_533,In_2843,In_4265);
and U534 (N_534,In_1359,In_440);
or U535 (N_535,In_2454,In_1271);
and U536 (N_536,In_3662,In_2797);
or U537 (N_537,In_1377,In_464);
and U538 (N_538,In_1042,In_2603);
or U539 (N_539,In_4784,In_145);
or U540 (N_540,In_3091,In_126);
nand U541 (N_541,In_2511,In_4308);
nor U542 (N_542,In_2198,In_1073);
nand U543 (N_543,In_3599,In_1865);
nand U544 (N_544,In_3135,In_3248);
or U545 (N_545,In_3399,In_2391);
xnor U546 (N_546,In_1704,In_4405);
and U547 (N_547,In_1638,In_819);
nand U548 (N_548,In_899,In_2534);
and U549 (N_549,In_4919,In_3131);
or U550 (N_550,In_722,In_4702);
or U551 (N_551,In_4753,In_1688);
or U552 (N_552,In_4129,In_4550);
nand U553 (N_553,In_967,In_3660);
nor U554 (N_554,In_2577,In_4829);
and U555 (N_555,In_836,In_2251);
and U556 (N_556,In_4856,In_371);
nand U557 (N_557,In_860,In_1872);
and U558 (N_558,In_4572,In_628);
nor U559 (N_559,In_4203,In_690);
nor U560 (N_560,In_826,In_3121);
xnor U561 (N_561,In_3149,In_352);
or U562 (N_562,In_3012,In_980);
nand U563 (N_563,In_3742,In_1292);
nor U564 (N_564,In_4775,In_1746);
or U565 (N_565,In_1345,In_2155);
or U566 (N_566,In_1677,In_2416);
or U567 (N_567,In_1414,In_2933);
and U568 (N_568,In_3329,In_3290);
or U569 (N_569,In_2320,In_1598);
and U570 (N_570,In_2835,In_680);
nand U571 (N_571,In_438,In_2354);
nor U572 (N_572,In_1612,In_414);
and U573 (N_573,In_63,In_3910);
nand U574 (N_574,In_4698,In_4323);
or U575 (N_575,In_1733,In_633);
or U576 (N_576,In_4902,In_1777);
or U577 (N_577,In_1707,In_927);
nor U578 (N_578,In_291,In_1661);
nand U579 (N_579,In_1572,In_1038);
nor U580 (N_580,In_3118,In_4015);
or U581 (N_581,In_4419,In_1261);
and U582 (N_582,In_1820,In_289);
nand U583 (N_583,In_2127,In_3692);
or U584 (N_584,In_3530,In_3523);
xor U585 (N_585,In_10,In_1106);
or U586 (N_586,In_3624,In_4921);
or U587 (N_587,In_2508,In_156);
or U588 (N_588,In_3005,In_1654);
nand U589 (N_589,In_1921,In_387);
nor U590 (N_590,In_2253,In_3821);
nand U591 (N_591,In_2317,In_4621);
nor U592 (N_592,In_4142,In_687);
nand U593 (N_593,In_2816,In_1894);
xor U594 (N_594,In_4248,In_2703);
nand U595 (N_595,In_2068,In_1866);
xnor U596 (N_596,In_2540,In_706);
or U597 (N_597,In_4734,In_1563);
xor U598 (N_598,In_3014,In_3385);
nor U599 (N_599,In_1338,In_905);
nand U600 (N_600,In_4534,In_3059);
or U601 (N_601,In_2080,In_4788);
or U602 (N_602,In_3651,In_3074);
nand U603 (N_603,In_283,In_3700);
or U604 (N_604,In_1330,In_4793);
xor U605 (N_605,In_2657,In_2120);
or U606 (N_606,In_4713,In_2076);
or U607 (N_607,In_866,In_2375);
nor U608 (N_608,In_1908,In_1172);
and U609 (N_609,In_2991,In_4264);
nor U610 (N_610,In_846,In_138);
nand U611 (N_611,In_1980,In_1312);
and U612 (N_612,In_4461,In_3076);
or U613 (N_613,In_3792,In_3263);
nor U614 (N_614,In_3010,In_2462);
nand U615 (N_615,In_2638,In_224);
nand U616 (N_616,In_3303,In_3287);
xnor U617 (N_617,In_4004,In_1020);
and U618 (N_618,In_3064,In_3509);
and U619 (N_619,In_4482,In_4997);
nor U620 (N_620,In_862,In_2878);
nor U621 (N_621,In_2021,In_987);
or U622 (N_622,In_4162,In_1430);
and U623 (N_623,In_1655,In_4774);
nor U624 (N_624,In_2767,In_923);
and U625 (N_625,In_4502,In_1465);
nor U626 (N_626,In_3237,In_3000);
or U627 (N_627,In_2456,In_1366);
xor U628 (N_628,In_441,In_1785);
xnor U629 (N_629,In_742,In_269);
and U630 (N_630,In_2190,In_1013);
and U631 (N_631,In_721,In_1125);
nor U632 (N_632,In_3610,In_3661);
xnor U633 (N_633,In_3067,In_4875);
or U634 (N_634,In_469,In_3874);
and U635 (N_635,In_2944,In_2858);
nor U636 (N_636,In_143,In_3820);
nand U637 (N_637,In_3052,In_1388);
nor U638 (N_638,In_2618,In_4398);
and U639 (N_639,In_2530,In_239);
nand U640 (N_640,In_2098,In_3346);
nand U641 (N_641,In_1126,In_978);
or U642 (N_642,In_2921,In_3857);
or U643 (N_643,In_3815,In_2450);
nand U644 (N_644,In_3071,In_4900);
and U645 (N_645,In_3163,In_648);
and U646 (N_646,In_1927,In_3877);
nand U647 (N_647,In_4942,In_491);
or U648 (N_648,In_271,In_2865);
nand U649 (N_649,In_2314,In_367);
and U650 (N_650,In_188,In_3103);
nor U651 (N_651,In_1001,In_4109);
and U652 (N_652,In_3092,In_4807);
and U653 (N_653,In_2135,In_4507);
or U654 (N_654,In_3050,In_3891);
nor U655 (N_655,In_1469,In_465);
or U656 (N_656,In_691,In_2780);
and U657 (N_657,In_580,In_95);
xnor U658 (N_658,In_685,In_4212);
nor U659 (N_659,In_3291,In_4804);
nor U660 (N_660,In_3996,In_2853);
or U661 (N_661,In_3062,In_4543);
nor U662 (N_662,In_326,In_3234);
or U663 (N_663,In_2412,In_273);
nor U664 (N_664,In_347,In_3684);
and U665 (N_665,In_635,In_4812);
or U666 (N_666,In_3162,In_991);
nand U667 (N_667,In_1804,In_1107);
nand U668 (N_668,In_1146,In_2046);
nand U669 (N_669,In_1973,In_279);
nand U670 (N_670,In_4681,In_4341);
xnor U671 (N_671,In_3337,In_2388);
and U672 (N_672,In_4629,In_708);
and U673 (N_673,In_1151,In_1758);
and U674 (N_674,In_682,In_3381);
or U675 (N_675,In_168,In_1701);
xnor U676 (N_676,In_2204,In_956);
and U677 (N_677,In_957,In_3492);
or U678 (N_678,In_4547,In_1180);
nor U679 (N_679,In_1810,In_1913);
or U680 (N_680,In_3023,In_1358);
and U681 (N_681,In_3379,In_2031);
or U682 (N_682,In_1438,In_1319);
nand U683 (N_683,In_69,In_2092);
and U684 (N_684,In_4776,In_432);
nor U685 (N_685,In_937,In_2160);
nand U686 (N_686,In_2074,In_4200);
nor U687 (N_687,In_4307,In_4275);
or U688 (N_688,In_1560,In_4261);
and U689 (N_689,In_2720,In_3253);
nand U690 (N_690,In_558,In_3471);
and U691 (N_691,In_3668,In_3414);
or U692 (N_692,In_2486,In_1381);
nor U693 (N_693,In_3218,In_1763);
nand U694 (N_694,In_21,In_2275);
nand U695 (N_695,In_834,In_1710);
nand U696 (N_696,In_4394,In_3758);
or U697 (N_697,In_2597,In_395);
nor U698 (N_698,In_3753,In_3494);
xnor U699 (N_699,In_3069,In_4371);
nand U700 (N_700,In_4619,In_278);
or U701 (N_701,In_1898,In_3497);
nand U702 (N_702,In_3500,In_1281);
nand U703 (N_703,In_47,In_2676);
xor U704 (N_704,In_4916,In_3081);
and U705 (N_705,In_3945,In_1564);
nand U706 (N_706,In_4865,In_3160);
xor U707 (N_707,In_1795,In_2418);
and U708 (N_708,In_4737,In_3265);
xor U709 (N_709,In_3403,In_1233);
or U710 (N_710,In_2810,In_801);
or U711 (N_711,In_1427,In_4881);
nor U712 (N_712,In_3883,In_3186);
or U713 (N_713,In_2866,In_228);
nor U714 (N_714,In_999,In_2473);
nor U715 (N_715,In_2435,In_1334);
nor U716 (N_716,In_1446,In_530);
nor U717 (N_717,In_4328,In_724);
nand U718 (N_718,In_793,In_950);
or U719 (N_719,In_2239,In_4259);
or U720 (N_720,In_88,In_2290);
nor U721 (N_721,In_3828,In_550);
and U722 (N_722,In_1211,In_1941);
nand U723 (N_723,In_700,In_637);
nand U724 (N_724,In_2564,In_677);
nand U725 (N_725,In_929,In_1511);
nand U726 (N_726,In_1287,In_4218);
nor U727 (N_727,In_4485,In_4131);
and U728 (N_728,In_2646,In_1398);
and U729 (N_729,In_2774,In_1558);
and U730 (N_730,In_3396,In_3574);
and U731 (N_731,In_601,In_658);
or U732 (N_732,In_940,In_1400);
nor U733 (N_733,In_2348,In_1284);
nand U734 (N_734,In_1270,In_1953);
xor U735 (N_735,In_3957,In_2973);
nor U736 (N_736,In_485,In_1610);
or U737 (N_737,In_4588,In_4719);
xnor U738 (N_738,In_590,In_615);
and U739 (N_739,In_4873,In_1213);
nand U740 (N_740,In_4365,In_4627);
or U741 (N_741,In_1719,In_738);
and U742 (N_742,In_1611,In_3377);
or U743 (N_743,In_1034,In_1504);
xnor U744 (N_744,In_1720,In_1411);
and U745 (N_745,In_1017,In_554);
nand U746 (N_746,In_2872,In_3188);
or U747 (N_747,In_2460,In_4850);
nor U748 (N_748,In_2437,In_2784);
or U749 (N_749,In_1428,In_4193);
nor U750 (N_750,In_3079,In_84);
xnor U751 (N_751,In_3173,In_2097);
nor U752 (N_752,In_4722,In_1622);
nand U753 (N_753,In_2518,In_4815);
or U754 (N_754,In_2292,In_1803);
or U755 (N_755,In_1070,In_4906);
or U756 (N_756,In_4894,In_4423);
or U757 (N_757,In_894,In_403);
or U758 (N_758,In_195,In_517);
or U759 (N_759,In_4683,In_2154);
nand U760 (N_760,In_4772,In_454);
xor U761 (N_761,In_4372,In_81);
or U762 (N_762,In_4143,In_3225);
and U763 (N_763,In_4088,In_4134);
nor U764 (N_764,In_1355,In_1548);
nor U765 (N_765,In_560,In_3953);
nor U766 (N_766,In_1774,In_1471);
nor U767 (N_767,In_3409,In_1988);
nor U768 (N_768,In_4453,In_51);
nand U769 (N_769,In_2813,In_1276);
or U770 (N_770,In_4392,In_3510);
or U771 (N_771,In_65,In_3466);
xor U772 (N_772,In_3360,In_537);
or U773 (N_773,In_4583,In_3146);
nand U774 (N_774,In_2255,In_2470);
nand U775 (N_775,In_1076,In_1000);
nor U776 (N_776,In_2256,In_4796);
nor U777 (N_777,In_276,In_4689);
or U778 (N_778,In_4078,In_3200);
and U779 (N_779,In_4768,In_184);
nand U780 (N_780,In_2115,In_1093);
or U781 (N_781,In_1293,In_1752);
nor U782 (N_782,In_2055,In_4286);
nor U783 (N_783,In_2381,In_1174);
and U784 (N_784,In_2681,In_4091);
or U785 (N_785,In_2211,In_215);
nor U786 (N_786,In_3001,In_2571);
nor U787 (N_787,In_2048,In_3280);
nor U788 (N_788,In_3210,In_3550);
or U789 (N_789,In_4001,In_1500);
and U790 (N_790,In_4634,In_2583);
nand U791 (N_791,In_1392,In_4096);
and U792 (N_792,In_379,In_455);
nand U793 (N_793,In_3648,In_2494);
or U794 (N_794,In_4066,In_1714);
and U795 (N_795,In_4434,In_3772);
nand U796 (N_796,In_4613,In_1829);
or U797 (N_797,In_3357,In_3950);
or U798 (N_798,In_2778,In_1524);
and U799 (N_799,In_3143,In_1410);
and U800 (N_800,In_2959,In_254);
or U801 (N_801,In_4725,In_1990);
nor U802 (N_802,In_1884,In_712);
nor U803 (N_803,In_436,In_3051);
nor U804 (N_804,In_4010,In_2876);
nand U805 (N_805,In_2722,In_3389);
and U806 (N_806,In_2662,In_150);
nor U807 (N_807,In_4039,In_2038);
nand U808 (N_808,In_4659,In_3472);
nand U809 (N_809,In_740,In_2379);
xor U810 (N_810,In_1530,In_4863);
nor U811 (N_811,In_1353,In_2478);
nand U812 (N_812,In_4045,In_592);
nand U813 (N_813,In_2644,In_3640);
and U814 (N_814,In_1647,In_3008);
nand U815 (N_815,In_4518,In_3596);
and U816 (N_816,In_1075,In_1773);
nor U817 (N_817,In_714,In_3439);
and U818 (N_818,In_4079,In_2398);
nand U819 (N_819,In_1051,In_2633);
and U820 (N_820,In_1104,In_4496);
nor U821 (N_821,In_4606,In_1520);
nand U822 (N_822,In_3281,In_4117);
or U823 (N_823,In_392,In_131);
nand U824 (N_824,In_174,In_4668);
nor U825 (N_825,In_3709,In_3557);
nor U826 (N_826,In_106,In_186);
nor U827 (N_827,In_2743,In_4374);
or U828 (N_828,In_1336,In_1814);
or U829 (N_829,In_2749,In_895);
xor U830 (N_830,In_1240,In_180);
nor U831 (N_831,In_907,In_1715);
nand U832 (N_832,In_3657,In_2565);
or U833 (N_833,In_3493,In_758);
nor U834 (N_834,In_3182,In_3203);
nand U835 (N_835,In_3388,In_4139);
nor U836 (N_836,In_1046,In_161);
nand U837 (N_837,In_4330,In_3645);
and U838 (N_838,In_2653,In_2401);
or U839 (N_839,In_840,In_917);
and U840 (N_840,In_2032,In_105);
nor U841 (N_841,In_2264,In_2236);
nand U842 (N_842,In_1900,In_2502);
nor U843 (N_843,In_4554,In_2312);
or U844 (N_844,In_3,In_503);
and U845 (N_845,In_645,In_1515);
or U846 (N_846,In_2163,In_4887);
nor U847 (N_847,In_4210,In_3032);
or U848 (N_848,In_2436,In_4973);
or U849 (N_849,In_4790,In_3279);
nand U850 (N_850,In_4885,In_4570);
nor U851 (N_851,In_813,In_3576);
nor U852 (N_852,In_2191,In_2187);
nand U853 (N_853,In_1753,In_3671);
nand U854 (N_854,In_3577,In_3835);
nor U855 (N_855,In_1529,In_4479);
nor U856 (N_856,In_4416,In_3138);
nand U857 (N_857,In_3765,In_3277);
nor U858 (N_858,In_4744,In_510);
xnor U859 (N_859,In_89,In_1477);
nand U860 (N_860,In_4441,In_1418);
nor U861 (N_861,In_1190,In_562);
xnor U862 (N_862,In_1755,In_1241);
and U863 (N_863,In_2145,In_459);
nor U864 (N_864,In_4439,In_4126);
nand U865 (N_865,In_3100,In_781);
nor U866 (N_866,In_130,In_3728);
or U867 (N_867,In_2812,In_3652);
nor U868 (N_868,In_3220,In_391);
and U869 (N_869,In_1698,In_3802);
or U870 (N_870,In_2214,In_4047);
and U871 (N_871,In_3954,In_461);
and U872 (N_872,In_1984,In_1116);
or U873 (N_873,In_3269,In_4991);
or U874 (N_874,In_2680,In_2700);
nor U875 (N_875,In_2286,In_2711);
nor U876 (N_876,In_948,In_3364);
nor U877 (N_877,In_1628,In_1082);
nor U878 (N_878,In_4148,In_1996);
nor U879 (N_879,In_3043,In_4112);
nand U880 (N_880,In_4229,In_3536);
xnor U881 (N_881,In_4537,In_3097);
nand U882 (N_882,In_3139,In_4651);
nand U883 (N_883,In_3794,In_4859);
nor U884 (N_884,In_2744,In_2981);
nor U885 (N_885,In_292,In_282);
or U886 (N_886,In_4108,In_3018);
nor U887 (N_887,In_730,In_3900);
or U888 (N_888,In_3428,In_2231);
and U889 (N_889,In_2232,In_2805);
and U890 (N_890,In_2605,In_489);
nand U891 (N_891,In_3105,In_3451);
or U892 (N_892,In_4946,In_1845);
nor U893 (N_893,In_4813,In_1881);
nor U894 (N_894,In_482,In_3818);
and U895 (N_895,In_4165,In_2781);
nand U896 (N_896,In_3916,In_1325);
nor U897 (N_897,In_2782,In_3993);
nor U898 (N_898,In_3284,In_1679);
nor U899 (N_899,In_4036,In_4809);
nand U900 (N_900,In_14,In_2740);
or U901 (N_901,In_1764,In_3881);
nand U902 (N_902,In_4792,In_2786);
or U903 (N_903,In_1468,In_4106);
and U904 (N_904,In_4448,In_2948);
nor U905 (N_905,In_3579,In_3563);
and U906 (N_906,In_4816,In_1417);
nand U907 (N_907,In_2988,In_2886);
or U908 (N_908,In_4043,In_1278);
or U909 (N_909,In_3007,In_3165);
and U910 (N_910,In_611,In_3862);
and U911 (N_911,In_56,In_4017);
and U912 (N_912,In_107,In_2122);
or U913 (N_913,In_1567,In_1579);
and U914 (N_914,In_2293,In_3595);
nand U915 (N_915,In_3585,In_3782);
or U916 (N_916,In_1420,In_811);
nor U917 (N_917,In_3830,In_4517);
nor U918 (N_918,In_423,In_377);
or U919 (N_919,In_2090,In_4878);
xnor U920 (N_920,In_824,In_1095);
or U921 (N_921,In_709,In_3174);
xnor U922 (N_922,In_1535,In_1544);
nand U923 (N_923,In_3324,In_3115);
nand U924 (N_924,In_4475,In_3971);
or U925 (N_925,In_1761,In_405);
xor U926 (N_926,In_4892,In_297);
nand U927 (N_927,In_3817,In_1682);
nand U928 (N_928,In_3450,In_1153);
nor U929 (N_929,In_4969,In_1109);
and U930 (N_930,In_4422,In_4686);
nor U931 (N_931,In_1590,In_2859);
nor U932 (N_932,In_1480,In_1003);
xor U933 (N_933,In_3984,In_1188);
nor U934 (N_934,In_3404,In_2487);
or U935 (N_935,In_1303,In_2554);
nand U936 (N_936,In_4234,In_3555);
and U937 (N_937,In_4983,In_3060);
nor U938 (N_938,In_1616,In_24);
and U939 (N_939,In_3630,In_148);
nor U940 (N_940,In_536,In_2630);
or U941 (N_941,In_426,In_2758);
nand U942 (N_942,In_280,In_336);
nor U943 (N_943,In_2690,In_2645);
nor U944 (N_944,In_3712,In_4414);
nand U945 (N_945,In_857,In_951);
nor U946 (N_946,In_1432,In_1122);
nand U947 (N_947,In_1021,In_4525);
and U948 (N_948,In_2049,In_2732);
and U949 (N_949,In_3607,In_1972);
and U950 (N_950,In_4945,In_93);
and U951 (N_951,In_4443,In_3814);
or U952 (N_952,In_4198,In_4718);
or U953 (N_953,In_746,In_256);
or U954 (N_954,In_838,In_1455);
nor U955 (N_955,In_652,In_4216);
nand U956 (N_956,In_57,In_399);
or U957 (N_957,In_4028,In_83);
nand U958 (N_958,In_4350,In_4982);
or U959 (N_959,In_4299,In_871);
nand U960 (N_960,In_144,In_4761);
nand U961 (N_961,In_2980,In_4400);
nor U962 (N_962,In_1910,In_1182);
xor U963 (N_963,In_3310,In_2785);
and U964 (N_964,In_2908,In_1505);
and U965 (N_965,In_2056,In_4256);
or U966 (N_966,In_2329,In_2604);
nand U967 (N_967,In_3304,In_437);
nand U968 (N_968,In_3810,In_2541);
and U969 (N_969,In_1978,In_3568);
xnor U970 (N_970,In_3619,In_2404);
and U971 (N_971,In_3975,In_1140);
nand U972 (N_972,In_3002,In_4569);
and U973 (N_973,In_1974,In_2532);
nor U974 (N_974,In_4729,In_736);
nor U975 (N_975,In_1201,In_2);
and U976 (N_976,In_2958,In_1102);
or U977 (N_977,In_472,In_1194);
or U978 (N_978,In_2965,In_4207);
and U979 (N_979,In_3147,In_55);
nand U980 (N_980,In_111,In_4553);
nor U981 (N_981,In_2342,In_2729);
or U982 (N_982,In_3569,In_3221);
or U983 (N_983,In_3056,In_2602);
and U984 (N_984,In_4389,In_4587);
or U985 (N_985,In_4488,In_1039);
and U986 (N_986,In_756,In_3816);
nand U987 (N_987,In_2413,In_4664);
and U988 (N_988,In_3664,In_745);
nand U989 (N_989,In_2962,In_4046);
and U990 (N_990,In_3659,In_4663);
or U991 (N_991,In_2258,In_1646);
nand U992 (N_992,In_3937,In_3370);
or U993 (N_993,In_4179,In_3856);
xnor U994 (N_994,In_115,In_4652);
nand U995 (N_995,In_394,In_4846);
nor U996 (N_996,In_4354,In_939);
and U997 (N_997,In_3292,In_833);
nor U998 (N_998,In_4738,In_1386);
xnor U999 (N_999,In_1,In_2685);
and U1000 (N_1000,In_2066,In_2240);
or U1001 (N_1001,In_4269,In_1288);
nor U1002 (N_1002,In_2304,In_4928);
nor U1003 (N_1003,In_3839,In_2016);
and U1004 (N_1004,In_3400,In_808);
and U1005 (N_1005,In_4287,In_1821);
and U1006 (N_1006,In_4172,In_3272);
and U1007 (N_1007,In_3833,In_1460);
and U1008 (N_1008,In_540,In_3117);
xnor U1009 (N_1009,In_1399,In_1149);
and U1010 (N_1010,In_3401,In_2580);
nor U1011 (N_1011,In_3099,In_4471);
or U1012 (N_1012,In_39,In_3233);
nor U1013 (N_1013,In_2770,In_2796);
or U1014 (N_1014,In_2710,In_2039);
or U1015 (N_1015,In_4970,In_4498);
nor U1016 (N_1016,In_4567,In_1556);
nor U1017 (N_1017,In_3724,In_2854);
and U1018 (N_1018,In_1043,In_4697);
nor U1019 (N_1019,In_4646,In_97);
and U1020 (N_1020,In_2880,In_4362);
nor U1021 (N_1021,In_2050,In_4490);
nor U1022 (N_1022,In_2914,In_1971);
or U1023 (N_1023,In_2689,In_3800);
and U1024 (N_1024,In_608,In_3011);
and U1025 (N_1025,In_1145,In_1269);
nor U1026 (N_1026,In_2828,In_4682);
and U1027 (N_1027,In_3970,In_3635);
or U1028 (N_1028,In_3201,In_785);
and U1029 (N_1029,In_3194,In_673);
or U1030 (N_1030,In_1632,In_2064);
or U1031 (N_1031,In_3517,In_262);
and U1032 (N_1032,In_2234,In_1891);
xor U1033 (N_1033,In_2072,In_3741);
nand U1034 (N_1034,In_874,In_1443);
nand U1035 (N_1035,In_339,In_2273);
or U1036 (N_1036,In_497,In_791);
nor U1037 (N_1037,In_4227,In_1279);
xnor U1038 (N_1038,In_553,In_3565);
and U1039 (N_1039,In_1137,In_3475);
xor U1040 (N_1040,In_3299,In_4500);
or U1041 (N_1041,In_4610,In_4510);
nor U1042 (N_1042,In_2977,In_4242);
nand U1043 (N_1043,In_4506,In_1630);
nor U1044 (N_1044,In_1929,In_1727);
or U1045 (N_1045,In_2242,In_3055);
nand U1046 (N_1046,In_2624,In_761);
nand U1047 (N_1047,In_743,In_68);
nand U1048 (N_1048,In_818,In_1656);
xnor U1049 (N_1049,In_3677,In_4417);
and U1050 (N_1050,In_3300,In_1748);
and U1051 (N_1051,In_28,In_3980);
or U1052 (N_1052,In_3801,In_318);
xnor U1053 (N_1053,In_625,In_2579);
nand U1054 (N_1054,In_2751,In_1487);
nor U1055 (N_1055,In_4293,In_3755);
and U1056 (N_1056,In_1834,In_2575);
nor U1057 (N_1057,In_3588,In_3537);
nand U1058 (N_1058,In_167,In_1840);
and U1059 (N_1059,In_244,In_1983);
nor U1060 (N_1060,In_2733,In_973);
nor U1061 (N_1061,In_1252,In_3608);
xor U1062 (N_1062,In_1263,In_419);
or U1063 (N_1063,In_366,In_1723);
and U1064 (N_1064,In_2795,In_401);
nor U1065 (N_1065,In_2663,In_1132);
and U1066 (N_1066,In_3086,In_844);
xor U1067 (N_1067,In_847,In_823);
and U1068 (N_1068,In_2990,In_3940);
and U1069 (N_1069,In_2367,In_2789);
nand U1070 (N_1070,In_2611,In_1749);
nor U1071 (N_1071,In_2890,In_2308);
and U1072 (N_1072,In_1436,In_1859);
and U1073 (N_1073,In_3239,In_330);
nand U1074 (N_1074,In_3969,In_158);
or U1075 (N_1075,In_1904,In_2667);
or U1076 (N_1076,In_926,In_400);
or U1077 (N_1077,In_1209,In_2996);
and U1078 (N_1078,In_1745,In_1711);
nor U1079 (N_1079,In_4359,In_4576);
or U1080 (N_1080,In_2114,In_3845);
nor U1081 (N_1081,In_3421,In_225);
nor U1082 (N_1082,In_763,In_4063);
nand U1083 (N_1083,In_2734,In_3559);
xnor U1084 (N_1084,In_3776,In_4204);
and U1085 (N_1085,In_3487,In_1670);
or U1086 (N_1086,In_3025,In_2295);
or U1087 (N_1087,In_1935,In_15);
nor U1088 (N_1088,In_2148,In_2975);
nand U1089 (N_1089,In_373,In_4624);
nor U1090 (N_1090,In_2851,In_1161);
xnor U1091 (N_1091,In_4635,In_2238);
xnor U1092 (N_1092,In_790,In_2058);
or U1093 (N_1093,In_340,In_3729);
nand U1094 (N_1094,In_3456,In_4018);
nor U1095 (N_1095,In_285,In_3554);
or U1096 (N_1096,In_1975,In_1464);
nand U1097 (N_1097,In_157,In_4548);
and U1098 (N_1098,In_1620,In_3098);
nand U1099 (N_1099,In_3452,In_2180);
xor U1100 (N_1100,In_1645,In_1117);
and U1101 (N_1101,In_1128,In_1542);
and U1102 (N_1102,In_1449,In_2207);
nor U1103 (N_1103,In_4596,In_1088);
nor U1104 (N_1104,In_4309,In_159);
and U1105 (N_1105,In_2769,In_3305);
nor U1106 (N_1106,In_3720,In_1060);
and U1107 (N_1107,In_1453,In_112);
xor U1108 (N_1108,In_1092,In_814);
nor U1109 (N_1109,In_2989,In_2162);
or U1110 (N_1110,In_4082,In_122);
nor U1111 (N_1111,In_4535,In_4037);
nand U1112 (N_1112,In_4630,In_4176);
xnor U1113 (N_1113,In_447,In_845);
nand U1114 (N_1114,In_3125,In_728);
nand U1115 (N_1115,In_3539,In_3804);
or U1116 (N_1116,In_4828,In_731);
and U1117 (N_1117,In_420,In_18);
nor U1118 (N_1118,In_210,In_3454);
nor U1119 (N_1119,In_4253,In_4384);
xnor U1120 (N_1120,In_4180,In_3947);
nand U1121 (N_1121,In_1344,In_3694);
nor U1122 (N_1122,In_2779,In_944);
xnor U1123 (N_1123,In_729,In_3780);
nand U1124 (N_1124,In_1450,In_842);
nand U1125 (N_1125,In_1875,In_223);
nor U1126 (N_1126,In_546,In_2108);
or U1127 (N_1127,In_696,In_780);
nor U1128 (N_1128,In_1262,In_3701);
and U1129 (N_1129,In_2832,In_4951);
nand U1130 (N_1130,In_4364,In_1683);
nor U1131 (N_1131,In_958,In_32);
nand U1132 (N_1132,In_1035,In_1350);
or U1133 (N_1133,In_4656,In_3527);
xor U1134 (N_1134,In_4493,In_3240);
nor U1135 (N_1135,In_4292,In_2325);
or U1136 (N_1136,In_4593,In_3369);
nand U1137 (N_1137,In_1337,In_2125);
and U1138 (N_1138,In_4118,In_4794);
nor U1139 (N_1139,In_4188,In_3406);
nor U1140 (N_1140,In_3951,In_11);
nand U1141 (N_1141,In_4068,In_2822);
and U1142 (N_1142,In_1769,In_3030);
and U1143 (N_1143,In_172,In_3057);
xnor U1144 (N_1144,In_1673,In_4342);
nand U1145 (N_1145,In_1867,In_2201);
or U1146 (N_1146,In_4748,In_23);
nand U1147 (N_1147,In_3952,In_1928);
xor U1148 (N_1148,In_4053,In_1272);
nor U1149 (N_1149,In_2830,In_2200);
or U1150 (N_1150,In_4303,In_3242);
and U1151 (N_1151,In_452,In_1552);
and U1152 (N_1152,In_1588,In_4853);
or U1153 (N_1153,In_2067,In_3672);
and U1154 (N_1154,In_1086,In_3089);
and U1155 (N_1155,In_3518,In_3353);
and U1156 (N_1156,In_3470,In_4190);
and U1157 (N_1157,In_1772,In_338);
nor U1158 (N_1158,In_1998,In_1985);
nor U1159 (N_1159,In_2953,In_298);
and U1160 (N_1160,In_2871,In_3016);
or U1161 (N_1161,In_2623,In_656);
nor U1162 (N_1162,In_2468,In_3416);
nand U1163 (N_1163,In_4263,In_3283);
xnor U1164 (N_1164,In_2702,In_3122);
nand U1165 (N_1165,In_1523,In_3561);
or U1166 (N_1166,In_1539,In_4571);
or U1167 (N_1167,In_216,In_2666);
and U1168 (N_1168,In_3622,In_581);
or U1169 (N_1169,In_4222,In_185);
or U1170 (N_1170,In_3787,In_2310);
nand U1171 (N_1171,In_1685,In_3707);
and U1172 (N_1172,In_2972,In_3243);
nand U1173 (N_1173,In_4489,In_2378);
or U1174 (N_1174,In_233,In_622);
nor U1175 (N_1175,In_2517,In_4608);
nor U1176 (N_1176,In_260,In_4561);
nor U1177 (N_1177,In_2557,In_4847);
or U1178 (N_1178,In_201,In_2230);
nor U1179 (N_1179,In_3943,In_568);
nor U1180 (N_1180,In_2861,In_820);
and U1181 (N_1181,In_3806,In_3336);
nor U1182 (N_1182,In_3144,In_1499);
or U1183 (N_1183,In_1313,In_3995);
or U1184 (N_1184,In_4345,In_4864);
nand U1185 (N_1185,In_1937,In_435);
and U1186 (N_1186,In_1893,In_3863);
nand U1187 (N_1187,In_2574,In_4628);
nand U1188 (N_1188,In_354,In_2697);
or U1189 (N_1189,In_3521,In_3294);
or U1190 (N_1190,In_4410,In_2520);
nor U1191 (N_1191,In_2684,In_1062);
or U1192 (N_1192,In_3250,In_120);
xnor U1193 (N_1193,In_457,In_1690);
or U1194 (N_1194,In_4300,In_1235);
nor U1195 (N_1195,In_2269,In_2147);
nand U1196 (N_1196,In_1778,In_3231);
or U1197 (N_1197,In_2669,In_3799);
nor U1198 (N_1198,In_3154,In_934);
nand U1199 (N_1199,In_4814,In_1421);
nand U1200 (N_1200,In_1202,In_2341);
nor U1201 (N_1201,In_1422,In_900);
nor U1202 (N_1202,In_4657,In_2444);
and U1203 (N_1203,In_2589,In_1349);
or U1204 (N_1204,In_646,In_1643);
or U1205 (N_1205,In_3888,In_3150);
nand U1206 (N_1206,In_3604,In_1314);
nor U1207 (N_1207,In_4460,In_4282);
or U1208 (N_1208,In_2111,In_4830);
nand U1209 (N_1209,In_4418,In_4285);
nor U1210 (N_1210,In_3697,In_386);
or U1211 (N_1211,In_832,In_2352);
nor U1212 (N_1212,In_4026,In_304);
or U1213 (N_1213,In_4810,In_732);
nand U1214 (N_1214,In_725,In_2984);
nand U1215 (N_1215,In_2884,In_4638);
nand U1216 (N_1216,In_389,In_3985);
or U1217 (N_1217,In_4963,In_4296);
or U1218 (N_1218,In_1830,In_1296);
nand U1219 (N_1219,In_1360,In_2060);
nand U1220 (N_1220,In_1961,In_3359);
xnor U1221 (N_1221,In_365,In_2894);
nor U1222 (N_1222,In_3254,In_509);
nor U1223 (N_1223,In_3580,In_4124);
or U1224 (N_1224,In_1273,In_4024);
or U1225 (N_1225,In_312,In_3967);
nor U1226 (N_1226,In_2423,In_2582);
nand U1227 (N_1227,In_4723,In_1575);
nor U1228 (N_1228,In_2402,In_3570);
xnor U1229 (N_1229,In_1120,In_3754);
or U1230 (N_1230,In_4655,In_364);
nand U1231 (N_1231,In_3892,In_2194);
or U1232 (N_1232,In_231,In_3841);
nand U1233 (N_1233,In_4765,In_1823);
or U1234 (N_1234,In_1015,In_2386);
xnor U1235 (N_1235,In_1614,In_966);
nor U1236 (N_1236,In_266,In_1224);
nor U1237 (N_1237,In_1119,In_2719);
or U1238 (N_1238,In_3615,In_1324);
nor U1239 (N_1239,In_2257,In_1071);
and U1240 (N_1240,In_2300,In_2102);
and U1241 (N_1241,In_1280,In_3691);
or U1242 (N_1242,In_4334,In_1333);
nand U1243 (N_1243,In_2082,In_2103);
nor U1244 (N_1244,In_651,In_4747);
nor U1245 (N_1245,In_4246,In_2426);
xnor U1246 (N_1246,In_3459,In_2054);
nand U1247 (N_1247,In_1223,In_852);
xor U1248 (N_1248,In_4832,In_1917);
or U1249 (N_1249,In_3338,In_2335);
nand U1250 (N_1250,In_2841,In_2909);
nor U1251 (N_1251,In_17,In_249);
nor U1252 (N_1252,In_4922,In_4833);
and U1253 (N_1253,In_3190,In_3587);
and U1254 (N_1254,In_3177,In_4769);
nor U1255 (N_1255,In_4728,In_2377);
nor U1256 (N_1256,In_3904,In_649);
nor U1257 (N_1257,In_4270,In_1074);
or U1258 (N_1258,In_1993,In_1861);
nand U1259 (N_1259,In_3687,In_4952);
and U1260 (N_1260,In_1739,In_1578);
and U1261 (N_1261,In_1096,In_137);
and U1262 (N_1262,In_2452,In_4644);
nand U1263 (N_1263,In_3443,In_3744);
nand U1264 (N_1264,In_928,In_1047);
and U1265 (N_1265,In_2936,In_311);
or U1266 (N_1266,In_2252,In_496);
nor U1267 (N_1267,In_4113,In_3127);
or U1268 (N_1268,In_2999,In_3274);
nor U1269 (N_1269,In_3387,In_2566);
xor U1270 (N_1270,In_4735,In_778);
and U1271 (N_1271,In_3003,In_2376);
nand U1272 (N_1272,In_1425,In_3734);
nand U1273 (N_1273,In_3412,In_1009);
and U1274 (N_1274,In_1163,In_4272);
xnor U1275 (N_1275,In_2387,In_3854);
nor U1276 (N_1276,In_3430,In_3666);
nor U1277 (N_1277,In_2837,In_3847);
nand U1278 (N_1278,In_3347,In_1914);
nand U1279 (N_1279,In_3779,In_1781);
or U1280 (N_1280,In_1849,In_431);
nor U1281 (N_1281,In_1452,In_3306);
xnor U1282 (N_1282,In_3549,In_2451);
nand U1283 (N_1283,In_3354,In_1317);
nand U1284 (N_1284,In_4590,In_4432);
xnor U1285 (N_1285,In_1547,In_2931);
nor U1286 (N_1286,In_4603,In_4860);
nand U1287 (N_1287,In_2403,In_1633);
or U1288 (N_1288,In_2087,In_970);
and U1289 (N_1289,In_2134,In_1926);
and U1290 (N_1290,In_383,In_3425);
and U1291 (N_1291,In_3853,In_4909);
nand U1292 (N_1292,In_128,In_4206);
or U1293 (N_1293,In_4199,In_2942);
nor U1294 (N_1294,In_512,In_2790);
nor U1295 (N_1295,In_1780,In_4375);
or U1296 (N_1296,In_2362,In_2651);
and U1297 (N_1297,In_1268,In_3956);
nor U1298 (N_1298,In_2480,In_261);
and U1299 (N_1299,In_2550,In_2104);
xor U1300 (N_1300,In_4914,In_4975);
and U1301 (N_1301,In_3245,In_1518);
xnor U1302 (N_1302,In_1905,In_4411);
and U1303 (N_1303,In_1882,In_98);
or U1304 (N_1304,In_1025,In_599);
nor U1305 (N_1305,In_3045,In_4779);
nor U1306 (N_1306,In_1793,In_4840);
xor U1307 (N_1307,In_2289,In_3987);
or U1308 (N_1308,In_4130,In_4332);
and U1309 (N_1309,In_4074,In_1222);
xnor U1310 (N_1310,In_2693,In_2189);
or U1311 (N_1311,In_3533,In_2433);
nor U1312 (N_1312,In_4757,In_1966);
xnor U1313 (N_1313,In_1295,In_1065);
and U1314 (N_1314,In_1111,In_3726);
nand U1315 (N_1315,In_4531,In_3545);
nand U1316 (N_1316,In_2493,In_1962);
nor U1317 (N_1317,In_307,In_2891);
or U1318 (N_1318,In_3981,In_2170);
xor U1319 (N_1319,In_3795,In_2441);
or U1320 (N_1320,In_3824,In_2787);
xnor U1321 (N_1321,In_1870,In_384);
xor U1322 (N_1322,In_1837,In_1939);
and U1323 (N_1323,In_397,In_2410);
and U1324 (N_1324,In_3851,In_3184);
and U1325 (N_1325,In_378,In_2919);
nand U1326 (N_1326,In_1404,In_2197);
nor U1327 (N_1327,In_2907,In_605);
nand U1328 (N_1328,In_3852,In_4484);
nand U1329 (N_1329,In_1310,In_1402);
nand U1330 (N_1330,In_2466,In_2044);
xor U1331 (N_1331,In_2062,In_337);
and U1332 (N_1332,In_2165,In_409);
nand U1333 (N_1333,In_3423,In_916);
nand U1334 (N_1334,In_4407,In_3885);
nand U1335 (N_1335,In_3321,In_3199);
nand U1336 (N_1336,In_4978,In_1999);
nor U1337 (N_1337,In_1676,In_52);
or U1338 (N_1338,In_4136,In_2970);
nand U1339 (N_1339,In_4343,In_1768);
nor U1340 (N_1340,In_3629,In_4452);
nor U1341 (N_1341,In_4981,In_3944);
xnor U1342 (N_1342,In_136,In_3583);
or U1343 (N_1343,In_936,In_3382);
nand U1344 (N_1344,In_1828,In_0);
and U1345 (N_1345,In_4626,In_2419);
and U1346 (N_1346,In_3159,In_147);
nor U1347 (N_1347,In_2935,In_572);
and U1348 (N_1348,In_979,In_4023);
or U1349 (N_1349,In_1285,In_4196);
nand U1350 (N_1350,In_771,In_2801);
or U1351 (N_1351,In_2615,In_3386);
xor U1352 (N_1352,In_3693,In_997);
nor U1353 (N_1353,In_4504,In_1321);
nand U1354 (N_1354,In_4665,In_1124);
and U1355 (N_1355,In_4030,In_3713);
or U1356 (N_1356,In_1987,In_368);
nand U1357 (N_1357,In_525,In_13);
and U1358 (N_1358,In_1871,In_2838);
and U1359 (N_1359,In_2608,In_3958);
xor U1360 (N_1360,In_1187,In_946);
and U1361 (N_1361,In_719,In_2920);
or U1362 (N_1362,In_3541,In_2168);
xnor U1363 (N_1363,In_1880,In_1930);
and U1364 (N_1364,In_1697,In_4361);
nor U1365 (N_1365,In_325,In_1507);
or U1366 (N_1366,In_3747,In_1108);
nand U1367 (N_1367,In_589,In_4831);
nand U1368 (N_1368,In_770,In_1982);
nor U1369 (N_1369,In_4527,In_2414);
xnor U1370 (N_1370,In_1819,In_2137);
nand U1371 (N_1371,In_443,In_2929);
nand U1372 (N_1372,In_3447,In_1846);
and U1373 (N_1373,In_3731,In_3004);
and U1374 (N_1374,In_3522,In_2303);
nand U1375 (N_1375,In_1674,In_4870);
nor U1376 (N_1376,In_3486,In_2213);
xnor U1377 (N_1377,In_3244,In_2085);
nor U1378 (N_1378,In_4173,In_4855);
xor U1379 (N_1379,In_809,In_4612);
nor U1380 (N_1380,In_2282,In_411);
or U1381 (N_1381,In_2764,In_1012);
xnor U1382 (N_1382,In_4985,In_1294);
nor U1383 (N_1383,In_1566,In_872);
and U1384 (N_1384,In_993,In_4758);
nand U1385 (N_1385,In_4965,In_3920);
and U1386 (N_1386,In_3968,In_4824);
or U1387 (N_1387,In_2763,In_2636);
or U1388 (N_1388,In_3417,In_1826);
or U1389 (N_1389,In_3351,In_4138);
and U1390 (N_1390,In_2868,In_3919);
nand U1391 (N_1391,In_1212,In_1061);
nand U1392 (N_1392,In_3495,In_1378);
nor U1393 (N_1393,In_3019,In_831);
and U1394 (N_1394,In_1014,In_3524);
nand U1395 (N_1395,In_2932,In_2714);
nand U1396 (N_1396,In_2241,In_499);
and U1397 (N_1397,In_576,In_1512);
or U1398 (N_1398,In_4986,In_2075);
nand U1399 (N_1399,In_3773,In_1403);
nand U1400 (N_1400,In_3571,In_668);
nor U1401 (N_1401,In_1607,In_909);
or U1402 (N_1402,In_4781,In_717);
xor U1403 (N_1403,In_2244,In_3318);
or U1404 (N_1404,In_2754,In_2898);
or U1405 (N_1405,In_4767,In_234);
nor U1406 (N_1406,In_4368,In_444);
nor U1407 (N_1407,In_2934,In_43);
or U1408 (N_1408,In_3893,In_1085);
xnor U1409 (N_1409,In_3609,In_2173);
xor U1410 (N_1410,In_4852,In_2671);
and U1411 (N_1411,In_3440,In_1668);
or U1412 (N_1412,In_4648,In_1634);
and U1413 (N_1413,In_2011,In_1551);
xor U1414 (N_1414,In_1706,In_2477);
nor U1415 (N_1415,In_3566,In_2216);
nand U1416 (N_1416,In_2546,In_681);
or U1417 (N_1417,In_2609,In_1127);
nor U1418 (N_1418,In_1694,In_363);
or U1419 (N_1419,In_4861,In_415);
and U1420 (N_1420,In_1457,In_4084);
or U1421 (N_1421,In_121,In_3072);
xnor U1422 (N_1422,In_888,In_3902);
nand U1423 (N_1423,In_2042,In_1561);
nand U1424 (N_1424,In_44,In_3164);
nor U1425 (N_1425,In_1969,In_1491);
and U1426 (N_1426,In_3889,In_1818);
nand U1427 (N_1427,In_1068,In_376);
or U1428 (N_1428,In_1853,In_3542);
or U1429 (N_1429,In_3914,In_3395);
and U1430 (N_1430,In_890,In_3344);
nand U1431 (N_1431,In_1008,In_3732);
or U1432 (N_1432,In_4791,In_42);
and U1433 (N_1433,In_3769,In_3334);
xor U1434 (N_1434,In_1797,In_4123);
and U1435 (N_1435,In_2018,In_2440);
xor U1436 (N_1436,In_220,In_3155);
or U1437 (N_1437,In_1461,In_674);
and U1438 (N_1438,In_1587,In_320);
nand U1439 (N_1439,In_2040,In_382);
and U1440 (N_1440,In_627,In_2950);
or U1441 (N_1441,In_3335,In_372);
or U1442 (N_1442,In_2438,In_2947);
nand U1443 (N_1443,In_2052,In_2824);
nand U1444 (N_1444,In_3922,In_2319);
and U1445 (N_1445,In_410,In_4060);
and U1446 (N_1446,In_1437,In_4174);
nor U1447 (N_1447,In_449,In_1144);
xor U1448 (N_1448,In_272,In_2363);
nand U1449 (N_1449,In_1580,In_1497);
nand U1450 (N_1450,In_1230,In_4353);
xnor U1451 (N_1451,In_1246,In_1185);
and U1452 (N_1452,In_4301,In_2366);
or U1453 (N_1453,In_1148,In_4605);
nor U1454 (N_1454,In_4127,In_2570);
nor U1455 (N_1455,In_4101,In_1799);
nand U1456 (N_1456,In_631,In_4033);
nor U1457 (N_1457,In_1078,In_4777);
or U1458 (N_1458,In_94,In_3235);
nor U1459 (N_1459,In_2652,In_2106);
or U1460 (N_1460,In_4929,In_2047);
or U1461 (N_1461,In_1631,In_3170);
and U1462 (N_1462,In_1429,In_4594);
or U1463 (N_1463,In_4771,In_2459);
xor U1464 (N_1464,In_49,In_3034);
nor U1465 (N_1465,In_2501,In_4609);
nor U1466 (N_1466,In_4746,In_3468);
nand U1467 (N_1467,In_2581,In_4022);
xor U1468 (N_1468,In_3698,In_3690);
and U1469 (N_1469,In_4393,In_1072);
nand U1470 (N_1470,In_2005,In_2617);
nand U1471 (N_1471,In_4169,In_3546);
xor U1472 (N_1472,In_2458,In_4566);
or U1473 (N_1473,In_1933,In_2955);
and U1474 (N_1474,In_2151,In_3977);
or U1475 (N_1475,In_3682,In_4201);
and U1476 (N_1476,In_1957,In_4085);
nor U1477 (N_1477,In_4563,In_665);
nor U1478 (N_1478,In_1604,In_1164);
or U1479 (N_1479,In_1301,In_1238);
or U1480 (N_1480,In_2998,In_1363);
or U1481 (N_1481,In_2107,In_2488);
nand U1482 (N_1482,In_117,In_4801);
or U1483 (N_1483,In_1625,In_4465);
nand U1484 (N_1484,In_398,In_1981);
or U1485 (N_1485,In_1650,In_1251);
nand U1486 (N_1486,In_2682,In_4450);
and U1487 (N_1487,In_3562,In_2261);
nor U1488 (N_1488,In_1526,In_2263);
xnor U1489 (N_1489,In_2182,In_3411);
or U1490 (N_1490,In_2621,In_2625);
xor U1491 (N_1491,In_494,In_2730);
nand U1492 (N_1492,In_3419,In_3846);
xor U1493 (N_1493,In_4225,In_2008);
and U1494 (N_1494,In_4041,In_2927);
nor U1495 (N_1495,In_1922,In_4841);
and U1496 (N_1496,In_80,In_1540);
and U1497 (N_1497,In_3267,In_739);
nor U1498 (N_1498,In_3063,In_555);
and U1499 (N_1499,In_3899,In_2612);
xor U1500 (N_1500,In_3994,In_300);
or U1501 (N_1501,In_313,In_910);
xor U1502 (N_1502,In_1253,In_3964);
and U1503 (N_1503,In_1387,In_2007);
nor U1504 (N_1504,In_1596,In_4167);
and U1505 (N_1505,In_2028,In_4825);
nand U1506 (N_1506,In_777,In_1766);
xor U1507 (N_1507,In_2101,In_2382);
and U1508 (N_1508,In_4992,In_1613);
or U1509 (N_1509,In_295,In_2209);
nand U1510 (N_1510,In_3761,In_1762);
nand U1511 (N_1511,In_2417,In_2698);
nand U1512 (N_1512,In_2563,In_3432);
nand U1513 (N_1513,In_932,In_4006);
nand U1514 (N_1514,In_193,In_3921);
nor U1515 (N_1515,In_2961,In_2000);
and U1516 (N_1516,In_2002,In_4390);
nand U1517 (N_1517,In_2298,In_2429);
or U1518 (N_1518,In_4277,In_3836);
nor U1519 (N_1519,In_3036,In_22);
or U1520 (N_1520,In_657,In_3434);
and U1521 (N_1521,In_1444,In_3077);
and U1522 (N_1522,In_2027,In_388);
xor U1523 (N_1523,In_4573,In_4568);
and U1524 (N_1524,In_3942,In_1371);
nor U1525 (N_1525,In_1770,In_109);
or U1526 (N_1526,In_1134,In_522);
nor U1527 (N_1527,In_1568,In_574);
and U1528 (N_1528,In_4175,In_2063);
nand U1529 (N_1529,In_349,In_4947);
nor U1530 (N_1530,In_4107,In_2274);
nor U1531 (N_1531,In_2701,In_3749);
nor U1532 (N_1532,In_3317,In_4338);
or U1533 (N_1533,In_1198,In_4467);
nand U1534 (N_1534,In_1105,In_678);
and U1535 (N_1535,In_753,In_3650);
and U1536 (N_1536,In_471,In_1858);
or U1537 (N_1537,In_858,In_3445);
nor U1538 (N_1538,In_4247,In_1033);
or U1539 (N_1539,In_160,In_4014);
xnor U1540 (N_1540,In_1519,In_693);
or U1541 (N_1541,In_1593,In_1225);
nand U1542 (N_1542,In_3649,In_2875);
xor U1543 (N_1543,In_1407,In_4505);
nor U1544 (N_1544,In_1049,In_4964);
nand U1545 (N_1545,In_4712,In_2807);
nand U1546 (N_1546,In_1374,In_3101);
nand U1547 (N_1547,In_4395,In_4260);
nor U1548 (N_1548,In_4838,In_458);
and U1549 (N_1549,In_4844,In_2024);
or U1550 (N_1550,In_4778,In_3503);
xor U1551 (N_1551,In_4540,In_417);
or U1552 (N_1552,In_2634,In_4477);
nand U1553 (N_1553,In_1031,In_2326);
and U1554 (N_1554,In_3054,In_3481);
nand U1555 (N_1555,In_4062,In_4896);
or U1556 (N_1556,In_316,In_2447);
and U1557 (N_1557,In_2964,In_2951);
nand U1558 (N_1558,In_4239,In_3238);
nor U1559 (N_1559,In_2639,In_2538);
xor U1560 (N_1560,In_2146,In_4121);
or U1561 (N_1561,In_726,In_3544);
and U1562 (N_1562,In_662,In_4760);
nor U1563 (N_1563,In_2307,In_4382);
or U1564 (N_1564,In_985,In_1439);
nor U1565 (N_1565,In_2059,In_2235);
nand U1566 (N_1566,In_2449,In_4503);
and U1567 (N_1567,In_1069,In_4401);
and U1568 (N_1568,In_4034,In_3774);
and U1569 (N_1569,In_74,In_4958);
nor U1570 (N_1570,In_3260,In_4020);
or U1571 (N_1571,In_2343,In_3625);
xor U1572 (N_1572,In_3332,In_1771);
and U1573 (N_1573,In_827,In_1824);
and U1574 (N_1574,In_3129,In_3333);
or U1575 (N_1575,In_4194,In_4972);
nand U1576 (N_1576,In_704,In_2945);
nand U1577 (N_1577,In_1362,In_1356);
or U1578 (N_1578,In_478,In_493);
or U1579 (N_1579,In_630,In_155);
nand U1580 (N_1580,In_965,In_3929);
xnor U1581 (N_1581,In_359,In_4019);
nand U1582 (N_1582,In_3183,In_848);
and U1583 (N_1583,In_2906,In_4002);
and U1584 (N_1584,In_3618,In_3232);
nor U1585 (N_1585,In_4238,In_4696);
or U1586 (N_1586,In_4714,In_1391);
and U1587 (N_1587,In_1968,In_3502);
nand U1588 (N_1588,In_3558,In_4160);
and U1589 (N_1589,In_1250,In_4670);
nand U1590 (N_1590,In_4907,In_569);
or U1591 (N_1591,In_2130,In_2206);
nor U1592 (N_1592,In_1143,In_4961);
or U1593 (N_1593,In_2100,In_4232);
xor U1594 (N_1594,In_2527,In_1426);
xnor U1595 (N_1595,In_153,In_1942);
nor U1596 (N_1596,In_1157,In_764);
nor U1597 (N_1597,In_4344,In_1379);
nor U1598 (N_1598,In_502,In_3153);
or U1599 (N_1599,In_3111,In_2179);
nand U1600 (N_1600,In_3227,In_1669);
xor U1601 (N_1601,In_4237,In_4910);
xnor U1602 (N_1602,In_1725,In_650);
xor U1603 (N_1603,In_4327,In_3797);
nor U1604 (N_1604,In_422,In_267);
xor U1605 (N_1605,In_570,In_4556);
nor U1606 (N_1606,In_3181,In_2691);
nor U1607 (N_1607,In_2845,In_2857);
nand U1608 (N_1608,In_2405,In_2392);
or U1609 (N_1609,In_519,In_1097);
xor U1610 (N_1610,In_3298,In_2370);
or U1611 (N_1611,In_727,In_3611);
nor U1612 (N_1612,In_4058,In_1236);
or U1613 (N_1613,In_3483,In_3743);
nor U1614 (N_1614,In_2777,In_3251);
nor U1615 (N_1615,In_614,In_1375);
nand U1616 (N_1616,In_4582,In_1543);
and U1617 (N_1617,In_2356,In_613);
nor U1618 (N_1618,In_1053,In_2792);
nand U1619 (N_1619,In_1485,In_1393);
nand U1620 (N_1620,In_4835,In_559);
and U1621 (N_1621,In_1315,In_2280);
and U1622 (N_1622,In_1026,In_500);
and U1623 (N_1623,In_445,In_3590);
or U1624 (N_1624,In_3080,In_4716);
nor U1625 (N_1625,In_2136,In_1549);
and U1626 (N_1626,In_4075,In_3197);
nor U1627 (N_1627,In_4995,In_4183);
and U1628 (N_1628,In_1765,In_1087);
or U1629 (N_1629,In_1835,In_476);
and U1630 (N_1630,In_448,In_4396);
nand U1631 (N_1631,In_1416,In_3230);
or U1632 (N_1632,In_1686,In_3832);
nor U1633 (N_1633,In_1369,In_1503);
xnor U1634 (N_1634,In_784,In_2910);
nor U1635 (N_1635,In_2529,In_3094);
xor U1636 (N_1636,In_1997,In_4295);
and U1637 (N_1637,In_381,In_2883);
nand U1638 (N_1638,In_3751,In_3479);
or U1639 (N_1639,In_2969,In_3087);
nor U1640 (N_1640,In_4100,In_4352);
and U1641 (N_1641,In_334,In_4480);
or U1642 (N_1642,In_3785,In_332);
and U1643 (N_1643,In_2475,In_2399);
nand U1644 (N_1644,In_2339,In_1887);
or U1645 (N_1645,In_2110,In_915);
nor U1646 (N_1646,In_4005,In_1574);
xnor U1647 (N_1647,In_3157,In_19);
nor U1648 (N_1648,In_1265,In_2772);
or U1649 (N_1649,In_3803,In_4673);
or U1650 (N_1650,In_240,In_2500);
or U1651 (N_1651,In_1951,In_3791);
nand U1652 (N_1652,In_1991,In_1304);
nor U1653 (N_1653,In_2641,In_2768);
nor U1654 (N_1654,In_1594,In_2587);
nand U1655 (N_1655,In_4397,In_4032);
and U1656 (N_1656,In_962,In_466);
xnor U1657 (N_1657,In_175,In_2051);
or U1658 (N_1658,In_1357,In_3617);
nor U1659 (N_1659,In_4463,In_2899);
nand U1660 (N_1660,In_524,In_4501);
and U1661 (N_1661,In_1441,In_3748);
nor U1662 (N_1662,In_1214,In_4536);
nand U1663 (N_1663,In_4420,In_3049);
nor U1664 (N_1664,In_2248,In_412);
or U1665 (N_1665,In_2873,In_3628);
and U1666 (N_1666,In_908,In_1947);
and U1667 (N_1667,In_4706,In_2522);
or U1668 (N_1668,In_3405,In_1956);
or U1669 (N_1669,In_2943,In_1794);
xnor U1670 (N_1670,In_1862,In_1592);
and U1671 (N_1671,In_4278,In_2773);
nor U1672 (N_1672,In_4370,In_3278);
nor U1673 (N_1673,In_3104,In_3505);
nor U1674 (N_1674,In_3865,In_4939);
and U1675 (N_1675,In_78,In_2629);
xor U1676 (N_1676,In_4944,In_4409);
nor U1677 (N_1677,In_4959,In_192);
or U1678 (N_1678,In_4273,In_2568);
nor U1679 (N_1679,In_2512,In_2420);
and U1680 (N_1680,In_4140,In_4128);
nor U1681 (N_1681,In_3474,In_2924);
and U1682 (N_1682,In_4483,In_4402);
or U1683 (N_1683,In_92,In_3960);
nand U1684 (N_1684,In_3669,In_3175);
nor U1685 (N_1685,In_566,In_335);
nor U1686 (N_1686,In_4660,In_3911);
nor U1687 (N_1687,In_1945,In_1305);
nand U1688 (N_1688,In_4512,In_2081);
and U1689 (N_1689,In_768,In_369);
nor U1690 (N_1690,In_1419,In_4637);
and U1691 (N_1691,In_76,In_2432);
xnor U1692 (N_1692,In_4366,In_639);
and U1693 (N_1693,In_3531,In_1653);
nand U1694 (N_1694,In_1902,In_2350);
and U1695 (N_1695,In_3308,In_2385);
or U1696 (N_1696,In_3905,In_830);
and U1697 (N_1697,In_247,In_3394);
nand U1698 (N_1698,In_2679,In_703);
nand U1699 (N_1699,In_4633,In_4459);
nor U1700 (N_1700,In_4064,In_2938);
nor U1701 (N_1701,In_3066,In_3345);
and U1702 (N_1702,In_4103,In_1915);
nand U1703 (N_1703,In_4166,In_2288);
nand U1704 (N_1704,In_270,In_4920);
nor U1705 (N_1705,In_4957,In_1058);
and U1706 (N_1706,In_2065,In_585);
nor U1707 (N_1707,In_3286,In_2306);
or U1708 (N_1708,In_2675,In_3838);
or U1709 (N_1709,In_3342,In_2658);
nor U1710 (N_1710,In_4891,In_2889);
nand U1711 (N_1711,In_6,In_2109);
or U1712 (N_1712,In_945,In_4499);
or U1713 (N_1713,In_3178,In_3315);
nand U1714 (N_1714,In_2203,In_1080);
or U1715 (N_1715,In_904,In_2539);
nor U1716 (N_1716,In_3614,In_4249);
or U1717 (N_1717,In_2053,In_1675);
nand U1718 (N_1718,In_2591,In_577);
nand U1719 (N_1719,In_4110,In_429);
nand U1720 (N_1720,In_2156,In_3191);
or U1721 (N_1721,In_1390,In_600);
nand U1722 (N_1722,In_3028,In_1964);
nand U1723 (N_1723,In_40,In_3021);
nand U1724 (N_1724,In_3675,In_2545);
nand U1725 (N_1725,In_1789,In_508);
xor U1726 (N_1726,In_2818,In_1165);
and U1727 (N_1727,In_3501,In_2766);
or U1728 (N_1728,In_2202,In_686);
nand U1729 (N_1729,In_3123,In_3616);
xnor U1730 (N_1730,In_3913,In_4966);
nor U1731 (N_1731,In_1986,In_1716);
and U1732 (N_1732,In_3793,In_4336);
nor U1733 (N_1733,In_4811,In_2762);
and U1734 (N_1734,In_1138,In_3085);
or U1735 (N_1735,In_142,In_1470);
nand U1736 (N_1736,In_1899,In_342);
xor U1737 (N_1737,In_4472,In_3398);
or U1738 (N_1738,In_3504,In_4823);
and U1739 (N_1739,In_1886,In_468);
or U1740 (N_1740,In_1490,In_407);
nand U1741 (N_1741,In_3444,In_3973);
and U1742 (N_1742,In_4640,In_1896);
nor U1743 (N_1743,In_380,In_483);
xor U1744 (N_1744,In_2268,In_1342);
and U1745 (N_1745,In_3621,In_4707);
and U1746 (N_1746,In_2088,In_1642);
nor U1747 (N_1747,In_3384,In_3455);
and U1748 (N_1748,In_176,In_1277);
xor U1749 (N_1749,In_3031,In_453);
nand U1750 (N_1750,In_4446,In_750);
nor U1751 (N_1751,In_4514,In_2157);
or U1752 (N_1752,In_2739,In_4031);
nand U1753 (N_1753,In_4319,In_3658);
nand U1754 (N_1754,In_1435,In_4444);
nand U1755 (N_1755,In_1848,In_2742);
and U1756 (N_1756,In_2073,In_2569);
xor U1757 (N_1757,In_3978,In_1413);
nand U1758 (N_1758,In_698,In_487);
and U1759 (N_1759,In_3259,In_3110);
or U1760 (N_1760,In_1045,In_4192);
or U1761 (N_1761,In_288,In_4283);
or U1762 (N_1762,In_434,In_3006);
nor U1763 (N_1763,In_1114,In_2001);
nand U1764 (N_1764,In_815,In_302);
nor U1765 (N_1765,In_477,In_2129);
nor U1766 (N_1766,In_3823,In_3654);
nand U1767 (N_1767,In_230,In_849);
nor U1768 (N_1768,In_4674,In_773);
and U1769 (N_1769,In_1878,In_511);
nor U1770 (N_1770,In_4071,In_1091);
xor U1771 (N_1771,In_1041,In_4508);
and U1772 (N_1772,In_2171,In_1559);
or U1773 (N_1773,In_361,In_4826);
nand U1774 (N_1774,In_1615,In_2708);
and U1775 (N_1775,In_87,In_4065);
or U1776 (N_1776,In_505,In_2879);
nor U1777 (N_1777,In_1940,In_4523);
or U1778 (N_1778,In_2506,In_3484);
and U1779 (N_1779,In_1297,In_3176);
nand U1780 (N_1780,In_3575,In_2328);
nand U1781 (N_1781,In_4562,In_1531);
nand U1782 (N_1782,In_4799,In_1640);
xnor U1783 (N_1783,In_3736,In_3187);
or U1784 (N_1784,In_3706,In_4956);
or U1785 (N_1785,In_4731,In_1318);
nor U1786 (N_1786,In_941,In_8);
or U1787 (N_1787,In_1447,In_1274);
or U1788 (N_1788,In_3158,In_1692);
nor U1789 (N_1789,In_498,In_891);
nor U1790 (N_1790,In_3275,In_1019);
or U1791 (N_1791,In_4072,In_3935);
and U1792 (N_1792,In_843,In_2723);
nor U1793 (N_1793,In_4797,In_2637);
or U1794 (N_1794,In_4669,In_2852);
nand U1795 (N_1795,In_1489,In_3998);
nand U1796 (N_1796,In_598,In_1175);
nand U1797 (N_1797,In_3044,In_4685);
xor U1798 (N_1798,In_3193,In_1599);
and U1799 (N_1799,In_1731,In_1291);
nand U1800 (N_1800,In_2923,In_2133);
or U1801 (N_1801,In_1266,In_644);
and U1802 (N_1802,In_1842,In_2491);
nand U1803 (N_1803,In_2262,In_2448);
nor U1804 (N_1804,In_1879,In_1513);
and U1805 (N_1805,In_2971,In_3151);
and U1806 (N_1806,In_3107,In_2359);
xor U1807 (N_1807,In_4602,In_3783);
or U1808 (N_1808,In_2226,In_48);
nand U1809 (N_1809,In_3725,In_4954);
nor U1810 (N_1810,In_396,In_4209);
nor U1811 (N_1811,In_2736,In_3375);
nand U1812 (N_1812,In_3378,In_324);
nand U1813 (N_1813,In_1555,In_428);
xor U1814 (N_1814,In_4936,In_2212);
xor U1815 (N_1815,In_2285,In_2284);
nor U1816 (N_1816,In_4149,In_4893);
xnor U1817 (N_1817,In_1906,In_3699);
and U1818 (N_1818,In_2937,In_2559);
nor U1819 (N_1819,In_4950,In_3809);
and U1820 (N_1820,In_4533,In_1254);
xor U1821 (N_1821,In_1660,In_578);
xnor U1822 (N_1822,In_4217,In_2121);
and U1823 (N_1823,In_2070,In_2877);
and U1824 (N_1824,In_3180,In_134);
xnor U1825 (N_1825,In_4642,In_177);
and U1826 (N_1826,In_1264,In_2464);
and U1827 (N_1827,In_807,In_1754);
nand U1828 (N_1828,In_3982,In_226);
and U1829 (N_1829,In_4090,In_654);
or U1830 (N_1830,In_579,In_4934);
nand U1831 (N_1831,In_1309,In_1323);
nand U1832 (N_1832,In_1216,In_1162);
xor U1833 (N_1833,In_2369,In_492);
or U1834 (N_1834,In_4877,In_196);
nor U1835 (N_1835,In_1644,In_1573);
or U1836 (N_1836,In_91,In_2322);
nand U1837 (N_1837,In_3520,In_4184);
nand U1838 (N_1838,In_4647,In_4546);
and U1839 (N_1839,In_3735,In_3988);
nand U1840 (N_1840,In_2834,In_710);
xor U1841 (N_1841,In_1423,In_4968);
xor U1842 (N_1842,In_3374,In_4559);
xor U1843 (N_1843,In_4000,In_4786);
and U1844 (N_1844,In_4542,In_3789);
nor U1845 (N_1845,In_1726,In_1626);
xnor U1846 (N_1846,In_989,In_802);
nand U1847 (N_1847,In_1569,In_2699);
and U1848 (N_1848,In_3639,In_2930);
nand U1849 (N_1849,In_2205,In_4267);
and U1850 (N_1850,In_424,In_4726);
nand U1851 (N_1851,In_618,In_4762);
or U1852 (N_1852,In_3325,In_1876);
and U1853 (N_1853,In_61,In_4974);
nand U1854 (N_1854,In_2017,In_1522);
nand U1855 (N_1855,In_1090,In_1197);
nand U1856 (N_1856,In_3840,In_2622);
nand U1857 (N_1857,In_2036,In_2913);
or U1858 (N_1858,In_385,In_3241);
nand U1859 (N_1859,In_609,In_3041);
nor U1860 (N_1860,In_67,In_859);
nand U1861 (N_1861,In_1170,In_58);
and U1862 (N_1862,In_1851,In_3266);
xor U1863 (N_1863,In_1775,In_3711);
nor U1864 (N_1864,In_3597,In_4541);
or U1865 (N_1865,In_2119,In_4182);
nor U1866 (N_1866,In_3356,In_3070);
nor U1867 (N_1867,In_3262,In_1586);
nand U1868 (N_1868,In_3209,In_1916);
nor U1869 (N_1869,In_1328,In_3790);
xor U1870 (N_1870,In_1583,In_1483);
or U1871 (N_1871,In_4105,In_943);
nand U1872 (N_1872,In_4054,In_672);
or U1873 (N_1873,In_1171,In_1747);
nor U1874 (N_1874,In_3112,In_2718);
nand U1875 (N_1875,In_969,In_4806);
or U1876 (N_1876,In_2324,In_3637);
nor U1877 (N_1877,In_1372,In_2309);
and U1878 (N_1878,In_3831,In_46);
nor U1879 (N_1879,In_1032,In_2660);
nor U1880 (N_1880,In_4358,In_2266);
nand U1881 (N_1881,In_1004,In_2788);
nor U1882 (N_1882,In_2817,In_2495);
nand U1883 (N_1883,In_3750,In_4009);
and U1884 (N_1884,In_924,In_2775);
and U1885 (N_1885,In_3402,In_3477);
nand U1886 (N_1886,In_4298,In_3252);
and U1887 (N_1887,In_2260,In_4680);
and U1888 (N_1888,In_3065,In_2411);
or U1889 (N_1889,In_3033,In_535);
nor U1890 (N_1890,In_3930,In_3525);
nand U1891 (N_1891,In_640,In_328);
or U1892 (N_1892,In_4086,In_788);
nor U1893 (N_1893,In_2123,In_1445);
or U1894 (N_1894,In_2840,In_1166);
xor U1895 (N_1895,In_4255,In_4363);
and U1896 (N_1896,In_274,In_3532);
nand U1897 (N_1897,In_2776,In_4457);
or U1898 (N_1898,In_4539,In_2848);
or U1899 (N_1899,In_3620,In_2771);
nand U1900 (N_1900,In_2635,In_1382);
and U1901 (N_1901,In_4574,In_4061);
or U1902 (N_1902,In_3219,In_3822);
nand U1903 (N_1903,In_2850,In_4524);
and U1904 (N_1904,In_563,In_1856);
and U1905 (N_1905,In_822,In_2484);
nand U1906 (N_1906,In_2086,In_4491);
and U1907 (N_1907,In_3141,In_3526);
and U1908 (N_1908,In_3721,In_3367);
xor U1909 (N_1909,In_296,In_4834);
nor U1910 (N_1910,In_1184,In_4219);
nand U1911 (N_1911,In_2338,In_360);
or U1912 (N_1912,In_4915,In_3560);
and U1913 (N_1913,In_2833,In_971);
or U1914 (N_1914,In_1936,In_3506);
or U1915 (N_1915,In_4442,In_4250);
or U1916 (N_1916,In_2360,In_3933);
xnor U1917 (N_1917,In_4661,In_4095);
nor U1918 (N_1918,In_257,In_4240);
and U1919 (N_1919,In_4532,In_3514);
or U1920 (N_1920,In_4607,In_911);
nand U1921 (N_1921,In_4331,In_3488);
nand U1922 (N_1922,In_4403,In_3778);
or U1923 (N_1923,In_3834,In_1493);
and U1924 (N_1924,In_898,In_3035);
and U1925 (N_1925,In_133,In_2957);
nand U1926 (N_1926,In_2199,In_3553);
and U1927 (N_1927,In_116,In_737);
nand U1928 (N_1928,In_3688,In_533);
nor U1929 (N_1929,In_2009,In_1750);
nand U1930 (N_1930,In_2091,In_998);
and U1931 (N_1931,In_4340,In_102);
or U1932 (N_1932,In_893,In_653);
and U1933 (N_1933,In_4998,In_1869);
and U1934 (N_1934,In_3979,In_2347);
nor U1935 (N_1935,In_2925,In_990);
or U1936 (N_1936,In_1724,In_880);
and U1937 (N_1937,In_3068,In_3632);
nor U1938 (N_1938,In_4705,In_3047);
nand U1939 (N_1939,In_250,In_3896);
nor U1940 (N_1940,In_12,In_2902);
nand U1941 (N_1941,In_3383,In_4406);
nand U1942 (N_1942,In_805,In_3264);
xor U1943 (N_1943,In_284,In_4867);
and U1944 (N_1944,In_3166,In_2505);
nand U1945 (N_1945,In_977,In_3161);
nor U1946 (N_1946,In_2757,In_4901);
nor U1947 (N_1947,In_3591,In_901);
nand U1948 (N_1948,In_4818,In_3473);
nand U1949 (N_1949,In_4980,In_2498);
nand U1950 (N_1950,In_2687,In_164);
nor U1951 (N_1951,In_817,In_2302);
nor U1952 (N_1952,In_2535,In_1977);
nand U1953 (N_1953,In_1649,In_245);
nor U1954 (N_1954,In_4168,In_1950);
and U1955 (N_1955,In_450,In_2221);
nand U1956 (N_1956,In_2820,In_451);
or U1957 (N_1957,In_734,In_3126);
nand U1958 (N_1958,In_4987,In_1247);
nor U1959 (N_1959,In_897,In_149);
or U1960 (N_1960,In_4555,In_2985);
and U1961 (N_1961,In_2755,In_4575);
and U1962 (N_1962,In_2311,In_3843);
or U1963 (N_1963,In_3876,In_3058);
and U1964 (N_1964,In_2917,In_2344);
nand U1965 (N_1965,In_4798,In_2481);
nor U1966 (N_1966,In_152,In_2613);
nor U1967 (N_1967,In_1448,In_66);
or U1968 (N_1968,In_779,In_3195);
or U1969 (N_1969,In_2217,In_3825);
xor U1970 (N_1970,In_1742,In_375);
or U1971 (N_1971,In_2692,In_1316);
xor U1972 (N_1972,In_2548,In_632);
nand U1973 (N_1973,In_1624,In_1708);
and U1974 (N_1974,In_4486,In_2842);
and U1975 (N_1975,In_1173,In_1576);
and U1976 (N_1976,In_3805,In_2616);
xnor U1977 (N_1977,In_3739,In_561);
or U1978 (N_1978,In_1808,In_4427);
and U1979 (N_1979,In_1458,In_3746);
or U1980 (N_1980,In_3879,In_4262);
nor U1981 (N_1981,In_994,In_4012);
nand U1982 (N_1982,In_2654,In_4622);
nor U1983 (N_1983,In_235,In_1181);
and U1984 (N_1984,In_3603,In_2351);
nand U1985 (N_1985,In_1652,In_1255);
nand U1986 (N_1986,In_348,In_930);
xnor U1987 (N_1987,In_4932,In_4782);
nor U1988 (N_1988,In_804,In_2728);
or U1989 (N_1989,In_189,In_1838);
or U1990 (N_1990,In_4750,In_1883);
nand U1991 (N_1991,In_2340,In_851);
nand U1992 (N_1992,In_2578,In_26);
or U1993 (N_1993,In_2821,In_1637);
nand U1994 (N_1994,In_3972,In_2077);
and U1995 (N_1995,In_4244,In_1695);
nor U1996 (N_1996,In_2270,In_1550);
and U1997 (N_1997,In_953,In_1290);
nand U1998 (N_1998,In_3642,In_2099);
nand U1999 (N_1999,In_4274,In_2738);
and U2000 (N_2000,In_4284,In_4667);
or U2001 (N_2001,In_4692,In_41);
and U2002 (N_2002,In_110,In_5);
nor U2003 (N_2003,In_1129,In_1219);
nor U2004 (N_2004,In_3819,In_3433);
or U2005 (N_2005,In_760,In_1994);
nor U2006 (N_2006,In_4821,In_129);
nor U2007 (N_2007,In_1208,In_1052);
nor U2008 (N_2008,In_108,In_2140);
nand U2009 (N_2009,In_1600,In_1479);
nand U2010 (N_2010,In_4897,In_1852);
and U2011 (N_2011,In_1002,In_4294);
and U2012 (N_2012,In_4297,In_2294);
nand U2013 (N_2013,In_2208,In_4848);
or U2014 (N_2014,In_1207,In_4055);
nand U2015 (N_2015,In_4025,In_2408);
nand U2016 (N_2016,In_3598,In_4654);
nand U2017 (N_2017,In_516,In_3873);
or U2018 (N_2018,In_1226,In_211);
xnor U2019 (N_2019,In_123,In_786);
nor U2020 (N_2020,In_1831,In_3136);
nand U2021 (N_2021,In_2963,In_3061);
xnor U2022 (N_2022,In_2648,In_3519);
and U2023 (N_2023,In_229,In_1396);
nand U2024 (N_2024,In_1283,In_118);
nor U2025 (N_2025,In_798,In_933);
nor U2026 (N_2026,In_4557,In_856);
or U2027 (N_2027,In_3327,In_3093);
nor U2028 (N_2028,In_882,In_584);
nand U2029 (N_2029,In_370,In_3766);
and U2030 (N_2030,In_2874,In_204);
and U2031 (N_2031,In_4857,In_194);
and U2032 (N_2032,In_4317,In_1486);
and U2033 (N_2033,In_1142,In_3907);
nor U2034 (N_2034,In_2061,In_960);
and U2035 (N_2035,In_3350,In_2724);
and U2036 (N_2036,In_2507,In_2422);
and U2037 (N_2037,In_2079,In_2952);
xor U2038 (N_2038,In_1110,In_641);
or U2039 (N_2039,In_2361,In_2393);
and U2040 (N_2040,In_2126,In_4720);
xnor U2041 (N_2041,In_1788,In_1079);
xor U2042 (N_2042,In_2673,In_2472);
and U2043 (N_2043,In_2022,In_520);
or U2044 (N_2044,In_1760,In_170);
or U2045 (N_2045,In_4214,In_3959);
and U2046 (N_2046,In_2465,In_4266);
nor U2047 (N_2047,In_4470,In_140);
and U2048 (N_2048,In_3715,In_427);
nor U2049 (N_2049,In_4228,In_165);
and U2050 (N_2050,In_1671,In_3714);
and U2051 (N_2051,In_3878,In_3870);
nand U2052 (N_2052,In_925,In_2037);
or U2053 (N_2053,In_4904,In_1385);
nand U2054 (N_2054,In_2144,In_4386);
nor U2055 (N_2055,In_1011,In_829);
nor U2056 (N_2056,In_1541,In_4171);
nor U2057 (N_2057,In_2313,In_191);
and U2058 (N_2058,In_1932,In_659);
or U2059 (N_2059,In_1100,In_3038);
nand U2060 (N_2060,In_1713,In_2562);
and U2061 (N_2061,In_90,In_209);
nand U2062 (N_2062,In_799,In_2463);
nor U2063 (N_2063,In_1311,In_3090);
nor U2064 (N_2064,In_3775,In_4069);
nand U2065 (N_2065,In_1629,In_490);
and U2066 (N_2066,In_4013,In_456);
nor U2067 (N_2067,In_2783,In_583);
and U2068 (N_2068,In_3880,In_1597);
and U2069 (N_2069,In_1960,In_701);
nand U2070 (N_2070,In_4977,In_841);
nor U2071 (N_2071,In_4040,In_1776);
nor U2072 (N_2072,In_3397,In_4691);
or U2073 (N_2073,In_2709,In_4888);
nor U2074 (N_2074,In_3460,In_1193);
and U2075 (N_2075,In_2093,In_3966);
or U2076 (N_2076,In_4337,In_2901);
nand U2077 (N_2077,In_3435,In_4955);
nor U2078 (N_2078,In_4752,In_3301);
nand U2079 (N_2079,In_3529,In_1938);
and U2080 (N_2080,In_4529,In_309);
and U2081 (N_2081,In_4454,In_4721);
or U2082 (N_2082,In_2572,In_2631);
and U2083 (N_2083,In_2811,In_513);
nand U2084 (N_2084,In_1689,In_4251);
and U2085 (N_2085,In_4960,In_902);
nor U2086 (N_2086,In_749,In_241);
nor U2087 (N_2087,In_1131,In_3991);
nand U2088 (N_2088,In_3887,In_1735);
or U2089 (N_2089,In_9,In_4151);
nor U2090 (N_2090,In_127,In_71);
nor U2091 (N_2091,In_796,In_2346);
and U2092 (N_2092,In_421,In_1952);
xnor U2093 (N_2093,In_390,In_3918);
and U2094 (N_2094,In_775,In_1098);
nand U2095 (N_2095,In_2012,In_4080);
xor U2096 (N_2096,In_504,In_3983);
nor U2097 (N_2097,In_4755,In_787);
or U2098 (N_2098,In_2870,In_1699);
xnor U2099 (N_2099,In_4513,In_1121);
and U2100 (N_2100,In_1094,In_1602);
or U2101 (N_2101,In_2735,In_3931);
nor U2102 (N_2102,In_3534,In_3665);
and U2103 (N_2103,In_545,In_4387);
nand U2104 (N_2104,In_676,In_286);
or U2105 (N_2105,In_2455,In_60);
or U2106 (N_2106,In_4842,In_1178);
or U2107 (N_2107,In_2297,In_1367);
nor U2108 (N_2108,In_4241,In_3767);
nor U2109 (N_2109,In_4839,In_4990);
nand U2110 (N_2110,In_2175,In_2688);
nand U2111 (N_2111,In_4114,In_582);
or U2112 (N_2112,In_479,In_3507);
and U2113 (N_2113,In_1584,In_1792);
nand U2114 (N_2114,In_1482,In_4425);
or U2115 (N_2115,In_2526,In_2867);
nand U2116 (N_2116,In_867,In_4144);
nand U2117 (N_2117,In_2966,In_1546);
or U2118 (N_2118,In_982,In_1083);
nand U2119 (N_2119,In_181,In_2471);
or U2120 (N_2120,In_794,In_179);
nand U2121 (N_2121,In_3343,In_692);
or U2122 (N_2122,In_4883,In_675);
or U2123 (N_2123,In_275,In_2078);
nor U2124 (N_2124,In_2138,In_3363);
nand U2125 (N_2125,In_2706,In_3932);
and U2126 (N_2126,In_1005,In_1150);
nor U2127 (N_2127,In_2141,In_4310);
nor U2128 (N_2128,In_1192,In_695);
and U2129 (N_2129,In_1384,In_4276);
nand U2130 (N_2130,In_1995,In_1791);
nand U2131 (N_2131,In_2004,In_3496);
nand U2132 (N_2132,In_290,In_835);
xor U2133 (N_2133,In_3293,In_643);
and U2134 (N_2134,In_2960,In_1832);
and U2135 (N_2135,In_1152,In_3020);
nand U2136 (N_2136,In_1018,In_2598);
nand U2137 (N_2137,In_2057,In_166);
xnor U2138 (N_2138,In_2128,In_3246);
or U2139 (N_2139,In_1965,In_3189);
nor U2140 (N_2140,In_4549,In_162);
or U2141 (N_2141,In_596,In_4736);
or U2142 (N_2142,In_1159,In_3686);
nand U2143 (N_2143,In_4741,In_2809);
and U2144 (N_2144,In_3826,In_2536);
nor U2145 (N_2145,In_1730,In_4604);
or U2146 (N_2146,In_4766,In_3955);
nor U2147 (N_2147,In_1063,In_3102);
and U2148 (N_2148,In_3026,In_1784);
nand U2149 (N_2149,In_3986,In_1463);
or U2150 (N_2150,In_1155,In_751);
nand U2151 (N_2151,In_214,In_1635);
nor U2152 (N_2152,In_135,In_4645);
nor U2153 (N_2153,In_3258,In_2510);
nor U2154 (N_2154,In_2555,In_4469);
or U2155 (N_2155,In_82,In_146);
or U2156 (N_2156,In_707,In_3543);
xor U2157 (N_2157,In_3022,In_4837);
nand U2158 (N_2158,In_2223,In_1242);
or U2159 (N_2159,In_1672,In_2741);
nand U2160 (N_2160,In_1380,In_1528);
and U2161 (N_2161,In_1538,In_2798);
nand U2162 (N_2162,In_3936,In_238);
nor U2163 (N_2163,In_3270,In_4903);
or U2164 (N_2164,In_1340,In_4565);
or U2165 (N_2165,In_2640,In_4617);
xor U2166 (N_2166,In_2626,In_2069);
or U2167 (N_2167,In_1329,In_4616);
nor U2168 (N_2168,In_3424,In_515);
nor U2169 (N_2169,In_4271,In_64);
nand U2170 (N_2170,In_2995,In_1249);
xor U2171 (N_2171,In_4133,In_3886);
nand U2172 (N_2172,In_4701,In_1067);
nand U2173 (N_2173,In_1010,In_4601);
or U2174 (N_2174,In_1577,In_4);
and U2175 (N_2175,In_3116,In_4869);
or U2176 (N_2176,In_4913,In_647);
xor U2177 (N_2177,In_3798,In_2186);
or U2178 (N_2178,In_3653,In_2490);
or U2179 (N_2179,In_1221,In_3427);
xnor U2180 (N_2180,In_2489,In_2804);
nand U2181 (N_2181,In_252,In_1084);
nor U2182 (N_2182,In_353,In_2727);
and U2183 (N_2183,In_99,In_1609);
and U2184 (N_2184,In_4067,In_425);
and U2185 (N_2185,In_3461,In_538);
or U2186 (N_2186,In_4658,In_4052);
or U2187 (N_2187,In_2516,In_3612);
and U2188 (N_2188,In_3319,In_2276);
or U2189 (N_2189,In_1805,In_2365);
nor U2190 (N_2190,In_3489,In_4759);
nor U2191 (N_2191,In_626,In_2014);
and U2192 (N_2192,In_3442,In_1963);
xnor U2193 (N_2193,In_207,In_604);
and U2194 (N_2194,In_2967,In_2826);
and U2195 (N_2195,In_3311,In_125);
and U2196 (N_2196,In_4224,In_4057);
nand U2197 (N_2197,In_864,In_1373);
and U2198 (N_2198,In_1565,In_610);
and U2199 (N_2199,In_1059,In_573);
or U2200 (N_2200,In_341,In_2143);
nor U2201 (N_2201,In_4191,In_2596);
nor U2202 (N_2202,In_3681,In_1130);
xor U2203 (N_2203,In_4099,In_4871);
nand U2204 (N_2204,In_839,In_2406);
or U2205 (N_2205,In_29,In_4170);
nand U2206 (N_2206,In_886,In_812);
and U2207 (N_2207,In_4421,In_3498);
or U2208 (N_2208,In_1705,In_199);
nand U2209 (N_2209,In_4324,In_1741);
or U2210 (N_2210,In_3578,In_2665);
or U2211 (N_2211,In_2979,In_3372);
nor U2212 (N_2212,In_2503,In_3013);
xor U2213 (N_2213,In_2250,In_4709);
nor U2214 (N_2214,In_4146,In_2043);
or U2215 (N_2215,In_4924,In_1322);
nor U2216 (N_2216,In_4211,In_4415);
nand U2217 (N_2217,In_3941,In_772);
nor U2218 (N_2218,In_797,In_762);
and U2219 (N_2219,In_3796,In_4666);
nand U2220 (N_2220,In_3137,In_4236);
nor U2221 (N_2221,In_4202,In_2761);
and U2222 (N_2222,In_3029,In_3634);
nor U2223 (N_2223,In_4943,In_1440);
or U2224 (N_2224,In_1244,In_4996);
or U2225 (N_2225,In_3289,In_4377);
nor U2226 (N_2226,In_1118,In_4598);
nand U2227 (N_2227,In_4620,In_3924);
nor U2228 (N_2228,In_3538,In_3564);
xor U2229 (N_2229,In_4820,In_2384);
and U2230 (N_2230,In_4413,In_542);
and U2231 (N_2231,In_3453,In_4008);
and U2232 (N_2232,In_544,In_3015);
or U2233 (N_2233,In_163,In_1459);
and U2234 (N_2234,In_912,In_2225);
and U2235 (N_2235,In_3073,In_4600);
nor U2236 (N_2236,In_1738,In_3600);
xnor U2237 (N_2237,In_3695,In_4650);
or U2238 (N_2238,In_4817,In_765);
or U2239 (N_2239,In_3482,In_1976);
or U2240 (N_2240,In_402,In_3760);
or U2241 (N_2241,In_1401,In_1205);
or U2242 (N_2242,In_2531,In_268);
and U2243 (N_2243,In_2911,In_1186);
or U2244 (N_2244,In_3046,In_1191);
xnor U2245 (N_2245,In_705,In_1215);
or U2246 (N_2246,In_683,In_4302);
or U2247 (N_2247,In_4125,In_2747);
nor U2248 (N_2248,In_3320,In_322);
nand U2249 (N_2249,In_2655,In_2030);
or U2250 (N_2250,In_2124,In_2586);
xor U2251 (N_2251,In_3548,In_1154);
and U2252 (N_2252,In_2745,In_1066);
and U2253 (N_2253,In_1354,In_1801);
or U2254 (N_2254,In_2237,In_4315);
xnor U2255 (N_2255,In_3623,In_2219);
or U2256 (N_2256,In_3119,In_4476);
xnor U2257 (N_2257,In_2885,In_1351);
or U2258 (N_2258,In_473,In_1040);
nor U2259 (N_2259,In_863,In_4745);
nor U2260 (N_2260,In_869,In_486);
nand U2261 (N_2261,In_2595,In_2218);
xnor U2262 (N_2262,In_548,In_3626);
and U2263 (N_2263,In_2994,In_344);
nor U2264 (N_2264,In_3348,In_319);
nor U2265 (N_2265,In_1501,In_702);
nand U2266 (N_2266,In_4070,In_3410);
nand U2267 (N_2267,In_4597,In_1081);
or U2268 (N_2268,In_1361,In_3592);
or U2269 (N_2269,In_2946,In_4451);
xor U2270 (N_2270,In_539,In_523);
or U2271 (N_2271,In_3024,In_4623);
or U2272 (N_2272,In_4152,In_2215);
nor U2273 (N_2273,In_2525,In_1667);
nor U2274 (N_2274,In_202,In_4073);
nor U2275 (N_2275,In_1112,In_1743);
nand U2276 (N_2276,In_868,In_96);
nand U2277 (N_2277,In_3145,In_3223);
nor U2278 (N_2278,In_1103,In_3864);
or U2279 (N_2279,In_854,In_3939);
or U2280 (N_2280,In_3551,In_299);
nor U2281 (N_2281,In_1415,In_3868);
xnor U2282 (N_2282,In_935,In_4715);
nand U2283 (N_2283,In_4367,In_2753);
nand U2284 (N_2284,In_3556,In_1167);
nand U2285 (N_2285,In_198,In_975);
nor U2286 (N_2286,In_3037,In_3148);
xnor U2287 (N_2287,In_870,In_1850);
and U2288 (N_2288,In_3302,In_663);
and U2289 (N_2289,In_3938,In_3547);
nand U2290 (N_2290,In_1341,In_3009);
or U2291 (N_2291,In_1658,In_541);
nand U2292 (N_2292,In_3605,In_2428);
nand U2293 (N_2293,In_3663,In_2233);
and U2294 (N_2294,In_3236,In_3807);
nand U2295 (N_2295,In_357,In_1844);
and U2296 (N_2296,In_1868,In_942);
and U2297 (N_2297,In_1700,In_2864);
xor U2298 (N_2298,In_206,In_4215);
nand U2299 (N_2299,In_2184,In_679);
or U2300 (N_2300,In_3441,In_1492);
and U2301 (N_2301,In_877,In_1718);
nand U2302 (N_2302,In_2301,In_2560);
nand U2303 (N_2303,In_4632,In_62);
nand U2304 (N_2304,In_1662,In_2746);
nand U2305 (N_2305,In_4381,In_1300);
or U2306 (N_2306,In_4895,In_3017);
or U2307 (N_2307,In_1267,In_2349);
and U2308 (N_2308,In_4558,In_619);
nand U2309 (N_2309,In_2013,In_355);
nand U2310 (N_2310,In_1895,In_2717);
nand U2311 (N_2311,In_264,In_4580);
nor U2312 (N_2312,In_3934,In_3314);
and U2313 (N_2313,In_629,In_4880);
nand U2314 (N_2314,In_1347,In_3224);
and U2315 (N_2315,In_2549,In_2829);
or U2316 (N_2316,In_3390,In_3312);
and U2317 (N_2317,In_2029,In_101);
nor U2318 (N_2318,In_4440,In_2174);
nand U2319 (N_2319,In_3683,In_2905);
or U2320 (N_2320,In_549,In_2533);
and U2321 (N_2321,In_2567,In_2799);
nand U2322 (N_2322,In_4326,In_3867);
nor U2323 (N_2323,In_1099,In_3762);
nor U2324 (N_2324,In_4158,In_3850);
nor U2325 (N_2325,In_2331,In_3457);
nor U2326 (N_2326,In_1306,In_4849);
nor U2327 (N_2327,In_752,In_4281);
nor U2328 (N_2328,In_1048,In_1757);
and U2329 (N_2329,In_3413,In_3855);
and U2330 (N_2330,In_1627,In_2337);
xor U2331 (N_2331,In_4369,In_1864);
and U2332 (N_2332,In_3133,In_1024);
or U2333 (N_2333,In_2721,In_3202);
nand U2334 (N_2334,In_4388,In_3192);
and U2335 (N_2335,In_1621,In_2552);
nor U2336 (N_2336,In_3463,In_4564);
nor U2337 (N_2337,In_151,In_2632);
xnor U2338 (N_2338,In_1509,In_3869);
xnor U2339 (N_2339,In_3567,In_2210);
nand U2340 (N_2340,In_1364,In_795);
nor U2341 (N_2341,In_4081,In_305);
and U2342 (N_2342,In_642,In_1331);
and U2343 (N_2343,In_4197,In_374);
nand U2344 (N_2344,In_124,In_3696);
nand U2345 (N_2345,In_3198,In_3646);
nor U2346 (N_2346,In_3296,In_735);
or U2347 (N_2347,In_1843,In_2661);
and U2348 (N_2348,In_1811,In_1582);
and U2349 (N_2349,In_4890,In_85);
nor U2350 (N_2350,In_2397,In_1873);
and U2351 (N_2351,In_4408,In_3355);
or U2352 (N_2352,In_4494,In_2383);
xnor U2353 (N_2353,In_1958,In_1618);
and U2354 (N_2354,In_4699,In_4711);
nand U2355 (N_2355,In_1812,In_1195);
nand U2356 (N_2356,In_1847,In_4679);
or U2357 (N_2357,In_3606,In_4560);
or U2358 (N_2358,In_755,In_3925);
nand U2359 (N_2359,In_2731,In_2542);
or U2360 (N_2360,In_4931,In_4288);
nand U2361 (N_2361,In_4732,In_4027);
and U2362 (N_2362,In_3040,In_4930);
xnor U2363 (N_2363,In_219,In_4289);
or U2364 (N_2364,In_4245,In_1946);
and U2365 (N_2365,In_3602,In_481);
nand U2366 (N_2366,In_2169,In_661);
nor U2367 (N_2367,In_2607,In_4438);
and U2368 (N_2368,In_265,In_4051);
and U2369 (N_2369,In_4424,In_2315);
and U2370 (N_2370,In_2149,In_855);
or U2371 (N_2371,In_3812,In_2020);
nand U2372 (N_2372,In_1779,In_879);
xnor U2373 (N_2373,In_4347,In_4949);
nor U2374 (N_2374,In_1948,In_4671);
nor U2375 (N_2375,In_314,In_1431);
and U2376 (N_2376,In_3513,In_1712);
and U2377 (N_2377,In_914,In_4805);
and U2378 (N_2378,In_4649,In_1782);
or U2379 (N_2379,In_2707,In_59);
or U2380 (N_2380,In_2380,In_3391);
nand U2381 (N_2381,In_1553,In_1681);
xor U2382 (N_2382,In_2846,In_3469);
or U2383 (N_2383,In_3140,In_4690);
or U2384 (N_2384,In_2164,In_3257);
nand U2385 (N_2385,In_2442,In_484);
and U2386 (N_2386,In_3586,In_4618);
or U2387 (N_2387,In_2803,In_218);
or U2388 (N_2388,In_2172,In_1841);
and U2389 (N_2389,In_2941,In_53);
nor U2390 (N_2390,In_2355,In_3884);
xnor U2391 (N_2391,In_1687,In_4412);
nand U2392 (N_2392,In_1571,In_3515);
xor U2393 (N_2393,In_4520,In_1751);
xnor U2394 (N_2394,In_670,In_227);
nor U2395 (N_2395,In_3601,In_3228);
and U2396 (N_2396,In_4050,In_141);
nor U2397 (N_2397,In_2896,In_591);
or U2398 (N_2398,In_1954,In_4836);
and U2399 (N_2399,In_3185,In_4822);
xor U2400 (N_2400,In_4795,In_4385);
or U2401 (N_2401,In_3786,In_2825);
and U2402 (N_2402,In_593,In_1570);
and U2403 (N_2403,In_2390,In_3573);
or U2404 (N_2404,In_4854,In_1557);
and U2405 (N_2405,In_45,In_4586);
xor U2406 (N_2406,In_4321,In_4233);
nand U2407 (N_2407,In_4094,In_2556);
nor U2408 (N_2408,In_3366,In_1346);
or U2409 (N_2409,In_4429,In_4097);
nor U2410 (N_2410,In_1659,In_4803);
nand U2411 (N_2411,In_79,In_393);
and U2412 (N_2412,In_1089,In_3415);
nor U2413 (N_2413,In_4695,In_1168);
and U2414 (N_2414,In_881,In_1258);
and U2415 (N_2415,In_4937,In_2446);
nand U2416 (N_2416,In_2573,In_2071);
xnor U2417 (N_2417,In_4984,In_2704);
xnor U2418 (N_2418,In_2694,In_4999);
nor U2419 (N_2419,In_4994,In_2368);
nand U2420 (N_2420,In_2912,In_3844);
nand U2421 (N_2421,In_1451,In_4694);
xnor U2422 (N_2422,In_3446,In_1890);
nor U2423 (N_2423,In_3927,In_1286);
nand U2424 (N_2424,In_1488,In_1925);
nor U2425 (N_2425,In_3788,In_1027);
or U2426 (N_2426,In_4428,In_4137);
xnor U2427 (N_2427,In_4436,In_4291);
nor U2428 (N_2428,In_1036,In_2296);
nor U2429 (N_2429,In_3949,In_4048);
nor U2430 (N_2430,In_3448,In_4516);
nor U2431 (N_2431,In_931,In_1732);
xor U2432 (N_2432,In_996,In_4770);
or U2433 (N_2433,In_2483,In_1787);
or U2434 (N_2434,In_837,In_4522);
and U2435 (N_2435,In_1023,In_3638);
or U2436 (N_2436,In_1210,In_2610);
or U2437 (N_2437,In_70,In_294);
nand U2438 (N_2438,In_187,In_1232);
nand U2439 (N_2439,In_4724,In_2278);
nand U2440 (N_2440,In_2831,In_467);
or U2441 (N_2441,In_3458,In_1806);
nand U2442 (N_2442,In_4077,In_1516);
xnor U2443 (N_2443,In_3643,In_1756);
and U2444 (N_2444,In_1737,In_2892);
nor U2445 (N_2445,In_1206,In_2430);
nor U2446 (N_2446,In_3923,In_1717);
or U2447 (N_2447,In_660,In_1585);
nand U2448 (N_2448,In_2178,In_3613);
nand U2449 (N_2449,In_4688,In_4905);
or U2450 (N_2450,In_1545,In_3572);
and U2451 (N_2451,In_4155,In_4329);
and U2452 (N_2452,In_343,In_531);
nand U2453 (N_2453,In_4495,In_1395);
or U2454 (N_2454,In_1243,In_2427);
xor U2455 (N_2455,In_667,In_4595);
nand U2456 (N_2456,In_1663,In_3207);
xor U2457 (N_2457,In_2524,In_3168);
xnor U2458 (N_2458,In_3702,In_2993);
or U2459 (N_2459,In_2649,In_4119);
nor U2460 (N_2460,In_3829,In_1665);
and U2461 (N_2461,In_3689,In_139);
nor U2462 (N_2462,In_3508,In_2808);
nand U2463 (N_2463,In_3516,In_4349);
or U2464 (N_2464,In_3349,In_362);
nor U2465 (N_2465,In_1796,In_37);
or U2466 (N_2466,In_2474,In_4933);
or U2467 (N_2467,In_3132,In_4938);
or U2468 (N_2468,In_50,In_4677);
and U2469 (N_2469,In_2793,In_638);
or U2470 (N_2470,In_3491,In_1562);
nand U2471 (N_2471,In_981,In_2628);
and U2472 (N_2472,In_602,In_1601);
nor U2473 (N_2473,In_501,In_2467);
nor U2474 (N_2474,In_3276,In_4235);
nand U2475 (N_2475,In_889,In_4708);
nor U2476 (N_2476,In_2585,In_3108);
nor U2477 (N_2477,In_2903,In_4404);
nand U2478 (N_2478,In_3859,In_2357);
nor U2479 (N_2479,In_3997,In_208);
nor U2480 (N_2480,In_2715,In_2855);
nor U2481 (N_2481,In_2421,In_4220);
nand U2482 (N_2482,In_1736,In_2034);
nand U2483 (N_2483,In_2485,In_4872);
and U2484 (N_2484,In_3678,In_213);
and U2485 (N_2485,In_2678,In_4122);
nand U2486 (N_2486,In_4918,In_1424);
and U2487 (N_2487,In_3271,In_4312);
nor U2488 (N_2488,In_2112,In_2229);
and U2489 (N_2489,In_3861,In_2695);
and U2490 (N_2490,In_154,In_1022);
or U2491 (N_2491,In_232,In_1786);
and U2492 (N_2492,In_3737,In_4181);
xnor U2493 (N_2493,In_4874,In_1064);
xnor U2494 (N_2494,In_961,In_416);
or U2495 (N_2495,In_1204,In_920);
or U2496 (N_2496,In_769,In_2791);
nor U2497 (N_2497,In_4912,In_3965);
and U2498 (N_2498,In_1903,In_3368);
or U2499 (N_2499,In_243,In_4717);
or U2500 (N_2500,In_2714,In_1181);
and U2501 (N_2501,In_4237,In_3672);
or U2502 (N_2502,In_4896,In_3263);
and U2503 (N_2503,In_3480,In_66);
or U2504 (N_2504,In_4754,In_117);
nand U2505 (N_2505,In_3259,In_4914);
and U2506 (N_2506,In_4934,In_1673);
or U2507 (N_2507,In_1274,In_2842);
and U2508 (N_2508,In_4300,In_3781);
and U2509 (N_2509,In_2136,In_2439);
nor U2510 (N_2510,In_213,In_1946);
and U2511 (N_2511,In_3562,In_568);
or U2512 (N_2512,In_770,In_4626);
nor U2513 (N_2513,In_1904,In_3107);
xnor U2514 (N_2514,In_2955,In_1027);
nor U2515 (N_2515,In_3215,In_3674);
or U2516 (N_2516,In_3689,In_2223);
nand U2517 (N_2517,In_4251,In_4830);
nand U2518 (N_2518,In_4021,In_1952);
or U2519 (N_2519,In_416,In_4235);
nor U2520 (N_2520,In_597,In_1039);
and U2521 (N_2521,In_3937,In_2332);
and U2522 (N_2522,In_4148,In_3655);
nor U2523 (N_2523,In_1868,In_296);
and U2524 (N_2524,In_4052,In_3456);
xor U2525 (N_2525,In_3609,In_4872);
xnor U2526 (N_2526,In_3960,In_2116);
nand U2527 (N_2527,In_1642,In_105);
or U2528 (N_2528,In_1793,In_2230);
or U2529 (N_2529,In_1593,In_294);
nor U2530 (N_2530,In_890,In_4745);
nand U2531 (N_2531,In_2771,In_2266);
and U2532 (N_2532,In_2029,In_3042);
or U2533 (N_2533,In_3162,In_1107);
or U2534 (N_2534,In_1997,In_1825);
and U2535 (N_2535,In_3626,In_813);
nor U2536 (N_2536,In_3982,In_4347);
and U2537 (N_2537,In_56,In_4490);
nor U2538 (N_2538,In_4209,In_3754);
and U2539 (N_2539,In_4848,In_1379);
and U2540 (N_2540,In_2530,In_1601);
and U2541 (N_2541,In_3290,In_4629);
nand U2542 (N_2542,In_2587,In_637);
or U2543 (N_2543,In_535,In_4822);
and U2544 (N_2544,In_1552,In_3377);
nor U2545 (N_2545,In_3789,In_4421);
nand U2546 (N_2546,In_3501,In_3007);
nor U2547 (N_2547,In_2055,In_4335);
and U2548 (N_2548,In_2460,In_1352);
or U2549 (N_2549,In_2684,In_2473);
nand U2550 (N_2550,In_2304,In_616);
and U2551 (N_2551,In_2455,In_984);
and U2552 (N_2552,In_1836,In_4705);
and U2553 (N_2553,In_3183,In_4670);
xor U2554 (N_2554,In_727,In_2646);
nand U2555 (N_2555,In_320,In_627);
nor U2556 (N_2556,In_2448,In_3478);
and U2557 (N_2557,In_4489,In_3006);
and U2558 (N_2558,In_3493,In_1387);
nand U2559 (N_2559,In_1434,In_3322);
nor U2560 (N_2560,In_3553,In_653);
xnor U2561 (N_2561,In_1610,In_2043);
nor U2562 (N_2562,In_1364,In_2599);
or U2563 (N_2563,In_1002,In_2721);
and U2564 (N_2564,In_1502,In_335);
nor U2565 (N_2565,In_2151,In_27);
or U2566 (N_2566,In_1687,In_4077);
and U2567 (N_2567,In_1340,In_89);
and U2568 (N_2568,In_2988,In_4168);
xor U2569 (N_2569,In_3558,In_4740);
nand U2570 (N_2570,In_3091,In_2047);
and U2571 (N_2571,In_1335,In_3382);
xor U2572 (N_2572,In_4022,In_3702);
nor U2573 (N_2573,In_3955,In_4883);
xnor U2574 (N_2574,In_1386,In_926);
or U2575 (N_2575,In_1506,In_2238);
nand U2576 (N_2576,In_4910,In_191);
nor U2577 (N_2577,In_2912,In_1776);
nand U2578 (N_2578,In_4376,In_1131);
xnor U2579 (N_2579,In_2860,In_1335);
nand U2580 (N_2580,In_1915,In_969);
nand U2581 (N_2581,In_3242,In_2433);
nand U2582 (N_2582,In_4974,In_4273);
nand U2583 (N_2583,In_3457,In_2155);
xnor U2584 (N_2584,In_1492,In_3772);
and U2585 (N_2585,In_757,In_4502);
nor U2586 (N_2586,In_2813,In_2211);
and U2587 (N_2587,In_3959,In_3522);
and U2588 (N_2588,In_2924,In_4307);
nand U2589 (N_2589,In_1693,In_1874);
and U2590 (N_2590,In_4903,In_2901);
nor U2591 (N_2591,In_173,In_2322);
and U2592 (N_2592,In_2608,In_2052);
nor U2593 (N_2593,In_3860,In_4525);
and U2594 (N_2594,In_4631,In_2613);
or U2595 (N_2595,In_1479,In_4539);
nor U2596 (N_2596,In_50,In_446);
or U2597 (N_2597,In_2474,In_4248);
nor U2598 (N_2598,In_1140,In_2373);
and U2599 (N_2599,In_4071,In_1344);
nor U2600 (N_2600,In_2655,In_173);
nand U2601 (N_2601,In_3064,In_3009);
nand U2602 (N_2602,In_2312,In_1);
nand U2603 (N_2603,In_1559,In_2816);
nor U2604 (N_2604,In_2607,In_4604);
and U2605 (N_2605,In_4819,In_638);
nor U2606 (N_2606,In_769,In_4563);
or U2607 (N_2607,In_4933,In_105);
and U2608 (N_2608,In_105,In_1972);
nor U2609 (N_2609,In_2433,In_838);
and U2610 (N_2610,In_958,In_556);
nor U2611 (N_2611,In_3575,In_3989);
and U2612 (N_2612,In_363,In_2937);
nand U2613 (N_2613,In_320,In_1573);
nor U2614 (N_2614,In_1944,In_3656);
nand U2615 (N_2615,In_3261,In_4764);
and U2616 (N_2616,In_4978,In_4785);
or U2617 (N_2617,In_1004,In_3971);
nor U2618 (N_2618,In_3970,In_2338);
or U2619 (N_2619,In_4390,In_1068);
and U2620 (N_2620,In_3383,In_3743);
or U2621 (N_2621,In_1421,In_4106);
or U2622 (N_2622,In_3627,In_2703);
nor U2623 (N_2623,In_3767,In_4770);
or U2624 (N_2624,In_4645,In_1081);
xor U2625 (N_2625,In_3091,In_4812);
nor U2626 (N_2626,In_4806,In_1330);
and U2627 (N_2627,In_1544,In_2719);
nand U2628 (N_2628,In_830,In_4616);
xor U2629 (N_2629,In_2809,In_4890);
or U2630 (N_2630,In_1996,In_1843);
and U2631 (N_2631,In_2059,In_4433);
nand U2632 (N_2632,In_4382,In_4136);
and U2633 (N_2633,In_1144,In_259);
xnor U2634 (N_2634,In_2156,In_751);
or U2635 (N_2635,In_1943,In_701);
nor U2636 (N_2636,In_4890,In_3796);
nand U2637 (N_2637,In_348,In_773);
and U2638 (N_2638,In_2139,In_2877);
nand U2639 (N_2639,In_4367,In_2998);
nor U2640 (N_2640,In_3341,In_920);
and U2641 (N_2641,In_4778,In_3081);
and U2642 (N_2642,In_2385,In_2189);
and U2643 (N_2643,In_1977,In_4517);
nand U2644 (N_2644,In_3887,In_1019);
nor U2645 (N_2645,In_949,In_2487);
or U2646 (N_2646,In_666,In_1934);
or U2647 (N_2647,In_2106,In_1756);
and U2648 (N_2648,In_4787,In_486);
nand U2649 (N_2649,In_2607,In_4367);
or U2650 (N_2650,In_1464,In_3666);
xor U2651 (N_2651,In_2085,In_1238);
or U2652 (N_2652,In_1884,In_3232);
xnor U2653 (N_2653,In_1144,In_189);
xnor U2654 (N_2654,In_826,In_417);
nand U2655 (N_2655,In_2303,In_4276);
nand U2656 (N_2656,In_341,In_1101);
and U2657 (N_2657,In_626,In_231);
and U2658 (N_2658,In_2927,In_134);
or U2659 (N_2659,In_1436,In_689);
nor U2660 (N_2660,In_4746,In_757);
or U2661 (N_2661,In_3812,In_1621);
nand U2662 (N_2662,In_2007,In_1505);
or U2663 (N_2663,In_1554,In_2004);
or U2664 (N_2664,In_1106,In_3097);
nand U2665 (N_2665,In_582,In_2267);
and U2666 (N_2666,In_1340,In_4323);
nand U2667 (N_2667,In_1764,In_916);
nand U2668 (N_2668,In_111,In_3427);
and U2669 (N_2669,In_2120,In_3137);
xor U2670 (N_2670,In_2306,In_1233);
or U2671 (N_2671,In_2669,In_2392);
and U2672 (N_2672,In_2891,In_1038);
or U2673 (N_2673,In_1781,In_3162);
and U2674 (N_2674,In_1611,In_2685);
and U2675 (N_2675,In_1909,In_3862);
xor U2676 (N_2676,In_545,In_4315);
nand U2677 (N_2677,In_2791,In_779);
nor U2678 (N_2678,In_1697,In_4032);
or U2679 (N_2679,In_4922,In_511);
and U2680 (N_2680,In_4924,In_4111);
nor U2681 (N_2681,In_1815,In_1285);
nand U2682 (N_2682,In_287,In_909);
or U2683 (N_2683,In_1876,In_4842);
nand U2684 (N_2684,In_2205,In_2299);
xor U2685 (N_2685,In_3406,In_3098);
nor U2686 (N_2686,In_4148,In_474);
and U2687 (N_2687,In_2444,In_2406);
nand U2688 (N_2688,In_1768,In_3689);
nand U2689 (N_2689,In_2058,In_1042);
or U2690 (N_2690,In_3012,In_160);
or U2691 (N_2691,In_4910,In_4336);
nand U2692 (N_2692,In_3176,In_3195);
or U2693 (N_2693,In_1028,In_2766);
nor U2694 (N_2694,In_1668,In_4161);
nor U2695 (N_2695,In_2015,In_4014);
or U2696 (N_2696,In_1258,In_4694);
and U2697 (N_2697,In_4052,In_1223);
or U2698 (N_2698,In_84,In_3109);
and U2699 (N_2699,In_1600,In_422);
and U2700 (N_2700,In_3259,In_2561);
and U2701 (N_2701,In_910,In_1584);
nand U2702 (N_2702,In_4971,In_4775);
or U2703 (N_2703,In_1375,In_2574);
and U2704 (N_2704,In_3542,In_1802);
nor U2705 (N_2705,In_1890,In_4535);
nand U2706 (N_2706,In_3994,In_2595);
nand U2707 (N_2707,In_2310,In_179);
and U2708 (N_2708,In_3589,In_2859);
xnor U2709 (N_2709,In_4101,In_4668);
nor U2710 (N_2710,In_2073,In_3898);
and U2711 (N_2711,In_4978,In_1177);
nor U2712 (N_2712,In_753,In_4033);
or U2713 (N_2713,In_4602,In_4663);
or U2714 (N_2714,In_1682,In_2471);
and U2715 (N_2715,In_3023,In_2946);
and U2716 (N_2716,In_1273,In_3571);
nor U2717 (N_2717,In_3638,In_4528);
and U2718 (N_2718,In_422,In_1807);
or U2719 (N_2719,In_1941,In_4585);
or U2720 (N_2720,In_2003,In_3014);
or U2721 (N_2721,In_936,In_3884);
or U2722 (N_2722,In_2274,In_4081);
nor U2723 (N_2723,In_1119,In_4613);
nand U2724 (N_2724,In_4380,In_325);
or U2725 (N_2725,In_3760,In_1995);
and U2726 (N_2726,In_34,In_1856);
and U2727 (N_2727,In_741,In_565);
and U2728 (N_2728,In_576,In_168);
nand U2729 (N_2729,In_3838,In_3268);
nand U2730 (N_2730,In_4350,In_4825);
and U2731 (N_2731,In_847,In_2032);
and U2732 (N_2732,In_1602,In_14);
nand U2733 (N_2733,In_1865,In_1586);
and U2734 (N_2734,In_4336,In_366);
xnor U2735 (N_2735,In_4905,In_4873);
nand U2736 (N_2736,In_3660,In_56);
xnor U2737 (N_2737,In_1519,In_3416);
xnor U2738 (N_2738,In_3393,In_4797);
nand U2739 (N_2739,In_4661,In_2416);
nor U2740 (N_2740,In_3452,In_2335);
nor U2741 (N_2741,In_3975,In_3130);
xnor U2742 (N_2742,In_4777,In_2367);
and U2743 (N_2743,In_2150,In_3532);
and U2744 (N_2744,In_4336,In_2682);
nand U2745 (N_2745,In_2070,In_2933);
xnor U2746 (N_2746,In_408,In_89);
or U2747 (N_2747,In_710,In_3404);
nor U2748 (N_2748,In_1717,In_964);
or U2749 (N_2749,In_3830,In_3465);
nor U2750 (N_2750,In_2209,In_608);
nor U2751 (N_2751,In_978,In_1181);
nor U2752 (N_2752,In_4182,In_2813);
nand U2753 (N_2753,In_1326,In_2553);
nor U2754 (N_2754,In_1434,In_3238);
and U2755 (N_2755,In_3958,In_283);
nor U2756 (N_2756,In_590,In_3654);
nor U2757 (N_2757,In_3329,In_4352);
nor U2758 (N_2758,In_3862,In_2688);
and U2759 (N_2759,In_3584,In_1811);
xnor U2760 (N_2760,In_955,In_4651);
or U2761 (N_2761,In_3493,In_622);
and U2762 (N_2762,In_3765,In_1832);
nor U2763 (N_2763,In_181,In_806);
nor U2764 (N_2764,In_4649,In_405);
or U2765 (N_2765,In_1493,In_1264);
and U2766 (N_2766,In_3871,In_2554);
nor U2767 (N_2767,In_1953,In_264);
or U2768 (N_2768,In_3559,In_943);
nand U2769 (N_2769,In_2755,In_4511);
or U2770 (N_2770,In_3947,In_1458);
nor U2771 (N_2771,In_3758,In_4415);
or U2772 (N_2772,In_3762,In_3675);
or U2773 (N_2773,In_292,In_2115);
and U2774 (N_2774,In_791,In_1052);
and U2775 (N_2775,In_2374,In_2187);
or U2776 (N_2776,In_1017,In_3721);
nor U2777 (N_2777,In_3934,In_3981);
and U2778 (N_2778,In_4947,In_4233);
or U2779 (N_2779,In_2469,In_297);
xor U2780 (N_2780,In_684,In_4276);
nand U2781 (N_2781,In_706,In_3553);
nand U2782 (N_2782,In_1776,In_358);
nor U2783 (N_2783,In_108,In_3236);
nand U2784 (N_2784,In_1032,In_2330);
and U2785 (N_2785,In_1708,In_2728);
xor U2786 (N_2786,In_2333,In_1526);
nor U2787 (N_2787,In_1574,In_1765);
or U2788 (N_2788,In_591,In_2824);
and U2789 (N_2789,In_2915,In_3569);
or U2790 (N_2790,In_968,In_1315);
and U2791 (N_2791,In_682,In_2149);
xnor U2792 (N_2792,In_1731,In_389);
and U2793 (N_2793,In_513,In_3994);
and U2794 (N_2794,In_3909,In_939);
and U2795 (N_2795,In_2123,In_4684);
and U2796 (N_2796,In_4375,In_2744);
nor U2797 (N_2797,In_3800,In_2577);
nor U2798 (N_2798,In_4567,In_3909);
or U2799 (N_2799,In_4510,In_2622);
nand U2800 (N_2800,In_906,In_513);
and U2801 (N_2801,In_4113,In_406);
and U2802 (N_2802,In_1530,In_637);
nand U2803 (N_2803,In_2973,In_3378);
or U2804 (N_2804,In_743,In_4196);
nor U2805 (N_2805,In_3563,In_2804);
or U2806 (N_2806,In_3778,In_3047);
and U2807 (N_2807,In_1869,In_4743);
or U2808 (N_2808,In_4275,In_1972);
and U2809 (N_2809,In_114,In_985);
or U2810 (N_2810,In_3357,In_1449);
nand U2811 (N_2811,In_1776,In_525);
xnor U2812 (N_2812,In_731,In_1041);
and U2813 (N_2813,In_3023,In_3912);
nand U2814 (N_2814,In_1540,In_200);
nor U2815 (N_2815,In_3379,In_4323);
or U2816 (N_2816,In_752,In_2798);
xnor U2817 (N_2817,In_1890,In_2705);
and U2818 (N_2818,In_796,In_2569);
nor U2819 (N_2819,In_4741,In_1990);
and U2820 (N_2820,In_2788,In_700);
and U2821 (N_2821,In_2708,In_2905);
nand U2822 (N_2822,In_2907,In_4163);
nand U2823 (N_2823,In_4501,In_2482);
and U2824 (N_2824,In_4193,In_3289);
xor U2825 (N_2825,In_648,In_4243);
nand U2826 (N_2826,In_614,In_2662);
xor U2827 (N_2827,In_655,In_4208);
nand U2828 (N_2828,In_2879,In_2863);
nor U2829 (N_2829,In_1674,In_1838);
nand U2830 (N_2830,In_2619,In_4673);
nor U2831 (N_2831,In_2595,In_1453);
or U2832 (N_2832,In_4361,In_3092);
and U2833 (N_2833,In_2679,In_137);
xnor U2834 (N_2834,In_734,In_2125);
and U2835 (N_2835,In_2870,In_2454);
and U2836 (N_2836,In_1186,In_3177);
nand U2837 (N_2837,In_2536,In_1013);
xor U2838 (N_2838,In_4651,In_3119);
nor U2839 (N_2839,In_2646,In_3331);
nand U2840 (N_2840,In_83,In_3261);
or U2841 (N_2841,In_2680,In_2983);
and U2842 (N_2842,In_2840,In_4124);
nor U2843 (N_2843,In_1764,In_900);
or U2844 (N_2844,In_4923,In_374);
and U2845 (N_2845,In_941,In_1652);
xor U2846 (N_2846,In_2258,In_2566);
or U2847 (N_2847,In_2020,In_3800);
nor U2848 (N_2848,In_2888,In_3893);
and U2849 (N_2849,In_1779,In_4637);
nor U2850 (N_2850,In_2030,In_2896);
nand U2851 (N_2851,In_827,In_544);
and U2852 (N_2852,In_4463,In_1721);
and U2853 (N_2853,In_355,In_878);
nand U2854 (N_2854,In_3830,In_3685);
nand U2855 (N_2855,In_1938,In_1591);
nand U2856 (N_2856,In_3083,In_54);
nand U2857 (N_2857,In_319,In_269);
or U2858 (N_2858,In_612,In_4509);
xor U2859 (N_2859,In_2106,In_1719);
nand U2860 (N_2860,In_3471,In_4842);
or U2861 (N_2861,In_2629,In_4884);
nand U2862 (N_2862,In_1747,In_1083);
and U2863 (N_2863,In_3311,In_2689);
xor U2864 (N_2864,In_3690,In_3432);
xnor U2865 (N_2865,In_1860,In_1681);
nand U2866 (N_2866,In_590,In_972);
or U2867 (N_2867,In_3695,In_1661);
nand U2868 (N_2868,In_3322,In_3119);
nor U2869 (N_2869,In_3012,In_2346);
or U2870 (N_2870,In_2332,In_4994);
nand U2871 (N_2871,In_3526,In_2971);
and U2872 (N_2872,In_311,In_2205);
and U2873 (N_2873,In_1579,In_2809);
nand U2874 (N_2874,In_2653,In_1537);
and U2875 (N_2875,In_1512,In_3802);
nand U2876 (N_2876,In_68,In_4738);
nand U2877 (N_2877,In_4069,In_1278);
nor U2878 (N_2878,In_782,In_3782);
and U2879 (N_2879,In_783,In_2481);
and U2880 (N_2880,In_2883,In_4861);
nor U2881 (N_2881,In_2438,In_2209);
nor U2882 (N_2882,In_3399,In_1896);
nor U2883 (N_2883,In_4772,In_1954);
nor U2884 (N_2884,In_733,In_1868);
or U2885 (N_2885,In_2189,In_2007);
and U2886 (N_2886,In_721,In_2975);
nor U2887 (N_2887,In_963,In_3648);
nand U2888 (N_2888,In_2442,In_2732);
or U2889 (N_2889,In_1577,In_3697);
nor U2890 (N_2890,In_2868,In_2657);
and U2891 (N_2891,In_64,In_1895);
xnor U2892 (N_2892,In_41,In_1629);
nand U2893 (N_2893,In_4426,In_1273);
nor U2894 (N_2894,In_876,In_306);
nand U2895 (N_2895,In_2054,In_272);
nor U2896 (N_2896,In_1576,In_3816);
nand U2897 (N_2897,In_3954,In_2388);
or U2898 (N_2898,In_598,In_3008);
nor U2899 (N_2899,In_4838,In_4152);
or U2900 (N_2900,In_1596,In_1078);
nor U2901 (N_2901,In_1126,In_1130);
nor U2902 (N_2902,In_3274,In_3033);
nor U2903 (N_2903,In_4743,In_2373);
xnor U2904 (N_2904,In_3681,In_1760);
or U2905 (N_2905,In_4030,In_2217);
or U2906 (N_2906,In_3499,In_2454);
nand U2907 (N_2907,In_1507,In_1133);
and U2908 (N_2908,In_4558,In_2323);
and U2909 (N_2909,In_1175,In_488);
or U2910 (N_2910,In_2607,In_4442);
and U2911 (N_2911,In_2138,In_505);
nor U2912 (N_2912,In_1049,In_2776);
and U2913 (N_2913,In_2415,In_2307);
xnor U2914 (N_2914,In_3192,In_1138);
xor U2915 (N_2915,In_759,In_323);
or U2916 (N_2916,In_2742,In_1299);
or U2917 (N_2917,In_987,In_2247);
and U2918 (N_2918,In_1368,In_820);
and U2919 (N_2919,In_1893,In_1925);
and U2920 (N_2920,In_2195,In_3248);
and U2921 (N_2921,In_158,In_4025);
or U2922 (N_2922,In_1376,In_3849);
xnor U2923 (N_2923,In_1550,In_3129);
nand U2924 (N_2924,In_2369,In_4088);
and U2925 (N_2925,In_54,In_1479);
nor U2926 (N_2926,In_4517,In_4013);
nor U2927 (N_2927,In_3719,In_3038);
xor U2928 (N_2928,In_2140,In_3304);
xor U2929 (N_2929,In_464,In_2327);
nor U2930 (N_2930,In_1222,In_4415);
nand U2931 (N_2931,In_2227,In_1714);
or U2932 (N_2932,In_1837,In_1176);
nor U2933 (N_2933,In_2574,In_2014);
nor U2934 (N_2934,In_552,In_3702);
and U2935 (N_2935,In_670,In_17);
and U2936 (N_2936,In_1819,In_4689);
nor U2937 (N_2937,In_2142,In_3119);
nor U2938 (N_2938,In_1183,In_4610);
or U2939 (N_2939,In_769,In_786);
and U2940 (N_2940,In_3824,In_4933);
and U2941 (N_2941,In_1461,In_576);
or U2942 (N_2942,In_760,In_2454);
and U2943 (N_2943,In_1520,In_2742);
or U2944 (N_2944,In_1548,In_172);
xnor U2945 (N_2945,In_4653,In_2767);
nor U2946 (N_2946,In_3144,In_2286);
and U2947 (N_2947,In_2432,In_2712);
nor U2948 (N_2948,In_102,In_606);
and U2949 (N_2949,In_2593,In_80);
nand U2950 (N_2950,In_1472,In_4585);
nor U2951 (N_2951,In_3869,In_1595);
nand U2952 (N_2952,In_186,In_2422);
or U2953 (N_2953,In_912,In_4912);
and U2954 (N_2954,In_3887,In_3479);
and U2955 (N_2955,In_4995,In_3663);
and U2956 (N_2956,In_3696,In_1787);
or U2957 (N_2957,In_3458,In_1980);
or U2958 (N_2958,In_4876,In_4864);
and U2959 (N_2959,In_993,In_4519);
or U2960 (N_2960,In_1759,In_1581);
nand U2961 (N_2961,In_2769,In_345);
and U2962 (N_2962,In_1342,In_646);
nor U2963 (N_2963,In_4433,In_3619);
nor U2964 (N_2964,In_3395,In_4146);
and U2965 (N_2965,In_156,In_2902);
xor U2966 (N_2966,In_446,In_1902);
nand U2967 (N_2967,In_1077,In_1514);
and U2968 (N_2968,In_2835,In_1478);
or U2969 (N_2969,In_2366,In_4789);
and U2970 (N_2970,In_2562,In_1951);
or U2971 (N_2971,In_1378,In_4309);
nand U2972 (N_2972,In_252,In_2017);
and U2973 (N_2973,In_3723,In_3961);
and U2974 (N_2974,In_4988,In_4182);
and U2975 (N_2975,In_3352,In_4680);
or U2976 (N_2976,In_4331,In_2346);
nand U2977 (N_2977,In_1826,In_4847);
and U2978 (N_2978,In_497,In_3160);
and U2979 (N_2979,In_2988,In_3690);
and U2980 (N_2980,In_3500,In_4329);
nand U2981 (N_2981,In_4357,In_148);
and U2982 (N_2982,In_4803,In_1513);
and U2983 (N_2983,In_4616,In_4848);
or U2984 (N_2984,In_3439,In_4499);
nor U2985 (N_2985,In_3515,In_4697);
xor U2986 (N_2986,In_1532,In_261);
nand U2987 (N_2987,In_2896,In_1199);
or U2988 (N_2988,In_619,In_1589);
nor U2989 (N_2989,In_535,In_3002);
and U2990 (N_2990,In_2490,In_4916);
or U2991 (N_2991,In_4835,In_4361);
nand U2992 (N_2992,In_2350,In_319);
xnor U2993 (N_2993,In_2272,In_4502);
or U2994 (N_2994,In_2995,In_568);
xor U2995 (N_2995,In_2821,In_4658);
nand U2996 (N_2996,In_2389,In_3961);
and U2997 (N_2997,In_205,In_2055);
nand U2998 (N_2998,In_3093,In_1854);
and U2999 (N_2999,In_3561,In_2842);
or U3000 (N_3000,In_3242,In_1914);
xnor U3001 (N_3001,In_4755,In_1458);
nand U3002 (N_3002,In_2340,In_694);
nand U3003 (N_3003,In_3009,In_3864);
nand U3004 (N_3004,In_2201,In_867);
xor U3005 (N_3005,In_1777,In_2531);
or U3006 (N_3006,In_2027,In_1524);
nor U3007 (N_3007,In_1733,In_4429);
nor U3008 (N_3008,In_4292,In_198);
and U3009 (N_3009,In_1550,In_633);
xor U3010 (N_3010,In_4584,In_1289);
or U3011 (N_3011,In_2306,In_2234);
nor U3012 (N_3012,In_1167,In_4151);
nor U3013 (N_3013,In_3076,In_2329);
or U3014 (N_3014,In_1232,In_4166);
or U3015 (N_3015,In_2217,In_2924);
and U3016 (N_3016,In_3455,In_2141);
or U3017 (N_3017,In_1401,In_2823);
and U3018 (N_3018,In_3342,In_3448);
xor U3019 (N_3019,In_792,In_4246);
nand U3020 (N_3020,In_1266,In_1495);
xor U3021 (N_3021,In_2379,In_2491);
and U3022 (N_3022,In_3568,In_4108);
nor U3023 (N_3023,In_1854,In_129);
and U3024 (N_3024,In_4132,In_3673);
nand U3025 (N_3025,In_1738,In_215);
xnor U3026 (N_3026,In_2534,In_1084);
nand U3027 (N_3027,In_112,In_2705);
nor U3028 (N_3028,In_829,In_120);
nand U3029 (N_3029,In_2914,In_2516);
and U3030 (N_3030,In_2389,In_2024);
or U3031 (N_3031,In_290,In_2769);
or U3032 (N_3032,In_2920,In_4144);
nand U3033 (N_3033,In_2351,In_806);
nand U3034 (N_3034,In_3973,In_3707);
and U3035 (N_3035,In_1275,In_3839);
nor U3036 (N_3036,In_1640,In_59);
and U3037 (N_3037,In_2823,In_657);
nor U3038 (N_3038,In_3927,In_733);
and U3039 (N_3039,In_4118,In_3087);
and U3040 (N_3040,In_1641,In_311);
nand U3041 (N_3041,In_230,In_1250);
nand U3042 (N_3042,In_2237,In_3599);
nor U3043 (N_3043,In_2414,In_3489);
or U3044 (N_3044,In_4450,In_1);
nand U3045 (N_3045,In_4756,In_2249);
nand U3046 (N_3046,In_4003,In_4105);
nand U3047 (N_3047,In_4299,In_3429);
nor U3048 (N_3048,In_897,In_4275);
nor U3049 (N_3049,In_1487,In_223);
nor U3050 (N_3050,In_2130,In_1097);
nor U3051 (N_3051,In_1512,In_608);
nor U3052 (N_3052,In_260,In_4601);
nand U3053 (N_3053,In_1271,In_4217);
and U3054 (N_3054,In_4876,In_3248);
or U3055 (N_3055,In_2187,In_1108);
nand U3056 (N_3056,In_3416,In_2197);
or U3057 (N_3057,In_4843,In_2011);
xor U3058 (N_3058,In_1429,In_3675);
nor U3059 (N_3059,In_4195,In_4682);
or U3060 (N_3060,In_2035,In_2979);
xor U3061 (N_3061,In_2874,In_4486);
nor U3062 (N_3062,In_3288,In_2288);
nor U3063 (N_3063,In_3666,In_3735);
or U3064 (N_3064,In_1734,In_4899);
and U3065 (N_3065,In_3952,In_4401);
nand U3066 (N_3066,In_1592,In_4839);
nand U3067 (N_3067,In_4673,In_1845);
or U3068 (N_3068,In_2386,In_2489);
nor U3069 (N_3069,In_2085,In_2516);
or U3070 (N_3070,In_2560,In_624);
nor U3071 (N_3071,In_4099,In_1055);
nand U3072 (N_3072,In_1088,In_4945);
and U3073 (N_3073,In_4552,In_839);
xor U3074 (N_3074,In_1860,In_1524);
xor U3075 (N_3075,In_533,In_2485);
and U3076 (N_3076,In_2173,In_1716);
nor U3077 (N_3077,In_1877,In_2844);
nor U3078 (N_3078,In_3986,In_2556);
nor U3079 (N_3079,In_2398,In_4847);
nand U3080 (N_3080,In_2424,In_2246);
or U3081 (N_3081,In_4417,In_68);
or U3082 (N_3082,In_4234,In_2274);
or U3083 (N_3083,In_3781,In_1042);
nand U3084 (N_3084,In_3384,In_350);
nor U3085 (N_3085,In_1949,In_3607);
nor U3086 (N_3086,In_45,In_2891);
nand U3087 (N_3087,In_2497,In_2583);
or U3088 (N_3088,In_2026,In_3630);
nand U3089 (N_3089,In_2816,In_4999);
xor U3090 (N_3090,In_2968,In_1854);
and U3091 (N_3091,In_849,In_731);
nand U3092 (N_3092,In_4164,In_2361);
or U3093 (N_3093,In_4401,In_1743);
nand U3094 (N_3094,In_971,In_1003);
and U3095 (N_3095,In_3249,In_2327);
and U3096 (N_3096,In_1068,In_1575);
nand U3097 (N_3097,In_755,In_553);
nor U3098 (N_3098,In_618,In_1766);
and U3099 (N_3099,In_4136,In_2962);
or U3100 (N_3100,In_4505,In_1375);
and U3101 (N_3101,In_3877,In_4363);
nor U3102 (N_3102,In_4487,In_3157);
nand U3103 (N_3103,In_1930,In_4705);
or U3104 (N_3104,In_4320,In_131);
nor U3105 (N_3105,In_4987,In_2435);
nor U3106 (N_3106,In_359,In_3497);
nor U3107 (N_3107,In_781,In_1937);
nand U3108 (N_3108,In_4236,In_1056);
nand U3109 (N_3109,In_3369,In_710);
or U3110 (N_3110,In_1131,In_2598);
and U3111 (N_3111,In_1156,In_2020);
xor U3112 (N_3112,In_27,In_4844);
xnor U3113 (N_3113,In_3813,In_4484);
nor U3114 (N_3114,In_3704,In_4993);
nor U3115 (N_3115,In_4117,In_2622);
nand U3116 (N_3116,In_4045,In_2354);
or U3117 (N_3117,In_859,In_153);
or U3118 (N_3118,In_217,In_107);
or U3119 (N_3119,In_445,In_4903);
and U3120 (N_3120,In_701,In_4759);
or U3121 (N_3121,In_596,In_744);
or U3122 (N_3122,In_203,In_2905);
nand U3123 (N_3123,In_4386,In_3566);
nand U3124 (N_3124,In_889,In_2795);
xor U3125 (N_3125,In_4594,In_3936);
and U3126 (N_3126,In_2547,In_4466);
nand U3127 (N_3127,In_3446,In_1681);
xnor U3128 (N_3128,In_3936,In_2211);
nor U3129 (N_3129,In_1700,In_3647);
and U3130 (N_3130,In_373,In_2904);
nor U3131 (N_3131,In_852,In_1194);
and U3132 (N_3132,In_1139,In_4989);
and U3133 (N_3133,In_1387,In_4810);
or U3134 (N_3134,In_332,In_1945);
and U3135 (N_3135,In_4607,In_2493);
xor U3136 (N_3136,In_3929,In_2189);
and U3137 (N_3137,In_1393,In_2723);
nand U3138 (N_3138,In_1018,In_917);
and U3139 (N_3139,In_21,In_2141);
nand U3140 (N_3140,In_602,In_3710);
nor U3141 (N_3141,In_1831,In_2637);
xor U3142 (N_3142,In_3087,In_2909);
or U3143 (N_3143,In_1775,In_4282);
nor U3144 (N_3144,In_1622,In_3199);
xnor U3145 (N_3145,In_3377,In_3519);
nand U3146 (N_3146,In_2999,In_2958);
nand U3147 (N_3147,In_3823,In_2354);
or U3148 (N_3148,In_4783,In_4789);
xnor U3149 (N_3149,In_803,In_2874);
xnor U3150 (N_3150,In_719,In_2964);
and U3151 (N_3151,In_1639,In_1638);
nor U3152 (N_3152,In_2018,In_3438);
nand U3153 (N_3153,In_1752,In_597);
and U3154 (N_3154,In_73,In_3146);
nor U3155 (N_3155,In_4181,In_2615);
or U3156 (N_3156,In_1870,In_684);
nand U3157 (N_3157,In_3195,In_2462);
nand U3158 (N_3158,In_4136,In_4792);
or U3159 (N_3159,In_4574,In_561);
and U3160 (N_3160,In_2223,In_2928);
nand U3161 (N_3161,In_2363,In_3745);
xor U3162 (N_3162,In_2587,In_2072);
nor U3163 (N_3163,In_2435,In_171);
and U3164 (N_3164,In_2187,In_1037);
or U3165 (N_3165,In_445,In_509);
and U3166 (N_3166,In_1376,In_3514);
xor U3167 (N_3167,In_3193,In_926);
xnor U3168 (N_3168,In_3738,In_3132);
nor U3169 (N_3169,In_4757,In_710);
and U3170 (N_3170,In_3249,In_2553);
and U3171 (N_3171,In_3738,In_2521);
or U3172 (N_3172,In_1356,In_4428);
and U3173 (N_3173,In_4315,In_3714);
nand U3174 (N_3174,In_2609,In_3622);
and U3175 (N_3175,In_273,In_3715);
and U3176 (N_3176,In_2395,In_2979);
xor U3177 (N_3177,In_99,In_4544);
nand U3178 (N_3178,In_4290,In_1266);
and U3179 (N_3179,In_3298,In_1598);
or U3180 (N_3180,In_83,In_2492);
nand U3181 (N_3181,In_4841,In_2510);
xor U3182 (N_3182,In_4305,In_1894);
and U3183 (N_3183,In_3362,In_2887);
nor U3184 (N_3184,In_3490,In_2385);
and U3185 (N_3185,In_740,In_3063);
nor U3186 (N_3186,In_4196,In_4896);
xnor U3187 (N_3187,In_3889,In_2715);
xor U3188 (N_3188,In_1533,In_2442);
and U3189 (N_3189,In_4841,In_2903);
nand U3190 (N_3190,In_342,In_1179);
or U3191 (N_3191,In_367,In_2944);
nand U3192 (N_3192,In_4624,In_408);
or U3193 (N_3193,In_1878,In_282);
and U3194 (N_3194,In_2008,In_1428);
nor U3195 (N_3195,In_1467,In_1453);
xnor U3196 (N_3196,In_869,In_4946);
or U3197 (N_3197,In_414,In_3218);
or U3198 (N_3198,In_4,In_1845);
nor U3199 (N_3199,In_4627,In_1652);
or U3200 (N_3200,In_1602,In_1521);
xnor U3201 (N_3201,In_2318,In_3963);
nand U3202 (N_3202,In_4489,In_4528);
and U3203 (N_3203,In_1036,In_2969);
or U3204 (N_3204,In_3700,In_3405);
nor U3205 (N_3205,In_4396,In_3298);
and U3206 (N_3206,In_4703,In_1963);
nor U3207 (N_3207,In_1091,In_4125);
nand U3208 (N_3208,In_2785,In_325);
and U3209 (N_3209,In_3640,In_1851);
nor U3210 (N_3210,In_4305,In_3578);
or U3211 (N_3211,In_2172,In_588);
and U3212 (N_3212,In_2585,In_2383);
nor U3213 (N_3213,In_2117,In_1015);
nor U3214 (N_3214,In_4478,In_525);
nor U3215 (N_3215,In_4211,In_2968);
and U3216 (N_3216,In_2734,In_828);
nor U3217 (N_3217,In_2271,In_4983);
and U3218 (N_3218,In_4047,In_4675);
and U3219 (N_3219,In_87,In_1118);
and U3220 (N_3220,In_1596,In_4721);
and U3221 (N_3221,In_323,In_3662);
and U3222 (N_3222,In_998,In_2731);
and U3223 (N_3223,In_3588,In_2843);
or U3224 (N_3224,In_4882,In_3488);
and U3225 (N_3225,In_2464,In_4221);
and U3226 (N_3226,In_3164,In_3747);
and U3227 (N_3227,In_1605,In_2004);
nand U3228 (N_3228,In_4578,In_2162);
nand U3229 (N_3229,In_285,In_2036);
nor U3230 (N_3230,In_1255,In_3315);
xnor U3231 (N_3231,In_1422,In_2908);
nand U3232 (N_3232,In_1050,In_664);
xnor U3233 (N_3233,In_3380,In_1854);
or U3234 (N_3234,In_1558,In_2383);
and U3235 (N_3235,In_3436,In_3750);
nor U3236 (N_3236,In_4429,In_3350);
nand U3237 (N_3237,In_703,In_4987);
nand U3238 (N_3238,In_2724,In_1896);
and U3239 (N_3239,In_1020,In_564);
nand U3240 (N_3240,In_4624,In_430);
and U3241 (N_3241,In_3685,In_522);
xnor U3242 (N_3242,In_4102,In_539);
or U3243 (N_3243,In_620,In_2483);
nor U3244 (N_3244,In_2118,In_2685);
nor U3245 (N_3245,In_396,In_4003);
nand U3246 (N_3246,In_3923,In_395);
nand U3247 (N_3247,In_3371,In_4707);
nor U3248 (N_3248,In_1692,In_2320);
nand U3249 (N_3249,In_1056,In_237);
and U3250 (N_3250,In_1757,In_4933);
or U3251 (N_3251,In_4343,In_617);
nand U3252 (N_3252,In_4755,In_2328);
and U3253 (N_3253,In_4886,In_4368);
xnor U3254 (N_3254,In_1364,In_3273);
nor U3255 (N_3255,In_1951,In_1590);
or U3256 (N_3256,In_3229,In_4958);
and U3257 (N_3257,In_2785,In_4302);
nor U3258 (N_3258,In_3054,In_1597);
nor U3259 (N_3259,In_1022,In_4836);
nand U3260 (N_3260,In_727,In_2510);
and U3261 (N_3261,In_4167,In_2421);
and U3262 (N_3262,In_4588,In_2223);
or U3263 (N_3263,In_4054,In_245);
or U3264 (N_3264,In_2302,In_4734);
nand U3265 (N_3265,In_4449,In_377);
and U3266 (N_3266,In_530,In_1507);
nand U3267 (N_3267,In_2183,In_2478);
nor U3268 (N_3268,In_833,In_144);
nand U3269 (N_3269,In_4637,In_3791);
xnor U3270 (N_3270,In_1472,In_3076);
nor U3271 (N_3271,In_2510,In_359);
nand U3272 (N_3272,In_4000,In_1980);
and U3273 (N_3273,In_3749,In_128);
nand U3274 (N_3274,In_4493,In_1486);
nand U3275 (N_3275,In_3574,In_499);
xnor U3276 (N_3276,In_170,In_922);
or U3277 (N_3277,In_3677,In_4703);
nand U3278 (N_3278,In_890,In_879);
nor U3279 (N_3279,In_3595,In_1773);
and U3280 (N_3280,In_2434,In_3052);
nor U3281 (N_3281,In_522,In_2958);
and U3282 (N_3282,In_3338,In_4069);
or U3283 (N_3283,In_2819,In_3169);
nand U3284 (N_3284,In_346,In_546);
or U3285 (N_3285,In_2957,In_1943);
xnor U3286 (N_3286,In_600,In_3709);
nand U3287 (N_3287,In_356,In_1811);
nand U3288 (N_3288,In_2550,In_857);
or U3289 (N_3289,In_4631,In_3324);
nor U3290 (N_3290,In_2296,In_2573);
xnor U3291 (N_3291,In_723,In_1849);
xor U3292 (N_3292,In_579,In_4749);
nor U3293 (N_3293,In_3898,In_4120);
and U3294 (N_3294,In_1302,In_3297);
nor U3295 (N_3295,In_11,In_1852);
xnor U3296 (N_3296,In_85,In_455);
nor U3297 (N_3297,In_1446,In_656);
or U3298 (N_3298,In_1607,In_2586);
nor U3299 (N_3299,In_4607,In_162);
or U3300 (N_3300,In_4742,In_2731);
nor U3301 (N_3301,In_2929,In_356);
nor U3302 (N_3302,In_261,In_4928);
nand U3303 (N_3303,In_1427,In_3461);
and U3304 (N_3304,In_463,In_1493);
nand U3305 (N_3305,In_198,In_1339);
nand U3306 (N_3306,In_74,In_1412);
and U3307 (N_3307,In_4619,In_4714);
nor U3308 (N_3308,In_4253,In_2661);
nor U3309 (N_3309,In_4630,In_4532);
nor U3310 (N_3310,In_4346,In_1198);
nor U3311 (N_3311,In_1921,In_2960);
or U3312 (N_3312,In_2043,In_2266);
nand U3313 (N_3313,In_1345,In_4602);
nand U3314 (N_3314,In_1825,In_2340);
or U3315 (N_3315,In_1933,In_3892);
or U3316 (N_3316,In_953,In_242);
or U3317 (N_3317,In_1627,In_2185);
nand U3318 (N_3318,In_3630,In_4174);
and U3319 (N_3319,In_4152,In_4143);
nor U3320 (N_3320,In_3191,In_2892);
nor U3321 (N_3321,In_2350,In_729);
and U3322 (N_3322,In_4996,In_747);
or U3323 (N_3323,In_2116,In_3175);
or U3324 (N_3324,In_1361,In_2932);
nor U3325 (N_3325,In_2027,In_3711);
or U3326 (N_3326,In_59,In_90);
nor U3327 (N_3327,In_897,In_1574);
or U3328 (N_3328,In_2215,In_4094);
nand U3329 (N_3329,In_310,In_3333);
nor U3330 (N_3330,In_2111,In_4258);
nor U3331 (N_3331,In_1111,In_735);
and U3332 (N_3332,In_4217,In_4141);
xnor U3333 (N_3333,In_4019,In_2239);
and U3334 (N_3334,In_827,In_2531);
nand U3335 (N_3335,In_70,In_1309);
and U3336 (N_3336,In_4617,In_2686);
nor U3337 (N_3337,In_1598,In_4724);
nand U3338 (N_3338,In_2619,In_3388);
nor U3339 (N_3339,In_4039,In_1025);
and U3340 (N_3340,In_2732,In_82);
and U3341 (N_3341,In_4622,In_2772);
nand U3342 (N_3342,In_1271,In_1664);
nor U3343 (N_3343,In_1480,In_4426);
and U3344 (N_3344,In_3394,In_3849);
or U3345 (N_3345,In_800,In_4997);
and U3346 (N_3346,In_3918,In_3194);
xor U3347 (N_3347,In_2360,In_3977);
nor U3348 (N_3348,In_2083,In_1691);
nor U3349 (N_3349,In_2887,In_3125);
and U3350 (N_3350,In_1442,In_3047);
nand U3351 (N_3351,In_3605,In_4619);
and U3352 (N_3352,In_2749,In_4019);
or U3353 (N_3353,In_3055,In_1156);
or U3354 (N_3354,In_4300,In_729);
nand U3355 (N_3355,In_3035,In_3490);
or U3356 (N_3356,In_2135,In_157);
and U3357 (N_3357,In_2969,In_4197);
and U3358 (N_3358,In_1865,In_3708);
and U3359 (N_3359,In_2480,In_4977);
nor U3360 (N_3360,In_528,In_4287);
and U3361 (N_3361,In_1786,In_1536);
nor U3362 (N_3362,In_3248,In_1676);
or U3363 (N_3363,In_2623,In_1527);
nand U3364 (N_3364,In_4144,In_2940);
xor U3365 (N_3365,In_3368,In_1425);
nor U3366 (N_3366,In_4768,In_4686);
nand U3367 (N_3367,In_3429,In_1641);
xor U3368 (N_3368,In_2532,In_1617);
or U3369 (N_3369,In_1466,In_3911);
nor U3370 (N_3370,In_1706,In_583);
or U3371 (N_3371,In_1151,In_4026);
nor U3372 (N_3372,In_2763,In_4890);
nor U3373 (N_3373,In_2242,In_2935);
and U3374 (N_3374,In_2237,In_2160);
or U3375 (N_3375,In_40,In_2133);
and U3376 (N_3376,In_4017,In_1619);
nand U3377 (N_3377,In_4901,In_623);
nand U3378 (N_3378,In_1553,In_3193);
nor U3379 (N_3379,In_3866,In_2137);
nor U3380 (N_3380,In_570,In_3438);
nor U3381 (N_3381,In_4483,In_2211);
and U3382 (N_3382,In_512,In_1984);
and U3383 (N_3383,In_4612,In_645);
and U3384 (N_3384,In_1512,In_1225);
nand U3385 (N_3385,In_2628,In_4378);
nor U3386 (N_3386,In_2057,In_672);
nor U3387 (N_3387,In_4500,In_3745);
and U3388 (N_3388,In_3272,In_4939);
or U3389 (N_3389,In_2663,In_4591);
nand U3390 (N_3390,In_1403,In_4693);
and U3391 (N_3391,In_2087,In_4203);
nand U3392 (N_3392,In_140,In_951);
and U3393 (N_3393,In_4117,In_1665);
nor U3394 (N_3394,In_3550,In_3259);
and U3395 (N_3395,In_3147,In_4815);
or U3396 (N_3396,In_308,In_2067);
nand U3397 (N_3397,In_303,In_4573);
nor U3398 (N_3398,In_2174,In_184);
or U3399 (N_3399,In_556,In_4917);
or U3400 (N_3400,In_575,In_2786);
nand U3401 (N_3401,In_4963,In_3334);
nand U3402 (N_3402,In_4791,In_1064);
and U3403 (N_3403,In_323,In_3587);
and U3404 (N_3404,In_2588,In_862);
or U3405 (N_3405,In_3597,In_4075);
nand U3406 (N_3406,In_2706,In_858);
xor U3407 (N_3407,In_1754,In_3732);
or U3408 (N_3408,In_4532,In_2177);
nor U3409 (N_3409,In_1709,In_608);
nor U3410 (N_3410,In_1316,In_1432);
nor U3411 (N_3411,In_4496,In_2664);
and U3412 (N_3412,In_4853,In_2609);
nand U3413 (N_3413,In_2135,In_2025);
nor U3414 (N_3414,In_1204,In_2687);
or U3415 (N_3415,In_1161,In_1277);
or U3416 (N_3416,In_1880,In_2299);
and U3417 (N_3417,In_1954,In_1788);
nor U3418 (N_3418,In_1069,In_4313);
nand U3419 (N_3419,In_3053,In_2052);
nor U3420 (N_3420,In_289,In_2302);
and U3421 (N_3421,In_395,In_4490);
and U3422 (N_3422,In_1234,In_3713);
or U3423 (N_3423,In_2556,In_3916);
and U3424 (N_3424,In_3480,In_4498);
nor U3425 (N_3425,In_4231,In_3992);
nand U3426 (N_3426,In_973,In_2492);
nand U3427 (N_3427,In_2967,In_1534);
or U3428 (N_3428,In_1850,In_492);
nand U3429 (N_3429,In_2140,In_4247);
and U3430 (N_3430,In_4611,In_1775);
and U3431 (N_3431,In_1450,In_578);
or U3432 (N_3432,In_1508,In_1128);
nand U3433 (N_3433,In_4338,In_563);
nand U3434 (N_3434,In_3768,In_2259);
nor U3435 (N_3435,In_4249,In_4391);
and U3436 (N_3436,In_22,In_2715);
xor U3437 (N_3437,In_2889,In_4285);
and U3438 (N_3438,In_1760,In_743);
nor U3439 (N_3439,In_4685,In_3660);
nor U3440 (N_3440,In_939,In_1450);
or U3441 (N_3441,In_1249,In_1924);
or U3442 (N_3442,In_3324,In_1341);
and U3443 (N_3443,In_398,In_2177);
nand U3444 (N_3444,In_4400,In_2845);
nand U3445 (N_3445,In_3638,In_3109);
nand U3446 (N_3446,In_2330,In_3568);
nand U3447 (N_3447,In_4543,In_2268);
nor U3448 (N_3448,In_3746,In_1812);
or U3449 (N_3449,In_4769,In_3290);
xor U3450 (N_3450,In_3595,In_4745);
and U3451 (N_3451,In_3864,In_3179);
nor U3452 (N_3452,In_1345,In_4892);
nand U3453 (N_3453,In_1765,In_4351);
nand U3454 (N_3454,In_3990,In_2015);
nand U3455 (N_3455,In_1367,In_1240);
xnor U3456 (N_3456,In_4023,In_709);
and U3457 (N_3457,In_2781,In_2350);
and U3458 (N_3458,In_4530,In_4201);
nand U3459 (N_3459,In_1487,In_3559);
or U3460 (N_3460,In_1920,In_4521);
nor U3461 (N_3461,In_3200,In_3154);
and U3462 (N_3462,In_4900,In_3035);
nand U3463 (N_3463,In_3460,In_3345);
nor U3464 (N_3464,In_312,In_3019);
or U3465 (N_3465,In_1625,In_4895);
nor U3466 (N_3466,In_2005,In_2647);
or U3467 (N_3467,In_2726,In_280);
nor U3468 (N_3468,In_3092,In_1018);
or U3469 (N_3469,In_369,In_4216);
and U3470 (N_3470,In_2845,In_1595);
and U3471 (N_3471,In_600,In_2549);
xnor U3472 (N_3472,In_4307,In_4688);
and U3473 (N_3473,In_4490,In_3775);
or U3474 (N_3474,In_650,In_97);
and U3475 (N_3475,In_4486,In_1239);
xor U3476 (N_3476,In_2169,In_776);
or U3477 (N_3477,In_3885,In_2016);
and U3478 (N_3478,In_4520,In_1349);
nor U3479 (N_3479,In_634,In_1118);
nor U3480 (N_3480,In_2455,In_527);
or U3481 (N_3481,In_2064,In_569);
nand U3482 (N_3482,In_2250,In_1645);
and U3483 (N_3483,In_370,In_3745);
and U3484 (N_3484,In_4289,In_3050);
nor U3485 (N_3485,In_1270,In_1582);
or U3486 (N_3486,In_1867,In_84);
or U3487 (N_3487,In_950,In_4865);
nand U3488 (N_3488,In_801,In_2112);
nor U3489 (N_3489,In_2364,In_3649);
xnor U3490 (N_3490,In_3536,In_4836);
and U3491 (N_3491,In_847,In_1369);
nand U3492 (N_3492,In_2796,In_4825);
and U3493 (N_3493,In_1069,In_137);
or U3494 (N_3494,In_764,In_1380);
nor U3495 (N_3495,In_857,In_363);
or U3496 (N_3496,In_4276,In_4284);
or U3497 (N_3497,In_4631,In_3676);
or U3498 (N_3498,In_3785,In_1359);
and U3499 (N_3499,In_852,In_4814);
nor U3500 (N_3500,In_1428,In_915);
and U3501 (N_3501,In_3020,In_750);
nand U3502 (N_3502,In_4380,In_2367);
and U3503 (N_3503,In_1505,In_1344);
nor U3504 (N_3504,In_56,In_3150);
or U3505 (N_3505,In_3783,In_472);
or U3506 (N_3506,In_3970,In_220);
nand U3507 (N_3507,In_4803,In_1158);
nor U3508 (N_3508,In_3590,In_794);
and U3509 (N_3509,In_1083,In_307);
or U3510 (N_3510,In_2367,In_3762);
xor U3511 (N_3511,In_1303,In_1725);
nand U3512 (N_3512,In_4886,In_247);
and U3513 (N_3513,In_380,In_2931);
or U3514 (N_3514,In_3472,In_2310);
xor U3515 (N_3515,In_782,In_755);
nand U3516 (N_3516,In_2368,In_4659);
nor U3517 (N_3517,In_280,In_4191);
and U3518 (N_3518,In_4996,In_4134);
and U3519 (N_3519,In_3349,In_4559);
or U3520 (N_3520,In_2748,In_4585);
or U3521 (N_3521,In_3752,In_4997);
or U3522 (N_3522,In_4784,In_4597);
and U3523 (N_3523,In_1962,In_1242);
nand U3524 (N_3524,In_513,In_4364);
nand U3525 (N_3525,In_977,In_1600);
and U3526 (N_3526,In_4469,In_797);
nand U3527 (N_3527,In_1634,In_1251);
or U3528 (N_3528,In_3108,In_286);
nor U3529 (N_3529,In_4883,In_2552);
nand U3530 (N_3530,In_4349,In_4050);
xor U3531 (N_3531,In_1449,In_2659);
nor U3532 (N_3532,In_1767,In_551);
nand U3533 (N_3533,In_4789,In_2110);
or U3534 (N_3534,In_3159,In_2775);
nor U3535 (N_3535,In_4090,In_1803);
nor U3536 (N_3536,In_3869,In_1645);
xor U3537 (N_3537,In_2805,In_2195);
and U3538 (N_3538,In_1812,In_2470);
or U3539 (N_3539,In_3001,In_2086);
nor U3540 (N_3540,In_4588,In_1137);
nand U3541 (N_3541,In_2003,In_287);
nor U3542 (N_3542,In_869,In_1929);
and U3543 (N_3543,In_1309,In_4923);
xnor U3544 (N_3544,In_891,In_2213);
nor U3545 (N_3545,In_1191,In_3112);
nand U3546 (N_3546,In_4266,In_1103);
nand U3547 (N_3547,In_4729,In_1825);
and U3548 (N_3548,In_3245,In_2020);
nor U3549 (N_3549,In_3885,In_2144);
xnor U3550 (N_3550,In_4387,In_4185);
and U3551 (N_3551,In_831,In_1844);
and U3552 (N_3552,In_155,In_3574);
or U3553 (N_3553,In_145,In_656);
nor U3554 (N_3554,In_1631,In_4739);
nor U3555 (N_3555,In_3549,In_3151);
nor U3556 (N_3556,In_1328,In_774);
or U3557 (N_3557,In_4779,In_2271);
or U3558 (N_3558,In_1386,In_17);
and U3559 (N_3559,In_3055,In_763);
nor U3560 (N_3560,In_4313,In_454);
and U3561 (N_3561,In_4114,In_1651);
or U3562 (N_3562,In_1163,In_4119);
and U3563 (N_3563,In_4958,In_4284);
and U3564 (N_3564,In_2530,In_1236);
and U3565 (N_3565,In_1059,In_4589);
nand U3566 (N_3566,In_3978,In_1958);
xor U3567 (N_3567,In_2953,In_2670);
nand U3568 (N_3568,In_2193,In_3250);
nand U3569 (N_3569,In_1507,In_3543);
nand U3570 (N_3570,In_3564,In_3848);
and U3571 (N_3571,In_569,In_2152);
nand U3572 (N_3572,In_3342,In_1855);
nor U3573 (N_3573,In_3718,In_2264);
nand U3574 (N_3574,In_2758,In_3756);
and U3575 (N_3575,In_1997,In_1079);
and U3576 (N_3576,In_3178,In_491);
nor U3577 (N_3577,In_4382,In_216);
and U3578 (N_3578,In_1785,In_3334);
xnor U3579 (N_3579,In_1685,In_4396);
nand U3580 (N_3580,In_439,In_2882);
nand U3581 (N_3581,In_268,In_837);
or U3582 (N_3582,In_4989,In_2861);
or U3583 (N_3583,In_3491,In_2673);
or U3584 (N_3584,In_3264,In_141);
nor U3585 (N_3585,In_599,In_4823);
and U3586 (N_3586,In_46,In_4674);
nor U3587 (N_3587,In_1263,In_4264);
nand U3588 (N_3588,In_1081,In_1781);
nand U3589 (N_3589,In_4324,In_3443);
nor U3590 (N_3590,In_201,In_1448);
or U3591 (N_3591,In_3236,In_3830);
or U3592 (N_3592,In_1400,In_3805);
nor U3593 (N_3593,In_4183,In_4668);
nand U3594 (N_3594,In_1378,In_4755);
nand U3595 (N_3595,In_2593,In_1945);
or U3596 (N_3596,In_779,In_997);
or U3597 (N_3597,In_4562,In_3503);
and U3598 (N_3598,In_1797,In_2280);
and U3599 (N_3599,In_1227,In_2881);
or U3600 (N_3600,In_698,In_1429);
nor U3601 (N_3601,In_3561,In_2521);
and U3602 (N_3602,In_3110,In_1988);
or U3603 (N_3603,In_4369,In_2502);
nand U3604 (N_3604,In_1274,In_1553);
nand U3605 (N_3605,In_3115,In_574);
xnor U3606 (N_3606,In_2369,In_3758);
or U3607 (N_3607,In_2888,In_4000);
or U3608 (N_3608,In_241,In_4302);
nor U3609 (N_3609,In_2401,In_1844);
nand U3610 (N_3610,In_3488,In_4353);
nor U3611 (N_3611,In_546,In_1707);
nor U3612 (N_3612,In_2248,In_329);
and U3613 (N_3613,In_2522,In_33);
or U3614 (N_3614,In_4615,In_4479);
or U3615 (N_3615,In_1051,In_98);
xor U3616 (N_3616,In_2509,In_3097);
or U3617 (N_3617,In_4265,In_4857);
nor U3618 (N_3618,In_4763,In_2574);
nand U3619 (N_3619,In_3385,In_1555);
nor U3620 (N_3620,In_1657,In_4461);
nor U3621 (N_3621,In_1188,In_1996);
nor U3622 (N_3622,In_3638,In_4024);
nor U3623 (N_3623,In_3200,In_1421);
nor U3624 (N_3624,In_993,In_2651);
and U3625 (N_3625,In_4430,In_2719);
nor U3626 (N_3626,In_3453,In_673);
nor U3627 (N_3627,In_4749,In_808);
or U3628 (N_3628,In_4027,In_3352);
or U3629 (N_3629,In_148,In_4349);
xnor U3630 (N_3630,In_10,In_1474);
and U3631 (N_3631,In_99,In_2439);
and U3632 (N_3632,In_3416,In_659);
nand U3633 (N_3633,In_407,In_2018);
or U3634 (N_3634,In_1587,In_2001);
nand U3635 (N_3635,In_1126,In_2982);
and U3636 (N_3636,In_579,In_2202);
or U3637 (N_3637,In_2100,In_2141);
or U3638 (N_3638,In_3077,In_1735);
nand U3639 (N_3639,In_4666,In_919);
nand U3640 (N_3640,In_3058,In_3194);
and U3641 (N_3641,In_3772,In_2736);
nand U3642 (N_3642,In_2531,In_578);
nor U3643 (N_3643,In_4646,In_3865);
or U3644 (N_3644,In_4477,In_509);
xnor U3645 (N_3645,In_1185,In_3114);
xor U3646 (N_3646,In_1606,In_1908);
or U3647 (N_3647,In_311,In_3054);
and U3648 (N_3648,In_4749,In_3240);
and U3649 (N_3649,In_3975,In_1800);
nand U3650 (N_3650,In_1035,In_288);
or U3651 (N_3651,In_2568,In_4680);
nor U3652 (N_3652,In_4946,In_3481);
or U3653 (N_3653,In_4465,In_4668);
nand U3654 (N_3654,In_1524,In_4634);
nor U3655 (N_3655,In_2810,In_885);
nor U3656 (N_3656,In_2475,In_2712);
nor U3657 (N_3657,In_2751,In_3857);
nand U3658 (N_3658,In_4781,In_4558);
nand U3659 (N_3659,In_3702,In_1706);
nor U3660 (N_3660,In_1905,In_979);
nor U3661 (N_3661,In_3861,In_3068);
nand U3662 (N_3662,In_4743,In_380);
nand U3663 (N_3663,In_2117,In_2115);
xor U3664 (N_3664,In_4167,In_3011);
nor U3665 (N_3665,In_156,In_4219);
and U3666 (N_3666,In_4678,In_1893);
and U3667 (N_3667,In_2069,In_3083);
and U3668 (N_3668,In_4690,In_1955);
xnor U3669 (N_3669,In_4627,In_4652);
xor U3670 (N_3670,In_1453,In_3642);
and U3671 (N_3671,In_3483,In_3158);
nor U3672 (N_3672,In_1626,In_3862);
nor U3673 (N_3673,In_2875,In_2684);
nand U3674 (N_3674,In_4165,In_4492);
and U3675 (N_3675,In_2319,In_4818);
xor U3676 (N_3676,In_216,In_4946);
and U3677 (N_3677,In_3977,In_3605);
xor U3678 (N_3678,In_3564,In_186);
and U3679 (N_3679,In_4816,In_2876);
nand U3680 (N_3680,In_1670,In_4554);
nor U3681 (N_3681,In_2137,In_2513);
nor U3682 (N_3682,In_2329,In_3498);
xor U3683 (N_3683,In_1016,In_4357);
and U3684 (N_3684,In_2902,In_2287);
and U3685 (N_3685,In_987,In_4286);
nor U3686 (N_3686,In_66,In_4539);
and U3687 (N_3687,In_4825,In_3029);
xnor U3688 (N_3688,In_2542,In_4730);
or U3689 (N_3689,In_2353,In_522);
or U3690 (N_3690,In_3407,In_3341);
and U3691 (N_3691,In_186,In_4097);
xor U3692 (N_3692,In_2981,In_1259);
or U3693 (N_3693,In_3392,In_3805);
nand U3694 (N_3694,In_2767,In_2387);
and U3695 (N_3695,In_2863,In_686);
and U3696 (N_3696,In_3522,In_4705);
and U3697 (N_3697,In_4282,In_1295);
xnor U3698 (N_3698,In_786,In_746);
nor U3699 (N_3699,In_427,In_4036);
or U3700 (N_3700,In_1724,In_3872);
and U3701 (N_3701,In_4513,In_2109);
or U3702 (N_3702,In_3807,In_3954);
xnor U3703 (N_3703,In_1827,In_4276);
or U3704 (N_3704,In_3009,In_2759);
and U3705 (N_3705,In_1946,In_1036);
or U3706 (N_3706,In_3002,In_510);
nand U3707 (N_3707,In_4731,In_2587);
and U3708 (N_3708,In_885,In_851);
xor U3709 (N_3709,In_1027,In_3632);
nand U3710 (N_3710,In_1251,In_4851);
nor U3711 (N_3711,In_248,In_4016);
nand U3712 (N_3712,In_4133,In_3694);
or U3713 (N_3713,In_1286,In_1797);
or U3714 (N_3714,In_2878,In_4387);
nor U3715 (N_3715,In_2326,In_63);
or U3716 (N_3716,In_4040,In_919);
or U3717 (N_3717,In_2322,In_185);
or U3718 (N_3718,In_691,In_1746);
or U3719 (N_3719,In_4898,In_4329);
or U3720 (N_3720,In_365,In_337);
nor U3721 (N_3721,In_522,In_2350);
and U3722 (N_3722,In_1686,In_2393);
or U3723 (N_3723,In_3572,In_2626);
or U3724 (N_3724,In_355,In_1238);
and U3725 (N_3725,In_2187,In_3941);
nor U3726 (N_3726,In_4655,In_1363);
nand U3727 (N_3727,In_2921,In_3999);
xnor U3728 (N_3728,In_2886,In_4446);
and U3729 (N_3729,In_1479,In_793);
nor U3730 (N_3730,In_1338,In_605);
and U3731 (N_3731,In_626,In_1618);
or U3732 (N_3732,In_2640,In_3085);
or U3733 (N_3733,In_398,In_3695);
nand U3734 (N_3734,In_1601,In_4650);
xor U3735 (N_3735,In_143,In_679);
or U3736 (N_3736,In_3,In_1876);
and U3737 (N_3737,In_3704,In_2806);
nand U3738 (N_3738,In_459,In_4460);
or U3739 (N_3739,In_720,In_3210);
or U3740 (N_3740,In_890,In_3505);
and U3741 (N_3741,In_2201,In_903);
and U3742 (N_3742,In_4154,In_2218);
nand U3743 (N_3743,In_4535,In_1874);
and U3744 (N_3744,In_193,In_1521);
and U3745 (N_3745,In_25,In_4816);
nand U3746 (N_3746,In_519,In_4523);
and U3747 (N_3747,In_4665,In_1491);
or U3748 (N_3748,In_431,In_791);
nor U3749 (N_3749,In_1842,In_1898);
nand U3750 (N_3750,In_4600,In_3370);
nand U3751 (N_3751,In_110,In_4091);
nand U3752 (N_3752,In_2771,In_4975);
nor U3753 (N_3753,In_4710,In_3057);
xnor U3754 (N_3754,In_1508,In_3140);
or U3755 (N_3755,In_1373,In_2642);
or U3756 (N_3756,In_4643,In_2054);
xor U3757 (N_3757,In_4332,In_2250);
nand U3758 (N_3758,In_921,In_181);
or U3759 (N_3759,In_3515,In_3281);
or U3760 (N_3760,In_4592,In_1313);
nand U3761 (N_3761,In_3852,In_589);
nor U3762 (N_3762,In_4903,In_333);
nor U3763 (N_3763,In_4506,In_622);
or U3764 (N_3764,In_599,In_2356);
nand U3765 (N_3765,In_4813,In_3847);
xor U3766 (N_3766,In_4945,In_2035);
or U3767 (N_3767,In_4804,In_3723);
nand U3768 (N_3768,In_4815,In_1688);
nand U3769 (N_3769,In_2347,In_1877);
xor U3770 (N_3770,In_1115,In_3604);
nor U3771 (N_3771,In_4150,In_2604);
or U3772 (N_3772,In_615,In_1429);
and U3773 (N_3773,In_4562,In_315);
nand U3774 (N_3774,In_2438,In_4214);
nor U3775 (N_3775,In_2129,In_3313);
nor U3776 (N_3776,In_2434,In_2626);
xnor U3777 (N_3777,In_736,In_2119);
and U3778 (N_3778,In_1426,In_4743);
and U3779 (N_3779,In_4489,In_143);
nor U3780 (N_3780,In_457,In_2127);
and U3781 (N_3781,In_4280,In_3342);
xor U3782 (N_3782,In_4784,In_2183);
nand U3783 (N_3783,In_4291,In_644);
or U3784 (N_3784,In_421,In_3177);
and U3785 (N_3785,In_566,In_632);
or U3786 (N_3786,In_4239,In_1224);
nor U3787 (N_3787,In_4160,In_4420);
nand U3788 (N_3788,In_4602,In_2615);
and U3789 (N_3789,In_1194,In_719);
nor U3790 (N_3790,In_1088,In_3894);
and U3791 (N_3791,In_2334,In_108);
nor U3792 (N_3792,In_1226,In_3236);
xnor U3793 (N_3793,In_2505,In_331);
nor U3794 (N_3794,In_4771,In_3165);
nand U3795 (N_3795,In_1012,In_1129);
nor U3796 (N_3796,In_3767,In_2050);
nor U3797 (N_3797,In_4426,In_2624);
or U3798 (N_3798,In_945,In_4219);
nor U3799 (N_3799,In_3708,In_4258);
nor U3800 (N_3800,In_4687,In_245);
nor U3801 (N_3801,In_4592,In_2512);
or U3802 (N_3802,In_4449,In_4004);
or U3803 (N_3803,In_4104,In_1582);
nand U3804 (N_3804,In_1507,In_2975);
nand U3805 (N_3805,In_957,In_602);
nand U3806 (N_3806,In_941,In_2767);
nand U3807 (N_3807,In_1123,In_3152);
nor U3808 (N_3808,In_831,In_2503);
and U3809 (N_3809,In_232,In_1774);
nand U3810 (N_3810,In_1742,In_4521);
nor U3811 (N_3811,In_4189,In_2);
or U3812 (N_3812,In_1486,In_1988);
nor U3813 (N_3813,In_4279,In_710);
xor U3814 (N_3814,In_1555,In_4701);
and U3815 (N_3815,In_1102,In_3566);
nor U3816 (N_3816,In_4767,In_2081);
or U3817 (N_3817,In_4667,In_2622);
and U3818 (N_3818,In_4203,In_3408);
nor U3819 (N_3819,In_3237,In_1955);
or U3820 (N_3820,In_3301,In_1330);
xor U3821 (N_3821,In_3034,In_2439);
or U3822 (N_3822,In_2049,In_2625);
or U3823 (N_3823,In_2447,In_311);
nand U3824 (N_3824,In_3554,In_882);
nand U3825 (N_3825,In_4484,In_254);
xor U3826 (N_3826,In_1360,In_3855);
nand U3827 (N_3827,In_2086,In_3429);
nor U3828 (N_3828,In_3200,In_4093);
nor U3829 (N_3829,In_3227,In_3910);
nand U3830 (N_3830,In_3123,In_4804);
and U3831 (N_3831,In_1268,In_4094);
or U3832 (N_3832,In_2275,In_2590);
or U3833 (N_3833,In_564,In_3652);
or U3834 (N_3834,In_4024,In_863);
nand U3835 (N_3835,In_1261,In_633);
nand U3836 (N_3836,In_1128,In_736);
nand U3837 (N_3837,In_1627,In_4281);
and U3838 (N_3838,In_3946,In_1755);
xnor U3839 (N_3839,In_3182,In_3980);
xnor U3840 (N_3840,In_2414,In_3486);
nand U3841 (N_3841,In_3876,In_589);
nand U3842 (N_3842,In_4514,In_4490);
xnor U3843 (N_3843,In_2887,In_3392);
and U3844 (N_3844,In_1187,In_4317);
and U3845 (N_3845,In_4541,In_4301);
or U3846 (N_3846,In_2794,In_856);
nand U3847 (N_3847,In_4070,In_4917);
nand U3848 (N_3848,In_2414,In_3885);
nand U3849 (N_3849,In_4112,In_2330);
nand U3850 (N_3850,In_3054,In_3123);
or U3851 (N_3851,In_1446,In_4791);
nor U3852 (N_3852,In_1601,In_4221);
or U3853 (N_3853,In_71,In_4486);
or U3854 (N_3854,In_995,In_1373);
nand U3855 (N_3855,In_3969,In_4401);
nor U3856 (N_3856,In_4980,In_1999);
nor U3857 (N_3857,In_454,In_3935);
and U3858 (N_3858,In_2760,In_4495);
and U3859 (N_3859,In_782,In_1736);
xnor U3860 (N_3860,In_2140,In_4606);
or U3861 (N_3861,In_745,In_3102);
or U3862 (N_3862,In_1211,In_3455);
xnor U3863 (N_3863,In_2225,In_1069);
nor U3864 (N_3864,In_571,In_459);
and U3865 (N_3865,In_4183,In_4447);
nor U3866 (N_3866,In_438,In_4030);
and U3867 (N_3867,In_4197,In_2628);
or U3868 (N_3868,In_2158,In_2541);
or U3869 (N_3869,In_4311,In_4599);
nand U3870 (N_3870,In_1244,In_1933);
xor U3871 (N_3871,In_1367,In_3606);
or U3872 (N_3872,In_709,In_1419);
nand U3873 (N_3873,In_1863,In_3523);
nor U3874 (N_3874,In_2550,In_3648);
or U3875 (N_3875,In_4079,In_3566);
nor U3876 (N_3876,In_3373,In_2489);
or U3877 (N_3877,In_269,In_2585);
nor U3878 (N_3878,In_2765,In_3628);
or U3879 (N_3879,In_4292,In_4508);
or U3880 (N_3880,In_333,In_4967);
nand U3881 (N_3881,In_1067,In_1133);
nor U3882 (N_3882,In_778,In_3348);
or U3883 (N_3883,In_3312,In_1636);
nand U3884 (N_3884,In_446,In_4753);
and U3885 (N_3885,In_3937,In_1751);
xor U3886 (N_3886,In_4612,In_1834);
nand U3887 (N_3887,In_3258,In_771);
or U3888 (N_3888,In_2435,In_1737);
and U3889 (N_3889,In_3127,In_1928);
nand U3890 (N_3890,In_2911,In_3592);
nor U3891 (N_3891,In_2527,In_176);
and U3892 (N_3892,In_2225,In_3773);
and U3893 (N_3893,In_3140,In_1042);
and U3894 (N_3894,In_4145,In_4920);
xor U3895 (N_3895,In_63,In_4975);
nand U3896 (N_3896,In_539,In_4873);
xnor U3897 (N_3897,In_1280,In_682);
nand U3898 (N_3898,In_1644,In_1727);
or U3899 (N_3899,In_2504,In_2074);
or U3900 (N_3900,In_349,In_1019);
nor U3901 (N_3901,In_600,In_2155);
xnor U3902 (N_3902,In_2549,In_1072);
nand U3903 (N_3903,In_3113,In_3597);
xor U3904 (N_3904,In_945,In_3338);
and U3905 (N_3905,In_1194,In_2853);
nor U3906 (N_3906,In_4906,In_3966);
and U3907 (N_3907,In_2354,In_3124);
nand U3908 (N_3908,In_4447,In_1939);
nand U3909 (N_3909,In_2860,In_1670);
and U3910 (N_3910,In_1361,In_1630);
nor U3911 (N_3911,In_4066,In_2172);
nand U3912 (N_3912,In_4818,In_15);
nor U3913 (N_3913,In_3579,In_4340);
nor U3914 (N_3914,In_2008,In_2892);
or U3915 (N_3915,In_803,In_1781);
nor U3916 (N_3916,In_3236,In_3417);
nand U3917 (N_3917,In_981,In_2801);
or U3918 (N_3918,In_2411,In_866);
nand U3919 (N_3919,In_3818,In_4276);
nand U3920 (N_3920,In_4673,In_1301);
or U3921 (N_3921,In_4529,In_4604);
nand U3922 (N_3922,In_1517,In_77);
and U3923 (N_3923,In_1851,In_2102);
or U3924 (N_3924,In_4563,In_179);
nor U3925 (N_3925,In_1618,In_2611);
nor U3926 (N_3926,In_4546,In_3704);
and U3927 (N_3927,In_299,In_4588);
and U3928 (N_3928,In_4224,In_3695);
xnor U3929 (N_3929,In_3060,In_4729);
nand U3930 (N_3930,In_2420,In_660);
and U3931 (N_3931,In_2760,In_2560);
nor U3932 (N_3932,In_3336,In_3850);
and U3933 (N_3933,In_40,In_2276);
nor U3934 (N_3934,In_2395,In_4702);
and U3935 (N_3935,In_4617,In_3892);
nor U3936 (N_3936,In_1060,In_1641);
xor U3937 (N_3937,In_3715,In_1557);
nor U3938 (N_3938,In_1605,In_3897);
and U3939 (N_3939,In_1115,In_391);
nor U3940 (N_3940,In_2521,In_1727);
nor U3941 (N_3941,In_4082,In_4732);
nor U3942 (N_3942,In_4334,In_3585);
and U3943 (N_3943,In_3964,In_4168);
and U3944 (N_3944,In_1112,In_4129);
nand U3945 (N_3945,In_4991,In_381);
or U3946 (N_3946,In_3062,In_1975);
and U3947 (N_3947,In_4512,In_2991);
nor U3948 (N_3948,In_2727,In_1700);
nand U3949 (N_3949,In_4581,In_3101);
and U3950 (N_3950,In_687,In_4298);
nor U3951 (N_3951,In_3215,In_1556);
and U3952 (N_3952,In_2998,In_3899);
or U3953 (N_3953,In_3500,In_4176);
or U3954 (N_3954,In_3774,In_4286);
xnor U3955 (N_3955,In_2980,In_2675);
nand U3956 (N_3956,In_233,In_3629);
and U3957 (N_3957,In_513,In_4029);
nor U3958 (N_3958,In_3468,In_2381);
or U3959 (N_3959,In_3678,In_3059);
nand U3960 (N_3960,In_3028,In_2760);
xor U3961 (N_3961,In_1913,In_3170);
nand U3962 (N_3962,In_1010,In_1748);
nor U3963 (N_3963,In_1697,In_3120);
and U3964 (N_3964,In_2195,In_4456);
nor U3965 (N_3965,In_3727,In_683);
nor U3966 (N_3966,In_1478,In_3549);
and U3967 (N_3967,In_2433,In_4817);
xor U3968 (N_3968,In_4432,In_3218);
xnor U3969 (N_3969,In_4316,In_4199);
nor U3970 (N_3970,In_2494,In_2189);
or U3971 (N_3971,In_2077,In_3800);
and U3972 (N_3972,In_3883,In_1497);
nor U3973 (N_3973,In_2344,In_2125);
nand U3974 (N_3974,In_4141,In_4963);
nor U3975 (N_3975,In_3275,In_3680);
and U3976 (N_3976,In_1241,In_4587);
nor U3977 (N_3977,In_3893,In_4335);
nor U3978 (N_3978,In_1157,In_1443);
nand U3979 (N_3979,In_1049,In_1631);
and U3980 (N_3980,In_3928,In_1664);
nor U3981 (N_3981,In_3828,In_867);
xnor U3982 (N_3982,In_3502,In_1894);
and U3983 (N_3983,In_1184,In_3552);
xor U3984 (N_3984,In_66,In_2564);
nand U3985 (N_3985,In_1150,In_457);
nor U3986 (N_3986,In_347,In_1385);
or U3987 (N_3987,In_1458,In_1650);
nor U3988 (N_3988,In_4354,In_2574);
nand U3989 (N_3989,In_4504,In_3962);
nand U3990 (N_3990,In_376,In_1545);
xor U3991 (N_3991,In_1314,In_3742);
nand U3992 (N_3992,In_2598,In_1811);
or U3993 (N_3993,In_4958,In_4374);
and U3994 (N_3994,In_4349,In_1453);
nor U3995 (N_3995,In_3072,In_1429);
nor U3996 (N_3996,In_3860,In_4575);
nand U3997 (N_3997,In_2935,In_3901);
nand U3998 (N_3998,In_3918,In_2468);
or U3999 (N_3999,In_4092,In_491);
nand U4000 (N_4000,In_2341,In_2329);
nor U4001 (N_4001,In_4307,In_1106);
and U4002 (N_4002,In_4026,In_3682);
and U4003 (N_4003,In_4299,In_1800);
nand U4004 (N_4004,In_877,In_949);
and U4005 (N_4005,In_1949,In_1797);
and U4006 (N_4006,In_2190,In_2076);
nand U4007 (N_4007,In_3794,In_4583);
or U4008 (N_4008,In_1945,In_1382);
and U4009 (N_4009,In_226,In_475);
nor U4010 (N_4010,In_4871,In_1079);
and U4011 (N_4011,In_3084,In_16);
nor U4012 (N_4012,In_1369,In_2179);
nor U4013 (N_4013,In_2643,In_1127);
xor U4014 (N_4014,In_2143,In_1512);
nand U4015 (N_4015,In_1133,In_4126);
or U4016 (N_4016,In_2654,In_124);
nor U4017 (N_4017,In_381,In_558);
or U4018 (N_4018,In_1862,In_2241);
xnor U4019 (N_4019,In_3657,In_805);
nand U4020 (N_4020,In_2841,In_4146);
nand U4021 (N_4021,In_3406,In_980);
and U4022 (N_4022,In_4100,In_2969);
and U4023 (N_4023,In_1488,In_1017);
nor U4024 (N_4024,In_2911,In_4936);
nor U4025 (N_4025,In_3613,In_155);
xnor U4026 (N_4026,In_3194,In_2627);
nand U4027 (N_4027,In_3147,In_2862);
nand U4028 (N_4028,In_2675,In_2776);
or U4029 (N_4029,In_750,In_844);
nor U4030 (N_4030,In_3722,In_4814);
or U4031 (N_4031,In_4653,In_1372);
or U4032 (N_4032,In_322,In_2026);
nor U4033 (N_4033,In_1412,In_719);
and U4034 (N_4034,In_983,In_1303);
or U4035 (N_4035,In_2323,In_1650);
nand U4036 (N_4036,In_1394,In_3005);
and U4037 (N_4037,In_2496,In_4952);
and U4038 (N_4038,In_594,In_1747);
or U4039 (N_4039,In_4517,In_1254);
and U4040 (N_4040,In_4242,In_3610);
nand U4041 (N_4041,In_1486,In_3726);
and U4042 (N_4042,In_2247,In_3822);
or U4043 (N_4043,In_4397,In_789);
or U4044 (N_4044,In_4312,In_2840);
nand U4045 (N_4045,In_4732,In_713);
xor U4046 (N_4046,In_4720,In_495);
or U4047 (N_4047,In_1947,In_4505);
or U4048 (N_4048,In_1066,In_1742);
or U4049 (N_4049,In_1979,In_3157);
xor U4050 (N_4050,In_3948,In_2033);
nor U4051 (N_4051,In_2539,In_2061);
and U4052 (N_4052,In_3936,In_1731);
nand U4053 (N_4053,In_2659,In_3795);
nand U4054 (N_4054,In_1235,In_3236);
xor U4055 (N_4055,In_1754,In_2001);
or U4056 (N_4056,In_4354,In_2969);
xor U4057 (N_4057,In_4942,In_3094);
xnor U4058 (N_4058,In_1789,In_771);
and U4059 (N_4059,In_4153,In_4830);
nand U4060 (N_4060,In_944,In_3288);
or U4061 (N_4061,In_2866,In_3416);
or U4062 (N_4062,In_2485,In_4702);
or U4063 (N_4063,In_4777,In_4740);
nand U4064 (N_4064,In_655,In_384);
nand U4065 (N_4065,In_3041,In_876);
xnor U4066 (N_4066,In_3667,In_3706);
nand U4067 (N_4067,In_4198,In_2451);
nand U4068 (N_4068,In_2398,In_643);
nand U4069 (N_4069,In_986,In_1369);
and U4070 (N_4070,In_4109,In_3238);
nand U4071 (N_4071,In_1557,In_238);
or U4072 (N_4072,In_101,In_329);
or U4073 (N_4073,In_2640,In_4449);
or U4074 (N_4074,In_3023,In_149);
nor U4075 (N_4075,In_3420,In_4432);
nor U4076 (N_4076,In_3252,In_1645);
nand U4077 (N_4077,In_3413,In_3876);
nor U4078 (N_4078,In_3555,In_1499);
xnor U4079 (N_4079,In_692,In_4083);
nand U4080 (N_4080,In_3061,In_4675);
or U4081 (N_4081,In_483,In_2457);
or U4082 (N_4082,In_80,In_497);
and U4083 (N_4083,In_1854,In_986);
or U4084 (N_4084,In_2373,In_2336);
and U4085 (N_4085,In_3084,In_2265);
nor U4086 (N_4086,In_3946,In_4655);
and U4087 (N_4087,In_2517,In_2761);
xor U4088 (N_4088,In_1700,In_3072);
nand U4089 (N_4089,In_3062,In_3199);
nand U4090 (N_4090,In_1422,In_3789);
or U4091 (N_4091,In_3319,In_3492);
or U4092 (N_4092,In_4313,In_4808);
nand U4093 (N_4093,In_2880,In_3973);
nor U4094 (N_4094,In_284,In_1890);
or U4095 (N_4095,In_4148,In_4648);
xor U4096 (N_4096,In_988,In_4358);
nor U4097 (N_4097,In_4578,In_4783);
nand U4098 (N_4098,In_2816,In_2461);
and U4099 (N_4099,In_2125,In_2381);
nor U4100 (N_4100,In_1035,In_1368);
and U4101 (N_4101,In_2057,In_549);
or U4102 (N_4102,In_4654,In_4993);
nor U4103 (N_4103,In_4585,In_4973);
or U4104 (N_4104,In_4081,In_61);
xor U4105 (N_4105,In_4780,In_4733);
nor U4106 (N_4106,In_4605,In_1778);
or U4107 (N_4107,In_4753,In_4421);
and U4108 (N_4108,In_3198,In_4272);
nand U4109 (N_4109,In_99,In_825);
nand U4110 (N_4110,In_2139,In_399);
or U4111 (N_4111,In_1681,In_4667);
nor U4112 (N_4112,In_4554,In_1922);
and U4113 (N_4113,In_3808,In_4952);
or U4114 (N_4114,In_3021,In_935);
and U4115 (N_4115,In_547,In_3903);
nand U4116 (N_4116,In_3001,In_2748);
or U4117 (N_4117,In_1277,In_485);
or U4118 (N_4118,In_881,In_3409);
or U4119 (N_4119,In_1970,In_2402);
or U4120 (N_4120,In_2403,In_4766);
nor U4121 (N_4121,In_3994,In_1666);
or U4122 (N_4122,In_2791,In_2778);
and U4123 (N_4123,In_337,In_3581);
nand U4124 (N_4124,In_3098,In_759);
nand U4125 (N_4125,In_1372,In_4546);
and U4126 (N_4126,In_875,In_2736);
or U4127 (N_4127,In_3943,In_58);
nand U4128 (N_4128,In_4486,In_2435);
xnor U4129 (N_4129,In_822,In_3121);
nor U4130 (N_4130,In_4464,In_4823);
or U4131 (N_4131,In_2333,In_1578);
nand U4132 (N_4132,In_1868,In_3436);
or U4133 (N_4133,In_374,In_330);
and U4134 (N_4134,In_4641,In_2414);
nor U4135 (N_4135,In_2453,In_1714);
and U4136 (N_4136,In_4502,In_1884);
nor U4137 (N_4137,In_3161,In_4490);
nor U4138 (N_4138,In_373,In_3941);
and U4139 (N_4139,In_4731,In_2854);
and U4140 (N_4140,In_245,In_2111);
and U4141 (N_4141,In_256,In_2022);
xor U4142 (N_4142,In_2404,In_3900);
nor U4143 (N_4143,In_1009,In_1445);
and U4144 (N_4144,In_3308,In_2066);
or U4145 (N_4145,In_1957,In_1314);
nor U4146 (N_4146,In_1383,In_3865);
nand U4147 (N_4147,In_984,In_597);
nor U4148 (N_4148,In_2962,In_3909);
or U4149 (N_4149,In_3693,In_1517);
nor U4150 (N_4150,In_624,In_2642);
or U4151 (N_4151,In_13,In_2543);
nand U4152 (N_4152,In_3261,In_4915);
nor U4153 (N_4153,In_1654,In_2564);
or U4154 (N_4154,In_129,In_715);
nand U4155 (N_4155,In_1187,In_2911);
nor U4156 (N_4156,In_438,In_1396);
or U4157 (N_4157,In_1521,In_3615);
nor U4158 (N_4158,In_3392,In_3659);
nor U4159 (N_4159,In_2514,In_3278);
nand U4160 (N_4160,In_4065,In_681);
and U4161 (N_4161,In_3407,In_4806);
nor U4162 (N_4162,In_2450,In_2272);
xor U4163 (N_4163,In_1298,In_2077);
nand U4164 (N_4164,In_2773,In_251);
nor U4165 (N_4165,In_4135,In_352);
or U4166 (N_4166,In_1635,In_3256);
and U4167 (N_4167,In_2207,In_3554);
and U4168 (N_4168,In_1013,In_3339);
nor U4169 (N_4169,In_2449,In_1772);
nor U4170 (N_4170,In_3846,In_3947);
nor U4171 (N_4171,In_3104,In_2341);
and U4172 (N_4172,In_4246,In_4324);
or U4173 (N_4173,In_2636,In_1151);
or U4174 (N_4174,In_3323,In_2890);
or U4175 (N_4175,In_1080,In_2326);
or U4176 (N_4176,In_172,In_3593);
nand U4177 (N_4177,In_3172,In_1497);
nor U4178 (N_4178,In_251,In_4877);
and U4179 (N_4179,In_4399,In_912);
nand U4180 (N_4180,In_220,In_518);
xor U4181 (N_4181,In_4677,In_3436);
xor U4182 (N_4182,In_3883,In_1783);
nand U4183 (N_4183,In_4965,In_2668);
and U4184 (N_4184,In_3323,In_2256);
xnor U4185 (N_4185,In_1262,In_3999);
xor U4186 (N_4186,In_1912,In_4236);
nor U4187 (N_4187,In_190,In_1280);
or U4188 (N_4188,In_3404,In_2275);
or U4189 (N_4189,In_4847,In_4355);
or U4190 (N_4190,In_2912,In_4856);
xor U4191 (N_4191,In_4481,In_1002);
and U4192 (N_4192,In_364,In_579);
xnor U4193 (N_4193,In_1369,In_208);
and U4194 (N_4194,In_1685,In_3107);
and U4195 (N_4195,In_1451,In_3754);
and U4196 (N_4196,In_3386,In_1788);
nand U4197 (N_4197,In_821,In_3479);
nor U4198 (N_4198,In_625,In_2944);
or U4199 (N_4199,In_3672,In_4842);
nor U4200 (N_4200,In_730,In_2481);
nand U4201 (N_4201,In_3587,In_366);
nand U4202 (N_4202,In_4996,In_3157);
nor U4203 (N_4203,In_3349,In_11);
or U4204 (N_4204,In_4933,In_2555);
or U4205 (N_4205,In_127,In_1534);
xor U4206 (N_4206,In_3417,In_791);
xnor U4207 (N_4207,In_1877,In_3773);
nor U4208 (N_4208,In_1074,In_647);
nor U4209 (N_4209,In_4099,In_4918);
and U4210 (N_4210,In_3215,In_3081);
nor U4211 (N_4211,In_1797,In_3098);
xnor U4212 (N_4212,In_3579,In_4601);
or U4213 (N_4213,In_4262,In_2093);
and U4214 (N_4214,In_3764,In_827);
or U4215 (N_4215,In_1599,In_1529);
nand U4216 (N_4216,In_1846,In_4090);
nand U4217 (N_4217,In_2238,In_2057);
and U4218 (N_4218,In_228,In_777);
nor U4219 (N_4219,In_672,In_3884);
and U4220 (N_4220,In_3611,In_131);
xor U4221 (N_4221,In_2663,In_1237);
nand U4222 (N_4222,In_2081,In_2683);
and U4223 (N_4223,In_1367,In_2087);
nand U4224 (N_4224,In_4273,In_2929);
nor U4225 (N_4225,In_2064,In_3090);
or U4226 (N_4226,In_565,In_4756);
or U4227 (N_4227,In_3721,In_3697);
nor U4228 (N_4228,In_1089,In_1224);
nand U4229 (N_4229,In_1223,In_2443);
xnor U4230 (N_4230,In_1998,In_3941);
and U4231 (N_4231,In_2346,In_412);
or U4232 (N_4232,In_841,In_3108);
xor U4233 (N_4233,In_1661,In_541);
or U4234 (N_4234,In_2131,In_274);
or U4235 (N_4235,In_105,In_1244);
nor U4236 (N_4236,In_3282,In_408);
and U4237 (N_4237,In_3888,In_4500);
and U4238 (N_4238,In_1518,In_1345);
and U4239 (N_4239,In_4643,In_4513);
nor U4240 (N_4240,In_1085,In_4103);
and U4241 (N_4241,In_740,In_3326);
and U4242 (N_4242,In_4278,In_246);
xnor U4243 (N_4243,In_898,In_4348);
nand U4244 (N_4244,In_2524,In_2671);
or U4245 (N_4245,In_1342,In_4696);
and U4246 (N_4246,In_2458,In_2109);
and U4247 (N_4247,In_4914,In_821);
nor U4248 (N_4248,In_4835,In_265);
nand U4249 (N_4249,In_738,In_1481);
nand U4250 (N_4250,In_663,In_3961);
nor U4251 (N_4251,In_1864,In_3034);
nand U4252 (N_4252,In_1407,In_1818);
or U4253 (N_4253,In_3043,In_2680);
xnor U4254 (N_4254,In_3673,In_47);
and U4255 (N_4255,In_1897,In_290);
nand U4256 (N_4256,In_674,In_1937);
nor U4257 (N_4257,In_3088,In_2176);
xnor U4258 (N_4258,In_2064,In_1599);
nand U4259 (N_4259,In_4613,In_4678);
and U4260 (N_4260,In_861,In_4498);
nor U4261 (N_4261,In_4500,In_124);
nand U4262 (N_4262,In_1593,In_77);
nor U4263 (N_4263,In_3080,In_1110);
or U4264 (N_4264,In_255,In_688);
nor U4265 (N_4265,In_717,In_1111);
or U4266 (N_4266,In_259,In_2320);
and U4267 (N_4267,In_4263,In_1780);
xor U4268 (N_4268,In_3265,In_2658);
and U4269 (N_4269,In_3820,In_1190);
nand U4270 (N_4270,In_3087,In_2735);
and U4271 (N_4271,In_2486,In_4221);
nor U4272 (N_4272,In_4195,In_2687);
nor U4273 (N_4273,In_1280,In_1020);
nor U4274 (N_4274,In_906,In_3644);
or U4275 (N_4275,In_3303,In_2810);
and U4276 (N_4276,In_2271,In_1274);
or U4277 (N_4277,In_2330,In_4796);
and U4278 (N_4278,In_2695,In_1761);
and U4279 (N_4279,In_89,In_168);
or U4280 (N_4280,In_2130,In_3125);
or U4281 (N_4281,In_4344,In_2082);
nand U4282 (N_4282,In_1611,In_3658);
nor U4283 (N_4283,In_3728,In_1151);
xnor U4284 (N_4284,In_3031,In_1566);
or U4285 (N_4285,In_2863,In_4183);
xnor U4286 (N_4286,In_890,In_1530);
or U4287 (N_4287,In_1809,In_1298);
nand U4288 (N_4288,In_3589,In_4683);
nor U4289 (N_4289,In_615,In_792);
nor U4290 (N_4290,In_1499,In_970);
or U4291 (N_4291,In_3626,In_1095);
or U4292 (N_4292,In_937,In_3919);
nor U4293 (N_4293,In_2023,In_1440);
and U4294 (N_4294,In_3109,In_742);
or U4295 (N_4295,In_3798,In_3886);
nand U4296 (N_4296,In_1508,In_4661);
nor U4297 (N_4297,In_4376,In_2119);
nand U4298 (N_4298,In_683,In_2696);
or U4299 (N_4299,In_1583,In_860);
or U4300 (N_4300,In_1409,In_1852);
or U4301 (N_4301,In_1579,In_638);
and U4302 (N_4302,In_1879,In_557);
or U4303 (N_4303,In_1572,In_4013);
xor U4304 (N_4304,In_2006,In_1898);
or U4305 (N_4305,In_2985,In_1798);
nand U4306 (N_4306,In_2447,In_1689);
or U4307 (N_4307,In_1600,In_3255);
and U4308 (N_4308,In_4964,In_1166);
nand U4309 (N_4309,In_1051,In_693);
nand U4310 (N_4310,In_336,In_1188);
xor U4311 (N_4311,In_5,In_4484);
nand U4312 (N_4312,In_3907,In_388);
nand U4313 (N_4313,In_84,In_1100);
or U4314 (N_4314,In_32,In_1723);
or U4315 (N_4315,In_1772,In_1963);
or U4316 (N_4316,In_1802,In_3916);
xor U4317 (N_4317,In_4176,In_1531);
or U4318 (N_4318,In_1638,In_2437);
or U4319 (N_4319,In_1571,In_3573);
nand U4320 (N_4320,In_1534,In_326);
nand U4321 (N_4321,In_545,In_3886);
nor U4322 (N_4322,In_455,In_2000);
and U4323 (N_4323,In_3002,In_1590);
and U4324 (N_4324,In_194,In_1235);
xnor U4325 (N_4325,In_3041,In_2390);
or U4326 (N_4326,In_3776,In_1029);
nand U4327 (N_4327,In_66,In_4673);
nand U4328 (N_4328,In_80,In_2465);
nor U4329 (N_4329,In_2200,In_2190);
xor U4330 (N_4330,In_3243,In_2061);
and U4331 (N_4331,In_4174,In_4504);
nor U4332 (N_4332,In_3249,In_2777);
nand U4333 (N_4333,In_3251,In_2400);
or U4334 (N_4334,In_1688,In_1187);
xor U4335 (N_4335,In_3182,In_4929);
nand U4336 (N_4336,In_238,In_1996);
and U4337 (N_4337,In_2130,In_4540);
xnor U4338 (N_4338,In_4686,In_488);
and U4339 (N_4339,In_1324,In_3891);
nand U4340 (N_4340,In_2029,In_504);
or U4341 (N_4341,In_4916,In_944);
nor U4342 (N_4342,In_273,In_2221);
and U4343 (N_4343,In_202,In_3199);
or U4344 (N_4344,In_1078,In_3521);
or U4345 (N_4345,In_2238,In_3827);
xor U4346 (N_4346,In_601,In_3052);
xor U4347 (N_4347,In_4684,In_1130);
or U4348 (N_4348,In_1221,In_3748);
and U4349 (N_4349,In_3245,In_4003);
and U4350 (N_4350,In_775,In_3811);
nand U4351 (N_4351,In_3426,In_3489);
and U4352 (N_4352,In_4354,In_979);
nand U4353 (N_4353,In_3320,In_2096);
xor U4354 (N_4354,In_648,In_1143);
and U4355 (N_4355,In_813,In_4379);
and U4356 (N_4356,In_471,In_1145);
nand U4357 (N_4357,In_3047,In_3617);
nand U4358 (N_4358,In_1280,In_3131);
nand U4359 (N_4359,In_4148,In_1977);
nand U4360 (N_4360,In_52,In_302);
nor U4361 (N_4361,In_3015,In_2057);
or U4362 (N_4362,In_3573,In_1638);
nand U4363 (N_4363,In_1051,In_2919);
or U4364 (N_4364,In_2492,In_1837);
nor U4365 (N_4365,In_1395,In_3797);
nand U4366 (N_4366,In_1797,In_1833);
and U4367 (N_4367,In_4270,In_831);
or U4368 (N_4368,In_4792,In_3950);
nand U4369 (N_4369,In_613,In_1522);
xnor U4370 (N_4370,In_403,In_1881);
and U4371 (N_4371,In_3915,In_2410);
and U4372 (N_4372,In_1977,In_2263);
and U4373 (N_4373,In_3110,In_3864);
nand U4374 (N_4374,In_4351,In_3349);
and U4375 (N_4375,In_1485,In_4952);
nor U4376 (N_4376,In_2488,In_1956);
or U4377 (N_4377,In_3323,In_303);
nand U4378 (N_4378,In_2342,In_1310);
or U4379 (N_4379,In_4402,In_2440);
and U4380 (N_4380,In_2760,In_3121);
nor U4381 (N_4381,In_4238,In_2114);
nand U4382 (N_4382,In_4211,In_2161);
xor U4383 (N_4383,In_1151,In_1926);
xor U4384 (N_4384,In_3772,In_21);
or U4385 (N_4385,In_4611,In_3275);
nor U4386 (N_4386,In_1697,In_4790);
or U4387 (N_4387,In_1151,In_2327);
and U4388 (N_4388,In_921,In_337);
nand U4389 (N_4389,In_4709,In_2946);
or U4390 (N_4390,In_4317,In_1056);
or U4391 (N_4391,In_577,In_2631);
nor U4392 (N_4392,In_4609,In_234);
nand U4393 (N_4393,In_1955,In_4955);
nor U4394 (N_4394,In_3191,In_1503);
xor U4395 (N_4395,In_1897,In_4395);
xnor U4396 (N_4396,In_2839,In_2272);
and U4397 (N_4397,In_3527,In_4569);
nand U4398 (N_4398,In_4402,In_1740);
and U4399 (N_4399,In_2575,In_2556);
and U4400 (N_4400,In_3516,In_2535);
or U4401 (N_4401,In_3224,In_2291);
xor U4402 (N_4402,In_123,In_4935);
nand U4403 (N_4403,In_4332,In_2333);
nand U4404 (N_4404,In_4997,In_2706);
and U4405 (N_4405,In_4795,In_3393);
or U4406 (N_4406,In_621,In_2369);
and U4407 (N_4407,In_1104,In_1961);
nor U4408 (N_4408,In_3783,In_2067);
nand U4409 (N_4409,In_1828,In_4066);
nor U4410 (N_4410,In_3012,In_790);
nor U4411 (N_4411,In_1255,In_4515);
nor U4412 (N_4412,In_3030,In_4608);
or U4413 (N_4413,In_4504,In_2901);
or U4414 (N_4414,In_1007,In_1491);
nand U4415 (N_4415,In_1188,In_4620);
nand U4416 (N_4416,In_4081,In_619);
nor U4417 (N_4417,In_1495,In_3686);
or U4418 (N_4418,In_2628,In_2275);
nand U4419 (N_4419,In_1753,In_4445);
nand U4420 (N_4420,In_2539,In_3913);
nor U4421 (N_4421,In_2196,In_2024);
nor U4422 (N_4422,In_4293,In_1019);
or U4423 (N_4423,In_1126,In_343);
xor U4424 (N_4424,In_4223,In_2372);
nand U4425 (N_4425,In_3874,In_2631);
and U4426 (N_4426,In_2755,In_2077);
nand U4427 (N_4427,In_4403,In_3913);
nand U4428 (N_4428,In_3877,In_3629);
nor U4429 (N_4429,In_1132,In_922);
or U4430 (N_4430,In_248,In_2993);
and U4431 (N_4431,In_4431,In_1867);
and U4432 (N_4432,In_263,In_4026);
nor U4433 (N_4433,In_644,In_4543);
and U4434 (N_4434,In_164,In_4375);
nand U4435 (N_4435,In_4467,In_4605);
nand U4436 (N_4436,In_1593,In_94);
or U4437 (N_4437,In_3498,In_3335);
or U4438 (N_4438,In_3599,In_2837);
or U4439 (N_4439,In_554,In_3180);
and U4440 (N_4440,In_3880,In_1326);
or U4441 (N_4441,In_4885,In_409);
nor U4442 (N_4442,In_450,In_1773);
xor U4443 (N_4443,In_402,In_338);
nand U4444 (N_4444,In_2090,In_4730);
xor U4445 (N_4445,In_2833,In_4286);
or U4446 (N_4446,In_1782,In_1072);
nand U4447 (N_4447,In_3581,In_3189);
and U4448 (N_4448,In_2654,In_4579);
nor U4449 (N_4449,In_794,In_4635);
xor U4450 (N_4450,In_2403,In_734);
and U4451 (N_4451,In_3619,In_3482);
and U4452 (N_4452,In_2332,In_1325);
nand U4453 (N_4453,In_2093,In_2051);
or U4454 (N_4454,In_4622,In_3120);
or U4455 (N_4455,In_2673,In_1583);
xor U4456 (N_4456,In_488,In_1564);
xor U4457 (N_4457,In_1799,In_2183);
nor U4458 (N_4458,In_1546,In_4075);
nand U4459 (N_4459,In_4675,In_3233);
and U4460 (N_4460,In_2045,In_288);
nand U4461 (N_4461,In_3282,In_2936);
and U4462 (N_4462,In_3853,In_212);
nor U4463 (N_4463,In_1859,In_2331);
and U4464 (N_4464,In_4792,In_3826);
nor U4465 (N_4465,In_3302,In_906);
nand U4466 (N_4466,In_579,In_3084);
xnor U4467 (N_4467,In_4256,In_3586);
nor U4468 (N_4468,In_3820,In_241);
or U4469 (N_4469,In_3610,In_3204);
nor U4470 (N_4470,In_3572,In_3921);
or U4471 (N_4471,In_729,In_4367);
nor U4472 (N_4472,In_2181,In_1118);
or U4473 (N_4473,In_1142,In_3744);
nor U4474 (N_4474,In_1318,In_4646);
nand U4475 (N_4475,In_3315,In_2286);
and U4476 (N_4476,In_2669,In_4951);
and U4477 (N_4477,In_346,In_3974);
nor U4478 (N_4478,In_1276,In_1138);
and U4479 (N_4479,In_3790,In_3983);
nor U4480 (N_4480,In_3257,In_1874);
and U4481 (N_4481,In_1958,In_2358);
nor U4482 (N_4482,In_3170,In_3883);
or U4483 (N_4483,In_1629,In_416);
or U4484 (N_4484,In_643,In_4769);
or U4485 (N_4485,In_1303,In_883);
nand U4486 (N_4486,In_1035,In_1290);
nor U4487 (N_4487,In_4092,In_1568);
nor U4488 (N_4488,In_2084,In_2028);
or U4489 (N_4489,In_750,In_756);
xor U4490 (N_4490,In_2095,In_3981);
nand U4491 (N_4491,In_1776,In_260);
and U4492 (N_4492,In_1943,In_2269);
nand U4493 (N_4493,In_840,In_1551);
nand U4494 (N_4494,In_2307,In_802);
or U4495 (N_4495,In_3323,In_3855);
nand U4496 (N_4496,In_2349,In_2954);
or U4497 (N_4497,In_4333,In_1622);
nand U4498 (N_4498,In_4840,In_3624);
nor U4499 (N_4499,In_4340,In_1564);
nor U4500 (N_4500,In_3178,In_348);
nor U4501 (N_4501,In_1866,In_1234);
xnor U4502 (N_4502,In_2664,In_1709);
nor U4503 (N_4503,In_4308,In_4930);
nor U4504 (N_4504,In_939,In_3199);
and U4505 (N_4505,In_1672,In_363);
nor U4506 (N_4506,In_4215,In_1558);
xor U4507 (N_4507,In_1895,In_4486);
nand U4508 (N_4508,In_4310,In_3663);
nor U4509 (N_4509,In_4600,In_3388);
and U4510 (N_4510,In_1860,In_2154);
or U4511 (N_4511,In_4774,In_1242);
and U4512 (N_4512,In_4370,In_500);
xor U4513 (N_4513,In_4187,In_3253);
xor U4514 (N_4514,In_2617,In_1515);
or U4515 (N_4515,In_4957,In_2232);
nand U4516 (N_4516,In_2743,In_4994);
or U4517 (N_4517,In_3884,In_264);
nor U4518 (N_4518,In_3913,In_3677);
or U4519 (N_4519,In_4933,In_2710);
nor U4520 (N_4520,In_938,In_951);
xnor U4521 (N_4521,In_4335,In_0);
and U4522 (N_4522,In_4240,In_2585);
nand U4523 (N_4523,In_1486,In_569);
nand U4524 (N_4524,In_1119,In_573);
nand U4525 (N_4525,In_3852,In_2744);
nand U4526 (N_4526,In_4983,In_2575);
nor U4527 (N_4527,In_1250,In_2313);
and U4528 (N_4528,In_270,In_2332);
nand U4529 (N_4529,In_1675,In_4799);
nor U4530 (N_4530,In_4024,In_1353);
xnor U4531 (N_4531,In_475,In_2794);
and U4532 (N_4532,In_659,In_79);
nand U4533 (N_4533,In_3053,In_1938);
or U4534 (N_4534,In_4750,In_4363);
nand U4535 (N_4535,In_3546,In_2764);
nand U4536 (N_4536,In_1356,In_3362);
xor U4537 (N_4537,In_150,In_4544);
and U4538 (N_4538,In_331,In_2658);
nand U4539 (N_4539,In_3479,In_2183);
nor U4540 (N_4540,In_1585,In_2493);
or U4541 (N_4541,In_1568,In_4113);
nor U4542 (N_4542,In_3370,In_2186);
nor U4543 (N_4543,In_1600,In_2678);
nand U4544 (N_4544,In_3232,In_991);
nand U4545 (N_4545,In_185,In_4051);
or U4546 (N_4546,In_915,In_646);
nand U4547 (N_4547,In_2334,In_1065);
and U4548 (N_4548,In_2081,In_474);
and U4549 (N_4549,In_2503,In_2572);
and U4550 (N_4550,In_1564,In_483);
nand U4551 (N_4551,In_1936,In_3002);
and U4552 (N_4552,In_509,In_3193);
or U4553 (N_4553,In_54,In_2469);
nor U4554 (N_4554,In_80,In_4448);
xor U4555 (N_4555,In_2336,In_1571);
or U4556 (N_4556,In_3180,In_2355);
and U4557 (N_4557,In_2416,In_102);
nor U4558 (N_4558,In_3201,In_2391);
nand U4559 (N_4559,In_4280,In_3407);
nor U4560 (N_4560,In_549,In_3181);
or U4561 (N_4561,In_529,In_3822);
nand U4562 (N_4562,In_3899,In_62);
and U4563 (N_4563,In_2949,In_4476);
nand U4564 (N_4564,In_4654,In_3508);
and U4565 (N_4565,In_4639,In_2736);
xor U4566 (N_4566,In_189,In_4639);
xor U4567 (N_4567,In_4781,In_4769);
nand U4568 (N_4568,In_4753,In_3435);
and U4569 (N_4569,In_1293,In_3046);
xor U4570 (N_4570,In_3633,In_3736);
and U4571 (N_4571,In_1907,In_4017);
nand U4572 (N_4572,In_4405,In_1899);
nor U4573 (N_4573,In_3311,In_4963);
or U4574 (N_4574,In_4289,In_1644);
or U4575 (N_4575,In_395,In_3261);
nor U4576 (N_4576,In_1014,In_4366);
and U4577 (N_4577,In_573,In_1424);
or U4578 (N_4578,In_3952,In_236);
and U4579 (N_4579,In_2594,In_76);
xor U4580 (N_4580,In_4646,In_3014);
xor U4581 (N_4581,In_3784,In_4520);
or U4582 (N_4582,In_1969,In_14);
nor U4583 (N_4583,In_4876,In_361);
nand U4584 (N_4584,In_2021,In_3743);
or U4585 (N_4585,In_846,In_3222);
and U4586 (N_4586,In_3071,In_4351);
or U4587 (N_4587,In_4202,In_1080);
or U4588 (N_4588,In_2126,In_1515);
or U4589 (N_4589,In_2408,In_3582);
and U4590 (N_4590,In_2785,In_57);
and U4591 (N_4591,In_3459,In_2878);
and U4592 (N_4592,In_84,In_3058);
nor U4593 (N_4593,In_1041,In_2022);
nor U4594 (N_4594,In_3869,In_2788);
nor U4595 (N_4595,In_1946,In_227);
nor U4596 (N_4596,In_4966,In_60);
and U4597 (N_4597,In_2121,In_204);
and U4598 (N_4598,In_2871,In_3970);
xor U4599 (N_4599,In_4589,In_4890);
or U4600 (N_4600,In_4820,In_4960);
and U4601 (N_4601,In_3335,In_4918);
and U4602 (N_4602,In_3014,In_3599);
and U4603 (N_4603,In_2062,In_819);
nor U4604 (N_4604,In_888,In_3448);
nor U4605 (N_4605,In_922,In_834);
xor U4606 (N_4606,In_2398,In_2592);
nor U4607 (N_4607,In_4102,In_367);
nand U4608 (N_4608,In_4505,In_534);
xor U4609 (N_4609,In_4966,In_1935);
xnor U4610 (N_4610,In_3910,In_2283);
xnor U4611 (N_4611,In_4431,In_4161);
nor U4612 (N_4612,In_4286,In_1551);
and U4613 (N_4613,In_2338,In_2118);
nor U4614 (N_4614,In_1571,In_2828);
nor U4615 (N_4615,In_236,In_3862);
nor U4616 (N_4616,In_4551,In_4695);
and U4617 (N_4617,In_3407,In_4640);
or U4618 (N_4618,In_4243,In_222);
nand U4619 (N_4619,In_1704,In_1139);
or U4620 (N_4620,In_2884,In_1121);
nor U4621 (N_4621,In_3632,In_3966);
nor U4622 (N_4622,In_1016,In_2745);
nand U4623 (N_4623,In_3076,In_833);
nor U4624 (N_4624,In_243,In_3207);
xor U4625 (N_4625,In_413,In_2519);
nand U4626 (N_4626,In_4574,In_1383);
or U4627 (N_4627,In_2384,In_4494);
nand U4628 (N_4628,In_844,In_2241);
or U4629 (N_4629,In_1321,In_2481);
nand U4630 (N_4630,In_4895,In_467);
or U4631 (N_4631,In_1999,In_4533);
nor U4632 (N_4632,In_975,In_1927);
or U4633 (N_4633,In_4336,In_3065);
nand U4634 (N_4634,In_1697,In_1157);
nand U4635 (N_4635,In_1224,In_2787);
nand U4636 (N_4636,In_3832,In_1577);
nor U4637 (N_4637,In_2721,In_145);
nor U4638 (N_4638,In_4651,In_2891);
and U4639 (N_4639,In_563,In_1863);
nor U4640 (N_4640,In_4764,In_1883);
or U4641 (N_4641,In_3928,In_2888);
nand U4642 (N_4642,In_1490,In_437);
nor U4643 (N_4643,In_150,In_1613);
or U4644 (N_4644,In_1256,In_1359);
nand U4645 (N_4645,In_4240,In_1897);
and U4646 (N_4646,In_2418,In_1517);
nand U4647 (N_4647,In_994,In_3046);
nand U4648 (N_4648,In_752,In_3879);
xnor U4649 (N_4649,In_109,In_1951);
and U4650 (N_4650,In_2412,In_1993);
or U4651 (N_4651,In_1512,In_4807);
nor U4652 (N_4652,In_2211,In_4248);
or U4653 (N_4653,In_2445,In_950);
nand U4654 (N_4654,In_1013,In_1528);
or U4655 (N_4655,In_516,In_668);
and U4656 (N_4656,In_4987,In_4410);
nor U4657 (N_4657,In_1148,In_1313);
nand U4658 (N_4658,In_435,In_2895);
and U4659 (N_4659,In_1746,In_819);
or U4660 (N_4660,In_4229,In_3534);
and U4661 (N_4661,In_2632,In_4105);
nor U4662 (N_4662,In_2555,In_3027);
nand U4663 (N_4663,In_3075,In_4518);
and U4664 (N_4664,In_1234,In_4169);
xor U4665 (N_4665,In_673,In_1223);
and U4666 (N_4666,In_3677,In_2340);
xor U4667 (N_4667,In_3091,In_3151);
and U4668 (N_4668,In_2912,In_2530);
nand U4669 (N_4669,In_1050,In_4998);
or U4670 (N_4670,In_2912,In_2748);
xor U4671 (N_4671,In_1012,In_3393);
and U4672 (N_4672,In_4588,In_1640);
and U4673 (N_4673,In_1331,In_1918);
nor U4674 (N_4674,In_4274,In_4243);
nor U4675 (N_4675,In_2984,In_4221);
nand U4676 (N_4676,In_2752,In_3117);
nand U4677 (N_4677,In_331,In_3664);
or U4678 (N_4678,In_756,In_2642);
nand U4679 (N_4679,In_732,In_4671);
nand U4680 (N_4680,In_3786,In_1248);
nor U4681 (N_4681,In_2769,In_841);
nor U4682 (N_4682,In_678,In_429);
nor U4683 (N_4683,In_3573,In_4694);
and U4684 (N_4684,In_2919,In_4179);
xor U4685 (N_4685,In_4251,In_4951);
and U4686 (N_4686,In_2822,In_1918);
and U4687 (N_4687,In_2160,In_2357);
nand U4688 (N_4688,In_1170,In_961);
and U4689 (N_4689,In_3534,In_906);
or U4690 (N_4690,In_4043,In_2051);
nor U4691 (N_4691,In_3824,In_803);
nand U4692 (N_4692,In_1946,In_288);
or U4693 (N_4693,In_3465,In_356);
nor U4694 (N_4694,In_1716,In_3454);
nand U4695 (N_4695,In_914,In_456);
or U4696 (N_4696,In_1354,In_3332);
or U4697 (N_4697,In_2464,In_2421);
nand U4698 (N_4698,In_3259,In_4508);
nor U4699 (N_4699,In_1382,In_4785);
and U4700 (N_4700,In_4681,In_1384);
and U4701 (N_4701,In_3382,In_2781);
nor U4702 (N_4702,In_4117,In_4175);
and U4703 (N_4703,In_622,In_4788);
and U4704 (N_4704,In_2115,In_3892);
and U4705 (N_4705,In_3556,In_602);
and U4706 (N_4706,In_4951,In_1480);
or U4707 (N_4707,In_3933,In_3185);
xor U4708 (N_4708,In_284,In_3893);
and U4709 (N_4709,In_1323,In_2108);
nor U4710 (N_4710,In_99,In_2160);
or U4711 (N_4711,In_1648,In_4737);
nor U4712 (N_4712,In_2322,In_1467);
nor U4713 (N_4713,In_2480,In_3055);
nor U4714 (N_4714,In_904,In_4947);
nand U4715 (N_4715,In_2028,In_2894);
and U4716 (N_4716,In_2304,In_4697);
or U4717 (N_4717,In_1233,In_3662);
nor U4718 (N_4718,In_115,In_1771);
nand U4719 (N_4719,In_4569,In_3976);
xnor U4720 (N_4720,In_4097,In_2942);
nor U4721 (N_4721,In_804,In_2117);
or U4722 (N_4722,In_4223,In_1096);
xor U4723 (N_4723,In_3587,In_4419);
nor U4724 (N_4724,In_2528,In_4186);
nand U4725 (N_4725,In_926,In_123);
nor U4726 (N_4726,In_4450,In_4316);
or U4727 (N_4727,In_3886,In_1386);
or U4728 (N_4728,In_2300,In_2069);
and U4729 (N_4729,In_102,In_1036);
nand U4730 (N_4730,In_1460,In_4839);
xor U4731 (N_4731,In_1588,In_1800);
xnor U4732 (N_4732,In_4408,In_3047);
nand U4733 (N_4733,In_4418,In_1079);
and U4734 (N_4734,In_1701,In_2672);
xnor U4735 (N_4735,In_3559,In_451);
and U4736 (N_4736,In_4463,In_585);
nor U4737 (N_4737,In_3787,In_1386);
nand U4738 (N_4738,In_1530,In_3706);
nor U4739 (N_4739,In_4166,In_3152);
nor U4740 (N_4740,In_4176,In_2352);
or U4741 (N_4741,In_1517,In_4885);
nor U4742 (N_4742,In_3021,In_1623);
and U4743 (N_4743,In_3649,In_3316);
or U4744 (N_4744,In_11,In_2862);
or U4745 (N_4745,In_2117,In_3049);
and U4746 (N_4746,In_872,In_3474);
nor U4747 (N_4747,In_627,In_37);
nand U4748 (N_4748,In_234,In_311);
nand U4749 (N_4749,In_3133,In_4724);
nor U4750 (N_4750,In_3009,In_3625);
or U4751 (N_4751,In_4645,In_2254);
and U4752 (N_4752,In_3080,In_126);
xnor U4753 (N_4753,In_4386,In_2641);
and U4754 (N_4754,In_2759,In_2682);
xnor U4755 (N_4755,In_709,In_1868);
nor U4756 (N_4756,In_1996,In_3813);
or U4757 (N_4757,In_3085,In_2452);
and U4758 (N_4758,In_1159,In_3419);
nand U4759 (N_4759,In_4341,In_3957);
and U4760 (N_4760,In_2718,In_1693);
and U4761 (N_4761,In_2579,In_3369);
or U4762 (N_4762,In_816,In_2864);
or U4763 (N_4763,In_3057,In_1825);
and U4764 (N_4764,In_783,In_4935);
xor U4765 (N_4765,In_1061,In_4268);
and U4766 (N_4766,In_3926,In_4816);
and U4767 (N_4767,In_1232,In_1412);
nor U4768 (N_4768,In_1792,In_2159);
and U4769 (N_4769,In_3814,In_425);
nor U4770 (N_4770,In_3478,In_952);
and U4771 (N_4771,In_3406,In_484);
nand U4772 (N_4772,In_2187,In_2893);
and U4773 (N_4773,In_12,In_1796);
and U4774 (N_4774,In_1998,In_616);
or U4775 (N_4775,In_1408,In_912);
and U4776 (N_4776,In_2127,In_867);
nand U4777 (N_4777,In_3087,In_912);
and U4778 (N_4778,In_587,In_2734);
xnor U4779 (N_4779,In_1896,In_2883);
nor U4780 (N_4780,In_2050,In_3595);
or U4781 (N_4781,In_460,In_4680);
or U4782 (N_4782,In_2623,In_1867);
nand U4783 (N_4783,In_2849,In_3391);
nand U4784 (N_4784,In_3805,In_1342);
nor U4785 (N_4785,In_313,In_4293);
nor U4786 (N_4786,In_3557,In_706);
or U4787 (N_4787,In_932,In_4929);
and U4788 (N_4788,In_4079,In_1039);
or U4789 (N_4789,In_1531,In_1364);
or U4790 (N_4790,In_1569,In_4186);
nor U4791 (N_4791,In_839,In_128);
and U4792 (N_4792,In_2669,In_2729);
or U4793 (N_4793,In_3214,In_3775);
and U4794 (N_4794,In_1006,In_3926);
nand U4795 (N_4795,In_3496,In_4411);
and U4796 (N_4796,In_385,In_2947);
nor U4797 (N_4797,In_4307,In_4193);
nor U4798 (N_4798,In_748,In_4047);
nand U4799 (N_4799,In_371,In_549);
xnor U4800 (N_4800,In_4019,In_4313);
and U4801 (N_4801,In_3071,In_28);
and U4802 (N_4802,In_579,In_1318);
or U4803 (N_4803,In_3262,In_2325);
or U4804 (N_4804,In_1588,In_4957);
xnor U4805 (N_4805,In_3210,In_127);
and U4806 (N_4806,In_2506,In_728);
nand U4807 (N_4807,In_617,In_2913);
and U4808 (N_4808,In_2141,In_1988);
and U4809 (N_4809,In_1003,In_2625);
nand U4810 (N_4810,In_3771,In_4173);
and U4811 (N_4811,In_3200,In_3043);
nand U4812 (N_4812,In_4089,In_3160);
nand U4813 (N_4813,In_3328,In_3751);
nor U4814 (N_4814,In_2571,In_1939);
or U4815 (N_4815,In_2939,In_3715);
and U4816 (N_4816,In_3271,In_4083);
xnor U4817 (N_4817,In_1152,In_3026);
nor U4818 (N_4818,In_542,In_2820);
nor U4819 (N_4819,In_2183,In_3083);
and U4820 (N_4820,In_3686,In_2092);
or U4821 (N_4821,In_1907,In_3630);
nor U4822 (N_4822,In_3103,In_762);
and U4823 (N_4823,In_3591,In_1907);
nand U4824 (N_4824,In_2180,In_2957);
nand U4825 (N_4825,In_1935,In_1824);
and U4826 (N_4826,In_2346,In_2764);
or U4827 (N_4827,In_3132,In_409);
and U4828 (N_4828,In_1332,In_2018);
or U4829 (N_4829,In_4606,In_2319);
nand U4830 (N_4830,In_3243,In_1378);
nor U4831 (N_4831,In_234,In_4571);
nor U4832 (N_4832,In_3424,In_3685);
xnor U4833 (N_4833,In_187,In_1794);
or U4834 (N_4834,In_4983,In_1631);
nor U4835 (N_4835,In_4627,In_1466);
or U4836 (N_4836,In_3886,In_4476);
and U4837 (N_4837,In_4905,In_577);
nor U4838 (N_4838,In_3332,In_3066);
and U4839 (N_4839,In_4030,In_1334);
xnor U4840 (N_4840,In_4586,In_2162);
and U4841 (N_4841,In_1353,In_2006);
and U4842 (N_4842,In_4270,In_4257);
nor U4843 (N_4843,In_3319,In_2199);
nand U4844 (N_4844,In_1720,In_1488);
nand U4845 (N_4845,In_1560,In_2064);
or U4846 (N_4846,In_4131,In_4977);
nor U4847 (N_4847,In_3130,In_4963);
and U4848 (N_4848,In_736,In_3371);
nand U4849 (N_4849,In_1547,In_2740);
or U4850 (N_4850,In_419,In_3925);
and U4851 (N_4851,In_3569,In_4924);
xnor U4852 (N_4852,In_1359,In_3557);
and U4853 (N_4853,In_97,In_269);
or U4854 (N_4854,In_144,In_3411);
xnor U4855 (N_4855,In_4768,In_258);
xnor U4856 (N_4856,In_2826,In_1498);
and U4857 (N_4857,In_3343,In_1203);
and U4858 (N_4858,In_4473,In_2825);
nand U4859 (N_4859,In_2091,In_3510);
nor U4860 (N_4860,In_1407,In_2239);
nor U4861 (N_4861,In_1827,In_206);
nor U4862 (N_4862,In_2004,In_881);
nor U4863 (N_4863,In_4801,In_1302);
nand U4864 (N_4864,In_4315,In_4577);
nand U4865 (N_4865,In_1570,In_4426);
nand U4866 (N_4866,In_2241,In_3403);
nor U4867 (N_4867,In_1632,In_1079);
nor U4868 (N_4868,In_798,In_1024);
nor U4869 (N_4869,In_990,In_3387);
nor U4870 (N_4870,In_2089,In_4562);
or U4871 (N_4871,In_1172,In_4744);
nand U4872 (N_4872,In_2081,In_2557);
and U4873 (N_4873,In_3992,In_1554);
and U4874 (N_4874,In_1280,In_4238);
nor U4875 (N_4875,In_3585,In_2993);
nand U4876 (N_4876,In_1723,In_4895);
nor U4877 (N_4877,In_179,In_4923);
xor U4878 (N_4878,In_4360,In_1859);
nand U4879 (N_4879,In_4282,In_2254);
or U4880 (N_4880,In_3363,In_2423);
and U4881 (N_4881,In_596,In_1300);
and U4882 (N_4882,In_565,In_908);
nor U4883 (N_4883,In_4649,In_302);
nor U4884 (N_4884,In_1508,In_1854);
nor U4885 (N_4885,In_2179,In_2141);
and U4886 (N_4886,In_4494,In_3582);
nand U4887 (N_4887,In_1779,In_1690);
nand U4888 (N_4888,In_4066,In_1123);
nor U4889 (N_4889,In_441,In_982);
or U4890 (N_4890,In_3149,In_3162);
and U4891 (N_4891,In_1068,In_3723);
nand U4892 (N_4892,In_2463,In_3252);
nand U4893 (N_4893,In_1207,In_2831);
nand U4894 (N_4894,In_1239,In_3346);
or U4895 (N_4895,In_429,In_1323);
or U4896 (N_4896,In_4056,In_2218);
xnor U4897 (N_4897,In_983,In_1979);
nand U4898 (N_4898,In_1875,In_4271);
or U4899 (N_4899,In_3585,In_2454);
nand U4900 (N_4900,In_18,In_2900);
and U4901 (N_4901,In_3986,In_3576);
and U4902 (N_4902,In_2821,In_771);
nand U4903 (N_4903,In_3190,In_2726);
nor U4904 (N_4904,In_3116,In_1114);
nor U4905 (N_4905,In_636,In_162);
or U4906 (N_4906,In_3717,In_199);
nor U4907 (N_4907,In_4413,In_2602);
nor U4908 (N_4908,In_2115,In_2017);
nor U4909 (N_4909,In_2488,In_622);
or U4910 (N_4910,In_3534,In_4055);
xor U4911 (N_4911,In_599,In_267);
and U4912 (N_4912,In_1099,In_4522);
and U4913 (N_4913,In_2118,In_4242);
or U4914 (N_4914,In_3906,In_839);
nor U4915 (N_4915,In_482,In_3309);
xnor U4916 (N_4916,In_1603,In_2215);
and U4917 (N_4917,In_2655,In_3731);
or U4918 (N_4918,In_4038,In_1528);
nand U4919 (N_4919,In_1862,In_4003);
and U4920 (N_4920,In_881,In_3856);
xnor U4921 (N_4921,In_4976,In_2738);
and U4922 (N_4922,In_3747,In_338);
and U4923 (N_4923,In_2400,In_1507);
nand U4924 (N_4924,In_2528,In_4204);
nand U4925 (N_4925,In_1382,In_871);
and U4926 (N_4926,In_3573,In_4465);
nand U4927 (N_4927,In_1126,In_4688);
and U4928 (N_4928,In_4587,In_3453);
or U4929 (N_4929,In_2542,In_4798);
nor U4930 (N_4930,In_4967,In_2432);
nand U4931 (N_4931,In_30,In_2623);
or U4932 (N_4932,In_475,In_4935);
and U4933 (N_4933,In_536,In_1618);
nor U4934 (N_4934,In_207,In_2893);
nand U4935 (N_4935,In_4870,In_1446);
nor U4936 (N_4936,In_4752,In_162);
nor U4937 (N_4937,In_1774,In_3972);
and U4938 (N_4938,In_3052,In_1134);
nand U4939 (N_4939,In_3472,In_4691);
nand U4940 (N_4940,In_4342,In_594);
or U4941 (N_4941,In_3500,In_4834);
nand U4942 (N_4942,In_3598,In_2626);
and U4943 (N_4943,In_2856,In_2484);
nor U4944 (N_4944,In_3554,In_3572);
or U4945 (N_4945,In_751,In_350);
xnor U4946 (N_4946,In_717,In_2142);
nand U4947 (N_4947,In_437,In_4523);
nor U4948 (N_4948,In_3710,In_2452);
nor U4949 (N_4949,In_3363,In_2515);
and U4950 (N_4950,In_2977,In_4813);
nand U4951 (N_4951,In_4920,In_1491);
or U4952 (N_4952,In_2045,In_4984);
nand U4953 (N_4953,In_1130,In_4242);
and U4954 (N_4954,In_3829,In_541);
xor U4955 (N_4955,In_4698,In_3020);
or U4956 (N_4956,In_2531,In_271);
xnor U4957 (N_4957,In_2707,In_2143);
nand U4958 (N_4958,In_2714,In_4860);
nor U4959 (N_4959,In_1208,In_1355);
or U4960 (N_4960,In_4386,In_3384);
and U4961 (N_4961,In_1017,In_3569);
nor U4962 (N_4962,In_321,In_2663);
nor U4963 (N_4963,In_3724,In_2934);
and U4964 (N_4964,In_1683,In_4001);
and U4965 (N_4965,In_1940,In_516);
and U4966 (N_4966,In_3020,In_1465);
and U4967 (N_4967,In_563,In_3313);
nor U4968 (N_4968,In_636,In_1884);
and U4969 (N_4969,In_3248,In_1512);
nand U4970 (N_4970,In_3123,In_1927);
nor U4971 (N_4971,In_1519,In_3242);
and U4972 (N_4972,In_1367,In_3293);
xor U4973 (N_4973,In_500,In_57);
nor U4974 (N_4974,In_2013,In_4209);
nor U4975 (N_4975,In_3602,In_4186);
or U4976 (N_4976,In_402,In_2487);
and U4977 (N_4977,In_4302,In_4143);
xor U4978 (N_4978,In_1511,In_367);
nor U4979 (N_4979,In_4954,In_1819);
nand U4980 (N_4980,In_3332,In_1984);
nor U4981 (N_4981,In_924,In_1749);
or U4982 (N_4982,In_2553,In_2209);
or U4983 (N_4983,In_955,In_4045);
nor U4984 (N_4984,In_363,In_434);
xnor U4985 (N_4985,In_2950,In_3460);
nor U4986 (N_4986,In_1089,In_3985);
and U4987 (N_4987,In_3438,In_2014);
and U4988 (N_4988,In_1287,In_3523);
and U4989 (N_4989,In_983,In_3979);
nand U4990 (N_4990,In_2176,In_4842);
or U4991 (N_4991,In_3309,In_946);
xor U4992 (N_4992,In_3046,In_3387);
nand U4993 (N_4993,In_3877,In_2470);
or U4994 (N_4994,In_1846,In_3548);
xor U4995 (N_4995,In_1448,In_1318);
and U4996 (N_4996,In_4655,In_2885);
xor U4997 (N_4997,In_1022,In_3578);
nor U4998 (N_4998,In_3268,In_1591);
or U4999 (N_4999,In_3160,In_1118);
or U5000 (N_5000,N_3728,N_2337);
and U5001 (N_5001,N_1368,N_3681);
and U5002 (N_5002,N_2201,N_1306);
and U5003 (N_5003,N_1071,N_1597);
nor U5004 (N_5004,N_4247,N_4980);
nand U5005 (N_5005,N_4619,N_3158);
or U5006 (N_5006,N_4204,N_3748);
and U5007 (N_5007,N_2407,N_3279);
and U5008 (N_5008,N_232,N_733);
or U5009 (N_5009,N_1120,N_4943);
or U5010 (N_5010,N_4040,N_3490);
nor U5011 (N_5011,N_2100,N_1802);
or U5012 (N_5012,N_2919,N_4085);
nor U5013 (N_5013,N_1105,N_1462);
or U5014 (N_5014,N_4344,N_502);
nor U5015 (N_5015,N_507,N_3166);
nand U5016 (N_5016,N_4759,N_2090);
nor U5017 (N_5017,N_473,N_214);
nand U5018 (N_5018,N_3356,N_1782);
and U5019 (N_5019,N_4604,N_1174);
xor U5020 (N_5020,N_4087,N_155);
nand U5021 (N_5021,N_1749,N_4186);
or U5022 (N_5022,N_674,N_3810);
and U5023 (N_5023,N_356,N_2755);
nor U5024 (N_5024,N_1121,N_4148);
nand U5025 (N_5025,N_625,N_3315);
xor U5026 (N_5026,N_3746,N_2845);
nand U5027 (N_5027,N_1407,N_1626);
xor U5028 (N_5028,N_1976,N_1442);
and U5029 (N_5029,N_2224,N_1046);
nor U5030 (N_5030,N_4799,N_2151);
nor U5031 (N_5031,N_1585,N_3779);
or U5032 (N_5032,N_4476,N_3030);
nor U5033 (N_5033,N_2029,N_1864);
nor U5034 (N_5034,N_2254,N_3107);
and U5035 (N_5035,N_4329,N_663);
xor U5036 (N_5036,N_4218,N_220);
nand U5037 (N_5037,N_1773,N_408);
xor U5038 (N_5038,N_3185,N_1033);
nand U5039 (N_5039,N_1087,N_3502);
nand U5040 (N_5040,N_654,N_3176);
and U5041 (N_5041,N_3248,N_998);
and U5042 (N_5042,N_2959,N_3685);
nor U5043 (N_5043,N_49,N_3578);
and U5044 (N_5044,N_4195,N_441);
xnor U5045 (N_5045,N_3684,N_542);
and U5046 (N_5046,N_2047,N_4539);
nand U5047 (N_5047,N_1834,N_2112);
nand U5048 (N_5048,N_3295,N_854);
and U5049 (N_5049,N_2764,N_4669);
nand U5050 (N_5050,N_1238,N_2610);
and U5051 (N_5051,N_2804,N_3117);
nand U5052 (N_5052,N_3686,N_3220);
or U5053 (N_5053,N_1662,N_1086);
or U5054 (N_5054,N_3568,N_3260);
nand U5055 (N_5055,N_397,N_1390);
and U5056 (N_5056,N_178,N_1798);
nand U5057 (N_5057,N_2376,N_3812);
nand U5058 (N_5058,N_223,N_2825);
or U5059 (N_5059,N_4910,N_544);
nand U5060 (N_5060,N_185,N_70);
and U5061 (N_5061,N_14,N_712);
or U5062 (N_5062,N_284,N_3980);
or U5063 (N_5063,N_688,N_4632);
or U5064 (N_5064,N_2396,N_817);
nand U5065 (N_5065,N_4133,N_2244);
nor U5066 (N_5066,N_3857,N_944);
and U5067 (N_5067,N_1661,N_1269);
nor U5068 (N_5068,N_254,N_2917);
or U5069 (N_5069,N_1088,N_60);
or U5070 (N_5070,N_3640,N_593);
or U5071 (N_5071,N_1399,N_3817);
and U5072 (N_5072,N_2937,N_1289);
nand U5073 (N_5073,N_3861,N_692);
or U5074 (N_5074,N_353,N_4831);
nand U5075 (N_5075,N_3522,N_1586);
nand U5076 (N_5076,N_4340,N_2135);
nand U5077 (N_5077,N_1781,N_2991);
and U5078 (N_5078,N_120,N_48);
nor U5079 (N_5079,N_4656,N_1673);
and U5080 (N_5080,N_4364,N_697);
nor U5081 (N_5081,N_447,N_3552);
or U5082 (N_5082,N_323,N_2631);
nand U5083 (N_5083,N_624,N_404);
or U5084 (N_5084,N_335,N_1867);
and U5085 (N_5085,N_1800,N_4228);
nand U5086 (N_5086,N_3702,N_1872);
nand U5087 (N_5087,N_3055,N_4473);
or U5088 (N_5088,N_971,N_4482);
and U5089 (N_5089,N_3112,N_4991);
or U5090 (N_5090,N_4298,N_3473);
xor U5091 (N_5091,N_4007,N_311);
nand U5092 (N_5092,N_2734,N_2036);
nand U5093 (N_5093,N_84,N_3078);
nand U5094 (N_5094,N_0,N_445);
nand U5095 (N_5095,N_583,N_2938);
nand U5096 (N_5096,N_3643,N_2699);
nand U5097 (N_5097,N_4966,N_1728);
nand U5098 (N_5098,N_551,N_18);
nor U5099 (N_5099,N_3447,N_3351);
nand U5100 (N_5100,N_4797,N_175);
nor U5101 (N_5101,N_1763,N_3137);
nand U5102 (N_5102,N_2505,N_3092);
or U5103 (N_5103,N_1665,N_3280);
xnor U5104 (N_5104,N_1326,N_4025);
or U5105 (N_5105,N_30,N_4917);
xnor U5106 (N_5106,N_2843,N_483);
nor U5107 (N_5107,N_1899,N_2163);
xnor U5108 (N_5108,N_302,N_2323);
and U5109 (N_5109,N_3270,N_1868);
nand U5110 (N_5110,N_55,N_3815);
or U5111 (N_5111,N_3478,N_2452);
xnor U5112 (N_5112,N_1658,N_1895);
nand U5113 (N_5113,N_2821,N_1829);
nand U5114 (N_5114,N_3754,N_1278);
or U5115 (N_5115,N_2936,N_4225);
and U5116 (N_5116,N_993,N_2609);
nor U5117 (N_5117,N_3836,N_3085);
nor U5118 (N_5118,N_2878,N_1841);
and U5119 (N_5119,N_3916,N_2183);
nand U5120 (N_5120,N_2598,N_3088);
nand U5121 (N_5121,N_1455,N_2908);
or U5122 (N_5122,N_3506,N_217);
or U5123 (N_5123,N_849,N_4230);
nand U5124 (N_5124,N_3480,N_1352);
xnor U5125 (N_5125,N_1489,N_2714);
or U5126 (N_5126,N_3093,N_672);
nand U5127 (N_5127,N_2654,N_2616);
nand U5128 (N_5128,N_2028,N_2421);
or U5129 (N_5129,N_2620,N_1051);
xor U5130 (N_5130,N_4872,N_609);
nand U5131 (N_5131,N_3307,N_4697);
nand U5132 (N_5132,N_1161,N_3637);
and U5133 (N_5133,N_2692,N_4821);
and U5134 (N_5134,N_1785,N_4594);
nand U5135 (N_5135,N_2241,N_4321);
nor U5136 (N_5136,N_3436,N_4946);
nand U5137 (N_5137,N_3846,N_29);
nor U5138 (N_5138,N_3658,N_4440);
or U5139 (N_5139,N_2984,N_3694);
nand U5140 (N_5140,N_4090,N_2374);
nand U5141 (N_5141,N_3387,N_4947);
and U5142 (N_5142,N_3050,N_2292);
nor U5143 (N_5143,N_201,N_3274);
or U5144 (N_5144,N_3291,N_3720);
nor U5145 (N_5145,N_2463,N_1073);
nand U5146 (N_5146,N_652,N_3284);
nand U5147 (N_5147,N_482,N_2689);
nand U5148 (N_5148,N_4516,N_2345);
nor U5149 (N_5149,N_3974,N_3268);
or U5150 (N_5150,N_1023,N_437);
and U5151 (N_5151,N_3427,N_1055);
xnor U5152 (N_5152,N_2205,N_4388);
nor U5153 (N_5153,N_600,N_2538);
and U5154 (N_5154,N_3074,N_16);
or U5155 (N_5155,N_2302,N_384);
and U5156 (N_5156,N_4505,N_386);
nor U5157 (N_5157,N_4242,N_3213);
and U5158 (N_5158,N_4731,N_3363);
nor U5159 (N_5159,N_1267,N_802);
xnor U5160 (N_5160,N_841,N_2999);
nor U5161 (N_5161,N_199,N_1446);
or U5162 (N_5162,N_1173,N_1754);
and U5163 (N_5163,N_4960,N_373);
nor U5164 (N_5164,N_2669,N_4652);
or U5165 (N_5165,N_4015,N_578);
nor U5166 (N_5166,N_2942,N_4716);
and U5167 (N_5167,N_1726,N_216);
nand U5168 (N_5168,N_166,N_4989);
or U5169 (N_5169,N_4955,N_4844);
or U5170 (N_5170,N_3992,N_91);
xnor U5171 (N_5171,N_4355,N_2574);
nand U5172 (N_5172,N_1149,N_582);
and U5173 (N_5173,N_2909,N_2852);
nor U5174 (N_5174,N_1048,N_4832);
nor U5175 (N_5175,N_533,N_3269);
nand U5176 (N_5176,N_2078,N_1984);
xnor U5177 (N_5177,N_2829,N_1905);
nand U5178 (N_5178,N_684,N_1224);
nor U5179 (N_5179,N_3532,N_446);
nor U5180 (N_5180,N_129,N_3513);
nand U5181 (N_5181,N_1472,N_4368);
nand U5182 (N_5182,N_1250,N_4415);
nand U5183 (N_5183,N_4501,N_2572);
nand U5184 (N_5184,N_3003,N_200);
nand U5185 (N_5185,N_4800,N_4219);
and U5186 (N_5186,N_823,N_2473);
nor U5187 (N_5187,N_1599,N_2954);
nor U5188 (N_5188,N_2270,N_4626);
and U5189 (N_5189,N_4926,N_3249);
xnor U5190 (N_5190,N_3182,N_862);
and U5191 (N_5191,N_4478,N_4411);
nand U5192 (N_5192,N_847,N_4264);
or U5193 (N_5193,N_3168,N_2043);
nor U5194 (N_5194,N_1060,N_2976);
nor U5195 (N_5195,N_3312,N_2710);
and U5196 (N_5196,N_3322,N_211);
nand U5197 (N_5197,N_3128,N_3125);
and U5198 (N_5198,N_2877,N_1491);
or U5199 (N_5199,N_248,N_2310);
and U5200 (N_5200,N_837,N_4235);
nand U5201 (N_5201,N_3521,N_2943);
and U5202 (N_5202,N_4681,N_1603);
and U5203 (N_5203,N_747,N_745);
and U5204 (N_5204,N_2176,N_4013);
and U5205 (N_5205,N_4083,N_3808);
nand U5206 (N_5206,N_4940,N_4142);
or U5207 (N_5207,N_576,N_4098);
xnor U5208 (N_5208,N_3965,N_1593);
or U5209 (N_5209,N_3350,N_3147);
and U5210 (N_5210,N_1194,N_3624);
xor U5211 (N_5211,N_1427,N_2202);
or U5212 (N_5212,N_283,N_2569);
nand U5213 (N_5213,N_2182,N_171);
and U5214 (N_5214,N_3566,N_3780);
xnor U5215 (N_5215,N_4746,N_340);
nand U5216 (N_5216,N_1428,N_846);
xor U5217 (N_5217,N_3082,N_4023);
nand U5218 (N_5218,N_259,N_2913);
or U5219 (N_5219,N_215,N_169);
nand U5220 (N_5220,N_4131,N_1254);
or U5221 (N_5221,N_1300,N_4965);
nor U5222 (N_5222,N_784,N_4734);
or U5223 (N_5223,N_1237,N_2060);
nand U5224 (N_5224,N_4804,N_4959);
nand U5225 (N_5225,N_3736,N_411);
or U5226 (N_5226,N_2304,N_2601);
and U5227 (N_5227,N_4294,N_931);
or U5228 (N_5228,N_1878,N_3947);
nor U5229 (N_5229,N_3641,N_308);
nand U5230 (N_5230,N_93,N_351);
or U5231 (N_5231,N_126,N_260);
nand U5232 (N_5232,N_4564,N_2299);
or U5233 (N_5233,N_1050,N_4082);
and U5234 (N_5234,N_4081,N_2419);
and U5235 (N_5235,N_3587,N_1476);
and U5236 (N_5236,N_1038,N_851);
or U5237 (N_5237,N_980,N_1053);
nand U5238 (N_5238,N_1447,N_2);
and U5239 (N_5239,N_3868,N_3978);
xor U5240 (N_5240,N_1002,N_1772);
or U5241 (N_5241,N_2216,N_152);
nand U5242 (N_5242,N_127,N_755);
nand U5243 (N_5243,N_4441,N_3120);
nand U5244 (N_5244,N_4413,N_33);
nand U5245 (N_5245,N_1738,N_4975);
and U5246 (N_5246,N_3494,N_3793);
and U5247 (N_5247,N_4471,N_2320);
or U5248 (N_5248,N_330,N_1978);
or U5249 (N_5249,N_4328,N_41);
nand U5250 (N_5250,N_858,N_3921);
or U5251 (N_5251,N_4969,N_218);
nand U5252 (N_5252,N_184,N_1153);
nand U5253 (N_5253,N_2827,N_2520);
or U5254 (N_5254,N_1499,N_1605);
and U5255 (N_5255,N_3994,N_2778);
nor U5256 (N_5256,N_2603,N_191);
and U5257 (N_5257,N_4707,N_342);
or U5258 (N_5258,N_4560,N_23);
or U5259 (N_5259,N_2243,N_396);
nand U5260 (N_5260,N_979,N_2793);
xor U5261 (N_5261,N_4189,N_1840);
xnor U5262 (N_5262,N_2548,N_4168);
or U5263 (N_5263,N_1724,N_1793);
nand U5264 (N_5264,N_1759,N_3452);
nor U5265 (N_5265,N_1275,N_3306);
nor U5266 (N_5266,N_1980,N_1618);
or U5267 (N_5267,N_2405,N_476);
nor U5268 (N_5268,N_2398,N_4951);
nor U5269 (N_5269,N_2651,N_1588);
or U5270 (N_5270,N_2808,N_1027);
nor U5271 (N_5271,N_3445,N_607);
nor U5272 (N_5272,N_2422,N_3930);
nand U5273 (N_5273,N_1104,N_454);
nor U5274 (N_5274,N_1495,N_2153);
or U5275 (N_5275,N_4693,N_1089);
and U5276 (N_5276,N_1676,N_4155);
and U5277 (N_5277,N_256,N_246);
nand U5278 (N_5278,N_4270,N_4791);
or U5279 (N_5279,N_3934,N_3617);
and U5280 (N_5280,N_264,N_4593);
nor U5281 (N_5281,N_4396,N_1939);
or U5282 (N_5282,N_795,N_367);
or U5283 (N_5283,N_810,N_160);
and U5284 (N_5284,N_503,N_575);
and U5285 (N_5285,N_4753,N_4934);
nand U5286 (N_5286,N_1682,N_1388);
or U5287 (N_5287,N_3028,N_4992);
nand U5288 (N_5288,N_4984,N_3497);
nor U5289 (N_5289,N_2291,N_4634);
nor U5290 (N_5290,N_51,N_560);
or U5291 (N_5291,N_3734,N_1412);
xor U5292 (N_5292,N_1896,N_3191);
and U5293 (N_5293,N_911,N_3842);
and U5294 (N_5294,N_3275,N_2789);
nand U5295 (N_5295,N_4589,N_4521);
nand U5296 (N_5296,N_2772,N_2638);
or U5297 (N_5297,N_3990,N_1144);
nand U5298 (N_5298,N_2663,N_388);
and U5299 (N_5299,N_227,N_1312);
nand U5300 (N_5300,N_3535,N_2040);
xor U5301 (N_5301,N_4572,N_2246);
and U5302 (N_5302,N_2066,N_2494);
nor U5303 (N_5303,N_2230,N_3998);
and U5304 (N_5304,N_3262,N_4367);
nor U5305 (N_5305,N_4404,N_2719);
nand U5306 (N_5306,N_3847,N_3241);
nand U5307 (N_5307,N_638,N_4034);
or U5308 (N_5308,N_2104,N_2171);
or U5309 (N_5309,N_3599,N_1703);
or U5310 (N_5310,N_1551,N_4937);
and U5311 (N_5311,N_213,N_3118);
nand U5312 (N_5312,N_4853,N_3848);
nand U5313 (N_5313,N_963,N_2904);
nand U5314 (N_5314,N_2615,N_2342);
nor U5315 (N_5315,N_2058,N_2543);
or U5316 (N_5316,N_1006,N_763);
and U5317 (N_5317,N_2306,N_3380);
or U5318 (N_5318,N_2626,N_1389);
nor U5319 (N_5319,N_4875,N_3486);
nand U5320 (N_5320,N_4672,N_929);
nand U5321 (N_5321,N_4324,N_973);
or U5322 (N_5322,N_2140,N_4256);
nand U5323 (N_5323,N_4153,N_3798);
and U5324 (N_5324,N_4874,N_2830);
or U5325 (N_5325,N_1404,N_2437);
or U5326 (N_5326,N_4483,N_4719);
nand U5327 (N_5327,N_1413,N_1965);
xor U5328 (N_5328,N_2354,N_130);
xor U5329 (N_5329,N_3931,N_3049);
and U5330 (N_5330,N_3972,N_2023);
and U5331 (N_5331,N_2257,N_1775);
or U5332 (N_5332,N_193,N_2633);
nand U5333 (N_5333,N_848,N_2081);
and U5334 (N_5334,N_875,N_2567);
nand U5335 (N_5335,N_1647,N_4703);
nor U5336 (N_5336,N_631,N_4453);
or U5337 (N_5337,N_2048,N_3923);
or U5338 (N_5338,N_904,N_4858);
nor U5339 (N_5339,N_298,N_183);
nor U5340 (N_5340,N_3619,N_2747);
nor U5341 (N_5341,N_4795,N_2436);
nand U5342 (N_5342,N_2737,N_2123);
nand U5343 (N_5343,N_4156,N_4467);
nand U5344 (N_5344,N_872,N_2497);
or U5345 (N_5345,N_3973,N_890);
or U5346 (N_5346,N_4709,N_1216);
xnor U5347 (N_5347,N_2953,N_3109);
and U5348 (N_5348,N_2739,N_901);
nor U5349 (N_5349,N_414,N_4750);
or U5350 (N_5350,N_737,N_210);
xor U5351 (N_5351,N_1982,N_3504);
or U5352 (N_5352,N_2196,N_4512);
or U5353 (N_5353,N_1203,N_4559);
nor U5354 (N_5354,N_2550,N_4954);
or U5355 (N_5355,N_759,N_2486);
or U5356 (N_5356,N_3906,N_3545);
and U5357 (N_5357,N_333,N_1745);
or U5358 (N_5358,N_1420,N_4140);
nor U5359 (N_5359,N_3007,N_4163);
nand U5360 (N_5360,N_4193,N_1953);
xor U5361 (N_5361,N_1094,N_1415);
and U5362 (N_5362,N_3046,N_1525);
and U5363 (N_5363,N_2898,N_3762);
and U5364 (N_5364,N_1102,N_641);
and U5365 (N_5365,N_2261,N_2540);
and U5366 (N_5366,N_3946,N_3154);
xnor U5367 (N_5367,N_3361,N_4525);
or U5368 (N_5368,N_4124,N_3448);
or U5369 (N_5369,N_3354,N_2442);
or U5370 (N_5370,N_4215,N_1125);
or U5371 (N_5371,N_4145,N_3570);
nor U5372 (N_5372,N_4456,N_2557);
nand U5373 (N_5373,N_3011,N_4576);
xor U5374 (N_5374,N_965,N_1609);
and U5375 (N_5375,N_681,N_1947);
and U5376 (N_5376,N_2792,N_1241);
xor U5377 (N_5377,N_1701,N_1493);
and U5378 (N_5378,N_668,N_250);
nand U5379 (N_5379,N_2316,N_2471);
nand U5380 (N_5380,N_2105,N_4177);
xor U5381 (N_5381,N_73,N_1496);
nand U5382 (N_5382,N_3381,N_4768);
and U5383 (N_5383,N_2381,N_2348);
nor U5384 (N_5384,N_2911,N_1253);
and U5385 (N_5385,N_3647,N_1721);
nand U5386 (N_5386,N_3612,N_3703);
or U5387 (N_5387,N_3613,N_1202);
or U5388 (N_5388,N_1284,N_635);
and U5389 (N_5389,N_1353,N_2264);
nand U5390 (N_5390,N_1314,N_4331);
or U5391 (N_5391,N_1434,N_518);
nand U5392 (N_5392,N_1068,N_3027);
and U5393 (N_5393,N_2659,N_3369);
nor U5394 (N_5394,N_4585,N_2915);
or U5395 (N_5395,N_2800,N_3051);
and U5396 (N_5396,N_1334,N_1906);
nor U5397 (N_5397,N_2847,N_1200);
nor U5398 (N_5398,N_2069,N_3124);
nor U5399 (N_5399,N_4674,N_1336);
or U5400 (N_5400,N_4210,N_1308);
and U5401 (N_5401,N_2042,N_657);
xor U5402 (N_5402,N_190,N_3608);
nor U5403 (N_5403,N_4487,N_866);
nor U5404 (N_5404,N_2880,N_4458);
or U5405 (N_5405,N_2231,N_1850);
and U5406 (N_5406,N_1667,N_1030);
and U5407 (N_5407,N_1163,N_2359);
nand U5408 (N_5408,N_3273,N_1329);
or U5409 (N_5409,N_1645,N_4182);
nor U5410 (N_5410,N_4406,N_2883);
nor U5411 (N_5411,N_4738,N_822);
and U5412 (N_5412,N_1123,N_1681);
or U5413 (N_5413,N_3707,N_4679);
and U5414 (N_5414,N_1715,N_1718);
nor U5415 (N_5415,N_2454,N_573);
xnor U5416 (N_5416,N_3598,N_4659);
nor U5417 (N_5417,N_4949,N_2109);
or U5418 (N_5418,N_2448,N_3485);
nand U5419 (N_5419,N_209,N_234);
xor U5420 (N_5420,N_2738,N_597);
nor U5421 (N_5421,N_2655,N_2079);
nor U5422 (N_5422,N_1522,N_2971);
xor U5423 (N_5423,N_141,N_3329);
or U5424 (N_5424,N_3537,N_4561);
or U5425 (N_5425,N_1583,N_3180);
nand U5426 (N_5426,N_3403,N_2614);
or U5427 (N_5427,N_1674,N_3477);
nand U5428 (N_5428,N_273,N_4260);
nor U5429 (N_5429,N_2696,N_3559);
nand U5430 (N_5430,N_1537,N_1350);
and U5431 (N_5431,N_147,N_4472);
and U5432 (N_5432,N_2977,N_4028);
xnor U5433 (N_5433,N_4115,N_4689);
nand U5434 (N_5434,N_1709,N_1204);
or U5435 (N_5435,N_4039,N_2677);
and U5436 (N_5436,N_3620,N_2077);
nor U5437 (N_5437,N_3706,N_24);
xor U5438 (N_5438,N_1543,N_774);
nor U5439 (N_5439,N_693,N_2427);
or U5440 (N_5440,N_1988,N_2203);
xor U5441 (N_5441,N_3903,N_964);
or U5442 (N_5442,N_4764,N_434);
nor U5443 (N_5443,N_2590,N_4664);
nor U5444 (N_5444,N_2673,N_2210);
or U5445 (N_5445,N_1807,N_2576);
nor U5446 (N_5446,N_3839,N_2145);
and U5447 (N_5447,N_188,N_344);
nand U5448 (N_5448,N_4392,N_1400);
and U5449 (N_5449,N_164,N_3272);
and U5450 (N_5450,N_196,N_722);
nor U5451 (N_5451,N_740,N_664);
nand U5452 (N_5452,N_241,N_1544);
xor U5453 (N_5453,N_3276,N_497);
nand U5454 (N_5454,N_38,N_2357);
or U5455 (N_5455,N_3386,N_2884);
nor U5456 (N_5456,N_3009,N_3717);
and U5457 (N_5457,N_288,N_878);
nor U5458 (N_5458,N_2392,N_559);
or U5459 (N_5459,N_3483,N_380);
and U5460 (N_5460,N_1419,N_2760);
nand U5461 (N_5461,N_4971,N_883);
xnor U5462 (N_5462,N_3753,N_2885);
and U5463 (N_5463,N_3806,N_124);
and U5464 (N_5464,N_3061,N_907);
or U5465 (N_5465,N_3621,N_4915);
and U5466 (N_5466,N_63,N_2649);
nor U5467 (N_5467,N_4578,N_4702);
nor U5468 (N_5468,N_28,N_4866);
and U5469 (N_5469,N_4773,N_4938);
nand U5470 (N_5470,N_3553,N_3708);
and U5471 (N_5471,N_1456,N_423);
nand U5472 (N_5472,N_2750,N_2950);
and U5473 (N_5473,N_3173,N_966);
xor U5474 (N_5474,N_1938,N_2508);
nor U5475 (N_5475,N_1600,N_3277);
or U5476 (N_5476,N_4810,N_1025);
and U5477 (N_5477,N_4823,N_4301);
nor U5478 (N_5478,N_2403,N_324);
nand U5479 (N_5479,N_4706,N_3374);
or U5480 (N_5480,N_4922,N_4784);
and U5481 (N_5481,N_1066,N_653);
nor U5482 (N_5482,N_1578,N_3100);
or U5483 (N_5483,N_1986,N_403);
or U5484 (N_5484,N_1915,N_2004);
nand U5485 (N_5485,N_422,N_3103);
and U5486 (N_5486,N_4387,N_2679);
nand U5487 (N_5487,N_1058,N_4653);
and U5488 (N_5488,N_144,N_546);
nor U5489 (N_5489,N_1171,N_3496);
nand U5490 (N_5490,N_3881,N_3984);
nand U5491 (N_5491,N_1340,N_1505);
nand U5492 (N_5492,N_244,N_1504);
or U5493 (N_5493,N_4451,N_4936);
and U5494 (N_5494,N_3075,N_4714);
or U5495 (N_5495,N_4586,N_2816);
xnor U5496 (N_5496,N_4121,N_2050);
nor U5497 (N_5497,N_3971,N_2686);
or U5498 (N_5498,N_2277,N_3673);
nand U5499 (N_5499,N_4597,N_4283);
or U5500 (N_5500,N_253,N_3775);
and U5501 (N_5501,N_2161,N_1826);
nor U5502 (N_5502,N_3081,N_440);
nand U5503 (N_5503,N_1127,N_3834);
and U5504 (N_5504,N_3663,N_2511);
nand U5505 (N_5505,N_4893,N_154);
or U5506 (N_5506,N_2838,N_3188);
nand U5507 (N_5507,N_159,N_4060);
or U5508 (N_5508,N_3451,N_4447);
nor U5509 (N_5509,N_721,N_2120);
and U5510 (N_5510,N_1235,N_831);
nand U5511 (N_5511,N_1507,N_212);
and U5512 (N_5512,N_1614,N_1677);
nor U5513 (N_5513,N_3246,N_1266);
nor U5514 (N_5514,N_2371,N_2003);
nor U5515 (N_5515,N_3651,N_1766);
nand U5516 (N_5516,N_4904,N_1625);
nand U5517 (N_5517,N_1783,N_3087);
xor U5518 (N_5518,N_1044,N_3951);
nand U5519 (N_5519,N_3750,N_1780);
xnor U5520 (N_5520,N_2790,N_3243);
nand U5521 (N_5521,N_4906,N_4263);
xor U5522 (N_5522,N_4818,N_3035);
nand U5523 (N_5523,N_1069,N_2276);
and U5524 (N_5524,N_4515,N_2629);
nand U5525 (N_5525,N_1748,N_2093);
nand U5526 (N_5526,N_3033,N_3152);
or U5527 (N_5527,N_1262,N_1441);
or U5528 (N_5528,N_1574,N_4918);
nor U5529 (N_5529,N_3628,N_4780);
nor U5530 (N_5530,N_4921,N_2758);
nor U5531 (N_5531,N_4920,N_3474);
or U5532 (N_5532,N_4164,N_4316);
and U5533 (N_5533,N_1811,N_1771);
or U5534 (N_5534,N_1932,N_1955);
nor U5535 (N_5535,N_1650,N_2844);
and U5536 (N_5536,N_715,N_1619);
xnor U5537 (N_5537,N_1887,N_3763);
xnor U5538 (N_5538,N_305,N_3597);
or U5539 (N_5539,N_163,N_612);
and U5540 (N_5540,N_3872,N_716);
xnor U5541 (N_5541,N_4851,N_413);
nor U5542 (N_5542,N_3743,N_4615);
and U5543 (N_5543,N_1711,N_394);
or U5544 (N_5544,N_969,N_2702);
or U5545 (N_5545,N_1467,N_432);
nand U5546 (N_5546,N_3674,N_1032);
xnor U5547 (N_5547,N_3852,N_1083);
nor U5548 (N_5548,N_678,N_2149);
xnor U5549 (N_5549,N_4907,N_494);
and U5550 (N_5550,N_842,N_2867);
nor U5551 (N_5551,N_4407,N_1663);
and U5552 (N_5552,N_1358,N_4510);
nor U5553 (N_5553,N_2068,N_608);
and U5554 (N_5554,N_1426,N_87);
nor U5555 (N_5555,N_3534,N_839);
nand U5556 (N_5556,N_4217,N_2637);
nand U5557 (N_5557,N_4437,N_97);
nor U5558 (N_5558,N_3023,N_4254);
or U5559 (N_5559,N_669,N_433);
or U5560 (N_5560,N_492,N_1917);
nand U5561 (N_5561,N_1236,N_4027);
nand U5562 (N_5562,N_4555,N_4911);
or U5563 (N_5563,N_4913,N_1192);
and U5564 (N_5564,N_4044,N_1519);
nor U5565 (N_5565,N_1375,N_3211);
nand U5566 (N_5566,N_1477,N_3993);
and U5567 (N_5567,N_4391,N_530);
nor U5568 (N_5568,N_2114,N_2228);
or U5569 (N_5569,N_2142,N_2715);
nand U5570 (N_5570,N_3096,N_1580);
and U5571 (N_5571,N_2672,N_903);
and U5572 (N_5572,N_2340,N_2771);
nand U5573 (N_5573,N_2317,N_917);
nand U5574 (N_5574,N_1344,N_3760);
nor U5575 (N_5575,N_3463,N_2478);
and U5576 (N_5576,N_2418,N_3136);
nor U5577 (N_5577,N_1996,N_2981);
nand U5578 (N_5578,N_1839,N_505);
and U5579 (N_5579,N_2940,N_2147);
and U5580 (N_5580,N_2155,N_4053);
and U5581 (N_5581,N_3943,N_331);
nor U5582 (N_5582,N_956,N_202);
and U5583 (N_5583,N_2424,N_359);
nor U5584 (N_5584,N_343,N_3070);
and U5585 (N_5585,N_4794,N_3044);
nor U5586 (N_5586,N_3484,N_4397);
nand U5587 (N_5587,N_3,N_2818);
nor U5588 (N_5588,N_1922,N_1299);
nor U5589 (N_5589,N_1734,N_4012);
nor U5590 (N_5590,N_4883,N_2385);
nand U5591 (N_5591,N_4502,N_327);
nand U5592 (N_5592,N_622,N_3704);
and U5593 (N_5593,N_1874,N_893);
nand U5594 (N_5594,N_54,N_3263);
or U5595 (N_5595,N_1430,N_4064);
and U5596 (N_5596,N_772,N_293);
nor U5597 (N_5597,N_3461,N_2618);
nand U5598 (N_5598,N_1685,N_4336);
and U5599 (N_5599,N_119,N_4212);
nor U5600 (N_5600,N_2656,N_1175);
or U5601 (N_5601,N_2958,N_4405);
nor U5602 (N_5602,N_4745,N_2439);
xor U5603 (N_5603,N_750,N_222);
nor U5604 (N_5604,N_3744,N_125);
nand U5605 (N_5605,N_3721,N_536);
nor U5606 (N_5606,N_2347,N_2070);
and U5607 (N_5607,N_1659,N_2237);
or U5608 (N_5608,N_2960,N_4887);
and U5609 (N_5609,N_270,N_894);
and U5610 (N_5610,N_1601,N_1852);
or U5611 (N_5611,N_4019,N_4531);
or U5612 (N_5612,N_312,N_646);
or U5613 (N_5613,N_2275,N_31);
and U5614 (N_5614,N_105,N_192);
nor U5615 (N_5615,N_1858,N_729);
or U5616 (N_5616,N_2493,N_1554);
and U5617 (N_5617,N_718,N_701);
nor U5618 (N_5618,N_4996,N_928);
nand U5619 (N_5619,N_4688,N_145);
and U5620 (N_5620,N_3149,N_2853);
nand U5621 (N_5621,N_2639,N_393);
xnor U5622 (N_5622,N_1095,N_3340);
nand U5623 (N_5623,N_4805,N_2444);
nor U5624 (N_5624,N_601,N_3252);
nor U5625 (N_5625,N_3862,N_4342);
or U5626 (N_5626,N_3104,N_4704);
or U5627 (N_5627,N_938,N_3475);
and U5628 (N_5628,N_1264,N_2858);
xnor U5629 (N_5629,N_3823,N_3829);
and U5630 (N_5630,N_262,N_1570);
or U5631 (N_5631,N_974,N_2130);
and U5632 (N_5632,N_1684,N_4488);
and U5633 (N_5633,N_2326,N_3879);
and U5634 (N_5634,N_2429,N_4608);
nor U5635 (N_5635,N_1387,N_900);
nor U5636 (N_5636,N_4354,N_1613);
and U5637 (N_5637,N_591,N_379);
nand U5638 (N_5638,N_4848,N_3095);
and U5639 (N_5639,N_82,N_3813);
nand U5640 (N_5640,N_832,N_2343);
nor U5641 (N_5641,N_2281,N_26);
nand U5642 (N_5642,N_2537,N_4378);
and U5643 (N_5643,N_3310,N_3863);
or U5644 (N_5644,N_1337,N_4629);
nand U5645 (N_5645,N_3979,N_1680);
and U5646 (N_5646,N_2288,N_1746);
nor U5647 (N_5647,N_66,N_836);
or U5648 (N_5648,N_1582,N_2514);
and U5649 (N_5649,N_2732,N_923);
xor U5650 (N_5650,N_4639,N_4941);
nor U5651 (N_5651,N_1015,N_3129);
nand U5652 (N_5652,N_377,N_2555);
nand U5653 (N_5653,N_512,N_3800);
nand U5654 (N_5654,N_3809,N_2887);
or U5655 (N_5655,N_1750,N_1806);
and U5656 (N_5656,N_3919,N_1569);
nand U5657 (N_5657,N_1672,N_3870);
and U5658 (N_5658,N_3454,N_3510);
and U5659 (N_5659,N_811,N_4132);
nor U5660 (N_5660,N_3505,N_4777);
nand U5661 (N_5661,N_4180,N_3245);
nand U5662 (N_5662,N_4169,N_2839);
nor U5663 (N_5663,N_1933,N_3170);
nand U5664 (N_5664,N_813,N_1621);
nor U5665 (N_5665,N_4330,N_3232);
or U5666 (N_5666,N_2187,N_2854);
and U5667 (N_5667,N_540,N_2466);
and U5668 (N_5668,N_2881,N_1903);
and U5669 (N_5669,N_3938,N_1178);
nand U5670 (N_5670,N_2435,N_3339);
nand U5671 (N_5671,N_975,N_4766);
nand U5672 (N_5672,N_605,N_2495);
nor U5673 (N_5673,N_4741,N_2681);
nor U5674 (N_5674,N_2240,N_3582);
xor U5675 (N_5675,N_4248,N_1245);
or U5676 (N_5676,N_2634,N_1425);
nand U5677 (N_5677,N_950,N_1444);
or U5678 (N_5678,N_744,N_3867);
nand U5679 (N_5679,N_2623,N_531);
nor U5680 (N_5680,N_2513,N_3208);
nand U5681 (N_5681,N_3342,N_2477);
and U5682 (N_5682,N_888,N_4360);
and U5683 (N_5683,N_4520,N_3169);
or U5684 (N_5684,N_4809,N_586);
and U5685 (N_5685,N_4251,N_3589);
and U5686 (N_5686,N_1884,N_2064);
and U5687 (N_5687,N_271,N_2076);
nand U5688 (N_5688,N_2897,N_2685);
and U5689 (N_5689,N_3966,N_1879);
nor U5690 (N_5690,N_4696,N_2091);
nand U5691 (N_5691,N_577,N_2362);
and U5692 (N_5692,N_1758,N_4657);
and U5693 (N_5693,N_3233,N_4568);
nor U5694 (N_5694,N_4811,N_1769);
or U5695 (N_5695,N_2660,N_3557);
nor U5696 (N_5696,N_1008,N_1220);
and U5697 (N_5697,N_4430,N_140);
or U5698 (N_5698,N_4722,N_1311);
xnor U5699 (N_5699,N_2087,N_231);
xnor U5700 (N_5700,N_3196,N_2731);
xor U5701 (N_5701,N_3412,N_2535);
nor U5702 (N_5702,N_421,N_2946);
nand U5703 (N_5703,N_3654,N_3797);
nor U5704 (N_5704,N_4043,N_2172);
nand U5705 (N_5705,N_3230,N_3201);
nand U5706 (N_5706,N_1824,N_2242);
or U5707 (N_5707,N_2723,N_1248);
nand U5708 (N_5708,N_611,N_4231);
or U5709 (N_5709,N_4057,N_4481);
and U5710 (N_5710,N_2586,N_856);
xor U5711 (N_5711,N_4187,N_1942);
and U5712 (N_5712,N_2134,N_1473);
nor U5713 (N_5713,N_2249,N_3514);
nor U5714 (N_5714,N_2413,N_2923);
or U5715 (N_5715,N_1309,N_4756);
and U5716 (N_5716,N_2263,N_475);
and U5717 (N_5717,N_1657,N_4486);
nor U5718 (N_5718,N_3837,N_4508);
and U5719 (N_5719,N_2918,N_3791);
nand U5720 (N_5720,N_3038,N_3160);
nand U5721 (N_5721,N_1927,N_267);
nor U5722 (N_5722,N_17,N_4575);
and U5723 (N_5723,N_1360,N_2945);
or U5724 (N_5724,N_4573,N_1931);
or U5725 (N_5725,N_2975,N_4269);
xor U5726 (N_5726,N_3388,N_876);
nor U5727 (N_5727,N_3649,N_2177);
nor U5728 (N_5728,N_2284,N_402);
and U5729 (N_5729,N_1137,N_4438);
and U5730 (N_5730,N_4201,N_4785);
and U5731 (N_5731,N_4617,N_4878);
nand U5732 (N_5732,N_444,N_296);
nor U5733 (N_5733,N_3820,N_4737);
nor U5734 (N_5734,N_1641,N_4982);
and U5735 (N_5735,N_3080,N_350);
nor U5736 (N_5736,N_2185,N_3650);
nand U5737 (N_5737,N_3278,N_3110);
or U5738 (N_5738,N_3037,N_3214);
nand U5739 (N_5739,N_1722,N_2260);
nor U5740 (N_5740,N_2630,N_1112);
or U5741 (N_5741,N_1921,N_1832);
nor U5742 (N_5742,N_619,N_2571);
and U5743 (N_5743,N_4757,N_2107);
nand U5744 (N_5744,N_4903,N_3712);
nand U5745 (N_5745,N_520,N_886);
and U5746 (N_5746,N_3345,N_2215);
nand U5747 (N_5747,N_3739,N_4429);
xnor U5748 (N_5748,N_4055,N_661);
or U5749 (N_5749,N_4606,N_4588);
nand U5750 (N_5750,N_2562,N_855);
nor U5751 (N_5751,N_3722,N_3668);
or U5752 (N_5752,N_2222,N_3579);
nor U5753 (N_5753,N_1279,N_4782);
or U5754 (N_5754,N_3773,N_1821);
nand U5755 (N_5755,N_3313,N_1920);
nand U5756 (N_5756,N_3442,N_3290);
nand U5757 (N_5757,N_236,N_3792);
xor U5758 (N_5758,N_1335,N_2744);
nand U5759 (N_5759,N_960,N_528);
nor U5760 (N_5760,N_4258,N_783);
nor U5761 (N_5761,N_4891,N_2777);
nand U5762 (N_5762,N_4489,N_1549);
or U5763 (N_5763,N_3177,N_4705);
xnor U5764 (N_5764,N_834,N_2225);
nand U5765 (N_5765,N_1689,N_2994);
nor U5766 (N_5766,N_970,N_3265);
or U5767 (N_5767,N_2727,N_2443);
nand U5768 (N_5768,N_3255,N_4016);
and U5769 (N_5769,N_617,N_1369);
nand U5770 (N_5770,N_1348,N_3615);
or U5771 (N_5771,N_1151,N_1752);
and U5772 (N_5772,N_1521,N_4747);
nand U5773 (N_5773,N_1968,N_4914);
and U5774 (N_5774,N_4598,N_3229);
and U5775 (N_5775,N_912,N_4221);
or U5776 (N_5776,N_2095,N_1789);
and U5777 (N_5777,N_2687,N_2122);
and U5778 (N_5778,N_1222,N_3332);
or U5779 (N_5779,N_2835,N_827);
or U5780 (N_5780,N_3648,N_4808);
xnor U5781 (N_5781,N_1741,N_529);
xor U5782 (N_5782,N_1837,N_3432);
nor U5783 (N_5783,N_4234,N_3556);
and U5784 (N_5784,N_2632,N_460);
and U5785 (N_5785,N_3600,N_2293);
or U5786 (N_5786,N_326,N_2542);
or U5787 (N_5787,N_3215,N_2740);
and U5788 (N_5788,N_3914,N_1860);
nand U5789 (N_5789,N_4088,N_64);
xnor U5790 (N_5790,N_4609,N_4078);
or U5791 (N_5791,N_2636,N_3167);
and U5792 (N_5792,N_99,N_3546);
or U5793 (N_5793,N_128,N_2901);
and U5794 (N_5794,N_902,N_3657);
nand U5795 (N_5795,N_4290,N_2465);
nand U5796 (N_5796,N_4661,N_1109);
nor U5797 (N_5797,N_2974,N_4790);
nand U5798 (N_5798,N_399,N_2559);
or U5799 (N_5799,N_2352,N_968);
or U5800 (N_5800,N_1562,N_1205);
and U5801 (N_5801,N_4830,N_4855);
nand U5802 (N_5802,N_3383,N_2321);
and U5803 (N_5803,N_3989,N_2148);
nand U5804 (N_5804,N_1801,N_2133);
nand U5805 (N_5805,N_1209,N_280);
nand U5806 (N_5806,N_3102,N_3789);
or U5807 (N_5807,N_4842,N_4026);
nand U5808 (N_5808,N_2767,N_4152);
or U5809 (N_5809,N_735,N_3457);
nand U5810 (N_5810,N_2515,N_4663);
nand U5811 (N_5811,N_1575,N_2695);
or U5812 (N_5812,N_746,N_2420);
and U5813 (N_5813,N_1908,N_930);
nand U5814 (N_5814,N_3219,N_1074);
nor U5815 (N_5815,N_752,N_2761);
or U5816 (N_5816,N_2703,N_4173);
and U5817 (N_5817,N_74,N_2552);
and U5818 (N_5818,N_821,N_1365);
and U5819 (N_5819,N_760,N_1230);
nor U5820 (N_5820,N_4658,N_4485);
or U5821 (N_5821,N_4030,N_4779);
nor U5822 (N_5822,N_1191,N_1469);
nor U5823 (N_5823,N_3016,N_3395);
and U5824 (N_5824,N_3202,N_4108);
or U5825 (N_5825,N_1888,N_1809);
nand U5826 (N_5826,N_4599,N_101);
nand U5827 (N_5827,N_1486,N_143);
nor U5828 (N_5828,N_4774,N_2252);
and U5829 (N_5829,N_4816,N_4460);
and U5830 (N_5830,N_4139,N_1702);
nand U5831 (N_5831,N_2289,N_3653);
nor U5832 (N_5832,N_187,N_2509);
nor U5833 (N_5833,N_3845,N_4712);
nor U5834 (N_5834,N_1179,N_4509);
xnor U5835 (N_5835,N_4812,N_1898);
or U5836 (N_5836,N_3226,N_1528);
or U5837 (N_5837,N_2138,N_467);
nor U5838 (N_5838,N_85,N_3690);
nand U5839 (N_5839,N_1158,N_2893);
nor U5840 (N_5840,N_149,N_4581);
or U5841 (N_5841,N_2390,N_4080);
nor U5842 (N_5842,N_4383,N_3398);
or U5843 (N_5843,N_4684,N_3066);
or U5844 (N_5844,N_3379,N_1319);
nor U5845 (N_5845,N_272,N_1776);
or U5846 (N_5846,N_3359,N_1902);
nand U5847 (N_5847,N_2962,N_3068);
nor U5848 (N_5848,N_1130,N_2025);
or U5849 (N_5849,N_1154,N_3880);
xor U5850 (N_5850,N_3844,N_1768);
and U5851 (N_5851,N_4333,N_37);
or U5852 (N_5852,N_1031,N_2470);
and U5853 (N_5853,N_2267,N_4223);
nand U5854 (N_5854,N_2178,N_2795);
nor U5855 (N_5855,N_1487,N_3604);
nand U5856 (N_5856,N_1481,N_392);
and U5857 (N_5857,N_3560,N_732);
or U5858 (N_5858,N_2146,N_4611);
nor U5859 (N_5859,N_2501,N_2724);
and U5860 (N_5860,N_2756,N_410);
nor U5861 (N_5861,N_2906,N_1111);
nor U5862 (N_5862,N_565,N_3853);
xor U5863 (N_5863,N_1453,N_1904);
xor U5864 (N_5864,N_4879,N_2939);
or U5865 (N_5865,N_2377,N_4837);
and U5866 (N_5866,N_3952,N_2871);
and U5867 (N_5867,N_3468,N_4897);
nor U5868 (N_5868,N_749,N_3716);
or U5869 (N_5869,N_3353,N_4445);
xor U5870 (N_5870,N_4677,N_1304);
nor U5871 (N_5871,N_317,N_4963);
nor U5872 (N_5872,N_4927,N_676);
nor U5873 (N_5873,N_4384,N_3122);
nand U5874 (N_5874,N_3758,N_4051);
or U5875 (N_5875,N_630,N_4427);
or U5876 (N_5876,N_3311,N_659);
and U5877 (N_5877,N_4229,N_4497);
and U5878 (N_5878,N_4170,N_1349);
xnor U5879 (N_5879,N_4551,N_1152);
xor U5880 (N_5880,N_2668,N_642);
and U5881 (N_5881,N_2368,N_121);
nor U5882 (N_5882,N_708,N_4739);
or U5883 (N_5883,N_1835,N_4983);
nand U5884 (N_5884,N_2127,N_4660);
or U5885 (N_5885,N_800,N_1255);
nor U5886 (N_5886,N_915,N_3382);
nand U5887 (N_5887,N_4846,N_3695);
nand U5888 (N_5888,N_1937,N_2084);
or U5889 (N_5889,N_2074,N_1515);
xnor U5890 (N_5890,N_2118,N_1556);
and U5891 (N_5891,N_3886,N_4902);
nand U5892 (N_5892,N_3364,N_4452);
nor U5893 (N_5893,N_4349,N_1339);
nand U5894 (N_5894,N_3488,N_3577);
nor U5895 (N_5895,N_1347,N_32);
or U5896 (N_5896,N_4500,N_958);
nor U5897 (N_5897,N_2914,N_4579);
nor U5898 (N_5898,N_949,N_1382);
and U5899 (N_5899,N_4461,N_1156);
nand U5900 (N_5900,N_1197,N_2313);
xor U5901 (N_5901,N_4350,N_2814);
or U5902 (N_5902,N_4761,N_2034);
nor U5903 (N_5903,N_2823,N_1168);
nand U5904 (N_5904,N_3539,N_910);
or U5905 (N_5905,N_1797,N_1201);
nand U5906 (N_5906,N_650,N_3079);
and U5907 (N_5907,N_4208,N_4718);
nand U5908 (N_5908,N_4059,N_645);
and U5909 (N_5909,N_3948,N_4856);
xor U5910 (N_5910,N_3164,N_3455);
or U5911 (N_5911,N_71,N_1463);
and U5912 (N_5912,N_1004,N_4628);
nand U5913 (N_5913,N_4976,N_1290);
nand U5914 (N_5914,N_2125,N_3814);
or U5915 (N_5915,N_1591,N_2266);
or U5916 (N_5916,N_1276,N_1206);
or U5917 (N_5917,N_2873,N_2459);
or U5918 (N_5918,N_3040,N_1636);
or U5919 (N_5919,N_3444,N_3828);
and U5920 (N_5920,N_2186,N_4105);
and U5921 (N_5921,N_3060,N_4183);
nand U5922 (N_5922,N_4713,N_1403);
nor U5923 (N_5923,N_1439,N_368);
and U5924 (N_5924,N_992,N_3221);
nor U5925 (N_5925,N_906,N_4434);
nor U5926 (N_5926,N_2500,N_1506);
nand U5927 (N_5927,N_136,N_2706);
nand U5928 (N_5928,N_4783,N_1945);
or U5929 (N_5929,N_1091,N_3983);
xnor U5930 (N_5930,N_3005,N_3250);
nor U5931 (N_5931,N_61,N_89);
nand U5932 (N_5932,N_1440,N_3561);
and U5933 (N_5933,N_1590,N_4244);
xor U5934 (N_5934,N_2430,N_4769);
or U5935 (N_5935,N_3968,N_2857);
nor U5936 (N_5936,N_3581,N_2604);
nand U5937 (N_5937,N_378,N_2268);
nand U5938 (N_5938,N_4570,N_1706);
nor U5939 (N_5939,N_4031,N_1162);
nand U5940 (N_5940,N_274,N_4433);
and U5941 (N_5941,N_4365,N_3193);
nor U5942 (N_5942,N_4479,N_2606);
nand U5943 (N_5943,N_620,N_1155);
nand U5944 (N_5944,N_2455,N_2850);
nor U5945 (N_5945,N_3940,N_3889);
xor U5946 (N_5946,N_3768,N_1592);
or U5947 (N_5947,N_1573,N_1770);
nor U5948 (N_5948,N_1788,N_1134);
or U5949 (N_5949,N_2507,N_67);
xnor U5950 (N_5950,N_3711,N_291);
nand U5951 (N_5951,N_4997,N_4544);
nand U5952 (N_5952,N_3802,N_4261);
nand U5953 (N_5953,N_2783,N_2754);
or U5954 (N_5954,N_1660,N_4860);
and U5955 (N_5955,N_2143,N_1990);
nand U5956 (N_5956,N_4363,N_1656);
nor U5957 (N_5957,N_1298,N_4762);
xnor U5958 (N_5958,N_4616,N_2990);
nor U5959 (N_5959,N_2279,N_629);
xor U5960 (N_5960,N_3148,N_4268);
nor U5961 (N_5961,N_36,N_176);
and U5962 (N_5962,N_4932,N_1666);
and U5963 (N_5963,N_4701,N_360);
and U5964 (N_5964,N_3507,N_3922);
nor U5965 (N_5965,N_1633,N_2965);
nor U5966 (N_5966,N_2080,N_527);
and U5967 (N_5967,N_4144,N_203);
or U5968 (N_5968,N_2258,N_3376);
and U5969 (N_5969,N_3926,N_156);
nor U5970 (N_5970,N_2156,N_1831);
nand U5971 (N_5971,N_468,N_4793);
nand U5972 (N_5972,N_1249,N_3462);
nand U5973 (N_5973,N_554,N_3418);
and U5974 (N_5974,N_3638,N_4066);
and U5975 (N_5975,N_3835,N_1886);
nor U5976 (N_5976,N_137,N_2697);
nand U5977 (N_5977,N_4534,N_626);
nand U5978 (N_5978,N_4207,N_1316);
xnor U5979 (N_5979,N_448,N_4491);
or U5980 (N_5980,N_4099,N_3614);
and U5981 (N_5981,N_1497,N_547);
and U5982 (N_5982,N_4786,N_2402);
xor U5983 (N_5983,N_3222,N_1885);
or U5984 (N_5984,N_3705,N_2955);
and U5985 (N_5985,N_355,N_2700);
nand U5986 (N_5986,N_4119,N_2799);
nand U5987 (N_5987,N_4197,N_4390);
nor U5988 (N_5988,N_1989,N_4035);
nand U5989 (N_5989,N_3161,N_4700);
nand U5990 (N_5990,N_2351,N_2683);
xor U5991 (N_5991,N_2229,N_983);
nand U5992 (N_5992,N_4454,N_465);
nor U5993 (N_5993,N_3237,N_3439);
nand U5994 (N_5994,N_2698,N_1538);
xor U5995 (N_5995,N_2504,N_1977);
and U5996 (N_5996,N_972,N_1513);
or U5997 (N_5997,N_1392,N_4143);
and U5998 (N_5998,N_3954,N_4257);
and U5999 (N_5999,N_4549,N_3130);
or U6000 (N_6000,N_1559,N_667);
nand U6001 (N_6001,N_2613,N_336);
or U6002 (N_6002,N_4295,N_2892);
nor U6003 (N_6003,N_4723,N_133);
nand U6004 (N_6004,N_3304,N_2033);
or U6005 (N_6005,N_2665,N_3091);
nand U6006 (N_6006,N_2652,N_3787);
nand U6007 (N_6007,N_3162,N_3121);
nor U6008 (N_6008,N_3183,N_2988);
nand U6009 (N_6009,N_477,N_3715);
and U6010 (N_6010,N_951,N_796);
and U6011 (N_6011,N_1196,N_2964);
nor U6012 (N_6012,N_2001,N_3319);
nor U6013 (N_6013,N_1410,N_3285);
and U6014 (N_6014,N_2441,N_1804);
nand U6015 (N_6015,N_4859,N_3877);
nor U6016 (N_6016,N_4246,N_52);
and U6017 (N_6017,N_2046,N_4767);
and U6018 (N_6018,N_2388,N_1305);
and U6019 (N_6019,N_1189,N_4671);
nor U6020 (N_6020,N_4638,N_2998);
and U6021 (N_6021,N_3207,N_3428);
and U6022 (N_6022,N_4928,N_132);
and U6023 (N_6023,N_4135,N_1343);
nor U6024 (N_6024,N_913,N_2479);
or U6025 (N_6025,N_4833,N_457);
and U6026 (N_6026,N_2308,N_2083);
and U6027 (N_6027,N_4046,N_1166);
nor U6028 (N_6028,N_4032,N_4202);
nor U6029 (N_6029,N_2819,N_4618);
nor U6030 (N_6030,N_1470,N_1790);
nor U6031 (N_6031,N_1376,N_4513);
nor U6032 (N_6032,N_2379,N_741);
and U6033 (N_6033,N_1764,N_1889);
xnor U6034 (N_6034,N_2966,N_1974);
or U6035 (N_6035,N_72,N_430);
and U6036 (N_6036,N_8,N_4463);
xnor U6037 (N_6037,N_541,N_3838);
nand U6038 (N_6038,N_4979,N_4346);
nand U6039 (N_6039,N_1846,N_4017);
nor U6040 (N_6040,N_2986,N_933);
and U6041 (N_6041,N_352,N_4103);
or U6042 (N_6042,N_3563,N_2644);
nand U6043 (N_6043,N_1853,N_4200);
nor U6044 (N_6044,N_1733,N_4288);
and U6045 (N_6045,N_1126,N_4072);
xor U6046 (N_6046,N_4326,N_161);
and U6047 (N_6047,N_455,N_1492);
nor U6048 (N_6048,N_412,N_4993);
and U6049 (N_6049,N_976,N_2693);
or U6050 (N_6050,N_334,N_4308);
or U6051 (N_6051,N_3761,N_4882);
or U6052 (N_6052,N_2019,N_2468);
nor U6053 (N_6053,N_515,N_2456);
nand U6054 (N_6054,N_2882,N_4436);
or U6055 (N_6055,N_2657,N_4038);
or U6056 (N_6056,N_1099,N_387);
nor U6057 (N_6057,N_717,N_2278);
or U6058 (N_6058,N_409,N_3228);
and U6059 (N_6059,N_2662,N_2595);
or U6060 (N_6060,N_1587,N_853);
nand U6061 (N_6061,N_2560,N_1649);
or U6062 (N_6062,N_3509,N_2432);
xnor U6063 (N_6063,N_3482,N_3424);
xor U6064 (N_6064,N_623,N_4503);
and U6065 (N_6065,N_3302,N_756);
nor U6066 (N_6066,N_2635,N_4870);
or U6067 (N_6067,N_1838,N_4580);
xnor U6068 (N_6068,N_539,N_3052);
nor U6069 (N_6069,N_1132,N_2717);
and U6070 (N_6070,N_2399,N_4359);
and U6071 (N_6071,N_3021,N_3141);
or U6072 (N_6072,N_1940,N_2417);
nor U6073 (N_6073,N_4282,N_4916);
xor U6074 (N_6074,N_3259,N_2716);
and U6075 (N_6075,N_2037,N_4425);
xor U6076 (N_6076,N_570,N_3700);
nand U6077 (N_6077,N_3056,N_3384);
nor U6078 (N_6078,N_4892,N_3240);
or U6079 (N_6079,N_3172,N_370);
or U6080 (N_6080,N_1700,N_2361);
xor U6081 (N_6081,N_3367,N_2931);
nand U6082 (N_6082,N_2128,N_1214);
xnor U6083 (N_6083,N_3165,N_4770);
nor U6084 (N_6084,N_1897,N_698);
nand U6085 (N_6085,N_3818,N_2336);
or U6086 (N_6086,N_2395,N_1411);
nor U6087 (N_6087,N_4306,N_3805);
nand U6088 (N_6088,N_1572,N_3212);
nor U6089 (N_6089,N_4744,N_1757);
nand U6090 (N_6090,N_2061,N_4967);
nand U6091 (N_6091,N_463,N_1664);
nand U6092 (N_6092,N_2707,N_1294);
nand U6093 (N_6093,N_868,N_4894);
nand U6094 (N_6094,N_4806,N_3131);
nand U6095 (N_6095,N_3286,N_2983);
nand U6096 (N_6096,N_2841,N_3735);
or U6097 (N_6097,N_2561,N_1655);
nand U6098 (N_6098,N_306,N_521);
and U6099 (N_6099,N_1468,N_3824);
nor U6100 (N_6100,N_2985,N_771);
and U6101 (N_6101,N_803,N_1296);
nand U6102 (N_6102,N_2341,N_1013);
nor U6103 (N_6103,N_9,N_4444);
nor U6104 (N_6104,N_1697,N_2022);
or U6105 (N_6105,N_3928,N_859);
and U6106 (N_6106,N_4335,N_792);
nor U6107 (N_6107,N_1517,N_2666);
nor U6108 (N_6108,N_281,N_4686);
nor U6109 (N_6109,N_1630,N_1891);
or U6110 (N_6110,N_561,N_2743);
or U6111 (N_6111,N_1914,N_3355);
nor U6112 (N_6112,N_3737,N_95);
nand U6113 (N_6113,N_4232,N_4596);
nand U6114 (N_6114,N_3244,N_3309);
and U6115 (N_6115,N_3324,N_2813);
nor U6116 (N_6116,N_1435,N_1966);
or U6117 (N_6117,N_1735,N_4889);
nand U6118 (N_6118,N_2016,N_1079);
nand U6119 (N_6119,N_2895,N_1170);
or U6120 (N_6120,N_429,N_3592);
and U6121 (N_6121,N_4382,N_4499);
xor U6122 (N_6122,N_3541,N_3822);
or U6123 (N_6123,N_255,N_2539);
nand U6124 (N_6124,N_2851,N_742);
nor U6125 (N_6125,N_2910,N_1696);
nand U6126 (N_6126,N_1186,N_2207);
and U6127 (N_6127,N_4873,N_731);
xor U6128 (N_6128,N_4631,N_1557);
nand U6129 (N_6129,N_3179,N_2935);
or U6130 (N_6130,N_2583,N_3910);
and U6131 (N_6131,N_4554,N_4584);
nand U6132 (N_6132,N_545,N_4898);
nand U6133 (N_6133,N_3596,N_2071);
nand U6134 (N_6134,N_3372,N_3586);
or U6135 (N_6135,N_2330,N_3588);
and U6136 (N_6136,N_2862,N_2328);
nand U6137 (N_6137,N_170,N_588);
or U6138 (N_6138,N_3727,N_2248);
and U6139 (N_6139,N_2428,N_2227);
xnor U6140 (N_6140,N_3631,N_2269);
nor U6141 (N_6141,N_4802,N_808);
or U6142 (N_6142,N_407,N_1648);
or U6143 (N_6143,N_3942,N_78);
and U6144 (N_6144,N_4571,N_2197);
nand U6145 (N_6145,N_780,N_643);
nor U6146 (N_6146,N_197,N_2580);
nor U6147 (N_6147,N_3520,N_4094);
nand U6148 (N_6148,N_4796,N_294);
and U6149 (N_6149,N_1393,N_2678);
or U6150 (N_6150,N_2062,N_1357);
nor U6151 (N_6151,N_689,N_4546);
and U6152 (N_6152,N_1893,N_4380);
xor U6153 (N_6153,N_3902,N_897);
nor U6154 (N_6154,N_4109,N_2803);
nor U6155 (N_6155,N_1078,N_4432);
or U6156 (N_6156,N_3019,N_303);
xnor U6157 (N_6157,N_4300,N_4052);
and U6158 (N_6158,N_4775,N_3316);
or U6159 (N_6159,N_1277,N_1627);
xor U6160 (N_6160,N_1067,N_2086);
nor U6161 (N_6161,N_816,N_4637);
nor U6162 (N_6162,N_2533,N_2993);
nor U6163 (N_6163,N_1526,N_289);
xnor U6164 (N_6164,N_3294,N_2784);
and U6165 (N_6165,N_920,N_3406);
or U6166 (N_6166,N_2741,N_1720);
or U6167 (N_6167,N_1755,N_1531);
and U6168 (N_6168,N_4562,N_2311);
xnor U6169 (N_6169,N_879,N_3767);
nand U6170 (N_6170,N_1596,N_1786);
nor U6171 (N_6171,N_825,N_1232);
nor U6172 (N_6172,N_3308,N_4003);
nor U6173 (N_6173,N_4319,N_4047);
xor U6174 (N_6174,N_2057,N_2691);
and U6175 (N_6175,N_1611,N_3726);
and U6176 (N_6176,N_2488,N_2729);
and U6177 (N_6177,N_2600,N_2768);
nor U6178 (N_6178,N_748,N_3554);
nor U6179 (N_6179,N_458,N_1272);
nor U6180 (N_6180,N_1564,N_1247);
and U6181 (N_6181,N_1792,N_4748);
and U6182 (N_6182,N_1034,N_319);
nand U6183 (N_6183,N_3358,N_610);
nor U6184 (N_6184,N_3192,N_2056);
and U6185 (N_6185,N_2353,N_198);
nor U6186 (N_6186,N_4715,N_1652);
and U6187 (N_6187,N_4250,N_2810);
or U6188 (N_6188,N_1019,N_2607);
nand U6189 (N_6189,N_2300,N_1558);
or U6190 (N_6190,N_2621,N_1925);
nor U6191 (N_6191,N_1713,N_1280);
nor U6192 (N_6192,N_2213,N_1188);
and U6193 (N_6193,N_3756,N_4760);
nor U6194 (N_6194,N_2386,N_4116);
nand U6195 (N_6195,N_1767,N_2169);
and U6196 (N_6196,N_4646,N_3305);
nor U6197 (N_6197,N_4216,N_3841);
nand U6198 (N_6198,N_2860,N_3231);
xnor U6199 (N_6199,N_2265,N_3065);
nor U6200 (N_6200,N_1260,N_899);
nor U6201 (N_6201,N_935,N_4253);
nor U6202 (N_6202,N_3205,N_3186);
nor U6203 (N_6203,N_3580,N_1383);
or U6204 (N_6204,N_2680,N_3209);
or U6205 (N_6205,N_2726,N_751);
nand U6206 (N_6206,N_252,N_4162);
or U6207 (N_6207,N_1576,N_3988);
nand U6208 (N_6208,N_2961,N_2578);
or U6209 (N_6209,N_4093,N_2124);
nor U6210 (N_6210,N_4541,N_1234);
or U6211 (N_6211,N_3119,N_3766);
or U6212 (N_6212,N_3511,N_1737);
xnor U6213 (N_6213,N_793,N_679);
nand U6214 (N_6214,N_1391,N_1195);
or U6215 (N_6215,N_3138,N_3336);
xor U6216 (N_6216,N_3292,N_2018);
nand U6217 (N_6217,N_3636,N_1998);
nand U6218 (N_6218,N_4765,N_1863);
xnor U6219 (N_6219,N_310,N_2054);
nand U6220 (N_6220,N_1207,N_4995);
and U6221 (N_6221,N_562,N_3572);
or U6222 (N_6222,N_1695,N_2926);
nand U6223 (N_6223,N_4613,N_618);
and U6224 (N_6224,N_1542,N_3423);
and U6225 (N_6225,N_3006,N_665);
nor U6226 (N_6226,N_3421,N_4567);
and U6227 (N_6227,N_4845,N_726);
and U6228 (N_6228,N_2855,N_3073);
and U6229 (N_6229,N_4623,N_2113);
nand U6230 (N_6230,N_3501,N_4643);
nand U6231 (N_6231,N_3900,N_4138);
nor U6232 (N_6232,N_699,N_925);
or U6233 (N_6233,N_167,N_4236);
nand U6234 (N_6234,N_1064,N_786);
and U6235 (N_6235,N_2762,N_3105);
or U6236 (N_6236,N_3331,N_1190);
and U6237 (N_6237,N_1371,N_4238);
xor U6238 (N_6238,N_3849,N_1820);
xor U6239 (N_6239,N_1900,N_11);
nand U6240 (N_6240,N_3682,N_4224);
nand U6241 (N_6241,N_984,N_297);
nand U6242 (N_6242,N_895,N_1536);
nand U6243 (N_6243,N_714,N_258);
nor U6244 (N_6244,N_3134,N_2856);
or U6245 (N_6245,N_797,N_4725);
and U6246 (N_6246,N_1328,N_1160);
xnor U6247 (N_6247,N_2773,N_4881);
and U6248 (N_6248,N_2870,N_4455);
nand U6249 (N_6249,N_3323,N_936);
or U6250 (N_6250,N_4582,N_3453);
or U6251 (N_6251,N_2262,N_3897);
or U6252 (N_6252,N_1317,N_1604);
nor U6253 (N_6253,N_613,N_235);
nor U6254 (N_6254,N_1313,N_2032);
nor U6255 (N_6255,N_4607,N_4428);
and U6256 (N_6256,N_2005,N_4423);
xor U6257 (N_6257,N_4307,N_861);
or U6258 (N_6258,N_535,N_2643);
nor U6259 (N_6259,N_2834,N_695);
nor U6260 (N_6260,N_3001,N_1116);
nand U6261 (N_6261,N_1070,N_4311);
nor U6262 (N_6262,N_4159,N_3008);
nand U6263 (N_6263,N_1948,N_1100);
xnor U6264 (N_6264,N_1227,N_3261);
nand U6265 (N_6265,N_2530,N_4185);
xnor U6266 (N_6266,N_1876,N_2640);
nand U6267 (N_6267,N_1084,N_1546);
nand U6268 (N_6268,N_4839,N_103);
xnor U6269 (N_6269,N_2383,N_1765);
and U6270 (N_6270,N_4113,N_4735);
nand U6271 (N_6271,N_4493,N_265);
nor U6272 (N_6272,N_869,N_204);
and U6273 (N_6273,N_1631,N_3171);
or U6274 (N_6274,N_418,N_566);
nor U6275 (N_6275,N_3794,N_787);
or U6276 (N_6276,N_3866,N_776);
and U6277 (N_6277,N_3022,N_905);
and U6278 (N_6278,N_4327,N_106);
or U6279 (N_6279,N_711,N_988);
or U6280 (N_6280,N_2527,N_117);
and U6281 (N_6281,N_3069,N_2573);
or U6282 (N_6282,N_1243,N_357);
or U6283 (N_6283,N_4896,N_4386);
nand U6284 (N_6284,N_2584,N_2200);
or U6285 (N_6285,N_249,N_1024);
or U6286 (N_6286,N_781,N_1414);
and U6287 (N_6287,N_2889,N_4351);
or U6288 (N_6288,N_3883,N_4591);
xnor U6289 (N_6289,N_4829,N_1779);
or U6290 (N_6290,N_2868,N_4421);
and U6291 (N_6291,N_1373,N_425);
nand U6292 (N_6292,N_3089,N_2579);
or U6293 (N_6293,N_852,N_295);
and U6294 (N_6294,N_3644,N_1740);
or U6295 (N_6295,N_361,N_1182);
or U6296 (N_6296,N_1639,N_4566);
nand U6297 (N_6297,N_2526,N_724);
xor U6298 (N_6298,N_3325,N_4511);
and U6299 (N_6299,N_2872,N_3206);
nor U6300 (N_6300,N_4227,N_1520);
nor U6301 (N_6301,N_4522,N_3785);
nor U6302 (N_6302,N_4953,N_1550);
nand U6303 (N_6303,N_337,N_4249);
nor U6304 (N_6304,N_514,N_1719);
or U6305 (N_6305,N_3142,N_4086);
nor U6306 (N_6306,N_2049,N_2807);
nand U6307 (N_6307,N_2694,N_4309);
and U6308 (N_6308,N_3562,N_1364);
nor U6309 (N_6309,N_2097,N_3855);
xor U6310 (N_6310,N_4849,N_3555);
nand U6311 (N_6311,N_2546,N_828);
and U6312 (N_6312,N_365,N_3826);
nand U6313 (N_6313,N_279,N_1199);
or U6314 (N_6314,N_4129,N_4347);
nand U6315 (N_6315,N_122,N_673);
or U6316 (N_6316,N_3042,N_3360);
or U6317 (N_6317,N_339,N_1712);
nand U6318 (N_6318,N_3696,N_4381);
nand U6319 (N_6319,N_1828,N_3320);
and U6320 (N_6320,N_590,N_3299);
or U6321 (N_6321,N_3660,N_2324);
or U6322 (N_6322,N_2779,N_3018);
nand U6323 (N_6323,N_1402,N_4824);
and U6324 (N_6324,N_65,N_2150);
nor U6325 (N_6325,N_277,N_3953);
and U6326 (N_6326,N_548,N_469);
nor U6327 (N_6327,N_4973,N_3958);
and U6328 (N_6328,N_2587,N_2836);
or U6329 (N_6329,N_1803,N_3437);
nand U6330 (N_6330,N_4826,N_1651);
or U6331 (N_6331,N_2995,N_4315);
nand U6332 (N_6332,N_251,N_2035);
and U6333 (N_6333,N_981,N_1552);
nand U6334 (N_6334,N_3199,N_1464);
nand U6335 (N_6335,N_2387,N_3429);
nor U6336 (N_6336,N_3574,N_2992);
or U6337 (N_6337,N_2220,N_269);
and U6338 (N_6338,N_3108,N_3890);
xnor U6339 (N_6339,N_2451,N_134);
nand U6340 (N_6340,N_300,N_1169);
or U6341 (N_6341,N_2296,N_2849);
and U6342 (N_6342,N_1005,N_2232);
or U6343 (N_6343,N_506,N_1516);
and U6344 (N_6344,N_1963,N_1301);
and U6345 (N_6345,N_3407,N_2489);
and U6346 (N_6346,N_2797,N_3731);
and U6347 (N_6347,N_1270,N_1366);
and U6348 (N_6348,N_2788,N_3719);
nor U6349 (N_6349,N_918,N_2445);
nand U6350 (N_6350,N_3908,N_3595);
nand U6351 (N_6351,N_4313,N_486);
and U6352 (N_6352,N_3865,N_2503);
nand U6353 (N_6353,N_3178,N_1256);
nand U6354 (N_6354,N_2928,N_4642);
nor U6355 (N_6355,N_2389,N_4366);
xor U6356 (N_6356,N_1242,N_1418);
nand U6357 (N_6357,N_4408,N_3869);
nand U6358 (N_6358,N_2874,N_3441);
and U6359 (N_6359,N_1233,N_439);
or U6360 (N_6360,N_2596,N_243);
nor U6361 (N_6361,N_4377,N_558);
nor U6362 (N_6362,N_2815,N_4994);
and U6363 (N_6363,N_4420,N_1862);
and U6364 (N_6364,N_4203,N_4998);
or U6365 (N_6365,N_4459,N_4633);
nand U6366 (N_6366,N_338,N_4243);
or U6367 (N_6367,N_1061,N_2209);
nor U6368 (N_6368,N_1791,N_3876);
nor U6369 (N_6369,N_3996,N_257);
nor U6370 (N_6370,N_3742,N_1210);
nor U6371 (N_6371,N_3957,N_4970);
xnor U6372 (N_6372,N_651,N_3525);
nor U6373 (N_6373,N_4863,N_3671);
or U6374 (N_6374,N_2221,N_1918);
and U6375 (N_6375,N_4595,N_3394);
nand U6376 (N_6376,N_4343,N_1509);
nor U6377 (N_6377,N_4565,N_1622);
nor U6378 (N_6378,N_2315,N_3851);
nor U6379 (N_6379,N_2521,N_4357);
nor U6380 (N_6380,N_3077,N_1503);
nor U6381 (N_6381,N_3014,N_490);
and U6382 (N_6382,N_4395,N_519);
nand U6383 (N_6383,N_1653,N_1016);
nand U6384 (N_6384,N_509,N_4788);
nand U6385 (N_6385,N_3672,N_809);
and U6386 (N_6386,N_4610,N_4220);
or U6387 (N_6387,N_4469,N_3783);
xnor U6388 (N_6388,N_4648,N_3330);
nand U6389 (N_6389,N_649,N_2671);
xnor U6390 (N_6390,N_1036,N_1075);
or U6391 (N_6391,N_2753,N_2366);
nor U6392 (N_6392,N_3782,N_702);
nor U6393 (N_6393,N_584,N_658);
and U6394 (N_6394,N_2674,N_4075);
or U6395 (N_6395,N_3774,N_96);
and U6396 (N_6396,N_452,N_4068);
nand U6397 (N_6397,N_3732,N_2294);
or U6398 (N_6398,N_1183,N_1096);
and U6399 (N_6399,N_1907,N_94);
or U6400 (N_6400,N_4114,N_4535);
nor U6401 (N_6401,N_3343,N_898);
and U6402 (N_6402,N_3913,N_3575);
and U6403 (N_6403,N_1103,N_3111);
nand U6404 (N_6404,N_2749,N_165);
and U6405 (N_6405,N_1421,N_180);
and U6406 (N_6406,N_4147,N_1916);
nor U6407 (N_6407,N_585,N_4136);
or U6408 (N_6408,N_2611,N_2980);
nand U6409 (N_6409,N_2701,N_1589);
nand U6410 (N_6410,N_4627,N_2052);
nand U6411 (N_6411,N_3530,N_3807);
nor U6412 (N_6412,N_1342,N_826);
nand U6413 (N_6413,N_1356,N_4371);
xnor U6414 (N_6414,N_606,N_3404);
nand U6415 (N_6415,N_3635,N_1475);
nand U6416 (N_6416,N_3157,N_1581);
nand U6417 (N_6417,N_4728,N_1146);
or U6418 (N_6418,N_4403,N_860);
xnor U6419 (N_6419,N_4110,N_567);
xor U6420 (N_6420,N_1408,N_1969);
nand U6421 (N_6421,N_3585,N_4305);
nand U6422 (N_6422,N_2008,N_4732);
nand U6423 (N_6423,N_2531,N_3524);
nor U6424 (N_6424,N_304,N_1119);
nor U6425 (N_6425,N_2218,N_1670);
or U6426 (N_6426,N_3770,N_1394);
nand U6427 (N_6427,N_4394,N_2360);
nand U6428 (N_6428,N_4475,N_4239);
and U6429 (N_6429,N_1263,N_4172);
and U6430 (N_6430,N_2787,N_1465);
nand U6431 (N_6431,N_1291,N_4612);
or U6432 (N_6432,N_4931,N_1363);
xor U6433 (N_6433,N_1459,N_1139);
xnor U6434 (N_6434,N_2905,N_1374);
and U6435 (N_6435,N_3976,N_1325);
nor U6436 (N_6436,N_2863,N_3289);
or U6437 (N_6437,N_4778,N_1778);
and U6438 (N_6438,N_1035,N_569);
nor U6439 (N_6439,N_3790,N_4063);
nor U6440 (N_6440,N_3603,N_2464);
and U6441 (N_6441,N_22,N_3481);
or U6442 (N_6442,N_871,N_2645);
and U6443 (N_6443,N_1535,N_4919);
and U6444 (N_6444,N_4733,N_3759);
nand U6445 (N_6445,N_4385,N_525);
xor U6446 (N_6446,N_2011,N_2811);
nand U6447 (N_6447,N_957,N_1460);
or U6448 (N_6448,N_2063,N_229);
nor U6449 (N_6449,N_4665,N_2181);
or U6450 (N_6450,N_205,N_4042);
nor U6451 (N_6451,N_4048,N_4422);
nand U6452 (N_6452,N_3949,N_3116);
nand U6453 (N_6453,N_3047,N_1934);
nor U6454 (N_6454,N_3045,N_594);
xnor U6455 (N_6455,N_2301,N_785);
nand U6456 (N_6456,N_943,N_115);
nor U6457 (N_6457,N_845,N_4518);
xnor U6458 (N_6458,N_173,N_3526);
nor U6459 (N_6459,N_92,N_3714);
nor U6460 (N_6460,N_2801,N_474);
nor U6461 (N_6461,N_942,N_3200);
and U6462 (N_6462,N_3127,N_989);
xnor U6463 (N_6463,N_2658,N_1445);
and U6464 (N_6464,N_3257,N_1361);
or U6465 (N_6465,N_4074,N_1743);
nor U6466 (N_6466,N_3781,N_4868);
nor U6467 (N_6467,N_1385,N_3755);
xor U6468 (N_6468,N_1355,N_2204);
nor U6469 (N_6469,N_1148,N_3548);
or U6470 (N_6470,N_2121,N_4556);
and U6471 (N_6471,N_47,N_3945);
or U6472 (N_6472,N_189,N_4400);
and U6473 (N_6473,N_2817,N_2233);
and U6474 (N_6474,N_3610,N_978);
nor U6475 (N_6475,N_687,N_1568);
nand U6476 (N_6476,N_3677,N_2101);
xnor U6477 (N_6477,N_4222,N_1405);
nor U6478 (N_6478,N_1756,N_1454);
nand U6479 (N_6479,N_1805,N_4682);
or U6480 (N_6480,N_4149,N_2627);
xnor U6481 (N_6481,N_3981,N_579);
nor U6482 (N_6482,N_1007,N_3873);
nor U6483 (N_6483,N_58,N_3713);
nor U6484 (N_6484,N_892,N_4827);
or U6485 (N_6485,N_3281,N_332);
nor U6486 (N_6486,N_3769,N_4742);
nand U6487 (N_6487,N_398,N_3487);
or U6488 (N_6488,N_1327,N_3256);
or U6489 (N_6489,N_4199,N_3646);
and U6490 (N_6490,N_2822,N_4819);
or U6491 (N_6491,N_4069,N_3784);
nand U6492 (N_6492,N_3469,N_1638);
and U6493 (N_6493,N_491,N_3675);
nand U6494 (N_6494,N_461,N_1961);
and U6495 (N_6495,N_2796,N_3601);
nor U6496 (N_6496,N_3519,N_4621);
or U6497 (N_6497,N_2314,N_363);
or U6498 (N_6498,N_110,N_3029);
nand U6499 (N_6499,N_3912,N_682);
xnor U6500 (N_6500,N_4464,N_644);
nor U6501 (N_6501,N_4803,N_3527);
nor U6502 (N_6502,N_4698,N_4196);
or U6503 (N_6503,N_4880,N_3997);
nand U6504 (N_6504,N_3297,N_632);
xor U6505 (N_6505,N_1511,N_3825);
xnor U6506 (N_6506,N_1198,N_1478);
nand U6507 (N_6507,N_1997,N_2733);
and U6508 (N_6508,N_2179,N_1164);
xnor U6509 (N_6509,N_364,N_3163);
nand U6510 (N_6510,N_3856,N_2866);
nor U6511 (N_6511,N_2170,N_2525);
nand U6512 (N_6512,N_2075,N_2136);
nor U6513 (N_6513,N_1579,N_3786);
nor U6514 (N_6514,N_2997,N_4304);
and U6515 (N_6515,N_2335,N_656);
nand U6516 (N_6516,N_4278,N_4154);
nand U6517 (N_6517,N_1623,N_2624);
or U6518 (N_6518,N_375,N_3626);
xor U6519 (N_6519,N_2886,N_2735);
and U6520 (N_6520,N_553,N_1634);
xor U6521 (N_6521,N_1707,N_4923);
xor U6522 (N_6522,N_172,N_4435);
nor U6523 (N_6523,N_4675,N_4558);
nand U6524 (N_6524,N_824,N_3135);
and U6525 (N_6525,N_4869,N_2303);
nor U6526 (N_6526,N_2188,N_1956);
and U6527 (N_6527,N_1021,N_1823);
nor U6528 (N_6528,N_1212,N_1602);
and U6529 (N_6529,N_3536,N_1398);
or U6530 (N_6530,N_1705,N_2307);
xor U6531 (N_6531,N_1825,N_98);
nand U6532 (N_6532,N_4877,N_2098);
nand U6533 (N_6533,N_1691,N_2256);
and U6534 (N_6534,N_3652,N_2820);
nor U6535 (N_6535,N_4213,N_3977);
and U6536 (N_6536,N_1810,N_926);
nor U6537 (N_6537,N_4097,N_1045);
or U6538 (N_6538,N_4010,N_3393);
xor U6539 (N_6539,N_1541,N_1185);
nand U6540 (N_6540,N_4850,N_15);
and U6541 (N_6541,N_1297,N_639);
and U6542 (N_6542,N_564,N_390);
xor U6543 (N_6543,N_4178,N_3195);
nor U6544 (N_6544,N_453,N_769);
nand U6545 (N_6545,N_3041,N_3396);
nor U6546 (N_6546,N_863,N_3238);
or U6547 (N_6547,N_627,N_4439);
or U6548 (N_6548,N_2397,N_3963);
nor U6549 (N_6549,N_3472,N_2144);
and U6550 (N_6550,N_3145,N_2190);
nand U6551 (N_6551,N_1612,N_3132);
or U6552 (N_6552,N_2318,N_4417);
or U6553 (N_6553,N_4822,N_997);
or U6554 (N_6554,N_2298,N_3871);
xor U6555 (N_6555,N_3987,N_1584);
nand U6556 (N_6556,N_522,N_4590);
xnor U6557 (N_6557,N_881,N_3344);
nor U6558 (N_6558,N_1396,N_4020);
and U6559 (N_6559,N_1378,N_3803);
and U6560 (N_6560,N_4533,N_961);
and U6561 (N_6561,N_4292,N_420);
or U6562 (N_6562,N_2499,N_3860);
nand U6563 (N_6563,N_3133,N_1106);
or U6564 (N_6564,N_2705,N_555);
xor U6565 (N_6565,N_2245,N_245);
and U6566 (N_6566,N_777,N_829);
or U6567 (N_6567,N_225,N_4798);
xor U6568 (N_6568,N_1488,N_4834);
nor U6569 (N_6569,N_4095,N_4601);
and U6570 (N_6570,N_1138,N_647);
or U6571 (N_6571,N_4930,N_766);
nor U6572 (N_6572,N_4006,N_4530);
nand U6573 (N_6573,N_391,N_4279);
or U6574 (N_6574,N_1704,N_538);
nand U6575 (N_6575,N_4271,N_1608);
nand U6576 (N_6576,N_1011,N_2367);
and U6577 (N_6577,N_2414,N_369);
nand U6578 (N_6578,N_719,N_4369);
nand U6579 (N_6579,N_909,N_3435);
nand U6580 (N_6580,N_4557,N_3438);
xnor U6581 (N_6581,N_346,N_2712);
and U6582 (N_6582,N_700,N_1815);
and U6583 (N_6583,N_587,N_3961);
xor U6584 (N_6584,N_4276,N_4755);
nor U6585 (N_6585,N_349,N_2021);
nor U6586 (N_6586,N_882,N_1261);
and U6587 (N_6587,N_779,N_2453);
or U6588 (N_6588,N_2745,N_348);
and U6589 (N_6589,N_2139,N_3086);
and U6590 (N_6590,N_1882,N_4956);
and U6591 (N_6591,N_4867,N_499);
nand U6592 (N_6592,N_3296,N_1372);
nand U6593 (N_6593,N_1946,N_4987);
or U6594 (N_6594,N_3194,N_4667);
and U6595 (N_6595,N_2661,N_2846);
or U6596 (N_6596,N_3071,N_1040);
nor U6597 (N_6597,N_2925,N_3709);
nand U6598 (N_6598,N_3602,N_4158);
xor U6599 (N_6599,N_1380,N_4574);
nor U6600 (N_6600,N_2115,N_4041);
and U6601 (N_6601,N_436,N_466);
and U6602 (N_6602,N_3450,N_3884);
xnor U6603 (N_6603,N_2718,N_896);
or U6604 (N_6604,N_4645,N_686);
and U6605 (N_6605,N_7,N_4776);
or U6606 (N_6606,N_1274,N_3827);
or U6607 (N_6607,N_921,N_1514);
nand U6608 (N_6608,N_3683,N_3959);
nor U6609 (N_6609,N_3057,N_1812);
xor U6610 (N_6610,N_4084,N_443);
xnor U6611 (N_6611,N_4524,N_2625);
nor U6612 (N_6612,N_3267,N_2528);
xor U6613 (N_6613,N_4647,N_633);
nand U6614 (N_6614,N_4092,N_1854);
nand U6615 (N_6615,N_2522,N_4676);
nand U6616 (N_6616,N_1668,N_4726);
and U6617 (N_6617,N_4418,N_4001);
nor U6618 (N_6618,N_2476,N_3150);
nor U6619 (N_6619,N_1501,N_4899);
nor U6620 (N_6620,N_1108,N_3084);
nor U6621 (N_6621,N_395,N_228);
nand U6622 (N_6622,N_4065,N_1646);
nand U6623 (N_6623,N_4651,N_1530);
xor U6624 (N_6624,N_3499,N_599);
and U6625 (N_6625,N_2235,N_1844);
or U6626 (N_6626,N_68,N_4484);
xor U6627 (N_6627,N_1181,N_3492);
and U6628 (N_6628,N_3833,N_4569);
nand U6629 (N_6629,N_1012,N_3099);
or U6630 (N_6630,N_3225,N_2759);
nand U6631 (N_6631,N_996,N_4176);
and U6632 (N_6632,N_4939,N_3002);
or U6633 (N_6633,N_4781,N_814);
or U6634 (N_6634,N_3899,N_2593);
nor U6635 (N_6635,N_345,N_3258);
nand U6636 (N_6636,N_2393,N_1999);
nor U6637 (N_6637,N_4668,N_798);
nand U6638 (N_6638,N_4211,N_1081);
nand U6639 (N_6639,N_3155,N_1231);
and U6640 (N_6640,N_3655,N_2941);
xor U6641 (N_6641,N_2394,N_4605);
or U6642 (N_6642,N_1090,N_321);
nand U6643 (N_6643,N_3516,N_3752);
and U6644 (N_6644,N_3048,N_2490);
and U6645 (N_6645,N_3017,N_1565);
nand U6646 (N_6646,N_3034,N_2484);
xnor U6647 (N_6647,N_4729,N_3370);
nand U6648 (N_6648,N_1926,N_2709);
and U6649 (N_6649,N_4167,N_3670);
and U6650 (N_6650,N_2363,N_470);
nor U6651 (N_6651,N_419,N_4325);
and U6652 (N_6652,N_3678,N_4);
or U6653 (N_6653,N_2349,N_568);
nor U6654 (N_6654,N_2247,N_4237);
or U6655 (N_6655,N_472,N_2160);
nor U6656 (N_6656,N_3235,N_4506);
nand U6657 (N_6657,N_1424,N_3189);
nand U6658 (N_6658,N_4861,N_2766);
and U6659 (N_6659,N_2806,N_1092);
nor U6660 (N_6660,N_2641,N_616);
or U6661 (N_6661,N_754,N_1502);
or U6662 (N_6662,N_3616,N_1288);
or U6663 (N_6663,N_1124,N_3094);
nand U6664 (N_6664,N_4772,N_2752);
nor U6665 (N_6665,N_2924,N_2780);
and U6666 (N_6666,N_4644,N_4536);
nor U6667 (N_6667,N_4504,N_1629);
or U6668 (N_6668,N_2164,N_3701);
or U6669 (N_6669,N_2055,N_1381);
nand U6670 (N_6670,N_112,N_2226);
nor U6671 (N_6671,N_4602,N_757);
or U6672 (N_6672,N_1332,N_3741);
or U6673 (N_6673,N_371,N_2014);
nand U6674 (N_6674,N_4988,N_3217);
xor U6675 (N_6675,N_1282,N_2116);
nor U6676 (N_6676,N_2223,N_962);
xnor U6677 (N_6677,N_3067,N_4100);
nand U6678 (N_6678,N_2890,N_3479);
and U6679 (N_6679,N_1000,N_2108);
nand U6680 (N_6680,N_34,N_2346);
nand U6681 (N_6681,N_4356,N_2622);
or U6682 (N_6682,N_438,N_801);
or U6683 (N_6683,N_4820,N_3203);
and U6684 (N_6684,N_3470,N_2404);
and U6685 (N_6685,N_366,N_4393);
xnor U6686 (N_6686,N_4293,N_1857);
and U6687 (N_6687,N_3547,N_4457);
and U6688 (N_6688,N_4004,N_3659);
nor U6689 (N_6689,N_3687,N_4958);
and U6690 (N_6690,N_1760,N_3253);
or U6691 (N_6691,N_4977,N_2879);
xor U6692 (N_6692,N_3888,N_3917);
or U6693 (N_6693,N_4284,N_81);
and U6694 (N_6694,N_2350,N_2757);
nor U6695 (N_6695,N_4895,N_75);
and U6696 (N_6696,N_3409,N_1063);
and U6697 (N_6697,N_1508,N_1730);
or U6698 (N_6698,N_571,N_1640);
and U6699 (N_6699,N_83,N_4273);
and U6700 (N_6700,N_3012,N_4942);
nor U6701 (N_6701,N_1598,N_4711);
and U6702 (N_6702,N_838,N_2812);
xor U6703 (N_6703,N_952,N_2864);
and U6704 (N_6704,N_595,N_3733);
nand U6705 (N_6705,N_1675,N_3101);
or U6706 (N_6706,N_4655,N_4310);
nand U6707 (N_6707,N_3239,N_3811);
or U6708 (N_6708,N_3283,N_2369);
nor U6709 (N_6709,N_479,N_3629);
nor U6710 (N_6710,N_1842,N_459);
or U6711 (N_6711,N_4553,N_4547);
and U6712 (N_6712,N_2676,N_1941);
and U6713 (N_6713,N_1995,N_2206);
nand U6714 (N_6714,N_1333,N_3465);
and U6715 (N_6715,N_4752,N_2212);
or U6716 (N_6716,N_4517,N_1732);
xnor U6717 (N_6717,N_4603,N_4649);
and U6718 (N_6718,N_2529,N_3909);
and U6719 (N_6719,N_1912,N_2234);
nor U6720 (N_6720,N_2457,N_2309);
or U6721 (N_6721,N_4624,N_3593);
or U6722 (N_6722,N_1122,N_4076);
and U6723 (N_6723,N_4101,N_108);
and U6724 (N_6724,N_3939,N_3565);
nand U6725 (N_6725,N_3642,N_1739);
and U6726 (N_6726,N_764,N_4160);
or U6727 (N_6727,N_967,N_1742);
nand U6728 (N_6728,N_1637,N_628);
xnor U6729 (N_6729,N_114,N_1180);
nand U6730 (N_6730,N_2682,N_341);
nand U6731 (N_6731,N_2728,N_3778);
and U6732 (N_6732,N_3515,N_4375);
nor U6733 (N_6733,N_4654,N_315);
and U6734 (N_6734,N_2894,N_88);
and U6735 (N_6735,N_57,N_1157);
or U6736 (N_6736,N_4680,N_1813);
nor U6737 (N_6737,N_4338,N_3962);
xor U6738 (N_6738,N_76,N_1944);
nor U6739 (N_6739,N_174,N_3242);
nor U6740 (N_6740,N_2713,N_1686);
nor U6741 (N_6741,N_790,N_4526);
nand U6742 (N_6742,N_3969,N_2194);
or U6743 (N_6743,N_1607,N_1548);
and U6744 (N_6744,N_3098,N_2769);
or U6745 (N_6745,N_4150,N_2664);
or U6746 (N_6746,N_2010,N_2217);
nor U6747 (N_6747,N_523,N_1529);
and U6748 (N_6748,N_1909,N_2482);
and U6749 (N_6749,N_2582,N_2842);
and U6750 (N_6750,N_3335,N_4112);
and U6751 (N_6751,N_4670,N_2059);
nand U6752 (N_6752,N_1452,N_934);
nor U6753 (N_6753,N_2372,N_4409);
and U6754 (N_6754,N_2152,N_761);
or U6755 (N_6755,N_680,N_1225);
or U6756 (N_6756,N_2462,N_3816);
and U6757 (N_6757,N_2903,N_2612);
or U6758 (N_6758,N_1057,N_2785);
nand U6759 (N_6759,N_194,N_2902);
nor U6760 (N_6760,N_955,N_3032);
nor U6761 (N_6761,N_1315,N_3334);
or U6762 (N_6762,N_603,N_2592);
or U6763 (N_6763,N_4968,N_485);
and U6764 (N_6764,N_2159,N_1678);
nor U6765 (N_6765,N_3634,N_1624);
and U6766 (N_6766,N_426,N_3043);
or U6767 (N_6767,N_857,N_3204);
nand U6768 (N_6768,N_3656,N_2688);
xor U6769 (N_6769,N_1577,N_471);
or U6770 (N_6770,N_1226,N_1451);
nor U6771 (N_6771,N_2876,N_4021);
and U6772 (N_6772,N_3623,N_4372);
nor U6773 (N_6773,N_4583,N_3058);
xor U6774 (N_6774,N_1547,N_3251);
nand U6775 (N_6775,N_2073,N_153);
nand U6776 (N_6776,N_4067,N_358);
and U6777 (N_6777,N_2280,N_157);
nor U6778 (N_6778,N_2208,N_2305);
or U6779 (N_6779,N_3271,N_3639);
nand U6780 (N_6780,N_1894,N_1679);
and U6781 (N_6781,N_867,N_953);
nor U6782 (N_6782,N_885,N_1443);
or U6783 (N_6783,N_1292,N_3935);
nand U6784 (N_6784,N_516,N_794);
and U6785 (N_6785,N_2111,N_3020);
and U6786 (N_6786,N_4431,N_3665);
nand U6787 (N_6787,N_1794,N_3357);
nor U6788 (N_6788,N_2027,N_4206);
nor U6789 (N_6789,N_563,N_4339);
nand U6790 (N_6790,N_3693,N_2173);
xnor U6791 (N_6791,N_328,N_1919);
and U6792 (N_6792,N_4710,N_2970);
or U6793 (N_6793,N_1911,N_1302);
and U6794 (N_6794,N_2746,N_2907);
or U6795 (N_6795,N_2563,N_4361);
or U6796 (N_6796,N_4972,N_2585);
nor U6797 (N_6797,N_2344,N_3618);
nand U6798 (N_6798,N_4465,N_1018);
xor U6799 (N_6799,N_2132,N_3413);
nor U6800 (N_6800,N_3015,N_3549);
nor U6801 (N_6801,N_2480,N_4587);
nand U6802 (N_6802,N_4537,N_1208);
or U6803 (N_6803,N_1351,N_3751);
nor U6804 (N_6804,N_833,N_2375);
and U6805 (N_6805,N_932,N_4789);
and U6806 (N_6806,N_3326,N_2338);
nor U6807 (N_6807,N_1432,N_2157);
xor U6808 (N_6808,N_504,N_532);
nor U6809 (N_6809,N_660,N_27);
and U6810 (N_6810,N_2329,N_1727);
nor U6811 (N_6811,N_3076,N_3298);
nor U6812 (N_6812,N_773,N_4161);
or U6813 (N_6813,N_4029,N_1527);
xor U6814 (N_6814,N_4838,N_4358);
or U6815 (N_6815,N_1251,N_3583);
nand U6816 (N_6816,N_4542,N_550);
or U6817 (N_6817,N_19,N_873);
nand U6818 (N_6818,N_1307,N_2534);
and U6819 (N_6819,N_2948,N_2072);
nor U6820 (N_6820,N_301,N_2272);
xor U6821 (N_6821,N_4814,N_1082);
nor U6822 (N_6822,N_238,N_53);
nand U6823 (N_6823,N_3924,N_79);
nand U6824 (N_6824,N_517,N_3489);
or U6825 (N_6825,N_62,N_691);
or U6826 (N_6826,N_758,N_2002);
nor U6827 (N_6827,N_524,N_1213);
nand U6828 (N_6828,N_80,N_1117);
and U6829 (N_6829,N_1386,N_4835);
and U6830 (N_6830,N_3995,N_3858);
nand U6831 (N_6831,N_1555,N_2517);
and U6832 (N_6832,N_3187,N_2832);
nor U6833 (N_6833,N_2930,N_3936);
and U6834 (N_6834,N_3730,N_4056);
or U6835 (N_6835,N_1861,N_4205);
nand U6836 (N_6836,N_2987,N_1303);
nor U6837 (N_6837,N_614,N_4362);
xor U6838 (N_6838,N_4514,N_2460);
and U6839 (N_6839,N_195,N_3287);
and U6840 (N_6840,N_4291,N_3146);
nand U6841 (N_6841,N_2167,N_325);
nand U6842 (N_6842,N_3937,N_1133);
nand U6843 (N_6843,N_4448,N_3352);
or U6844 (N_6844,N_1873,N_3691);
nor U6845 (N_6845,N_3402,N_3991);
and U6846 (N_6846,N_142,N_2007);
nand U6847 (N_6847,N_1056,N_4600);
nor U6848 (N_6848,N_3540,N_480);
or U6849 (N_6849,N_4414,N_1991);
nor U6850 (N_6850,N_1635,N_40);
nand U6851 (N_6851,N_2775,N_999);
nor U6852 (N_6852,N_1518,N_753);
nand U6853 (N_6853,N_3964,N_4037);
nand U6854 (N_6854,N_2411,N_4126);
nor U6855 (N_6855,N_282,N_4690);
or U6856 (N_6856,N_4468,N_2006);
and U6857 (N_6857,N_2030,N_3584);
xnor U6858 (N_6858,N_3385,N_4908);
and U6859 (N_6859,N_1458,N_1833);
nand U6860 (N_6860,N_4171,N_2588);
or U6861 (N_6861,N_4073,N_1690);
nor U6862 (N_6862,N_2012,N_3126);
and U6863 (N_6863,N_986,N_4009);
or U6864 (N_6864,N_2358,N_1943);
nor U6865 (N_6865,N_1848,N_4061);
or U6866 (N_6866,N_1494,N_3666);
and U6867 (N_6867,N_3039,N_4477);
xnor U6868 (N_6868,N_1107,N_2782);
and U6869 (N_6869,N_1281,N_4490);
nand U6870 (N_6870,N_4625,N_4801);
nand U6871 (N_6871,N_1883,N_940);
nand U6872 (N_6872,N_690,N_168);
nor U6873 (N_6873,N_799,N_1901);
or U6874 (N_6874,N_4245,N_4948);
or U6875 (N_6875,N_400,N_3569);
or U6876 (N_6876,N_592,N_4901);
nand U6877 (N_6877,N_1318,N_424);
and U6878 (N_6878,N_987,N_1085);
xnor U6879 (N_6879,N_1971,N_1992);
and U6880 (N_6880,N_372,N_478);
or U6881 (N_6881,N_1341,N_818);
or U6882 (N_6882,N_508,N_1449);
xor U6883 (N_6883,N_1973,N_1784);
and U6884 (N_6884,N_86,N_1688);
nor U6885 (N_6885,N_4412,N_2039);
and U6886 (N_6886,N_637,N_927);
nand U6887 (N_6887,N_3933,N_1563);
nand U6888 (N_6888,N_4817,N_3197);
xor U6889 (N_6889,N_739,N_3321);
nor U6890 (N_6890,N_1377,N_709);
nor U6891 (N_6891,N_3956,N_3567);
and U6892 (N_6892,N_2619,N_3422);
nand U6893 (N_6893,N_382,N_4077);
nor U6894 (N_6894,N_990,N_3440);
xnor U6895 (N_6895,N_3293,N_3975);
and U6896 (N_6896,N_3414,N_1271);
nand U6897 (N_6897,N_4192,N_4836);
xor U6898 (N_6898,N_4662,N_2617);
nor U6899 (N_6899,N_2952,N_4280);
nand U6900 (N_6900,N_3929,N_59);
or U6901 (N_6901,N_4402,N_602);
nor U6902 (N_6902,N_4277,N_685);
or U6903 (N_6903,N_556,N_1534);
and U6904 (N_6904,N_456,N_3927);
or U6905 (N_6905,N_3341,N_2129);
nand U6906 (N_6906,N_268,N_131);
nor U6907 (N_6907,N_598,N_1080);
nand U6908 (N_6908,N_3210,N_4137);
nor U6909 (N_6909,N_946,N_2646);
or U6910 (N_6910,N_995,N_1483);
or U6911 (N_6911,N_3664,N_4944);
nor U6912 (N_6912,N_727,N_1330);
or U6913 (N_6913,N_4815,N_3904);
or U6914 (N_6914,N_1699,N_1985);
and U6915 (N_6915,N_2219,N_4828);
xnor U6916 (N_6916,N_1751,N_1098);
xor U6917 (N_6917,N_1433,N_2791);
and U6918 (N_6918,N_549,N_3198);
or U6919 (N_6919,N_2446,N_2099);
nor U6920 (N_6920,N_1524,N_2794);
xor U6921 (N_6921,N_3625,N_922);
or U6922 (N_6922,N_1047,N_179);
or U6923 (N_6923,N_4274,N_1244);
xor U6924 (N_6924,N_1949,N_4749);
nand U6925 (N_6925,N_2828,N_2978);
nand U6926 (N_6926,N_1211,N_4011);
nor U6927 (N_6927,N_39,N_4096);
nand U6928 (N_6928,N_1762,N_4014);
and U6929 (N_6929,N_1145,N_3967);
nor U6930 (N_6930,N_1644,N_4323);
and U6931 (N_6931,N_2566,N_3025);
nand U6932 (N_6932,N_3944,N_4045);
nand U6933 (N_6933,N_1184,N_1545);
nor U6934 (N_6934,N_820,N_1338);
or U6935 (N_6935,N_1176,N_730);
or U6936 (N_6936,N_3417,N_4123);
nand U6937 (N_6937,N_2554,N_3533);
and U6938 (N_6938,N_207,N_2670);
nor U6939 (N_6939,N_2781,N_292);
nor U6940 (N_6940,N_3531,N_401);
nand U6941 (N_6941,N_4337,N_354);
nor U6942 (N_6942,N_3911,N_2973);
or U6943 (N_6943,N_3898,N_3328);
and U6944 (N_6944,N_3821,N_266);
or U6945 (N_6945,N_4529,N_1110);
or U6946 (N_6946,N_318,N_1324);
nor U6947 (N_6947,N_675,N_3662);
nor U6948 (N_6948,N_417,N_4111);
and U6949 (N_6949,N_427,N_1731);
nand U6950 (N_6950,N_4151,N_4259);
and U6951 (N_6951,N_1438,N_3804);
nand U6952 (N_6952,N_1054,N_3493);
and U6953 (N_6953,N_2933,N_2502);
nand U6954 (N_6954,N_3106,N_3013);
and U6955 (N_6955,N_2356,N_2492);
nand U6956 (N_6956,N_385,N_4498);
and U6957 (N_6957,N_4492,N_1683);
nand U6958 (N_6958,N_2096,N_2378);
nand U6959 (N_6959,N_4127,N_3400);
or U6960 (N_6960,N_4332,N_1037);
or U6961 (N_6961,N_945,N_4758);
and U6962 (N_6962,N_3819,N_4106);
or U6963 (N_6963,N_1498,N_3371);
and U6964 (N_6964,N_406,N_3795);
or U6965 (N_6965,N_3303,N_4062);
or U6966 (N_6966,N_3282,N_240);
and U6967 (N_6967,N_3571,N_4683);
xnor U6968 (N_6968,N_1147,N_1972);
nor U6969 (N_6969,N_3955,N_206);
or U6970 (N_6970,N_574,N_3699);
xor U6971 (N_6971,N_1819,N_791);
nor U6972 (N_6972,N_770,N_1397);
nand U6973 (N_6973,N_1620,N_4233);
or U6974 (N_6974,N_2180,N_3698);
xor U6975 (N_6975,N_2382,N_100);
and U6976 (N_6976,N_1817,N_4978);
nand U6977 (N_6977,N_3301,N_1436);
xnor U6978 (N_6978,N_1814,N_2475);
nor U6979 (N_6979,N_3375,N_3605);
or U6980 (N_6980,N_2597,N_2648);
or U6981 (N_6981,N_3431,N_2996);
or U6982 (N_6982,N_1310,N_4058);
nor U6983 (N_6983,N_2512,N_4620);
nand U6984 (N_6984,N_3925,N_865);
or U6985 (N_6985,N_2467,N_2774);
and U6986 (N_6986,N_1851,N_1257);
nand U6987 (N_6987,N_916,N_1935);
nand U6988 (N_6988,N_4519,N_1367);
nor U6989 (N_6989,N_1135,N_4181);
and U6990 (N_6990,N_3878,N_4240);
xor U6991 (N_6991,N_2506,N_2553);
and U6992 (N_6992,N_2295,N_2406);
nor U6993 (N_6993,N_1265,N_4754);
nand U6994 (N_6994,N_481,N_4166);
or U6995 (N_6995,N_1020,N_1960);
nor U6996 (N_6996,N_10,N_694);
xnor U6997 (N_6997,N_488,N_1847);
and U6998 (N_6998,N_2391,N_615);
nor U6999 (N_6999,N_4962,N_45);
nand U7000 (N_7000,N_4401,N_1561);
xnor U7001 (N_7001,N_2409,N_177);
and U7002 (N_7002,N_4424,N_2009);
nand U7003 (N_7003,N_3679,N_812);
xnor U7004 (N_7004,N_1039,N_43);
or U7005 (N_7005,N_3854,N_4398);
and U7006 (N_7006,N_13,N_3543);
nand U7007 (N_7007,N_464,N_725);
or U7008 (N_7008,N_4462,N_1975);
nand U7009 (N_7009,N_1594,N_4630);
or U7010 (N_7010,N_3218,N_4691);
or U7011 (N_7011,N_46,N_3114);
nor U7012 (N_7012,N_3749,N_2053);
and U7013 (N_7013,N_4281,N_4538);
nor U7014 (N_7014,N_3433,N_1240);
nor U7015 (N_7015,N_2896,N_908);
and U7016 (N_7016,N_1787,N_4345);
nor U7017 (N_7017,N_2044,N_543);
or U7018 (N_7018,N_1401,N_4470);
or U7019 (N_7019,N_493,N_1172);
nand U7020 (N_7020,N_4104,N_844);
or U7021 (N_7021,N_3718,N_102);
nor U7022 (N_7022,N_2805,N_275);
nand U7023 (N_7023,N_4592,N_69);
nand U7024 (N_7024,N_383,N_3144);
and U7025 (N_7025,N_3512,N_914);
or U7026 (N_7026,N_2748,N_4945);
nand U7027 (N_7027,N_1140,N_4070);
nand U7028 (N_7028,N_4685,N_2045);
or U7029 (N_7029,N_2137,N_2536);
nor U7030 (N_7030,N_877,N_2861);
nand U7031 (N_7031,N_1409,N_2979);
nor U7032 (N_7032,N_3113,N_1692);
nor U7033 (N_7033,N_487,N_3288);
and U7034 (N_7034,N_118,N_495);
nor U7035 (N_7035,N_1698,N_1936);
or U7036 (N_7036,N_3776,N_3405);
nor U7037 (N_7037,N_1022,N_3458);
nand U7038 (N_7038,N_3391,N_1761);
and U7039 (N_7039,N_3159,N_4320);
nand U7040 (N_7040,N_3495,N_1150);
xnor U7041 (N_7041,N_3460,N_3723);
xor U7042 (N_7042,N_1370,N_3832);
nand U7043 (N_7043,N_3503,N_1799);
or U7044 (N_7044,N_56,N_3449);
nand U7045 (N_7045,N_1395,N_4285);
or U7046 (N_7046,N_4717,N_3590);
nand U7047 (N_7047,N_4876,N_2736);
nand U7048 (N_7048,N_720,N_670);
nor U7049 (N_7049,N_2725,N_2110);
or U7050 (N_7050,N_2720,N_2472);
xor U7051 (N_7051,N_2722,N_2085);
nand U7052 (N_7052,N_6,N_4054);
nand U7053 (N_7053,N_2947,N_4317);
nor U7054 (N_7054,N_4724,N_450);
and U7055 (N_7055,N_3905,N_4678);
nor U7056 (N_7056,N_2024,N_2117);
nor U7057 (N_7057,N_4272,N_2972);
nand U7058 (N_7058,N_3932,N_4130);
and U7059 (N_7059,N_4974,N_1830);
and U7060 (N_7060,N_25,N_552);
and U7061 (N_7061,N_4466,N_4102);
and U7062 (N_7062,N_4289,N_3528);
nand U7063 (N_7063,N_1866,N_2684);
nand U7064 (N_7064,N_230,N_1431);
nand U7065 (N_7065,N_604,N_4267);
nor U7066 (N_7066,N_2013,N_3368);
or U7067 (N_7067,N_1890,N_991);
xor U7068 (N_7068,N_864,N_44);
and U7069 (N_7069,N_2092,N_4736);
or U7070 (N_7070,N_3885,N_3950);
nand U7071 (N_7071,N_3059,N_3729);
nor U7072 (N_7072,N_501,N_4957);
nor U7073 (N_7073,N_2000,N_3630);
and U7074 (N_7074,N_2106,N_3338);
xor U7075 (N_7075,N_2250,N_3500);
nand U7076 (N_7076,N_496,N_3576);
or U7077 (N_7077,N_2570,N_3542);
or U7078 (N_7078,N_636,N_1118);
nor U7079 (N_7079,N_2474,N_775);
nand U7080 (N_7080,N_1193,N_1167);
or U7081 (N_7081,N_182,N_683);
or U7082 (N_7082,N_4450,N_939);
or U7083 (N_7083,N_329,N_2921);
nand U7084 (N_7084,N_3611,N_1285);
xnor U7085 (N_7085,N_1323,N_2449);
and U7086 (N_7086,N_1571,N_1818);
and U7087 (N_7087,N_1177,N_4000);
xnor U7088 (N_7088,N_2589,N_2763);
and U7089 (N_7089,N_2401,N_1028);
nor U7090 (N_7090,N_219,N_2599);
or U7091 (N_7091,N_2015,N_3895);
nand U7092 (N_7092,N_4050,N_3550);
nand U7093 (N_7093,N_2331,N_4024);
nor U7094 (N_7094,N_1429,N_462);
nand U7095 (N_7095,N_242,N_1049);
nand U7096 (N_7096,N_2891,N_2297);
or U7097 (N_7097,N_3777,N_3999);
or U7098 (N_7098,N_278,N_2089);
and U7099 (N_7099,N_2416,N_3591);
nor U7100 (N_7100,N_4933,N_2082);
xnor U7101 (N_7101,N_1113,N_1532);
and U7102 (N_7102,N_2426,N_2848);
and U7103 (N_7103,N_830,N_4743);
or U7104 (N_7104,N_3390,N_3317);
nor U7105 (N_7105,N_2485,N_2195);
or U7106 (N_7106,N_4986,N_843);
or U7107 (N_7107,N_2577,N_3411);
or U7108 (N_7108,N_416,N_4841);
xnor U7109 (N_7109,N_3139,N_2384);
nor U7110 (N_7110,N_3892,N_4952);
nand U7111 (N_7111,N_2831,N_442);
and U7112 (N_7112,N_4548,N_381);
xnor U7113 (N_7113,N_4507,N_1736);
and U7114 (N_7114,N_1929,N_4157);
nor U7115 (N_7115,N_3801,N_3443);
xnor U7116 (N_7116,N_4379,N_158);
or U7117 (N_7117,N_1979,N_2837);
and U7118 (N_7118,N_3799,N_2199);
nand U7119 (N_7119,N_2450,N_3887);
and U7120 (N_7120,N_2565,N_1448);
nand U7121 (N_7121,N_2650,N_431);
nand U7122 (N_7122,N_285,N_2239);
nor U7123 (N_7123,N_4474,N_840);
and U7124 (N_7124,N_1097,N_4540);
nand U7125 (N_7125,N_1628,N_3529);
nand U7126 (N_7126,N_1077,N_4033);
xnor U7127 (N_7127,N_1930,N_4787);
or U7128 (N_7128,N_947,N_2487);
or U7129 (N_7129,N_3153,N_2425);
and U7130 (N_7130,N_3740,N_20);
xor U7131 (N_7131,N_713,N_2158);
and U7132 (N_7132,N_3874,N_3236);
nand U7133 (N_7133,N_2765,N_4695);
or U7134 (N_7134,N_1970,N_1859);
nor U7135 (N_7135,N_4886,N_2339);
and U7136 (N_7136,N_2496,N_1052);
or U7137 (N_7137,N_4563,N_4191);
or U7138 (N_7138,N_2544,N_2020);
and U7139 (N_7139,N_2968,N_1560);
or U7140 (N_7140,N_1010,N_2602);
and U7141 (N_7141,N_484,N_226);
nand U7142 (N_7142,N_1913,N_3764);
or U7143 (N_7143,N_3558,N_498);
nor U7144 (N_7144,N_2899,N_2365);
nor U7145 (N_7145,N_2564,N_1484);
xnor U7146 (N_7146,N_1268,N_1610);
nor U7147 (N_7147,N_3986,N_1);
nand U7148 (N_7148,N_2556,N_4852);
nand U7149 (N_7149,N_1950,N_186);
nor U7150 (N_7150,N_941,N_3408);
and U7151 (N_7151,N_287,N_4912);
nor U7152 (N_7152,N_807,N_2088);
nor U7153 (N_7153,N_3224,N_3622);
nand U7154 (N_7154,N_3346,N_2274);
and U7155 (N_7155,N_3175,N_3366);
and U7156 (N_7156,N_765,N_4141);
and U7157 (N_7157,N_3632,N_1967);
nand U7158 (N_7158,N_2364,N_707);
or U7159 (N_7159,N_1482,N_1881);
nor U7160 (N_7160,N_4091,N_1687);
or U7161 (N_7161,N_4399,N_4049);
nand U7162 (N_7162,N_3688,N_4299);
and U7163 (N_7163,N_1322,N_1959);
or U7164 (N_7164,N_1796,N_4175);
nand U7165 (N_7165,N_1510,N_1849);
and U7166 (N_7166,N_723,N_3392);
or U7167 (N_7167,N_4813,N_3692);
xnor U7168 (N_7168,N_314,N_2312);
nor U7169 (N_7169,N_3907,N_2969);
nor U7170 (N_7170,N_1774,N_1043);
nor U7171 (N_7171,N_1252,N_4985);
or U7172 (N_7172,N_1827,N_489);
and U7173 (N_7173,N_2017,N_891);
xnor U7174 (N_7174,N_634,N_977);
and U7175 (N_7175,N_4266,N_4265);
nor U7176 (N_7176,N_850,N_4550);
xnor U7177 (N_7177,N_2433,N_1822);
and U7178 (N_7178,N_3054,N_3333);
nor U7179 (N_7179,N_4125,N_146);
or U7180 (N_7180,N_4302,N_4410);
and U7181 (N_7181,N_107,N_1321);
nor U7182 (N_7182,N_3456,N_2253);
and U7183 (N_7183,N_2875,N_2824);
or U7184 (N_7184,N_4341,N_3915);
nor U7185 (N_7185,N_3864,N_1362);
nor U7186 (N_7186,N_948,N_307);
nand U7187 (N_7187,N_3216,N_2989);
xnor U7188 (N_7188,N_3725,N_2786);
and U7189 (N_7189,N_2174,N_4252);
nand U7190 (N_7190,N_3697,N_924);
or U7191 (N_7191,N_4871,N_4146);
or U7192 (N_7192,N_1009,N_2166);
or U7193 (N_7193,N_1406,N_2929);
or U7194 (N_7194,N_3143,N_181);
nand U7195 (N_7195,N_2809,N_2912);
and U7196 (N_7196,N_3264,N_42);
or U7197 (N_7197,N_677,N_3633);
nand U7198 (N_7198,N_4543,N_4909);
nor U7199 (N_7199,N_3348,N_1136);
nor U7200 (N_7200,N_4296,N_1229);
nand U7201 (N_7201,N_2038,N_1026);
xor U7202 (N_7202,N_4950,N_233);
nand U7203 (N_7203,N_3036,N_889);
nor U7204 (N_7204,N_767,N_2957);
or U7205 (N_7205,N_806,N_572);
nor U7206 (N_7206,N_4640,N_1957);
or U7207 (N_7207,N_2963,N_1539);
or U7208 (N_7208,N_1870,N_1215);
xor U7209 (N_7209,N_1128,N_2742);
or U7210 (N_7210,N_1142,N_1924);
nand U7211 (N_7211,N_1983,N_247);
nor U7212 (N_7212,N_2184,N_4673);
or U7213 (N_7213,N_2168,N_3064);
or U7214 (N_7214,N_3606,N_4389);
nor U7215 (N_7215,N_162,N_3430);
or U7216 (N_7216,N_2236,N_1246);
and U7217 (N_7217,N_3772,N_1259);
or U7218 (N_7218,N_534,N_1717);
or U7219 (N_7219,N_1595,N_819);
nor U7220 (N_7220,N_1865,N_1065);
or U7221 (N_7221,N_2833,N_4843);
nand U7222 (N_7222,N_4122,N_4523);
nand U7223 (N_7223,N_874,N_4036);
nand U7224 (N_7224,N_789,N_1354);
or U7225 (N_7225,N_239,N_2410);
nand U7226 (N_7226,N_1490,N_4862);
and U7227 (N_7227,N_2370,N_3724);
or U7228 (N_7228,N_1072,N_4751);
nor U7229 (N_7229,N_1540,N_3538);
nor U7230 (N_7230,N_2859,N_3788);
xnor U7231 (N_7231,N_4348,N_3026);
and U7232 (N_7232,N_703,N_2545);
nor U7233 (N_7233,N_4376,N_2273);
nor U7234 (N_7234,N_2498,N_1617);
nand U7235 (N_7235,N_3850,N_2798);
or U7236 (N_7236,N_919,N_4318);
or U7237 (N_7237,N_1293,N_3234);
nor U7238 (N_7238,N_2431,N_736);
nand U7239 (N_7239,N_2408,N_4807);
nor U7240 (N_7240,N_1003,N_2667);
nand U7241 (N_7241,N_1283,N_290);
nand U7242 (N_7242,N_2423,N_4188);
nor U7243 (N_7243,N_3676,N_2285);
xor U7244 (N_7244,N_4174,N_2271);
nor U7245 (N_7245,N_3551,N_104);
xor U7246 (N_7246,N_2041,N_804);
or U7247 (N_7247,N_3609,N_704);
nand U7248 (N_7248,N_2400,N_1479);
or U7249 (N_7249,N_4198,N_4303);
and U7250 (N_7250,N_3415,N_2373);
nor U7251 (N_7251,N_1845,N_1331);
or U7252 (N_7252,N_3318,N_4190);
nor U7253 (N_7253,N_1062,N_3517);
or U7254 (N_7254,N_3471,N_3416);
and U7255 (N_7255,N_1141,N_3738);
nor U7256 (N_7256,N_4884,N_1417);
and U7257 (N_7257,N_2094,N_4374);
xor U7258 (N_7258,N_1964,N_4740);
nor U7259 (N_7259,N_3446,N_4214);
nor U7260 (N_7260,N_1014,N_77);
or U7261 (N_7261,N_3544,N_2916);
nand U7262 (N_7262,N_1533,N_4699);
or U7263 (N_7263,N_3190,N_4496);
nand U7264 (N_7264,N_3710,N_3498);
nor U7265 (N_7265,N_1346,N_320);
nand U7266 (N_7266,N_4900,N_1345);
xnor U7267 (N_7267,N_3347,N_3564);
nand U7268 (N_7268,N_2519,N_4005);
or U7269 (N_7269,N_3896,N_3669);
xor U7270 (N_7270,N_666,N_3123);
or U7271 (N_7271,N_3115,N_389);
xor U7272 (N_7272,N_449,N_1856);
xor U7273 (N_7273,N_3831,N_3523);
nand U7274 (N_7274,N_2932,N_4262);
nor U7275 (N_7275,N_526,N_2568);
or U7276 (N_7276,N_1379,N_3397);
or U7277 (N_7277,N_3508,N_1131);
nand U7278 (N_7278,N_2469,N_2888);
xor U7279 (N_7279,N_994,N_1566);
nand U7280 (N_7280,N_513,N_1958);
xor U7281 (N_7281,N_1694,N_4002);
and U7282 (N_7282,N_2826,N_4118);
or U7283 (N_7283,N_2162,N_1643);
nor U7284 (N_7284,N_1500,N_35);
nand U7285 (N_7285,N_738,N_2518);
nor U7286 (N_7286,N_2840,N_4935);
or U7287 (N_7287,N_835,N_1258);
nor U7288 (N_7288,N_2653,N_4089);
or U7289 (N_7289,N_2711,N_728);
and U7290 (N_7290,N_3985,N_870);
or U7291 (N_7291,N_4495,N_2524);
and U7292 (N_7292,N_1669,N_3181);
xor U7293 (N_7293,N_589,N_4614);
nand U7294 (N_7294,N_2119,N_299);
nor U7295 (N_7295,N_208,N_1437);
xor U7296 (N_7296,N_696,N_1485);
nand U7297 (N_7297,N_1228,N_1114);
xnor U7298 (N_7298,N_3004,N_743);
nand U7299 (N_7299,N_3083,N_1041);
or U7300 (N_7300,N_4687,N_90);
and U7301 (N_7301,N_1816,N_1871);
and U7302 (N_7302,N_2949,N_4771);
and U7303 (N_7303,N_884,N_3327);
and U7304 (N_7304,N_557,N_2628);
and U7305 (N_7305,N_3389,N_1744);
nand U7306 (N_7306,N_4847,N_4419);
or U7307 (N_7307,N_1115,N_2647);
or U7308 (N_7308,N_2865,N_1295);
xor U7309 (N_7309,N_3053,N_3097);
or U7310 (N_7310,N_805,N_2102);
and U7311 (N_7311,N_4727,N_880);
nand U7312 (N_7312,N_1017,N_1320);
nand U7313 (N_7313,N_2922,N_1747);
xnor U7314 (N_7314,N_4545,N_4079);
or U7315 (N_7315,N_3745,N_1606);
or U7316 (N_7316,N_768,N_1843);
and U7317 (N_7317,N_510,N_4999);
or U7318 (N_7318,N_3594,N_4107);
nor U7319 (N_7319,N_4636,N_4449);
nor U7320 (N_7320,N_139,N_3970);
and U7321 (N_7321,N_148,N_3377);
nand U7322 (N_7322,N_3156,N_2690);
nand U7323 (N_7323,N_2549,N_1855);
nand U7324 (N_7324,N_2214,N_710);
nand U7325 (N_7325,N_3941,N_4890);
or U7326 (N_7326,N_2770,N_276);
xnor U7327 (N_7327,N_1795,N_2051);
nand U7328 (N_7328,N_4312,N_4825);
nor U7329 (N_7329,N_4370,N_4622);
nand U7330 (N_7330,N_4022,N_1869);
and U7331 (N_7331,N_2141,N_2251);
nor U7332 (N_7332,N_3920,N_2175);
nor U7333 (N_7333,N_1457,N_982);
nor U7334 (N_7334,N_4708,N_2065);
or U7335 (N_7335,N_2067,N_4226);
and U7336 (N_7336,N_2721,N_3300);
xnor U7337 (N_7337,N_4730,N_309);
nor U7338 (N_7338,N_3254,N_887);
nor U7339 (N_7339,N_1952,N_4494);
or U7340 (N_7340,N_4071,N_451);
or U7341 (N_7341,N_2287,N_3266);
nand U7342 (N_7342,N_1059,N_2198);
nand U7343 (N_7343,N_376,N_1218);
or U7344 (N_7344,N_2380,N_4255);
or U7345 (N_7345,N_3000,N_3247);
nor U7346 (N_7346,N_1384,N_2708);
or U7347 (N_7347,N_3491,N_4865);
nand U7348 (N_7348,N_3419,N_1461);
and U7349 (N_7349,N_3859,N_4287);
nand U7350 (N_7350,N_1716,N_734);
nor U7351 (N_7351,N_648,N_3362);
and U7352 (N_7352,N_985,N_3420);
and U7353 (N_7353,N_3072,N_4179);
xor U7354 (N_7354,N_1654,N_1616);
nand U7355 (N_7355,N_640,N_3771);
nor U7356 (N_7356,N_2481,N_2751);
nor U7357 (N_7357,N_4721,N_5);
or U7358 (N_7358,N_313,N_1981);
nor U7359 (N_7359,N_2776,N_3918);
or U7360 (N_7360,N_3223,N_2412);
xnor U7361 (N_7361,N_3140,N_2642);
xnor U7362 (N_7362,N_316,N_2031);
xnor U7363 (N_7363,N_3893,N_2131);
or U7364 (N_7364,N_1273,N_1217);
nand U7365 (N_7365,N_4692,N_3627);
xor U7366 (N_7366,N_778,N_3960);
xnor U7367 (N_7367,N_2327,N_4117);
or U7368 (N_7368,N_4241,N_4426);
and U7369 (N_7369,N_3796,N_596);
nand U7370 (N_7370,N_1553,N_4275);
and U7371 (N_7371,N_1359,N_4446);
or U7372 (N_7372,N_2458,N_2730);
and U7373 (N_7373,N_4128,N_1159);
nand U7374 (N_7374,N_2900,N_2211);
xor U7375 (N_7375,N_1708,N_3425);
xnor U7376 (N_7376,N_762,N_2541);
nor U7377 (N_7377,N_705,N_2608);
xnor U7378 (N_7378,N_3378,N_3757);
nor U7379 (N_7379,N_3573,N_2581);
and U7380 (N_7380,N_4134,N_4528);
nor U7381 (N_7381,N_2334,N_1286);
and U7382 (N_7382,N_3184,N_4322);
or U7383 (N_7383,N_3090,N_21);
and U7384 (N_7384,N_4885,N_621);
and U7385 (N_7385,N_2447,N_2575);
and U7386 (N_7386,N_2255,N_3607);
nand U7387 (N_7387,N_224,N_374);
nor U7388 (N_7388,N_1450,N_4857);
nand U7389 (N_7389,N_1287,N_263);
nor U7390 (N_7390,N_954,N_1693);
nor U7391 (N_7391,N_1165,N_2704);
nor U7392 (N_7392,N_1877,N_580);
nor U7393 (N_7393,N_1987,N_4442);
or U7394 (N_7394,N_2026,N_435);
nand U7395 (N_7395,N_4990,N_1143);
or U7396 (N_7396,N_2956,N_1753);
or U7397 (N_7397,N_2189,N_4297);
nand U7398 (N_7398,N_4532,N_3661);
nor U7399 (N_7399,N_1723,N_2193);
and U7400 (N_7400,N_788,N_4120);
xor U7401 (N_7401,N_3024,N_3365);
or U7402 (N_7402,N_4925,N_1076);
nor U7403 (N_7403,N_2355,N_405);
nand U7404 (N_7404,N_3227,N_1808);
and U7405 (N_7405,N_2558,N_1729);
and U7406 (N_7406,N_581,N_1001);
and U7407 (N_7407,N_3843,N_511);
xor U7408 (N_7408,N_2415,N_2286);
or U7409 (N_7409,N_1875,N_4929);
nand U7410 (N_7410,N_2491,N_123);
and U7411 (N_7411,N_1671,N_1993);
nor U7412 (N_7412,N_2438,N_3434);
nor U7413 (N_7413,N_3765,N_1777);
or U7414 (N_7414,N_1928,N_1836);
nand U7415 (N_7415,N_4964,N_111);
or U7416 (N_7416,N_4840,N_2967);
and U7417 (N_7417,N_3349,N_2591);
and U7418 (N_7418,N_1223,N_4165);
or U7419 (N_7419,N_4480,N_3151);
nand U7420 (N_7420,N_3459,N_3891);
and U7421 (N_7421,N_1416,N_4018);
nand U7422 (N_7422,N_4635,N_4352);
and U7423 (N_7423,N_2483,N_261);
and U7424 (N_7424,N_2126,N_1219);
nor U7425 (N_7425,N_3747,N_12);
xor U7426 (N_7426,N_2322,N_347);
nand U7427 (N_7427,N_2547,N_2802);
nand U7428 (N_7428,N_3426,N_3401);
and U7429 (N_7429,N_1221,N_2191);
or U7430 (N_7430,N_2332,N_4763);
nand U7431 (N_7431,N_815,N_3464);
or U7432 (N_7432,N_151,N_4184);
and U7433 (N_7433,N_1239,N_1029);
and U7434 (N_7434,N_286,N_4008);
or U7435 (N_7435,N_4443,N_1101);
or U7436 (N_7436,N_4854,N_3174);
and U7437 (N_7437,N_2982,N_1632);
or U7438 (N_7438,N_237,N_2238);
nand U7439 (N_7439,N_4373,N_2551);
or U7440 (N_7440,N_3031,N_1962);
or U7441 (N_7441,N_3063,N_655);
or U7442 (N_7442,N_2532,N_2510);
xor U7443 (N_7443,N_4314,N_662);
nor U7444 (N_7444,N_937,N_4334);
nor U7445 (N_7445,N_1480,N_4720);
or U7446 (N_7446,N_2103,N_3875);
and U7447 (N_7447,N_2283,N_3467);
and U7448 (N_7448,N_113,N_428);
nor U7449 (N_7449,N_537,N_2259);
xnor U7450 (N_7450,N_4864,N_322);
nor U7451 (N_7451,N_706,N_4527);
or U7452 (N_7452,N_1892,N_2434);
or U7453 (N_7453,N_50,N_138);
or U7454 (N_7454,N_1042,N_3373);
or U7455 (N_7455,N_2461,N_2594);
and U7456 (N_7456,N_959,N_116);
xor U7457 (N_7457,N_1994,N_4961);
xor U7458 (N_7458,N_1466,N_415);
nor U7459 (N_7459,N_3010,N_1910);
nor U7460 (N_7460,N_150,N_1725);
or U7461 (N_7461,N_2154,N_3667);
and U7462 (N_7462,N_500,N_4577);
or U7463 (N_7463,N_3882,N_3410);
and U7464 (N_7464,N_1474,N_2523);
nor U7465 (N_7465,N_2192,N_3466);
nand U7466 (N_7466,N_2516,N_2605);
nand U7467 (N_7467,N_3062,N_2282);
nand U7468 (N_7468,N_4888,N_4981);
nor U7469 (N_7469,N_4792,N_1642);
xnor U7470 (N_7470,N_2325,N_2165);
xnor U7471 (N_7471,N_1512,N_1615);
xor U7472 (N_7472,N_1880,N_3399);
nand U7473 (N_7473,N_2951,N_1093);
nand U7474 (N_7474,N_1954,N_2333);
and U7475 (N_7475,N_362,N_1471);
xor U7476 (N_7476,N_2319,N_1567);
or U7477 (N_7477,N_1714,N_3645);
and U7478 (N_7478,N_3901,N_2920);
and U7479 (N_7479,N_782,N_4694);
or U7480 (N_7480,N_4552,N_2675);
nand U7481 (N_7481,N_1951,N_2440);
and U7482 (N_7482,N_3982,N_1710);
nand U7483 (N_7483,N_4353,N_1423);
nor U7484 (N_7484,N_3518,N_3680);
and U7485 (N_7485,N_2944,N_4416);
or U7486 (N_7486,N_671,N_221);
and U7487 (N_7487,N_4194,N_2869);
or U7488 (N_7488,N_4209,N_3476);
and U7489 (N_7489,N_1187,N_3894);
nor U7490 (N_7490,N_109,N_4924);
and U7491 (N_7491,N_3314,N_3689);
nor U7492 (N_7492,N_1923,N_3840);
or U7493 (N_7493,N_3830,N_1422);
nor U7494 (N_7494,N_135,N_2290);
nand U7495 (N_7495,N_4286,N_2927);
nand U7496 (N_7496,N_4905,N_1129);
or U7497 (N_7497,N_1523,N_4666);
or U7498 (N_7498,N_2934,N_3337);
or U7499 (N_7499,N_4641,N_4650);
nand U7500 (N_7500,N_2043,N_99);
nand U7501 (N_7501,N_2280,N_4015);
nand U7502 (N_7502,N_308,N_742);
nor U7503 (N_7503,N_756,N_4592);
and U7504 (N_7504,N_1067,N_2172);
or U7505 (N_7505,N_4400,N_1774);
nor U7506 (N_7506,N_500,N_2795);
xor U7507 (N_7507,N_4167,N_4052);
or U7508 (N_7508,N_296,N_4108);
and U7509 (N_7509,N_993,N_2453);
xnor U7510 (N_7510,N_4352,N_238);
and U7511 (N_7511,N_1146,N_2355);
or U7512 (N_7512,N_629,N_3980);
or U7513 (N_7513,N_4400,N_1654);
or U7514 (N_7514,N_2591,N_272);
xor U7515 (N_7515,N_343,N_212);
and U7516 (N_7516,N_247,N_2433);
and U7517 (N_7517,N_746,N_3925);
nor U7518 (N_7518,N_2615,N_1962);
xnor U7519 (N_7519,N_389,N_408);
and U7520 (N_7520,N_4482,N_1750);
and U7521 (N_7521,N_1507,N_4208);
nand U7522 (N_7522,N_4517,N_4387);
or U7523 (N_7523,N_2418,N_2277);
and U7524 (N_7524,N_1247,N_3769);
nor U7525 (N_7525,N_1677,N_2664);
nor U7526 (N_7526,N_3943,N_2254);
nand U7527 (N_7527,N_3025,N_858);
nand U7528 (N_7528,N_3026,N_4291);
nor U7529 (N_7529,N_4670,N_1939);
nor U7530 (N_7530,N_1603,N_4466);
nor U7531 (N_7531,N_4988,N_4016);
or U7532 (N_7532,N_3323,N_992);
or U7533 (N_7533,N_70,N_1456);
xor U7534 (N_7534,N_1637,N_4204);
nor U7535 (N_7535,N_2047,N_1827);
or U7536 (N_7536,N_3969,N_718);
nor U7537 (N_7537,N_4629,N_253);
and U7538 (N_7538,N_2353,N_2306);
and U7539 (N_7539,N_2217,N_464);
xor U7540 (N_7540,N_160,N_1276);
and U7541 (N_7541,N_3690,N_1279);
or U7542 (N_7542,N_326,N_2570);
and U7543 (N_7543,N_3881,N_2043);
nor U7544 (N_7544,N_786,N_2471);
or U7545 (N_7545,N_65,N_4420);
nor U7546 (N_7546,N_23,N_3679);
or U7547 (N_7547,N_1181,N_2548);
or U7548 (N_7548,N_3663,N_1699);
or U7549 (N_7549,N_3489,N_180);
nor U7550 (N_7550,N_2748,N_43);
or U7551 (N_7551,N_2717,N_2280);
or U7552 (N_7552,N_4888,N_1770);
nor U7553 (N_7553,N_2371,N_3376);
xor U7554 (N_7554,N_246,N_916);
and U7555 (N_7555,N_4047,N_3785);
xor U7556 (N_7556,N_680,N_647);
nand U7557 (N_7557,N_2344,N_4579);
nor U7558 (N_7558,N_679,N_3017);
and U7559 (N_7559,N_136,N_1338);
nand U7560 (N_7560,N_1261,N_3971);
xnor U7561 (N_7561,N_4345,N_2062);
nand U7562 (N_7562,N_2524,N_1214);
nand U7563 (N_7563,N_212,N_823);
nand U7564 (N_7564,N_2562,N_3743);
or U7565 (N_7565,N_3558,N_3038);
nor U7566 (N_7566,N_4163,N_283);
nor U7567 (N_7567,N_269,N_4827);
or U7568 (N_7568,N_1241,N_2548);
or U7569 (N_7569,N_1197,N_2728);
or U7570 (N_7570,N_3539,N_2009);
nand U7571 (N_7571,N_3035,N_2371);
nand U7572 (N_7572,N_2385,N_3504);
and U7573 (N_7573,N_809,N_4650);
nor U7574 (N_7574,N_1581,N_4252);
xor U7575 (N_7575,N_3518,N_428);
nand U7576 (N_7576,N_22,N_1633);
nor U7577 (N_7577,N_2192,N_4324);
or U7578 (N_7578,N_3219,N_2718);
and U7579 (N_7579,N_4940,N_3712);
or U7580 (N_7580,N_4484,N_3817);
or U7581 (N_7581,N_2064,N_3897);
or U7582 (N_7582,N_1065,N_3834);
nand U7583 (N_7583,N_1691,N_3577);
and U7584 (N_7584,N_4568,N_3931);
and U7585 (N_7585,N_2833,N_1714);
and U7586 (N_7586,N_4116,N_3920);
nand U7587 (N_7587,N_654,N_4980);
nor U7588 (N_7588,N_184,N_1359);
nand U7589 (N_7589,N_521,N_4296);
and U7590 (N_7590,N_2193,N_493);
nand U7591 (N_7591,N_3025,N_1665);
nand U7592 (N_7592,N_2372,N_2301);
or U7593 (N_7593,N_239,N_2617);
nor U7594 (N_7594,N_4769,N_1524);
and U7595 (N_7595,N_2606,N_2468);
nor U7596 (N_7596,N_670,N_4344);
nor U7597 (N_7597,N_2051,N_614);
nor U7598 (N_7598,N_3031,N_4782);
and U7599 (N_7599,N_921,N_3919);
or U7600 (N_7600,N_3050,N_1788);
and U7601 (N_7601,N_711,N_4913);
xnor U7602 (N_7602,N_2794,N_2251);
nand U7603 (N_7603,N_4334,N_342);
nor U7604 (N_7604,N_1191,N_4285);
xor U7605 (N_7605,N_3269,N_4925);
nand U7606 (N_7606,N_1481,N_3293);
or U7607 (N_7607,N_4763,N_4796);
nor U7608 (N_7608,N_4187,N_4011);
nand U7609 (N_7609,N_4406,N_1466);
nor U7610 (N_7610,N_186,N_3626);
and U7611 (N_7611,N_2908,N_640);
nor U7612 (N_7612,N_3815,N_61);
xnor U7613 (N_7613,N_1282,N_2944);
or U7614 (N_7614,N_4836,N_4273);
nor U7615 (N_7615,N_937,N_360);
nand U7616 (N_7616,N_4474,N_4819);
nor U7617 (N_7617,N_2547,N_100);
nor U7618 (N_7618,N_1230,N_2664);
nor U7619 (N_7619,N_1135,N_4853);
nor U7620 (N_7620,N_3474,N_1193);
and U7621 (N_7621,N_4703,N_3561);
nand U7622 (N_7622,N_331,N_3124);
nor U7623 (N_7623,N_2995,N_964);
nand U7624 (N_7624,N_2487,N_2430);
and U7625 (N_7625,N_4867,N_4811);
or U7626 (N_7626,N_3781,N_57);
and U7627 (N_7627,N_4042,N_4364);
nor U7628 (N_7628,N_3791,N_3568);
nand U7629 (N_7629,N_3432,N_4022);
nand U7630 (N_7630,N_3331,N_3951);
nor U7631 (N_7631,N_4580,N_2278);
xor U7632 (N_7632,N_3755,N_4531);
or U7633 (N_7633,N_56,N_1763);
nand U7634 (N_7634,N_677,N_1850);
nand U7635 (N_7635,N_1595,N_4414);
or U7636 (N_7636,N_4406,N_2486);
nand U7637 (N_7637,N_4167,N_3085);
nand U7638 (N_7638,N_3865,N_2310);
nor U7639 (N_7639,N_1331,N_517);
or U7640 (N_7640,N_589,N_4339);
xor U7641 (N_7641,N_1754,N_2412);
and U7642 (N_7642,N_454,N_429);
nand U7643 (N_7643,N_1215,N_2707);
nand U7644 (N_7644,N_980,N_2269);
nand U7645 (N_7645,N_4869,N_3900);
nand U7646 (N_7646,N_3569,N_67);
xnor U7647 (N_7647,N_4735,N_1895);
and U7648 (N_7648,N_3991,N_1858);
or U7649 (N_7649,N_4046,N_1704);
or U7650 (N_7650,N_4343,N_4616);
and U7651 (N_7651,N_2463,N_4460);
nand U7652 (N_7652,N_2,N_637);
or U7653 (N_7653,N_3479,N_2938);
and U7654 (N_7654,N_211,N_2333);
nor U7655 (N_7655,N_4688,N_2372);
and U7656 (N_7656,N_3417,N_3103);
xor U7657 (N_7657,N_3006,N_1206);
or U7658 (N_7658,N_4708,N_4264);
nor U7659 (N_7659,N_4245,N_2797);
xnor U7660 (N_7660,N_2060,N_3412);
or U7661 (N_7661,N_1221,N_504);
nor U7662 (N_7662,N_1508,N_2872);
or U7663 (N_7663,N_1052,N_4131);
nor U7664 (N_7664,N_3351,N_4443);
nand U7665 (N_7665,N_1111,N_1756);
nor U7666 (N_7666,N_3520,N_2677);
nor U7667 (N_7667,N_82,N_513);
or U7668 (N_7668,N_2755,N_2104);
or U7669 (N_7669,N_3692,N_4425);
nand U7670 (N_7670,N_3707,N_2715);
and U7671 (N_7671,N_1696,N_270);
nor U7672 (N_7672,N_2821,N_1340);
nand U7673 (N_7673,N_1669,N_3532);
and U7674 (N_7674,N_2611,N_2111);
and U7675 (N_7675,N_1698,N_511);
nand U7676 (N_7676,N_1128,N_3937);
nor U7677 (N_7677,N_142,N_3518);
or U7678 (N_7678,N_3078,N_3289);
and U7679 (N_7679,N_2523,N_453);
nand U7680 (N_7680,N_4292,N_549);
nor U7681 (N_7681,N_1134,N_803);
nand U7682 (N_7682,N_1644,N_535);
or U7683 (N_7683,N_1906,N_4812);
nand U7684 (N_7684,N_3544,N_2479);
nand U7685 (N_7685,N_1653,N_3440);
nand U7686 (N_7686,N_2991,N_2603);
xor U7687 (N_7687,N_3895,N_3836);
nor U7688 (N_7688,N_1201,N_3953);
nand U7689 (N_7689,N_492,N_4782);
or U7690 (N_7690,N_4267,N_3485);
nand U7691 (N_7691,N_920,N_171);
nand U7692 (N_7692,N_4204,N_4367);
nor U7693 (N_7693,N_2021,N_3297);
and U7694 (N_7694,N_679,N_1970);
nand U7695 (N_7695,N_3135,N_877);
xnor U7696 (N_7696,N_2876,N_667);
nand U7697 (N_7697,N_4333,N_232);
nor U7698 (N_7698,N_3540,N_701);
nor U7699 (N_7699,N_3261,N_3615);
and U7700 (N_7700,N_205,N_4340);
xnor U7701 (N_7701,N_4438,N_893);
or U7702 (N_7702,N_469,N_2487);
or U7703 (N_7703,N_3735,N_4571);
xor U7704 (N_7704,N_4372,N_1785);
or U7705 (N_7705,N_4157,N_274);
nor U7706 (N_7706,N_3568,N_3095);
nand U7707 (N_7707,N_4523,N_4785);
nor U7708 (N_7708,N_65,N_4067);
nand U7709 (N_7709,N_4523,N_3381);
and U7710 (N_7710,N_3261,N_3376);
and U7711 (N_7711,N_4944,N_4645);
or U7712 (N_7712,N_3855,N_1257);
or U7713 (N_7713,N_4609,N_1255);
xnor U7714 (N_7714,N_705,N_4268);
xor U7715 (N_7715,N_2101,N_1095);
nand U7716 (N_7716,N_1659,N_1926);
nand U7717 (N_7717,N_881,N_1992);
and U7718 (N_7718,N_3585,N_3561);
or U7719 (N_7719,N_143,N_3481);
xor U7720 (N_7720,N_4518,N_733);
nand U7721 (N_7721,N_1603,N_2078);
xor U7722 (N_7722,N_4325,N_3044);
nand U7723 (N_7723,N_3966,N_4440);
nand U7724 (N_7724,N_595,N_1121);
and U7725 (N_7725,N_155,N_4847);
and U7726 (N_7726,N_2084,N_102);
or U7727 (N_7727,N_1121,N_969);
nor U7728 (N_7728,N_2037,N_487);
or U7729 (N_7729,N_1092,N_4139);
nand U7730 (N_7730,N_779,N_4533);
or U7731 (N_7731,N_1950,N_3062);
or U7732 (N_7732,N_4908,N_3497);
or U7733 (N_7733,N_2581,N_2982);
and U7734 (N_7734,N_3,N_4160);
nor U7735 (N_7735,N_4471,N_2536);
or U7736 (N_7736,N_708,N_1076);
and U7737 (N_7737,N_3300,N_71);
and U7738 (N_7738,N_4883,N_3806);
and U7739 (N_7739,N_1740,N_4487);
or U7740 (N_7740,N_2282,N_4620);
xnor U7741 (N_7741,N_925,N_1769);
and U7742 (N_7742,N_4940,N_248);
nand U7743 (N_7743,N_4662,N_1632);
nand U7744 (N_7744,N_34,N_1715);
nor U7745 (N_7745,N_4308,N_2281);
nand U7746 (N_7746,N_1852,N_1631);
xor U7747 (N_7747,N_4718,N_531);
nor U7748 (N_7748,N_1242,N_3591);
and U7749 (N_7749,N_1044,N_2495);
nor U7750 (N_7750,N_1425,N_361);
and U7751 (N_7751,N_85,N_4622);
xor U7752 (N_7752,N_311,N_2276);
and U7753 (N_7753,N_3884,N_388);
xnor U7754 (N_7754,N_3365,N_2956);
nand U7755 (N_7755,N_4033,N_2637);
nor U7756 (N_7756,N_4073,N_810);
nor U7757 (N_7757,N_2958,N_2613);
nor U7758 (N_7758,N_3813,N_1909);
nor U7759 (N_7759,N_875,N_4379);
nand U7760 (N_7760,N_2140,N_1660);
or U7761 (N_7761,N_1740,N_566);
or U7762 (N_7762,N_461,N_4580);
nand U7763 (N_7763,N_4207,N_2300);
xnor U7764 (N_7764,N_3948,N_1934);
xor U7765 (N_7765,N_1575,N_3331);
xnor U7766 (N_7766,N_2973,N_154);
and U7767 (N_7767,N_2774,N_4352);
nor U7768 (N_7768,N_347,N_3092);
xor U7769 (N_7769,N_2667,N_2474);
nor U7770 (N_7770,N_3274,N_4892);
or U7771 (N_7771,N_4104,N_1635);
or U7772 (N_7772,N_2935,N_289);
or U7773 (N_7773,N_570,N_1810);
and U7774 (N_7774,N_215,N_1135);
nand U7775 (N_7775,N_4794,N_2647);
nand U7776 (N_7776,N_2771,N_3403);
or U7777 (N_7777,N_4876,N_2239);
and U7778 (N_7778,N_4795,N_4208);
or U7779 (N_7779,N_4649,N_539);
nand U7780 (N_7780,N_2183,N_3562);
or U7781 (N_7781,N_3422,N_3319);
xor U7782 (N_7782,N_4630,N_1720);
nand U7783 (N_7783,N_2106,N_903);
nand U7784 (N_7784,N_3089,N_2374);
or U7785 (N_7785,N_2755,N_3468);
or U7786 (N_7786,N_620,N_211);
or U7787 (N_7787,N_2254,N_766);
and U7788 (N_7788,N_1372,N_2217);
nand U7789 (N_7789,N_1859,N_1353);
or U7790 (N_7790,N_3654,N_444);
and U7791 (N_7791,N_2872,N_3912);
xnor U7792 (N_7792,N_4281,N_4286);
nand U7793 (N_7793,N_1725,N_4761);
nor U7794 (N_7794,N_3216,N_2375);
nor U7795 (N_7795,N_1267,N_1491);
xor U7796 (N_7796,N_3134,N_4947);
or U7797 (N_7797,N_996,N_3178);
or U7798 (N_7798,N_2948,N_370);
and U7799 (N_7799,N_3838,N_799);
or U7800 (N_7800,N_4455,N_3870);
and U7801 (N_7801,N_2355,N_4387);
or U7802 (N_7802,N_2909,N_1630);
or U7803 (N_7803,N_894,N_1741);
nor U7804 (N_7804,N_1568,N_2565);
nand U7805 (N_7805,N_2404,N_4079);
nor U7806 (N_7806,N_1827,N_2904);
or U7807 (N_7807,N_2662,N_2896);
nor U7808 (N_7808,N_2527,N_3320);
nor U7809 (N_7809,N_234,N_1577);
nor U7810 (N_7810,N_4694,N_4451);
or U7811 (N_7811,N_4238,N_3454);
nor U7812 (N_7812,N_1117,N_3427);
xnor U7813 (N_7813,N_1681,N_826);
and U7814 (N_7814,N_4935,N_1156);
or U7815 (N_7815,N_3191,N_4352);
or U7816 (N_7816,N_3279,N_1928);
or U7817 (N_7817,N_2053,N_4899);
nor U7818 (N_7818,N_1319,N_1451);
xor U7819 (N_7819,N_577,N_255);
and U7820 (N_7820,N_4101,N_1876);
nor U7821 (N_7821,N_2919,N_820);
or U7822 (N_7822,N_3030,N_1232);
nor U7823 (N_7823,N_263,N_4905);
xnor U7824 (N_7824,N_1326,N_4312);
nor U7825 (N_7825,N_2314,N_1892);
or U7826 (N_7826,N_3682,N_1186);
xor U7827 (N_7827,N_3224,N_467);
xor U7828 (N_7828,N_2148,N_4310);
and U7829 (N_7829,N_3072,N_2120);
nor U7830 (N_7830,N_2081,N_4687);
nand U7831 (N_7831,N_3693,N_2151);
and U7832 (N_7832,N_2238,N_4039);
nor U7833 (N_7833,N_4514,N_2692);
or U7834 (N_7834,N_1613,N_783);
nand U7835 (N_7835,N_1800,N_3366);
and U7836 (N_7836,N_1092,N_3540);
xor U7837 (N_7837,N_39,N_2602);
nor U7838 (N_7838,N_1645,N_3623);
nor U7839 (N_7839,N_3974,N_680);
nand U7840 (N_7840,N_4670,N_3413);
and U7841 (N_7841,N_4920,N_3987);
and U7842 (N_7842,N_1982,N_3156);
xnor U7843 (N_7843,N_1576,N_1420);
or U7844 (N_7844,N_1326,N_648);
nor U7845 (N_7845,N_1242,N_807);
and U7846 (N_7846,N_3876,N_4877);
nor U7847 (N_7847,N_992,N_4906);
nor U7848 (N_7848,N_1663,N_2816);
and U7849 (N_7849,N_3022,N_2408);
and U7850 (N_7850,N_1651,N_1294);
or U7851 (N_7851,N_1062,N_580);
or U7852 (N_7852,N_4970,N_1633);
nand U7853 (N_7853,N_1726,N_2199);
xnor U7854 (N_7854,N_4439,N_1197);
xnor U7855 (N_7855,N_4004,N_3535);
nor U7856 (N_7856,N_1233,N_3361);
nand U7857 (N_7857,N_475,N_1501);
nor U7858 (N_7858,N_3174,N_3134);
and U7859 (N_7859,N_717,N_2941);
nor U7860 (N_7860,N_3944,N_4888);
or U7861 (N_7861,N_1290,N_2536);
nand U7862 (N_7862,N_871,N_3609);
nor U7863 (N_7863,N_4909,N_2120);
or U7864 (N_7864,N_1935,N_2303);
or U7865 (N_7865,N_3008,N_4286);
nor U7866 (N_7866,N_3951,N_2335);
or U7867 (N_7867,N_666,N_1683);
or U7868 (N_7868,N_4002,N_4657);
or U7869 (N_7869,N_2530,N_665);
nand U7870 (N_7870,N_2860,N_3733);
or U7871 (N_7871,N_3058,N_692);
or U7872 (N_7872,N_4920,N_3475);
and U7873 (N_7873,N_2629,N_1095);
xnor U7874 (N_7874,N_4262,N_2635);
nand U7875 (N_7875,N_3261,N_206);
nand U7876 (N_7876,N_271,N_1361);
or U7877 (N_7877,N_4342,N_1448);
xnor U7878 (N_7878,N_574,N_1811);
nand U7879 (N_7879,N_4670,N_2978);
and U7880 (N_7880,N_2038,N_2945);
nor U7881 (N_7881,N_4250,N_3452);
and U7882 (N_7882,N_2874,N_4630);
and U7883 (N_7883,N_2383,N_4962);
and U7884 (N_7884,N_4625,N_2186);
or U7885 (N_7885,N_4708,N_1934);
nand U7886 (N_7886,N_2636,N_3140);
nor U7887 (N_7887,N_3556,N_1815);
nand U7888 (N_7888,N_2038,N_1974);
or U7889 (N_7889,N_989,N_1594);
nand U7890 (N_7890,N_1013,N_2665);
and U7891 (N_7891,N_2552,N_1690);
and U7892 (N_7892,N_57,N_1136);
nor U7893 (N_7893,N_4014,N_4566);
and U7894 (N_7894,N_4193,N_2768);
nand U7895 (N_7895,N_3230,N_144);
nor U7896 (N_7896,N_1929,N_2797);
xnor U7897 (N_7897,N_2592,N_3297);
or U7898 (N_7898,N_306,N_10);
or U7899 (N_7899,N_1841,N_1245);
or U7900 (N_7900,N_2627,N_4928);
nor U7901 (N_7901,N_880,N_4726);
or U7902 (N_7902,N_4781,N_744);
and U7903 (N_7903,N_2403,N_2089);
or U7904 (N_7904,N_466,N_2920);
and U7905 (N_7905,N_2022,N_4214);
and U7906 (N_7906,N_2388,N_1662);
nand U7907 (N_7907,N_942,N_2465);
or U7908 (N_7908,N_3530,N_4257);
or U7909 (N_7909,N_2891,N_4772);
nand U7910 (N_7910,N_1877,N_387);
nor U7911 (N_7911,N_1094,N_2197);
nor U7912 (N_7912,N_791,N_1386);
and U7913 (N_7913,N_2503,N_4746);
xnor U7914 (N_7914,N_1505,N_4682);
nand U7915 (N_7915,N_565,N_4550);
and U7916 (N_7916,N_2448,N_3820);
or U7917 (N_7917,N_2016,N_4171);
nor U7918 (N_7918,N_1909,N_2006);
or U7919 (N_7919,N_689,N_2569);
or U7920 (N_7920,N_143,N_144);
xnor U7921 (N_7921,N_1751,N_4751);
and U7922 (N_7922,N_3835,N_2808);
nand U7923 (N_7923,N_134,N_220);
or U7924 (N_7924,N_3614,N_3527);
nor U7925 (N_7925,N_3995,N_2659);
nor U7926 (N_7926,N_2348,N_2622);
xnor U7927 (N_7927,N_895,N_1091);
nor U7928 (N_7928,N_3504,N_2568);
nand U7929 (N_7929,N_1842,N_1623);
or U7930 (N_7930,N_4317,N_4380);
nand U7931 (N_7931,N_4974,N_2083);
nor U7932 (N_7932,N_2312,N_1486);
nor U7933 (N_7933,N_532,N_3107);
and U7934 (N_7934,N_1826,N_2441);
xnor U7935 (N_7935,N_2126,N_4852);
xor U7936 (N_7936,N_3260,N_2491);
or U7937 (N_7937,N_4260,N_192);
and U7938 (N_7938,N_4488,N_3848);
and U7939 (N_7939,N_3712,N_1235);
nand U7940 (N_7940,N_3050,N_1301);
and U7941 (N_7941,N_3795,N_4415);
and U7942 (N_7942,N_2076,N_2462);
or U7943 (N_7943,N_1450,N_201);
nor U7944 (N_7944,N_1470,N_3361);
and U7945 (N_7945,N_2713,N_2491);
and U7946 (N_7946,N_3238,N_1604);
nor U7947 (N_7947,N_4474,N_4261);
and U7948 (N_7948,N_3017,N_1060);
or U7949 (N_7949,N_4591,N_2180);
and U7950 (N_7950,N_2242,N_1522);
nor U7951 (N_7951,N_3779,N_2687);
nor U7952 (N_7952,N_36,N_3696);
nor U7953 (N_7953,N_4294,N_4933);
nand U7954 (N_7954,N_565,N_465);
and U7955 (N_7955,N_4127,N_4028);
nand U7956 (N_7956,N_4545,N_2315);
nor U7957 (N_7957,N_3279,N_4595);
or U7958 (N_7958,N_3095,N_1447);
nand U7959 (N_7959,N_4166,N_2619);
or U7960 (N_7960,N_80,N_3867);
or U7961 (N_7961,N_2957,N_3826);
or U7962 (N_7962,N_4269,N_1428);
nor U7963 (N_7963,N_2557,N_2110);
nand U7964 (N_7964,N_2712,N_571);
or U7965 (N_7965,N_322,N_2442);
nor U7966 (N_7966,N_4708,N_2952);
or U7967 (N_7967,N_3540,N_3352);
nor U7968 (N_7968,N_4051,N_754);
and U7969 (N_7969,N_1666,N_4512);
nor U7970 (N_7970,N_160,N_819);
or U7971 (N_7971,N_1969,N_871);
nor U7972 (N_7972,N_2708,N_3109);
nand U7973 (N_7973,N_1064,N_3210);
or U7974 (N_7974,N_4881,N_4191);
nand U7975 (N_7975,N_4223,N_1587);
xnor U7976 (N_7976,N_3878,N_4453);
nor U7977 (N_7977,N_3635,N_2418);
nand U7978 (N_7978,N_2159,N_4612);
nor U7979 (N_7979,N_1240,N_444);
or U7980 (N_7980,N_3440,N_4930);
and U7981 (N_7981,N_1659,N_4936);
nor U7982 (N_7982,N_4345,N_97);
nor U7983 (N_7983,N_1645,N_4696);
nor U7984 (N_7984,N_4985,N_987);
and U7985 (N_7985,N_849,N_3286);
and U7986 (N_7986,N_2722,N_1384);
and U7987 (N_7987,N_4864,N_3393);
and U7988 (N_7988,N_4489,N_3508);
or U7989 (N_7989,N_4948,N_1086);
nor U7990 (N_7990,N_3375,N_3863);
nand U7991 (N_7991,N_2664,N_4813);
nand U7992 (N_7992,N_3286,N_3824);
nor U7993 (N_7993,N_4468,N_4291);
and U7994 (N_7994,N_1025,N_3028);
nor U7995 (N_7995,N_4513,N_844);
and U7996 (N_7996,N_2455,N_3534);
xnor U7997 (N_7997,N_1175,N_938);
nand U7998 (N_7998,N_2447,N_4085);
xor U7999 (N_7999,N_1862,N_2195);
or U8000 (N_8000,N_546,N_296);
nand U8001 (N_8001,N_1832,N_4824);
or U8002 (N_8002,N_2033,N_2626);
or U8003 (N_8003,N_1120,N_3752);
or U8004 (N_8004,N_2625,N_163);
xor U8005 (N_8005,N_4294,N_4512);
nor U8006 (N_8006,N_4684,N_3424);
xnor U8007 (N_8007,N_48,N_3392);
and U8008 (N_8008,N_4414,N_3912);
or U8009 (N_8009,N_4136,N_559);
nor U8010 (N_8010,N_1785,N_3720);
xor U8011 (N_8011,N_1718,N_4853);
and U8012 (N_8012,N_319,N_3228);
nor U8013 (N_8013,N_3646,N_2239);
and U8014 (N_8014,N_2589,N_4806);
nor U8015 (N_8015,N_232,N_2142);
and U8016 (N_8016,N_2909,N_4406);
nand U8017 (N_8017,N_3902,N_1760);
xor U8018 (N_8018,N_3536,N_842);
nor U8019 (N_8019,N_2575,N_1489);
nand U8020 (N_8020,N_3745,N_1172);
nand U8021 (N_8021,N_3423,N_200);
nor U8022 (N_8022,N_4665,N_2072);
nor U8023 (N_8023,N_1102,N_918);
and U8024 (N_8024,N_1789,N_588);
xnor U8025 (N_8025,N_197,N_3095);
or U8026 (N_8026,N_3802,N_4467);
and U8027 (N_8027,N_4789,N_1074);
nand U8028 (N_8028,N_4573,N_3524);
and U8029 (N_8029,N_3069,N_1177);
nand U8030 (N_8030,N_2470,N_2629);
xnor U8031 (N_8031,N_2965,N_2833);
or U8032 (N_8032,N_3043,N_179);
and U8033 (N_8033,N_2296,N_3062);
nand U8034 (N_8034,N_3676,N_604);
nor U8035 (N_8035,N_1159,N_3631);
nor U8036 (N_8036,N_113,N_4874);
nor U8037 (N_8037,N_1102,N_4278);
or U8038 (N_8038,N_4910,N_774);
nand U8039 (N_8039,N_4020,N_2457);
xnor U8040 (N_8040,N_4451,N_3613);
nor U8041 (N_8041,N_4688,N_1456);
nor U8042 (N_8042,N_269,N_1027);
nor U8043 (N_8043,N_57,N_498);
xor U8044 (N_8044,N_2099,N_698);
nand U8045 (N_8045,N_4131,N_2629);
or U8046 (N_8046,N_3250,N_2782);
or U8047 (N_8047,N_4436,N_432);
or U8048 (N_8048,N_2845,N_3135);
nand U8049 (N_8049,N_3210,N_3395);
nor U8050 (N_8050,N_234,N_3361);
or U8051 (N_8051,N_839,N_2174);
or U8052 (N_8052,N_1953,N_2279);
nand U8053 (N_8053,N_675,N_2893);
nor U8054 (N_8054,N_4528,N_4985);
nand U8055 (N_8055,N_475,N_130);
or U8056 (N_8056,N_3290,N_2050);
or U8057 (N_8057,N_3379,N_254);
nor U8058 (N_8058,N_2377,N_2704);
and U8059 (N_8059,N_1318,N_2346);
nor U8060 (N_8060,N_2114,N_466);
or U8061 (N_8061,N_2848,N_2203);
nand U8062 (N_8062,N_3680,N_1125);
nor U8063 (N_8063,N_2465,N_121);
or U8064 (N_8064,N_787,N_4284);
nand U8065 (N_8065,N_3821,N_2500);
xnor U8066 (N_8066,N_4391,N_972);
and U8067 (N_8067,N_2541,N_928);
nor U8068 (N_8068,N_182,N_881);
nand U8069 (N_8069,N_3919,N_1584);
nor U8070 (N_8070,N_1666,N_2297);
nand U8071 (N_8071,N_4517,N_919);
and U8072 (N_8072,N_1732,N_331);
or U8073 (N_8073,N_3180,N_2348);
and U8074 (N_8074,N_684,N_4879);
and U8075 (N_8075,N_823,N_2114);
nor U8076 (N_8076,N_2781,N_3829);
and U8077 (N_8077,N_3246,N_328);
and U8078 (N_8078,N_1029,N_4434);
and U8079 (N_8079,N_477,N_2055);
or U8080 (N_8080,N_4364,N_1089);
or U8081 (N_8081,N_328,N_4179);
nand U8082 (N_8082,N_3132,N_222);
or U8083 (N_8083,N_2113,N_1202);
nand U8084 (N_8084,N_4073,N_30);
nand U8085 (N_8085,N_4578,N_710);
nor U8086 (N_8086,N_3569,N_1849);
nand U8087 (N_8087,N_4643,N_2538);
nand U8088 (N_8088,N_1542,N_439);
or U8089 (N_8089,N_3062,N_1660);
or U8090 (N_8090,N_1882,N_2571);
and U8091 (N_8091,N_4999,N_1915);
and U8092 (N_8092,N_1362,N_1960);
and U8093 (N_8093,N_445,N_1327);
nor U8094 (N_8094,N_2266,N_1136);
or U8095 (N_8095,N_500,N_4790);
or U8096 (N_8096,N_3606,N_916);
nand U8097 (N_8097,N_2295,N_4563);
or U8098 (N_8098,N_3083,N_2173);
nand U8099 (N_8099,N_4776,N_4727);
and U8100 (N_8100,N_293,N_4220);
nor U8101 (N_8101,N_2515,N_138);
nor U8102 (N_8102,N_1981,N_3009);
nand U8103 (N_8103,N_3042,N_4731);
and U8104 (N_8104,N_3598,N_4319);
and U8105 (N_8105,N_3801,N_772);
nor U8106 (N_8106,N_4691,N_4611);
nor U8107 (N_8107,N_3612,N_2725);
nor U8108 (N_8108,N_2235,N_2016);
nand U8109 (N_8109,N_2892,N_2292);
or U8110 (N_8110,N_4954,N_3715);
or U8111 (N_8111,N_3416,N_2705);
nor U8112 (N_8112,N_874,N_4932);
nor U8113 (N_8113,N_461,N_1136);
or U8114 (N_8114,N_3338,N_1227);
nor U8115 (N_8115,N_123,N_3429);
and U8116 (N_8116,N_1425,N_1423);
nand U8117 (N_8117,N_2701,N_2047);
nor U8118 (N_8118,N_1097,N_4350);
nand U8119 (N_8119,N_2651,N_2646);
xor U8120 (N_8120,N_2424,N_3543);
or U8121 (N_8121,N_963,N_4036);
or U8122 (N_8122,N_1137,N_22);
nand U8123 (N_8123,N_192,N_1343);
and U8124 (N_8124,N_1667,N_1196);
xnor U8125 (N_8125,N_3189,N_2471);
nor U8126 (N_8126,N_2426,N_2729);
xor U8127 (N_8127,N_187,N_2184);
or U8128 (N_8128,N_531,N_3877);
or U8129 (N_8129,N_4725,N_3851);
xor U8130 (N_8130,N_1718,N_3508);
and U8131 (N_8131,N_4968,N_4943);
xnor U8132 (N_8132,N_617,N_4440);
nor U8133 (N_8133,N_4240,N_1966);
nor U8134 (N_8134,N_1897,N_1758);
or U8135 (N_8135,N_4561,N_2896);
or U8136 (N_8136,N_3025,N_4319);
and U8137 (N_8137,N_3676,N_1963);
or U8138 (N_8138,N_1753,N_2499);
and U8139 (N_8139,N_606,N_4669);
nor U8140 (N_8140,N_3573,N_3344);
nand U8141 (N_8141,N_1371,N_3757);
nand U8142 (N_8142,N_4778,N_725);
and U8143 (N_8143,N_2150,N_368);
and U8144 (N_8144,N_3840,N_1075);
nor U8145 (N_8145,N_4516,N_3353);
and U8146 (N_8146,N_3967,N_862);
nand U8147 (N_8147,N_2331,N_3492);
nand U8148 (N_8148,N_4543,N_3129);
xor U8149 (N_8149,N_1364,N_4284);
nand U8150 (N_8150,N_1644,N_2350);
and U8151 (N_8151,N_590,N_1965);
or U8152 (N_8152,N_1654,N_249);
nor U8153 (N_8153,N_2729,N_3847);
and U8154 (N_8154,N_3005,N_4918);
nor U8155 (N_8155,N_1624,N_4023);
and U8156 (N_8156,N_4710,N_2842);
nor U8157 (N_8157,N_3041,N_1517);
and U8158 (N_8158,N_3976,N_3337);
nand U8159 (N_8159,N_421,N_1516);
or U8160 (N_8160,N_1582,N_252);
and U8161 (N_8161,N_3736,N_865);
or U8162 (N_8162,N_1912,N_1705);
nand U8163 (N_8163,N_149,N_1486);
and U8164 (N_8164,N_3624,N_4609);
or U8165 (N_8165,N_3586,N_3264);
nand U8166 (N_8166,N_1871,N_2771);
or U8167 (N_8167,N_1425,N_4400);
or U8168 (N_8168,N_1608,N_4693);
nor U8169 (N_8169,N_1517,N_1315);
or U8170 (N_8170,N_4819,N_3530);
xnor U8171 (N_8171,N_2248,N_1410);
nor U8172 (N_8172,N_4554,N_4615);
nor U8173 (N_8173,N_2328,N_410);
or U8174 (N_8174,N_1296,N_3173);
xor U8175 (N_8175,N_720,N_4530);
xnor U8176 (N_8176,N_3965,N_49);
and U8177 (N_8177,N_4071,N_719);
nor U8178 (N_8178,N_3374,N_872);
or U8179 (N_8179,N_4171,N_3566);
or U8180 (N_8180,N_3155,N_594);
xor U8181 (N_8181,N_2630,N_4655);
or U8182 (N_8182,N_553,N_391);
and U8183 (N_8183,N_1460,N_3863);
and U8184 (N_8184,N_181,N_3567);
nand U8185 (N_8185,N_345,N_1033);
xnor U8186 (N_8186,N_3515,N_2696);
nand U8187 (N_8187,N_1720,N_262);
xor U8188 (N_8188,N_4751,N_3946);
and U8189 (N_8189,N_2760,N_1708);
nand U8190 (N_8190,N_3393,N_3125);
nand U8191 (N_8191,N_518,N_629);
xnor U8192 (N_8192,N_4908,N_251);
and U8193 (N_8193,N_4822,N_558);
nand U8194 (N_8194,N_4076,N_2459);
or U8195 (N_8195,N_2152,N_2865);
nand U8196 (N_8196,N_861,N_2521);
nor U8197 (N_8197,N_2521,N_3487);
nor U8198 (N_8198,N_4992,N_3671);
and U8199 (N_8199,N_900,N_3402);
and U8200 (N_8200,N_2080,N_2422);
nand U8201 (N_8201,N_1352,N_1131);
or U8202 (N_8202,N_3544,N_667);
nor U8203 (N_8203,N_1730,N_3388);
nor U8204 (N_8204,N_2163,N_2779);
nor U8205 (N_8205,N_4782,N_3755);
and U8206 (N_8206,N_2872,N_2642);
nor U8207 (N_8207,N_1853,N_64);
and U8208 (N_8208,N_2052,N_3566);
or U8209 (N_8209,N_3714,N_724);
or U8210 (N_8210,N_4853,N_2398);
and U8211 (N_8211,N_2753,N_4244);
nand U8212 (N_8212,N_2689,N_3556);
or U8213 (N_8213,N_324,N_3732);
or U8214 (N_8214,N_850,N_2557);
and U8215 (N_8215,N_4298,N_4873);
nor U8216 (N_8216,N_2438,N_2787);
xor U8217 (N_8217,N_1124,N_742);
xnor U8218 (N_8218,N_3187,N_2277);
nor U8219 (N_8219,N_1280,N_2668);
and U8220 (N_8220,N_2399,N_3314);
nor U8221 (N_8221,N_1180,N_4364);
nor U8222 (N_8222,N_1795,N_4448);
nor U8223 (N_8223,N_1529,N_1634);
nor U8224 (N_8224,N_410,N_232);
nor U8225 (N_8225,N_1636,N_1383);
or U8226 (N_8226,N_2891,N_3360);
or U8227 (N_8227,N_2960,N_1122);
or U8228 (N_8228,N_2987,N_2211);
nor U8229 (N_8229,N_2337,N_3029);
and U8230 (N_8230,N_3526,N_3728);
or U8231 (N_8231,N_1409,N_4095);
nand U8232 (N_8232,N_3619,N_2307);
and U8233 (N_8233,N_2422,N_4914);
nand U8234 (N_8234,N_4190,N_4183);
nor U8235 (N_8235,N_227,N_4914);
and U8236 (N_8236,N_2223,N_1082);
nand U8237 (N_8237,N_872,N_1333);
or U8238 (N_8238,N_3212,N_4222);
nand U8239 (N_8239,N_3811,N_3252);
nor U8240 (N_8240,N_350,N_2748);
or U8241 (N_8241,N_3542,N_4684);
or U8242 (N_8242,N_4983,N_3117);
nand U8243 (N_8243,N_1018,N_2622);
xnor U8244 (N_8244,N_3784,N_586);
nand U8245 (N_8245,N_2818,N_4655);
and U8246 (N_8246,N_1769,N_3842);
or U8247 (N_8247,N_1280,N_3418);
xnor U8248 (N_8248,N_2454,N_311);
or U8249 (N_8249,N_1564,N_517);
or U8250 (N_8250,N_577,N_4931);
nand U8251 (N_8251,N_1335,N_2277);
nand U8252 (N_8252,N_653,N_1867);
or U8253 (N_8253,N_4314,N_3450);
and U8254 (N_8254,N_2975,N_535);
nor U8255 (N_8255,N_301,N_3952);
nand U8256 (N_8256,N_642,N_1347);
or U8257 (N_8257,N_3125,N_2228);
nor U8258 (N_8258,N_4264,N_2724);
and U8259 (N_8259,N_4756,N_1932);
and U8260 (N_8260,N_122,N_2529);
nor U8261 (N_8261,N_4797,N_8);
xor U8262 (N_8262,N_2516,N_91);
nor U8263 (N_8263,N_3287,N_4209);
or U8264 (N_8264,N_4435,N_2763);
xor U8265 (N_8265,N_3531,N_2468);
and U8266 (N_8266,N_4905,N_592);
or U8267 (N_8267,N_1637,N_3827);
or U8268 (N_8268,N_1533,N_4368);
and U8269 (N_8269,N_3899,N_1491);
xnor U8270 (N_8270,N_1694,N_505);
nand U8271 (N_8271,N_3935,N_2148);
xnor U8272 (N_8272,N_4910,N_2556);
or U8273 (N_8273,N_4762,N_2758);
and U8274 (N_8274,N_3851,N_1721);
nor U8275 (N_8275,N_2275,N_224);
nand U8276 (N_8276,N_2408,N_4761);
xnor U8277 (N_8277,N_2557,N_196);
nand U8278 (N_8278,N_3851,N_4552);
nor U8279 (N_8279,N_906,N_2932);
nor U8280 (N_8280,N_3957,N_4513);
nand U8281 (N_8281,N_1242,N_4288);
nand U8282 (N_8282,N_3544,N_4127);
nor U8283 (N_8283,N_3309,N_1133);
or U8284 (N_8284,N_3821,N_4400);
nand U8285 (N_8285,N_3255,N_4377);
and U8286 (N_8286,N_745,N_2951);
or U8287 (N_8287,N_1119,N_242);
nor U8288 (N_8288,N_2307,N_1232);
and U8289 (N_8289,N_1284,N_1941);
and U8290 (N_8290,N_2587,N_1084);
nor U8291 (N_8291,N_2693,N_3376);
and U8292 (N_8292,N_1588,N_3010);
nor U8293 (N_8293,N_231,N_4748);
and U8294 (N_8294,N_4216,N_3358);
and U8295 (N_8295,N_4718,N_773);
and U8296 (N_8296,N_972,N_4810);
nor U8297 (N_8297,N_2769,N_364);
and U8298 (N_8298,N_1385,N_4404);
nor U8299 (N_8299,N_1794,N_2927);
and U8300 (N_8300,N_2114,N_2729);
and U8301 (N_8301,N_3920,N_539);
nor U8302 (N_8302,N_277,N_3559);
xor U8303 (N_8303,N_2827,N_1228);
nand U8304 (N_8304,N_4436,N_1743);
nand U8305 (N_8305,N_3092,N_72);
or U8306 (N_8306,N_2762,N_4643);
xor U8307 (N_8307,N_2201,N_1963);
nand U8308 (N_8308,N_4911,N_2041);
and U8309 (N_8309,N_4197,N_3059);
and U8310 (N_8310,N_2208,N_3723);
nor U8311 (N_8311,N_2447,N_2491);
nand U8312 (N_8312,N_1744,N_358);
and U8313 (N_8313,N_4040,N_3968);
or U8314 (N_8314,N_1681,N_3469);
nand U8315 (N_8315,N_1607,N_2381);
or U8316 (N_8316,N_527,N_1129);
and U8317 (N_8317,N_1170,N_4510);
nor U8318 (N_8318,N_3139,N_1866);
xnor U8319 (N_8319,N_3674,N_345);
nor U8320 (N_8320,N_3288,N_2728);
and U8321 (N_8321,N_1380,N_541);
nand U8322 (N_8322,N_1261,N_608);
and U8323 (N_8323,N_2547,N_4880);
nor U8324 (N_8324,N_4780,N_3970);
nand U8325 (N_8325,N_2523,N_2163);
nor U8326 (N_8326,N_2721,N_4641);
nor U8327 (N_8327,N_1965,N_4218);
nand U8328 (N_8328,N_3255,N_558);
or U8329 (N_8329,N_2604,N_1093);
nor U8330 (N_8330,N_3878,N_4946);
nand U8331 (N_8331,N_3048,N_3292);
or U8332 (N_8332,N_655,N_2239);
and U8333 (N_8333,N_3670,N_1541);
nand U8334 (N_8334,N_4024,N_3206);
and U8335 (N_8335,N_1598,N_2525);
and U8336 (N_8336,N_4850,N_1638);
nand U8337 (N_8337,N_2200,N_1922);
or U8338 (N_8338,N_4953,N_2860);
or U8339 (N_8339,N_737,N_4233);
or U8340 (N_8340,N_4453,N_70);
xor U8341 (N_8341,N_2191,N_2853);
nor U8342 (N_8342,N_1401,N_3285);
nor U8343 (N_8343,N_627,N_541);
nand U8344 (N_8344,N_3541,N_3396);
and U8345 (N_8345,N_1662,N_367);
and U8346 (N_8346,N_1702,N_2662);
and U8347 (N_8347,N_1444,N_4013);
nor U8348 (N_8348,N_2797,N_2057);
and U8349 (N_8349,N_4359,N_3309);
nand U8350 (N_8350,N_3507,N_2098);
nand U8351 (N_8351,N_1276,N_3731);
nand U8352 (N_8352,N_3068,N_2548);
nor U8353 (N_8353,N_2758,N_4179);
nand U8354 (N_8354,N_2780,N_3703);
and U8355 (N_8355,N_1971,N_1562);
nor U8356 (N_8356,N_3832,N_1146);
nor U8357 (N_8357,N_1554,N_1794);
or U8358 (N_8358,N_1853,N_1823);
xnor U8359 (N_8359,N_3017,N_2101);
and U8360 (N_8360,N_307,N_1972);
nand U8361 (N_8361,N_4320,N_3604);
and U8362 (N_8362,N_4394,N_3275);
nor U8363 (N_8363,N_2158,N_1828);
nor U8364 (N_8364,N_2593,N_4591);
or U8365 (N_8365,N_1336,N_3970);
nor U8366 (N_8366,N_1635,N_1976);
and U8367 (N_8367,N_2738,N_4079);
or U8368 (N_8368,N_221,N_964);
or U8369 (N_8369,N_3080,N_1685);
nor U8370 (N_8370,N_888,N_2309);
nor U8371 (N_8371,N_1294,N_494);
nand U8372 (N_8372,N_837,N_2952);
nand U8373 (N_8373,N_3326,N_2223);
nor U8374 (N_8374,N_2736,N_357);
nor U8375 (N_8375,N_4141,N_1892);
or U8376 (N_8376,N_866,N_3957);
and U8377 (N_8377,N_2307,N_4079);
and U8378 (N_8378,N_4803,N_3536);
xor U8379 (N_8379,N_4834,N_1352);
and U8380 (N_8380,N_2349,N_1136);
and U8381 (N_8381,N_180,N_1511);
or U8382 (N_8382,N_546,N_2216);
and U8383 (N_8383,N_1487,N_838);
or U8384 (N_8384,N_2952,N_1035);
nand U8385 (N_8385,N_3435,N_3100);
xnor U8386 (N_8386,N_1692,N_4556);
xnor U8387 (N_8387,N_272,N_450);
nand U8388 (N_8388,N_4323,N_1953);
or U8389 (N_8389,N_696,N_197);
nand U8390 (N_8390,N_4634,N_1093);
nor U8391 (N_8391,N_3660,N_1575);
nor U8392 (N_8392,N_2806,N_857);
nand U8393 (N_8393,N_4859,N_1848);
and U8394 (N_8394,N_3008,N_1760);
and U8395 (N_8395,N_2026,N_4169);
nand U8396 (N_8396,N_660,N_4023);
nand U8397 (N_8397,N_529,N_3197);
nand U8398 (N_8398,N_3774,N_3877);
or U8399 (N_8399,N_4645,N_214);
xnor U8400 (N_8400,N_4868,N_3152);
and U8401 (N_8401,N_2495,N_4566);
nand U8402 (N_8402,N_3979,N_1423);
or U8403 (N_8403,N_2501,N_2386);
or U8404 (N_8404,N_1184,N_535);
and U8405 (N_8405,N_1397,N_4796);
nand U8406 (N_8406,N_4256,N_197);
and U8407 (N_8407,N_1013,N_1175);
nand U8408 (N_8408,N_4006,N_1692);
nand U8409 (N_8409,N_1260,N_1207);
xnor U8410 (N_8410,N_145,N_244);
and U8411 (N_8411,N_3178,N_3877);
and U8412 (N_8412,N_4084,N_4726);
xor U8413 (N_8413,N_3193,N_27);
or U8414 (N_8414,N_200,N_4463);
and U8415 (N_8415,N_2957,N_871);
nor U8416 (N_8416,N_3752,N_740);
and U8417 (N_8417,N_2964,N_3549);
and U8418 (N_8418,N_2597,N_3386);
xor U8419 (N_8419,N_2487,N_4258);
and U8420 (N_8420,N_1447,N_2668);
and U8421 (N_8421,N_1603,N_645);
or U8422 (N_8422,N_957,N_1652);
and U8423 (N_8423,N_872,N_585);
or U8424 (N_8424,N_233,N_2565);
nor U8425 (N_8425,N_694,N_2833);
or U8426 (N_8426,N_4522,N_3987);
nor U8427 (N_8427,N_3357,N_86);
and U8428 (N_8428,N_4505,N_702);
nand U8429 (N_8429,N_3026,N_964);
nand U8430 (N_8430,N_1737,N_2728);
and U8431 (N_8431,N_2309,N_1207);
nand U8432 (N_8432,N_4856,N_1318);
and U8433 (N_8433,N_3715,N_4959);
or U8434 (N_8434,N_3454,N_344);
or U8435 (N_8435,N_3799,N_2934);
nor U8436 (N_8436,N_4650,N_1933);
nand U8437 (N_8437,N_1789,N_1177);
or U8438 (N_8438,N_141,N_1225);
nor U8439 (N_8439,N_818,N_1137);
or U8440 (N_8440,N_3220,N_2920);
and U8441 (N_8441,N_3338,N_4642);
and U8442 (N_8442,N_288,N_1585);
nand U8443 (N_8443,N_533,N_439);
nand U8444 (N_8444,N_2250,N_4958);
and U8445 (N_8445,N_3136,N_1693);
or U8446 (N_8446,N_2349,N_3319);
nand U8447 (N_8447,N_4786,N_4828);
nand U8448 (N_8448,N_2248,N_407);
nor U8449 (N_8449,N_1288,N_1190);
nand U8450 (N_8450,N_4284,N_2377);
nand U8451 (N_8451,N_3190,N_4338);
nand U8452 (N_8452,N_737,N_1931);
nor U8453 (N_8453,N_926,N_3078);
xnor U8454 (N_8454,N_88,N_4628);
and U8455 (N_8455,N_3331,N_2582);
nor U8456 (N_8456,N_3428,N_1606);
nand U8457 (N_8457,N_185,N_3214);
xnor U8458 (N_8458,N_3526,N_1151);
and U8459 (N_8459,N_4075,N_1452);
or U8460 (N_8460,N_1061,N_2317);
nand U8461 (N_8461,N_2248,N_2849);
nor U8462 (N_8462,N_126,N_1200);
or U8463 (N_8463,N_338,N_697);
or U8464 (N_8464,N_597,N_283);
nand U8465 (N_8465,N_1795,N_2145);
nor U8466 (N_8466,N_2334,N_4542);
nor U8467 (N_8467,N_3828,N_2399);
nand U8468 (N_8468,N_4770,N_2566);
or U8469 (N_8469,N_3405,N_4064);
xnor U8470 (N_8470,N_3529,N_4326);
nand U8471 (N_8471,N_3694,N_1187);
and U8472 (N_8472,N_3320,N_2973);
nand U8473 (N_8473,N_2481,N_4828);
nand U8474 (N_8474,N_3922,N_49);
or U8475 (N_8475,N_4037,N_3502);
xor U8476 (N_8476,N_14,N_890);
and U8477 (N_8477,N_1290,N_1217);
nor U8478 (N_8478,N_2074,N_4746);
nand U8479 (N_8479,N_2632,N_4176);
or U8480 (N_8480,N_4437,N_2624);
nor U8481 (N_8481,N_2999,N_74);
and U8482 (N_8482,N_2832,N_869);
and U8483 (N_8483,N_1528,N_910);
and U8484 (N_8484,N_414,N_2847);
nand U8485 (N_8485,N_3648,N_4608);
or U8486 (N_8486,N_853,N_3039);
nand U8487 (N_8487,N_795,N_2055);
nor U8488 (N_8488,N_2750,N_4717);
nor U8489 (N_8489,N_3042,N_2166);
or U8490 (N_8490,N_2878,N_1062);
and U8491 (N_8491,N_2292,N_4924);
nand U8492 (N_8492,N_439,N_3935);
nor U8493 (N_8493,N_4842,N_1841);
nand U8494 (N_8494,N_169,N_4233);
nand U8495 (N_8495,N_755,N_2278);
and U8496 (N_8496,N_3991,N_4208);
nor U8497 (N_8497,N_4934,N_668);
nand U8498 (N_8498,N_1592,N_608);
nor U8499 (N_8499,N_3562,N_58);
nand U8500 (N_8500,N_4719,N_4306);
nor U8501 (N_8501,N_4427,N_2217);
nor U8502 (N_8502,N_3192,N_2951);
or U8503 (N_8503,N_2323,N_531);
nor U8504 (N_8504,N_2693,N_1589);
or U8505 (N_8505,N_1949,N_3207);
nand U8506 (N_8506,N_54,N_2846);
and U8507 (N_8507,N_1080,N_3503);
or U8508 (N_8508,N_345,N_1928);
or U8509 (N_8509,N_1616,N_2900);
nand U8510 (N_8510,N_1815,N_1748);
and U8511 (N_8511,N_3949,N_1282);
and U8512 (N_8512,N_3830,N_2239);
nor U8513 (N_8513,N_1746,N_2440);
and U8514 (N_8514,N_4229,N_688);
nor U8515 (N_8515,N_4386,N_2295);
and U8516 (N_8516,N_631,N_125);
nor U8517 (N_8517,N_3701,N_865);
xnor U8518 (N_8518,N_400,N_3230);
or U8519 (N_8519,N_2471,N_25);
xnor U8520 (N_8520,N_4294,N_2519);
and U8521 (N_8521,N_699,N_2859);
xnor U8522 (N_8522,N_3708,N_1894);
and U8523 (N_8523,N_1865,N_1416);
xnor U8524 (N_8524,N_3686,N_1492);
nand U8525 (N_8525,N_1126,N_3776);
and U8526 (N_8526,N_734,N_4485);
and U8527 (N_8527,N_3377,N_1286);
xnor U8528 (N_8528,N_4715,N_2754);
xnor U8529 (N_8529,N_980,N_3983);
nand U8530 (N_8530,N_4868,N_1231);
xor U8531 (N_8531,N_2659,N_487);
and U8532 (N_8532,N_2390,N_3077);
nand U8533 (N_8533,N_4494,N_2990);
and U8534 (N_8534,N_1517,N_1836);
or U8535 (N_8535,N_3144,N_2484);
or U8536 (N_8536,N_2608,N_2116);
and U8537 (N_8537,N_2302,N_1473);
xnor U8538 (N_8538,N_1311,N_2939);
and U8539 (N_8539,N_3826,N_1882);
and U8540 (N_8540,N_4235,N_2458);
or U8541 (N_8541,N_1751,N_62);
and U8542 (N_8542,N_2585,N_241);
nand U8543 (N_8543,N_4894,N_3224);
or U8544 (N_8544,N_1365,N_4450);
nor U8545 (N_8545,N_928,N_1066);
nor U8546 (N_8546,N_2055,N_56);
nor U8547 (N_8547,N_1318,N_1665);
and U8548 (N_8548,N_129,N_1073);
or U8549 (N_8549,N_956,N_1118);
and U8550 (N_8550,N_2068,N_2699);
nor U8551 (N_8551,N_3820,N_1738);
or U8552 (N_8552,N_3221,N_2726);
nor U8553 (N_8553,N_1528,N_3260);
or U8554 (N_8554,N_4741,N_3472);
or U8555 (N_8555,N_785,N_4818);
nand U8556 (N_8556,N_1594,N_1452);
and U8557 (N_8557,N_1813,N_3611);
xor U8558 (N_8558,N_1088,N_1339);
and U8559 (N_8559,N_4834,N_272);
nand U8560 (N_8560,N_2789,N_4058);
nand U8561 (N_8561,N_1571,N_2659);
nand U8562 (N_8562,N_4641,N_261);
or U8563 (N_8563,N_2555,N_3743);
nor U8564 (N_8564,N_4502,N_3934);
nor U8565 (N_8565,N_3245,N_2431);
nand U8566 (N_8566,N_4933,N_8);
and U8567 (N_8567,N_1153,N_3011);
xor U8568 (N_8568,N_4397,N_105);
and U8569 (N_8569,N_4035,N_1783);
or U8570 (N_8570,N_3357,N_3526);
and U8571 (N_8571,N_1582,N_127);
nor U8572 (N_8572,N_3819,N_2424);
or U8573 (N_8573,N_4797,N_1004);
nand U8574 (N_8574,N_2116,N_2400);
nor U8575 (N_8575,N_204,N_3462);
nor U8576 (N_8576,N_3157,N_2042);
nor U8577 (N_8577,N_994,N_4405);
xor U8578 (N_8578,N_4530,N_2619);
nor U8579 (N_8579,N_1821,N_524);
and U8580 (N_8580,N_4896,N_4588);
nor U8581 (N_8581,N_1968,N_3860);
and U8582 (N_8582,N_3644,N_4630);
or U8583 (N_8583,N_2402,N_3370);
and U8584 (N_8584,N_4790,N_4984);
nor U8585 (N_8585,N_4924,N_503);
nor U8586 (N_8586,N_3660,N_1316);
nand U8587 (N_8587,N_4736,N_2364);
nor U8588 (N_8588,N_946,N_4197);
nand U8589 (N_8589,N_1261,N_4565);
nand U8590 (N_8590,N_4745,N_1951);
or U8591 (N_8591,N_1163,N_2445);
nand U8592 (N_8592,N_1702,N_1135);
nor U8593 (N_8593,N_2966,N_2980);
and U8594 (N_8594,N_1992,N_475);
or U8595 (N_8595,N_2295,N_533);
nand U8596 (N_8596,N_3764,N_4907);
or U8597 (N_8597,N_1375,N_1737);
nor U8598 (N_8598,N_1538,N_4475);
nand U8599 (N_8599,N_3998,N_4567);
or U8600 (N_8600,N_238,N_1663);
nor U8601 (N_8601,N_1870,N_1893);
and U8602 (N_8602,N_1366,N_527);
and U8603 (N_8603,N_883,N_4078);
or U8604 (N_8604,N_2363,N_453);
or U8605 (N_8605,N_3164,N_4093);
and U8606 (N_8606,N_3733,N_946);
nor U8607 (N_8607,N_1702,N_4625);
or U8608 (N_8608,N_1697,N_456);
nor U8609 (N_8609,N_3223,N_4576);
or U8610 (N_8610,N_2566,N_1407);
xor U8611 (N_8611,N_1948,N_1337);
and U8612 (N_8612,N_4982,N_524);
nor U8613 (N_8613,N_2235,N_2038);
or U8614 (N_8614,N_290,N_2652);
or U8615 (N_8615,N_3640,N_490);
nand U8616 (N_8616,N_2591,N_4400);
nand U8617 (N_8617,N_4507,N_161);
or U8618 (N_8618,N_459,N_2680);
nor U8619 (N_8619,N_3417,N_693);
or U8620 (N_8620,N_2709,N_2313);
xor U8621 (N_8621,N_3300,N_870);
nor U8622 (N_8622,N_1399,N_4518);
or U8623 (N_8623,N_3120,N_3199);
nand U8624 (N_8624,N_672,N_1976);
nor U8625 (N_8625,N_2444,N_4307);
and U8626 (N_8626,N_1704,N_1113);
nor U8627 (N_8627,N_722,N_156);
or U8628 (N_8628,N_4567,N_4768);
or U8629 (N_8629,N_11,N_3358);
nand U8630 (N_8630,N_3097,N_2142);
and U8631 (N_8631,N_3625,N_4032);
xor U8632 (N_8632,N_418,N_249);
or U8633 (N_8633,N_3984,N_2236);
nor U8634 (N_8634,N_3214,N_3597);
or U8635 (N_8635,N_1281,N_1844);
or U8636 (N_8636,N_4633,N_853);
nor U8637 (N_8637,N_1981,N_2325);
or U8638 (N_8638,N_3780,N_1774);
nand U8639 (N_8639,N_4219,N_991);
nor U8640 (N_8640,N_4106,N_1987);
nor U8641 (N_8641,N_3779,N_932);
xnor U8642 (N_8642,N_3090,N_424);
and U8643 (N_8643,N_2748,N_3584);
nand U8644 (N_8644,N_2516,N_235);
and U8645 (N_8645,N_2246,N_2203);
or U8646 (N_8646,N_510,N_1579);
or U8647 (N_8647,N_3964,N_828);
and U8648 (N_8648,N_1982,N_3779);
nand U8649 (N_8649,N_152,N_3528);
or U8650 (N_8650,N_1409,N_889);
nor U8651 (N_8651,N_1524,N_4654);
nor U8652 (N_8652,N_1613,N_2744);
and U8653 (N_8653,N_2662,N_3140);
and U8654 (N_8654,N_463,N_2138);
or U8655 (N_8655,N_3635,N_3571);
and U8656 (N_8656,N_4583,N_2084);
and U8657 (N_8657,N_3987,N_1672);
nand U8658 (N_8658,N_1302,N_1731);
and U8659 (N_8659,N_1967,N_2726);
nand U8660 (N_8660,N_1416,N_4980);
and U8661 (N_8661,N_3198,N_643);
nand U8662 (N_8662,N_359,N_2423);
xor U8663 (N_8663,N_573,N_4142);
nand U8664 (N_8664,N_524,N_523);
nand U8665 (N_8665,N_1935,N_3763);
and U8666 (N_8666,N_4973,N_878);
and U8667 (N_8667,N_3703,N_485);
nand U8668 (N_8668,N_906,N_3937);
or U8669 (N_8669,N_4668,N_2337);
or U8670 (N_8670,N_3065,N_4886);
nand U8671 (N_8671,N_1309,N_2828);
or U8672 (N_8672,N_3199,N_88);
nor U8673 (N_8673,N_4359,N_2779);
nor U8674 (N_8674,N_4475,N_4023);
nor U8675 (N_8675,N_55,N_2213);
or U8676 (N_8676,N_1365,N_3781);
nand U8677 (N_8677,N_4134,N_3157);
and U8678 (N_8678,N_2220,N_1434);
nand U8679 (N_8679,N_619,N_506);
or U8680 (N_8680,N_4870,N_419);
xnor U8681 (N_8681,N_2088,N_501);
nor U8682 (N_8682,N_3637,N_474);
xor U8683 (N_8683,N_4383,N_4194);
nand U8684 (N_8684,N_3925,N_598);
nor U8685 (N_8685,N_2556,N_4819);
and U8686 (N_8686,N_2252,N_3032);
nor U8687 (N_8687,N_2433,N_1459);
or U8688 (N_8688,N_419,N_1802);
xor U8689 (N_8689,N_4667,N_4340);
nand U8690 (N_8690,N_4147,N_1320);
nand U8691 (N_8691,N_1957,N_585);
nor U8692 (N_8692,N_314,N_459);
nand U8693 (N_8693,N_4761,N_229);
nor U8694 (N_8694,N_280,N_4321);
nor U8695 (N_8695,N_4088,N_790);
nand U8696 (N_8696,N_496,N_1797);
nand U8697 (N_8697,N_4485,N_4007);
nor U8698 (N_8698,N_431,N_2480);
nor U8699 (N_8699,N_3837,N_441);
or U8700 (N_8700,N_1238,N_499);
nor U8701 (N_8701,N_502,N_3947);
nor U8702 (N_8702,N_3593,N_3172);
or U8703 (N_8703,N_148,N_2436);
nand U8704 (N_8704,N_4688,N_331);
and U8705 (N_8705,N_3097,N_4853);
or U8706 (N_8706,N_3115,N_4637);
or U8707 (N_8707,N_1581,N_4061);
nor U8708 (N_8708,N_3472,N_3875);
nand U8709 (N_8709,N_2826,N_3061);
nor U8710 (N_8710,N_3992,N_479);
nand U8711 (N_8711,N_4827,N_3806);
nand U8712 (N_8712,N_1558,N_928);
nand U8713 (N_8713,N_3711,N_3348);
nand U8714 (N_8714,N_3152,N_3091);
or U8715 (N_8715,N_1843,N_757);
and U8716 (N_8716,N_1000,N_1651);
or U8717 (N_8717,N_1205,N_1667);
nand U8718 (N_8718,N_4633,N_1707);
or U8719 (N_8719,N_2448,N_4801);
xnor U8720 (N_8720,N_581,N_3230);
nand U8721 (N_8721,N_2194,N_369);
nor U8722 (N_8722,N_1541,N_539);
nor U8723 (N_8723,N_3765,N_3300);
nor U8724 (N_8724,N_3068,N_1444);
nand U8725 (N_8725,N_4819,N_3616);
nand U8726 (N_8726,N_4661,N_1853);
or U8727 (N_8727,N_443,N_342);
and U8728 (N_8728,N_3618,N_3599);
xnor U8729 (N_8729,N_1915,N_593);
or U8730 (N_8730,N_4187,N_4137);
nand U8731 (N_8731,N_2617,N_4528);
nand U8732 (N_8732,N_2047,N_3279);
nand U8733 (N_8733,N_2782,N_4675);
nand U8734 (N_8734,N_1054,N_158);
nor U8735 (N_8735,N_2849,N_609);
nand U8736 (N_8736,N_2714,N_1074);
nor U8737 (N_8737,N_4392,N_4233);
nor U8738 (N_8738,N_696,N_3649);
nand U8739 (N_8739,N_3153,N_1949);
nand U8740 (N_8740,N_2649,N_1472);
xor U8741 (N_8741,N_463,N_285);
and U8742 (N_8742,N_4448,N_3821);
nand U8743 (N_8743,N_1738,N_2454);
nand U8744 (N_8744,N_3727,N_1363);
nand U8745 (N_8745,N_3217,N_2968);
and U8746 (N_8746,N_995,N_1114);
xnor U8747 (N_8747,N_1319,N_22);
nor U8748 (N_8748,N_3903,N_1305);
and U8749 (N_8749,N_2235,N_4665);
nor U8750 (N_8750,N_1574,N_3399);
xnor U8751 (N_8751,N_2442,N_3187);
or U8752 (N_8752,N_4822,N_2421);
nor U8753 (N_8753,N_1964,N_1250);
nor U8754 (N_8754,N_4418,N_94);
or U8755 (N_8755,N_3162,N_1381);
or U8756 (N_8756,N_3760,N_545);
nor U8757 (N_8757,N_1197,N_3276);
and U8758 (N_8758,N_145,N_4061);
or U8759 (N_8759,N_651,N_1587);
xnor U8760 (N_8760,N_1802,N_2623);
xor U8761 (N_8761,N_4252,N_806);
nand U8762 (N_8762,N_530,N_4256);
nor U8763 (N_8763,N_310,N_1020);
or U8764 (N_8764,N_2620,N_1982);
or U8765 (N_8765,N_2540,N_3349);
or U8766 (N_8766,N_2022,N_1067);
or U8767 (N_8767,N_3794,N_4308);
and U8768 (N_8768,N_2489,N_2643);
nand U8769 (N_8769,N_1604,N_1791);
or U8770 (N_8770,N_4939,N_583);
nand U8771 (N_8771,N_1355,N_3166);
nand U8772 (N_8772,N_1144,N_1053);
nor U8773 (N_8773,N_110,N_355);
xnor U8774 (N_8774,N_1950,N_2136);
nand U8775 (N_8775,N_1707,N_3102);
and U8776 (N_8776,N_2449,N_836);
or U8777 (N_8777,N_922,N_2325);
xnor U8778 (N_8778,N_2851,N_3355);
and U8779 (N_8779,N_1745,N_622);
xor U8780 (N_8780,N_4603,N_3630);
nor U8781 (N_8781,N_2106,N_54);
nand U8782 (N_8782,N_1408,N_3267);
nor U8783 (N_8783,N_4113,N_2831);
xor U8784 (N_8784,N_3378,N_4472);
and U8785 (N_8785,N_1425,N_1878);
xor U8786 (N_8786,N_4885,N_2741);
xnor U8787 (N_8787,N_536,N_141);
nand U8788 (N_8788,N_2519,N_3248);
and U8789 (N_8789,N_1309,N_858);
nand U8790 (N_8790,N_3200,N_2013);
nand U8791 (N_8791,N_4436,N_3930);
and U8792 (N_8792,N_3826,N_3184);
nor U8793 (N_8793,N_2733,N_4466);
or U8794 (N_8794,N_274,N_3786);
and U8795 (N_8795,N_767,N_28);
nor U8796 (N_8796,N_4216,N_2457);
and U8797 (N_8797,N_1395,N_2725);
or U8798 (N_8798,N_96,N_1050);
nand U8799 (N_8799,N_3362,N_300);
nor U8800 (N_8800,N_2263,N_1159);
nand U8801 (N_8801,N_4077,N_341);
xor U8802 (N_8802,N_3135,N_4571);
nor U8803 (N_8803,N_1941,N_1625);
nand U8804 (N_8804,N_2712,N_1651);
or U8805 (N_8805,N_4075,N_4462);
or U8806 (N_8806,N_4310,N_3056);
or U8807 (N_8807,N_2235,N_228);
or U8808 (N_8808,N_4926,N_4424);
nor U8809 (N_8809,N_2860,N_4575);
nand U8810 (N_8810,N_3190,N_3454);
nor U8811 (N_8811,N_2576,N_2435);
nand U8812 (N_8812,N_2049,N_3262);
and U8813 (N_8813,N_2507,N_3438);
xor U8814 (N_8814,N_1747,N_690);
and U8815 (N_8815,N_1959,N_4848);
nand U8816 (N_8816,N_3523,N_1674);
or U8817 (N_8817,N_4271,N_3885);
and U8818 (N_8818,N_3919,N_4971);
nor U8819 (N_8819,N_3509,N_3761);
nand U8820 (N_8820,N_3631,N_573);
xnor U8821 (N_8821,N_944,N_3287);
and U8822 (N_8822,N_2302,N_3331);
nand U8823 (N_8823,N_1963,N_2415);
and U8824 (N_8824,N_120,N_1130);
xor U8825 (N_8825,N_152,N_4248);
and U8826 (N_8826,N_1122,N_4950);
nand U8827 (N_8827,N_2624,N_3995);
nand U8828 (N_8828,N_2485,N_3570);
and U8829 (N_8829,N_2513,N_540);
and U8830 (N_8830,N_1165,N_1141);
and U8831 (N_8831,N_1162,N_3748);
or U8832 (N_8832,N_2812,N_1243);
or U8833 (N_8833,N_1443,N_4749);
nor U8834 (N_8834,N_2338,N_3893);
nor U8835 (N_8835,N_1420,N_2391);
or U8836 (N_8836,N_1418,N_4823);
and U8837 (N_8837,N_3272,N_2761);
nand U8838 (N_8838,N_212,N_4403);
or U8839 (N_8839,N_2409,N_4187);
nor U8840 (N_8840,N_610,N_3762);
or U8841 (N_8841,N_2477,N_4760);
nand U8842 (N_8842,N_4279,N_1460);
nor U8843 (N_8843,N_1114,N_3608);
nand U8844 (N_8844,N_3631,N_4247);
or U8845 (N_8845,N_3403,N_2199);
xor U8846 (N_8846,N_219,N_3583);
or U8847 (N_8847,N_3659,N_2796);
and U8848 (N_8848,N_1750,N_1359);
and U8849 (N_8849,N_2367,N_286);
and U8850 (N_8850,N_3927,N_3536);
nand U8851 (N_8851,N_3273,N_2952);
and U8852 (N_8852,N_1479,N_4888);
xnor U8853 (N_8853,N_4428,N_3307);
or U8854 (N_8854,N_2208,N_125);
or U8855 (N_8855,N_1789,N_2077);
nand U8856 (N_8856,N_3113,N_1612);
nand U8857 (N_8857,N_2520,N_1054);
and U8858 (N_8858,N_4259,N_401);
nor U8859 (N_8859,N_3876,N_4976);
or U8860 (N_8860,N_70,N_430);
or U8861 (N_8861,N_876,N_4899);
or U8862 (N_8862,N_3446,N_3611);
nand U8863 (N_8863,N_4305,N_2952);
or U8864 (N_8864,N_331,N_4458);
nor U8865 (N_8865,N_1100,N_2914);
xnor U8866 (N_8866,N_4198,N_556);
and U8867 (N_8867,N_1460,N_4876);
and U8868 (N_8868,N_4558,N_1518);
or U8869 (N_8869,N_3747,N_3219);
or U8870 (N_8870,N_2553,N_208);
and U8871 (N_8871,N_4674,N_3106);
nor U8872 (N_8872,N_3603,N_2998);
or U8873 (N_8873,N_4827,N_1284);
nor U8874 (N_8874,N_1806,N_1312);
or U8875 (N_8875,N_681,N_1086);
and U8876 (N_8876,N_4996,N_638);
or U8877 (N_8877,N_4774,N_242);
and U8878 (N_8878,N_828,N_4734);
or U8879 (N_8879,N_2196,N_963);
nand U8880 (N_8880,N_475,N_4503);
nor U8881 (N_8881,N_4145,N_4219);
xor U8882 (N_8882,N_2554,N_3917);
nand U8883 (N_8883,N_4645,N_4078);
or U8884 (N_8884,N_3242,N_2359);
nand U8885 (N_8885,N_3771,N_3682);
nand U8886 (N_8886,N_3896,N_4760);
nor U8887 (N_8887,N_4322,N_492);
nand U8888 (N_8888,N_0,N_2028);
nor U8889 (N_8889,N_1698,N_238);
xnor U8890 (N_8890,N_196,N_4138);
nor U8891 (N_8891,N_2228,N_736);
nand U8892 (N_8892,N_4499,N_717);
nand U8893 (N_8893,N_3652,N_4149);
nor U8894 (N_8894,N_2280,N_3353);
and U8895 (N_8895,N_2413,N_3219);
and U8896 (N_8896,N_2870,N_1767);
nor U8897 (N_8897,N_4396,N_2822);
or U8898 (N_8898,N_3588,N_4246);
and U8899 (N_8899,N_2724,N_2550);
or U8900 (N_8900,N_3191,N_1677);
nor U8901 (N_8901,N_3231,N_4092);
nand U8902 (N_8902,N_3071,N_2258);
nand U8903 (N_8903,N_3590,N_1248);
xor U8904 (N_8904,N_2952,N_4550);
nand U8905 (N_8905,N_2390,N_1754);
and U8906 (N_8906,N_3344,N_689);
nand U8907 (N_8907,N_2769,N_4693);
and U8908 (N_8908,N_32,N_4613);
nand U8909 (N_8909,N_3246,N_2992);
nand U8910 (N_8910,N_4036,N_443);
xnor U8911 (N_8911,N_3826,N_4314);
or U8912 (N_8912,N_51,N_251);
nand U8913 (N_8913,N_2418,N_4494);
or U8914 (N_8914,N_1115,N_186);
or U8915 (N_8915,N_1418,N_697);
nand U8916 (N_8916,N_538,N_2953);
and U8917 (N_8917,N_2779,N_3242);
xnor U8918 (N_8918,N_3188,N_1513);
nand U8919 (N_8919,N_4680,N_113);
and U8920 (N_8920,N_3878,N_1633);
or U8921 (N_8921,N_430,N_3599);
nor U8922 (N_8922,N_920,N_3484);
nand U8923 (N_8923,N_3077,N_3007);
nand U8924 (N_8924,N_1310,N_1916);
or U8925 (N_8925,N_2100,N_4416);
nor U8926 (N_8926,N_1508,N_1758);
or U8927 (N_8927,N_2428,N_4679);
nand U8928 (N_8928,N_2135,N_550);
and U8929 (N_8929,N_4081,N_1365);
nand U8930 (N_8930,N_2190,N_4881);
nand U8931 (N_8931,N_4577,N_2705);
nor U8932 (N_8932,N_2635,N_563);
nand U8933 (N_8933,N_2468,N_4358);
nand U8934 (N_8934,N_4020,N_1145);
nand U8935 (N_8935,N_1068,N_183);
xor U8936 (N_8936,N_3930,N_520);
nor U8937 (N_8937,N_3694,N_1387);
or U8938 (N_8938,N_3775,N_1372);
nand U8939 (N_8939,N_581,N_3201);
or U8940 (N_8940,N_2398,N_793);
or U8941 (N_8941,N_4647,N_1738);
nand U8942 (N_8942,N_3899,N_4072);
and U8943 (N_8943,N_2638,N_3573);
nand U8944 (N_8944,N_2595,N_3173);
or U8945 (N_8945,N_1578,N_458);
and U8946 (N_8946,N_3700,N_1566);
nor U8947 (N_8947,N_3548,N_4722);
and U8948 (N_8948,N_4100,N_2249);
nor U8949 (N_8949,N_1213,N_663);
and U8950 (N_8950,N_4598,N_2510);
nor U8951 (N_8951,N_4882,N_3844);
nor U8952 (N_8952,N_443,N_4258);
xnor U8953 (N_8953,N_828,N_3185);
nor U8954 (N_8954,N_3605,N_3094);
nand U8955 (N_8955,N_171,N_262);
nand U8956 (N_8956,N_4425,N_1846);
and U8957 (N_8957,N_2812,N_3942);
and U8958 (N_8958,N_1009,N_3460);
nor U8959 (N_8959,N_4859,N_4701);
and U8960 (N_8960,N_1700,N_750);
and U8961 (N_8961,N_181,N_969);
or U8962 (N_8962,N_922,N_1503);
and U8963 (N_8963,N_189,N_4623);
nor U8964 (N_8964,N_3915,N_4992);
xnor U8965 (N_8965,N_2378,N_2526);
and U8966 (N_8966,N_1788,N_4663);
nand U8967 (N_8967,N_4631,N_1057);
nand U8968 (N_8968,N_98,N_3849);
nand U8969 (N_8969,N_2900,N_4462);
nand U8970 (N_8970,N_609,N_1705);
or U8971 (N_8971,N_3891,N_100);
and U8972 (N_8972,N_2561,N_3383);
and U8973 (N_8973,N_371,N_658);
xor U8974 (N_8974,N_1385,N_593);
nand U8975 (N_8975,N_3925,N_3028);
and U8976 (N_8976,N_1605,N_665);
or U8977 (N_8977,N_4596,N_2894);
or U8978 (N_8978,N_3495,N_4927);
or U8979 (N_8979,N_2981,N_3813);
nand U8980 (N_8980,N_4466,N_3334);
nand U8981 (N_8981,N_4445,N_3848);
nor U8982 (N_8982,N_2338,N_3956);
and U8983 (N_8983,N_3281,N_683);
nor U8984 (N_8984,N_3890,N_302);
xnor U8985 (N_8985,N_1204,N_3708);
nand U8986 (N_8986,N_867,N_4586);
xor U8987 (N_8987,N_4523,N_783);
nor U8988 (N_8988,N_3000,N_2368);
nor U8989 (N_8989,N_631,N_1438);
nor U8990 (N_8990,N_3362,N_3199);
and U8991 (N_8991,N_1197,N_2719);
xnor U8992 (N_8992,N_3811,N_3642);
and U8993 (N_8993,N_1261,N_1501);
nand U8994 (N_8994,N_2845,N_4689);
and U8995 (N_8995,N_2752,N_3607);
and U8996 (N_8996,N_3303,N_140);
nand U8997 (N_8997,N_1314,N_169);
or U8998 (N_8998,N_1098,N_3004);
or U8999 (N_8999,N_2090,N_3922);
or U9000 (N_9000,N_1607,N_2620);
nor U9001 (N_9001,N_2876,N_3393);
and U9002 (N_9002,N_2242,N_3855);
or U9003 (N_9003,N_2118,N_3165);
nor U9004 (N_9004,N_3971,N_1735);
or U9005 (N_9005,N_104,N_3846);
nand U9006 (N_9006,N_3045,N_3498);
or U9007 (N_9007,N_4888,N_4920);
nor U9008 (N_9008,N_1041,N_1944);
or U9009 (N_9009,N_1335,N_1279);
or U9010 (N_9010,N_985,N_4233);
and U9011 (N_9011,N_4627,N_1171);
and U9012 (N_9012,N_1574,N_4611);
xor U9013 (N_9013,N_469,N_220);
or U9014 (N_9014,N_2904,N_3413);
and U9015 (N_9015,N_4527,N_2395);
nor U9016 (N_9016,N_1923,N_3299);
nor U9017 (N_9017,N_2523,N_4744);
and U9018 (N_9018,N_3141,N_3856);
nand U9019 (N_9019,N_780,N_3861);
xor U9020 (N_9020,N_2688,N_4724);
and U9021 (N_9021,N_1727,N_524);
nor U9022 (N_9022,N_1434,N_782);
or U9023 (N_9023,N_2505,N_2936);
and U9024 (N_9024,N_4687,N_407);
or U9025 (N_9025,N_883,N_2154);
or U9026 (N_9026,N_1302,N_750);
nor U9027 (N_9027,N_3233,N_1169);
or U9028 (N_9028,N_4772,N_4082);
nand U9029 (N_9029,N_1620,N_2413);
nor U9030 (N_9030,N_3527,N_1932);
nor U9031 (N_9031,N_4634,N_1113);
nor U9032 (N_9032,N_1787,N_1561);
and U9033 (N_9033,N_4914,N_119);
and U9034 (N_9034,N_2678,N_4651);
nor U9035 (N_9035,N_2044,N_4662);
or U9036 (N_9036,N_1072,N_3161);
or U9037 (N_9037,N_4203,N_551);
and U9038 (N_9038,N_1794,N_2989);
and U9039 (N_9039,N_4954,N_4632);
and U9040 (N_9040,N_3360,N_293);
nor U9041 (N_9041,N_4180,N_338);
or U9042 (N_9042,N_468,N_3391);
or U9043 (N_9043,N_426,N_4425);
nand U9044 (N_9044,N_861,N_1265);
and U9045 (N_9045,N_848,N_3542);
and U9046 (N_9046,N_1170,N_2027);
and U9047 (N_9047,N_97,N_950);
xnor U9048 (N_9048,N_256,N_2851);
or U9049 (N_9049,N_2275,N_2780);
or U9050 (N_9050,N_4406,N_4099);
xor U9051 (N_9051,N_3151,N_114);
or U9052 (N_9052,N_1795,N_1162);
nand U9053 (N_9053,N_3655,N_3213);
nand U9054 (N_9054,N_2366,N_197);
and U9055 (N_9055,N_3654,N_2629);
or U9056 (N_9056,N_3164,N_4809);
xor U9057 (N_9057,N_3736,N_4522);
nand U9058 (N_9058,N_1666,N_3894);
and U9059 (N_9059,N_2104,N_1064);
xor U9060 (N_9060,N_2965,N_1998);
and U9061 (N_9061,N_1022,N_107);
or U9062 (N_9062,N_1890,N_287);
nand U9063 (N_9063,N_2603,N_1451);
or U9064 (N_9064,N_1512,N_1630);
or U9065 (N_9065,N_3573,N_3140);
and U9066 (N_9066,N_4343,N_2033);
nor U9067 (N_9067,N_2383,N_994);
nand U9068 (N_9068,N_2901,N_4118);
and U9069 (N_9069,N_4622,N_1726);
and U9070 (N_9070,N_2080,N_2892);
or U9071 (N_9071,N_3104,N_3485);
xor U9072 (N_9072,N_2254,N_4890);
nor U9073 (N_9073,N_3988,N_2439);
xor U9074 (N_9074,N_2784,N_4501);
nand U9075 (N_9075,N_3086,N_1323);
xnor U9076 (N_9076,N_4293,N_2895);
nor U9077 (N_9077,N_3849,N_4513);
or U9078 (N_9078,N_996,N_1477);
nand U9079 (N_9079,N_2402,N_1445);
xnor U9080 (N_9080,N_1039,N_3605);
nor U9081 (N_9081,N_1471,N_4403);
nor U9082 (N_9082,N_4024,N_2580);
nor U9083 (N_9083,N_3956,N_1431);
nor U9084 (N_9084,N_1100,N_3313);
nor U9085 (N_9085,N_2458,N_1460);
nor U9086 (N_9086,N_1688,N_3110);
xnor U9087 (N_9087,N_3924,N_80);
nand U9088 (N_9088,N_3559,N_2153);
nand U9089 (N_9089,N_1677,N_1243);
xnor U9090 (N_9090,N_2027,N_2704);
or U9091 (N_9091,N_1847,N_3327);
nand U9092 (N_9092,N_4129,N_3770);
nor U9093 (N_9093,N_15,N_4209);
nor U9094 (N_9094,N_2664,N_2268);
nor U9095 (N_9095,N_1780,N_1542);
and U9096 (N_9096,N_1165,N_3261);
or U9097 (N_9097,N_441,N_4291);
and U9098 (N_9098,N_74,N_3236);
nor U9099 (N_9099,N_294,N_3657);
xnor U9100 (N_9100,N_252,N_2756);
or U9101 (N_9101,N_2640,N_12);
or U9102 (N_9102,N_2255,N_4251);
nand U9103 (N_9103,N_3895,N_2041);
nand U9104 (N_9104,N_2303,N_1092);
xnor U9105 (N_9105,N_1273,N_1110);
or U9106 (N_9106,N_1483,N_1105);
nand U9107 (N_9107,N_4416,N_3834);
and U9108 (N_9108,N_1357,N_4322);
nor U9109 (N_9109,N_2910,N_2664);
or U9110 (N_9110,N_2338,N_314);
nand U9111 (N_9111,N_2351,N_2429);
nand U9112 (N_9112,N_288,N_1739);
and U9113 (N_9113,N_4266,N_2545);
or U9114 (N_9114,N_3902,N_4316);
xor U9115 (N_9115,N_594,N_1075);
nor U9116 (N_9116,N_4402,N_1098);
nand U9117 (N_9117,N_387,N_1832);
nor U9118 (N_9118,N_2586,N_4356);
xnor U9119 (N_9119,N_1089,N_3014);
and U9120 (N_9120,N_4154,N_3135);
nand U9121 (N_9121,N_4811,N_1532);
and U9122 (N_9122,N_3299,N_4666);
nand U9123 (N_9123,N_1811,N_2731);
nor U9124 (N_9124,N_3600,N_2267);
or U9125 (N_9125,N_234,N_4831);
nor U9126 (N_9126,N_487,N_1016);
nand U9127 (N_9127,N_2045,N_671);
nor U9128 (N_9128,N_4873,N_1036);
nand U9129 (N_9129,N_2331,N_835);
or U9130 (N_9130,N_3381,N_2522);
and U9131 (N_9131,N_4156,N_209);
or U9132 (N_9132,N_3032,N_2794);
or U9133 (N_9133,N_4182,N_2101);
xor U9134 (N_9134,N_2626,N_995);
nand U9135 (N_9135,N_2867,N_4817);
or U9136 (N_9136,N_3841,N_1450);
or U9137 (N_9137,N_469,N_853);
xor U9138 (N_9138,N_4133,N_4916);
and U9139 (N_9139,N_28,N_3850);
nor U9140 (N_9140,N_4100,N_1059);
and U9141 (N_9141,N_3219,N_2035);
or U9142 (N_9142,N_1939,N_1801);
or U9143 (N_9143,N_3486,N_4770);
nor U9144 (N_9144,N_2198,N_3199);
nor U9145 (N_9145,N_3613,N_3274);
and U9146 (N_9146,N_3657,N_2467);
xnor U9147 (N_9147,N_1929,N_1697);
nor U9148 (N_9148,N_4431,N_3299);
xor U9149 (N_9149,N_2609,N_4485);
nor U9150 (N_9150,N_2805,N_3904);
or U9151 (N_9151,N_3913,N_3541);
nor U9152 (N_9152,N_4172,N_769);
and U9153 (N_9153,N_571,N_2357);
nor U9154 (N_9154,N_2293,N_1712);
nand U9155 (N_9155,N_318,N_1983);
or U9156 (N_9156,N_2899,N_642);
and U9157 (N_9157,N_4992,N_300);
or U9158 (N_9158,N_2550,N_3676);
nand U9159 (N_9159,N_488,N_4075);
and U9160 (N_9160,N_4726,N_3974);
and U9161 (N_9161,N_1217,N_3543);
nor U9162 (N_9162,N_4355,N_3305);
and U9163 (N_9163,N_2414,N_2871);
xnor U9164 (N_9164,N_2979,N_1314);
nor U9165 (N_9165,N_1207,N_3261);
nor U9166 (N_9166,N_1393,N_2680);
or U9167 (N_9167,N_1907,N_365);
and U9168 (N_9168,N_4233,N_1981);
nand U9169 (N_9169,N_4007,N_88);
nor U9170 (N_9170,N_2631,N_3979);
nand U9171 (N_9171,N_1216,N_4692);
and U9172 (N_9172,N_4063,N_2649);
nand U9173 (N_9173,N_2979,N_3826);
nand U9174 (N_9174,N_1622,N_4073);
and U9175 (N_9175,N_1444,N_4542);
and U9176 (N_9176,N_1010,N_244);
or U9177 (N_9177,N_3016,N_4501);
or U9178 (N_9178,N_489,N_1650);
or U9179 (N_9179,N_914,N_177);
nor U9180 (N_9180,N_1210,N_1024);
and U9181 (N_9181,N_1148,N_672);
and U9182 (N_9182,N_1252,N_165);
xnor U9183 (N_9183,N_4694,N_4507);
or U9184 (N_9184,N_1918,N_2300);
nor U9185 (N_9185,N_1945,N_972);
nand U9186 (N_9186,N_782,N_2875);
or U9187 (N_9187,N_3350,N_3640);
nor U9188 (N_9188,N_3672,N_2175);
and U9189 (N_9189,N_2025,N_1146);
or U9190 (N_9190,N_1668,N_3587);
nor U9191 (N_9191,N_2094,N_2433);
and U9192 (N_9192,N_3889,N_3643);
and U9193 (N_9193,N_2955,N_374);
or U9194 (N_9194,N_3199,N_3394);
and U9195 (N_9195,N_3820,N_625);
nor U9196 (N_9196,N_3867,N_1899);
nand U9197 (N_9197,N_1324,N_2418);
or U9198 (N_9198,N_3744,N_2603);
nor U9199 (N_9199,N_2874,N_638);
and U9200 (N_9200,N_3202,N_3704);
nand U9201 (N_9201,N_3080,N_3051);
xor U9202 (N_9202,N_4885,N_1859);
or U9203 (N_9203,N_841,N_2441);
or U9204 (N_9204,N_4019,N_89);
nor U9205 (N_9205,N_3508,N_4673);
nand U9206 (N_9206,N_966,N_4139);
nor U9207 (N_9207,N_3320,N_1369);
and U9208 (N_9208,N_4424,N_467);
nor U9209 (N_9209,N_984,N_1764);
or U9210 (N_9210,N_4058,N_4309);
nor U9211 (N_9211,N_4383,N_4663);
nor U9212 (N_9212,N_4838,N_1044);
or U9213 (N_9213,N_4208,N_2483);
nor U9214 (N_9214,N_61,N_480);
nor U9215 (N_9215,N_839,N_4568);
and U9216 (N_9216,N_242,N_517);
nand U9217 (N_9217,N_3103,N_3104);
and U9218 (N_9218,N_299,N_3590);
nand U9219 (N_9219,N_535,N_934);
nand U9220 (N_9220,N_663,N_7);
nor U9221 (N_9221,N_15,N_1381);
or U9222 (N_9222,N_3783,N_4116);
and U9223 (N_9223,N_506,N_286);
and U9224 (N_9224,N_970,N_4994);
xor U9225 (N_9225,N_668,N_696);
nand U9226 (N_9226,N_603,N_3015);
nand U9227 (N_9227,N_878,N_2298);
nor U9228 (N_9228,N_210,N_4041);
nor U9229 (N_9229,N_4850,N_2655);
or U9230 (N_9230,N_1023,N_4032);
xor U9231 (N_9231,N_3619,N_2690);
or U9232 (N_9232,N_4107,N_4502);
or U9233 (N_9233,N_2488,N_989);
or U9234 (N_9234,N_3936,N_3260);
and U9235 (N_9235,N_4310,N_3335);
nand U9236 (N_9236,N_2246,N_1417);
or U9237 (N_9237,N_1369,N_4538);
xor U9238 (N_9238,N_3347,N_3722);
or U9239 (N_9239,N_3528,N_3047);
nor U9240 (N_9240,N_3254,N_2320);
nand U9241 (N_9241,N_3816,N_2844);
or U9242 (N_9242,N_417,N_2282);
nand U9243 (N_9243,N_1770,N_1128);
and U9244 (N_9244,N_3038,N_4927);
and U9245 (N_9245,N_2457,N_2225);
nand U9246 (N_9246,N_4328,N_1780);
nor U9247 (N_9247,N_223,N_613);
and U9248 (N_9248,N_1258,N_659);
or U9249 (N_9249,N_1141,N_87);
nand U9250 (N_9250,N_4320,N_1564);
nor U9251 (N_9251,N_1333,N_579);
nand U9252 (N_9252,N_4851,N_3749);
nand U9253 (N_9253,N_3001,N_67);
and U9254 (N_9254,N_2240,N_2647);
and U9255 (N_9255,N_3291,N_995);
nor U9256 (N_9256,N_4413,N_235);
nand U9257 (N_9257,N_4533,N_3821);
and U9258 (N_9258,N_4598,N_1403);
or U9259 (N_9259,N_4130,N_720);
xor U9260 (N_9260,N_3788,N_806);
nand U9261 (N_9261,N_3100,N_3866);
and U9262 (N_9262,N_4463,N_554);
and U9263 (N_9263,N_1198,N_4575);
and U9264 (N_9264,N_1842,N_3820);
and U9265 (N_9265,N_119,N_1291);
and U9266 (N_9266,N_1619,N_309);
and U9267 (N_9267,N_839,N_3772);
or U9268 (N_9268,N_737,N_1528);
nor U9269 (N_9269,N_2622,N_2842);
nand U9270 (N_9270,N_4931,N_2284);
xnor U9271 (N_9271,N_486,N_3609);
nor U9272 (N_9272,N_2283,N_1865);
and U9273 (N_9273,N_365,N_290);
nor U9274 (N_9274,N_4097,N_2445);
nor U9275 (N_9275,N_2653,N_3404);
or U9276 (N_9276,N_3707,N_610);
nor U9277 (N_9277,N_774,N_4774);
and U9278 (N_9278,N_930,N_3214);
or U9279 (N_9279,N_3763,N_2270);
xor U9280 (N_9280,N_1198,N_3984);
nand U9281 (N_9281,N_3337,N_2502);
nand U9282 (N_9282,N_4870,N_1458);
or U9283 (N_9283,N_4780,N_765);
and U9284 (N_9284,N_4419,N_608);
nand U9285 (N_9285,N_2337,N_676);
and U9286 (N_9286,N_1328,N_1256);
nor U9287 (N_9287,N_922,N_1346);
xnor U9288 (N_9288,N_4778,N_440);
nor U9289 (N_9289,N_2382,N_3698);
nand U9290 (N_9290,N_1038,N_2856);
nand U9291 (N_9291,N_554,N_1803);
and U9292 (N_9292,N_4817,N_2469);
nand U9293 (N_9293,N_3111,N_1027);
nand U9294 (N_9294,N_2399,N_4773);
nand U9295 (N_9295,N_2501,N_4242);
and U9296 (N_9296,N_2186,N_1707);
nor U9297 (N_9297,N_410,N_4945);
nand U9298 (N_9298,N_1682,N_754);
nand U9299 (N_9299,N_4503,N_2331);
and U9300 (N_9300,N_61,N_2036);
nand U9301 (N_9301,N_1620,N_1025);
or U9302 (N_9302,N_2996,N_4830);
nand U9303 (N_9303,N_1173,N_1027);
and U9304 (N_9304,N_1506,N_3503);
or U9305 (N_9305,N_3174,N_2167);
or U9306 (N_9306,N_1634,N_2419);
or U9307 (N_9307,N_3624,N_405);
nand U9308 (N_9308,N_3903,N_2330);
nor U9309 (N_9309,N_2052,N_1687);
or U9310 (N_9310,N_2772,N_3913);
and U9311 (N_9311,N_3790,N_4209);
nand U9312 (N_9312,N_4702,N_4873);
nand U9313 (N_9313,N_1447,N_3254);
xnor U9314 (N_9314,N_3803,N_4009);
and U9315 (N_9315,N_847,N_1492);
and U9316 (N_9316,N_4924,N_3619);
or U9317 (N_9317,N_3775,N_4007);
and U9318 (N_9318,N_1382,N_4772);
or U9319 (N_9319,N_782,N_3046);
and U9320 (N_9320,N_4659,N_2156);
and U9321 (N_9321,N_3634,N_2986);
or U9322 (N_9322,N_2286,N_1182);
or U9323 (N_9323,N_3200,N_3382);
xnor U9324 (N_9324,N_2663,N_25);
and U9325 (N_9325,N_550,N_207);
and U9326 (N_9326,N_377,N_3377);
xor U9327 (N_9327,N_2515,N_4317);
and U9328 (N_9328,N_2560,N_947);
nand U9329 (N_9329,N_3470,N_4753);
nor U9330 (N_9330,N_2360,N_306);
nand U9331 (N_9331,N_2579,N_827);
or U9332 (N_9332,N_1420,N_1024);
nor U9333 (N_9333,N_3385,N_2102);
and U9334 (N_9334,N_4262,N_1180);
and U9335 (N_9335,N_2123,N_1346);
nand U9336 (N_9336,N_4605,N_1695);
or U9337 (N_9337,N_3124,N_1586);
nand U9338 (N_9338,N_1729,N_3744);
nand U9339 (N_9339,N_4438,N_3236);
and U9340 (N_9340,N_1617,N_4943);
or U9341 (N_9341,N_2471,N_666);
and U9342 (N_9342,N_4880,N_3914);
nor U9343 (N_9343,N_1746,N_4797);
nor U9344 (N_9344,N_3717,N_2763);
or U9345 (N_9345,N_4426,N_1538);
or U9346 (N_9346,N_2892,N_1341);
nand U9347 (N_9347,N_1276,N_4017);
and U9348 (N_9348,N_27,N_4547);
and U9349 (N_9349,N_1954,N_599);
xor U9350 (N_9350,N_1817,N_4024);
and U9351 (N_9351,N_3517,N_708);
and U9352 (N_9352,N_657,N_517);
nand U9353 (N_9353,N_2761,N_470);
and U9354 (N_9354,N_2390,N_122);
nand U9355 (N_9355,N_2783,N_2262);
nor U9356 (N_9356,N_4480,N_4645);
and U9357 (N_9357,N_2532,N_2299);
and U9358 (N_9358,N_870,N_4938);
or U9359 (N_9359,N_39,N_3880);
xnor U9360 (N_9360,N_3086,N_4534);
nor U9361 (N_9361,N_3460,N_1191);
xor U9362 (N_9362,N_1742,N_1374);
and U9363 (N_9363,N_1524,N_2317);
or U9364 (N_9364,N_2182,N_4713);
and U9365 (N_9365,N_2050,N_3702);
and U9366 (N_9366,N_139,N_1416);
and U9367 (N_9367,N_2538,N_1358);
nor U9368 (N_9368,N_1447,N_2613);
and U9369 (N_9369,N_2406,N_2968);
or U9370 (N_9370,N_4046,N_1580);
nand U9371 (N_9371,N_3081,N_478);
nand U9372 (N_9372,N_2318,N_3600);
or U9373 (N_9373,N_1932,N_4228);
nand U9374 (N_9374,N_2461,N_4366);
and U9375 (N_9375,N_4866,N_3535);
and U9376 (N_9376,N_1530,N_1199);
nand U9377 (N_9377,N_4554,N_3324);
and U9378 (N_9378,N_4465,N_2005);
and U9379 (N_9379,N_4256,N_1558);
or U9380 (N_9380,N_2891,N_2919);
nor U9381 (N_9381,N_1789,N_989);
and U9382 (N_9382,N_3886,N_4361);
nand U9383 (N_9383,N_1734,N_649);
nor U9384 (N_9384,N_4380,N_850);
and U9385 (N_9385,N_4859,N_2490);
or U9386 (N_9386,N_2212,N_2249);
nor U9387 (N_9387,N_4978,N_635);
nand U9388 (N_9388,N_1507,N_911);
nor U9389 (N_9389,N_3018,N_3274);
nand U9390 (N_9390,N_2197,N_971);
xor U9391 (N_9391,N_1031,N_4187);
nand U9392 (N_9392,N_3620,N_750);
nor U9393 (N_9393,N_3700,N_259);
nor U9394 (N_9394,N_4639,N_4134);
nor U9395 (N_9395,N_1711,N_1158);
xor U9396 (N_9396,N_634,N_3372);
and U9397 (N_9397,N_757,N_4719);
nand U9398 (N_9398,N_1538,N_79);
and U9399 (N_9399,N_2440,N_326);
and U9400 (N_9400,N_4138,N_2202);
or U9401 (N_9401,N_2126,N_2023);
nor U9402 (N_9402,N_392,N_1236);
or U9403 (N_9403,N_2461,N_1537);
or U9404 (N_9404,N_856,N_4336);
nor U9405 (N_9405,N_2619,N_3276);
nand U9406 (N_9406,N_3963,N_1132);
nor U9407 (N_9407,N_2122,N_683);
xnor U9408 (N_9408,N_3466,N_949);
and U9409 (N_9409,N_4020,N_1031);
xor U9410 (N_9410,N_1546,N_1788);
and U9411 (N_9411,N_2230,N_949);
nor U9412 (N_9412,N_2730,N_3404);
and U9413 (N_9413,N_3224,N_4941);
and U9414 (N_9414,N_4825,N_2747);
and U9415 (N_9415,N_3967,N_1274);
nor U9416 (N_9416,N_2707,N_960);
nor U9417 (N_9417,N_2386,N_2926);
or U9418 (N_9418,N_375,N_1235);
nand U9419 (N_9419,N_27,N_4012);
nor U9420 (N_9420,N_3200,N_3712);
nand U9421 (N_9421,N_1788,N_771);
nor U9422 (N_9422,N_587,N_4653);
nand U9423 (N_9423,N_2725,N_1226);
nor U9424 (N_9424,N_2185,N_1993);
xor U9425 (N_9425,N_1628,N_2714);
or U9426 (N_9426,N_3419,N_2593);
nand U9427 (N_9427,N_3679,N_3172);
nand U9428 (N_9428,N_2760,N_3510);
or U9429 (N_9429,N_618,N_3327);
nand U9430 (N_9430,N_4742,N_4109);
nor U9431 (N_9431,N_532,N_3947);
and U9432 (N_9432,N_2985,N_3207);
and U9433 (N_9433,N_454,N_2655);
nand U9434 (N_9434,N_2169,N_3515);
and U9435 (N_9435,N_1303,N_1509);
nand U9436 (N_9436,N_1544,N_3099);
and U9437 (N_9437,N_3897,N_4313);
nand U9438 (N_9438,N_4952,N_2365);
nor U9439 (N_9439,N_4606,N_2681);
nor U9440 (N_9440,N_2412,N_4377);
or U9441 (N_9441,N_1060,N_694);
or U9442 (N_9442,N_4217,N_4778);
xor U9443 (N_9443,N_4567,N_2499);
nand U9444 (N_9444,N_3378,N_3879);
and U9445 (N_9445,N_1430,N_3828);
and U9446 (N_9446,N_2658,N_4790);
nor U9447 (N_9447,N_1619,N_2329);
nor U9448 (N_9448,N_4827,N_2839);
nor U9449 (N_9449,N_4929,N_3244);
nor U9450 (N_9450,N_2148,N_834);
and U9451 (N_9451,N_3606,N_1659);
or U9452 (N_9452,N_2471,N_260);
nand U9453 (N_9453,N_4885,N_2429);
nor U9454 (N_9454,N_1342,N_111);
nor U9455 (N_9455,N_4343,N_4948);
nor U9456 (N_9456,N_927,N_3251);
nor U9457 (N_9457,N_2449,N_2710);
and U9458 (N_9458,N_3533,N_562);
nand U9459 (N_9459,N_633,N_1353);
nand U9460 (N_9460,N_1202,N_3547);
nand U9461 (N_9461,N_2488,N_927);
xnor U9462 (N_9462,N_4281,N_2693);
and U9463 (N_9463,N_1731,N_1755);
nand U9464 (N_9464,N_3239,N_4610);
and U9465 (N_9465,N_2215,N_930);
nor U9466 (N_9466,N_625,N_2518);
or U9467 (N_9467,N_4678,N_2985);
nand U9468 (N_9468,N_4366,N_278);
or U9469 (N_9469,N_3367,N_4465);
nand U9470 (N_9470,N_1853,N_2654);
xor U9471 (N_9471,N_1768,N_4624);
and U9472 (N_9472,N_3452,N_4296);
nor U9473 (N_9473,N_1316,N_4103);
nand U9474 (N_9474,N_2777,N_2345);
nand U9475 (N_9475,N_4887,N_1614);
nand U9476 (N_9476,N_4384,N_1697);
or U9477 (N_9477,N_2041,N_2706);
or U9478 (N_9478,N_3298,N_578);
nand U9479 (N_9479,N_1040,N_221);
and U9480 (N_9480,N_4746,N_2643);
xor U9481 (N_9481,N_4812,N_4992);
nand U9482 (N_9482,N_3816,N_276);
nand U9483 (N_9483,N_551,N_4418);
nor U9484 (N_9484,N_3445,N_348);
or U9485 (N_9485,N_3481,N_3203);
nor U9486 (N_9486,N_2699,N_1324);
or U9487 (N_9487,N_271,N_2327);
nand U9488 (N_9488,N_3881,N_1836);
or U9489 (N_9489,N_1668,N_3370);
or U9490 (N_9490,N_2236,N_4361);
nor U9491 (N_9491,N_1451,N_4484);
xnor U9492 (N_9492,N_1346,N_4953);
xnor U9493 (N_9493,N_2105,N_1872);
nand U9494 (N_9494,N_3893,N_3190);
and U9495 (N_9495,N_4954,N_2519);
and U9496 (N_9496,N_109,N_589);
and U9497 (N_9497,N_4132,N_1661);
xor U9498 (N_9498,N_2858,N_3374);
nor U9499 (N_9499,N_4307,N_3010);
or U9500 (N_9500,N_3819,N_2898);
nor U9501 (N_9501,N_254,N_1992);
or U9502 (N_9502,N_4741,N_1073);
nand U9503 (N_9503,N_863,N_67);
and U9504 (N_9504,N_1144,N_3968);
and U9505 (N_9505,N_4652,N_3229);
or U9506 (N_9506,N_1531,N_3114);
xor U9507 (N_9507,N_1001,N_3566);
nand U9508 (N_9508,N_2740,N_4013);
nor U9509 (N_9509,N_1297,N_4509);
and U9510 (N_9510,N_636,N_715);
or U9511 (N_9511,N_4386,N_1469);
xnor U9512 (N_9512,N_714,N_3300);
nand U9513 (N_9513,N_427,N_3253);
and U9514 (N_9514,N_3927,N_3550);
or U9515 (N_9515,N_4640,N_404);
xnor U9516 (N_9516,N_403,N_4756);
xor U9517 (N_9517,N_976,N_4031);
and U9518 (N_9518,N_4248,N_1482);
or U9519 (N_9519,N_2983,N_4079);
nor U9520 (N_9520,N_1382,N_3595);
nand U9521 (N_9521,N_68,N_3621);
and U9522 (N_9522,N_4248,N_1962);
nor U9523 (N_9523,N_186,N_4303);
xnor U9524 (N_9524,N_485,N_2907);
and U9525 (N_9525,N_3487,N_886);
and U9526 (N_9526,N_560,N_3080);
nor U9527 (N_9527,N_4067,N_468);
or U9528 (N_9528,N_4641,N_4682);
and U9529 (N_9529,N_4859,N_3161);
or U9530 (N_9530,N_50,N_708);
or U9531 (N_9531,N_4389,N_2104);
and U9532 (N_9532,N_2255,N_4063);
and U9533 (N_9533,N_482,N_3476);
nor U9534 (N_9534,N_3674,N_4217);
nand U9535 (N_9535,N_4766,N_3359);
nand U9536 (N_9536,N_4592,N_3807);
nor U9537 (N_9537,N_3926,N_3588);
or U9538 (N_9538,N_2593,N_3774);
or U9539 (N_9539,N_4238,N_3408);
or U9540 (N_9540,N_873,N_2414);
nand U9541 (N_9541,N_991,N_2601);
and U9542 (N_9542,N_1104,N_4084);
or U9543 (N_9543,N_4828,N_1410);
nor U9544 (N_9544,N_166,N_4421);
nand U9545 (N_9545,N_108,N_3095);
or U9546 (N_9546,N_3474,N_1956);
and U9547 (N_9547,N_172,N_4398);
or U9548 (N_9548,N_3876,N_3805);
or U9549 (N_9549,N_957,N_2112);
or U9550 (N_9550,N_1723,N_2885);
or U9551 (N_9551,N_4448,N_944);
nand U9552 (N_9552,N_1332,N_1897);
nor U9553 (N_9553,N_4464,N_348);
or U9554 (N_9554,N_260,N_4560);
nand U9555 (N_9555,N_3062,N_2984);
nand U9556 (N_9556,N_768,N_3608);
nor U9557 (N_9557,N_3246,N_1483);
xor U9558 (N_9558,N_2737,N_572);
nor U9559 (N_9559,N_1631,N_1917);
or U9560 (N_9560,N_1888,N_1096);
nor U9561 (N_9561,N_2518,N_3757);
or U9562 (N_9562,N_2426,N_1628);
nor U9563 (N_9563,N_2499,N_195);
nor U9564 (N_9564,N_881,N_3263);
or U9565 (N_9565,N_3131,N_1215);
nor U9566 (N_9566,N_3102,N_4112);
or U9567 (N_9567,N_1696,N_2008);
and U9568 (N_9568,N_2649,N_2070);
or U9569 (N_9569,N_733,N_2986);
nor U9570 (N_9570,N_1627,N_1440);
or U9571 (N_9571,N_2694,N_2984);
nor U9572 (N_9572,N_4268,N_2952);
or U9573 (N_9573,N_2033,N_3775);
or U9574 (N_9574,N_176,N_3764);
or U9575 (N_9575,N_1555,N_1035);
nor U9576 (N_9576,N_2580,N_3458);
nand U9577 (N_9577,N_4147,N_4135);
nand U9578 (N_9578,N_1705,N_352);
xor U9579 (N_9579,N_1130,N_1431);
nor U9580 (N_9580,N_1696,N_3442);
nand U9581 (N_9581,N_685,N_3775);
and U9582 (N_9582,N_901,N_4467);
or U9583 (N_9583,N_3691,N_1761);
and U9584 (N_9584,N_236,N_4691);
and U9585 (N_9585,N_4757,N_2089);
nor U9586 (N_9586,N_2273,N_2988);
and U9587 (N_9587,N_2624,N_2860);
xnor U9588 (N_9588,N_1591,N_2594);
and U9589 (N_9589,N_668,N_412);
nand U9590 (N_9590,N_4273,N_2766);
nor U9591 (N_9591,N_3662,N_831);
nor U9592 (N_9592,N_857,N_303);
xnor U9593 (N_9593,N_146,N_2211);
nor U9594 (N_9594,N_3108,N_609);
nand U9595 (N_9595,N_505,N_685);
nor U9596 (N_9596,N_709,N_883);
or U9597 (N_9597,N_43,N_3464);
and U9598 (N_9598,N_2535,N_185);
or U9599 (N_9599,N_819,N_4331);
and U9600 (N_9600,N_4088,N_20);
or U9601 (N_9601,N_4110,N_728);
or U9602 (N_9602,N_2173,N_1027);
nand U9603 (N_9603,N_1560,N_3471);
and U9604 (N_9604,N_1646,N_4770);
xnor U9605 (N_9605,N_1478,N_4619);
and U9606 (N_9606,N_3682,N_3308);
nor U9607 (N_9607,N_413,N_1317);
nand U9608 (N_9608,N_4648,N_538);
nand U9609 (N_9609,N_1821,N_997);
and U9610 (N_9610,N_1245,N_4172);
nor U9611 (N_9611,N_376,N_848);
nand U9612 (N_9612,N_2322,N_655);
nand U9613 (N_9613,N_4276,N_535);
nand U9614 (N_9614,N_65,N_4659);
nor U9615 (N_9615,N_3370,N_890);
and U9616 (N_9616,N_2728,N_3631);
or U9617 (N_9617,N_2344,N_1075);
or U9618 (N_9618,N_810,N_3897);
and U9619 (N_9619,N_4614,N_1383);
or U9620 (N_9620,N_2659,N_734);
and U9621 (N_9621,N_2833,N_2105);
nor U9622 (N_9622,N_4200,N_2525);
and U9623 (N_9623,N_1430,N_507);
xnor U9624 (N_9624,N_387,N_3708);
or U9625 (N_9625,N_4738,N_2267);
xnor U9626 (N_9626,N_4591,N_4216);
or U9627 (N_9627,N_2656,N_2004);
or U9628 (N_9628,N_490,N_2684);
or U9629 (N_9629,N_4388,N_4884);
and U9630 (N_9630,N_835,N_2197);
xor U9631 (N_9631,N_36,N_2113);
nor U9632 (N_9632,N_774,N_2240);
and U9633 (N_9633,N_3577,N_3982);
or U9634 (N_9634,N_1319,N_4606);
nand U9635 (N_9635,N_805,N_4506);
xor U9636 (N_9636,N_1558,N_1118);
and U9637 (N_9637,N_3543,N_4853);
and U9638 (N_9638,N_2559,N_3342);
or U9639 (N_9639,N_2730,N_2326);
xor U9640 (N_9640,N_1965,N_3214);
and U9641 (N_9641,N_609,N_1193);
and U9642 (N_9642,N_1945,N_149);
xor U9643 (N_9643,N_969,N_806);
nand U9644 (N_9644,N_2885,N_283);
nand U9645 (N_9645,N_3985,N_55);
and U9646 (N_9646,N_2323,N_3996);
or U9647 (N_9647,N_2960,N_1499);
xnor U9648 (N_9648,N_3693,N_824);
nand U9649 (N_9649,N_1958,N_1263);
nor U9650 (N_9650,N_4333,N_3887);
nor U9651 (N_9651,N_1756,N_3499);
and U9652 (N_9652,N_1036,N_1837);
and U9653 (N_9653,N_3673,N_914);
and U9654 (N_9654,N_354,N_3320);
xnor U9655 (N_9655,N_2631,N_2153);
and U9656 (N_9656,N_4090,N_2494);
or U9657 (N_9657,N_117,N_1722);
or U9658 (N_9658,N_2930,N_1950);
and U9659 (N_9659,N_2465,N_3505);
or U9660 (N_9660,N_35,N_4570);
and U9661 (N_9661,N_512,N_4169);
nand U9662 (N_9662,N_4968,N_2071);
nor U9663 (N_9663,N_4606,N_4948);
or U9664 (N_9664,N_3807,N_2482);
nor U9665 (N_9665,N_3697,N_1126);
nand U9666 (N_9666,N_2069,N_3863);
or U9667 (N_9667,N_938,N_2659);
nand U9668 (N_9668,N_3291,N_3369);
or U9669 (N_9669,N_1873,N_3375);
and U9670 (N_9670,N_548,N_3895);
nor U9671 (N_9671,N_4550,N_3238);
and U9672 (N_9672,N_2844,N_1489);
and U9673 (N_9673,N_324,N_876);
and U9674 (N_9674,N_4063,N_4007);
and U9675 (N_9675,N_1280,N_316);
nand U9676 (N_9676,N_4264,N_2323);
xnor U9677 (N_9677,N_3557,N_3539);
nor U9678 (N_9678,N_50,N_1472);
nand U9679 (N_9679,N_1275,N_2637);
and U9680 (N_9680,N_2350,N_1859);
and U9681 (N_9681,N_446,N_4178);
nand U9682 (N_9682,N_1246,N_3649);
nand U9683 (N_9683,N_4256,N_4553);
or U9684 (N_9684,N_2348,N_3509);
nand U9685 (N_9685,N_1289,N_1114);
nand U9686 (N_9686,N_2804,N_2785);
nand U9687 (N_9687,N_200,N_3280);
and U9688 (N_9688,N_3446,N_2964);
and U9689 (N_9689,N_16,N_671);
and U9690 (N_9690,N_762,N_1898);
nand U9691 (N_9691,N_184,N_4075);
nor U9692 (N_9692,N_2630,N_3222);
or U9693 (N_9693,N_3644,N_4813);
or U9694 (N_9694,N_2166,N_1393);
and U9695 (N_9695,N_283,N_3494);
and U9696 (N_9696,N_2481,N_1989);
or U9697 (N_9697,N_259,N_4779);
xor U9698 (N_9698,N_4237,N_3726);
or U9699 (N_9699,N_3973,N_4574);
nor U9700 (N_9700,N_4518,N_1360);
nor U9701 (N_9701,N_4325,N_4250);
or U9702 (N_9702,N_4617,N_1365);
and U9703 (N_9703,N_2433,N_1958);
nand U9704 (N_9704,N_2482,N_1479);
nor U9705 (N_9705,N_4455,N_3319);
or U9706 (N_9706,N_4956,N_2360);
nand U9707 (N_9707,N_4451,N_4083);
or U9708 (N_9708,N_3085,N_2135);
nor U9709 (N_9709,N_3465,N_3278);
nand U9710 (N_9710,N_2403,N_1681);
and U9711 (N_9711,N_4080,N_1557);
or U9712 (N_9712,N_1531,N_3091);
and U9713 (N_9713,N_4848,N_1860);
and U9714 (N_9714,N_3138,N_2089);
xnor U9715 (N_9715,N_2092,N_579);
nand U9716 (N_9716,N_3016,N_4285);
and U9717 (N_9717,N_3074,N_4316);
xnor U9718 (N_9718,N_1504,N_2222);
and U9719 (N_9719,N_317,N_1135);
nand U9720 (N_9720,N_4131,N_3041);
nand U9721 (N_9721,N_4696,N_1167);
or U9722 (N_9722,N_3401,N_3400);
or U9723 (N_9723,N_3811,N_1821);
nand U9724 (N_9724,N_2136,N_2311);
nand U9725 (N_9725,N_3112,N_1578);
nor U9726 (N_9726,N_2965,N_4020);
or U9727 (N_9727,N_4802,N_3565);
nor U9728 (N_9728,N_4602,N_2484);
nand U9729 (N_9729,N_2130,N_86);
and U9730 (N_9730,N_906,N_1719);
nor U9731 (N_9731,N_3858,N_2839);
or U9732 (N_9732,N_2753,N_3753);
nor U9733 (N_9733,N_3770,N_4501);
nand U9734 (N_9734,N_3535,N_2843);
or U9735 (N_9735,N_2597,N_2122);
nand U9736 (N_9736,N_1138,N_2042);
nand U9737 (N_9737,N_2274,N_2687);
nand U9738 (N_9738,N_4101,N_4674);
or U9739 (N_9739,N_3351,N_3464);
nand U9740 (N_9740,N_2835,N_1262);
nor U9741 (N_9741,N_3697,N_2254);
and U9742 (N_9742,N_2944,N_2059);
xnor U9743 (N_9743,N_4291,N_178);
nor U9744 (N_9744,N_53,N_2471);
nor U9745 (N_9745,N_4913,N_3793);
nor U9746 (N_9746,N_562,N_4086);
and U9747 (N_9747,N_3364,N_3292);
nand U9748 (N_9748,N_1098,N_3732);
nand U9749 (N_9749,N_279,N_2103);
nand U9750 (N_9750,N_1188,N_3094);
nor U9751 (N_9751,N_4014,N_3298);
or U9752 (N_9752,N_136,N_1466);
nand U9753 (N_9753,N_378,N_3878);
and U9754 (N_9754,N_2722,N_1932);
and U9755 (N_9755,N_3987,N_676);
nand U9756 (N_9756,N_1552,N_3485);
nand U9757 (N_9757,N_2456,N_3891);
nand U9758 (N_9758,N_1379,N_1066);
xnor U9759 (N_9759,N_2644,N_2997);
and U9760 (N_9760,N_4856,N_3017);
nand U9761 (N_9761,N_2738,N_4744);
and U9762 (N_9762,N_995,N_1889);
nor U9763 (N_9763,N_4211,N_4257);
nor U9764 (N_9764,N_3889,N_2271);
nor U9765 (N_9765,N_2722,N_3087);
or U9766 (N_9766,N_1464,N_1052);
or U9767 (N_9767,N_3910,N_3219);
nor U9768 (N_9768,N_3603,N_3534);
and U9769 (N_9769,N_3407,N_2835);
and U9770 (N_9770,N_4110,N_2531);
nand U9771 (N_9771,N_1642,N_2325);
or U9772 (N_9772,N_844,N_2476);
nor U9773 (N_9773,N_481,N_928);
or U9774 (N_9774,N_2749,N_1136);
and U9775 (N_9775,N_3965,N_4187);
xor U9776 (N_9776,N_356,N_2197);
xnor U9777 (N_9777,N_1471,N_1463);
or U9778 (N_9778,N_192,N_2379);
nand U9779 (N_9779,N_1018,N_4722);
and U9780 (N_9780,N_3574,N_48);
xor U9781 (N_9781,N_4704,N_1308);
nor U9782 (N_9782,N_2591,N_4238);
nand U9783 (N_9783,N_1627,N_1679);
nand U9784 (N_9784,N_2404,N_912);
and U9785 (N_9785,N_4976,N_85);
nand U9786 (N_9786,N_3930,N_1612);
or U9787 (N_9787,N_2585,N_2237);
or U9788 (N_9788,N_1502,N_2430);
xnor U9789 (N_9789,N_2778,N_3517);
xnor U9790 (N_9790,N_3483,N_4294);
or U9791 (N_9791,N_1043,N_2686);
and U9792 (N_9792,N_4028,N_978);
nand U9793 (N_9793,N_2577,N_2089);
and U9794 (N_9794,N_3078,N_1728);
or U9795 (N_9795,N_3263,N_3168);
nand U9796 (N_9796,N_346,N_3285);
nand U9797 (N_9797,N_3384,N_1334);
xnor U9798 (N_9798,N_4995,N_3333);
and U9799 (N_9799,N_3913,N_4838);
nand U9800 (N_9800,N_3309,N_1238);
or U9801 (N_9801,N_989,N_4809);
and U9802 (N_9802,N_4708,N_4838);
xnor U9803 (N_9803,N_4551,N_4262);
nand U9804 (N_9804,N_3151,N_1345);
or U9805 (N_9805,N_153,N_434);
xnor U9806 (N_9806,N_189,N_222);
xor U9807 (N_9807,N_2796,N_143);
nor U9808 (N_9808,N_3743,N_3389);
nand U9809 (N_9809,N_4385,N_4478);
nand U9810 (N_9810,N_2299,N_1901);
and U9811 (N_9811,N_3460,N_4586);
nor U9812 (N_9812,N_127,N_4336);
and U9813 (N_9813,N_3195,N_3804);
and U9814 (N_9814,N_1955,N_4035);
and U9815 (N_9815,N_2232,N_300);
and U9816 (N_9816,N_226,N_2102);
xor U9817 (N_9817,N_3672,N_3218);
and U9818 (N_9818,N_4394,N_1308);
or U9819 (N_9819,N_4457,N_2698);
or U9820 (N_9820,N_3254,N_1459);
or U9821 (N_9821,N_2689,N_4974);
or U9822 (N_9822,N_2274,N_2018);
and U9823 (N_9823,N_3306,N_583);
and U9824 (N_9824,N_1570,N_4308);
nor U9825 (N_9825,N_3162,N_2301);
nor U9826 (N_9826,N_3701,N_4919);
or U9827 (N_9827,N_2353,N_397);
nor U9828 (N_9828,N_87,N_4051);
and U9829 (N_9829,N_977,N_1979);
xnor U9830 (N_9830,N_1586,N_1165);
nand U9831 (N_9831,N_1412,N_552);
nor U9832 (N_9832,N_778,N_1395);
or U9833 (N_9833,N_4604,N_1027);
and U9834 (N_9834,N_3224,N_1645);
nand U9835 (N_9835,N_4343,N_2429);
nor U9836 (N_9836,N_3186,N_2271);
and U9837 (N_9837,N_4682,N_3519);
nor U9838 (N_9838,N_3672,N_4295);
nand U9839 (N_9839,N_3992,N_194);
or U9840 (N_9840,N_4750,N_1424);
nand U9841 (N_9841,N_485,N_3185);
xor U9842 (N_9842,N_1722,N_3369);
or U9843 (N_9843,N_1655,N_4114);
xnor U9844 (N_9844,N_3056,N_2922);
nor U9845 (N_9845,N_752,N_903);
and U9846 (N_9846,N_561,N_1056);
nor U9847 (N_9847,N_3639,N_3839);
nor U9848 (N_9848,N_4079,N_2081);
and U9849 (N_9849,N_1806,N_4074);
and U9850 (N_9850,N_1584,N_2101);
nor U9851 (N_9851,N_1859,N_4277);
nor U9852 (N_9852,N_431,N_641);
and U9853 (N_9853,N_3070,N_1098);
or U9854 (N_9854,N_3381,N_520);
or U9855 (N_9855,N_3176,N_3331);
xor U9856 (N_9856,N_1449,N_2225);
and U9857 (N_9857,N_3859,N_342);
nand U9858 (N_9858,N_3612,N_2184);
nor U9859 (N_9859,N_1028,N_3532);
and U9860 (N_9860,N_2205,N_1107);
xnor U9861 (N_9861,N_4197,N_1932);
nand U9862 (N_9862,N_417,N_1786);
or U9863 (N_9863,N_4073,N_4187);
and U9864 (N_9864,N_1102,N_2183);
nand U9865 (N_9865,N_2584,N_1332);
nor U9866 (N_9866,N_4012,N_3809);
or U9867 (N_9867,N_2338,N_633);
nand U9868 (N_9868,N_2862,N_4973);
nor U9869 (N_9869,N_3922,N_1845);
or U9870 (N_9870,N_1213,N_2083);
xor U9871 (N_9871,N_3565,N_4396);
and U9872 (N_9872,N_4295,N_4654);
or U9873 (N_9873,N_1364,N_2181);
nor U9874 (N_9874,N_36,N_2362);
xor U9875 (N_9875,N_375,N_4598);
nand U9876 (N_9876,N_1496,N_4530);
nand U9877 (N_9877,N_1381,N_4477);
or U9878 (N_9878,N_2092,N_3497);
nand U9879 (N_9879,N_4128,N_2217);
nand U9880 (N_9880,N_532,N_38);
nand U9881 (N_9881,N_1831,N_155);
or U9882 (N_9882,N_3010,N_3964);
nand U9883 (N_9883,N_1588,N_4188);
or U9884 (N_9884,N_2969,N_4374);
or U9885 (N_9885,N_3336,N_1035);
nor U9886 (N_9886,N_2046,N_2072);
and U9887 (N_9887,N_4990,N_1511);
nor U9888 (N_9888,N_1129,N_3381);
or U9889 (N_9889,N_4044,N_132);
nand U9890 (N_9890,N_3759,N_1861);
and U9891 (N_9891,N_4994,N_3272);
nor U9892 (N_9892,N_4710,N_3142);
or U9893 (N_9893,N_2549,N_2654);
and U9894 (N_9894,N_4455,N_1119);
and U9895 (N_9895,N_2789,N_4229);
or U9896 (N_9896,N_708,N_2130);
nor U9897 (N_9897,N_1299,N_893);
or U9898 (N_9898,N_2731,N_2875);
nor U9899 (N_9899,N_2215,N_1622);
nor U9900 (N_9900,N_4545,N_2988);
and U9901 (N_9901,N_2350,N_1681);
nand U9902 (N_9902,N_4923,N_3962);
nor U9903 (N_9903,N_2393,N_2297);
xnor U9904 (N_9904,N_3829,N_827);
and U9905 (N_9905,N_3226,N_2463);
or U9906 (N_9906,N_1637,N_4858);
and U9907 (N_9907,N_3103,N_2015);
and U9908 (N_9908,N_1105,N_3922);
and U9909 (N_9909,N_3107,N_4730);
or U9910 (N_9910,N_4264,N_2317);
nand U9911 (N_9911,N_3285,N_2043);
xnor U9912 (N_9912,N_433,N_3589);
xor U9913 (N_9913,N_3482,N_130);
nor U9914 (N_9914,N_529,N_2770);
nand U9915 (N_9915,N_3933,N_4609);
nor U9916 (N_9916,N_1655,N_4447);
nor U9917 (N_9917,N_1026,N_4658);
xor U9918 (N_9918,N_3859,N_2448);
nor U9919 (N_9919,N_4589,N_3807);
and U9920 (N_9920,N_3805,N_4304);
nor U9921 (N_9921,N_3910,N_2650);
nand U9922 (N_9922,N_3005,N_2835);
xor U9923 (N_9923,N_2543,N_3976);
and U9924 (N_9924,N_4485,N_4530);
and U9925 (N_9925,N_1287,N_3649);
or U9926 (N_9926,N_1577,N_4581);
or U9927 (N_9927,N_1009,N_1543);
or U9928 (N_9928,N_1781,N_1031);
nand U9929 (N_9929,N_2605,N_3707);
or U9930 (N_9930,N_1224,N_1473);
nor U9931 (N_9931,N_1592,N_853);
nand U9932 (N_9932,N_1232,N_1979);
nor U9933 (N_9933,N_363,N_1633);
xnor U9934 (N_9934,N_420,N_1373);
or U9935 (N_9935,N_491,N_2031);
nand U9936 (N_9936,N_4824,N_2593);
nand U9937 (N_9937,N_636,N_2161);
nor U9938 (N_9938,N_3961,N_2774);
nand U9939 (N_9939,N_1392,N_790);
or U9940 (N_9940,N_3088,N_4889);
and U9941 (N_9941,N_1669,N_2219);
nand U9942 (N_9942,N_3848,N_1458);
or U9943 (N_9943,N_2133,N_4059);
and U9944 (N_9944,N_4214,N_995);
or U9945 (N_9945,N_1273,N_4997);
nand U9946 (N_9946,N_1206,N_2174);
or U9947 (N_9947,N_1080,N_586);
or U9948 (N_9948,N_4938,N_897);
nand U9949 (N_9949,N_1877,N_3842);
and U9950 (N_9950,N_231,N_1299);
and U9951 (N_9951,N_4857,N_1432);
nor U9952 (N_9952,N_114,N_2112);
nand U9953 (N_9953,N_3778,N_4362);
and U9954 (N_9954,N_3716,N_4125);
nor U9955 (N_9955,N_2879,N_2833);
or U9956 (N_9956,N_1194,N_3245);
nand U9957 (N_9957,N_4684,N_4121);
and U9958 (N_9958,N_1577,N_1653);
or U9959 (N_9959,N_4211,N_4805);
or U9960 (N_9960,N_2612,N_3397);
and U9961 (N_9961,N_4541,N_4673);
nor U9962 (N_9962,N_4695,N_864);
xor U9963 (N_9963,N_3285,N_360);
nand U9964 (N_9964,N_312,N_1084);
nor U9965 (N_9965,N_4939,N_222);
or U9966 (N_9966,N_1186,N_3610);
nor U9967 (N_9967,N_3454,N_107);
or U9968 (N_9968,N_2181,N_2913);
or U9969 (N_9969,N_347,N_2162);
xor U9970 (N_9970,N_1373,N_3548);
and U9971 (N_9971,N_586,N_3757);
and U9972 (N_9972,N_4913,N_4102);
nand U9973 (N_9973,N_848,N_355);
and U9974 (N_9974,N_1308,N_3388);
nor U9975 (N_9975,N_4556,N_3942);
xor U9976 (N_9976,N_1566,N_4286);
xnor U9977 (N_9977,N_4639,N_3098);
nand U9978 (N_9978,N_3917,N_3014);
nand U9979 (N_9979,N_1996,N_922);
nand U9980 (N_9980,N_3590,N_1859);
xnor U9981 (N_9981,N_2622,N_2436);
nor U9982 (N_9982,N_2141,N_2703);
or U9983 (N_9983,N_4309,N_3996);
and U9984 (N_9984,N_1921,N_3297);
nor U9985 (N_9985,N_51,N_3067);
nor U9986 (N_9986,N_4950,N_3962);
or U9987 (N_9987,N_15,N_1678);
nand U9988 (N_9988,N_2706,N_3145);
nor U9989 (N_9989,N_2917,N_3220);
or U9990 (N_9990,N_3138,N_2826);
and U9991 (N_9991,N_3014,N_320);
and U9992 (N_9992,N_3001,N_4671);
xor U9993 (N_9993,N_3009,N_4347);
or U9994 (N_9994,N_2704,N_1819);
or U9995 (N_9995,N_3408,N_4477);
or U9996 (N_9996,N_2948,N_4636);
xnor U9997 (N_9997,N_1106,N_1571);
and U9998 (N_9998,N_1285,N_3313);
nor U9999 (N_9999,N_473,N_235);
or U10000 (N_10000,N_5416,N_8087);
nor U10001 (N_10001,N_7265,N_5478);
or U10002 (N_10002,N_7529,N_7532);
xnor U10003 (N_10003,N_5870,N_7995);
nor U10004 (N_10004,N_7562,N_7494);
nand U10005 (N_10005,N_7343,N_5538);
xnor U10006 (N_10006,N_6929,N_7695);
nand U10007 (N_10007,N_5394,N_7415);
and U10008 (N_10008,N_8336,N_5088);
xor U10009 (N_10009,N_7476,N_5085);
nor U10010 (N_10010,N_8757,N_9224);
nor U10011 (N_10011,N_9949,N_8086);
nor U10012 (N_10012,N_7635,N_8775);
nor U10013 (N_10013,N_7647,N_7353);
nand U10014 (N_10014,N_5931,N_8293);
xor U10015 (N_10015,N_8463,N_6387);
xnor U10016 (N_10016,N_7675,N_7161);
nor U10017 (N_10017,N_7637,N_6550);
or U10018 (N_10018,N_7214,N_6925);
or U10019 (N_10019,N_5695,N_5632);
nand U10020 (N_10020,N_7766,N_8445);
and U10021 (N_10021,N_8203,N_9380);
nor U10022 (N_10022,N_6760,N_5249);
nor U10023 (N_10023,N_8827,N_8172);
or U10024 (N_10024,N_9447,N_9132);
or U10025 (N_10025,N_8930,N_5516);
and U10026 (N_10026,N_8672,N_5823);
nor U10027 (N_10027,N_5841,N_5649);
nor U10028 (N_10028,N_9106,N_5990);
xor U10029 (N_10029,N_8936,N_7734);
nand U10030 (N_10030,N_7979,N_6032);
nor U10031 (N_10031,N_8297,N_7765);
and U10032 (N_10032,N_7318,N_9461);
and U10033 (N_10033,N_9620,N_7609);
xor U10034 (N_10034,N_5889,N_6307);
and U10035 (N_10035,N_5878,N_8423);
or U10036 (N_10036,N_6084,N_7806);
nand U10037 (N_10037,N_7571,N_9173);
nor U10038 (N_10038,N_7955,N_5701);
nand U10039 (N_10039,N_8374,N_9963);
nor U10040 (N_10040,N_6858,N_8130);
xor U10041 (N_10041,N_8019,N_6682);
or U10042 (N_10042,N_5869,N_8529);
and U10043 (N_10043,N_8716,N_8359);
nor U10044 (N_10044,N_5945,N_5329);
nor U10045 (N_10045,N_5156,N_9752);
and U10046 (N_10046,N_9467,N_8266);
xnor U10047 (N_10047,N_6904,N_6822);
or U10048 (N_10048,N_5722,N_8344);
nor U10049 (N_10049,N_7491,N_6060);
nor U10050 (N_10050,N_9408,N_7338);
nand U10051 (N_10051,N_5831,N_8058);
or U10052 (N_10052,N_8243,N_5832);
or U10053 (N_10053,N_5456,N_9144);
nor U10054 (N_10054,N_7266,N_7255);
xnor U10055 (N_10055,N_7431,N_6248);
nor U10056 (N_10056,N_5699,N_8235);
or U10057 (N_10057,N_9974,N_5983);
nor U10058 (N_10058,N_6305,N_8139);
xnor U10059 (N_10059,N_6848,N_9354);
xnor U10060 (N_10060,N_9785,N_5370);
nor U10061 (N_10061,N_6978,N_8953);
nor U10062 (N_10062,N_7309,N_7194);
nand U10063 (N_10063,N_5477,N_5365);
nand U10064 (N_10064,N_6277,N_9057);
nand U10065 (N_10065,N_9210,N_8586);
or U10066 (N_10066,N_5586,N_7282);
and U10067 (N_10067,N_6488,N_8316);
nor U10068 (N_10068,N_5187,N_8310);
and U10069 (N_10069,N_8785,N_9585);
nor U10070 (N_10070,N_7911,N_5308);
nand U10071 (N_10071,N_6231,N_8343);
xor U10072 (N_10072,N_5042,N_5549);
or U10073 (N_10073,N_5497,N_6385);
or U10074 (N_10074,N_6404,N_9778);
and U10075 (N_10075,N_6532,N_9232);
and U10076 (N_10076,N_5279,N_9377);
and U10077 (N_10077,N_9270,N_7404);
nand U10078 (N_10078,N_9693,N_6196);
nor U10079 (N_10079,N_9172,N_8789);
nor U10080 (N_10080,N_9061,N_9250);
or U10081 (N_10081,N_8431,N_7264);
and U10082 (N_10082,N_9962,N_9274);
nor U10083 (N_10083,N_8324,N_9715);
nand U10084 (N_10084,N_8962,N_8511);
nor U10085 (N_10085,N_5916,N_5114);
nand U10086 (N_10086,N_7681,N_9947);
nand U10087 (N_10087,N_7783,N_5648);
nand U10088 (N_10088,N_7200,N_7542);
nand U10089 (N_10089,N_9049,N_5979);
nand U10090 (N_10090,N_7463,N_8915);
nor U10091 (N_10091,N_5471,N_5524);
nor U10092 (N_10092,N_5882,N_5509);
nand U10093 (N_10093,N_9235,N_6308);
or U10094 (N_10094,N_6371,N_6734);
xnor U10095 (N_10095,N_8003,N_8864);
or U10096 (N_10096,N_5034,N_5215);
xor U10097 (N_10097,N_7201,N_8302);
or U10098 (N_10098,N_5025,N_6664);
and U10099 (N_10099,N_7894,N_7380);
nor U10100 (N_10100,N_8528,N_7367);
xnor U10101 (N_10101,N_5313,N_6045);
and U10102 (N_10102,N_9737,N_9100);
or U10103 (N_10103,N_7347,N_5977);
nand U10104 (N_10104,N_5418,N_5715);
or U10105 (N_10105,N_8972,N_7888);
nand U10106 (N_10106,N_8661,N_9112);
or U10107 (N_10107,N_5071,N_5432);
nand U10108 (N_10108,N_9148,N_8066);
and U10109 (N_10109,N_9951,N_5667);
or U10110 (N_10110,N_5324,N_8729);
nand U10111 (N_10111,N_7379,N_5559);
or U10112 (N_10112,N_5158,N_9720);
and U10113 (N_10113,N_5295,N_9293);
and U10114 (N_10114,N_8387,N_8487);
or U10115 (N_10115,N_8613,N_7611);
or U10116 (N_10116,N_5293,N_8121);
and U10117 (N_10117,N_9137,N_8014);
or U10118 (N_10118,N_8060,N_5792);
xnor U10119 (N_10119,N_8724,N_9941);
or U10120 (N_10120,N_6028,N_6101);
and U10121 (N_10121,N_7554,N_8308);
nor U10122 (N_10122,N_7396,N_9826);
and U10123 (N_10123,N_6518,N_6033);
nor U10124 (N_10124,N_5198,N_6436);
or U10125 (N_10125,N_5556,N_6278);
or U10126 (N_10126,N_8568,N_7411);
nand U10127 (N_10127,N_9272,N_5590);
nor U10128 (N_10128,N_8170,N_9560);
or U10129 (N_10129,N_6506,N_8550);
xnor U10130 (N_10130,N_6762,N_8726);
xnor U10131 (N_10131,N_8645,N_7285);
nand U10132 (N_10132,N_7076,N_6431);
and U10133 (N_10133,N_9739,N_7622);
and U10134 (N_10134,N_7909,N_6411);
nand U10135 (N_10135,N_5510,N_7508);
xnor U10136 (N_10136,N_5018,N_6031);
and U10137 (N_10137,N_9557,N_8195);
nand U10138 (N_10138,N_6208,N_7493);
or U10139 (N_10139,N_8345,N_8559);
nor U10140 (N_10140,N_8774,N_9413);
and U10141 (N_10141,N_9656,N_8328);
nand U10142 (N_10142,N_7213,N_9959);
and U10143 (N_10143,N_6568,N_5589);
nand U10144 (N_10144,N_8975,N_5696);
and U10145 (N_10145,N_8959,N_5472);
xor U10146 (N_10146,N_8960,N_6146);
or U10147 (N_10147,N_5875,N_9625);
or U10148 (N_10148,N_6928,N_9289);
nor U10149 (N_10149,N_7921,N_5218);
nor U10150 (N_10150,N_8725,N_8231);
or U10151 (N_10151,N_5512,N_9328);
and U10152 (N_10152,N_8080,N_6519);
nor U10153 (N_10153,N_8106,N_8630);
nand U10154 (N_10154,N_9165,N_5747);
or U10155 (N_10155,N_7925,N_6464);
nor U10156 (N_10156,N_6498,N_6093);
nor U10157 (N_10157,N_5132,N_7427);
nor U10158 (N_10158,N_8268,N_7312);
nand U10159 (N_10159,N_9008,N_5397);
or U10160 (N_10160,N_8815,N_6451);
nand U10161 (N_10161,N_7078,N_7124);
or U10162 (N_10162,N_5730,N_8094);
nand U10163 (N_10163,N_8224,N_8867);
nor U10164 (N_10164,N_8833,N_7277);
and U10165 (N_10165,N_5453,N_7940);
and U10166 (N_10166,N_7485,N_7149);
or U10167 (N_10167,N_9842,N_6956);
or U10168 (N_10168,N_5656,N_7503);
and U10169 (N_10169,N_6441,N_9318);
nand U10170 (N_10170,N_6918,N_8841);
and U10171 (N_10171,N_8180,N_8322);
or U10172 (N_10172,N_8033,N_5716);
and U10173 (N_10173,N_9174,N_9127);
or U10174 (N_10174,N_8746,N_6180);
nand U10175 (N_10175,N_6794,N_5450);
nor U10176 (N_10176,N_9020,N_8146);
nand U10177 (N_10177,N_8593,N_9643);
or U10178 (N_10178,N_9637,N_8194);
and U10179 (N_10179,N_8444,N_8872);
or U10180 (N_10180,N_6748,N_9357);
and U10181 (N_10181,N_6399,N_9138);
and U10182 (N_10182,N_5281,N_5443);
and U10183 (N_10183,N_8028,N_6742);
and U10184 (N_10184,N_8545,N_8142);
nor U10185 (N_10185,N_8440,N_9624);
nor U10186 (N_10186,N_6966,N_8587);
nor U10187 (N_10187,N_7119,N_5751);
nand U10188 (N_10188,N_9911,N_8256);
nor U10189 (N_10189,N_5974,N_5988);
nand U10190 (N_10190,N_8191,N_7794);
or U10191 (N_10191,N_9308,N_9079);
or U10192 (N_10192,N_9869,N_9655);
nor U10193 (N_10193,N_8780,N_5410);
nand U10194 (N_10194,N_8184,N_7280);
nor U10195 (N_10195,N_9830,N_8114);
nand U10196 (N_10196,N_9683,N_7398);
nor U10197 (N_10197,N_9341,N_6988);
and U10198 (N_10198,N_6573,N_8212);
nand U10199 (N_10199,N_6138,N_7292);
or U10200 (N_10200,N_6288,N_8213);
nand U10201 (N_10201,N_7307,N_5464);
or U10202 (N_10202,N_5953,N_8307);
nor U10203 (N_10203,N_6214,N_9012);
or U10204 (N_10204,N_8326,N_7707);
nor U10205 (N_10205,N_5822,N_6998);
or U10206 (N_10206,N_8435,N_7646);
or U10207 (N_10207,N_8412,N_5372);
nor U10208 (N_10208,N_8311,N_6166);
nor U10209 (N_10209,N_9086,N_9381);
or U10210 (N_10210,N_8886,N_5790);
or U10211 (N_10211,N_9511,N_5588);
and U10212 (N_10212,N_6738,N_7448);
xor U10213 (N_10213,N_6358,N_9847);
and U10214 (N_10214,N_7570,N_9829);
xor U10215 (N_10215,N_5054,N_6425);
and U10216 (N_10216,N_6100,N_9298);
nor U10217 (N_10217,N_8022,N_6336);
nor U10218 (N_10218,N_5045,N_6434);
nor U10219 (N_10219,N_8032,N_7024);
or U10220 (N_10220,N_9595,N_9769);
or U10221 (N_10221,N_8116,N_5725);
nor U10222 (N_10222,N_9969,N_6206);
or U10223 (N_10223,N_9915,N_8134);
nand U10224 (N_10224,N_5234,N_9777);
nand U10225 (N_10225,N_8946,N_5617);
or U10226 (N_10226,N_7949,N_9553);
or U10227 (N_10227,N_6598,N_6781);
and U10228 (N_10228,N_8874,N_8442);
and U10229 (N_10229,N_6144,N_5024);
and U10230 (N_10230,N_8222,N_5735);
nor U10231 (N_10231,N_5845,N_6261);
and U10232 (N_10232,N_5333,N_9406);
xnor U10233 (N_10233,N_6731,N_8834);
nor U10234 (N_10234,N_6798,N_9288);
and U10235 (N_10235,N_5669,N_9464);
nand U10236 (N_10236,N_8734,N_8402);
and U10237 (N_10237,N_8095,N_7043);
and U10238 (N_10238,N_9848,N_5741);
nand U10239 (N_10239,N_8736,N_6744);
and U10240 (N_10240,N_7417,N_9577);
nor U10241 (N_10241,N_5978,N_8609);
nor U10242 (N_10242,N_6194,N_8051);
nand U10243 (N_10243,N_5660,N_7030);
nand U10244 (N_10244,N_8039,N_5886);
nand U10245 (N_10245,N_9796,N_5206);
nand U10246 (N_10246,N_8031,N_8395);
xor U10247 (N_10247,N_9741,N_7501);
or U10248 (N_10248,N_8935,N_9054);
or U10249 (N_10249,N_7403,N_9260);
or U10250 (N_10250,N_7163,N_9729);
or U10251 (N_10251,N_5278,N_8457);
nand U10252 (N_10252,N_7199,N_5193);
nor U10253 (N_10253,N_7833,N_9918);
and U10254 (N_10254,N_5448,N_7091);
or U10255 (N_10255,N_7120,N_6068);
xor U10256 (N_10256,N_7770,N_5221);
and U10257 (N_10257,N_6330,N_7639);
xor U10258 (N_10258,N_9980,N_7295);
nand U10259 (N_10259,N_9208,N_9305);
nand U10260 (N_10260,N_7405,N_5186);
nor U10261 (N_10261,N_6792,N_7581);
nand U10262 (N_10262,N_7327,N_6125);
xnor U10263 (N_10263,N_9822,N_9714);
nand U10264 (N_10264,N_7364,N_6927);
or U10265 (N_10265,N_9122,N_9835);
or U10266 (N_10266,N_9823,N_9297);
nor U10267 (N_10267,N_6478,N_7289);
or U10268 (N_10268,N_9202,N_6538);
nand U10269 (N_10269,N_5361,N_8223);
nand U10270 (N_10270,N_6723,N_7769);
nor U10271 (N_10271,N_7942,N_5619);
or U10272 (N_10272,N_8965,N_6793);
and U10273 (N_10273,N_9561,N_5343);
nand U10274 (N_10274,N_5754,N_7222);
or U10275 (N_10275,N_8763,N_7775);
or U10276 (N_10276,N_6656,N_5010);
and U10277 (N_10277,N_6765,N_8770);
nand U10278 (N_10278,N_9030,N_7310);
or U10279 (N_10279,N_9244,N_8073);
or U10280 (N_10280,N_6235,N_8955);
or U10281 (N_10281,N_5943,N_6730);
nor U10282 (N_10282,N_9209,N_8688);
nand U10283 (N_10283,N_5251,N_8744);
or U10284 (N_10284,N_7479,N_9649);
xor U10285 (N_10285,N_5314,N_8629);
nor U10286 (N_10286,N_7230,N_6761);
xnor U10287 (N_10287,N_9178,N_7469);
or U10288 (N_10288,N_7226,N_8931);
and U10289 (N_10289,N_9458,N_7477);
or U10290 (N_10290,N_9105,N_7710);
or U10291 (N_10291,N_8853,N_7095);
or U10292 (N_10292,N_9103,N_8105);
and U10293 (N_10293,N_5801,N_7514);
nor U10294 (N_10294,N_6572,N_6565);
and U10295 (N_10295,N_9440,N_9364);
nand U10296 (N_10296,N_7492,N_9880);
nand U10297 (N_10297,N_7385,N_8888);
xnor U10298 (N_10298,N_5220,N_6771);
and U10299 (N_10299,N_9253,N_5828);
nor U10300 (N_10300,N_9038,N_7607);
nor U10301 (N_10301,N_7610,N_6139);
nand U10302 (N_10302,N_5993,N_9587);
or U10303 (N_10303,N_6768,N_8475);
and U10304 (N_10304,N_7966,N_8173);
and U10305 (N_10305,N_6361,N_6696);
and U10306 (N_10306,N_9230,N_8221);
nand U10307 (N_10307,N_6666,N_7679);
and U10308 (N_10308,N_8706,N_7100);
nand U10309 (N_10309,N_7473,N_7549);
or U10310 (N_10310,N_5561,N_7767);
nor U10311 (N_10311,N_8216,N_8786);
nor U10312 (N_10312,N_5315,N_7598);
and U10313 (N_10313,N_6800,N_9372);
and U10314 (N_10314,N_7480,N_9363);
xnor U10315 (N_10315,N_5697,N_5047);
nor U10316 (N_10316,N_8535,N_6735);
or U10317 (N_10317,N_9727,N_9700);
nor U10318 (N_10318,N_5655,N_6926);
or U10319 (N_10319,N_9039,N_8971);
xor U10320 (N_10320,N_9825,N_5140);
and U10321 (N_10321,N_9286,N_5066);
nand U10322 (N_10322,N_8875,N_5224);
nand U10323 (N_10323,N_5640,N_7158);
nor U10324 (N_10324,N_9586,N_9043);
or U10325 (N_10325,N_8378,N_6609);
xor U10326 (N_10326,N_7730,N_9107);
or U10327 (N_10327,N_9499,N_5082);
nor U10328 (N_10328,N_6611,N_8265);
xor U10329 (N_10329,N_8468,N_9939);
or U10330 (N_10330,N_7962,N_8742);
and U10331 (N_10331,N_5992,N_8649);
or U10332 (N_10332,N_5355,N_8490);
xor U10333 (N_10333,N_7743,N_9688);
xnor U10334 (N_10334,N_6680,N_6616);
nor U10335 (N_10335,N_5166,N_7634);
xor U10336 (N_10336,N_9011,N_6945);
nor U10337 (N_10337,N_8560,N_8079);
and U10338 (N_10338,N_7442,N_7764);
nor U10339 (N_10339,N_9125,N_9453);
nand U10340 (N_10340,N_9021,N_5767);
nand U10341 (N_10341,N_7657,N_5188);
xnor U10342 (N_10342,N_5233,N_8509);
nand U10343 (N_10343,N_7854,N_6037);
nor U10344 (N_10344,N_6165,N_9075);
nand U10345 (N_10345,N_7300,N_5217);
nor U10346 (N_10346,N_6462,N_9110);
or U10347 (N_10347,N_7333,N_9696);
or U10348 (N_10348,N_5543,N_6246);
nand U10349 (N_10349,N_8289,N_7920);
or U10350 (N_10350,N_7875,N_5069);
or U10351 (N_10351,N_5661,N_5731);
and U10352 (N_10352,N_6593,N_8981);
nand U10353 (N_10353,N_7552,N_6564);
and U10354 (N_10354,N_5567,N_8461);
or U10355 (N_10355,N_9887,N_7221);
nand U10356 (N_10356,N_9793,N_6801);
and U10357 (N_10357,N_8694,N_5444);
nor U10358 (N_10358,N_9950,N_8899);
or U10359 (N_10359,N_7850,N_6319);
nand U10360 (N_10360,N_7653,N_6027);
or U10361 (N_10361,N_5710,N_8800);
nand U10362 (N_10362,N_8150,N_6947);
xnor U10363 (N_10363,N_6948,N_6684);
and U10364 (N_10364,N_7516,N_5582);
or U10365 (N_10365,N_9074,N_5548);
xnor U10366 (N_10366,N_8129,N_8466);
or U10367 (N_10367,N_9373,N_7207);
and U10368 (N_10368,N_8835,N_5603);
or U10369 (N_10369,N_7040,N_6547);
nor U10370 (N_10370,N_7899,N_7470);
xor U10371 (N_10371,N_6839,N_7414);
nand U10372 (N_10372,N_5342,N_7615);
nor U10373 (N_10373,N_6296,N_7690);
nor U10374 (N_10374,N_7774,N_9954);
and U10375 (N_10375,N_5998,N_5853);
and U10376 (N_10376,N_6335,N_8348);
nand U10377 (N_10377,N_8104,N_8281);
or U10378 (N_10378,N_9634,N_9243);
nand U10379 (N_10379,N_7540,N_9819);
and U10380 (N_10380,N_8283,N_8558);
xor U10381 (N_10381,N_7902,N_7438);
xor U10382 (N_10382,N_9884,N_8838);
or U10383 (N_10383,N_6900,N_7069);
nand U10384 (N_10384,N_8260,N_6600);
nand U10385 (N_10385,N_5605,N_6698);
nor U10386 (N_10386,N_8227,N_8335);
and U10387 (N_10387,N_7771,N_5176);
or U10388 (N_10388,N_7901,N_9680);
or U10389 (N_10389,N_9588,N_5402);
nor U10390 (N_10390,N_8499,N_8515);
nand U10391 (N_10391,N_9150,N_9261);
xor U10392 (N_10392,N_5636,N_9047);
nor U10393 (N_10393,N_6784,N_7314);
nor U10394 (N_10394,N_7644,N_7686);
or U10395 (N_10395,N_5141,N_9559);
nand U10396 (N_10396,N_8131,N_7410);
nand U10397 (N_10397,N_8561,N_8240);
and U10398 (N_10398,N_9903,N_6683);
nand U10399 (N_10399,N_8452,N_6201);
xor U10400 (N_10400,N_6252,N_9285);
nor U10401 (N_10401,N_9734,N_6154);
nand U10402 (N_10402,N_5824,N_6615);
and U10403 (N_10403,N_5932,N_7271);
nor U10404 (N_10404,N_8088,N_7430);
or U10405 (N_10405,N_6006,N_8148);
nor U10406 (N_10406,N_8948,N_6405);
nand U10407 (N_10407,N_8048,N_9984);
nand U10408 (N_10408,N_6938,N_5608);
or U10409 (N_10409,N_6934,N_9600);
and U10410 (N_10410,N_6646,N_7614);
and U10411 (N_10411,N_8369,N_6675);
or U10412 (N_10412,N_8332,N_6957);
xnor U10413 (N_10413,N_5732,N_8384);
or U10414 (N_10414,N_9761,N_9598);
nand U10415 (N_10415,N_9568,N_5785);
nor U10416 (N_10416,N_8333,N_8507);
nor U10417 (N_10417,N_7071,N_5379);
nand U10418 (N_10418,N_8171,N_6418);
or U10419 (N_10419,N_8846,N_7656);
nand U10420 (N_10420,N_7144,N_6749);
nand U10421 (N_10421,N_8917,N_7796);
nand U10422 (N_10422,N_5191,N_9776);
and U10423 (N_10423,N_5766,N_8421);
and U10424 (N_10424,N_7326,N_9046);
or U10425 (N_10425,N_8364,N_9489);
and U10426 (N_10426,N_7683,N_8027);
or U10427 (N_10427,N_8237,N_5760);
nor U10428 (N_10428,N_5285,N_7084);
xnor U10429 (N_10429,N_7781,N_5687);
or U10430 (N_10430,N_5645,N_7075);
or U10431 (N_10431,N_9311,N_5087);
xnor U10432 (N_10432,N_6013,N_5316);
or U10433 (N_10433,N_5599,N_7887);
nand U10434 (N_10434,N_5266,N_6229);
and U10435 (N_10435,N_6244,N_8665);
nand U10436 (N_10436,N_5486,N_6217);
nor U10437 (N_10437,N_8623,N_7851);
nor U10438 (N_10438,N_9626,N_5147);
nand U10439 (N_10439,N_7424,N_5255);
nand U10440 (N_10440,N_5143,N_6541);
and U10441 (N_10441,N_7591,N_5976);
nor U10442 (N_10442,N_9817,N_7714);
nand U10443 (N_10443,N_9449,N_8933);
nand U10444 (N_10444,N_5523,N_7801);
nand U10445 (N_10445,N_7951,N_7046);
nand U10446 (N_10446,N_7179,N_5435);
or U10447 (N_10447,N_9721,N_5681);
xor U10448 (N_10448,N_7928,N_6979);
and U10449 (N_10449,N_5129,N_7917);
nor U10450 (N_10450,N_7702,N_8866);
and U10451 (N_10451,N_7203,N_9498);
or U10452 (N_10452,N_6222,N_5781);
or U10453 (N_10453,N_6204,N_9438);
xor U10454 (N_10454,N_6141,N_5247);
and U10455 (N_10455,N_5750,N_9758);
nand U10456 (N_10456,N_8493,N_8054);
xor U10457 (N_10457,N_9602,N_8627);
or U10458 (N_10458,N_6840,N_7874);
or U10459 (N_10459,N_7628,N_6112);
nand U10460 (N_10460,N_6704,N_8296);
xnor U10461 (N_10461,N_8084,N_8318);
and U10462 (N_10462,N_5713,N_6525);
and U10463 (N_10463,N_8745,N_5043);
nand U10464 (N_10464,N_8824,N_6827);
and U10465 (N_10465,N_5610,N_6406);
and U10466 (N_10466,N_6409,N_5489);
nand U10467 (N_10467,N_6401,N_9033);
nand U10468 (N_10468,N_6604,N_8602);
and U10469 (N_10469,N_9989,N_9611);
xor U10470 (N_10470,N_9913,N_8233);
and U10471 (N_10471,N_8143,N_5057);
nor U10472 (N_10472,N_5246,N_6607);
nand U10473 (N_10473,N_9581,N_9471);
and U10474 (N_10474,N_8059,N_8840);
and U10475 (N_10475,N_7219,N_7478);
and U10476 (N_10476,N_9468,N_5201);
and U10477 (N_10477,N_8920,N_9827);
nor U10478 (N_10478,N_9436,N_6838);
or U10479 (N_10479,N_6352,N_5294);
xnor U10480 (N_10480,N_8436,N_7777);
and U10481 (N_10481,N_5482,N_7426);
nor U10482 (N_10482,N_5185,N_7356);
nor U10483 (N_10483,N_6211,N_7114);
or U10484 (N_10484,N_6083,N_9325);
nand U10485 (N_10485,N_6536,N_7694);
and U10486 (N_10486,N_9349,N_6443);
nand U10487 (N_10487,N_8247,N_8749);
nand U10488 (N_10488,N_7402,N_6981);
and U10489 (N_10489,N_8455,N_6339);
nor U10490 (N_10490,N_5629,N_8844);
nand U10491 (N_10491,N_8020,N_5683);
nor U10492 (N_10492,N_8347,N_9271);
and U10493 (N_10493,N_5055,N_5578);
nand U10494 (N_10494,N_5458,N_9184);
nor U10495 (N_10495,N_9213,N_9279);
nand U10496 (N_10496,N_9630,N_6514);
and U10497 (N_10497,N_7804,N_5651);
nor U10498 (N_10498,N_8471,N_6935);
or U10499 (N_10499,N_5228,N_6177);
or U10500 (N_10500,N_9537,N_5970);
xnor U10501 (N_10501,N_5376,N_6876);
and U10502 (N_10502,N_7400,N_6483);
nor U10503 (N_10503,N_6057,N_8773);
and U10504 (N_10504,N_7297,N_9723);
nor U10505 (N_10505,N_7423,N_5904);
nor U10506 (N_10506,N_6831,N_6342);
and U10507 (N_10507,N_7969,N_7539);
and U10508 (N_10508,N_9928,N_9348);
nand U10509 (N_10509,N_6531,N_7968);
nor U10510 (N_10510,N_7212,N_6143);
nor U10511 (N_10511,N_7696,N_8622);
and U10512 (N_10512,N_6752,N_6561);
nand U10513 (N_10513,N_7699,N_8783);
or U10514 (N_10514,N_9862,N_8635);
nor U10515 (N_10515,N_9536,N_8366);
nand U10516 (N_10516,N_5480,N_5672);
and U10517 (N_10517,N_8705,N_5070);
nand U10518 (N_10518,N_9525,N_8103);
nor U10519 (N_10519,N_9182,N_5427);
or U10520 (N_10520,N_5783,N_7394);
nand U10521 (N_10521,N_5056,N_5759);
nor U10522 (N_10522,N_9873,N_9569);
and U10523 (N_10523,N_6736,N_9323);
or U10524 (N_10524,N_9385,N_8398);
xor U10525 (N_10525,N_9565,N_5720);
nor U10526 (N_10526,N_8006,N_9035);
nor U10527 (N_10527,N_5929,N_5338);
or U10528 (N_10528,N_8393,N_9302);
nand U10529 (N_10529,N_7597,N_9136);
or U10530 (N_10530,N_8710,N_7990);
nor U10531 (N_10531,N_9425,N_9864);
nor U10532 (N_10532,N_7449,N_8997);
xnor U10533 (N_10533,N_7650,N_9399);
and U10534 (N_10534,N_7872,N_8368);
and U10535 (N_10535,N_8158,N_5462);
nor U10536 (N_10536,N_5866,N_7465);
and U10537 (N_10537,N_6359,N_5226);
or U10538 (N_10538,N_6024,N_7215);
and U10539 (N_10539,N_7234,N_9098);
nand U10540 (N_10540,N_8081,N_6174);
or U10541 (N_10541,N_6987,N_5357);
nand U10542 (N_10542,N_8594,N_8034);
nor U10543 (N_10543,N_7843,N_7531);
and U10544 (N_10544,N_6344,N_5320);
and U10545 (N_10545,N_7316,N_6274);
nand U10546 (N_10546,N_6845,N_7815);
and U10547 (N_10547,N_7257,N_5028);
nor U10548 (N_10548,N_8430,N_8621);
or U10549 (N_10549,N_9840,N_9398);
nand U10550 (N_10550,N_7283,N_8921);
nor U10551 (N_10551,N_7527,N_5814);
nor U10552 (N_10552,N_7056,N_5584);
and U10553 (N_10553,N_8999,N_5504);
and U10554 (N_10554,N_7189,N_6552);
nand U10555 (N_10555,N_9882,N_7982);
and U10556 (N_10556,N_9452,N_9731);
and U10557 (N_10557,N_6787,N_9390);
nor U10558 (N_10558,N_7520,N_5284);
xnor U10559 (N_10559,N_7439,N_9316);
and U10560 (N_10560,N_7620,N_6905);
nand U10561 (N_10561,N_8598,N_9571);
xnor U10562 (N_10562,N_5653,N_6124);
nor U10563 (N_10563,N_8353,N_6426);
or U10564 (N_10564,N_8122,N_6059);
xnor U10565 (N_10565,N_5485,N_8730);
nor U10566 (N_10566,N_5075,N_8244);
nor U10567 (N_10567,N_9483,N_5833);
nor U10568 (N_10568,N_7298,N_9163);
and U10569 (N_10569,N_6468,N_8188);
nor U10570 (N_10570,N_8415,N_6906);
or U10571 (N_10571,N_6895,N_5729);
and U10572 (N_10572,N_5269,N_6652);
or U10573 (N_10573,N_5968,N_5941);
and U10574 (N_10574,N_6559,N_6903);
or U10575 (N_10575,N_9104,N_8182);
or U10576 (N_10576,N_7908,N_9712);
nand U10577 (N_10577,N_6281,N_7228);
and U10578 (N_10578,N_7789,N_9116);
or U10579 (N_10579,N_7079,N_9401);
nand U10580 (N_10580,N_7739,N_5270);
and U10581 (N_10581,N_9687,N_7704);
nand U10582 (N_10582,N_6091,N_5287);
nand U10583 (N_10583,N_6994,N_7337);
xor U10584 (N_10584,N_9804,N_6435);
or U10585 (N_10585,N_7254,N_8477);
nand U10586 (N_10586,N_6467,N_6314);
and U10587 (N_10587,N_7728,N_6757);
or U10588 (N_10588,N_7536,N_6829);
nand U10589 (N_10589,N_9050,N_5368);
or U10590 (N_10590,N_5230,N_5309);
nor U10591 (N_10591,N_8601,N_5110);
nor U10592 (N_10592,N_5242,N_6632);
and U10593 (N_10593,N_8313,N_9494);
and U10594 (N_10594,N_5312,N_7864);
and U10595 (N_10595,N_6875,N_6658);
and U10596 (N_10596,N_9332,N_6164);
nor U10597 (N_10597,N_6290,N_5409);
and U10598 (N_10598,N_6570,N_6188);
xnor U10599 (N_10599,N_7588,N_5074);
xnor U10600 (N_10600,N_7365,N_8990);
nor U10601 (N_10601,N_7374,N_9640);
nor U10602 (N_10602,N_9192,N_8831);
nor U10603 (N_10603,N_6179,N_6679);
nand U10604 (N_10604,N_7059,N_9371);
and U10605 (N_10605,N_8372,N_6931);
nand U10606 (N_10606,N_7814,N_9570);
nand U10607 (N_10607,N_6745,N_7346);
xor U10608 (N_10608,N_7841,N_8044);
and U10609 (N_10609,N_9800,N_6692);
nor U10610 (N_10610,N_5468,N_6973);
nor U10611 (N_10611,N_9916,N_9659);
or U10612 (N_10612,N_6152,N_5810);
and U10613 (N_10613,N_6400,N_5620);
or U10614 (N_10614,N_5288,N_9226);
xor U10615 (N_10615,N_6907,N_7893);
or U10616 (N_10616,N_5483,N_8175);
nand U10617 (N_10617,N_8793,N_8074);
or U10618 (N_10618,N_6944,N_5015);
or U10619 (N_10619,N_6168,N_6087);
xnor U10620 (N_10620,N_6597,N_5890);
or U10621 (N_10621,N_9924,N_8396);
or U10622 (N_10622,N_9416,N_9048);
nand U10623 (N_10623,N_8226,N_7382);
nor U10624 (N_10624,N_8225,N_7583);
nand U10625 (N_10625,N_5614,N_9780);
nand U10626 (N_10626,N_7164,N_9663);
nor U10627 (N_10627,N_5552,N_9526);
nor U10628 (N_10628,N_7308,N_5854);
or U10629 (N_10629,N_7484,N_8036);
and U10630 (N_10630,N_5133,N_6114);
nand U10631 (N_10631,N_8234,N_7421);
nand U10632 (N_10632,N_7007,N_5684);
and U10633 (N_10633,N_9073,N_6148);
nor U10634 (N_10634,N_5262,N_9576);
or U10635 (N_10635,N_7565,N_8963);
and U10636 (N_10636,N_7475,N_5076);
nand U10637 (N_10637,N_7919,N_9324);
or U10638 (N_10638,N_9684,N_7537);
nand U10639 (N_10639,N_8969,N_5857);
nand U10640 (N_10640,N_9351,N_7236);
nor U10641 (N_10641,N_7320,N_7971);
xor U10642 (N_10642,N_7383,N_6688);
or U10643 (N_10643,N_7466,N_8061);
nor U10644 (N_10644,N_5787,N_9019);
and U10645 (N_10645,N_7759,N_7306);
or U10646 (N_10646,N_9402,N_5688);
and U10647 (N_10647,N_6090,N_5802);
nand U10648 (N_10648,N_7999,N_5289);
and U10649 (N_10649,N_8427,N_5300);
and U10650 (N_10650,N_7196,N_7758);
xor U10651 (N_10651,N_5189,N_9200);
xor U10652 (N_10652,N_7904,N_9343);
nand U10653 (N_10653,N_9786,N_7209);
nor U10654 (N_10654,N_7393,N_6799);
and U10655 (N_10655,N_5880,N_9251);
and U10656 (N_10656,N_5146,N_7459);
nand U10657 (N_10657,N_8938,N_8443);
or U10658 (N_10658,N_6029,N_7593);
or U10659 (N_10659,N_8612,N_9249);
nor U10660 (N_10660,N_6304,N_6712);
and U10661 (N_10661,N_9166,N_9881);
and U10662 (N_10662,N_9558,N_7606);
and U10663 (N_10663,N_6779,N_7519);
nor U10664 (N_10664,N_8057,N_7602);
or U10665 (N_10665,N_9459,N_7182);
and U10666 (N_10666,N_8458,N_6834);
or U10667 (N_10667,N_5771,N_7468);
or U10668 (N_10668,N_9930,N_8577);
nand U10669 (N_10669,N_9856,N_8715);
or U10670 (N_10670,N_8514,N_5160);
or U10671 (N_10671,N_6475,N_6967);
nor U10672 (N_10672,N_9344,N_5290);
and U10673 (N_10673,N_8682,N_7773);
or U10674 (N_10674,N_8634,N_9375);
or U10675 (N_10675,N_7102,N_9514);
nand U10676 (N_10676,N_6880,N_8794);
and U10677 (N_10677,N_5306,N_8210);
nor U10678 (N_10678,N_8913,N_8982);
nor U10679 (N_10679,N_7181,N_9518);
nor U10680 (N_10680,N_7827,N_5493);
or U10681 (N_10681,N_9201,N_7397);
nor U10682 (N_10682,N_6109,N_6729);
and U10683 (N_10683,N_6303,N_5291);
and U10684 (N_10684,N_8570,N_7900);
nand U10685 (N_10685,N_8413,N_9146);
nand U10686 (N_10686,N_9010,N_6558);
nand U10687 (N_10687,N_7706,N_7217);
nor U10688 (N_10688,N_9534,N_5535);
or U10689 (N_10689,N_5454,N_5131);
nand U10690 (N_10690,N_6102,N_6841);
nand U10691 (N_10691,N_6224,N_7837);
xor U10692 (N_10692,N_5753,N_9631);
or U10693 (N_10693,N_7997,N_8041);
or U10694 (N_10694,N_8922,N_7287);
xor U10695 (N_10695,N_8470,N_6785);
nand U10696 (N_10696,N_9031,N_5635);
nor U10697 (N_10697,N_9533,N_6094);
and U10698 (N_10698,N_8739,N_6513);
or U10699 (N_10699,N_5261,N_5029);
and U10700 (N_10700,N_8258,N_8015);
and U10701 (N_10701,N_9342,N_9556);
or U10702 (N_10702,N_6471,N_9092);
nand U10703 (N_10703,N_7574,N_5116);
and U10704 (N_10704,N_9259,N_6238);
xor U10705 (N_10705,N_6892,N_5078);
and U10706 (N_10706,N_6693,N_7141);
and U10707 (N_10707,N_8541,N_7334);
nor U10708 (N_10708,N_6321,N_9852);
nand U10709 (N_10709,N_7344,N_9597);
or U10710 (N_10710,N_7268,N_7852);
xor U10711 (N_10711,N_8994,N_8701);
and U10712 (N_10712,N_6654,N_7321);
or U10713 (N_10713,N_7559,N_8788);
nand U10714 (N_10714,N_8976,N_5846);
nor U10715 (N_10715,N_7462,N_7170);
or U10716 (N_10716,N_6445,N_7819);
or U10717 (N_10717,N_9672,N_5745);
nand U10718 (N_10718,N_8607,N_7440);
nand U10719 (N_10719,N_6920,N_6644);
nand U10720 (N_10720,N_6423,N_8397);
nand U10721 (N_10721,N_9088,N_7839);
xnor U10722 (N_10722,N_8685,N_7907);
nor U10723 (N_10723,N_8828,N_9330);
xor U10724 (N_10724,N_5579,N_6601);
nor U10725 (N_10725,N_7756,N_6687);
and U10726 (N_10726,N_9740,N_5473);
nand U10727 (N_10727,N_5638,N_7147);
nand U10728 (N_10728,N_9060,N_5803);
nor U10729 (N_10729,N_8731,N_6285);
nor U10730 (N_10730,N_7446,N_8439);
or U10731 (N_10731,N_8751,N_9410);
xnor U10732 (N_10732,N_8217,N_9563);
nand U10733 (N_10733,N_5881,N_7377);
nand U10734 (N_10734,N_6470,N_7019);
and U10735 (N_10735,N_9133,N_8383);
nand U10736 (N_10736,N_8858,N_6510);
nand U10737 (N_10737,N_9473,N_8923);
or U10738 (N_10738,N_9532,N_8524);
nor U10739 (N_10739,N_9904,N_9068);
and U10740 (N_10740,N_7640,N_9794);
and U10741 (N_10741,N_8494,N_6192);
nor U10742 (N_10742,N_5949,N_5367);
or U10743 (N_10743,N_6887,N_8657);
nor U10744 (N_10744,N_8974,N_9515);
nand U10745 (N_10745,N_9496,N_9053);
nor U10746 (N_10746,N_9177,N_6549);
nand U10747 (N_10747,N_5469,N_5212);
or U10748 (N_10748,N_7031,N_8787);
or U10749 (N_10749,N_9605,N_9488);
or U10750 (N_10750,N_8179,N_5712);
and U10751 (N_10751,N_6954,N_8951);
nor U10752 (N_10752,N_9345,N_6908);
nor U10753 (N_10753,N_9787,N_9240);
nand U10754 (N_10754,N_7453,N_5296);
or U10755 (N_10755,N_7068,N_5818);
and U10756 (N_10756,N_8610,N_8837);
or U10757 (N_10757,N_8943,N_9442);
nor U10758 (N_10758,N_5292,N_6974);
or U10759 (N_10759,N_5484,N_7094);
nor U10760 (N_10760,N_7303,N_8363);
or U10761 (N_10761,N_6457,N_9666);
and U10762 (N_10762,N_8894,N_6873);
nand U10763 (N_10763,N_8530,N_9395);
nor U10764 (N_10764,N_9594,N_7020);
and U10765 (N_10765,N_5236,N_9703);
and U10766 (N_10766,N_6612,N_8686);
nand U10767 (N_10767,N_8270,N_8164);
and U10768 (N_10768,N_5700,N_9193);
or U10769 (N_10769,N_7360,N_5036);
nand U10770 (N_10770,N_5905,N_8377);
or U10771 (N_10771,N_5470,N_7525);
or U10772 (N_10772,N_5374,N_5389);
nand U10773 (N_10773,N_7744,N_5809);
or U10774 (N_10774,N_9891,N_7805);
and U10775 (N_10775,N_5999,N_7244);
and U10776 (N_10776,N_5769,N_7051);
or U10777 (N_10777,N_7433,N_6098);
and U10778 (N_10778,N_5044,N_6630);
or U10779 (N_10779,N_5352,N_6159);
and U10780 (N_10780,N_5004,N_6725);
or U10781 (N_10781,N_6271,N_6324);
nand U10782 (N_10782,N_7080,N_5602);
xnor U10783 (N_10783,N_7472,N_7381);
or U10784 (N_10784,N_5679,N_8910);
nor U10785 (N_10785,N_9109,N_8218);
nor U10786 (N_10786,N_6884,N_8769);
nor U10787 (N_10787,N_5774,N_8389);
nor U10788 (N_10788,N_8619,N_6251);
and U10789 (N_10789,N_5714,N_7856);
nor U10790 (N_10790,N_5237,N_5772);
or U10791 (N_10791,N_7322,N_5817);
or U10792 (N_10792,N_6484,N_7608);
or U10793 (N_10793,N_9327,N_6790);
nand U10794 (N_10794,N_7248,N_5501);
xor U10795 (N_10795,N_6021,N_5159);
and U10796 (N_10796,N_7162,N_7922);
or U10797 (N_10797,N_7787,N_6041);
or U10798 (N_10798,N_9129,N_5184);
nand U10799 (N_10799,N_5690,N_7157);
or U10800 (N_10800,N_8748,N_9225);
or U10801 (N_10801,N_6254,N_8267);
and U10802 (N_10802,N_9616,N_6820);
nor U10803 (N_10803,N_5165,N_5844);
or U10804 (N_10804,N_9195,N_5328);
xnor U10805 (N_10805,N_8305,N_7240);
nand U10806 (N_10806,N_6136,N_7813);
nand U10807 (N_10807,N_8162,N_7032);
or U10808 (N_10808,N_9004,N_9797);
nand U10809 (N_10809,N_7047,N_9067);
or U10810 (N_10810,N_7135,N_9382);
nor U10811 (N_10811,N_7220,N_6171);
or U10812 (N_10812,N_8700,N_6959);
nand U10813 (N_10813,N_6381,N_6313);
or U10814 (N_10814,N_6708,N_8554);
nand U10815 (N_10815,N_6455,N_9407);
or U10816 (N_10816,N_6857,N_6061);
and U10817 (N_10817,N_9159,N_8292);
and U10818 (N_10818,N_6586,N_9728);
or U10819 (N_10819,N_7339,N_7061);
or U10820 (N_10820,N_5299,N_5083);
and U10821 (N_10821,N_9975,N_8573);
and U10822 (N_10822,N_9833,N_8481);
nor U10823 (N_10823,N_6740,N_5008);
nand U10824 (N_10824,N_5001,N_7941);
nor U10825 (N_10825,N_8185,N_9966);
nor U10826 (N_10826,N_8653,N_6527);
and U10827 (N_10827,N_6444,N_8735);
nor U10828 (N_10828,N_8119,N_7972);
or U10829 (N_10829,N_5213,N_8520);
nor U10830 (N_10830,N_8197,N_8264);
xnor U10831 (N_10831,N_6889,N_6701);
nand U10832 (N_10832,N_9519,N_6384);
or U10833 (N_10833,N_7093,N_7830);
and U10834 (N_10834,N_5798,N_8596);
and U10835 (N_10835,N_5694,N_5848);
and U10836 (N_10836,N_5954,N_6039);
and U10837 (N_10837,N_9018,N_6198);
nor U10838 (N_10838,N_7210,N_8024);
or U10839 (N_10839,N_9942,N_7315);
nor U10840 (N_10840,N_9623,N_9065);
or U10841 (N_10841,N_9196,N_8693);
or U10842 (N_10842,N_7541,N_6286);
nor U10843 (N_10843,N_9430,N_5739);
and U10844 (N_10844,N_6207,N_9858);
or U10845 (N_10845,N_8288,N_7953);
nor U10846 (N_10846,N_8380,N_8428);
nand U10847 (N_10847,N_9055,N_5386);
and U10848 (N_10848,N_7252,N_7780);
or U10849 (N_10849,N_9015,N_7530);
or U10850 (N_10850,N_5258,N_9255);
nand U10851 (N_10851,N_8488,N_5495);
nor U10852 (N_10852,N_6050,N_7110);
and U10853 (N_10853,N_5377,N_5899);
and U10854 (N_10854,N_9562,N_7003);
xor U10855 (N_10855,N_6591,N_8654);
and U10856 (N_10856,N_5546,N_6402);
nor U10857 (N_10857,N_6833,N_9495);
nand U10858 (N_10858,N_9698,N_7868);
or U10859 (N_10859,N_7748,N_6496);
nand U10860 (N_10860,N_7954,N_9077);
nand U10861 (N_10861,N_5799,N_5921);
and U10862 (N_10862,N_7669,N_9114);
or U10863 (N_10863,N_7489,N_5898);
and U10864 (N_10864,N_5463,N_5900);
or U10865 (N_10865,N_6940,N_9340);
nor U10866 (N_10866,N_7361,N_8482);
nand U10867 (N_10867,N_6092,N_9062);
nor U10868 (N_10868,N_7857,N_9792);
nand U10869 (N_10869,N_8597,N_5108);
nand U10870 (N_10870,N_5346,N_7260);
xnor U10871 (N_10871,N_5839,N_8885);
nand U10872 (N_10872,N_8123,N_9844);
and U10873 (N_10873,N_7370,N_6504);
and U10874 (N_10874,N_8196,N_7098);
xnor U10875 (N_10875,N_9922,N_8631);
or U10876 (N_10876,N_8198,N_8382);
or U10877 (N_10877,N_6364,N_7171);
and U10878 (N_10878,N_6380,N_5793);
or U10879 (N_10879,N_6117,N_7986);
nor U10880 (N_10880,N_5514,N_5161);
or U10881 (N_10881,N_7677,N_6428);
xor U10882 (N_10882,N_8360,N_7281);
nor U10883 (N_10883,N_8968,N_5304);
or U10884 (N_10884,N_8940,N_5371);
and U10885 (N_10885,N_6719,N_8896);
and U10886 (N_10886,N_6355,N_5518);
or U10887 (N_10887,N_5488,N_8927);
nand U10888 (N_10888,N_5360,N_7858);
and U10889 (N_10889,N_5181,N_9629);
or U10890 (N_10890,N_5476,N_5671);
and U10891 (N_10891,N_6289,N_8284);
nand U10892 (N_10892,N_7099,N_7803);
and U10893 (N_10893,N_9434,N_6422);
or U10894 (N_10894,N_6689,N_6958);
nand U10895 (N_10895,N_5326,N_7458);
nor U10896 (N_10896,N_8892,N_7535);
nor U10897 (N_10897,N_5837,N_9953);
and U10898 (N_10898,N_6969,N_6200);
and U10899 (N_10899,N_8762,N_7961);
and U10900 (N_10900,N_9176,N_9567);
nand U10901 (N_10901,N_9242,N_5946);
and U10902 (N_10902,N_8916,N_5982);
xor U10903 (N_10903,N_5286,N_5390);
and U10904 (N_10904,N_8242,N_7010);
or U10905 (N_10905,N_7505,N_8755);
and U10906 (N_10906,N_5544,N_6249);
nand U10907 (N_10907,N_6879,N_6438);
nor U10908 (N_10908,N_6637,N_7021);
nor U10909 (N_10909,N_7568,N_5689);
nand U10910 (N_10910,N_8459,N_7993);
xor U10911 (N_10911,N_6713,N_8854);
xor U10912 (N_10912,N_6477,N_6351);
nor U10913 (N_10913,N_7797,N_5530);
and U10914 (N_10914,N_7822,N_5691);
nand U10915 (N_10915,N_7988,N_8329);
nand U10916 (N_10916,N_7782,N_7227);
and U10917 (N_10917,N_6678,N_7932);
and U10918 (N_10918,N_8232,N_6132);
nor U10919 (N_10919,N_5175,N_5742);
xnor U10920 (N_10920,N_8450,N_5706);
nor U10921 (N_10921,N_8252,N_7332);
nand U10922 (N_10922,N_9713,N_6493);
nor U10923 (N_10923,N_6913,N_9524);
nand U10924 (N_10924,N_6257,N_7437);
or U10925 (N_10925,N_8381,N_9347);
xor U10926 (N_10926,N_5872,N_8069);
and U10927 (N_10927,N_6982,N_9755);
or U10928 (N_10928,N_5467,N_8907);
nand U10929 (N_10929,N_6474,N_6172);
and U10930 (N_10930,N_6886,N_6999);
or U10931 (N_10931,N_9744,N_8865);
nand U10932 (N_10932,N_6546,N_9905);
or U10933 (N_10933,N_9014,N_8849);
or U10934 (N_10934,N_5933,N_7892);
nor U10935 (N_10935,N_8663,N_5428);
nor U10936 (N_10936,N_6412,N_5081);
nor U10937 (N_10937,N_7945,N_9774);
nand U10938 (N_10938,N_5575,N_9609);
nand U10939 (N_10939,N_9089,N_9066);
xnor U10940 (N_10940,N_5171,N_7420);
nand U10941 (N_10941,N_6458,N_8880);
xnor U10942 (N_10942,N_6427,N_5138);
nand U10943 (N_10943,N_5317,N_8572);
nand U10944 (N_10944,N_6329,N_7626);
nor U10945 (N_10945,N_5303,N_6516);
xnor U10946 (N_10946,N_8479,N_6315);
nand U10947 (N_10947,N_7001,N_8549);
nand U10948 (N_10948,N_9396,N_6273);
nand U10949 (N_10949,N_5644,N_9017);
nand U10950 (N_10950,N_9238,N_8272);
nand U10951 (N_10951,N_8388,N_9169);
and U10952 (N_10952,N_9591,N_7667);
nand U10953 (N_10953,N_5311,N_6796);
xor U10954 (N_10954,N_6508,N_5838);
and U10955 (N_10955,N_7408,N_7861);
nand U10956 (N_10956,N_7447,N_8406);
and U10957 (N_10957,N_6542,N_8053);
nand U10958 (N_10958,N_6530,N_5086);
nor U10959 (N_10959,N_9868,N_6843);
nand U10960 (N_10960,N_9154,N_9523);
xnor U10961 (N_10961,N_8120,N_6183);
nand U10962 (N_10962,N_5035,N_6287);
nor U10963 (N_10963,N_7176,N_9748);
nand U10964 (N_10964,N_6012,N_9427);
nor U10965 (N_10965,N_5536,N_5887);
nand U10966 (N_10966,N_8052,N_7630);
and U10967 (N_10967,N_7106,N_8199);
nand U10968 (N_10968,N_9360,N_8262);
and U10969 (N_10969,N_9513,N_9628);
nand U10970 (N_10970,N_5779,N_7490);
or U10971 (N_10971,N_8967,N_8984);
and U10972 (N_10972,N_8285,N_9228);
or U10973 (N_10973,N_7727,N_6003);
nand U10974 (N_10974,N_9618,N_5940);
or U10975 (N_10975,N_5425,N_5498);
nor U10976 (N_10976,N_5852,N_9064);
or U10977 (N_10977,N_7973,N_7964);
nand U10978 (N_10978,N_9101,N_8924);
nand U10979 (N_10979,N_5922,N_9171);
nand U10980 (N_10980,N_8462,N_8168);
nand U10981 (N_10981,N_7616,N_7167);
and U10982 (N_10982,N_5229,N_5971);
xnor U10983 (N_10983,N_8004,N_6046);
nand U10984 (N_10984,N_9763,N_8096);
and U10985 (N_10985,N_9153,N_9485);
and U10986 (N_10986,N_7757,N_5120);
or U10987 (N_10987,N_5404,N_8998);
xor U10988 (N_10988,N_5235,N_7229);
nor U10989 (N_10989,N_6215,N_6081);
or U10990 (N_10990,N_9199,N_5830);
nor U10991 (N_10991,N_9157,N_6860);
and U10992 (N_10992,N_8802,N_7467);
or U10993 (N_10993,N_8432,N_9044);
nand U10994 (N_10994,N_9221,N_5153);
or U10995 (N_10995,N_7778,N_9529);
nand U10996 (N_10996,N_5437,N_7906);
nand U10997 (N_10997,N_5113,N_9756);
xor U10998 (N_10998,N_6686,N_9789);
or U10999 (N_10999,N_6259,N_9460);
or U11000 (N_11000,N_7599,N_8717);
nand U11001 (N_11001,N_8604,N_5863);
or U11002 (N_11002,N_8050,N_9808);
xor U11003 (N_11003,N_9268,N_8898);
nand U11004 (N_11004,N_7963,N_5157);
nand U11005 (N_11005,N_6078,N_5728);
or U11006 (N_11006,N_7811,N_5666);
nor U11007 (N_11007,N_9875,N_5633);
nor U11008 (N_11008,N_8934,N_6587);
and U11009 (N_11009,N_5918,N_6556);
xor U11010 (N_11010,N_7233,N_5135);
or U11011 (N_11011,N_8767,N_8147);
nor U11012 (N_11012,N_7074,N_7808);
and U11013 (N_11013,N_9475,N_9198);
nand U11014 (N_11014,N_5762,N_9299);
and U11015 (N_11015,N_5913,N_9123);
and U11016 (N_11016,N_5362,N_7726);
and U11017 (N_11017,N_8042,N_6743);
nor U11018 (N_11018,N_8437,N_7576);
nor U11019 (N_11019,N_5023,N_9056);
nand U11020 (N_11020,N_5500,N_8433);
nand U11021 (N_11021,N_8371,N_9967);
or U11022 (N_11022,N_5906,N_6403);
and U11023 (N_11023,N_9411,N_6226);
nor U11024 (N_11024,N_7905,N_8189);
and U11025 (N_11025,N_7567,N_8349);
nor U11026 (N_11026,N_8650,N_6421);
nor U11027 (N_11027,N_5021,N_8002);
or U11028 (N_11028,N_7112,N_9300);
xnor U11029 (N_11029,N_8961,N_8817);
or U11030 (N_11030,N_9331,N_5545);
nand U11031 (N_11031,N_8544,N_9940);
xnor U11032 (N_11032,N_9681,N_6193);
or U11033 (N_11033,N_5915,N_6420);
nand U11034 (N_11034,N_9992,N_6173);
nor U11035 (N_11035,N_9674,N_5616);
and U11036 (N_11036,N_6653,N_9026);
or U11037 (N_11037,N_6720,N_8407);
and U11038 (N_11038,N_9846,N_5583);
nand U11039 (N_11039,N_6219,N_6837);
nor U11040 (N_11040,N_5566,N_5973);
and U11041 (N_11041,N_8109,N_9614);
and U11042 (N_11042,N_8993,N_8241);
or U11043 (N_11043,N_5642,N_7866);
nor U11044 (N_11044,N_7812,N_7261);
nor U11045 (N_11045,N_6733,N_5969);
xor U11046 (N_11046,N_7717,N_6473);
and U11047 (N_11047,N_9134,N_6337);
or U11048 (N_11048,N_9424,N_5248);
xor U11049 (N_11049,N_8778,N_9866);
or U11050 (N_11050,N_6870,N_7688);
nor U11051 (N_11051,N_9162,N_6133);
nand U11052 (N_11052,N_9803,N_5873);
or U11053 (N_11053,N_7641,N_8669);
and U11054 (N_11054,N_8416,N_8043);
and U11055 (N_11055,N_7148,N_8228);
nand U11056 (N_11056,N_6366,N_8643);
nand U11057 (N_11057,N_7014,N_5763);
or U11058 (N_11058,N_9516,N_7474);
or U11059 (N_11059,N_7073,N_8903);
and U11060 (N_11060,N_6022,N_8502);
nor U11061 (N_11061,N_6044,N_8918);
xnor U11062 (N_11062,N_8186,N_8467);
xnor U11063 (N_11063,N_5127,N_7755);
nand U11064 (N_11064,N_5813,N_7601);
nor U11065 (N_11065,N_7832,N_7733);
or U11066 (N_11066,N_8720,N_6863);
xor U11067 (N_11067,N_5253,N_7225);
nand U11068 (N_11068,N_6009,N_8637);
nor U11069 (N_11069,N_7569,N_8441);
or U11070 (N_11070,N_8300,N_8732);
and U11071 (N_11071,N_6603,N_6082);
nand U11072 (N_11072,N_8595,N_8708);
xor U11073 (N_11073,N_9885,N_6617);
nand U11074 (N_11074,N_5939,N_6763);
xor U11075 (N_11075,N_7625,N_7528);
nand U11076 (N_11076,N_8399,N_6578);
nand U11077 (N_11077,N_7224,N_9215);
or U11078 (N_11078,N_5244,N_7121);
and U11079 (N_11079,N_8055,N_6463);
xor U11080 (N_11080,N_6849,N_7590);
nor U11081 (N_11081,N_5506,N_7009);
and U11082 (N_11082,N_9802,N_7204);
and U11083 (N_11083,N_9045,N_8848);
nor U11084 (N_11084,N_6569,N_5912);
nand U11085 (N_11085,N_5795,N_5569);
or U11086 (N_11086,N_7152,N_7253);
nand U11087 (N_11087,N_6638,N_9032);
and U11088 (N_11088,N_9078,N_6312);
nor U11089 (N_11089,N_6777,N_8469);
nand U11090 (N_11090,N_7154,N_8405);
and U11091 (N_11091,N_9615,N_9606);
nand U11092 (N_11092,N_9102,N_7747);
nand U11093 (N_11093,N_5322,N_8334);
and U11094 (N_11094,N_6852,N_5302);
nand U11095 (N_11095,N_5937,N_8618);
nor U11096 (N_11096,N_8711,N_7202);
nor U11097 (N_11097,N_5095,N_6714);
nand U11098 (N_11098,N_8290,N_8832);
nor U11099 (N_11099,N_8257,N_5112);
nand U11100 (N_11100,N_6485,N_8842);
xnor U11101 (N_11101,N_5734,N_5265);
or U11102 (N_11102,N_6023,N_5808);
nand U11103 (N_11103,N_6338,N_8155);
and U11104 (N_11104,N_8000,N_5791);
xor U11105 (N_11105,N_6129,N_8230);
nand U11106 (N_11106,N_8277,N_7435);
nor U11107 (N_11107,N_8187,N_9278);
nand U11108 (N_11108,N_7390,N_6825);
and U11109 (N_11109,N_6461,N_6103);
or U11110 (N_11110,N_8424,N_7720);
or U11111 (N_11111,N_8647,N_7425);
nor U11112 (N_11112,N_9987,N_9543);
nand U11113 (N_11113,N_8491,N_6576);
and U11114 (N_11114,N_6108,N_9502);
nand U11115 (N_11115,N_5891,N_9384);
and U11116 (N_11116,N_5851,N_8531);
nor U11117 (N_11117,N_8996,N_9531);
and U11118 (N_11118,N_5128,N_9717);
xnor U11119 (N_11119,N_5654,N_9472);
nor U11120 (N_11120,N_5094,N_9705);
nor U11121 (N_11121,N_5459,N_7125);
nor U11122 (N_11122,N_7190,N_6705);
or U11123 (N_11123,N_6047,N_5911);
nor U11124 (N_11124,N_6891,N_9287);
nand U11125 (N_11125,N_5172,N_7369);
nand U11126 (N_11126,N_7286,N_7974);
or U11127 (N_11127,N_5124,N_7085);
and U11128 (N_11128,N_8871,N_5321);
nor U11129 (N_11129,N_5996,N_5593);
nand U11130 (N_11130,N_5104,N_6480);
nand U11131 (N_11131,N_5718,N_8820);
or U11132 (N_11132,N_6465,N_5907);
nand U11133 (N_11133,N_6718,N_7551);
nor U11134 (N_11134,N_6002,N_6575);
or U11135 (N_11135,N_8056,N_5490);
or U11136 (N_11136,N_5513,N_9917);
or U11137 (N_11137,N_8689,N_9246);
or U11138 (N_11138,N_9596,N_7487);
nand U11139 (N_11139,N_5405,N_6985);
or U11140 (N_11140,N_9063,N_8255);
and U11141 (N_11141,N_9481,N_7488);
and U11142 (N_11142,N_5664,N_7697);
nand U11143 (N_11143,N_6417,N_7891);
nor U11144 (N_11144,N_8483,N_6276);
nor U11145 (N_11145,N_6454,N_6960);
or U11146 (N_11146,N_8025,N_7471);
nand U11147 (N_11147,N_5491,N_5573);
nand U11148 (N_11148,N_5356,N_8331);
or U11149 (N_11149,N_8484,N_9197);
nor U11150 (N_11150,N_7105,N_8236);
and U11151 (N_11151,N_5177,N_8901);
nor U11152 (N_11152,N_9773,N_8354);
and U11153 (N_11153,N_9386,N_9590);
nor U11154 (N_11154,N_6662,N_6203);
nor U11155 (N_11155,N_8246,N_6645);
xor U11156 (N_11156,N_9592,N_8365);
or U11157 (N_11157,N_5180,N_8149);
or U11158 (N_11158,N_7482,N_7235);
or U11159 (N_11159,N_6717,N_7603);
nand U11160 (N_11160,N_7645,N_8707);
xnor U11161 (N_11161,N_6660,N_7258);
and U11162 (N_11162,N_5446,N_8966);
or U11163 (N_11163,N_8306,N_9653);
nand U11164 (N_11164,N_8426,N_8206);
and U11165 (N_11165,N_6367,N_5400);
nor U11166 (N_11166,N_8989,N_9115);
or U11167 (N_11167,N_7692,N_7927);
nand U11168 (N_11168,N_9708,N_6566);
nand U11169 (N_11169,N_8460,N_6140);
and U11170 (N_11170,N_9108,N_6659);
or U11171 (N_11171,N_7975,N_9874);
nor U11172 (N_11172,N_8527,N_5511);
and U11173 (N_11173,N_7317,N_9952);
nor U11174 (N_11174,N_6491,N_9541);
or U11175 (N_11175,N_8884,N_7090);
nand U11176 (N_11176,N_5197,N_6320);
and U11177 (N_11177,N_9111,N_8097);
and U11178 (N_11178,N_5609,N_5431);
or U11179 (N_11179,N_9432,N_6916);
nor U11180 (N_11180,N_8030,N_8287);
or U11181 (N_11181,N_8771,N_5319);
and U11182 (N_11182,N_7660,N_5692);
and U11183 (N_11183,N_7461,N_9870);
and U11184 (N_11184,N_7175,N_7831);
and U11185 (N_11185,N_6816,N_9899);
and U11186 (N_11186,N_7246,N_8862);
nand U11187 (N_11187,N_8077,N_5987);
xnor U11188 (N_11188,N_5914,N_9042);
and U11189 (N_11189,N_6853,N_8072);
or U11190 (N_11190,N_6529,N_6323);
xnor U11191 (N_11191,N_8692,N_6828);
nand U11192 (N_11192,N_7378,N_9431);
xor U11193 (N_11193,N_7223,N_5520);
nor U11194 (N_11194,N_6951,N_9839);
or U11195 (N_11195,N_6111,N_7724);
xnor U11196 (N_11196,N_5272,N_6489);
nand U11197 (N_11197,N_6011,N_5426);
and U11198 (N_11198,N_9119,N_8132);
and U11199 (N_11199,N_8385,N_9403);
xnor U11200 (N_11200,N_9257,N_6939);
and U11201 (N_11201,N_7802,N_5412);
nand U11202 (N_11202,N_7406,N_5883);
nor U11203 (N_11203,N_7218,N_9772);
or U11204 (N_11204,N_5332,N_5550);
xor U11205 (N_11205,N_9838,N_6065);
nor U11206 (N_11206,N_8680,N_9212);
nand U11207 (N_11207,N_5927,N_8339);
nor U11208 (N_11208,N_5991,N_6353);
xor U11209 (N_11209,N_9006,N_7655);
nand U11210 (N_11210,N_7267,N_7930);
nand U11211 (N_11211,N_6775,N_5892);
and U11212 (N_11212,N_8790,N_8101);
nor U11213 (N_11213,N_8906,N_6515);
and U11214 (N_11214,N_7066,N_7412);
nand U11215 (N_11215,N_9517,N_5677);
nor U11216 (N_11216,N_7810,N_5951);
nor U11217 (N_11217,N_8603,N_6923);
and U11218 (N_11218,N_6000,N_5222);
nor U11219 (N_11219,N_9365,N_9751);
and U11220 (N_11220,N_7273,N_5000);
nor U11221 (N_11221,N_7082,N_7104);
and U11222 (N_11222,N_7809,N_8562);
and U11223 (N_11223,N_5622,N_5037);
xnor U11224 (N_11224,N_5930,N_6668);
nand U11225 (N_11225,N_6150,N_9806);
xor U11226 (N_11226,N_9143,N_6481);
xor U11227 (N_11227,N_7741,N_7048);
xnor U11228 (N_11228,N_8248,N_5183);
and U11229 (N_11229,N_8063,N_9418);
and U11230 (N_11230,N_9538,N_9923);
or U11231 (N_11231,N_5777,N_8589);
xnor U11232 (N_11232,N_8633,N_6376);
and U11233 (N_11233,N_7914,N_5038);
nand U11234 (N_11234,N_5012,N_9009);
or U11235 (N_11235,N_6955,N_6676);
nor U11236 (N_11236,N_8681,N_5053);
nand U11237 (N_11237,N_5440,N_8696);
and U11238 (N_11238,N_9901,N_8250);
or U11239 (N_11239,N_6579,N_5107);
and U11240 (N_11240,N_9315,N_7564);
and U11241 (N_11241,N_9943,N_9771);
nor U11242 (N_11242,N_9971,N_9443);
or U11243 (N_11243,N_7389,N_5200);
nand U11244 (N_11244,N_6691,N_7621);
xnor U11245 (N_11245,N_6256,N_6432);
nor U11246 (N_11246,N_5475,N_5562);
and U11247 (N_11247,N_7008,N_6490);
and U11248 (N_11248,N_6014,N_5541);
and U11249 (N_11249,N_5686,N_8897);
nor U11250 (N_11250,N_8722,N_5474);
nor U11251 (N_11251,N_5553,N_9760);
nand U11252 (N_11252,N_9770,N_7348);
or U11253 (N_11253,N_5540,N_7274);
or U11254 (N_11254,N_6574,N_5935);
xor U11255 (N_11255,N_9836,N_8453);
and U11256 (N_11256,N_9167,N_8615);
nor U11257 (N_11257,N_9414,N_8417);
or U11258 (N_11258,N_8517,N_8280);
nand U11259 (N_11259,N_8273,N_8465);
and U11260 (N_11260,N_7991,N_5909);
nor U11261 (N_11261,N_9539,N_5950);
xnor U11262 (N_11262,N_9564,N_8314);
or U11263 (N_11263,N_6846,N_9809);
nor U11264 (N_11264,N_8505,N_9131);
nand U11265 (N_11265,N_8741,N_9849);
nand U11266 (N_11266,N_6823,N_5105);
xor U11267 (N_11267,N_8401,N_9155);
or U11268 (N_11268,N_5577,N_7793);
nor U11269 (N_11269,N_9376,N_5560);
nand U11270 (N_11270,N_9747,N_7627);
xnor U11271 (N_11271,N_6225,N_8181);
nor U11272 (N_11272,N_6864,N_6922);
nand U11273 (N_11273,N_9183,N_8355);
and U11274 (N_11274,N_8029,N_9781);
and U11275 (N_11275,N_6071,N_8902);
or U11276 (N_11276,N_9582,N_6808);
nor U11277 (N_11277,N_8684,N_7980);
nor U11278 (N_11278,N_7823,N_5051);
nand U11279 (N_11279,N_6162,N_6562);
nor U11280 (N_11280,N_8599,N_8919);
nand U11281 (N_11281,N_9446,N_6128);
nand U11282 (N_11282,N_8229,N_8617);
or U11283 (N_11283,N_9369,N_5148);
and U11284 (N_11284,N_5901,N_5430);
or U11285 (N_11285,N_8418,N_5049);
xor U11286 (N_11286,N_7936,N_8881);
and U11287 (N_11287,N_5145,N_6663);
or U11288 (N_11288,N_8219,N_5721);
nor U11289 (N_11289,N_9575,N_9222);
and U11290 (N_11290,N_6588,N_5986);
nand U11291 (N_11291,N_7842,N_9338);
and U11292 (N_11292,N_5040,N_7915);
nor U11293 (N_11293,N_5994,N_7623);
nor U11294 (N_11294,N_7678,N_9378);
xor U11295 (N_11295,N_6452,N_9356);
nand U11296 (N_11296,N_7455,N_5879);
nor U11297 (N_11297,N_5196,N_7651);
nand U11298 (N_11298,N_9189,N_6472);
nand U11299 (N_11299,N_5563,N_6571);
nand U11300 (N_11300,N_9099,N_9572);
and U11301 (N_11301,N_6049,N_9664);
nor U11302 (N_11302,N_8192,N_8579);
nor U11303 (N_11303,N_6054,N_6522);
nor U11304 (N_11304,N_6390,N_8518);
nand U11305 (N_11305,N_9642,N_8608);
nand U11306 (N_11306,N_6595,N_5429);
nor U11307 (N_11307,N_6517,N_5758);
or U11308 (N_11308,N_5630,N_5850);
nand U11309 (N_11309,N_6062,N_5657);
or U11310 (N_11310,N_8887,N_9912);
nor U11311 (N_11311,N_6230,N_8522);
or U11312 (N_11312,N_7950,N_9258);
or U11313 (N_11313,N_7371,N_8165);
nand U11314 (N_11314,N_7208,N_6309);
and U11315 (N_11315,N_6476,N_7127);
or U11316 (N_11316,N_6992,N_6835);
nand U11317 (N_11317,N_8954,N_5658);
xor U11318 (N_11318,N_9859,N_7504);
nor U11319 (N_11319,N_8215,N_5547);
or U11320 (N_11320,N_5373,N_9976);
nor U11321 (N_11321,N_8480,N_5439);
xor U11322 (N_11322,N_8492,N_6520);
or U11323 (N_11323,N_8782,N_6153);
and U11324 (N_11324,N_5685,N_9633);
or U11325 (N_11325,N_7083,N_5178);
and U11326 (N_11326,N_7057,N_6807);
xnor U11327 (N_11327,N_6085,N_6115);
nor U11328 (N_11328,N_9892,N_8508);
or U11329 (N_11329,N_6501,N_7325);
and U11330 (N_11330,N_5871,N_5856);
and U11331 (N_11331,N_7115,N_6332);
and U11332 (N_11332,N_7604,N_9650);
nor U11333 (N_11333,N_6619,N_5170);
or U11334 (N_11334,N_5122,N_6996);
and U11335 (N_11335,N_7584,N_6099);
or U11336 (N_11336,N_8392,N_5243);
and U11337 (N_11337,N_7958,N_5564);
nor U11338 (N_11338,N_8583,N_5144);
and U11339 (N_11339,N_6694,N_9733);
nand U11340 (N_11340,N_8945,N_5452);
nor U11341 (N_11341,N_6747,N_6016);
nand U11342 (N_11342,N_9051,N_6818);
nor U11343 (N_11343,N_5952,N_8115);
nor U11344 (N_11344,N_9374,N_8220);
xnor U11345 (N_11345,N_5020,N_9180);
or U11346 (N_11346,N_9983,N_6284);
and U11347 (N_11347,N_5908,N_6543);
or U11348 (N_11348,N_5865,N_7873);
or U11349 (N_11349,N_5967,N_9437);
or U11350 (N_11350,N_8911,N_9352);
xnor U11351 (N_11351,N_6810,N_9775);
nor U11352 (N_11352,N_5805,N_9707);
nor U11353 (N_11353,N_8309,N_7238);
or U11354 (N_11354,N_6347,N_7335);
and U11355 (N_11355,N_7524,N_8703);
nor U11356 (N_11356,N_7247,N_5411);
and U11357 (N_11357,N_6859,N_9554);
nand U11358 (N_11358,N_5531,N_6555);
nor U11359 (N_11359,N_8163,N_7160);
nor U11360 (N_11360,N_5621,N_9301);
and U11361 (N_11361,N_9782,N_5707);
nor U11362 (N_11362,N_5307,N_9675);
and U11363 (N_11363,N_6759,N_9646);
nand U11364 (N_11364,N_6241,N_7772);
nor U11365 (N_11365,N_8082,N_6672);
nand U11366 (N_11366,N_9191,N_6322);
nor U11367 (N_11367,N_8851,N_5717);
nor U11368 (N_11368,N_8137,N_9419);
nor U11369 (N_11369,N_5917,N_5800);
xnor U11370 (N_11370,N_8988,N_9906);
and U11371 (N_11371,N_5027,N_6764);
nor U11372 (N_11372,N_7737,N_6910);
nand U11373 (N_11373,N_5330,N_9441);
nand U11374 (N_11374,N_8611,N_6968);
or U11375 (N_11375,N_6772,N_8294);
or U11376 (N_11376,N_7483,N_6137);
nor U11377 (N_11377,N_8438,N_8126);
xor U11378 (N_11378,N_9851,N_8850);
nor U11379 (N_11379,N_7543,N_8737);
nor U11380 (N_11380,N_8819,N_8956);
nand U11381 (N_11381,N_6753,N_9493);
xnor U11382 (N_11382,N_5245,N_6950);
nor U11383 (N_11383,N_7785,N_6356);
or U11384 (N_11384,N_7682,N_8868);
and U11385 (N_11385,N_9937,N_8970);
nand U11386 (N_11386,N_7122,N_5347);
nand U11387 (N_11387,N_6854,N_8449);
nand U11388 (N_11388,N_7409,N_5033);
and U11389 (N_11389,N_6716,N_5154);
or U11390 (N_11390,N_7557,N_9845);
nor U11391 (N_11391,N_5874,N_9925);
and U11392 (N_11392,N_8341,N_5505);
or U11393 (N_11393,N_5395,N_9001);
and U11394 (N_11394,N_7729,N_9281);
or U11395 (N_11395,N_9970,N_8183);
nand U11396 (N_11396,N_6370,N_9578);
and U11397 (N_11397,N_6836,N_8668);
nand U11398 (N_11398,N_7585,N_9284);
nand U11399 (N_11399,N_6291,N_7107);
and U11400 (N_11400,N_8702,N_8843);
nand U11401 (N_11401,N_5920,N_5363);
xnor U11402 (N_11402,N_6667,N_5834);
nor U11403 (N_11403,N_5465,N_8792);
or U11404 (N_11404,N_5344,N_5925);
nor U11405 (N_11405,N_9872,N_8361);
nand U11406 (N_11406,N_9457,N_9263);
nand U11407 (N_11407,N_8576,N_6056);
nand U11408 (N_11408,N_6413,N_8805);
nor U11409 (N_11409,N_8675,N_5058);
and U11410 (N_11410,N_9814,N_5835);
xnor U11411 (N_11411,N_7065,N_7740);
nand U11412 (N_11412,N_5460,N_9282);
xor U11413 (N_11413,N_6797,N_5383);
or U11414 (N_11414,N_5962,N_9497);
and U11415 (N_11415,N_9152,N_5073);
and U11416 (N_11416,N_8691,N_7436);
or U11417 (N_11417,N_5819,N_6824);
nand U11418 (N_11418,N_8671,N_8765);
nor U11419 (N_11419,N_6237,N_9482);
or U11420 (N_11420,N_7652,N_5192);
nor U11421 (N_11421,N_7178,N_6345);
nand U11422 (N_11422,N_5663,N_9522);
and U11423 (N_11423,N_7198,N_8485);
and U11424 (N_11424,N_7017,N_8174);
nand U11425 (N_11425,N_9546,N_8446);
nor U11426 (N_11426,N_6317,N_8616);
or U11427 (N_11427,N_6512,N_8836);
nor U11428 (N_11428,N_6210,N_7136);
nand U11429 (N_11429,N_5030,N_6788);
nand U11430 (N_11430,N_6813,N_9029);
and U11431 (N_11431,N_6149,N_5585);
nand U11432 (N_11432,N_6051,N_5811);
or U11433 (N_11433,N_5119,N_5433);
nor U11434 (N_11434,N_5276,N_9005);
xnor U11435 (N_11435,N_7636,N_5264);
nand U11436 (N_11436,N_7735,N_9993);
nand U11437 (N_11437,N_5142,N_8291);
or U11438 (N_11438,N_8648,N_9990);
and U11439 (N_11439,N_7705,N_6670);
nand U11440 (N_11440,N_7375,N_6298);
nand U11441 (N_11441,N_8519,N_6453);
and U11442 (N_11442,N_7750,N_8895);
or U11443 (N_11443,N_8276,N_9175);
xnor U11444 (N_11444,N_5227,N_5613);
and U11445 (N_11445,N_5415,N_8408);
or U11446 (N_11446,N_9933,N_9816);
and U11447 (N_11447,N_6469,N_7388);
and U11448 (N_11448,N_9938,N_8768);
and U11449 (N_11449,N_9448,N_6017);
nor U11450 (N_11450,N_5525,N_9306);
and U11451 (N_11451,N_7111,N_9764);
nor U11452 (N_11452,N_7947,N_5626);
or U11453 (N_11453,N_6343,N_6369);
nand U11454 (N_11454,N_9277,N_9023);
nand U11455 (N_11455,N_9701,N_7399);
or U11456 (N_11456,N_5348,N_6157);
and U11457 (N_11457,N_8208,N_5682);
nor U11458 (N_11458,N_9638,N_5225);
and U11459 (N_11459,N_6741,N_9028);
nor U11460 (N_11460,N_5257,N_5702);
nand U11461 (N_11461,N_6635,N_6067);
nor U11462 (N_11462,N_8699,N_5981);
and U11463 (N_11463,N_8394,N_7151);
xnor U11464 (N_11464,N_6885,N_7418);
xor U11465 (N_11465,N_8628,N_8784);
xnor U11466 (N_11466,N_5820,N_9478);
nand U11467 (N_11467,N_9314,N_8592);
xnor U11468 (N_11468,N_8547,N_7754);
nand U11469 (N_11469,N_7241,N_8473);
and U11470 (N_11470,N_7513,N_5345);
nand U11471 (N_11471,N_9387,N_8567);
and U11472 (N_11472,N_7847,N_8992);
or U11473 (N_11473,N_9968,N_5726);
or U11474 (N_11474,N_7577,N_5195);
xor U11475 (N_11475,N_6275,N_5052);
nand U11476 (N_11476,N_5576,N_8251);
nand U11477 (N_11477,N_7000,N_7510);
xnor U11478 (N_11478,N_9400,N_8893);
xor U11479 (N_11479,N_9898,N_7981);
nor U11480 (N_11480,N_5884,N_5419);
xnor U11481 (N_11481,N_9229,N_5652);
or U11482 (N_11482,N_7276,N_5364);
nand U11483 (N_11483,N_9639,N_9818);
and U11484 (N_11484,N_5349,N_8806);
nand U11485 (N_11485,N_5098,N_7985);
nand U11486 (N_11486,N_6197,N_5434);
xnor U11487 (N_11487,N_6972,N_7133);
nor U11488 (N_11488,N_8626,N_5050);
or U11489 (N_11489,N_7738,N_6205);
or U11490 (N_11490,N_8409,N_8543);
and U11491 (N_11491,N_8808,N_5858);
and U11492 (N_11492,N_8510,N_8656);
nand U11493 (N_11493,N_6610,N_5016);
nor U11494 (N_11494,N_9130,N_8727);
nand U11495 (N_11495,N_7262,N_7342);
and U11496 (N_11496,N_7245,N_7341);
or U11497 (N_11497,N_8958,N_6700);
or U11498 (N_11498,N_5399,N_7924);
or U11499 (N_11499,N_8807,N_6233);
nand U11500 (N_11500,N_8367,N_8557);
or U11501 (N_11501,N_8721,N_6160);
nor U11502 (N_11502,N_5821,N_6751);
and U11503 (N_11503,N_6282,N_7648);
and U11504 (N_11504,N_9504,N_9946);
or U11505 (N_11505,N_6872,N_5336);
nor U11506 (N_11506,N_9907,N_9041);
nand U11507 (N_11507,N_9671,N_5499);
nor U11508 (N_11508,N_9254,N_6004);
xor U11509 (N_11509,N_9072,N_5323);
or U11510 (N_11510,N_8193,N_8177);
xnor U11511 (N_11511,N_9580,N_8078);
and U11512 (N_11512,N_9878,N_9926);
and U11513 (N_11513,N_8157,N_6043);
nand U11514 (N_11514,N_6641,N_5283);
xor U11515 (N_11515,N_6020,N_8712);
or U11516 (N_11516,N_7387,N_8315);
xnor U11517 (N_11517,N_7715,N_6035);
or U11518 (N_11518,N_6526,N_5102);
nor U11519 (N_11519,N_5604,N_6118);
nor U11520 (N_11520,N_7977,N_5358);
nand U11521 (N_11521,N_6299,N_6861);
or U11522 (N_11522,N_6325,N_7883);
and U11523 (N_11523,N_5062,N_6901);
and U11524 (N_11524,N_6449,N_6983);
or U11525 (N_11525,N_7898,N_9194);
or U11526 (N_11526,N_8253,N_6814);
and U11527 (N_11527,N_7846,N_6069);
nand U11528 (N_11528,N_9544,N_7553);
and U11529 (N_11529,N_7128,N_8625);
nor U11530 (N_11530,N_6216,N_9711);
or U11531 (N_11531,N_7033,N_7594);
and U11532 (N_11532,N_5855,N_5002);
nor U11533 (N_11533,N_6346,N_9978);
and U11534 (N_11534,N_6774,N_7673);
nand U11535 (N_11535,N_5816,N_6673);
nand U11536 (N_11536,N_7172,N_9548);
nand U11537 (N_11537,N_9027,N_6181);
nor U11538 (N_11538,N_7486,N_9505);
xnor U11539 (N_11539,N_5606,N_6584);
or U11540 (N_11540,N_7913,N_7779);
and U11541 (N_11541,N_8040,N_7330);
nand U11542 (N_11542,N_7560,N_8986);
and U11543 (N_11543,N_7191,N_8501);
nand U11544 (N_11544,N_5384,N_7118);
or U11545 (N_11545,N_9692,N_5208);
nand U11546 (N_11546,N_5067,N_5207);
nor U11547 (N_11547,N_5351,N_5587);
or U11548 (N_11548,N_8141,N_8245);
or U11549 (N_11549,N_8679,N_8098);
or U11550 (N_11550,N_5090,N_6754);
or U11551 (N_11551,N_8614,N_6817);
and U11552 (N_11552,N_7670,N_5574);
nand U11553 (N_11553,N_6267,N_8533);
nor U11554 (N_11554,N_8581,N_7792);
nor U11555 (N_11555,N_6326,N_5639);
and U11556 (N_11556,N_7401,N_6991);
nand U11557 (N_11557,N_8274,N_6415);
or U11558 (N_11558,N_7165,N_7835);
nand U11559 (N_11559,N_9507,N_8145);
and U11560 (N_11560,N_7443,N_9988);
or U11561 (N_11561,N_6795,N_7992);
or U11562 (N_11562,N_5611,N_9085);
nor U11563 (N_11563,N_5738,N_7044);
and U11564 (N_11564,N_8476,N_6268);
or U11565 (N_11565,N_5100,N_7288);
nand U11566 (N_11566,N_6893,N_6524);
and U11567 (N_11567,N_7716,N_8709);
nor U11568 (N_11568,N_5241,N_5600);
and U11569 (N_11569,N_9336,N_9219);
nor U11570 (N_11570,N_9320,N_8565);
and U11571 (N_11571,N_5232,N_7323);
and U11572 (N_11572,N_7251,N_9312);
xor U11573 (N_11573,N_7663,N_6806);
nor U11574 (N_11574,N_9037,N_5749);
nor U11575 (N_11575,N_9366,N_7366);
nor U11576 (N_11576,N_6590,N_9574);
or U11577 (N_11577,N_8812,N_8124);
and U11578 (N_11578,N_5972,N_7526);
nand U11579 (N_11579,N_9422,N_8904);
and U11580 (N_11580,N_7026,N_5551);
nand U11581 (N_11581,N_9608,N_9236);
xnor U11582 (N_11582,N_7522,N_7058);
and U11583 (N_11583,N_5031,N_8889);
xnor U11584 (N_11584,N_8728,N_5164);
or U11585 (N_11585,N_5205,N_6416);
or U11586 (N_11586,N_5631,N_6316);
or U11587 (N_11587,N_9528,N_7269);
or U11588 (N_11588,N_6382,N_8135);
nor U11589 (N_11589,N_5554,N_7168);
and U11590 (N_11590,N_9231,N_6500);
nor U11591 (N_11591,N_7134,N_8655);
and U11592 (N_11592,N_5413,N_9635);
and U11593 (N_11593,N_7495,N_9455);
xor U11594 (N_11594,N_5634,N_7860);
xnor U11595 (N_11595,N_6001,N_8536);
and U11596 (N_11596,N_9584,N_9745);
and U11597 (N_11597,N_7159,N_9444);
nand U11598 (N_11598,N_5101,N_6856);
and U11599 (N_11599,N_6350,N_5392);
nand U11600 (N_11600,N_7432,N_8271);
xnor U11601 (N_11601,N_7762,N_6665);
or U11602 (N_11602,N_9117,N_6702);
or U11603 (N_11603,N_6245,N_8496);
nand U11604 (N_11604,N_6410,N_6419);
nor U11605 (N_11605,N_8552,N_6269);
nor U11606 (N_11606,N_7613,N_7013);
or U11607 (N_11607,N_9894,N_6270);
nand U11608 (N_11608,N_7838,N_8651);
and U11609 (N_11609,N_7934,N_5678);
nand U11610 (N_11610,N_5957,N_5481);
and U11611 (N_11611,N_8351,N_7790);
or U11612 (N_11612,N_9660,N_8275);
nor U11613 (N_11613,N_5039,N_7624);
or U11614 (N_11614,N_8005,N_7067);
and U11615 (N_11615,N_7331,N_5179);
xnor U11616 (N_11616,N_8883,N_7012);
or U11617 (N_11617,N_7272,N_6176);
nand U11618 (N_11618,N_9216,N_6311);
nor U11619 (N_11619,N_7849,N_6263);
or U11620 (N_11620,N_6534,N_8521);
and U11621 (N_11621,N_7870,N_6373);
xnor U11622 (N_11622,N_6328,N_5768);
nor U11623 (N_11623,N_8740,N_8987);
xnor U11624 (N_11624,N_6080,N_8159);
and U11625 (N_11625,N_8991,N_8719);
xor U11626 (N_11626,N_6391,N_5719);
and U11627 (N_11627,N_6378,N_5650);
or U11628 (N_11628,N_8798,N_6847);
nand U11629 (N_11629,N_5867,N_7828);
nand U11630 (N_11630,N_8422,N_9294);
nor U11631 (N_11631,N_8632,N_5936);
nor U11632 (N_11632,N_9490,N_7825);
nand U11633 (N_11633,N_9545,N_5442);
and U11634 (N_11634,N_8891,N_9405);
xnor U11635 (N_11635,N_9831,N_7002);
nand U11636 (N_11636,N_8357,N_5210);
and U11637 (N_11637,N_8376,N_5273);
nor U11638 (N_11638,N_7931,N_7037);
or U11639 (N_11639,N_9333,N_7575);
or U11640 (N_11640,N_9239,N_9682);
xnor U11641 (N_11641,N_8464,N_5492);
nor U11642 (N_11642,N_7967,N_9979);
nor U11643 (N_11643,N_6633,N_6495);
nand U11644 (N_11644,N_5840,N_9603);
nor U11645 (N_11645,N_9694,N_6450);
nand U11646 (N_11646,N_9326,N_5080);
xnor U11647 (N_11647,N_6970,N_8537);
or U11648 (N_11648,N_6437,N_5534);
or U11649 (N_11649,N_7496,N_7784);
nand U11650 (N_11650,N_8870,N_8498);
or U11651 (N_11651,N_7358,N_9156);
nor U11652 (N_11652,N_9120,N_5592);
nor U11653 (N_11653,N_7910,N_9791);
or U11654 (N_11654,N_5203,N_6077);
nand U11655 (N_11655,N_8620,N_5877);
or U11656 (N_11656,N_9893,N_9071);
nand U11657 (N_11657,N_8128,N_8772);
nand U11658 (N_11658,N_7441,N_6398);
nand U11659 (N_11659,N_5137,N_7239);
and U11660 (N_11660,N_9982,N_6912);
nor U11661 (N_11661,N_6629,N_7146);
xor U11662 (N_11662,N_8825,N_9841);
nand U11663 (N_11663,N_6260,N_7821);
nand U11664 (N_11664,N_8673,N_8107);
nand U11665 (N_11665,N_7886,N_6919);
xnor U11666 (N_11666,N_9828,N_6715);
xor U11667 (N_11667,N_8503,N_5934);
nor U11668 (N_11668,N_9583,N_7373);
nor U11669 (N_11669,N_9486,N_5748);
and U11670 (N_11670,N_7983,N_6583);
nor U11671 (N_11671,N_9837,N_9965);
nor U11672 (N_11672,N_7045,N_9810);
or U11673 (N_11673,N_8697,N_8375);
or U11674 (N_11674,N_5382,N_9234);
xor U11675 (N_11675,N_9503,N_6300);
or U11676 (N_11676,N_6301,N_9292);
xnor U11677 (N_11677,N_7138,N_6952);
or U11678 (N_11678,N_8238,N_8876);
xor U11679 (N_11679,N_9304,N_8690);
nand U11680 (N_11680,N_7340,N_9857);
nand U11681 (N_11681,N_6158,N_6868);
nand U11682 (N_11682,N_8325,N_6079);
nand U11683 (N_11683,N_7848,N_9566);
xnor U11684 (N_11684,N_9759,N_8064);
nand U11685 (N_11685,N_9439,N_6657);
nand U11686 (N_11686,N_8677,N_6602);
or U11687 (N_11687,N_8995,N_5944);
nor U11688 (N_11688,N_7452,N_9139);
nor U11689 (N_11689,N_7658,N_9573);
nand U11690 (N_11690,N_7713,N_9960);
or U11691 (N_11691,N_9648,N_5893);
and U11692 (N_11692,N_9492,N_5438);
xnor U11693 (N_11693,N_9290,N_5641);
and U11694 (N_11694,N_6756,N_6221);
nor U11695 (N_11695,N_7521,N_6990);
or U11696 (N_11696,N_6008,N_9313);
or U11697 (N_11697,N_9083,N_6123);
nand U11698 (N_11698,N_7662,N_9766);
nor U11699 (N_11699,N_9670,N_6042);
xor U11700 (N_11700,N_9735,N_5740);
and U11701 (N_11701,N_8553,N_8639);
and U11702 (N_11702,N_5825,N_8636);
nor U11703 (N_11703,N_8752,N_5457);
or U11704 (N_11704,N_5507,N_9879);
nand U11705 (N_11705,N_5615,N_7050);
nor U11706 (N_11706,N_6505,N_8733);
and U11707 (N_11707,N_9765,N_9058);
and U11708 (N_11708,N_6902,N_9860);
and U11709 (N_11709,N_5568,N_9746);
or U11710 (N_11710,N_8754,N_9706);
xor U11711 (N_11711,N_8695,N_6896);
and U11712 (N_11712,N_8979,N_8799);
nand U11713 (N_11713,N_7041,N_9749);
and U11714 (N_11714,N_7689,N_9685);
and U11715 (N_11715,N_8723,N_5659);
and U11716 (N_11716,N_8133,N_9346);
xor U11717 (N_11717,N_9476,N_7725);
nor U11718 (N_11718,N_9007,N_9501);
and U11719 (N_11719,N_7548,N_8304);
nor U11720 (N_11720,N_7685,N_6874);
nor U11721 (N_11721,N_6134,N_9750);
or U11722 (N_11722,N_6649,N_9267);
nand U11723 (N_11723,N_5674,N_6869);
and U11724 (N_11724,N_9909,N_8957);
and U11725 (N_11725,N_6121,N_7359);
xor U11726 (N_11726,N_6878,N_9551);
and U11727 (N_11727,N_8666,N_6671);
nand U11728 (N_11728,N_7395,N_7445);
and U11729 (N_11729,N_7392,N_7664);
nand U11730 (N_11730,N_8261,N_7556);
nor U11731 (N_11731,N_5378,N_6058);
nand U11732 (N_11732,N_6898,N_7984);
and U11733 (N_11733,N_9394,N_6577);
nor U11734 (N_11734,N_8026,N_6459);
nor U11735 (N_11735,N_6340,N_8584);
and U11736 (N_11736,N_7064,N_7368);
nor U11737 (N_11737,N_9725,N_5938);
and U11738 (N_11738,N_8516,N_8386);
nand U11739 (N_11739,N_6596,N_7029);
and U11740 (N_11740,N_5876,N_8678);
and U11741 (N_11741,N_9362,N_6360);
nand U11742 (N_11742,N_6674,N_5252);
nand U11743 (N_11743,N_6178,N_8269);
nand U11744 (N_11744,N_5401,N_7206);
or U11745 (N_11745,N_8813,N_8926);
or U11746 (N_11746,N_7555,N_8676);
xnor U11747 (N_11747,N_9227,N_5117);
xnor U11748 (N_11748,N_5896,N_6492);
nand U11749 (N_11749,N_9379,N_7578);
or U11750 (N_11750,N_5151,N_5806);
or U11751 (N_11751,N_7062,N_8667);
xnor U11752 (N_11752,N_6503,N_6446);
xnor U11753 (N_11753,N_6010,N_9855);
or U11754 (N_11754,N_8574,N_6063);
or U11755 (N_11755,N_6625,N_9491);
xnor U11756 (N_11756,N_6116,N_8013);
xnor U11757 (N_11757,N_7185,N_6782);
nand U11758 (N_11758,N_9593,N_8539);
xor U11759 (N_11759,N_6695,N_8001);
xor U11760 (N_11760,N_7155,N_7742);
or U11761 (N_11761,N_6075,N_5966);
or U11762 (N_11762,N_5570,N_7666);
nor U11763 (N_11763,N_9527,N_9955);
nand U11764 (N_11764,N_9094,N_8390);
nand U11765 (N_11765,N_5736,N_5910);
nand U11766 (N_11766,N_5381,N_6147);
xor U11767 (N_11767,N_7672,N_9811);
nand U11768 (N_11768,N_6018,N_6844);
or U11769 (N_11769,N_7649,N_7632);
and U11770 (N_11770,N_7592,N_8319);
nand U11771 (N_11771,N_9919,N_6877);
or U11772 (N_11772,N_5919,N_9821);
nor U11773 (N_11773,N_5219,N_7587);
nand U11774 (N_11774,N_8652,N_8176);
nor U11775 (N_11775,N_9090,N_7502);
nor U11776 (N_11776,N_7745,N_7880);
nand U11777 (N_11777,N_7113,N_9275);
or U11778 (N_11778,N_5369,N_7558);
nor U11779 (N_11779,N_5580,N_6899);
nand U11780 (N_11780,N_7498,N_9929);
nand U11781 (N_11781,N_7454,N_6936);
and U11782 (N_11782,N_6606,N_6721);
nor U11783 (N_11783,N_6821,N_5526);
nor U11784 (N_11784,N_9480,N_6388);
nand U11785 (N_11785,N_6690,N_7054);
or U11786 (N_11786,N_5761,N_9370);
nand U11787 (N_11787,N_7413,N_6375);
or U11788 (N_11788,N_6331,N_5975);
or U11789 (N_11789,N_5194,N_7180);
or U11790 (N_11790,N_6528,N_9211);
nand U11791 (N_11791,N_6119,N_5282);
or U11792 (N_11792,N_9784,N_9187);
and U11793 (N_11793,N_9391,N_9920);
nor U11794 (N_11794,N_9612,N_7428);
or U11795 (N_11795,N_7386,N_5902);
and U11796 (N_11796,N_5947,N_5708);
and U11797 (N_11797,N_9264,N_8908);
nor U11798 (N_11798,N_6589,N_5842);
nand U11799 (N_11799,N_5093,N_9081);
and U11800 (N_11800,N_8513,N_6791);
and U11801 (N_11801,N_9147,N_8049);
and U11802 (N_11802,N_8816,N_7192);
and U11803 (N_11803,N_9767,N_6122);
nor U11804 (N_11804,N_7177,N_8878);
nor U11805 (N_11805,N_5709,N_5420);
xor U11806 (N_11806,N_7512,N_7731);
and U11807 (N_11807,N_5508,N_9589);
or U11808 (N_11808,N_9247,N_9757);
nor U11809 (N_11809,N_7878,N_5903);
and U11810 (N_11810,N_7879,N_7237);
and U11811 (N_11811,N_7142,N_5354);
nand U11812 (N_11812,N_9730,N_5353);
and U11813 (N_11813,N_5072,N_8950);
xnor U11814 (N_11814,N_7089,N_9932);
nand U11815 (N_11815,N_7751,N_7055);
nand U11816 (N_11816,N_9367,N_8068);
nand U11817 (N_11817,N_8821,N_8980);
or U11818 (N_11818,N_9149,N_5406);
xnor U11819 (N_11819,N_6963,N_7507);
and U11820 (N_11820,N_9309,N_9834);
nand U11821 (N_11821,N_6131,N_8542);
nor U11822 (N_11822,N_7661,N_9091);
nand U11823 (N_11823,N_7126,N_7232);
and U11824 (N_11824,N_7680,N_5503);
nor U11825 (N_11825,N_9080,N_5466);
or U11826 (N_11826,N_6127,N_8538);
or U11827 (N_11827,N_6647,N_5646);
and U11828 (N_11828,N_6620,N_6354);
and U11829 (N_11829,N_6941,N_7916);
nor U11830 (N_11830,N_8571,N_9428);
nand U11831 (N_11831,N_5337,N_9732);
and U11832 (N_11832,N_5797,N_7959);
or U11833 (N_11833,N_6866,N_9280);
nor U11834 (N_11834,N_7676,N_7419);
or U11835 (N_11835,N_9087,N_7137);
xnor U11836 (N_11836,N_9214,N_5089);
xor U11837 (N_11837,N_7533,N_8282);
or U11838 (N_11838,N_6850,N_9742);
or U11839 (N_11839,N_6377,N_6019);
or U11840 (N_11840,N_7193,N_5733);
xnor U11841 (N_11841,N_8546,N_7946);
and U11842 (N_11842,N_7444,N_5662);
and U11843 (N_11843,N_9269,N_6053);
nand U11844 (N_11844,N_9450,N_8949);
or U11845 (N_11845,N_6383,N_8100);
xor U11846 (N_11846,N_7703,N_9168);
nand U11847 (N_11847,N_5984,N_5408);
or U11848 (N_11848,N_7231,N_8590);
nor U11849 (N_11849,N_5624,N_9295);
or U11850 (N_11850,N_9179,N_8556);
and U11851 (N_11851,N_5673,N_7687);
and U11852 (N_11852,N_9241,N_6227);
or U11853 (N_11853,N_5259,N_6349);
nor U11854 (N_11854,N_9652,N_7643);
nand U11855 (N_11855,N_6773,N_9927);
nor U11856 (N_11856,N_9957,N_6190);
xnor U11857 (N_11857,N_6628,N_7550);
nor U11858 (N_11858,N_9188,N_6486);
nand U11859 (N_11859,N_6830,N_7903);
and U11860 (N_11860,N_7788,N_6107);
nor U11861 (N_11861,N_8350,N_9931);
nand U11862 (N_11862,N_8525,N_7824);
or U11863 (N_11863,N_6293,N_9359);
or U11864 (N_11864,N_8201,N_7844);
or U11865 (N_11865,N_7586,N_6581);
or U11866 (N_11866,N_5079,N_6842);
xor U11867 (N_11867,N_8909,N_6297);
nand U11868 (N_11868,N_7884,N_9632);
or U11869 (N_11869,N_9977,N_7284);
nor U11870 (N_11870,N_8857,N_5985);
or U11871 (N_11871,N_7711,N_5868);
nand U11872 (N_11872,N_7305,N_9181);
and U11873 (N_11873,N_8156,N_5423);
or U11874 (N_11874,N_8641,N_7242);
or U11875 (N_11875,N_6327,N_6614);
nor U11876 (N_11876,N_9619,N_5827);
and U11877 (N_11877,N_5746,N_9890);
and U11878 (N_11878,N_6170,N_7311);
nor U11879 (N_11879,N_5417,N_6634);
or U11880 (N_11880,N_5711,N_5571);
nand U11881 (N_11881,N_8144,N_7544);
or U11882 (N_11882,N_6292,N_6120);
nand U11883 (N_11883,N_7156,N_5260);
nand U11884 (N_11884,N_9991,N_5130);
nand U11885 (N_11885,N_6151,N_6949);
or U11886 (N_11886,N_7188,N_8890);
or U11887 (N_11887,N_7053,N_5169);
and U11888 (N_11888,N_6072,N_7869);
and U11889 (N_11889,N_6439,N_7063);
or U11890 (N_11890,N_5862,N_7108);
nand U11891 (N_11891,N_8662,N_8358);
nor U11892 (N_11892,N_7460,N_9679);
nor U11893 (N_11893,N_9743,N_9644);
nand U11894 (N_11894,N_8205,N_9824);
nand U11895 (N_11895,N_6142,N_9865);
or U11896 (N_11896,N_9668,N_7691);
or U11897 (N_11897,N_5150,N_9003);
nor U11898 (N_11898,N_8420,N_7826);
and U11899 (N_11899,N_9815,N_6189);
nand U11900 (N_11900,N_8978,N_7853);
nand U11901 (N_11901,N_5424,N_6026);
and U11902 (N_11902,N_5403,N_6113);
or U11903 (N_11903,N_7077,N_8670);
and U11904 (N_11904,N_9397,N_6961);
xor U11905 (N_11905,N_8580,N_9936);
or U11906 (N_11906,N_6279,N_7761);
nor U11907 (N_11907,N_8985,N_6862);
nand U11908 (N_11908,N_9040,N_5298);
nor U11909 (N_11909,N_9702,N_8154);
nor U11910 (N_11910,N_5752,N_8814);
or U11911 (N_11911,N_9466,N_5558);
xnor U11912 (N_11912,N_9069,N_8352);
and U11913 (N_11913,N_7174,N_8211);
nand U11914 (N_11914,N_8301,N_5815);
xor U11915 (N_11915,N_9724,N_6599);
and U11916 (N_11916,N_8687,N_9599);
nand U11917 (N_11917,N_9096,N_9669);
nor U11918 (N_11918,N_5704,N_5980);
nand U11919 (N_11919,N_5301,N_5254);
and U11920 (N_11920,N_6855,N_9463);
nand U11921 (N_11921,N_9161,N_8939);
nand U11922 (N_11922,N_6348,N_7197);
nor U11923 (N_11923,N_8403,N_6499);
xnor U11924 (N_11924,N_6621,N_6804);
or U11925 (N_11925,N_5529,N_8575);
nor U11926 (N_11926,N_8478,N_7596);
or U11927 (N_11927,N_9339,N_5014);
and U11928 (N_11928,N_5539,N_7978);
or U11929 (N_11929,N_6460,N_5022);
nand U11930 (N_11930,N_9025,N_8472);
and U11931 (N_11931,N_8112,N_6169);
nand U11932 (N_11932,N_6545,N_8021);
nor U11933 (N_11933,N_7582,N_8303);
and U11934 (N_11934,N_5665,N_8847);
nand U11935 (N_11935,N_8127,N_7038);
nor U11936 (N_11936,N_8047,N_7131);
or U11937 (N_11937,N_9871,N_7357);
or U11938 (N_11938,N_8075,N_7998);
and U11939 (N_11939,N_7760,N_9795);
xor U11940 (N_11940,N_5064,N_7270);
or U11941 (N_11941,N_6187,N_6272);
nor U11942 (N_11942,N_7561,N_5341);
nand U11943 (N_11943,N_9995,N_5623);
nor U11944 (N_11944,N_6096,N_5705);
and U11945 (N_11945,N_7304,N_6507);
nand U11946 (N_11946,N_5006,N_5414);
nand U11947 (N_11947,N_9392,N_8964);
nor U11948 (N_11948,N_9716,N_7291);
xnor U11949 (N_11949,N_9393,N_6088);
nor U11950 (N_11950,N_8877,N_8582);
nand U11951 (N_11951,N_6769,N_5618);
or U11952 (N_11952,N_8777,N_6218);
and U11953 (N_11953,N_9798,N_8861);
nand U11954 (N_11954,N_6089,N_8791);
or U11955 (N_11955,N_8153,N_5385);
xor U11956 (N_11956,N_5895,N_8045);
and U11957 (N_11957,N_9076,N_6105);
nand U11958 (N_11958,N_7897,N_5829);
xnor U11959 (N_11959,N_5396,N_8811);
xor U11960 (N_11960,N_8642,N_6608);
and U11961 (N_11961,N_6703,N_9358);
and U11962 (N_11962,N_7143,N_6448);
or U11963 (N_11963,N_5861,N_6126);
nor U11964 (N_11964,N_9621,N_5155);
or U11965 (N_11965,N_6803,N_6930);
nand U11966 (N_11966,N_5555,N_6294);
xor U11967 (N_11967,N_6618,N_9678);
and U11968 (N_11968,N_8489,N_6433);
nand U11969 (N_11969,N_8914,N_6890);
nand U11970 (N_11970,N_6379,N_6867);
and U11971 (N_11971,N_9454,N_9266);
or U11972 (N_11972,N_6915,N_6456);
and U11973 (N_11973,N_6264,N_9097);
nand U11974 (N_11974,N_9550,N_8952);
nor U11975 (N_11975,N_9896,N_8373);
nor U11976 (N_11976,N_6677,N_5627);
nor U11977 (N_11977,N_7933,N_6440);
xnor U11978 (N_11978,N_7072,N_7052);
nor U11979 (N_11979,N_6394,N_5494);
xnor U11980 (N_11980,N_6365,N_5084);
nand U11981 (N_11981,N_6247,N_7456);
and U11982 (N_11982,N_7795,N_5011);
or U11983 (N_11983,N_7350,N_9673);
nor U11984 (N_11984,N_7345,N_7976);
and U11985 (N_11985,N_6811,N_7642);
and U11986 (N_11986,N_5888,N_7039);
nand U11987 (N_11987,N_8249,N_8429);
nor U11988 (N_11988,N_8646,N_5026);
nand U11989 (N_11989,N_6651,N_5019);
nor U11990 (N_11990,N_9510,N_7328);
nand U11991 (N_11991,N_7845,N_8410);
xnor U11992 (N_11992,N_8337,N_5997);
xnor U11993 (N_11993,N_8356,N_6407);
and U11994 (N_11994,N_8818,N_6234);
nor U11995 (N_11995,N_8346,N_7671);
nor U11996 (N_11996,N_8035,N_9535);
nand U11997 (N_11997,N_6946,N_9695);
or U11998 (N_11998,N_6213,N_7719);
nor U11999 (N_11999,N_7960,N_8451);
nor U12000 (N_12000,N_5422,N_5387);
nor U12001 (N_12001,N_5693,N_9321);
nor U12002 (N_12002,N_5923,N_9876);
and U12003 (N_12003,N_6953,N_7589);
nor U12004 (N_12004,N_5961,N_7518);
and U12005 (N_12005,N_7855,N_8743);
nor U12006 (N_12006,N_9435,N_8391);
and U12007 (N_12007,N_9999,N_6191);
nor U12008 (N_12008,N_7109,N_7896);
or U12009 (N_12009,N_6185,N_9207);
nand U12010 (N_12010,N_7349,N_9861);
nor U12011 (N_12011,N_6539,N_6212);
nand U12012 (N_12012,N_9604,N_8046);
and U12013 (N_12013,N_5103,N_5238);
nand U12014 (N_12014,N_6104,N_7674);
nand U12015 (N_12015,N_5670,N_7799);
xnor U12016 (N_12016,N_5782,N_9910);
or U12017 (N_12017,N_9738,N_7407);
nor U12018 (N_12018,N_5765,N_9530);
and U12019 (N_12019,N_7768,N_5956);
or U12020 (N_12020,N_9233,N_6917);
and U12021 (N_12021,N_9456,N_9024);
or U12022 (N_12022,N_7011,N_5612);
or U12023 (N_12023,N_8434,N_7081);
nand U12024 (N_12024,N_5274,N_7654);
or U12025 (N_12025,N_9699,N_7817);
and U12026 (N_12026,N_7935,N_5109);
or U12027 (N_12027,N_7036,N_9555);
and U12028 (N_12028,N_7173,N_9812);
nor U12029 (N_12029,N_6997,N_8822);
nor U12030 (N_12030,N_7354,N_9248);
xnor U12031 (N_12031,N_8136,N_8759);
or U12032 (N_12032,N_7299,N_7863);
and U12033 (N_12033,N_7293,N_8202);
nor U12034 (N_12034,N_7618,N_8564);
nand U12035 (N_12035,N_5032,N_8624);
nand U12036 (N_12036,N_5959,N_9262);
and U12037 (N_12037,N_5340,N_7329);
and U12038 (N_12038,N_8555,N_7263);
nand U12039 (N_12039,N_7515,N_9704);
nor U12040 (N_12040,N_9160,N_6155);
nor U12041 (N_12041,N_5123,N_9934);
or U12042 (N_12042,N_8089,N_5849);
and U12043 (N_12043,N_7545,N_7970);
nand U12044 (N_12044,N_9801,N_5325);
nor U12045 (N_12045,N_9016,N_8698);
and U12046 (N_12046,N_9451,N_6582);
or U12047 (N_12047,N_5216,N_9220);
and U12048 (N_12048,N_9843,N_7701);
xor U12049 (N_12049,N_8973,N_7746);
xnor U12050 (N_12050,N_6533,N_8644);
or U12051 (N_12051,N_9283,N_7416);
xnor U12052 (N_12052,N_6699,N_9296);
xor U12053 (N_12053,N_5380,N_5807);
nor U12054 (N_12054,N_9052,N_8362);
nand U12055 (N_12055,N_9151,N_5250);
nor U12056 (N_12056,N_7800,N_7132);
or U12057 (N_12057,N_7546,N_9423);
nor U12058 (N_12058,N_7352,N_6253);
and U12059 (N_12059,N_9223,N_8929);
or U12060 (N_12060,N_9409,N_6815);
or U12061 (N_12061,N_9273,N_5163);
nor U12062 (N_12062,N_5366,N_8900);
xnor U12063 (N_12063,N_7422,N_7097);
xnor U12064 (N_12064,N_9417,N_9854);
nor U12065 (N_12065,N_9790,N_7130);
nand U12066 (N_12066,N_6386,N_6414);
xnor U12067 (N_12067,N_6086,N_5231);
and U12068 (N_12068,N_5864,N_7938);
or U12069 (N_12069,N_9474,N_9762);
and U12070 (N_12070,N_8795,N_7698);
nand U12071 (N_12071,N_6368,N_6220);
nor U12072 (N_12072,N_7807,N_7096);
or U12073 (N_12073,N_7028,N_8404);
nor U12074 (N_12074,N_8659,N_6357);
or U12075 (N_12075,N_5502,N_6971);
nand U12076 (N_12076,N_6182,N_5755);
or U12077 (N_12077,N_9118,N_6362);
xnor U12078 (N_12078,N_5963,N_5162);
or U12079 (N_12079,N_5533,N_6897);
nand U12080 (N_12080,N_8941,N_5111);
or U12081 (N_12081,N_6223,N_6479);
xnor U12082 (N_12082,N_6964,N_9203);
nor U12083 (N_12083,N_5202,N_5190);
nand U12084 (N_12084,N_9082,N_8151);
nand U12085 (N_12085,N_5007,N_5063);
nor U12086 (N_12086,N_9307,N_5005);
nand U12087 (N_12087,N_5277,N_8071);
nand U12088 (N_12088,N_7566,N_9265);
xor U12089 (N_12089,N_9552,N_9141);
or U12090 (N_12090,N_6888,N_6040);
nor U12091 (N_12091,N_5449,N_9651);
xnor U12092 (N_12092,N_6395,N_8125);
nand U12093 (N_12093,N_5041,N_6295);
and U12094 (N_12094,N_5318,N_9813);
xnor U12095 (N_12095,N_6036,N_8585);
nor U12096 (N_12096,N_5773,N_6766);
and U12097 (N_12097,N_9877,N_9093);
nor U12098 (N_12098,N_6557,N_7573);
nand U12099 (N_12099,N_7547,N_8713);
and U12100 (N_12100,N_9686,N_8330);
or U12101 (N_12101,N_9736,N_6812);
nand U12102 (N_12102,N_8076,N_5591);
and U12103 (N_12103,N_9914,N_8747);
or U12104 (N_12104,N_6865,N_6487);
nand U12105 (N_12105,N_8286,N_8204);
and U12106 (N_12106,N_8092,N_5214);
nor U12107 (N_12107,N_9142,N_7834);
nand U12108 (N_12108,N_6767,N_8411);
nor U12109 (N_12109,N_6025,N_8563);
nand U12110 (N_12110,N_7619,N_8160);
nor U12111 (N_12111,N_9658,N_6882);
or U12112 (N_12112,N_7336,N_9657);
xor U12113 (N_12113,N_5517,N_5597);
and U12114 (N_12114,N_9521,N_6393);
or U12115 (N_12115,N_7877,N_6554);
and U12116 (N_12116,N_8873,N_6937);
or U12117 (N_12117,N_9719,N_6697);
nor U12118 (N_12118,N_9022,N_9256);
nand U12119 (N_12119,N_7006,N_6655);
nand U12120 (N_12120,N_8928,N_7249);
xnor U12121 (N_12121,N_6007,N_8830);
nand U12122 (N_12122,N_5174,N_9206);
xor U12123 (N_12123,N_6442,N_8414);
and U12124 (N_12124,N_5106,N_8658);
or U12125 (N_12125,N_6560,N_7836);
nor U12126 (N_12126,N_7579,N_6661);
or U12127 (N_12127,N_7612,N_5375);
or U12128 (N_12128,N_7025,N_9335);
or U12129 (N_12129,N_7363,N_8588);
or U12130 (N_12130,N_9361,N_5995);
xnor U12131 (N_12131,N_5451,N_5594);
or U12132 (N_12132,N_6038,N_5788);
or U12133 (N_12133,N_5812,N_9888);
and U12134 (N_12134,N_7889,N_6255);
and U12135 (N_12135,N_9627,N_9677);
xnor U12136 (N_12136,N_5924,N_8138);
nor U12137 (N_12137,N_6447,N_6266);
xor U12138 (N_12138,N_7256,N_7987);
nor U12139 (N_12139,N_7088,N_7749);
or U12140 (N_12140,N_7829,N_6135);
xor U12141 (N_12141,N_7184,N_8342);
nand U12142 (N_12142,N_5637,N_6199);
nand U12143 (N_12143,N_9164,N_9948);
or U12144 (N_12144,N_6755,N_7659);
nor U12145 (N_12145,N_5173,N_9647);
nor U12146 (N_12146,N_8038,N_8937);
and U12147 (N_12147,N_9245,N_6592);
or U12148 (N_12148,N_9412,N_7965);
or U12149 (N_12149,N_6163,N_7580);
nand U12150 (N_12150,N_7517,N_8852);
nand U12151 (N_12151,N_5331,N_6497);
nor U12152 (N_12152,N_7140,N_9322);
or U12153 (N_12153,N_9998,N_7798);
xor U12154 (N_12154,N_7294,N_8117);
nand U12155 (N_12155,N_8207,N_9508);
or U12156 (N_12156,N_5776,N_8083);
and U12157 (N_12157,N_6636,N_7355);
nor U12158 (N_12158,N_9329,N_6363);
and U12159 (N_12159,N_6167,N_6095);
or U12160 (N_12160,N_6429,N_8169);
and U12161 (N_12161,N_7034,N_6750);
and U12162 (N_12162,N_6306,N_8839);
and U12163 (N_12163,N_7027,N_6551);
and U12164 (N_12164,N_8606,N_5826);
nor U12165 (N_12165,N_6397,N_7169);
and U12166 (N_12166,N_5784,N_6066);
and U12167 (N_12167,N_7279,N_6921);
nor U12168 (N_12168,N_9368,N_7882);
nand U12169 (N_12169,N_6585,N_7595);
nor U12170 (N_12170,N_5675,N_8660);
xnor U12171 (N_12171,N_8067,N_5118);
xnor U12172 (N_12172,N_9487,N_6924);
or U12173 (N_12173,N_8776,N_6724);
or U12174 (N_12174,N_6627,N_7103);
and U12175 (N_12175,N_6685,N_7087);
or U12176 (N_12176,N_6805,N_6540);
nand U12177 (N_12177,N_7275,N_7499);
or U12178 (N_12178,N_5334,N_9429);
nand U12179 (N_12179,N_6739,N_5271);
and U12180 (N_12180,N_8209,N_6523);
nor U12181 (N_12181,N_9985,N_9973);
nand U12182 (N_12182,N_9549,N_6052);
nor U12183 (N_12183,N_6746,N_9404);
and U12184 (N_12184,N_5240,N_6613);
nor U12185 (N_12185,N_5521,N_9013);
or U12186 (N_12186,N_9958,N_8983);
nor U12187 (N_12187,N_7708,N_5625);
nand U12188 (N_12188,N_7994,N_6706);
xor U12189 (N_12189,N_5595,N_5860);
or U12190 (N_12190,N_7859,N_7187);
xnor U12191 (N_12191,N_9204,N_6494);
nand U12192 (N_12192,N_5359,N_9170);
or U12193 (N_12193,N_5167,N_9622);
nand U12194 (N_12194,N_9722,N_8664);
and U12195 (N_12195,N_7668,N_8140);
or U12196 (N_12196,N_9994,N_5126);
and U12197 (N_12197,N_6145,N_8534);
and U12198 (N_12198,N_7117,N_5280);
and U12199 (N_12199,N_5115,N_7572);
xor U12200 (N_12200,N_6262,N_5268);
and U12201 (N_12201,N_8758,N_6914);
or U12202 (N_12202,N_5775,N_7457);
nor U12203 (N_12203,N_6709,N_7722);
nor U12204 (N_12204,N_9334,N_6055);
xnor U12205 (N_12205,N_9059,N_9867);
or U12206 (N_12206,N_7867,N_9002);
and U12207 (N_12207,N_7150,N_7302);
nor U12208 (N_12208,N_7885,N_5199);
nand U12209 (N_12209,N_8704,N_8295);
xor U12210 (N_12210,N_7183,N_8497);
xnor U12211 (N_12211,N_8017,N_9520);
nor U12212 (N_12212,N_9415,N_9217);
nor U12213 (N_12213,N_9303,N_9124);
nor U12214 (N_12214,N_7721,N_9726);
or U12215 (N_12215,N_6732,N_5099);
nand U12216 (N_12216,N_9820,N_6975);
or U12217 (N_12217,N_6156,N_9190);
nand U12218 (N_12218,N_9433,N_9908);
nand U12219 (N_12219,N_6993,N_6310);
nand U12220 (N_12220,N_6726,N_8932);
nand U12221 (N_12221,N_5256,N_9036);
xor U12222 (N_12222,N_6334,N_7205);
and U12223 (N_12223,N_9445,N_7876);
xor U12224 (N_12224,N_8506,N_5796);
nor U12225 (N_12225,N_7506,N_5607);
nor U12226 (N_12226,N_8856,N_6986);
nand U12227 (N_12227,N_9421,N_8532);
or U12228 (N_12228,N_8091,N_8321);
nor U12229 (N_12229,N_8500,N_7890);
nor U12230 (N_12230,N_6242,N_9547);
or U12231 (N_12231,N_8512,N_6232);
nand U12232 (N_12232,N_7391,N_5061);
or U12233 (N_12233,N_5305,N_7752);
or U12234 (N_12234,N_8425,N_8714);
nor U12235 (N_12235,N_8108,N_5060);
nand U12236 (N_12236,N_9645,N_7996);
and U12237 (N_12237,N_6783,N_8942);
nand U12238 (N_12238,N_7538,N_6048);
nor U12239 (N_12239,N_5643,N_6789);
nor U12240 (N_12240,N_8011,N_5445);
nor U12241 (N_12241,N_6015,N_5847);
and U12242 (N_12242,N_7865,N_8259);
or U12243 (N_12243,N_5496,N_5527);
nor U12244 (N_12244,N_5894,N_8448);
or U12245 (N_12245,N_8845,N_6239);
or U12246 (N_12246,N_5965,N_6711);
nor U12247 (N_12247,N_8578,N_8419);
xor U12248 (N_12248,N_5310,N_8753);
xor U12249 (N_12249,N_5335,N_7693);
nand U12250 (N_12250,N_7723,N_6535);
nand U12251 (N_12251,N_9470,N_7523);
nor U12252 (N_12252,N_6776,N_7605);
or U12253 (N_12253,N_5676,N_9145);
nor U12254 (N_12254,N_9469,N_6537);
and U12255 (N_12255,N_5097,N_8750);
and U12256 (N_12256,N_9084,N_7631);
nand U12257 (N_12257,N_6482,N_9601);
nand U12258 (N_12258,N_7786,N_8023);
nand U12259 (N_12259,N_7939,N_5804);
and U12260 (N_12260,N_8756,N_9710);
xor U12261 (N_12261,N_9070,N_9996);
nor U12262 (N_12262,N_8338,N_9113);
nor U12263 (N_12263,N_6770,N_7700);
nand U12264 (N_12264,N_9617,N_7464);
and U12265 (N_12265,N_8111,N_5139);
xor U12266 (N_12266,N_8947,N_9986);
and U12267 (N_12267,N_5068,N_8526);
nand U12268 (N_12268,N_7362,N_6650);
or U12269 (N_12269,N_6106,N_9034);
nor U12270 (N_12270,N_9805,N_5668);
nor U12271 (N_12271,N_6933,N_7023);
or U12272 (N_12272,N_7926,N_6070);
and U12273 (N_12273,N_6710,N_5350);
nand U12274 (N_12274,N_9886,N_6064);
and U12275 (N_12275,N_9935,N_5121);
nor U12276 (N_12276,N_7957,N_5421);
nor U12277 (N_12277,N_8323,N_8320);
nand U12278 (N_12278,N_6511,N_9921);
xnor U12279 (N_12279,N_9997,N_9350);
and U12280 (N_12280,N_9462,N_9186);
xor U12281 (N_12281,N_5077,N_7250);
xnor U12282 (N_12282,N_8944,N_7534);
and U12283 (N_12283,N_5598,N_8190);
and U12284 (N_12284,N_8099,N_5204);
or U12285 (N_12285,N_6786,N_9900);
and U12286 (N_12286,N_9121,N_9883);
nor U12287 (N_12287,N_9484,N_5572);
nand U12288 (N_12288,N_9477,N_7684);
or U12289 (N_12289,N_7912,N_5960);
and U12290 (N_12290,N_5703,N_7004);
and U12291 (N_12291,N_5211,N_7243);
xnor U12292 (N_12292,N_7948,N_5149);
or U12293 (N_12293,N_5743,N_5724);
and U12294 (N_12294,N_7776,N_7018);
nand U12295 (N_12295,N_5778,N_8214);
xor U12296 (N_12296,N_8683,N_7259);
xnor U12297 (N_12297,N_6110,N_8761);
or U12298 (N_12298,N_9972,N_6341);
nand U12299 (N_12299,N_6521,N_8085);
or U12300 (N_12300,N_7816,N_8486);
xnor U12301 (N_12301,N_6548,N_8797);
nand U12302 (N_12302,N_7451,N_9158);
nor U12303 (N_12303,N_6984,N_5628);
nand U12304 (N_12304,N_8855,N_9895);
or U12305 (N_12305,N_5757,N_8638);
nand U12306 (N_12306,N_8110,N_9512);
and U12307 (N_12307,N_7129,N_9337);
nor U12308 (N_12308,N_6228,N_8551);
xor U12309 (N_12309,N_9956,N_7139);
nor U12310 (N_12310,N_6737,N_6624);
and U12311 (N_12311,N_6250,N_5046);
nand U12312 (N_12312,N_7509,N_7943);
xor U12313 (N_12313,N_9095,N_9889);
nor U12314 (N_12314,N_5744,N_9479);
xnor U12315 (N_12315,N_6871,N_5017);
and U12316 (N_12316,N_6727,N_8279);
nor U12317 (N_12317,N_7718,N_7500);
xor U12318 (N_12318,N_5209,N_6943);
nor U12319 (N_12319,N_9709,N_6883);
nor U12320 (N_12320,N_8456,N_8591);
nand U12321 (N_12321,N_6605,N_5727);
nand U12322 (N_12322,N_6396,N_9000);
xor U12323 (N_12323,N_7429,N_6389);
and U12324 (N_12324,N_6186,N_6622);
nor U12325 (N_12325,N_6408,N_7871);
and U12326 (N_12326,N_5092,N_6631);
and U12327 (N_12327,N_5003,N_7016);
nand U12328 (N_12328,N_5885,N_9961);
nand U12329 (N_12329,N_7005,N_7450);
nand U12330 (N_12330,N_8600,N_8764);
and U12331 (N_12331,N_9783,N_7918);
and U12332 (N_12332,N_9355,N_8495);
and U12333 (N_12333,N_9128,N_9676);
nand U12334 (N_12334,N_8803,N_6989);
nor U12335 (N_12335,N_5780,N_6283);
nand U12336 (N_12336,N_7116,N_9310);
nor U12337 (N_12337,N_9788,N_8810);
nand U12338 (N_12338,N_5182,N_8829);
nand U12339 (N_12339,N_8809,N_6030);
xnor U12340 (N_12340,N_9388,N_9689);
xnor U12341 (N_12341,N_6909,N_9135);
nor U12342 (N_12342,N_5859,N_8718);
nand U12343 (N_12343,N_9718,N_5388);
nand U12344 (N_12344,N_7709,N_6623);
nand U12345 (N_12345,N_5596,N_8569);
nor U12346 (N_12346,N_5519,N_8254);
nor U12347 (N_12347,N_5786,N_6962);
or U12348 (N_12348,N_7820,N_8504);
nand U12349 (N_12349,N_6161,N_6076);
or U12350 (N_12350,N_6809,N_8118);
nand U12351 (N_12351,N_7296,N_6005);
nand U12352 (N_12352,N_9218,N_9754);
or U12353 (N_12353,N_5091,N_8298);
nand U12354 (N_12354,N_5532,N_5125);
and U12355 (N_12355,N_8869,N_9276);
nand U12356 (N_12356,N_8102,N_5136);
or U12357 (N_12357,N_7944,N_8801);
or U12358 (N_12358,N_9662,N_7481);
nand U12359 (N_12359,N_9185,N_6074);
or U12360 (N_12360,N_7319,N_6374);
nand U12361 (N_12361,N_5487,N_9237);
and U12362 (N_12362,N_6567,N_6209);
nor U12363 (N_12363,N_5407,N_6258);
and U12364 (N_12364,N_5152,N_8166);
and U12365 (N_12365,N_9850,N_8018);
xor U12366 (N_12366,N_5479,N_8779);
nand U12367 (N_12367,N_5447,N_5223);
xor U12368 (N_12368,N_8263,N_6073);
nand U12369 (N_12369,N_7035,N_6648);
nor U12370 (N_12370,N_5327,N_7372);
nor U12371 (N_12371,N_5461,N_7633);
or U12372 (N_12372,N_9691,N_9697);
nand U12373 (N_12373,N_6175,N_9945);
nor U12374 (N_12374,N_6832,N_6130);
nand U12375 (N_12375,N_6184,N_5515);
nand U12376 (N_12376,N_7895,N_7015);
and U12377 (N_12377,N_5565,N_9807);
or U12378 (N_12378,N_6942,N_8093);
nand U12379 (N_12379,N_6280,N_8070);
and U12380 (N_12380,N_7376,N_7665);
and U12381 (N_12381,N_5393,N_6430);
or U12382 (N_12382,N_8278,N_8447);
nor U12383 (N_12383,N_9607,N_6563);
nor U12384 (N_12384,N_8738,N_7753);
nor U12385 (N_12385,N_7862,N_5770);
or U12386 (N_12386,N_7195,N_9317);
or U12387 (N_12387,N_5764,N_5958);
nand U12388 (N_12388,N_8152,N_7600);
nand U12389 (N_12389,N_8766,N_8113);
or U12390 (N_12390,N_6881,N_6466);
nand U12391 (N_12391,N_6707,N_5009);
nand U12392 (N_12392,N_6778,N_5601);
nor U12393 (N_12393,N_6851,N_9542);
nor U12394 (N_12394,N_5942,N_7956);
nor U12395 (N_12395,N_9319,N_5756);
and U12396 (N_12396,N_9853,N_5168);
nor U12397 (N_12397,N_8548,N_6580);
or U12398 (N_12398,N_6265,N_8090);
nand U12399 (N_12399,N_7301,N_8540);
or U12400 (N_12400,N_5964,N_8860);
nand U12401 (N_12401,N_7929,N_7123);
and U12402 (N_12402,N_5537,N_5297);
nand U12403 (N_12403,N_5059,N_6728);
xor U12404 (N_12404,N_9665,N_6911);
and U12405 (N_12405,N_8016,N_9291);
or U12406 (N_12406,N_9579,N_7022);
nor U12407 (N_12407,N_7313,N_5455);
nor U12408 (N_12408,N_7351,N_9383);
and U12409 (N_12409,N_6034,N_6642);
and U12410 (N_12410,N_5723,N_6780);
nor U12411 (N_12411,N_8474,N_9252);
nor U12412 (N_12412,N_6243,N_6669);
nand U12413 (N_12413,N_7629,N_9509);
and U12414 (N_12414,N_5263,N_6976);
nand U12415 (N_12415,N_7042,N_5134);
or U12416 (N_12416,N_7937,N_8400);
nor U12417 (N_12417,N_6681,N_8879);
or U12418 (N_12418,N_6626,N_8178);
nand U12419 (N_12419,N_8523,N_9636);
nor U12420 (N_12420,N_5955,N_7497);
nand U12421 (N_12421,N_7511,N_9641);
nor U12422 (N_12422,N_7060,N_5013);
nor U12423 (N_12423,N_5096,N_9540);
or U12424 (N_12424,N_6236,N_8062);
xor U12425 (N_12425,N_6894,N_7434);
and U12426 (N_12426,N_6977,N_9897);
nor U12427 (N_12427,N_7145,N_5391);
nand U12428 (N_12428,N_8796,N_7211);
and U12429 (N_12429,N_7086,N_5843);
nand U12430 (N_12430,N_8010,N_7166);
or U12431 (N_12431,N_8340,N_6643);
nand U12432 (N_12432,N_9667,N_8008);
nand U12433 (N_12433,N_6302,N_8760);
or U12434 (N_12434,N_7818,N_5239);
or U12435 (N_12435,N_8925,N_9140);
nand U12436 (N_12436,N_6826,N_7384);
nand U12437 (N_12437,N_8327,N_8454);
or U12438 (N_12438,N_6392,N_6553);
or U12439 (N_12439,N_6802,N_5698);
and U12440 (N_12440,N_8012,N_8161);
nand U12441 (N_12441,N_8566,N_5581);
and U12442 (N_12442,N_7216,N_7617);
or U12443 (N_12443,N_5789,N_9389);
and U12444 (N_12444,N_9610,N_7563);
nor U12445 (N_12445,N_8167,N_9690);
and U12446 (N_12446,N_9126,N_6502);
nor U12447 (N_12447,N_7732,N_5065);
and U12448 (N_12448,N_5836,N_7881);
or U12449 (N_12449,N_6318,N_8905);
or U12450 (N_12450,N_5794,N_7290);
nor U12451 (N_12451,N_7638,N_9981);
nand U12452 (N_12452,N_8804,N_7840);
or U12453 (N_12453,N_7763,N_9420);
nor U12454 (N_12454,N_8977,N_8605);
nand U12455 (N_12455,N_5275,N_9832);
or U12456 (N_12456,N_9768,N_5339);
and U12457 (N_12457,N_6594,N_8912);
or U12458 (N_12458,N_9753,N_6240);
and U12459 (N_12459,N_8826,N_6932);
nor U12460 (N_12460,N_7278,N_8823);
nor U12461 (N_12461,N_6333,N_9654);
xnor U12462 (N_12462,N_6372,N_8379);
nand U12463 (N_12463,N_9205,N_8674);
xor U12464 (N_12464,N_5989,N_8009);
and U12465 (N_12465,N_8239,N_5680);
nor U12466 (N_12466,N_5647,N_8007);
nor U12467 (N_12467,N_6097,N_6424);
xnor U12468 (N_12468,N_7153,N_6195);
and U12469 (N_12469,N_8317,N_7324);
and U12470 (N_12470,N_5542,N_9779);
xor U12471 (N_12471,N_5436,N_5267);
nand U12472 (N_12472,N_6980,N_9863);
nor U12473 (N_12473,N_9964,N_8859);
nand U12474 (N_12474,N_8312,N_6995);
and U12475 (N_12475,N_7049,N_7923);
nor U12476 (N_12476,N_7186,N_5926);
or U12477 (N_12477,N_6544,N_6758);
or U12478 (N_12478,N_8370,N_9902);
or U12479 (N_12479,N_6202,N_8640);
xnor U12480 (N_12480,N_8037,N_8882);
nand U12481 (N_12481,N_7101,N_9799);
or U12482 (N_12482,N_6965,N_6509);
nand U12483 (N_12483,N_9661,N_9500);
nand U12484 (N_12484,N_5928,N_8781);
xnor U12485 (N_12485,N_9353,N_7092);
or U12486 (N_12486,N_9613,N_8065);
or U12487 (N_12487,N_7791,N_5557);
xor U12488 (N_12488,N_5441,N_5398);
or U12489 (N_12489,N_7712,N_7736);
or U12490 (N_12490,N_9426,N_7070);
and U12491 (N_12491,N_6722,N_8863);
xnor U12492 (N_12492,N_5522,N_5897);
and U12493 (N_12493,N_6640,N_8200);
and U12494 (N_12494,N_5528,N_5737);
or U12495 (N_12495,N_7952,N_9465);
nor U12496 (N_12496,N_8299,N_5048);
and U12497 (N_12497,N_7989,N_9506);
nor U12498 (N_12498,N_9944,N_6819);
and U12499 (N_12499,N_6639,N_5948);
or U12500 (N_12500,N_6489,N_7308);
nand U12501 (N_12501,N_5841,N_7824);
nand U12502 (N_12502,N_8421,N_7544);
nor U12503 (N_12503,N_9519,N_8902);
and U12504 (N_12504,N_6953,N_9466);
xor U12505 (N_12505,N_9148,N_9546);
nor U12506 (N_12506,N_5340,N_5234);
nor U12507 (N_12507,N_5684,N_7953);
and U12508 (N_12508,N_9868,N_5776);
and U12509 (N_12509,N_9343,N_7926);
nand U12510 (N_12510,N_5487,N_9298);
nand U12511 (N_12511,N_5306,N_8441);
nand U12512 (N_12512,N_8427,N_8067);
or U12513 (N_12513,N_5092,N_6153);
nand U12514 (N_12514,N_6876,N_5792);
and U12515 (N_12515,N_5158,N_6392);
nor U12516 (N_12516,N_5145,N_8988);
nor U12517 (N_12517,N_5154,N_8932);
and U12518 (N_12518,N_8993,N_8874);
and U12519 (N_12519,N_5067,N_5197);
and U12520 (N_12520,N_8284,N_5006);
and U12521 (N_12521,N_8343,N_7026);
and U12522 (N_12522,N_8034,N_7568);
nand U12523 (N_12523,N_9049,N_7924);
nor U12524 (N_12524,N_9741,N_5458);
or U12525 (N_12525,N_6757,N_6522);
xnor U12526 (N_12526,N_8018,N_8859);
or U12527 (N_12527,N_6481,N_9228);
nor U12528 (N_12528,N_8633,N_8383);
nand U12529 (N_12529,N_9101,N_7717);
or U12530 (N_12530,N_6955,N_8564);
or U12531 (N_12531,N_9177,N_6678);
or U12532 (N_12532,N_9966,N_9167);
nand U12533 (N_12533,N_9551,N_9033);
nor U12534 (N_12534,N_7637,N_9189);
or U12535 (N_12535,N_8521,N_9544);
and U12536 (N_12536,N_7713,N_6513);
xnor U12537 (N_12537,N_6925,N_6869);
nand U12538 (N_12538,N_6489,N_7920);
nor U12539 (N_12539,N_8254,N_8865);
or U12540 (N_12540,N_8236,N_8962);
xnor U12541 (N_12541,N_6412,N_8444);
or U12542 (N_12542,N_8534,N_8103);
and U12543 (N_12543,N_8186,N_9920);
nand U12544 (N_12544,N_5854,N_6921);
xnor U12545 (N_12545,N_6130,N_6054);
nor U12546 (N_12546,N_6812,N_5544);
xnor U12547 (N_12547,N_7656,N_7806);
or U12548 (N_12548,N_5823,N_9970);
nand U12549 (N_12549,N_8410,N_6778);
and U12550 (N_12550,N_5655,N_6374);
nor U12551 (N_12551,N_9839,N_7222);
or U12552 (N_12552,N_6211,N_8513);
nand U12553 (N_12553,N_7687,N_8627);
nor U12554 (N_12554,N_8545,N_9496);
nor U12555 (N_12555,N_9992,N_6568);
and U12556 (N_12556,N_9122,N_8620);
nand U12557 (N_12557,N_7383,N_6147);
nand U12558 (N_12558,N_6710,N_9871);
nand U12559 (N_12559,N_5525,N_9215);
and U12560 (N_12560,N_5330,N_5555);
or U12561 (N_12561,N_7046,N_6728);
or U12562 (N_12562,N_8236,N_9000);
nand U12563 (N_12563,N_8245,N_9911);
or U12564 (N_12564,N_5976,N_5066);
nor U12565 (N_12565,N_9001,N_5210);
nand U12566 (N_12566,N_8676,N_9662);
or U12567 (N_12567,N_8928,N_6096);
xor U12568 (N_12568,N_6206,N_6907);
or U12569 (N_12569,N_5388,N_6558);
or U12570 (N_12570,N_9049,N_8647);
and U12571 (N_12571,N_8419,N_8133);
nand U12572 (N_12572,N_7388,N_5097);
and U12573 (N_12573,N_7070,N_9258);
or U12574 (N_12574,N_8818,N_7791);
nor U12575 (N_12575,N_7318,N_6401);
and U12576 (N_12576,N_9546,N_9052);
or U12577 (N_12577,N_8503,N_5938);
or U12578 (N_12578,N_8668,N_7278);
nand U12579 (N_12579,N_6739,N_7007);
nor U12580 (N_12580,N_9717,N_9048);
and U12581 (N_12581,N_7880,N_7932);
nor U12582 (N_12582,N_6154,N_5347);
nand U12583 (N_12583,N_9090,N_7791);
nor U12584 (N_12584,N_5831,N_8946);
nor U12585 (N_12585,N_5940,N_5094);
xor U12586 (N_12586,N_6145,N_9467);
nor U12587 (N_12587,N_5049,N_8314);
and U12588 (N_12588,N_6552,N_7701);
and U12589 (N_12589,N_7980,N_6503);
and U12590 (N_12590,N_7668,N_8696);
nor U12591 (N_12591,N_6941,N_8749);
nand U12592 (N_12592,N_6754,N_6115);
and U12593 (N_12593,N_8578,N_5829);
and U12594 (N_12594,N_7696,N_7441);
or U12595 (N_12595,N_6968,N_9171);
and U12596 (N_12596,N_7759,N_5201);
nand U12597 (N_12597,N_7283,N_9285);
nor U12598 (N_12598,N_8185,N_7608);
xor U12599 (N_12599,N_6423,N_5725);
or U12600 (N_12600,N_9700,N_7998);
or U12601 (N_12601,N_8645,N_5526);
nor U12602 (N_12602,N_9691,N_5303);
nand U12603 (N_12603,N_6213,N_9096);
nand U12604 (N_12604,N_9900,N_6380);
and U12605 (N_12605,N_9561,N_6096);
nand U12606 (N_12606,N_8766,N_7480);
nor U12607 (N_12607,N_9329,N_7420);
or U12608 (N_12608,N_7806,N_5561);
nor U12609 (N_12609,N_5018,N_6528);
xor U12610 (N_12610,N_7514,N_6289);
xnor U12611 (N_12611,N_7362,N_5603);
and U12612 (N_12612,N_8230,N_6970);
nand U12613 (N_12613,N_6836,N_7760);
or U12614 (N_12614,N_5467,N_6529);
nor U12615 (N_12615,N_5924,N_6190);
and U12616 (N_12616,N_7992,N_7563);
nor U12617 (N_12617,N_5436,N_8965);
and U12618 (N_12618,N_7349,N_9402);
and U12619 (N_12619,N_5323,N_7017);
and U12620 (N_12620,N_7358,N_5360);
nand U12621 (N_12621,N_5240,N_7289);
nand U12622 (N_12622,N_8600,N_9005);
or U12623 (N_12623,N_8251,N_8843);
nand U12624 (N_12624,N_7078,N_6867);
xor U12625 (N_12625,N_7888,N_9776);
and U12626 (N_12626,N_9672,N_9514);
or U12627 (N_12627,N_5662,N_7857);
and U12628 (N_12628,N_5230,N_8294);
nor U12629 (N_12629,N_7845,N_8542);
nor U12630 (N_12630,N_7441,N_6532);
or U12631 (N_12631,N_8264,N_5079);
nor U12632 (N_12632,N_9097,N_5298);
or U12633 (N_12633,N_6998,N_6579);
nor U12634 (N_12634,N_6758,N_5992);
or U12635 (N_12635,N_8328,N_8159);
or U12636 (N_12636,N_9048,N_5140);
or U12637 (N_12637,N_7341,N_9517);
and U12638 (N_12638,N_5479,N_8695);
or U12639 (N_12639,N_7062,N_8518);
and U12640 (N_12640,N_9824,N_6005);
nand U12641 (N_12641,N_9127,N_5695);
or U12642 (N_12642,N_7799,N_9661);
xnor U12643 (N_12643,N_7991,N_6081);
and U12644 (N_12644,N_8911,N_7100);
nand U12645 (N_12645,N_5694,N_5927);
xor U12646 (N_12646,N_9449,N_8429);
or U12647 (N_12647,N_8159,N_8878);
nor U12648 (N_12648,N_7507,N_7020);
nand U12649 (N_12649,N_6427,N_9120);
or U12650 (N_12650,N_5386,N_9621);
or U12651 (N_12651,N_5712,N_5793);
nand U12652 (N_12652,N_9413,N_8228);
nor U12653 (N_12653,N_8308,N_6503);
nor U12654 (N_12654,N_6403,N_8441);
nor U12655 (N_12655,N_6852,N_8746);
nand U12656 (N_12656,N_7008,N_8047);
xor U12657 (N_12657,N_5044,N_6741);
nor U12658 (N_12658,N_9516,N_8589);
nand U12659 (N_12659,N_8503,N_5392);
nor U12660 (N_12660,N_6485,N_6326);
nor U12661 (N_12661,N_5168,N_5085);
or U12662 (N_12662,N_5804,N_7960);
or U12663 (N_12663,N_5057,N_6240);
and U12664 (N_12664,N_8285,N_6781);
or U12665 (N_12665,N_9784,N_7880);
nand U12666 (N_12666,N_6545,N_5753);
nor U12667 (N_12667,N_7519,N_9425);
nor U12668 (N_12668,N_5322,N_5140);
or U12669 (N_12669,N_7981,N_9369);
or U12670 (N_12670,N_5545,N_5212);
nor U12671 (N_12671,N_9457,N_8555);
nand U12672 (N_12672,N_8385,N_5389);
xnor U12673 (N_12673,N_5036,N_5392);
or U12674 (N_12674,N_5417,N_6453);
nand U12675 (N_12675,N_7284,N_9407);
or U12676 (N_12676,N_9487,N_6971);
or U12677 (N_12677,N_5458,N_7861);
nand U12678 (N_12678,N_5391,N_9871);
or U12679 (N_12679,N_8100,N_5893);
nor U12680 (N_12680,N_8509,N_6153);
or U12681 (N_12681,N_5423,N_8219);
xor U12682 (N_12682,N_9946,N_5108);
and U12683 (N_12683,N_6504,N_9699);
nor U12684 (N_12684,N_6802,N_9416);
and U12685 (N_12685,N_5788,N_6848);
and U12686 (N_12686,N_8350,N_9385);
and U12687 (N_12687,N_7247,N_6859);
and U12688 (N_12688,N_9127,N_8482);
and U12689 (N_12689,N_8342,N_5451);
nand U12690 (N_12690,N_6847,N_7955);
or U12691 (N_12691,N_6647,N_9123);
or U12692 (N_12692,N_8937,N_8039);
and U12693 (N_12693,N_5816,N_9545);
and U12694 (N_12694,N_9335,N_8642);
and U12695 (N_12695,N_6877,N_8571);
nand U12696 (N_12696,N_8117,N_9298);
and U12697 (N_12697,N_7939,N_6156);
xnor U12698 (N_12698,N_9056,N_9931);
nor U12699 (N_12699,N_8839,N_9295);
nand U12700 (N_12700,N_8449,N_7596);
or U12701 (N_12701,N_9092,N_9366);
nand U12702 (N_12702,N_7593,N_7749);
nand U12703 (N_12703,N_9859,N_5854);
xor U12704 (N_12704,N_6827,N_9702);
and U12705 (N_12705,N_5560,N_7925);
nor U12706 (N_12706,N_8641,N_9445);
or U12707 (N_12707,N_9756,N_6129);
nor U12708 (N_12708,N_8304,N_8650);
nor U12709 (N_12709,N_8397,N_5678);
nor U12710 (N_12710,N_8150,N_5816);
and U12711 (N_12711,N_9711,N_7726);
and U12712 (N_12712,N_7878,N_9020);
or U12713 (N_12713,N_6251,N_6159);
nor U12714 (N_12714,N_6196,N_7407);
nor U12715 (N_12715,N_9493,N_6329);
and U12716 (N_12716,N_6828,N_5954);
and U12717 (N_12717,N_6343,N_9966);
xor U12718 (N_12718,N_9350,N_9443);
nand U12719 (N_12719,N_7011,N_8671);
and U12720 (N_12720,N_9829,N_5946);
nand U12721 (N_12721,N_9156,N_5438);
xnor U12722 (N_12722,N_9109,N_8526);
nor U12723 (N_12723,N_6981,N_9921);
and U12724 (N_12724,N_9692,N_8587);
nand U12725 (N_12725,N_8733,N_9991);
nand U12726 (N_12726,N_8970,N_6427);
xor U12727 (N_12727,N_8064,N_6845);
or U12728 (N_12728,N_8383,N_9676);
nand U12729 (N_12729,N_9320,N_9036);
nor U12730 (N_12730,N_6779,N_5060);
or U12731 (N_12731,N_7886,N_9619);
nand U12732 (N_12732,N_5707,N_9941);
nand U12733 (N_12733,N_5046,N_7181);
or U12734 (N_12734,N_5741,N_6306);
or U12735 (N_12735,N_6134,N_9454);
nor U12736 (N_12736,N_7336,N_7702);
and U12737 (N_12737,N_7835,N_5251);
nand U12738 (N_12738,N_8359,N_7643);
nor U12739 (N_12739,N_7750,N_9856);
or U12740 (N_12740,N_7855,N_7032);
nand U12741 (N_12741,N_9462,N_9123);
nand U12742 (N_12742,N_6600,N_5751);
nand U12743 (N_12743,N_7966,N_7362);
nor U12744 (N_12744,N_5381,N_7497);
or U12745 (N_12745,N_7263,N_8444);
or U12746 (N_12746,N_7876,N_7689);
and U12747 (N_12747,N_6231,N_8240);
nor U12748 (N_12748,N_9516,N_9492);
or U12749 (N_12749,N_9718,N_8130);
nand U12750 (N_12750,N_9407,N_5726);
xnor U12751 (N_12751,N_9591,N_9718);
xor U12752 (N_12752,N_6082,N_9595);
or U12753 (N_12753,N_6990,N_5640);
nand U12754 (N_12754,N_5645,N_9883);
nor U12755 (N_12755,N_7446,N_6500);
xnor U12756 (N_12756,N_8693,N_9301);
or U12757 (N_12757,N_8181,N_9387);
and U12758 (N_12758,N_9670,N_8688);
and U12759 (N_12759,N_9357,N_6306);
or U12760 (N_12760,N_6437,N_7786);
nor U12761 (N_12761,N_5998,N_8369);
xor U12762 (N_12762,N_5705,N_7966);
nor U12763 (N_12763,N_5919,N_8048);
or U12764 (N_12764,N_8981,N_7516);
nor U12765 (N_12765,N_8742,N_9905);
nor U12766 (N_12766,N_5570,N_8667);
or U12767 (N_12767,N_7142,N_9267);
xnor U12768 (N_12768,N_8761,N_6470);
or U12769 (N_12769,N_6580,N_5911);
or U12770 (N_12770,N_9975,N_7560);
and U12771 (N_12771,N_7773,N_7702);
nor U12772 (N_12772,N_8358,N_9551);
and U12773 (N_12773,N_8772,N_9335);
and U12774 (N_12774,N_9222,N_6244);
xnor U12775 (N_12775,N_7069,N_7638);
nand U12776 (N_12776,N_5701,N_6439);
nand U12777 (N_12777,N_5608,N_8940);
nand U12778 (N_12778,N_9736,N_5958);
nand U12779 (N_12779,N_8457,N_6721);
nand U12780 (N_12780,N_8810,N_8774);
nand U12781 (N_12781,N_7538,N_7587);
and U12782 (N_12782,N_5686,N_8558);
nor U12783 (N_12783,N_8109,N_7340);
nor U12784 (N_12784,N_9871,N_5411);
and U12785 (N_12785,N_8038,N_8012);
nor U12786 (N_12786,N_9189,N_5335);
nand U12787 (N_12787,N_5450,N_7360);
and U12788 (N_12788,N_6358,N_8079);
nand U12789 (N_12789,N_9676,N_8694);
nand U12790 (N_12790,N_7108,N_8059);
and U12791 (N_12791,N_7585,N_6660);
nor U12792 (N_12792,N_8603,N_9006);
or U12793 (N_12793,N_8133,N_9651);
or U12794 (N_12794,N_8501,N_8859);
nor U12795 (N_12795,N_8741,N_7418);
nor U12796 (N_12796,N_5291,N_9119);
nor U12797 (N_12797,N_8190,N_8343);
xor U12798 (N_12798,N_9104,N_9814);
and U12799 (N_12799,N_9828,N_5091);
xnor U12800 (N_12800,N_9209,N_7088);
and U12801 (N_12801,N_9039,N_6751);
xnor U12802 (N_12802,N_9353,N_7782);
xor U12803 (N_12803,N_8789,N_6990);
nor U12804 (N_12804,N_5745,N_7794);
nand U12805 (N_12805,N_7875,N_5678);
xor U12806 (N_12806,N_5053,N_5816);
and U12807 (N_12807,N_9492,N_6214);
nand U12808 (N_12808,N_8993,N_9694);
nand U12809 (N_12809,N_9645,N_5503);
or U12810 (N_12810,N_6190,N_7294);
and U12811 (N_12811,N_7174,N_6384);
or U12812 (N_12812,N_7707,N_6028);
nand U12813 (N_12813,N_9526,N_8960);
xnor U12814 (N_12814,N_8965,N_7596);
nand U12815 (N_12815,N_5765,N_6398);
nor U12816 (N_12816,N_7071,N_6093);
nor U12817 (N_12817,N_5603,N_7794);
or U12818 (N_12818,N_5466,N_8531);
or U12819 (N_12819,N_5005,N_5784);
nand U12820 (N_12820,N_6437,N_5776);
xnor U12821 (N_12821,N_7098,N_7058);
and U12822 (N_12822,N_8738,N_5952);
and U12823 (N_12823,N_5167,N_9047);
nand U12824 (N_12824,N_6179,N_7865);
nand U12825 (N_12825,N_7110,N_9014);
or U12826 (N_12826,N_7800,N_9646);
nor U12827 (N_12827,N_5095,N_8655);
and U12828 (N_12828,N_9796,N_9066);
or U12829 (N_12829,N_9982,N_9247);
nand U12830 (N_12830,N_7930,N_8427);
and U12831 (N_12831,N_7991,N_6758);
or U12832 (N_12832,N_8817,N_8126);
nand U12833 (N_12833,N_7538,N_8797);
xor U12834 (N_12834,N_9803,N_9943);
nand U12835 (N_12835,N_9179,N_8534);
and U12836 (N_12836,N_5086,N_8992);
nand U12837 (N_12837,N_8414,N_9841);
nand U12838 (N_12838,N_7268,N_6126);
or U12839 (N_12839,N_7210,N_6694);
and U12840 (N_12840,N_5244,N_7065);
nand U12841 (N_12841,N_8474,N_8757);
nand U12842 (N_12842,N_9539,N_6577);
xor U12843 (N_12843,N_6588,N_6273);
nor U12844 (N_12844,N_8640,N_5993);
nor U12845 (N_12845,N_9885,N_9513);
or U12846 (N_12846,N_6120,N_8922);
nor U12847 (N_12847,N_7644,N_8461);
or U12848 (N_12848,N_9948,N_9595);
nor U12849 (N_12849,N_7339,N_7729);
nor U12850 (N_12850,N_7312,N_7816);
nor U12851 (N_12851,N_9325,N_8065);
nand U12852 (N_12852,N_8406,N_7722);
nand U12853 (N_12853,N_8835,N_6080);
or U12854 (N_12854,N_6357,N_5657);
nor U12855 (N_12855,N_7438,N_9859);
nand U12856 (N_12856,N_6263,N_5341);
or U12857 (N_12857,N_9551,N_6793);
xor U12858 (N_12858,N_6706,N_6120);
or U12859 (N_12859,N_8797,N_8699);
nand U12860 (N_12860,N_8236,N_6613);
nand U12861 (N_12861,N_5804,N_9472);
nor U12862 (N_12862,N_7369,N_5640);
nor U12863 (N_12863,N_7417,N_9001);
nor U12864 (N_12864,N_5838,N_5624);
or U12865 (N_12865,N_9674,N_7006);
or U12866 (N_12866,N_5849,N_6659);
and U12867 (N_12867,N_8575,N_8349);
nor U12868 (N_12868,N_6331,N_9181);
and U12869 (N_12869,N_8360,N_5087);
and U12870 (N_12870,N_6492,N_8644);
and U12871 (N_12871,N_8873,N_7727);
and U12872 (N_12872,N_6397,N_7910);
or U12873 (N_12873,N_9527,N_8978);
or U12874 (N_12874,N_7785,N_9017);
and U12875 (N_12875,N_8651,N_6687);
or U12876 (N_12876,N_6920,N_5833);
nor U12877 (N_12877,N_5623,N_6042);
nor U12878 (N_12878,N_7094,N_9693);
and U12879 (N_12879,N_6210,N_5119);
or U12880 (N_12880,N_5681,N_9729);
nor U12881 (N_12881,N_7127,N_5646);
nor U12882 (N_12882,N_5238,N_5278);
and U12883 (N_12883,N_9116,N_6611);
xor U12884 (N_12884,N_8994,N_8241);
xor U12885 (N_12885,N_6663,N_9068);
and U12886 (N_12886,N_5283,N_5649);
or U12887 (N_12887,N_9633,N_7225);
nor U12888 (N_12888,N_9237,N_9735);
or U12889 (N_12889,N_6902,N_6612);
nand U12890 (N_12890,N_5869,N_7979);
nand U12891 (N_12891,N_9621,N_6472);
nor U12892 (N_12892,N_7414,N_9300);
or U12893 (N_12893,N_6662,N_9724);
or U12894 (N_12894,N_8769,N_7575);
nand U12895 (N_12895,N_6288,N_9794);
nand U12896 (N_12896,N_5549,N_9870);
nand U12897 (N_12897,N_6507,N_5404);
nor U12898 (N_12898,N_7788,N_5897);
nand U12899 (N_12899,N_5525,N_5955);
and U12900 (N_12900,N_6662,N_7185);
nand U12901 (N_12901,N_9244,N_8477);
nor U12902 (N_12902,N_5819,N_8420);
nor U12903 (N_12903,N_7140,N_9487);
and U12904 (N_12904,N_5912,N_9954);
and U12905 (N_12905,N_5859,N_5885);
nor U12906 (N_12906,N_6197,N_6687);
nand U12907 (N_12907,N_6036,N_6754);
or U12908 (N_12908,N_7559,N_8089);
nand U12909 (N_12909,N_6225,N_8391);
nor U12910 (N_12910,N_8502,N_5279);
nand U12911 (N_12911,N_7235,N_7508);
or U12912 (N_12912,N_7797,N_8162);
and U12913 (N_12913,N_5087,N_6228);
or U12914 (N_12914,N_9144,N_8716);
or U12915 (N_12915,N_7598,N_5752);
nand U12916 (N_12916,N_7316,N_7568);
nand U12917 (N_12917,N_9668,N_5989);
nor U12918 (N_12918,N_9858,N_6500);
or U12919 (N_12919,N_6546,N_7717);
and U12920 (N_12920,N_9424,N_6784);
nor U12921 (N_12921,N_8453,N_9459);
nor U12922 (N_12922,N_9864,N_9195);
or U12923 (N_12923,N_7260,N_8839);
or U12924 (N_12924,N_5880,N_5784);
nor U12925 (N_12925,N_9955,N_6054);
nand U12926 (N_12926,N_7202,N_6720);
or U12927 (N_12927,N_6035,N_5906);
and U12928 (N_12928,N_8144,N_9843);
xor U12929 (N_12929,N_6388,N_6373);
and U12930 (N_12930,N_8695,N_7780);
or U12931 (N_12931,N_9647,N_7491);
or U12932 (N_12932,N_7978,N_5677);
nand U12933 (N_12933,N_8078,N_6613);
or U12934 (N_12934,N_5081,N_9191);
and U12935 (N_12935,N_6057,N_6634);
nor U12936 (N_12936,N_6626,N_6768);
or U12937 (N_12937,N_9788,N_6757);
xnor U12938 (N_12938,N_6746,N_5878);
and U12939 (N_12939,N_6271,N_7361);
nand U12940 (N_12940,N_7375,N_6384);
xor U12941 (N_12941,N_5880,N_7280);
xor U12942 (N_12942,N_9813,N_8268);
nor U12943 (N_12943,N_5804,N_5387);
xnor U12944 (N_12944,N_9460,N_7312);
or U12945 (N_12945,N_9586,N_7168);
nor U12946 (N_12946,N_6082,N_5100);
nor U12947 (N_12947,N_5939,N_7001);
xnor U12948 (N_12948,N_7973,N_6359);
and U12949 (N_12949,N_8767,N_5152);
and U12950 (N_12950,N_7244,N_5414);
nand U12951 (N_12951,N_6613,N_7495);
and U12952 (N_12952,N_6503,N_6316);
and U12953 (N_12953,N_8352,N_6583);
nand U12954 (N_12954,N_8668,N_8772);
and U12955 (N_12955,N_9084,N_8987);
nand U12956 (N_12956,N_9164,N_9269);
or U12957 (N_12957,N_5616,N_7879);
nand U12958 (N_12958,N_9930,N_7780);
or U12959 (N_12959,N_7708,N_7429);
xor U12960 (N_12960,N_6204,N_5504);
nor U12961 (N_12961,N_7267,N_8065);
or U12962 (N_12962,N_8910,N_8657);
or U12963 (N_12963,N_8782,N_5551);
or U12964 (N_12964,N_5357,N_6895);
nand U12965 (N_12965,N_5810,N_5469);
and U12966 (N_12966,N_5012,N_6377);
nand U12967 (N_12967,N_6053,N_6605);
and U12968 (N_12968,N_5713,N_6077);
and U12969 (N_12969,N_6190,N_5153);
and U12970 (N_12970,N_5880,N_6755);
and U12971 (N_12971,N_5190,N_5249);
or U12972 (N_12972,N_8820,N_6536);
nor U12973 (N_12973,N_9944,N_9972);
xnor U12974 (N_12974,N_9940,N_6086);
and U12975 (N_12975,N_6244,N_6595);
nand U12976 (N_12976,N_5841,N_5046);
and U12977 (N_12977,N_9414,N_9478);
nor U12978 (N_12978,N_5212,N_9281);
nor U12979 (N_12979,N_6714,N_8602);
and U12980 (N_12980,N_9637,N_6498);
and U12981 (N_12981,N_7949,N_5106);
nand U12982 (N_12982,N_8428,N_9940);
or U12983 (N_12983,N_7883,N_6580);
xnor U12984 (N_12984,N_7034,N_6994);
or U12985 (N_12985,N_6664,N_6767);
or U12986 (N_12986,N_6231,N_8625);
nand U12987 (N_12987,N_5316,N_9227);
nor U12988 (N_12988,N_6942,N_6587);
nor U12989 (N_12989,N_8312,N_6338);
nor U12990 (N_12990,N_7239,N_8082);
nand U12991 (N_12991,N_9674,N_5845);
nor U12992 (N_12992,N_8757,N_7859);
nor U12993 (N_12993,N_5934,N_6695);
or U12994 (N_12994,N_5381,N_5995);
nor U12995 (N_12995,N_6020,N_5248);
nor U12996 (N_12996,N_5696,N_9653);
nor U12997 (N_12997,N_8975,N_6626);
nand U12998 (N_12998,N_6230,N_9283);
nand U12999 (N_12999,N_8472,N_6012);
nand U13000 (N_13000,N_7760,N_8686);
or U13001 (N_13001,N_6398,N_5953);
or U13002 (N_13002,N_6465,N_7010);
nor U13003 (N_13003,N_9755,N_5463);
nand U13004 (N_13004,N_6953,N_7902);
xor U13005 (N_13005,N_7770,N_9513);
and U13006 (N_13006,N_9721,N_9490);
nor U13007 (N_13007,N_7659,N_8447);
nor U13008 (N_13008,N_5655,N_6061);
xnor U13009 (N_13009,N_9535,N_5903);
nand U13010 (N_13010,N_9196,N_7125);
and U13011 (N_13011,N_9556,N_8789);
nand U13012 (N_13012,N_9628,N_8027);
and U13013 (N_13013,N_6983,N_7639);
and U13014 (N_13014,N_5322,N_5585);
xor U13015 (N_13015,N_8771,N_9286);
nand U13016 (N_13016,N_8549,N_5044);
and U13017 (N_13017,N_5752,N_5879);
nand U13018 (N_13018,N_8150,N_8412);
nor U13019 (N_13019,N_5251,N_9587);
nand U13020 (N_13020,N_5876,N_5110);
nand U13021 (N_13021,N_5521,N_5718);
and U13022 (N_13022,N_9472,N_7173);
nand U13023 (N_13023,N_6585,N_5555);
nor U13024 (N_13024,N_7744,N_6636);
and U13025 (N_13025,N_6117,N_6915);
nor U13026 (N_13026,N_8248,N_9848);
nand U13027 (N_13027,N_7718,N_7115);
and U13028 (N_13028,N_8471,N_7532);
and U13029 (N_13029,N_8045,N_5865);
nor U13030 (N_13030,N_5535,N_9766);
nor U13031 (N_13031,N_7564,N_8436);
or U13032 (N_13032,N_8041,N_7928);
xnor U13033 (N_13033,N_7453,N_6776);
and U13034 (N_13034,N_6443,N_5806);
nand U13035 (N_13035,N_5361,N_7580);
or U13036 (N_13036,N_9904,N_5832);
nand U13037 (N_13037,N_6307,N_5588);
nor U13038 (N_13038,N_6284,N_6047);
or U13039 (N_13039,N_9646,N_6086);
nor U13040 (N_13040,N_9074,N_7584);
nand U13041 (N_13041,N_5963,N_5761);
nand U13042 (N_13042,N_7289,N_9699);
and U13043 (N_13043,N_9429,N_7938);
xor U13044 (N_13044,N_5175,N_7420);
or U13045 (N_13045,N_7937,N_7793);
or U13046 (N_13046,N_9613,N_7085);
nor U13047 (N_13047,N_9697,N_7650);
or U13048 (N_13048,N_5338,N_6107);
nor U13049 (N_13049,N_8071,N_8005);
and U13050 (N_13050,N_8135,N_7112);
or U13051 (N_13051,N_7949,N_8775);
nand U13052 (N_13052,N_5634,N_8305);
nand U13053 (N_13053,N_6910,N_5066);
nor U13054 (N_13054,N_6906,N_7944);
or U13055 (N_13055,N_5845,N_7211);
and U13056 (N_13056,N_5903,N_5902);
nor U13057 (N_13057,N_6847,N_6580);
nor U13058 (N_13058,N_9465,N_7708);
nor U13059 (N_13059,N_7785,N_8366);
nor U13060 (N_13060,N_9418,N_6013);
nor U13061 (N_13061,N_6299,N_8941);
nand U13062 (N_13062,N_7732,N_7161);
nor U13063 (N_13063,N_7986,N_9336);
and U13064 (N_13064,N_5657,N_7458);
or U13065 (N_13065,N_5248,N_6824);
and U13066 (N_13066,N_8606,N_9320);
nor U13067 (N_13067,N_8178,N_7036);
nand U13068 (N_13068,N_5582,N_5977);
nor U13069 (N_13069,N_8521,N_7724);
or U13070 (N_13070,N_5225,N_5151);
and U13071 (N_13071,N_8622,N_9298);
xnor U13072 (N_13072,N_7804,N_9439);
or U13073 (N_13073,N_6793,N_9695);
and U13074 (N_13074,N_7428,N_9567);
nand U13075 (N_13075,N_9449,N_7809);
nor U13076 (N_13076,N_9758,N_9985);
nor U13077 (N_13077,N_6931,N_8168);
or U13078 (N_13078,N_6656,N_9678);
and U13079 (N_13079,N_5724,N_9096);
nor U13080 (N_13080,N_7135,N_8625);
and U13081 (N_13081,N_9980,N_8670);
nor U13082 (N_13082,N_8254,N_9054);
or U13083 (N_13083,N_7587,N_8544);
or U13084 (N_13084,N_5241,N_6760);
or U13085 (N_13085,N_8817,N_6643);
nand U13086 (N_13086,N_7556,N_5952);
or U13087 (N_13087,N_5182,N_8758);
xnor U13088 (N_13088,N_7740,N_9773);
or U13089 (N_13089,N_9103,N_5869);
xnor U13090 (N_13090,N_5837,N_9589);
nor U13091 (N_13091,N_8305,N_7523);
xor U13092 (N_13092,N_6752,N_7096);
and U13093 (N_13093,N_6634,N_6042);
nor U13094 (N_13094,N_6278,N_7898);
and U13095 (N_13095,N_5801,N_8944);
or U13096 (N_13096,N_8288,N_6047);
nor U13097 (N_13097,N_8524,N_6542);
and U13098 (N_13098,N_5814,N_6460);
nor U13099 (N_13099,N_9561,N_6494);
nor U13100 (N_13100,N_5109,N_6475);
xnor U13101 (N_13101,N_7926,N_8853);
and U13102 (N_13102,N_6943,N_9637);
and U13103 (N_13103,N_7952,N_9410);
or U13104 (N_13104,N_7332,N_8482);
nor U13105 (N_13105,N_8376,N_6974);
nor U13106 (N_13106,N_5767,N_5134);
and U13107 (N_13107,N_6449,N_7309);
nand U13108 (N_13108,N_9381,N_9324);
and U13109 (N_13109,N_9538,N_6820);
nor U13110 (N_13110,N_5506,N_9086);
nand U13111 (N_13111,N_5423,N_5822);
and U13112 (N_13112,N_7972,N_6100);
nor U13113 (N_13113,N_7585,N_6759);
nand U13114 (N_13114,N_9592,N_5301);
or U13115 (N_13115,N_7867,N_9088);
nor U13116 (N_13116,N_8142,N_7572);
and U13117 (N_13117,N_6360,N_7621);
or U13118 (N_13118,N_5910,N_5296);
and U13119 (N_13119,N_5720,N_8593);
nand U13120 (N_13120,N_9949,N_6434);
nor U13121 (N_13121,N_8971,N_8720);
or U13122 (N_13122,N_9143,N_8305);
nor U13123 (N_13123,N_8618,N_8809);
or U13124 (N_13124,N_6750,N_5226);
or U13125 (N_13125,N_8128,N_7935);
and U13126 (N_13126,N_7226,N_7171);
and U13127 (N_13127,N_6692,N_8587);
or U13128 (N_13128,N_5235,N_6988);
xnor U13129 (N_13129,N_5799,N_7681);
nand U13130 (N_13130,N_5047,N_9455);
or U13131 (N_13131,N_6587,N_5589);
nor U13132 (N_13132,N_7143,N_9202);
nor U13133 (N_13133,N_9395,N_8024);
nand U13134 (N_13134,N_9491,N_5215);
or U13135 (N_13135,N_6050,N_9787);
nand U13136 (N_13136,N_8547,N_7096);
nand U13137 (N_13137,N_7273,N_5355);
nand U13138 (N_13138,N_7303,N_8043);
or U13139 (N_13139,N_5361,N_6604);
nor U13140 (N_13140,N_5263,N_8564);
nor U13141 (N_13141,N_8975,N_7494);
and U13142 (N_13142,N_8785,N_5249);
and U13143 (N_13143,N_6692,N_6263);
or U13144 (N_13144,N_7784,N_5939);
or U13145 (N_13145,N_9936,N_6235);
nand U13146 (N_13146,N_9199,N_8158);
and U13147 (N_13147,N_6324,N_8591);
nand U13148 (N_13148,N_5424,N_8414);
nor U13149 (N_13149,N_8923,N_5874);
and U13150 (N_13150,N_8185,N_6461);
and U13151 (N_13151,N_8363,N_9689);
and U13152 (N_13152,N_6708,N_6971);
or U13153 (N_13153,N_9009,N_6021);
or U13154 (N_13154,N_7987,N_6233);
or U13155 (N_13155,N_8141,N_6198);
or U13156 (N_13156,N_6119,N_8580);
nor U13157 (N_13157,N_7586,N_7798);
nand U13158 (N_13158,N_5954,N_7177);
or U13159 (N_13159,N_5250,N_9232);
nand U13160 (N_13160,N_6978,N_5190);
nand U13161 (N_13161,N_5227,N_7462);
and U13162 (N_13162,N_5162,N_8026);
nor U13163 (N_13163,N_8284,N_9029);
and U13164 (N_13164,N_8182,N_6103);
and U13165 (N_13165,N_7144,N_8156);
and U13166 (N_13166,N_8935,N_5920);
or U13167 (N_13167,N_9504,N_8775);
nor U13168 (N_13168,N_9654,N_5518);
xor U13169 (N_13169,N_8645,N_8763);
nand U13170 (N_13170,N_6159,N_9724);
and U13171 (N_13171,N_9017,N_9876);
nor U13172 (N_13172,N_6190,N_7146);
and U13173 (N_13173,N_8754,N_8460);
nand U13174 (N_13174,N_5328,N_8403);
nor U13175 (N_13175,N_7058,N_5234);
and U13176 (N_13176,N_9752,N_9305);
or U13177 (N_13177,N_8885,N_5798);
or U13178 (N_13178,N_6187,N_5793);
nor U13179 (N_13179,N_5742,N_6906);
xnor U13180 (N_13180,N_6427,N_6070);
nor U13181 (N_13181,N_8436,N_9417);
and U13182 (N_13182,N_7127,N_5371);
and U13183 (N_13183,N_6379,N_5488);
nand U13184 (N_13184,N_6299,N_6398);
nand U13185 (N_13185,N_6702,N_6146);
or U13186 (N_13186,N_5350,N_5363);
and U13187 (N_13187,N_8831,N_6785);
and U13188 (N_13188,N_9838,N_5437);
nor U13189 (N_13189,N_7666,N_7702);
or U13190 (N_13190,N_8976,N_8204);
nor U13191 (N_13191,N_7724,N_8120);
nand U13192 (N_13192,N_7632,N_6338);
or U13193 (N_13193,N_7014,N_9929);
or U13194 (N_13194,N_7854,N_7113);
nor U13195 (N_13195,N_7478,N_8799);
nor U13196 (N_13196,N_7889,N_8111);
xor U13197 (N_13197,N_8788,N_5070);
or U13198 (N_13198,N_9787,N_6672);
nor U13199 (N_13199,N_5620,N_5767);
xor U13200 (N_13200,N_5295,N_5392);
and U13201 (N_13201,N_5372,N_9239);
xnor U13202 (N_13202,N_8137,N_6439);
or U13203 (N_13203,N_6101,N_6624);
xnor U13204 (N_13204,N_6634,N_9293);
nor U13205 (N_13205,N_7834,N_5529);
or U13206 (N_13206,N_6855,N_9981);
and U13207 (N_13207,N_5871,N_8337);
or U13208 (N_13208,N_9864,N_8670);
xnor U13209 (N_13209,N_6247,N_7258);
nand U13210 (N_13210,N_9963,N_5730);
or U13211 (N_13211,N_5310,N_7195);
or U13212 (N_13212,N_7598,N_7904);
nor U13213 (N_13213,N_9753,N_6751);
or U13214 (N_13214,N_9863,N_5462);
or U13215 (N_13215,N_6917,N_9285);
xor U13216 (N_13216,N_6022,N_5185);
nand U13217 (N_13217,N_9812,N_6782);
nand U13218 (N_13218,N_6556,N_5809);
or U13219 (N_13219,N_5254,N_6340);
or U13220 (N_13220,N_9983,N_6438);
nor U13221 (N_13221,N_8354,N_8438);
xor U13222 (N_13222,N_9355,N_7750);
xor U13223 (N_13223,N_7179,N_6139);
and U13224 (N_13224,N_6561,N_8840);
nand U13225 (N_13225,N_5500,N_6060);
nor U13226 (N_13226,N_9417,N_6152);
nor U13227 (N_13227,N_6104,N_8440);
or U13228 (N_13228,N_7160,N_5489);
nor U13229 (N_13229,N_8166,N_6499);
or U13230 (N_13230,N_6578,N_5265);
xor U13231 (N_13231,N_6267,N_6325);
or U13232 (N_13232,N_9644,N_7948);
and U13233 (N_13233,N_8213,N_9567);
and U13234 (N_13234,N_9645,N_8648);
or U13235 (N_13235,N_8455,N_7068);
or U13236 (N_13236,N_9495,N_7954);
nor U13237 (N_13237,N_5586,N_9687);
and U13238 (N_13238,N_9294,N_8247);
nor U13239 (N_13239,N_9482,N_6520);
and U13240 (N_13240,N_7772,N_5302);
xnor U13241 (N_13241,N_7832,N_5481);
and U13242 (N_13242,N_7611,N_8544);
or U13243 (N_13243,N_9067,N_7294);
and U13244 (N_13244,N_9598,N_9212);
or U13245 (N_13245,N_6560,N_7531);
nand U13246 (N_13246,N_8092,N_5038);
nor U13247 (N_13247,N_5912,N_7963);
or U13248 (N_13248,N_9551,N_8741);
or U13249 (N_13249,N_8856,N_5772);
and U13250 (N_13250,N_5099,N_6554);
nand U13251 (N_13251,N_5234,N_6628);
xor U13252 (N_13252,N_6966,N_5992);
nand U13253 (N_13253,N_9904,N_6504);
nor U13254 (N_13254,N_8493,N_6919);
and U13255 (N_13255,N_5819,N_7534);
nand U13256 (N_13256,N_9099,N_9866);
or U13257 (N_13257,N_6262,N_6626);
nand U13258 (N_13258,N_7485,N_7561);
and U13259 (N_13259,N_8407,N_9652);
nand U13260 (N_13260,N_8539,N_5319);
nand U13261 (N_13261,N_7391,N_5042);
xor U13262 (N_13262,N_8351,N_6000);
xor U13263 (N_13263,N_9065,N_8522);
nor U13264 (N_13264,N_8778,N_6204);
or U13265 (N_13265,N_7349,N_6788);
xor U13266 (N_13266,N_5044,N_5643);
and U13267 (N_13267,N_6563,N_7854);
and U13268 (N_13268,N_7008,N_7912);
nor U13269 (N_13269,N_9633,N_5087);
or U13270 (N_13270,N_9333,N_5708);
nand U13271 (N_13271,N_6311,N_9623);
or U13272 (N_13272,N_9239,N_9256);
nand U13273 (N_13273,N_9760,N_8867);
and U13274 (N_13274,N_9082,N_9462);
nor U13275 (N_13275,N_9888,N_7087);
nor U13276 (N_13276,N_8379,N_7673);
nand U13277 (N_13277,N_5598,N_9784);
nand U13278 (N_13278,N_9273,N_6137);
nand U13279 (N_13279,N_6158,N_8697);
nand U13280 (N_13280,N_7148,N_5216);
and U13281 (N_13281,N_6561,N_6169);
nand U13282 (N_13282,N_5650,N_6142);
or U13283 (N_13283,N_5167,N_8419);
and U13284 (N_13284,N_9742,N_9288);
and U13285 (N_13285,N_8031,N_6596);
nand U13286 (N_13286,N_9117,N_8973);
nand U13287 (N_13287,N_6059,N_8808);
or U13288 (N_13288,N_7868,N_6362);
nand U13289 (N_13289,N_5576,N_6904);
nor U13290 (N_13290,N_5194,N_7895);
or U13291 (N_13291,N_9940,N_7516);
and U13292 (N_13292,N_7216,N_5194);
xnor U13293 (N_13293,N_9064,N_9515);
nand U13294 (N_13294,N_6842,N_8251);
and U13295 (N_13295,N_9527,N_7468);
nor U13296 (N_13296,N_8970,N_7993);
and U13297 (N_13297,N_7769,N_8155);
or U13298 (N_13298,N_7758,N_5441);
nand U13299 (N_13299,N_9555,N_8616);
and U13300 (N_13300,N_5448,N_5256);
or U13301 (N_13301,N_7292,N_6644);
or U13302 (N_13302,N_9225,N_8971);
and U13303 (N_13303,N_7075,N_7595);
and U13304 (N_13304,N_7301,N_7125);
nand U13305 (N_13305,N_7356,N_5832);
and U13306 (N_13306,N_8497,N_7240);
nand U13307 (N_13307,N_8734,N_5399);
nand U13308 (N_13308,N_9454,N_5067);
or U13309 (N_13309,N_7977,N_9141);
or U13310 (N_13310,N_9798,N_9084);
or U13311 (N_13311,N_6680,N_7073);
xor U13312 (N_13312,N_8454,N_7483);
xor U13313 (N_13313,N_6854,N_5428);
nand U13314 (N_13314,N_6860,N_9213);
nor U13315 (N_13315,N_9588,N_6403);
nor U13316 (N_13316,N_8344,N_6049);
nor U13317 (N_13317,N_5472,N_5053);
and U13318 (N_13318,N_6659,N_7421);
nor U13319 (N_13319,N_6489,N_7498);
or U13320 (N_13320,N_7785,N_8195);
nor U13321 (N_13321,N_6675,N_9859);
and U13322 (N_13322,N_7527,N_7902);
nor U13323 (N_13323,N_7110,N_5572);
or U13324 (N_13324,N_5959,N_5531);
nand U13325 (N_13325,N_9712,N_6505);
and U13326 (N_13326,N_5206,N_5335);
nor U13327 (N_13327,N_8089,N_6499);
nand U13328 (N_13328,N_6691,N_8380);
or U13329 (N_13329,N_5076,N_6604);
or U13330 (N_13330,N_9371,N_7994);
or U13331 (N_13331,N_8116,N_9791);
and U13332 (N_13332,N_8166,N_6194);
nand U13333 (N_13333,N_7792,N_8622);
nand U13334 (N_13334,N_5994,N_7739);
or U13335 (N_13335,N_5914,N_5712);
nor U13336 (N_13336,N_8607,N_5235);
xnor U13337 (N_13337,N_5232,N_6059);
nor U13338 (N_13338,N_6356,N_7175);
and U13339 (N_13339,N_6081,N_7770);
nor U13340 (N_13340,N_9442,N_9866);
nor U13341 (N_13341,N_6860,N_8355);
and U13342 (N_13342,N_8214,N_9154);
or U13343 (N_13343,N_6229,N_7168);
nor U13344 (N_13344,N_5706,N_9223);
or U13345 (N_13345,N_6425,N_6722);
nor U13346 (N_13346,N_9695,N_8901);
and U13347 (N_13347,N_9707,N_9706);
nand U13348 (N_13348,N_6469,N_9690);
nand U13349 (N_13349,N_7899,N_9485);
or U13350 (N_13350,N_6778,N_6760);
nand U13351 (N_13351,N_7991,N_5058);
nor U13352 (N_13352,N_9110,N_8482);
nor U13353 (N_13353,N_9508,N_5109);
or U13354 (N_13354,N_8316,N_8989);
nor U13355 (N_13355,N_7712,N_5362);
nand U13356 (N_13356,N_5890,N_9676);
xor U13357 (N_13357,N_9698,N_9594);
or U13358 (N_13358,N_9723,N_9493);
nand U13359 (N_13359,N_9379,N_5825);
nand U13360 (N_13360,N_8666,N_9877);
or U13361 (N_13361,N_9068,N_5637);
xor U13362 (N_13362,N_9999,N_6210);
and U13363 (N_13363,N_8626,N_6951);
nor U13364 (N_13364,N_8236,N_7508);
nor U13365 (N_13365,N_7207,N_5722);
and U13366 (N_13366,N_9752,N_7962);
or U13367 (N_13367,N_8929,N_9630);
or U13368 (N_13368,N_9258,N_6905);
nor U13369 (N_13369,N_5381,N_9450);
or U13370 (N_13370,N_7473,N_5074);
or U13371 (N_13371,N_8451,N_8994);
nand U13372 (N_13372,N_7468,N_8664);
nand U13373 (N_13373,N_7768,N_7559);
nor U13374 (N_13374,N_8462,N_7826);
nor U13375 (N_13375,N_6246,N_5400);
and U13376 (N_13376,N_5607,N_5528);
nor U13377 (N_13377,N_5293,N_9050);
and U13378 (N_13378,N_7511,N_9425);
or U13379 (N_13379,N_7306,N_5236);
or U13380 (N_13380,N_8183,N_7816);
xnor U13381 (N_13381,N_7684,N_9959);
or U13382 (N_13382,N_6957,N_6811);
nor U13383 (N_13383,N_8602,N_5193);
or U13384 (N_13384,N_7308,N_5602);
and U13385 (N_13385,N_5566,N_8094);
nor U13386 (N_13386,N_5008,N_6563);
nand U13387 (N_13387,N_5511,N_9356);
nand U13388 (N_13388,N_7496,N_8636);
and U13389 (N_13389,N_7645,N_7424);
or U13390 (N_13390,N_8529,N_8621);
xnor U13391 (N_13391,N_5861,N_5457);
and U13392 (N_13392,N_5119,N_5769);
and U13393 (N_13393,N_8603,N_7256);
nor U13394 (N_13394,N_7166,N_5958);
and U13395 (N_13395,N_9822,N_5895);
nor U13396 (N_13396,N_8871,N_6067);
nor U13397 (N_13397,N_5280,N_6495);
nor U13398 (N_13398,N_5780,N_9741);
nor U13399 (N_13399,N_5133,N_9067);
nand U13400 (N_13400,N_9202,N_6618);
nand U13401 (N_13401,N_7852,N_5222);
and U13402 (N_13402,N_5171,N_5800);
or U13403 (N_13403,N_9188,N_6777);
nor U13404 (N_13404,N_9649,N_5470);
and U13405 (N_13405,N_7059,N_8239);
nand U13406 (N_13406,N_6183,N_9821);
xnor U13407 (N_13407,N_9333,N_8385);
xnor U13408 (N_13408,N_5829,N_9391);
nor U13409 (N_13409,N_8508,N_5782);
or U13410 (N_13410,N_5090,N_7418);
and U13411 (N_13411,N_8051,N_5682);
and U13412 (N_13412,N_9960,N_5083);
xor U13413 (N_13413,N_9307,N_7918);
or U13414 (N_13414,N_6614,N_9840);
nor U13415 (N_13415,N_8836,N_7208);
or U13416 (N_13416,N_9167,N_8000);
or U13417 (N_13417,N_7081,N_9894);
nand U13418 (N_13418,N_6675,N_7572);
nor U13419 (N_13419,N_8076,N_7157);
or U13420 (N_13420,N_8149,N_8448);
and U13421 (N_13421,N_8116,N_7434);
nand U13422 (N_13422,N_8017,N_7234);
nor U13423 (N_13423,N_8278,N_9145);
or U13424 (N_13424,N_8902,N_8038);
nand U13425 (N_13425,N_6729,N_8356);
or U13426 (N_13426,N_9802,N_8743);
or U13427 (N_13427,N_6264,N_8072);
or U13428 (N_13428,N_9042,N_7673);
and U13429 (N_13429,N_6266,N_6984);
nand U13430 (N_13430,N_8056,N_9357);
nor U13431 (N_13431,N_8166,N_6852);
and U13432 (N_13432,N_6508,N_8037);
xnor U13433 (N_13433,N_6340,N_9091);
xnor U13434 (N_13434,N_5781,N_8585);
nand U13435 (N_13435,N_9321,N_7304);
nand U13436 (N_13436,N_6776,N_6332);
nand U13437 (N_13437,N_5606,N_8486);
nand U13438 (N_13438,N_9874,N_8511);
or U13439 (N_13439,N_5646,N_9530);
nand U13440 (N_13440,N_6388,N_6473);
nand U13441 (N_13441,N_9152,N_7069);
nor U13442 (N_13442,N_7768,N_6902);
xnor U13443 (N_13443,N_5933,N_5140);
and U13444 (N_13444,N_8880,N_7065);
nand U13445 (N_13445,N_5132,N_8894);
nor U13446 (N_13446,N_8192,N_5953);
or U13447 (N_13447,N_5141,N_8426);
or U13448 (N_13448,N_8753,N_6223);
nand U13449 (N_13449,N_6406,N_5675);
or U13450 (N_13450,N_7691,N_8906);
nor U13451 (N_13451,N_9701,N_5670);
xor U13452 (N_13452,N_7247,N_5378);
or U13453 (N_13453,N_5811,N_6005);
and U13454 (N_13454,N_6996,N_7841);
nand U13455 (N_13455,N_6780,N_5543);
and U13456 (N_13456,N_6725,N_6991);
and U13457 (N_13457,N_8808,N_6466);
xnor U13458 (N_13458,N_7275,N_7972);
and U13459 (N_13459,N_5344,N_7772);
nor U13460 (N_13460,N_5075,N_7186);
nor U13461 (N_13461,N_6622,N_8049);
nor U13462 (N_13462,N_7537,N_9494);
and U13463 (N_13463,N_9482,N_8923);
and U13464 (N_13464,N_5963,N_5603);
and U13465 (N_13465,N_9060,N_8328);
nand U13466 (N_13466,N_8015,N_5207);
nand U13467 (N_13467,N_5189,N_5967);
nor U13468 (N_13468,N_6249,N_6506);
or U13469 (N_13469,N_9142,N_5869);
or U13470 (N_13470,N_8679,N_5195);
nor U13471 (N_13471,N_5661,N_5236);
nand U13472 (N_13472,N_5597,N_9720);
xor U13473 (N_13473,N_6917,N_8385);
or U13474 (N_13474,N_9887,N_5118);
nor U13475 (N_13475,N_6692,N_8276);
or U13476 (N_13476,N_6281,N_9305);
and U13477 (N_13477,N_5348,N_5709);
and U13478 (N_13478,N_5066,N_7082);
nand U13479 (N_13479,N_5227,N_9453);
or U13480 (N_13480,N_7089,N_7301);
and U13481 (N_13481,N_9406,N_6692);
or U13482 (N_13482,N_7368,N_6473);
nand U13483 (N_13483,N_5550,N_5480);
and U13484 (N_13484,N_6283,N_9137);
or U13485 (N_13485,N_9651,N_8596);
or U13486 (N_13486,N_8367,N_6409);
or U13487 (N_13487,N_8239,N_8625);
nor U13488 (N_13488,N_5068,N_6680);
and U13489 (N_13489,N_5848,N_5685);
and U13490 (N_13490,N_7478,N_7416);
and U13491 (N_13491,N_5326,N_9055);
nor U13492 (N_13492,N_6130,N_8589);
nand U13493 (N_13493,N_7439,N_9046);
and U13494 (N_13494,N_7939,N_7140);
and U13495 (N_13495,N_9135,N_5891);
nor U13496 (N_13496,N_9564,N_9983);
or U13497 (N_13497,N_8613,N_8042);
nand U13498 (N_13498,N_5168,N_9411);
xnor U13499 (N_13499,N_6069,N_7223);
and U13500 (N_13500,N_8598,N_7773);
nand U13501 (N_13501,N_7948,N_9742);
nand U13502 (N_13502,N_8264,N_9680);
nor U13503 (N_13503,N_5043,N_9675);
or U13504 (N_13504,N_5100,N_6161);
or U13505 (N_13505,N_8786,N_9384);
and U13506 (N_13506,N_6738,N_5019);
nor U13507 (N_13507,N_8897,N_7573);
nand U13508 (N_13508,N_7347,N_7171);
xnor U13509 (N_13509,N_9195,N_5447);
nor U13510 (N_13510,N_5396,N_9848);
nor U13511 (N_13511,N_9142,N_6511);
nand U13512 (N_13512,N_6990,N_6858);
nor U13513 (N_13513,N_8445,N_9829);
xor U13514 (N_13514,N_5292,N_6220);
and U13515 (N_13515,N_9838,N_9447);
nand U13516 (N_13516,N_5748,N_7065);
nand U13517 (N_13517,N_6033,N_9871);
or U13518 (N_13518,N_9873,N_5081);
and U13519 (N_13519,N_7811,N_7764);
nand U13520 (N_13520,N_5854,N_7649);
xnor U13521 (N_13521,N_8318,N_7676);
nor U13522 (N_13522,N_8804,N_5130);
xnor U13523 (N_13523,N_5037,N_8272);
or U13524 (N_13524,N_8787,N_8124);
and U13525 (N_13525,N_7115,N_9193);
nor U13526 (N_13526,N_8966,N_9109);
or U13527 (N_13527,N_9908,N_5653);
nor U13528 (N_13528,N_9362,N_9967);
nand U13529 (N_13529,N_8987,N_9910);
and U13530 (N_13530,N_5777,N_7390);
nor U13531 (N_13531,N_9074,N_5341);
nor U13532 (N_13532,N_6123,N_9511);
nor U13533 (N_13533,N_8280,N_6746);
or U13534 (N_13534,N_9503,N_5076);
nand U13535 (N_13535,N_9377,N_5486);
nand U13536 (N_13536,N_5755,N_7756);
nor U13537 (N_13537,N_5318,N_7768);
and U13538 (N_13538,N_7221,N_6508);
nand U13539 (N_13539,N_9730,N_7399);
nor U13540 (N_13540,N_8241,N_7350);
nor U13541 (N_13541,N_8468,N_8015);
or U13542 (N_13542,N_8293,N_7895);
xnor U13543 (N_13543,N_8863,N_9233);
nor U13544 (N_13544,N_8196,N_9903);
and U13545 (N_13545,N_8558,N_6276);
and U13546 (N_13546,N_5021,N_7267);
nand U13547 (N_13547,N_8201,N_5604);
nor U13548 (N_13548,N_7297,N_6794);
and U13549 (N_13549,N_8563,N_7896);
and U13550 (N_13550,N_9397,N_5622);
nand U13551 (N_13551,N_7875,N_9156);
or U13552 (N_13552,N_7649,N_9505);
nor U13553 (N_13553,N_9602,N_5845);
nand U13554 (N_13554,N_7969,N_6303);
and U13555 (N_13555,N_9764,N_6015);
and U13556 (N_13556,N_6643,N_6670);
and U13557 (N_13557,N_9838,N_6404);
xnor U13558 (N_13558,N_6155,N_5431);
and U13559 (N_13559,N_7537,N_6705);
and U13560 (N_13560,N_8492,N_5417);
or U13561 (N_13561,N_7867,N_9003);
xor U13562 (N_13562,N_7078,N_9566);
nand U13563 (N_13563,N_9905,N_9281);
and U13564 (N_13564,N_5790,N_6546);
nand U13565 (N_13565,N_7119,N_5540);
nor U13566 (N_13566,N_5017,N_6234);
and U13567 (N_13567,N_6581,N_9414);
or U13568 (N_13568,N_7835,N_8231);
xor U13569 (N_13569,N_7810,N_6593);
nor U13570 (N_13570,N_6088,N_5529);
and U13571 (N_13571,N_5680,N_7522);
nand U13572 (N_13572,N_7853,N_5831);
and U13573 (N_13573,N_9065,N_7192);
or U13574 (N_13574,N_9589,N_7455);
nand U13575 (N_13575,N_7310,N_6951);
or U13576 (N_13576,N_5540,N_7379);
and U13577 (N_13577,N_6831,N_8548);
and U13578 (N_13578,N_6495,N_7985);
or U13579 (N_13579,N_9069,N_8932);
nand U13580 (N_13580,N_7372,N_8176);
or U13581 (N_13581,N_8344,N_7404);
nand U13582 (N_13582,N_7646,N_7451);
or U13583 (N_13583,N_9766,N_6608);
and U13584 (N_13584,N_6984,N_5077);
or U13585 (N_13585,N_9146,N_9454);
or U13586 (N_13586,N_8151,N_8004);
and U13587 (N_13587,N_6615,N_8575);
nand U13588 (N_13588,N_9256,N_7498);
and U13589 (N_13589,N_5826,N_7596);
xnor U13590 (N_13590,N_9350,N_5970);
and U13591 (N_13591,N_7229,N_9108);
xor U13592 (N_13592,N_8185,N_9594);
nor U13593 (N_13593,N_5406,N_7156);
nor U13594 (N_13594,N_5782,N_5767);
xor U13595 (N_13595,N_6623,N_7828);
or U13596 (N_13596,N_8750,N_7522);
nor U13597 (N_13597,N_8050,N_9399);
nand U13598 (N_13598,N_7156,N_6265);
xnor U13599 (N_13599,N_9893,N_7501);
nand U13600 (N_13600,N_5291,N_6418);
and U13601 (N_13601,N_6670,N_7986);
or U13602 (N_13602,N_7392,N_8952);
nand U13603 (N_13603,N_5157,N_8934);
xnor U13604 (N_13604,N_5873,N_5276);
xnor U13605 (N_13605,N_7463,N_6561);
xnor U13606 (N_13606,N_9973,N_6273);
xnor U13607 (N_13607,N_9180,N_5677);
or U13608 (N_13608,N_8127,N_9246);
nand U13609 (N_13609,N_6333,N_7853);
xnor U13610 (N_13610,N_8192,N_5698);
or U13611 (N_13611,N_7490,N_7702);
nor U13612 (N_13612,N_6374,N_7573);
nand U13613 (N_13613,N_9157,N_6070);
and U13614 (N_13614,N_5335,N_9754);
nand U13615 (N_13615,N_5225,N_6593);
nor U13616 (N_13616,N_6922,N_5846);
and U13617 (N_13617,N_8422,N_7924);
nor U13618 (N_13618,N_5041,N_9327);
nand U13619 (N_13619,N_8968,N_7002);
xnor U13620 (N_13620,N_5718,N_9577);
or U13621 (N_13621,N_6611,N_7433);
nand U13622 (N_13622,N_5536,N_5344);
or U13623 (N_13623,N_7643,N_5584);
or U13624 (N_13624,N_9833,N_6019);
and U13625 (N_13625,N_6942,N_6210);
xor U13626 (N_13626,N_5159,N_6649);
or U13627 (N_13627,N_5108,N_5503);
or U13628 (N_13628,N_6755,N_8347);
xor U13629 (N_13629,N_5283,N_6783);
nand U13630 (N_13630,N_8750,N_8851);
nor U13631 (N_13631,N_9000,N_6310);
nand U13632 (N_13632,N_8574,N_9450);
or U13633 (N_13633,N_7726,N_6696);
and U13634 (N_13634,N_8535,N_7007);
and U13635 (N_13635,N_7570,N_6671);
or U13636 (N_13636,N_7933,N_9315);
or U13637 (N_13637,N_8455,N_5209);
or U13638 (N_13638,N_6415,N_5376);
nand U13639 (N_13639,N_9671,N_8608);
and U13640 (N_13640,N_6347,N_5386);
nor U13641 (N_13641,N_6054,N_6649);
xor U13642 (N_13642,N_7667,N_7230);
and U13643 (N_13643,N_7108,N_7061);
and U13644 (N_13644,N_5652,N_6572);
xor U13645 (N_13645,N_5920,N_9436);
nand U13646 (N_13646,N_6036,N_8043);
nand U13647 (N_13647,N_5917,N_7094);
and U13648 (N_13648,N_6474,N_5217);
and U13649 (N_13649,N_9172,N_5337);
nand U13650 (N_13650,N_6417,N_8689);
nor U13651 (N_13651,N_7804,N_9712);
and U13652 (N_13652,N_9856,N_7005);
xnor U13653 (N_13653,N_6920,N_6612);
nand U13654 (N_13654,N_9952,N_9419);
nor U13655 (N_13655,N_8186,N_9598);
and U13656 (N_13656,N_9969,N_7219);
or U13657 (N_13657,N_8378,N_9135);
nand U13658 (N_13658,N_6775,N_9645);
nand U13659 (N_13659,N_9850,N_8518);
or U13660 (N_13660,N_6323,N_8346);
and U13661 (N_13661,N_5930,N_7831);
and U13662 (N_13662,N_8684,N_9386);
and U13663 (N_13663,N_7604,N_6527);
nand U13664 (N_13664,N_5858,N_9194);
and U13665 (N_13665,N_8498,N_8313);
nand U13666 (N_13666,N_7356,N_5857);
or U13667 (N_13667,N_9755,N_5563);
or U13668 (N_13668,N_9123,N_8725);
and U13669 (N_13669,N_7335,N_6131);
xor U13670 (N_13670,N_8566,N_5187);
nand U13671 (N_13671,N_9381,N_5909);
and U13672 (N_13672,N_9475,N_5417);
nand U13673 (N_13673,N_8670,N_8555);
and U13674 (N_13674,N_8814,N_6733);
nor U13675 (N_13675,N_6080,N_9448);
nor U13676 (N_13676,N_6484,N_5810);
xor U13677 (N_13677,N_7717,N_7020);
nor U13678 (N_13678,N_9277,N_8609);
and U13679 (N_13679,N_9688,N_9807);
nand U13680 (N_13680,N_7958,N_7870);
and U13681 (N_13681,N_5931,N_5334);
or U13682 (N_13682,N_6229,N_9195);
and U13683 (N_13683,N_5911,N_5612);
and U13684 (N_13684,N_8828,N_6753);
and U13685 (N_13685,N_5684,N_8770);
nand U13686 (N_13686,N_6777,N_5370);
nor U13687 (N_13687,N_7270,N_6238);
nand U13688 (N_13688,N_5174,N_8690);
nor U13689 (N_13689,N_7276,N_8367);
and U13690 (N_13690,N_6366,N_5187);
and U13691 (N_13691,N_5958,N_8682);
or U13692 (N_13692,N_9903,N_7089);
nor U13693 (N_13693,N_6652,N_5404);
and U13694 (N_13694,N_9577,N_7814);
and U13695 (N_13695,N_7397,N_7991);
nand U13696 (N_13696,N_8240,N_7784);
nor U13697 (N_13697,N_6691,N_8103);
and U13698 (N_13698,N_8709,N_5027);
or U13699 (N_13699,N_6286,N_6390);
nand U13700 (N_13700,N_7284,N_9838);
and U13701 (N_13701,N_9298,N_8576);
and U13702 (N_13702,N_8997,N_5638);
nor U13703 (N_13703,N_9403,N_8367);
nand U13704 (N_13704,N_7437,N_9063);
or U13705 (N_13705,N_7736,N_8475);
and U13706 (N_13706,N_9238,N_7167);
nand U13707 (N_13707,N_6210,N_8872);
nor U13708 (N_13708,N_7642,N_7353);
nor U13709 (N_13709,N_6338,N_9437);
nand U13710 (N_13710,N_7501,N_7246);
or U13711 (N_13711,N_8798,N_6777);
nand U13712 (N_13712,N_7348,N_7466);
xnor U13713 (N_13713,N_8306,N_8895);
or U13714 (N_13714,N_9225,N_9992);
nor U13715 (N_13715,N_9944,N_5842);
nand U13716 (N_13716,N_9002,N_8135);
nor U13717 (N_13717,N_9595,N_5078);
xnor U13718 (N_13718,N_7436,N_5435);
or U13719 (N_13719,N_5812,N_6845);
xnor U13720 (N_13720,N_9675,N_8563);
or U13721 (N_13721,N_7297,N_6779);
and U13722 (N_13722,N_6267,N_9591);
nor U13723 (N_13723,N_9562,N_7101);
nor U13724 (N_13724,N_8216,N_8361);
nand U13725 (N_13725,N_6823,N_9179);
and U13726 (N_13726,N_5729,N_6504);
xor U13727 (N_13727,N_8908,N_6129);
or U13728 (N_13728,N_6618,N_5903);
nor U13729 (N_13729,N_6290,N_9499);
nand U13730 (N_13730,N_6297,N_9672);
nor U13731 (N_13731,N_8543,N_6590);
nand U13732 (N_13732,N_9444,N_8921);
and U13733 (N_13733,N_6821,N_7778);
nand U13734 (N_13734,N_9341,N_8148);
nand U13735 (N_13735,N_6205,N_6304);
nor U13736 (N_13736,N_9169,N_9942);
or U13737 (N_13737,N_5812,N_6231);
nand U13738 (N_13738,N_8785,N_6135);
nand U13739 (N_13739,N_5945,N_8271);
xnor U13740 (N_13740,N_8893,N_5243);
nor U13741 (N_13741,N_8642,N_8645);
nor U13742 (N_13742,N_5912,N_6761);
or U13743 (N_13743,N_8412,N_9600);
and U13744 (N_13744,N_7874,N_8174);
nand U13745 (N_13745,N_5916,N_7242);
xnor U13746 (N_13746,N_6657,N_5280);
and U13747 (N_13747,N_8732,N_7443);
and U13748 (N_13748,N_9704,N_8648);
nand U13749 (N_13749,N_6877,N_6413);
nand U13750 (N_13750,N_5700,N_9363);
nand U13751 (N_13751,N_6435,N_9342);
and U13752 (N_13752,N_9550,N_7449);
nor U13753 (N_13753,N_9609,N_6918);
nor U13754 (N_13754,N_8960,N_6365);
nand U13755 (N_13755,N_7298,N_6859);
and U13756 (N_13756,N_5103,N_8189);
xnor U13757 (N_13757,N_7625,N_9496);
nor U13758 (N_13758,N_8253,N_9712);
nor U13759 (N_13759,N_8614,N_5914);
nand U13760 (N_13760,N_7492,N_5497);
and U13761 (N_13761,N_5958,N_8681);
nor U13762 (N_13762,N_7990,N_5311);
xor U13763 (N_13763,N_9932,N_7631);
and U13764 (N_13764,N_8034,N_7829);
and U13765 (N_13765,N_9738,N_6735);
nor U13766 (N_13766,N_5721,N_6014);
nor U13767 (N_13767,N_5182,N_6820);
and U13768 (N_13768,N_5656,N_9559);
or U13769 (N_13769,N_6246,N_9470);
nand U13770 (N_13770,N_7366,N_8964);
or U13771 (N_13771,N_5901,N_6942);
nand U13772 (N_13772,N_9122,N_7755);
or U13773 (N_13773,N_5037,N_8472);
nor U13774 (N_13774,N_8040,N_5929);
nand U13775 (N_13775,N_5748,N_8552);
xnor U13776 (N_13776,N_6418,N_8453);
or U13777 (N_13777,N_7889,N_7906);
and U13778 (N_13778,N_7772,N_8953);
and U13779 (N_13779,N_9188,N_8942);
or U13780 (N_13780,N_9984,N_7287);
xnor U13781 (N_13781,N_7710,N_9914);
nor U13782 (N_13782,N_8843,N_7707);
or U13783 (N_13783,N_9567,N_8253);
and U13784 (N_13784,N_7036,N_5907);
nor U13785 (N_13785,N_7046,N_5264);
or U13786 (N_13786,N_5386,N_5884);
nor U13787 (N_13787,N_5173,N_5743);
nand U13788 (N_13788,N_7575,N_6066);
or U13789 (N_13789,N_9135,N_8335);
nand U13790 (N_13790,N_7554,N_8709);
and U13791 (N_13791,N_6652,N_5721);
and U13792 (N_13792,N_9052,N_6886);
and U13793 (N_13793,N_7467,N_5109);
nor U13794 (N_13794,N_9810,N_9633);
or U13795 (N_13795,N_9939,N_6908);
or U13796 (N_13796,N_9994,N_5086);
xnor U13797 (N_13797,N_6804,N_8028);
nor U13798 (N_13798,N_8519,N_6275);
nor U13799 (N_13799,N_6199,N_6901);
nor U13800 (N_13800,N_9132,N_6245);
nor U13801 (N_13801,N_9605,N_5009);
nor U13802 (N_13802,N_8340,N_7147);
nor U13803 (N_13803,N_5551,N_7345);
or U13804 (N_13804,N_6055,N_7970);
and U13805 (N_13805,N_6349,N_9219);
or U13806 (N_13806,N_7476,N_7868);
and U13807 (N_13807,N_6857,N_8101);
or U13808 (N_13808,N_7610,N_8756);
nand U13809 (N_13809,N_6512,N_8461);
nand U13810 (N_13810,N_5971,N_9412);
nand U13811 (N_13811,N_8170,N_5538);
and U13812 (N_13812,N_8727,N_9623);
and U13813 (N_13813,N_9416,N_7973);
or U13814 (N_13814,N_9875,N_5292);
nor U13815 (N_13815,N_6255,N_5346);
or U13816 (N_13816,N_6081,N_5273);
and U13817 (N_13817,N_7794,N_9494);
or U13818 (N_13818,N_8611,N_6764);
nand U13819 (N_13819,N_6720,N_8461);
xor U13820 (N_13820,N_9629,N_5466);
and U13821 (N_13821,N_8017,N_6777);
nand U13822 (N_13822,N_7979,N_7827);
or U13823 (N_13823,N_5471,N_5309);
and U13824 (N_13824,N_7576,N_7743);
nor U13825 (N_13825,N_7258,N_6086);
nand U13826 (N_13826,N_5403,N_7155);
or U13827 (N_13827,N_8586,N_6622);
nor U13828 (N_13828,N_8909,N_6062);
or U13829 (N_13829,N_9802,N_6355);
nor U13830 (N_13830,N_7579,N_9212);
or U13831 (N_13831,N_5215,N_5314);
nor U13832 (N_13832,N_5322,N_7581);
xor U13833 (N_13833,N_9779,N_6788);
and U13834 (N_13834,N_8955,N_8457);
nand U13835 (N_13835,N_5259,N_7844);
or U13836 (N_13836,N_9650,N_9607);
or U13837 (N_13837,N_5618,N_7063);
nand U13838 (N_13838,N_9042,N_7105);
or U13839 (N_13839,N_9397,N_5106);
nor U13840 (N_13840,N_5478,N_6761);
nand U13841 (N_13841,N_5653,N_5161);
nor U13842 (N_13842,N_7399,N_6882);
xor U13843 (N_13843,N_8469,N_7373);
or U13844 (N_13844,N_8711,N_5775);
nand U13845 (N_13845,N_7010,N_9657);
or U13846 (N_13846,N_9810,N_7360);
or U13847 (N_13847,N_8065,N_6345);
or U13848 (N_13848,N_7928,N_6423);
and U13849 (N_13849,N_8205,N_7146);
xnor U13850 (N_13850,N_6799,N_8586);
or U13851 (N_13851,N_9464,N_5148);
and U13852 (N_13852,N_9952,N_6225);
nor U13853 (N_13853,N_5952,N_8639);
nor U13854 (N_13854,N_8351,N_7301);
nand U13855 (N_13855,N_5623,N_5280);
or U13856 (N_13856,N_9260,N_9830);
nand U13857 (N_13857,N_7179,N_9562);
nor U13858 (N_13858,N_9292,N_8203);
and U13859 (N_13859,N_8684,N_7758);
xor U13860 (N_13860,N_7421,N_7034);
and U13861 (N_13861,N_9938,N_6748);
or U13862 (N_13862,N_6656,N_5686);
or U13863 (N_13863,N_5775,N_8918);
nand U13864 (N_13864,N_7152,N_8432);
nand U13865 (N_13865,N_6661,N_6285);
nor U13866 (N_13866,N_5174,N_5688);
and U13867 (N_13867,N_5676,N_9765);
nor U13868 (N_13868,N_9553,N_7543);
nand U13869 (N_13869,N_8009,N_7717);
and U13870 (N_13870,N_9504,N_8179);
or U13871 (N_13871,N_8293,N_7827);
nor U13872 (N_13872,N_7593,N_7943);
xnor U13873 (N_13873,N_7367,N_8949);
or U13874 (N_13874,N_7907,N_9135);
or U13875 (N_13875,N_5163,N_8500);
and U13876 (N_13876,N_8515,N_8722);
xor U13877 (N_13877,N_8539,N_6868);
nand U13878 (N_13878,N_9287,N_6083);
nor U13879 (N_13879,N_8188,N_7238);
nor U13880 (N_13880,N_8419,N_7954);
or U13881 (N_13881,N_5427,N_7056);
or U13882 (N_13882,N_8502,N_9423);
nand U13883 (N_13883,N_7519,N_8624);
nor U13884 (N_13884,N_9930,N_6789);
xor U13885 (N_13885,N_8114,N_6420);
nor U13886 (N_13886,N_8957,N_8709);
and U13887 (N_13887,N_6403,N_9188);
nand U13888 (N_13888,N_8321,N_7784);
or U13889 (N_13889,N_9848,N_9099);
or U13890 (N_13890,N_5736,N_5864);
nor U13891 (N_13891,N_9795,N_8392);
and U13892 (N_13892,N_8237,N_9961);
or U13893 (N_13893,N_5887,N_5668);
or U13894 (N_13894,N_5159,N_6544);
nor U13895 (N_13895,N_8221,N_6979);
xnor U13896 (N_13896,N_7632,N_8084);
nand U13897 (N_13897,N_5369,N_8681);
and U13898 (N_13898,N_7952,N_5923);
nand U13899 (N_13899,N_7706,N_9938);
and U13900 (N_13900,N_5425,N_5265);
nor U13901 (N_13901,N_8298,N_8375);
xor U13902 (N_13902,N_6286,N_6092);
xor U13903 (N_13903,N_6879,N_9833);
and U13904 (N_13904,N_9332,N_7389);
and U13905 (N_13905,N_7157,N_6883);
nor U13906 (N_13906,N_9913,N_8119);
nand U13907 (N_13907,N_8972,N_7776);
nor U13908 (N_13908,N_7989,N_7114);
nand U13909 (N_13909,N_9791,N_5545);
nand U13910 (N_13910,N_8550,N_6631);
and U13911 (N_13911,N_8832,N_5545);
nor U13912 (N_13912,N_7749,N_9804);
nand U13913 (N_13913,N_8139,N_5418);
and U13914 (N_13914,N_7463,N_9677);
nor U13915 (N_13915,N_8148,N_8309);
nor U13916 (N_13916,N_5221,N_5180);
and U13917 (N_13917,N_6675,N_9737);
nand U13918 (N_13918,N_6936,N_9234);
or U13919 (N_13919,N_5629,N_6543);
xnor U13920 (N_13920,N_7351,N_6163);
and U13921 (N_13921,N_8598,N_9350);
or U13922 (N_13922,N_9829,N_5628);
nand U13923 (N_13923,N_6633,N_6555);
or U13924 (N_13924,N_9636,N_8833);
or U13925 (N_13925,N_5505,N_6358);
or U13926 (N_13926,N_7626,N_5774);
and U13927 (N_13927,N_5512,N_7791);
xor U13928 (N_13928,N_9723,N_8837);
nand U13929 (N_13929,N_5764,N_8724);
and U13930 (N_13930,N_8476,N_7559);
nor U13931 (N_13931,N_8297,N_6016);
nand U13932 (N_13932,N_5050,N_5984);
nand U13933 (N_13933,N_6874,N_6083);
and U13934 (N_13934,N_9817,N_9931);
and U13935 (N_13935,N_7667,N_7041);
and U13936 (N_13936,N_9930,N_6798);
nor U13937 (N_13937,N_5581,N_9305);
nor U13938 (N_13938,N_5047,N_9778);
and U13939 (N_13939,N_9684,N_5621);
nor U13940 (N_13940,N_7838,N_7624);
or U13941 (N_13941,N_8304,N_5928);
nand U13942 (N_13942,N_6244,N_8651);
nand U13943 (N_13943,N_8309,N_7519);
and U13944 (N_13944,N_7677,N_6224);
or U13945 (N_13945,N_6339,N_8924);
nand U13946 (N_13946,N_5093,N_8134);
or U13947 (N_13947,N_5530,N_5939);
nor U13948 (N_13948,N_7130,N_6439);
or U13949 (N_13949,N_9225,N_9938);
nand U13950 (N_13950,N_5099,N_7471);
or U13951 (N_13951,N_7490,N_5774);
nor U13952 (N_13952,N_5103,N_8706);
xnor U13953 (N_13953,N_5399,N_9502);
nor U13954 (N_13954,N_8484,N_9036);
nand U13955 (N_13955,N_6158,N_6736);
nor U13956 (N_13956,N_6573,N_7506);
nand U13957 (N_13957,N_5539,N_9205);
or U13958 (N_13958,N_7452,N_8835);
nor U13959 (N_13959,N_8113,N_7220);
nor U13960 (N_13960,N_8794,N_8174);
nor U13961 (N_13961,N_5292,N_5886);
or U13962 (N_13962,N_6556,N_5091);
or U13963 (N_13963,N_7891,N_6267);
nand U13964 (N_13964,N_8344,N_5295);
nand U13965 (N_13965,N_8514,N_8454);
nand U13966 (N_13966,N_5878,N_5136);
xor U13967 (N_13967,N_7856,N_9866);
or U13968 (N_13968,N_9981,N_7224);
nand U13969 (N_13969,N_9501,N_9459);
and U13970 (N_13970,N_9480,N_9885);
nand U13971 (N_13971,N_6625,N_6790);
nor U13972 (N_13972,N_7783,N_7489);
and U13973 (N_13973,N_7438,N_9590);
and U13974 (N_13974,N_6995,N_6683);
or U13975 (N_13975,N_5965,N_7562);
nor U13976 (N_13976,N_7440,N_9184);
and U13977 (N_13977,N_9613,N_7591);
or U13978 (N_13978,N_9501,N_7000);
nand U13979 (N_13979,N_9068,N_8596);
nor U13980 (N_13980,N_5601,N_6228);
nor U13981 (N_13981,N_7357,N_5930);
or U13982 (N_13982,N_8680,N_7730);
or U13983 (N_13983,N_5480,N_9043);
and U13984 (N_13984,N_9756,N_6890);
nor U13985 (N_13985,N_6322,N_8266);
nand U13986 (N_13986,N_8283,N_8296);
or U13987 (N_13987,N_6881,N_6487);
nand U13988 (N_13988,N_5058,N_6397);
or U13989 (N_13989,N_6648,N_6870);
or U13990 (N_13990,N_7257,N_8727);
or U13991 (N_13991,N_5693,N_6712);
nand U13992 (N_13992,N_9777,N_6740);
or U13993 (N_13993,N_8831,N_6573);
nand U13994 (N_13994,N_9790,N_5285);
or U13995 (N_13995,N_5162,N_7476);
and U13996 (N_13996,N_6591,N_6492);
nor U13997 (N_13997,N_6201,N_6654);
and U13998 (N_13998,N_6300,N_7114);
xnor U13999 (N_13999,N_9115,N_6623);
or U14000 (N_14000,N_9715,N_8084);
and U14001 (N_14001,N_6129,N_7100);
nor U14002 (N_14002,N_6589,N_9909);
nor U14003 (N_14003,N_7925,N_8130);
and U14004 (N_14004,N_6704,N_7326);
nand U14005 (N_14005,N_9678,N_9804);
or U14006 (N_14006,N_7252,N_5108);
xnor U14007 (N_14007,N_8428,N_9723);
xnor U14008 (N_14008,N_6503,N_5366);
nor U14009 (N_14009,N_9261,N_6821);
or U14010 (N_14010,N_8115,N_7690);
nor U14011 (N_14011,N_9613,N_8420);
or U14012 (N_14012,N_8363,N_6978);
nor U14013 (N_14013,N_6886,N_7089);
xor U14014 (N_14014,N_6850,N_5743);
and U14015 (N_14015,N_9002,N_6094);
nor U14016 (N_14016,N_8198,N_7729);
nor U14017 (N_14017,N_7088,N_7005);
nor U14018 (N_14018,N_5058,N_9838);
nand U14019 (N_14019,N_7434,N_9015);
xnor U14020 (N_14020,N_9946,N_8475);
xor U14021 (N_14021,N_9359,N_9973);
nor U14022 (N_14022,N_9375,N_6921);
or U14023 (N_14023,N_8118,N_5414);
or U14024 (N_14024,N_8773,N_5058);
nand U14025 (N_14025,N_9831,N_7936);
nand U14026 (N_14026,N_6914,N_7854);
and U14027 (N_14027,N_8505,N_6296);
and U14028 (N_14028,N_8667,N_9383);
nand U14029 (N_14029,N_5558,N_6484);
or U14030 (N_14030,N_8600,N_7430);
xor U14031 (N_14031,N_9514,N_7336);
and U14032 (N_14032,N_8710,N_7983);
nor U14033 (N_14033,N_9130,N_8332);
nand U14034 (N_14034,N_7102,N_8189);
or U14035 (N_14035,N_7365,N_8581);
and U14036 (N_14036,N_9411,N_9166);
xor U14037 (N_14037,N_9439,N_8336);
and U14038 (N_14038,N_9399,N_8597);
and U14039 (N_14039,N_9244,N_6966);
nand U14040 (N_14040,N_8762,N_6171);
or U14041 (N_14041,N_5356,N_7592);
and U14042 (N_14042,N_7617,N_5315);
nor U14043 (N_14043,N_9965,N_6474);
or U14044 (N_14044,N_7908,N_7910);
nor U14045 (N_14045,N_6751,N_6871);
nor U14046 (N_14046,N_7889,N_7204);
xor U14047 (N_14047,N_7791,N_8367);
and U14048 (N_14048,N_7803,N_6379);
or U14049 (N_14049,N_5671,N_7659);
or U14050 (N_14050,N_7518,N_9369);
xnor U14051 (N_14051,N_5749,N_7941);
nor U14052 (N_14052,N_9238,N_6751);
xor U14053 (N_14053,N_5666,N_6619);
and U14054 (N_14054,N_8285,N_6324);
or U14055 (N_14055,N_7995,N_9461);
xnor U14056 (N_14056,N_5385,N_8723);
nand U14057 (N_14057,N_5158,N_7360);
and U14058 (N_14058,N_9036,N_6716);
and U14059 (N_14059,N_7937,N_6717);
xor U14060 (N_14060,N_8141,N_6919);
nand U14061 (N_14061,N_7926,N_7241);
and U14062 (N_14062,N_6641,N_6648);
or U14063 (N_14063,N_9919,N_5762);
nand U14064 (N_14064,N_5272,N_5643);
or U14065 (N_14065,N_6140,N_6014);
nand U14066 (N_14066,N_7016,N_8639);
nand U14067 (N_14067,N_6805,N_5890);
and U14068 (N_14068,N_9694,N_6247);
nor U14069 (N_14069,N_9848,N_5343);
or U14070 (N_14070,N_6623,N_6899);
nand U14071 (N_14071,N_9189,N_7448);
or U14072 (N_14072,N_9117,N_6762);
and U14073 (N_14073,N_7802,N_6722);
and U14074 (N_14074,N_7973,N_6593);
or U14075 (N_14075,N_6124,N_9765);
and U14076 (N_14076,N_5592,N_7311);
xor U14077 (N_14077,N_8637,N_8812);
or U14078 (N_14078,N_7189,N_9647);
or U14079 (N_14079,N_6197,N_7814);
or U14080 (N_14080,N_9731,N_5345);
xnor U14081 (N_14081,N_8910,N_7332);
nor U14082 (N_14082,N_8854,N_5287);
xnor U14083 (N_14083,N_6209,N_6469);
and U14084 (N_14084,N_8379,N_5670);
xnor U14085 (N_14085,N_9453,N_8822);
and U14086 (N_14086,N_6431,N_8079);
xor U14087 (N_14087,N_8693,N_8703);
nand U14088 (N_14088,N_8680,N_6078);
nand U14089 (N_14089,N_5755,N_8910);
or U14090 (N_14090,N_9630,N_8986);
nor U14091 (N_14091,N_8219,N_9025);
xnor U14092 (N_14092,N_5678,N_5042);
or U14093 (N_14093,N_6166,N_9628);
nand U14094 (N_14094,N_7018,N_5786);
nor U14095 (N_14095,N_5097,N_6474);
or U14096 (N_14096,N_5041,N_6867);
and U14097 (N_14097,N_5613,N_8154);
xnor U14098 (N_14098,N_8360,N_9118);
nand U14099 (N_14099,N_6187,N_5429);
nor U14100 (N_14100,N_6079,N_6776);
nor U14101 (N_14101,N_8332,N_9178);
xor U14102 (N_14102,N_8379,N_7179);
xor U14103 (N_14103,N_7751,N_7943);
nor U14104 (N_14104,N_9555,N_6937);
xor U14105 (N_14105,N_5437,N_8841);
nand U14106 (N_14106,N_6014,N_9967);
and U14107 (N_14107,N_5221,N_6775);
nand U14108 (N_14108,N_8460,N_7664);
nor U14109 (N_14109,N_7084,N_5893);
and U14110 (N_14110,N_9842,N_8552);
nand U14111 (N_14111,N_6380,N_6059);
and U14112 (N_14112,N_8579,N_5433);
and U14113 (N_14113,N_6548,N_6492);
nor U14114 (N_14114,N_5308,N_5044);
or U14115 (N_14115,N_7479,N_9052);
xnor U14116 (N_14116,N_8784,N_8262);
or U14117 (N_14117,N_8971,N_9615);
nor U14118 (N_14118,N_6557,N_7042);
nand U14119 (N_14119,N_5045,N_8544);
or U14120 (N_14120,N_6631,N_9418);
nor U14121 (N_14121,N_7027,N_9091);
or U14122 (N_14122,N_7519,N_9402);
or U14123 (N_14123,N_7037,N_7632);
xnor U14124 (N_14124,N_7228,N_7625);
nor U14125 (N_14125,N_8293,N_8721);
or U14126 (N_14126,N_6122,N_5673);
nand U14127 (N_14127,N_6321,N_5638);
and U14128 (N_14128,N_7836,N_9245);
or U14129 (N_14129,N_6408,N_5077);
and U14130 (N_14130,N_7192,N_5736);
xnor U14131 (N_14131,N_8849,N_7809);
nor U14132 (N_14132,N_8676,N_7976);
and U14133 (N_14133,N_8550,N_5417);
nor U14134 (N_14134,N_6655,N_7204);
nand U14135 (N_14135,N_7811,N_8034);
xnor U14136 (N_14136,N_8937,N_5255);
and U14137 (N_14137,N_8312,N_5119);
xor U14138 (N_14138,N_8483,N_8657);
nand U14139 (N_14139,N_5001,N_7964);
nor U14140 (N_14140,N_9890,N_5632);
or U14141 (N_14141,N_5227,N_6800);
nor U14142 (N_14142,N_6249,N_8528);
xnor U14143 (N_14143,N_5606,N_8498);
nand U14144 (N_14144,N_6550,N_7612);
or U14145 (N_14145,N_7808,N_8392);
nor U14146 (N_14146,N_5502,N_8624);
nand U14147 (N_14147,N_6748,N_6103);
and U14148 (N_14148,N_9918,N_7079);
nor U14149 (N_14149,N_5096,N_5498);
nor U14150 (N_14150,N_6389,N_9037);
nand U14151 (N_14151,N_7816,N_5912);
nor U14152 (N_14152,N_7953,N_7369);
nand U14153 (N_14153,N_8911,N_6324);
and U14154 (N_14154,N_6644,N_9368);
and U14155 (N_14155,N_7477,N_7237);
nor U14156 (N_14156,N_9118,N_8825);
nand U14157 (N_14157,N_8133,N_8763);
or U14158 (N_14158,N_8992,N_9987);
and U14159 (N_14159,N_8129,N_8311);
nand U14160 (N_14160,N_8810,N_9049);
or U14161 (N_14161,N_5612,N_7614);
nand U14162 (N_14162,N_5770,N_8994);
or U14163 (N_14163,N_8876,N_6828);
and U14164 (N_14164,N_7495,N_8853);
nor U14165 (N_14165,N_7361,N_6632);
xnor U14166 (N_14166,N_8378,N_9221);
nand U14167 (N_14167,N_8941,N_7753);
nand U14168 (N_14168,N_9864,N_5352);
or U14169 (N_14169,N_5935,N_6933);
nor U14170 (N_14170,N_9948,N_8005);
nand U14171 (N_14171,N_8560,N_8022);
or U14172 (N_14172,N_7720,N_6292);
or U14173 (N_14173,N_5608,N_6421);
nor U14174 (N_14174,N_5887,N_6695);
and U14175 (N_14175,N_7817,N_6765);
or U14176 (N_14176,N_5830,N_7131);
nand U14177 (N_14177,N_8927,N_9213);
nor U14178 (N_14178,N_7106,N_9448);
or U14179 (N_14179,N_9306,N_7669);
or U14180 (N_14180,N_5086,N_8998);
or U14181 (N_14181,N_9427,N_6561);
nor U14182 (N_14182,N_8941,N_5923);
nand U14183 (N_14183,N_5925,N_9201);
or U14184 (N_14184,N_6504,N_5657);
nor U14185 (N_14185,N_8637,N_8463);
or U14186 (N_14186,N_8777,N_5442);
nor U14187 (N_14187,N_9348,N_6971);
or U14188 (N_14188,N_7210,N_9665);
and U14189 (N_14189,N_5601,N_7450);
nand U14190 (N_14190,N_7959,N_8675);
nor U14191 (N_14191,N_8870,N_8584);
or U14192 (N_14192,N_8628,N_6155);
xor U14193 (N_14193,N_6700,N_5297);
xnor U14194 (N_14194,N_5765,N_6013);
and U14195 (N_14195,N_6155,N_9431);
nor U14196 (N_14196,N_6715,N_7197);
and U14197 (N_14197,N_8557,N_7853);
nor U14198 (N_14198,N_9877,N_7202);
or U14199 (N_14199,N_8319,N_9150);
nor U14200 (N_14200,N_6566,N_8466);
nor U14201 (N_14201,N_7479,N_5805);
or U14202 (N_14202,N_8665,N_6633);
or U14203 (N_14203,N_5636,N_9488);
and U14204 (N_14204,N_8743,N_6931);
xnor U14205 (N_14205,N_9355,N_8626);
and U14206 (N_14206,N_9308,N_5535);
and U14207 (N_14207,N_6640,N_6942);
nand U14208 (N_14208,N_5046,N_6988);
or U14209 (N_14209,N_6975,N_5420);
nor U14210 (N_14210,N_6298,N_8495);
and U14211 (N_14211,N_5716,N_6696);
and U14212 (N_14212,N_7085,N_7692);
or U14213 (N_14213,N_8874,N_9702);
nor U14214 (N_14214,N_9799,N_8357);
nor U14215 (N_14215,N_7937,N_9101);
xnor U14216 (N_14216,N_5925,N_9414);
nor U14217 (N_14217,N_5124,N_7925);
nand U14218 (N_14218,N_9675,N_8348);
nand U14219 (N_14219,N_9724,N_8320);
nand U14220 (N_14220,N_7388,N_9723);
or U14221 (N_14221,N_5693,N_6739);
nand U14222 (N_14222,N_5470,N_5580);
nor U14223 (N_14223,N_8952,N_6197);
nand U14224 (N_14224,N_8980,N_5908);
nor U14225 (N_14225,N_8704,N_9061);
nor U14226 (N_14226,N_7370,N_9167);
or U14227 (N_14227,N_5487,N_6887);
nor U14228 (N_14228,N_9494,N_5497);
xor U14229 (N_14229,N_9391,N_9302);
nand U14230 (N_14230,N_8152,N_9105);
and U14231 (N_14231,N_7375,N_9871);
or U14232 (N_14232,N_5364,N_6825);
nand U14233 (N_14233,N_5162,N_6794);
xnor U14234 (N_14234,N_7699,N_6262);
or U14235 (N_14235,N_6622,N_7912);
or U14236 (N_14236,N_8555,N_8200);
nor U14237 (N_14237,N_5246,N_6482);
and U14238 (N_14238,N_7959,N_8873);
nor U14239 (N_14239,N_9354,N_8015);
nand U14240 (N_14240,N_8952,N_9006);
and U14241 (N_14241,N_5065,N_7911);
nand U14242 (N_14242,N_9647,N_6775);
or U14243 (N_14243,N_9960,N_6494);
nor U14244 (N_14244,N_5367,N_8113);
nand U14245 (N_14245,N_8906,N_7002);
and U14246 (N_14246,N_7480,N_7817);
nand U14247 (N_14247,N_6503,N_6470);
nor U14248 (N_14248,N_7852,N_9395);
nand U14249 (N_14249,N_5433,N_9783);
and U14250 (N_14250,N_8083,N_5411);
or U14251 (N_14251,N_5147,N_6280);
nand U14252 (N_14252,N_6827,N_5265);
nand U14253 (N_14253,N_9011,N_9482);
and U14254 (N_14254,N_9493,N_5393);
or U14255 (N_14255,N_5935,N_9996);
and U14256 (N_14256,N_8834,N_9556);
nand U14257 (N_14257,N_9300,N_8357);
nor U14258 (N_14258,N_7341,N_5065);
nor U14259 (N_14259,N_8912,N_5166);
nor U14260 (N_14260,N_9539,N_9949);
nor U14261 (N_14261,N_7262,N_9635);
nand U14262 (N_14262,N_7887,N_8756);
or U14263 (N_14263,N_9063,N_7586);
nor U14264 (N_14264,N_7122,N_7132);
and U14265 (N_14265,N_5024,N_9947);
nand U14266 (N_14266,N_7082,N_9126);
and U14267 (N_14267,N_5933,N_5416);
nor U14268 (N_14268,N_8500,N_9884);
or U14269 (N_14269,N_6966,N_5672);
and U14270 (N_14270,N_8723,N_6448);
and U14271 (N_14271,N_8974,N_9401);
nand U14272 (N_14272,N_7599,N_9464);
nand U14273 (N_14273,N_9936,N_8022);
and U14274 (N_14274,N_8695,N_8940);
or U14275 (N_14275,N_5770,N_6471);
nand U14276 (N_14276,N_5089,N_8195);
nand U14277 (N_14277,N_7114,N_6389);
xor U14278 (N_14278,N_8692,N_7956);
nor U14279 (N_14279,N_8574,N_6794);
or U14280 (N_14280,N_9308,N_6706);
nor U14281 (N_14281,N_7282,N_7888);
and U14282 (N_14282,N_5669,N_8465);
or U14283 (N_14283,N_8273,N_8184);
or U14284 (N_14284,N_7321,N_5232);
nor U14285 (N_14285,N_8260,N_9588);
nand U14286 (N_14286,N_7343,N_8339);
or U14287 (N_14287,N_9218,N_6594);
nand U14288 (N_14288,N_8247,N_8809);
and U14289 (N_14289,N_9240,N_9340);
and U14290 (N_14290,N_6613,N_9911);
or U14291 (N_14291,N_6221,N_8172);
xnor U14292 (N_14292,N_8723,N_8178);
nand U14293 (N_14293,N_5273,N_5288);
or U14294 (N_14294,N_9625,N_7170);
nand U14295 (N_14295,N_7157,N_7989);
or U14296 (N_14296,N_9657,N_6817);
or U14297 (N_14297,N_6160,N_7111);
or U14298 (N_14298,N_9484,N_5293);
and U14299 (N_14299,N_6672,N_7130);
nand U14300 (N_14300,N_9739,N_9875);
or U14301 (N_14301,N_7318,N_5474);
and U14302 (N_14302,N_7203,N_8597);
xnor U14303 (N_14303,N_5598,N_9561);
and U14304 (N_14304,N_5530,N_7179);
and U14305 (N_14305,N_9613,N_5369);
or U14306 (N_14306,N_5053,N_8204);
nor U14307 (N_14307,N_9229,N_5847);
nor U14308 (N_14308,N_7381,N_5809);
and U14309 (N_14309,N_9683,N_9143);
and U14310 (N_14310,N_6514,N_7718);
nand U14311 (N_14311,N_5545,N_5131);
nand U14312 (N_14312,N_8311,N_6134);
xor U14313 (N_14313,N_6635,N_8925);
xor U14314 (N_14314,N_5413,N_6714);
nand U14315 (N_14315,N_8268,N_8575);
xnor U14316 (N_14316,N_5573,N_6975);
nor U14317 (N_14317,N_8550,N_6267);
nand U14318 (N_14318,N_7736,N_7770);
nand U14319 (N_14319,N_9441,N_6289);
nor U14320 (N_14320,N_5823,N_6459);
and U14321 (N_14321,N_7226,N_6297);
xnor U14322 (N_14322,N_7724,N_5030);
nor U14323 (N_14323,N_6463,N_6120);
and U14324 (N_14324,N_8373,N_5514);
and U14325 (N_14325,N_9715,N_6376);
nand U14326 (N_14326,N_6884,N_8447);
and U14327 (N_14327,N_7848,N_7168);
nand U14328 (N_14328,N_6814,N_8238);
and U14329 (N_14329,N_7113,N_6467);
and U14330 (N_14330,N_6530,N_8781);
nor U14331 (N_14331,N_9407,N_8332);
and U14332 (N_14332,N_8800,N_8571);
and U14333 (N_14333,N_6432,N_8831);
xor U14334 (N_14334,N_9101,N_5766);
or U14335 (N_14335,N_9877,N_7455);
and U14336 (N_14336,N_9659,N_5181);
nor U14337 (N_14337,N_7153,N_9281);
nor U14338 (N_14338,N_9503,N_6026);
nand U14339 (N_14339,N_8761,N_6587);
nor U14340 (N_14340,N_7388,N_6357);
nand U14341 (N_14341,N_5245,N_9084);
or U14342 (N_14342,N_9338,N_5875);
nor U14343 (N_14343,N_5587,N_6174);
and U14344 (N_14344,N_6528,N_8022);
or U14345 (N_14345,N_5003,N_9830);
nor U14346 (N_14346,N_6810,N_5628);
or U14347 (N_14347,N_8129,N_9811);
and U14348 (N_14348,N_6033,N_8595);
or U14349 (N_14349,N_8770,N_7984);
nand U14350 (N_14350,N_7639,N_7895);
or U14351 (N_14351,N_8698,N_6852);
nor U14352 (N_14352,N_9071,N_6157);
or U14353 (N_14353,N_9634,N_5153);
nand U14354 (N_14354,N_6099,N_6159);
and U14355 (N_14355,N_8557,N_9162);
nand U14356 (N_14356,N_5969,N_9957);
nor U14357 (N_14357,N_8575,N_5437);
and U14358 (N_14358,N_8656,N_6374);
or U14359 (N_14359,N_6263,N_5788);
or U14360 (N_14360,N_8885,N_6153);
or U14361 (N_14361,N_8120,N_9414);
or U14362 (N_14362,N_8314,N_7669);
nand U14363 (N_14363,N_8862,N_5806);
xnor U14364 (N_14364,N_8835,N_5139);
and U14365 (N_14365,N_9491,N_6824);
nand U14366 (N_14366,N_6805,N_7471);
nor U14367 (N_14367,N_5001,N_7286);
nand U14368 (N_14368,N_8571,N_8869);
or U14369 (N_14369,N_8246,N_6356);
and U14370 (N_14370,N_9527,N_5625);
xnor U14371 (N_14371,N_5566,N_9251);
or U14372 (N_14372,N_7615,N_6426);
nand U14373 (N_14373,N_9598,N_6293);
nand U14374 (N_14374,N_8291,N_9690);
and U14375 (N_14375,N_9310,N_7669);
nor U14376 (N_14376,N_6422,N_9069);
or U14377 (N_14377,N_5693,N_7620);
or U14378 (N_14378,N_8230,N_8825);
nand U14379 (N_14379,N_5849,N_9551);
and U14380 (N_14380,N_7061,N_7185);
nor U14381 (N_14381,N_6846,N_8453);
and U14382 (N_14382,N_6566,N_9201);
nor U14383 (N_14383,N_6773,N_9575);
nand U14384 (N_14384,N_8720,N_6747);
and U14385 (N_14385,N_5923,N_6479);
or U14386 (N_14386,N_5377,N_6842);
xor U14387 (N_14387,N_8492,N_6742);
and U14388 (N_14388,N_8093,N_9739);
nand U14389 (N_14389,N_8782,N_5320);
or U14390 (N_14390,N_7786,N_6030);
xnor U14391 (N_14391,N_8528,N_8421);
nand U14392 (N_14392,N_6085,N_8308);
or U14393 (N_14393,N_5122,N_5824);
nor U14394 (N_14394,N_6553,N_7379);
xor U14395 (N_14395,N_7021,N_8241);
nor U14396 (N_14396,N_9593,N_5764);
nor U14397 (N_14397,N_9190,N_7835);
xor U14398 (N_14398,N_5820,N_6186);
nor U14399 (N_14399,N_5506,N_9310);
or U14400 (N_14400,N_7173,N_5098);
nand U14401 (N_14401,N_9446,N_8546);
or U14402 (N_14402,N_8171,N_6373);
nor U14403 (N_14403,N_9542,N_6134);
nor U14404 (N_14404,N_5174,N_6513);
or U14405 (N_14405,N_9644,N_7783);
nand U14406 (N_14406,N_7668,N_8837);
nor U14407 (N_14407,N_9510,N_9771);
nand U14408 (N_14408,N_7066,N_6680);
nor U14409 (N_14409,N_7636,N_5395);
nand U14410 (N_14410,N_9091,N_7411);
and U14411 (N_14411,N_7581,N_5399);
nand U14412 (N_14412,N_8215,N_8472);
and U14413 (N_14413,N_5297,N_9551);
nor U14414 (N_14414,N_6923,N_8775);
or U14415 (N_14415,N_6155,N_7563);
and U14416 (N_14416,N_6189,N_6004);
and U14417 (N_14417,N_6746,N_7662);
nand U14418 (N_14418,N_5637,N_8637);
and U14419 (N_14419,N_5606,N_7694);
nand U14420 (N_14420,N_9704,N_9490);
nor U14421 (N_14421,N_5075,N_7363);
and U14422 (N_14422,N_9156,N_9976);
nor U14423 (N_14423,N_5324,N_7489);
or U14424 (N_14424,N_8528,N_6839);
and U14425 (N_14425,N_5843,N_9754);
and U14426 (N_14426,N_7167,N_5972);
or U14427 (N_14427,N_9055,N_7232);
nor U14428 (N_14428,N_5458,N_8468);
and U14429 (N_14429,N_5811,N_8762);
and U14430 (N_14430,N_8650,N_6147);
nand U14431 (N_14431,N_6601,N_5042);
xnor U14432 (N_14432,N_9617,N_9538);
or U14433 (N_14433,N_7091,N_5028);
and U14434 (N_14434,N_6790,N_7515);
nand U14435 (N_14435,N_6920,N_7737);
nor U14436 (N_14436,N_5426,N_7332);
nor U14437 (N_14437,N_6875,N_6271);
nor U14438 (N_14438,N_9740,N_8343);
or U14439 (N_14439,N_8107,N_8761);
or U14440 (N_14440,N_8437,N_8017);
or U14441 (N_14441,N_8303,N_9633);
or U14442 (N_14442,N_7519,N_7512);
nor U14443 (N_14443,N_8788,N_7640);
and U14444 (N_14444,N_9488,N_7434);
or U14445 (N_14445,N_6570,N_9255);
and U14446 (N_14446,N_8841,N_6781);
and U14447 (N_14447,N_7076,N_7510);
and U14448 (N_14448,N_5601,N_7111);
and U14449 (N_14449,N_7175,N_9508);
or U14450 (N_14450,N_6018,N_9365);
or U14451 (N_14451,N_6796,N_9379);
or U14452 (N_14452,N_5773,N_7543);
nand U14453 (N_14453,N_8156,N_9829);
and U14454 (N_14454,N_7072,N_7218);
nor U14455 (N_14455,N_9099,N_9653);
or U14456 (N_14456,N_9561,N_7620);
and U14457 (N_14457,N_7079,N_5157);
nor U14458 (N_14458,N_5870,N_5347);
and U14459 (N_14459,N_6808,N_8371);
and U14460 (N_14460,N_6283,N_9416);
nor U14461 (N_14461,N_9861,N_9214);
or U14462 (N_14462,N_9375,N_9633);
nor U14463 (N_14463,N_5221,N_6325);
and U14464 (N_14464,N_7338,N_6774);
nor U14465 (N_14465,N_6466,N_8027);
xnor U14466 (N_14466,N_6373,N_6181);
or U14467 (N_14467,N_5163,N_7289);
nand U14468 (N_14468,N_8809,N_7653);
or U14469 (N_14469,N_9763,N_8328);
and U14470 (N_14470,N_6428,N_9013);
nand U14471 (N_14471,N_6622,N_5058);
nor U14472 (N_14472,N_5665,N_5009);
or U14473 (N_14473,N_9620,N_6300);
nand U14474 (N_14474,N_8571,N_7129);
nand U14475 (N_14475,N_8659,N_7460);
or U14476 (N_14476,N_5857,N_8131);
nand U14477 (N_14477,N_6153,N_9964);
nor U14478 (N_14478,N_5846,N_7540);
and U14479 (N_14479,N_8328,N_8226);
xnor U14480 (N_14480,N_7963,N_5127);
xnor U14481 (N_14481,N_8138,N_7019);
nor U14482 (N_14482,N_9919,N_6968);
nor U14483 (N_14483,N_8380,N_7880);
and U14484 (N_14484,N_7970,N_5879);
xnor U14485 (N_14485,N_5011,N_5983);
and U14486 (N_14486,N_9563,N_9206);
nand U14487 (N_14487,N_7558,N_7541);
or U14488 (N_14488,N_6900,N_8861);
or U14489 (N_14489,N_8244,N_7720);
nand U14490 (N_14490,N_9497,N_6171);
and U14491 (N_14491,N_9325,N_9032);
xor U14492 (N_14492,N_6601,N_8908);
nor U14493 (N_14493,N_9904,N_9373);
nor U14494 (N_14494,N_7507,N_6720);
nor U14495 (N_14495,N_5715,N_9801);
or U14496 (N_14496,N_7790,N_7734);
nand U14497 (N_14497,N_6675,N_7643);
xnor U14498 (N_14498,N_7774,N_6036);
nor U14499 (N_14499,N_8722,N_9175);
and U14500 (N_14500,N_8518,N_9671);
nor U14501 (N_14501,N_8505,N_5962);
nor U14502 (N_14502,N_7968,N_7497);
xnor U14503 (N_14503,N_5988,N_9552);
and U14504 (N_14504,N_6706,N_7026);
nor U14505 (N_14505,N_5070,N_6006);
or U14506 (N_14506,N_6625,N_8514);
xor U14507 (N_14507,N_8711,N_6624);
or U14508 (N_14508,N_8291,N_8992);
xnor U14509 (N_14509,N_9673,N_5326);
or U14510 (N_14510,N_6908,N_6821);
nand U14511 (N_14511,N_9712,N_8397);
nand U14512 (N_14512,N_5050,N_6820);
and U14513 (N_14513,N_8507,N_7722);
nand U14514 (N_14514,N_7387,N_9437);
or U14515 (N_14515,N_7297,N_7388);
nand U14516 (N_14516,N_5213,N_6350);
and U14517 (N_14517,N_7619,N_9771);
xor U14518 (N_14518,N_9553,N_8879);
nand U14519 (N_14519,N_7132,N_6553);
nor U14520 (N_14520,N_7237,N_8467);
or U14521 (N_14521,N_6716,N_8029);
and U14522 (N_14522,N_5293,N_8530);
and U14523 (N_14523,N_9934,N_8218);
or U14524 (N_14524,N_9453,N_9533);
nand U14525 (N_14525,N_6413,N_5922);
nand U14526 (N_14526,N_6351,N_5175);
or U14527 (N_14527,N_7442,N_9125);
xor U14528 (N_14528,N_9588,N_9159);
or U14529 (N_14529,N_9791,N_7797);
xor U14530 (N_14530,N_8594,N_6820);
xnor U14531 (N_14531,N_5819,N_5715);
or U14532 (N_14532,N_8431,N_7361);
nor U14533 (N_14533,N_5536,N_9886);
nor U14534 (N_14534,N_9882,N_5888);
and U14535 (N_14535,N_5659,N_8498);
xor U14536 (N_14536,N_5475,N_7357);
and U14537 (N_14537,N_9667,N_6348);
xnor U14538 (N_14538,N_6938,N_9469);
nor U14539 (N_14539,N_5761,N_9437);
nor U14540 (N_14540,N_7937,N_9635);
nand U14541 (N_14541,N_8903,N_8417);
nor U14542 (N_14542,N_5682,N_9981);
nor U14543 (N_14543,N_8734,N_8483);
nor U14544 (N_14544,N_5897,N_5067);
or U14545 (N_14545,N_8004,N_5574);
and U14546 (N_14546,N_7995,N_8331);
and U14547 (N_14547,N_7823,N_7605);
nand U14548 (N_14548,N_8795,N_6765);
and U14549 (N_14549,N_6848,N_5560);
and U14550 (N_14550,N_6963,N_6774);
and U14551 (N_14551,N_9115,N_8581);
nand U14552 (N_14552,N_8639,N_5125);
and U14553 (N_14553,N_7478,N_7493);
or U14554 (N_14554,N_9689,N_6151);
and U14555 (N_14555,N_8804,N_6405);
or U14556 (N_14556,N_8523,N_9081);
nand U14557 (N_14557,N_7780,N_6772);
nand U14558 (N_14558,N_5176,N_8068);
nand U14559 (N_14559,N_9859,N_8733);
nand U14560 (N_14560,N_9009,N_9970);
nand U14561 (N_14561,N_8745,N_8303);
nand U14562 (N_14562,N_9811,N_8453);
and U14563 (N_14563,N_6295,N_6860);
and U14564 (N_14564,N_9501,N_7544);
and U14565 (N_14565,N_5567,N_6880);
nor U14566 (N_14566,N_9398,N_7136);
or U14567 (N_14567,N_8229,N_9391);
and U14568 (N_14568,N_6334,N_8809);
and U14569 (N_14569,N_6697,N_8728);
nand U14570 (N_14570,N_9119,N_9857);
nand U14571 (N_14571,N_8906,N_8212);
nand U14572 (N_14572,N_6996,N_9088);
and U14573 (N_14573,N_8164,N_6187);
and U14574 (N_14574,N_8186,N_8667);
or U14575 (N_14575,N_9722,N_5479);
nand U14576 (N_14576,N_9766,N_8956);
nor U14577 (N_14577,N_9058,N_8292);
xor U14578 (N_14578,N_9018,N_7707);
nor U14579 (N_14579,N_9417,N_6857);
or U14580 (N_14580,N_9624,N_8876);
nand U14581 (N_14581,N_9235,N_8759);
or U14582 (N_14582,N_9319,N_6117);
nor U14583 (N_14583,N_5805,N_6337);
or U14584 (N_14584,N_9743,N_8329);
nand U14585 (N_14585,N_8845,N_6897);
nand U14586 (N_14586,N_6686,N_5539);
xor U14587 (N_14587,N_5928,N_8419);
nand U14588 (N_14588,N_9946,N_9071);
and U14589 (N_14589,N_7582,N_5051);
xnor U14590 (N_14590,N_8145,N_7842);
or U14591 (N_14591,N_8387,N_5063);
or U14592 (N_14592,N_8318,N_5279);
nor U14593 (N_14593,N_6090,N_9475);
nand U14594 (N_14594,N_5281,N_5392);
or U14595 (N_14595,N_9607,N_5277);
xnor U14596 (N_14596,N_8225,N_7578);
nand U14597 (N_14597,N_8457,N_7481);
nor U14598 (N_14598,N_9640,N_8773);
or U14599 (N_14599,N_5268,N_8017);
xor U14600 (N_14600,N_7210,N_6448);
nor U14601 (N_14601,N_6547,N_5084);
nand U14602 (N_14602,N_6514,N_8469);
or U14603 (N_14603,N_5073,N_8296);
nor U14604 (N_14604,N_5144,N_7767);
nor U14605 (N_14605,N_5728,N_5701);
xor U14606 (N_14606,N_6876,N_6262);
nand U14607 (N_14607,N_7462,N_9639);
nand U14608 (N_14608,N_5882,N_8477);
nand U14609 (N_14609,N_9712,N_5181);
nor U14610 (N_14610,N_5565,N_5826);
nor U14611 (N_14611,N_9278,N_5891);
or U14612 (N_14612,N_9088,N_7407);
nand U14613 (N_14613,N_9070,N_5232);
xor U14614 (N_14614,N_5171,N_7969);
or U14615 (N_14615,N_9007,N_9878);
nor U14616 (N_14616,N_6657,N_7627);
xnor U14617 (N_14617,N_5871,N_5389);
nor U14618 (N_14618,N_8757,N_8187);
or U14619 (N_14619,N_5756,N_7637);
and U14620 (N_14620,N_5723,N_6452);
and U14621 (N_14621,N_9154,N_5007);
nor U14622 (N_14622,N_9048,N_8411);
or U14623 (N_14623,N_7335,N_9677);
nor U14624 (N_14624,N_8613,N_5322);
nand U14625 (N_14625,N_8771,N_6726);
xnor U14626 (N_14626,N_7825,N_9963);
and U14627 (N_14627,N_6610,N_7578);
and U14628 (N_14628,N_8923,N_9324);
and U14629 (N_14629,N_7597,N_8901);
and U14630 (N_14630,N_8656,N_5842);
or U14631 (N_14631,N_7520,N_9973);
or U14632 (N_14632,N_7988,N_5439);
or U14633 (N_14633,N_6871,N_5521);
or U14634 (N_14634,N_8195,N_8342);
or U14635 (N_14635,N_6607,N_9211);
and U14636 (N_14636,N_7932,N_9420);
xnor U14637 (N_14637,N_6692,N_7097);
or U14638 (N_14638,N_6733,N_8709);
nor U14639 (N_14639,N_8870,N_9127);
nand U14640 (N_14640,N_6254,N_9249);
nor U14641 (N_14641,N_5367,N_5114);
and U14642 (N_14642,N_5920,N_7044);
and U14643 (N_14643,N_5303,N_7481);
or U14644 (N_14644,N_5143,N_6715);
nor U14645 (N_14645,N_6938,N_8866);
nor U14646 (N_14646,N_7682,N_5389);
and U14647 (N_14647,N_5153,N_5836);
or U14648 (N_14648,N_8774,N_7395);
and U14649 (N_14649,N_6686,N_8901);
or U14650 (N_14650,N_9993,N_7970);
xor U14651 (N_14651,N_7652,N_8232);
and U14652 (N_14652,N_8198,N_6224);
and U14653 (N_14653,N_7601,N_6958);
nor U14654 (N_14654,N_7041,N_5853);
nand U14655 (N_14655,N_5094,N_9883);
xor U14656 (N_14656,N_5927,N_9801);
or U14657 (N_14657,N_5649,N_9015);
xnor U14658 (N_14658,N_5624,N_9738);
xor U14659 (N_14659,N_5327,N_9276);
nor U14660 (N_14660,N_8110,N_8477);
nor U14661 (N_14661,N_5301,N_6275);
or U14662 (N_14662,N_8289,N_7365);
xor U14663 (N_14663,N_8814,N_9405);
or U14664 (N_14664,N_5872,N_6262);
nor U14665 (N_14665,N_5094,N_5653);
xor U14666 (N_14666,N_9592,N_6341);
nand U14667 (N_14667,N_8935,N_9793);
nand U14668 (N_14668,N_7899,N_9079);
xnor U14669 (N_14669,N_5024,N_8362);
nor U14670 (N_14670,N_9297,N_7315);
nand U14671 (N_14671,N_8136,N_5212);
or U14672 (N_14672,N_6661,N_5060);
and U14673 (N_14673,N_8227,N_5625);
nand U14674 (N_14674,N_9244,N_5096);
nand U14675 (N_14675,N_9522,N_5734);
xnor U14676 (N_14676,N_6897,N_9579);
nand U14677 (N_14677,N_7719,N_5263);
nor U14678 (N_14678,N_8451,N_6509);
and U14679 (N_14679,N_7220,N_7184);
nor U14680 (N_14680,N_7823,N_8835);
nand U14681 (N_14681,N_6676,N_8370);
nand U14682 (N_14682,N_5552,N_6060);
nor U14683 (N_14683,N_7563,N_5025);
nor U14684 (N_14684,N_7612,N_5677);
and U14685 (N_14685,N_7442,N_8373);
xnor U14686 (N_14686,N_5684,N_8718);
or U14687 (N_14687,N_6271,N_5132);
nand U14688 (N_14688,N_7202,N_9048);
nor U14689 (N_14689,N_5729,N_9768);
xor U14690 (N_14690,N_8068,N_6367);
and U14691 (N_14691,N_9765,N_8066);
xnor U14692 (N_14692,N_9596,N_6055);
xnor U14693 (N_14693,N_5268,N_5045);
nor U14694 (N_14694,N_8180,N_7251);
and U14695 (N_14695,N_7210,N_5991);
nor U14696 (N_14696,N_9935,N_7983);
or U14697 (N_14697,N_5112,N_8955);
nor U14698 (N_14698,N_5979,N_8871);
nor U14699 (N_14699,N_5364,N_7063);
or U14700 (N_14700,N_8243,N_8635);
nand U14701 (N_14701,N_5257,N_6265);
and U14702 (N_14702,N_6616,N_7507);
and U14703 (N_14703,N_6155,N_7912);
and U14704 (N_14704,N_5780,N_7743);
or U14705 (N_14705,N_9089,N_9193);
nor U14706 (N_14706,N_6186,N_9124);
nor U14707 (N_14707,N_6406,N_5422);
nor U14708 (N_14708,N_6982,N_6083);
or U14709 (N_14709,N_9217,N_8699);
xor U14710 (N_14710,N_7870,N_7026);
and U14711 (N_14711,N_7718,N_6731);
nand U14712 (N_14712,N_7468,N_6937);
nand U14713 (N_14713,N_8428,N_5798);
nand U14714 (N_14714,N_7540,N_6718);
nor U14715 (N_14715,N_5769,N_6023);
nor U14716 (N_14716,N_6551,N_5106);
and U14717 (N_14717,N_7582,N_9766);
nand U14718 (N_14718,N_8033,N_6610);
and U14719 (N_14719,N_7459,N_6395);
nand U14720 (N_14720,N_6827,N_7385);
nand U14721 (N_14721,N_7044,N_7629);
xnor U14722 (N_14722,N_7819,N_5621);
or U14723 (N_14723,N_8929,N_6292);
xor U14724 (N_14724,N_7560,N_6774);
xnor U14725 (N_14725,N_6503,N_5583);
nand U14726 (N_14726,N_7277,N_8319);
and U14727 (N_14727,N_5281,N_9992);
nor U14728 (N_14728,N_6966,N_9951);
and U14729 (N_14729,N_7073,N_8543);
nand U14730 (N_14730,N_6603,N_8191);
nand U14731 (N_14731,N_9265,N_6399);
nand U14732 (N_14732,N_5250,N_8404);
nand U14733 (N_14733,N_6145,N_8002);
xor U14734 (N_14734,N_5102,N_9733);
or U14735 (N_14735,N_7590,N_8782);
and U14736 (N_14736,N_6865,N_8624);
nor U14737 (N_14737,N_6881,N_9147);
nor U14738 (N_14738,N_9776,N_5828);
nor U14739 (N_14739,N_9315,N_5664);
or U14740 (N_14740,N_6425,N_9037);
nand U14741 (N_14741,N_9653,N_8694);
and U14742 (N_14742,N_7702,N_9011);
or U14743 (N_14743,N_7742,N_7313);
nor U14744 (N_14744,N_5748,N_9755);
nor U14745 (N_14745,N_8837,N_8718);
or U14746 (N_14746,N_6479,N_9861);
and U14747 (N_14747,N_9942,N_6387);
or U14748 (N_14748,N_5183,N_6653);
nor U14749 (N_14749,N_8363,N_9766);
or U14750 (N_14750,N_6884,N_5410);
or U14751 (N_14751,N_8566,N_8021);
or U14752 (N_14752,N_8483,N_9724);
xnor U14753 (N_14753,N_5922,N_9903);
nand U14754 (N_14754,N_7711,N_8948);
or U14755 (N_14755,N_5440,N_7231);
nor U14756 (N_14756,N_8484,N_9597);
xnor U14757 (N_14757,N_8001,N_8800);
nor U14758 (N_14758,N_5493,N_5405);
and U14759 (N_14759,N_9090,N_9274);
and U14760 (N_14760,N_5749,N_5383);
nor U14761 (N_14761,N_5755,N_8795);
and U14762 (N_14762,N_7963,N_5861);
nor U14763 (N_14763,N_6500,N_7631);
and U14764 (N_14764,N_5401,N_5291);
and U14765 (N_14765,N_9445,N_5926);
nor U14766 (N_14766,N_9674,N_8359);
nor U14767 (N_14767,N_8439,N_7163);
or U14768 (N_14768,N_7637,N_5090);
nor U14769 (N_14769,N_9159,N_7068);
xor U14770 (N_14770,N_8401,N_7187);
nor U14771 (N_14771,N_9828,N_6437);
nand U14772 (N_14772,N_7902,N_7088);
nor U14773 (N_14773,N_7736,N_7675);
xnor U14774 (N_14774,N_8210,N_5551);
and U14775 (N_14775,N_6344,N_5965);
nor U14776 (N_14776,N_8259,N_6654);
and U14777 (N_14777,N_8494,N_9215);
nand U14778 (N_14778,N_7070,N_8521);
or U14779 (N_14779,N_7029,N_6563);
nor U14780 (N_14780,N_8332,N_9330);
and U14781 (N_14781,N_8881,N_6440);
and U14782 (N_14782,N_7535,N_9446);
xnor U14783 (N_14783,N_6957,N_7462);
and U14784 (N_14784,N_7380,N_7203);
and U14785 (N_14785,N_8733,N_8392);
nor U14786 (N_14786,N_5059,N_6773);
nor U14787 (N_14787,N_5980,N_8079);
or U14788 (N_14788,N_9114,N_9159);
or U14789 (N_14789,N_9443,N_9163);
or U14790 (N_14790,N_5843,N_6947);
and U14791 (N_14791,N_8065,N_8214);
nor U14792 (N_14792,N_6281,N_5633);
or U14793 (N_14793,N_9677,N_6399);
nand U14794 (N_14794,N_6325,N_9192);
or U14795 (N_14795,N_7538,N_9869);
and U14796 (N_14796,N_9583,N_5374);
nand U14797 (N_14797,N_5540,N_7476);
nand U14798 (N_14798,N_7499,N_9415);
nand U14799 (N_14799,N_6895,N_8289);
nand U14800 (N_14800,N_7749,N_6360);
xor U14801 (N_14801,N_6850,N_6613);
and U14802 (N_14802,N_9731,N_5404);
xnor U14803 (N_14803,N_5364,N_7952);
and U14804 (N_14804,N_7593,N_7273);
or U14805 (N_14805,N_9339,N_8464);
or U14806 (N_14806,N_9567,N_7649);
and U14807 (N_14807,N_8604,N_9629);
nand U14808 (N_14808,N_8812,N_7084);
nor U14809 (N_14809,N_5952,N_5624);
nor U14810 (N_14810,N_5102,N_9412);
or U14811 (N_14811,N_9411,N_5333);
nand U14812 (N_14812,N_5610,N_8822);
nor U14813 (N_14813,N_8907,N_5214);
or U14814 (N_14814,N_6606,N_5863);
nand U14815 (N_14815,N_8485,N_8637);
or U14816 (N_14816,N_8738,N_6129);
or U14817 (N_14817,N_8679,N_9076);
or U14818 (N_14818,N_7363,N_8688);
or U14819 (N_14819,N_7225,N_8426);
or U14820 (N_14820,N_9172,N_5902);
and U14821 (N_14821,N_8171,N_8709);
xnor U14822 (N_14822,N_7357,N_9231);
and U14823 (N_14823,N_9291,N_6456);
and U14824 (N_14824,N_9753,N_5000);
nand U14825 (N_14825,N_8606,N_9067);
or U14826 (N_14826,N_9488,N_6749);
xnor U14827 (N_14827,N_7933,N_6991);
nand U14828 (N_14828,N_7752,N_5219);
nand U14829 (N_14829,N_5641,N_7919);
nand U14830 (N_14830,N_8083,N_5714);
xor U14831 (N_14831,N_7387,N_7974);
nor U14832 (N_14832,N_6931,N_7309);
nand U14833 (N_14833,N_9837,N_5146);
or U14834 (N_14834,N_9645,N_7760);
and U14835 (N_14835,N_5751,N_5187);
and U14836 (N_14836,N_9471,N_8783);
or U14837 (N_14837,N_6154,N_5928);
nand U14838 (N_14838,N_9338,N_7728);
and U14839 (N_14839,N_8423,N_8757);
and U14840 (N_14840,N_5626,N_8285);
or U14841 (N_14841,N_8149,N_8284);
or U14842 (N_14842,N_5561,N_9172);
nor U14843 (N_14843,N_7006,N_6016);
and U14844 (N_14844,N_7996,N_5367);
nor U14845 (N_14845,N_7948,N_8057);
or U14846 (N_14846,N_7428,N_6084);
nand U14847 (N_14847,N_7626,N_6385);
nand U14848 (N_14848,N_7164,N_7299);
xor U14849 (N_14849,N_9714,N_6207);
or U14850 (N_14850,N_9553,N_8559);
xnor U14851 (N_14851,N_7093,N_8244);
and U14852 (N_14852,N_5488,N_6832);
or U14853 (N_14853,N_8519,N_9262);
nor U14854 (N_14854,N_9394,N_6586);
or U14855 (N_14855,N_5189,N_8898);
xor U14856 (N_14856,N_9929,N_6585);
nand U14857 (N_14857,N_7279,N_5479);
nand U14858 (N_14858,N_8750,N_5894);
nand U14859 (N_14859,N_9987,N_6623);
or U14860 (N_14860,N_5953,N_8744);
or U14861 (N_14861,N_6735,N_9991);
or U14862 (N_14862,N_5268,N_6830);
and U14863 (N_14863,N_6762,N_9589);
or U14864 (N_14864,N_8820,N_9786);
nand U14865 (N_14865,N_9135,N_6157);
nand U14866 (N_14866,N_6285,N_8676);
and U14867 (N_14867,N_7895,N_7968);
or U14868 (N_14868,N_8844,N_6750);
and U14869 (N_14869,N_8336,N_9623);
and U14870 (N_14870,N_5569,N_9165);
xnor U14871 (N_14871,N_7315,N_7577);
and U14872 (N_14872,N_8644,N_8426);
nor U14873 (N_14873,N_5626,N_7781);
nor U14874 (N_14874,N_5535,N_7130);
and U14875 (N_14875,N_5050,N_6195);
and U14876 (N_14876,N_9064,N_6282);
nand U14877 (N_14877,N_6256,N_5474);
nand U14878 (N_14878,N_8311,N_7452);
nand U14879 (N_14879,N_9649,N_6980);
nor U14880 (N_14880,N_5426,N_9969);
and U14881 (N_14881,N_5930,N_7851);
and U14882 (N_14882,N_5703,N_7185);
nor U14883 (N_14883,N_8170,N_8196);
nand U14884 (N_14884,N_9705,N_7886);
or U14885 (N_14885,N_9974,N_7192);
nand U14886 (N_14886,N_7103,N_9086);
or U14887 (N_14887,N_7288,N_5451);
nor U14888 (N_14888,N_9884,N_6201);
and U14889 (N_14889,N_5947,N_8256);
nor U14890 (N_14890,N_8013,N_7810);
nand U14891 (N_14891,N_9361,N_7038);
xor U14892 (N_14892,N_5140,N_5962);
nor U14893 (N_14893,N_9816,N_8476);
and U14894 (N_14894,N_9937,N_8264);
nor U14895 (N_14895,N_7766,N_8941);
nand U14896 (N_14896,N_7553,N_9464);
and U14897 (N_14897,N_9302,N_5766);
xor U14898 (N_14898,N_6287,N_5878);
and U14899 (N_14899,N_5336,N_5474);
nor U14900 (N_14900,N_7492,N_5424);
xor U14901 (N_14901,N_5584,N_5451);
nor U14902 (N_14902,N_5884,N_8493);
nand U14903 (N_14903,N_9501,N_5823);
and U14904 (N_14904,N_5323,N_7686);
xnor U14905 (N_14905,N_5694,N_8120);
or U14906 (N_14906,N_6527,N_8557);
or U14907 (N_14907,N_9072,N_8708);
nor U14908 (N_14908,N_6437,N_6357);
nor U14909 (N_14909,N_7816,N_7602);
nand U14910 (N_14910,N_6036,N_9079);
and U14911 (N_14911,N_6136,N_6913);
nor U14912 (N_14912,N_5053,N_5677);
or U14913 (N_14913,N_6606,N_5496);
and U14914 (N_14914,N_7912,N_6859);
or U14915 (N_14915,N_7926,N_5074);
and U14916 (N_14916,N_7488,N_7356);
or U14917 (N_14917,N_8104,N_9411);
and U14918 (N_14918,N_6756,N_6677);
or U14919 (N_14919,N_9217,N_7306);
nor U14920 (N_14920,N_8246,N_7171);
nand U14921 (N_14921,N_9338,N_9429);
xor U14922 (N_14922,N_9139,N_8545);
xor U14923 (N_14923,N_7423,N_9101);
and U14924 (N_14924,N_6878,N_9986);
and U14925 (N_14925,N_8913,N_7750);
or U14926 (N_14926,N_7361,N_9082);
or U14927 (N_14927,N_5254,N_6316);
xnor U14928 (N_14928,N_6210,N_5127);
nor U14929 (N_14929,N_6869,N_8795);
or U14930 (N_14930,N_8598,N_7905);
xnor U14931 (N_14931,N_8144,N_6435);
nor U14932 (N_14932,N_5934,N_8175);
nand U14933 (N_14933,N_6980,N_9044);
or U14934 (N_14934,N_8113,N_7941);
or U14935 (N_14935,N_8255,N_9070);
or U14936 (N_14936,N_8763,N_7045);
nor U14937 (N_14937,N_6721,N_6333);
nor U14938 (N_14938,N_8488,N_5791);
and U14939 (N_14939,N_9411,N_9031);
xnor U14940 (N_14940,N_7637,N_6065);
xnor U14941 (N_14941,N_6010,N_8630);
and U14942 (N_14942,N_5385,N_6303);
xor U14943 (N_14943,N_8130,N_9788);
nor U14944 (N_14944,N_8442,N_8683);
and U14945 (N_14945,N_6305,N_5542);
and U14946 (N_14946,N_5684,N_5749);
nand U14947 (N_14947,N_9141,N_9579);
nor U14948 (N_14948,N_9914,N_5033);
and U14949 (N_14949,N_7506,N_7988);
nor U14950 (N_14950,N_5088,N_9862);
or U14951 (N_14951,N_7683,N_6857);
or U14952 (N_14952,N_8709,N_6708);
or U14953 (N_14953,N_5681,N_6365);
or U14954 (N_14954,N_6361,N_6981);
and U14955 (N_14955,N_6230,N_8131);
and U14956 (N_14956,N_6894,N_9732);
nand U14957 (N_14957,N_8215,N_7661);
and U14958 (N_14958,N_6373,N_7666);
nor U14959 (N_14959,N_6358,N_5037);
nor U14960 (N_14960,N_6058,N_7655);
nor U14961 (N_14961,N_9639,N_7543);
or U14962 (N_14962,N_6671,N_5999);
or U14963 (N_14963,N_6506,N_9725);
nor U14964 (N_14964,N_5587,N_5494);
nor U14965 (N_14965,N_8218,N_8255);
nand U14966 (N_14966,N_8065,N_9395);
nand U14967 (N_14967,N_7786,N_5435);
or U14968 (N_14968,N_9953,N_8185);
and U14969 (N_14969,N_6801,N_5970);
or U14970 (N_14970,N_5063,N_7240);
xor U14971 (N_14971,N_5356,N_5078);
and U14972 (N_14972,N_8572,N_7914);
and U14973 (N_14973,N_7121,N_5304);
or U14974 (N_14974,N_5992,N_8959);
and U14975 (N_14975,N_8323,N_8694);
nand U14976 (N_14976,N_6397,N_5390);
nor U14977 (N_14977,N_9784,N_7993);
xor U14978 (N_14978,N_7072,N_8941);
and U14979 (N_14979,N_7889,N_7976);
nor U14980 (N_14980,N_6887,N_9691);
and U14981 (N_14981,N_6304,N_9052);
nand U14982 (N_14982,N_5484,N_6342);
and U14983 (N_14983,N_7142,N_5854);
and U14984 (N_14984,N_5817,N_9159);
xnor U14985 (N_14985,N_7706,N_9175);
nand U14986 (N_14986,N_6476,N_8882);
nand U14987 (N_14987,N_9810,N_9911);
or U14988 (N_14988,N_7776,N_9492);
nor U14989 (N_14989,N_6317,N_5900);
xnor U14990 (N_14990,N_7431,N_5425);
and U14991 (N_14991,N_7003,N_8916);
nor U14992 (N_14992,N_8098,N_7333);
nor U14993 (N_14993,N_6962,N_8492);
xnor U14994 (N_14994,N_9433,N_9029);
or U14995 (N_14995,N_6362,N_6700);
xnor U14996 (N_14996,N_7956,N_5889);
and U14997 (N_14997,N_5080,N_5806);
nand U14998 (N_14998,N_8101,N_5050);
and U14999 (N_14999,N_8900,N_8198);
nand U15000 (N_15000,N_14963,N_11235);
nand U15001 (N_15001,N_12880,N_13668);
or U15002 (N_15002,N_11613,N_14786);
and U15003 (N_15003,N_11776,N_12430);
nand U15004 (N_15004,N_13949,N_10582);
and U15005 (N_15005,N_10803,N_11171);
and U15006 (N_15006,N_14376,N_14273);
nor U15007 (N_15007,N_13682,N_12686);
and U15008 (N_15008,N_12107,N_11579);
xnor U15009 (N_15009,N_13223,N_12033);
and U15010 (N_15010,N_12230,N_10387);
or U15011 (N_15011,N_11580,N_11395);
or U15012 (N_15012,N_12283,N_10594);
nand U15013 (N_15013,N_10519,N_12339);
nor U15014 (N_15014,N_12372,N_11017);
and U15015 (N_15015,N_10413,N_10913);
xnor U15016 (N_15016,N_11011,N_14325);
nand U15017 (N_15017,N_11994,N_10540);
nor U15018 (N_15018,N_14600,N_11967);
nand U15019 (N_15019,N_12597,N_10742);
and U15020 (N_15020,N_11899,N_10168);
nor U15021 (N_15021,N_13732,N_14167);
or U15022 (N_15022,N_11115,N_10672);
and U15023 (N_15023,N_14380,N_13192);
nand U15024 (N_15024,N_14636,N_14206);
or U15025 (N_15025,N_11114,N_14406);
nor U15026 (N_15026,N_10897,N_14005);
or U15027 (N_15027,N_12215,N_14491);
nor U15028 (N_15028,N_11005,N_10308);
and U15029 (N_15029,N_13888,N_13032);
nor U15030 (N_15030,N_14441,N_10202);
xor U15031 (N_15031,N_12444,N_10025);
nor U15032 (N_15032,N_10376,N_13391);
xnor U15033 (N_15033,N_14387,N_12598);
nor U15034 (N_15034,N_11667,N_10045);
or U15035 (N_15035,N_10883,N_10736);
nor U15036 (N_15036,N_12236,N_14945);
or U15037 (N_15037,N_11687,N_14829);
nand U15038 (N_15038,N_11990,N_12287);
or U15039 (N_15039,N_13859,N_14013);
and U15040 (N_15040,N_12785,N_11020);
nand U15041 (N_15041,N_14552,N_10088);
and U15042 (N_15042,N_13741,N_10920);
or U15043 (N_15043,N_12987,N_13801);
nor U15044 (N_15044,N_11264,N_12140);
nand U15045 (N_15045,N_11311,N_12949);
and U15046 (N_15046,N_11714,N_12012);
and U15047 (N_15047,N_13768,N_12040);
and U15048 (N_15048,N_12886,N_12151);
xor U15049 (N_15049,N_14088,N_14578);
or U15050 (N_15050,N_10942,N_13739);
and U15051 (N_15051,N_12931,N_13012);
or U15052 (N_15052,N_11462,N_11051);
and U15053 (N_15053,N_13471,N_13658);
nand U15054 (N_15054,N_12836,N_13092);
nand U15055 (N_15055,N_14535,N_10411);
and U15056 (N_15056,N_10801,N_13652);
nand U15057 (N_15057,N_12994,N_14256);
nor U15058 (N_15058,N_10463,N_14310);
nor U15059 (N_15059,N_14052,N_10646);
or U15060 (N_15060,N_10676,N_13514);
nor U15061 (N_15061,N_14550,N_10812);
and U15062 (N_15062,N_12270,N_10490);
xor U15063 (N_15063,N_14344,N_12299);
xor U15064 (N_15064,N_14332,N_10944);
nor U15065 (N_15065,N_11417,N_12326);
or U15066 (N_15066,N_12711,N_14936);
and U15067 (N_15067,N_13592,N_12835);
nor U15068 (N_15068,N_13114,N_14754);
and U15069 (N_15069,N_10633,N_11228);
and U15070 (N_15070,N_13078,N_12629);
nand U15071 (N_15071,N_12014,N_12344);
or U15072 (N_15072,N_12684,N_11841);
and U15073 (N_15073,N_13014,N_14248);
and U15074 (N_15074,N_14937,N_11009);
and U15075 (N_15075,N_11262,N_11980);
nor U15076 (N_15076,N_13762,N_11824);
and U15077 (N_15077,N_14008,N_11645);
and U15078 (N_15078,N_13957,N_14860);
nand U15079 (N_15079,N_13438,N_12352);
and U15080 (N_15080,N_14217,N_11291);
and U15081 (N_15081,N_13774,N_13319);
or U15082 (N_15082,N_10237,N_12761);
nor U15083 (N_15083,N_12557,N_11304);
and U15084 (N_15084,N_11297,N_13634);
nor U15085 (N_15085,N_14446,N_13182);
and U15086 (N_15086,N_10833,N_13393);
nand U15087 (N_15087,N_10631,N_14927);
or U15088 (N_15088,N_12313,N_12417);
xor U15089 (N_15089,N_10453,N_13996);
nor U15090 (N_15090,N_10969,N_13889);
or U15091 (N_15091,N_10161,N_14382);
nand U15092 (N_15092,N_12055,N_13545);
xor U15093 (N_15093,N_13089,N_10694);
and U15094 (N_15094,N_14479,N_11289);
and U15095 (N_15095,N_11024,N_13353);
nand U15096 (N_15096,N_10776,N_11198);
nor U15097 (N_15097,N_13646,N_13262);
and U15098 (N_15098,N_11674,N_12185);
xnor U15099 (N_15099,N_14843,N_12722);
nand U15100 (N_15100,N_14677,N_11340);
nor U15101 (N_15101,N_14244,N_10125);
nand U15102 (N_15102,N_12022,N_13409);
nor U15103 (N_15103,N_14463,N_14683);
nor U15104 (N_15104,N_14658,N_13776);
nand U15105 (N_15105,N_11438,N_13745);
or U15106 (N_15106,N_10137,N_10034);
nand U15107 (N_15107,N_12092,N_14793);
and U15108 (N_15108,N_14951,N_13523);
and U15109 (N_15109,N_11138,N_10768);
and U15110 (N_15110,N_11661,N_10654);
and U15111 (N_15111,N_10362,N_13168);
nand U15112 (N_15112,N_10759,N_12455);
nand U15113 (N_15113,N_12616,N_10628);
or U15114 (N_15114,N_13371,N_12580);
nor U15115 (N_15115,N_14169,N_14852);
nand U15116 (N_15116,N_13218,N_11883);
and U15117 (N_15117,N_14000,N_10323);
nor U15118 (N_15118,N_14947,N_11528);
nor U15119 (N_15119,N_13659,N_13157);
and U15120 (N_15120,N_10854,N_12291);
or U15121 (N_15121,N_13043,N_10170);
or U15122 (N_15122,N_11632,N_10128);
or U15123 (N_15123,N_12803,N_14823);
and U15124 (N_15124,N_13351,N_11493);
nor U15125 (N_15125,N_10689,N_12190);
nor U15126 (N_15126,N_11895,N_13664);
or U15127 (N_15127,N_13992,N_14520);
or U15128 (N_15128,N_14121,N_14242);
nor U15129 (N_15129,N_10139,N_13425);
and U15130 (N_15130,N_10896,N_13788);
and U15131 (N_15131,N_14370,N_10075);
nor U15132 (N_15132,N_13470,N_11520);
nor U15133 (N_15133,N_14366,N_13017);
or U15134 (N_15134,N_14897,N_12209);
and U15135 (N_15135,N_10947,N_12727);
nor U15136 (N_15136,N_12519,N_12969);
or U15137 (N_15137,N_11180,N_11902);
nand U15138 (N_15138,N_10747,N_12654);
xor U15139 (N_15139,N_14498,N_11445);
nand U15140 (N_15140,N_11174,N_12936);
and U15141 (N_15141,N_10781,N_12567);
and U15142 (N_15142,N_11955,N_11224);
nor U15143 (N_15143,N_14471,N_11779);
nor U15144 (N_15144,N_13317,N_13093);
and U15145 (N_15145,N_10871,N_14627);
and U15146 (N_15146,N_12590,N_10817);
nand U15147 (N_15147,N_13210,N_10114);
nand U15148 (N_15148,N_10013,N_11656);
or U15149 (N_15149,N_11606,N_13326);
nand U15150 (N_15150,N_13656,N_10219);
or U15151 (N_15151,N_10467,N_13424);
xor U15152 (N_15152,N_11775,N_14926);
nor U15153 (N_15153,N_10405,N_11001);
xnor U15154 (N_15154,N_13618,N_12638);
or U15155 (N_15155,N_14270,N_13099);
xnor U15156 (N_15156,N_11513,N_10032);
and U15157 (N_15157,N_11874,N_11164);
xnor U15158 (N_15158,N_10906,N_11079);
nor U15159 (N_15159,N_10158,N_10234);
nand U15160 (N_15160,N_14718,N_12661);
xnor U15161 (N_15161,N_14371,N_11388);
or U15162 (N_15162,N_10398,N_14745);
and U15163 (N_15163,N_14315,N_10189);
or U15164 (N_15164,N_13428,N_11322);
xor U15165 (N_15165,N_14224,N_10243);
or U15166 (N_15166,N_14306,N_13253);
and U15167 (N_15167,N_12625,N_12111);
or U15168 (N_15168,N_10451,N_14971);
nand U15169 (N_15169,N_12691,N_11599);
nand U15170 (N_15170,N_14053,N_12581);
nand U15171 (N_15171,N_11999,N_10936);
nor U15172 (N_15172,N_10002,N_10910);
xnor U15173 (N_15173,N_12792,N_13242);
and U15174 (N_15174,N_12436,N_11589);
and U15175 (N_15175,N_11879,N_12043);
or U15176 (N_15176,N_14343,N_11244);
nor U15177 (N_15177,N_12345,N_12830);
or U15178 (N_15178,N_14379,N_10632);
and U15179 (N_15179,N_14831,N_11352);
nand U15180 (N_15180,N_14226,N_12447);
nor U15181 (N_15181,N_13819,N_11536);
and U15182 (N_15182,N_10573,N_10613);
xor U15183 (N_15183,N_13665,N_12930);
nand U15184 (N_15184,N_11214,N_10699);
xnor U15185 (N_15185,N_14395,N_13565);
or U15186 (N_15186,N_11184,N_11862);
xor U15187 (N_15187,N_14028,N_14676);
nor U15188 (N_15188,N_10392,N_14782);
or U15189 (N_15189,N_13626,N_13164);
nand U15190 (N_15190,N_13288,N_14254);
nor U15191 (N_15191,N_12582,N_13976);
nor U15192 (N_15192,N_14015,N_13132);
nor U15193 (N_15193,N_10012,N_11468);
nand U15194 (N_15194,N_12958,N_10069);
nor U15195 (N_15195,N_12524,N_10863);
nor U15196 (N_15196,N_12462,N_10439);
and U15197 (N_15197,N_14445,N_10063);
xnor U15198 (N_15198,N_10474,N_10769);
nand U15199 (N_15199,N_11006,N_14483);
nand U15200 (N_15200,N_11491,N_10064);
nor U15201 (N_15201,N_12646,N_10132);
nand U15202 (N_15202,N_12309,N_11399);
nand U15203 (N_15203,N_10119,N_14122);
xnor U15204 (N_15204,N_11756,N_14609);
or U15205 (N_15205,N_13296,N_14650);
nand U15206 (N_15206,N_12532,N_14796);
nand U15207 (N_15207,N_12009,N_12214);
nand U15208 (N_15208,N_13632,N_10008);
nor U15209 (N_15209,N_11713,N_10765);
and U15210 (N_15210,N_12319,N_13874);
or U15211 (N_15211,N_14223,N_12391);
and U15212 (N_15212,N_13767,N_14126);
and U15213 (N_15213,N_14302,N_13850);
nand U15214 (N_15214,N_12708,N_13953);
nand U15215 (N_15215,N_12117,N_11007);
nand U15216 (N_15216,N_13098,N_14918);
and U15217 (N_15217,N_11849,N_10369);
and U15218 (N_15218,N_12186,N_12704);
nor U15219 (N_15219,N_11105,N_11487);
xor U15220 (N_15220,N_13400,N_10917);
nor U15221 (N_15221,N_10987,N_12474);
or U15222 (N_15222,N_10180,N_14418);
and U15223 (N_15223,N_12995,N_12863);
and U15224 (N_15224,N_10698,N_13449);
nor U15225 (N_15225,N_10253,N_11199);
nor U15226 (N_15226,N_10328,N_10186);
nor U15227 (N_15227,N_12047,N_11031);
and U15228 (N_15228,N_13841,N_12731);
nor U15229 (N_15229,N_11927,N_13936);
or U15230 (N_15230,N_12498,N_13406);
xor U15231 (N_15231,N_14443,N_12149);
or U15232 (N_15232,N_13142,N_11316);
or U15233 (N_15233,N_13230,N_14727);
nor U15234 (N_15234,N_12351,N_12817);
or U15235 (N_15235,N_11312,N_11757);
nor U15236 (N_15236,N_14345,N_12207);
xor U15237 (N_15237,N_14935,N_10214);
nor U15238 (N_15238,N_11590,N_13323);
or U15239 (N_15239,N_12978,N_14208);
xor U15240 (N_15240,N_10737,N_11193);
and U15241 (N_15241,N_12053,N_14378);
nor U15242 (N_15242,N_12470,N_10465);
nand U15243 (N_15243,N_10607,N_13267);
and U15244 (N_15244,N_13381,N_14697);
xor U15245 (N_15245,N_11550,N_13231);
and U15246 (N_15246,N_10228,N_10819);
and U15247 (N_15247,N_11238,N_10574);
nand U15248 (N_15248,N_12039,N_11030);
nand U15249 (N_15249,N_12080,N_10049);
xnor U15250 (N_15250,N_11851,N_13589);
or U15251 (N_15251,N_11778,N_12926);
nand U15252 (N_15252,N_12805,N_11586);
or U15253 (N_15253,N_11906,N_13868);
or U15254 (N_15254,N_10815,N_13131);
nand U15255 (N_15255,N_12899,N_13412);
and U15256 (N_15256,N_10146,N_11231);
nand U15257 (N_15257,N_14836,N_12979);
and U15258 (N_15258,N_11053,N_13085);
xnor U15259 (N_15259,N_12689,N_12405);
or U15260 (N_15260,N_13102,N_12184);
or U15261 (N_15261,N_13985,N_10591);
or U15262 (N_15262,N_14139,N_12095);
or U15263 (N_15263,N_14847,N_11975);
xor U15264 (N_15264,N_12776,N_13981);
or U15265 (N_15265,N_14191,N_14098);
nand U15266 (N_15266,N_13537,N_10301);
or U15267 (N_15267,N_13224,N_13336);
nor U15268 (N_15268,N_12705,N_10276);
or U15269 (N_15269,N_12915,N_10060);
nand U15270 (N_15270,N_12892,N_14881);
and U15271 (N_15271,N_11887,N_14173);
nor U15272 (N_15272,N_11648,N_12228);
and U15273 (N_15273,N_10325,N_13150);
nand U15274 (N_15274,N_12538,N_12983);
nand U15275 (N_15275,N_11939,N_13706);
or U15276 (N_15276,N_14725,N_11113);
nand U15277 (N_15277,N_13310,N_13019);
nand U15278 (N_15278,N_11518,N_13485);
nor U15279 (N_15279,N_11591,N_14844);
nor U15280 (N_15280,N_14726,N_13766);
or U15281 (N_15281,N_12707,N_10611);
or U15282 (N_15282,N_10696,N_11160);
nand U15283 (N_15283,N_14879,N_10233);
nor U15284 (N_15284,N_12693,N_12278);
xnor U15285 (N_15285,N_12710,N_11637);
nand U15286 (N_15286,N_12136,N_11966);
xor U15287 (N_15287,N_14925,N_14915);
nor U15288 (N_15288,N_14615,N_11456);
or U15289 (N_15289,N_10391,N_10796);
nor U15290 (N_15290,N_11000,N_14282);
xnor U15291 (N_15291,N_10533,N_14335);
nor U15292 (N_15292,N_11993,N_10305);
or U15293 (N_15293,N_14225,N_10966);
or U15294 (N_15294,N_14081,N_10394);
nand U15295 (N_15295,N_13349,N_10856);
nand U15296 (N_15296,N_14175,N_12725);
and U15297 (N_15297,N_12993,N_12196);
nand U15298 (N_15298,N_14978,N_14626);
and U15299 (N_15299,N_14564,N_13360);
nor U15300 (N_15300,N_11646,N_13081);
xnor U15301 (N_15301,N_10360,N_14172);
and U15302 (N_15302,N_11155,N_13713);
and U15303 (N_15303,N_10210,N_12082);
and U15304 (N_15304,N_12148,N_12102);
xor U15305 (N_15305,N_13603,N_12595);
nand U15306 (N_15306,N_13550,N_14194);
or U15307 (N_15307,N_14522,N_11732);
or U15308 (N_15308,N_10581,N_11542);
nand U15309 (N_15309,N_14965,N_12697);
xnor U15310 (N_15310,N_11486,N_14505);
nor U15311 (N_15311,N_11205,N_12531);
or U15312 (N_15312,N_11149,N_11544);
nor U15313 (N_15313,N_13559,N_14944);
xor U15314 (N_15314,N_12211,N_11547);
or U15315 (N_15315,N_10426,N_11744);
and U15316 (N_15316,N_10030,N_11769);
and U15317 (N_15317,N_14108,N_14514);
xor U15318 (N_15318,N_10414,N_10761);
or U15319 (N_15319,N_14065,N_12850);
and U15320 (N_15320,N_10144,N_12063);
or U15321 (N_15321,N_11626,N_11791);
nand U15322 (N_15322,N_14704,N_13174);
nand U15323 (N_15323,N_14436,N_13029);
nand U15324 (N_15324,N_14792,N_11504);
nand U15325 (N_15325,N_11039,N_11797);
or U15326 (N_15326,N_11658,N_11943);
nor U15327 (N_15327,N_13293,N_12801);
and U15328 (N_15328,N_14930,N_14914);
or U15329 (N_15329,N_14261,N_13392);
nor U15330 (N_15330,N_13905,N_10015);
nand U15331 (N_15331,N_12876,N_12073);
and U15332 (N_15332,N_14818,N_13923);
or U15333 (N_15333,N_11961,N_12879);
nor U15334 (N_15334,N_14692,N_10436);
nor U15335 (N_15335,N_10123,N_12833);
nor U15336 (N_15336,N_11915,N_10230);
nor U15337 (N_15337,N_10355,N_12586);
and U15338 (N_15338,N_13667,N_11204);
nand U15339 (N_15339,N_13964,N_12489);
nand U15340 (N_15340,N_12611,N_14712);
nor U15341 (N_15341,N_14889,N_12651);
nand U15342 (N_15342,N_12399,N_13049);
nor U15343 (N_15343,N_12700,N_13640);
nand U15344 (N_15344,N_10371,N_12052);
and U15345 (N_15345,N_12624,N_13271);
nand U15346 (N_15346,N_10750,N_10011);
nand U15347 (N_15347,N_11963,N_14482);
nand U15348 (N_15348,N_13802,N_10232);
and U15349 (N_15349,N_10455,N_10337);
and U15350 (N_15350,N_12675,N_12045);
and U15351 (N_15351,N_11087,N_12974);
nor U15352 (N_15352,N_14815,N_14460);
and U15353 (N_15353,N_13484,N_14828);
nor U15354 (N_15354,N_10480,N_12181);
and U15355 (N_15355,N_12127,N_11329);
and U15356 (N_15356,N_10708,N_11837);
nand U15357 (N_15357,N_11634,N_11376);
nor U15358 (N_15358,N_14317,N_14574);
nand U15359 (N_15359,N_14504,N_11790);
xor U15360 (N_15360,N_14907,N_11046);
nor U15361 (N_15361,N_13307,N_12160);
and U15362 (N_15362,N_14706,N_14213);
and U15363 (N_15363,N_13095,N_11907);
nand U15364 (N_15364,N_10062,N_10444);
or U15365 (N_15365,N_12367,N_14608);
and U15366 (N_15366,N_14582,N_12086);
and U15367 (N_15367,N_14865,N_14234);
nand U15368 (N_15368,N_14526,N_13987);
nand U15369 (N_15369,N_12395,N_11481);
xor U15370 (N_15370,N_14746,N_11263);
xor U15371 (N_15371,N_13045,N_13502);
nor U15372 (N_15372,N_12274,N_11097);
nor U15373 (N_15373,N_13605,N_14975);
nor U15374 (N_15374,N_12240,N_10657);
xor U15375 (N_15375,N_11764,N_14761);
nor U15376 (N_15376,N_13920,N_11134);
nor U15377 (N_15377,N_12887,N_12766);
nor U15378 (N_15378,N_12205,N_12530);
xor U15379 (N_15379,N_11888,N_10127);
nor U15380 (N_15380,N_10194,N_11737);
and U15381 (N_15381,N_11361,N_12303);
or U15382 (N_15382,N_10499,N_12026);
and U15383 (N_15383,N_11770,N_14846);
nand U15384 (N_15384,N_12613,N_10932);
or U15385 (N_15385,N_10712,N_13035);
nor U15386 (N_15386,N_12459,N_14778);
nand U15387 (N_15387,N_13770,N_11440);
or U15388 (N_15388,N_12607,N_10904);
xnor U15389 (N_15389,N_10602,N_13619);
nand U15390 (N_15390,N_11704,N_10524);
nor U15391 (N_15391,N_12975,N_11912);
nand U15392 (N_15392,N_11317,N_12795);
nand U15393 (N_15393,N_11552,N_10227);
nand U15394 (N_15394,N_13365,N_10535);
xor U15395 (N_15395,N_12787,N_13480);
xnor U15396 (N_15396,N_10683,N_14643);
or U15397 (N_15397,N_14328,N_13477);
xnor U15398 (N_15398,N_13651,N_10789);
nor U15399 (N_15399,N_12554,N_11476);
and U15400 (N_15400,N_11302,N_10575);
nand U15401 (N_15401,N_14323,N_12408);
nor U15402 (N_15402,N_10929,N_12756);
or U15403 (N_15403,N_11609,N_14034);
and U15404 (N_15404,N_13729,N_12201);
nand U15405 (N_15405,N_10007,N_11633);
nor U15406 (N_15406,N_12241,N_12672);
nand U15407 (N_15407,N_10724,N_10251);
or U15408 (N_15408,N_14592,N_13512);
and U15409 (N_15409,N_10685,N_14838);
nand U15410 (N_15410,N_14050,N_12384);
xor U15411 (N_15411,N_11353,N_12502);
nand U15412 (N_15412,N_10622,N_10131);
or U15413 (N_15413,N_12985,N_10018);
or U15414 (N_15414,N_10621,N_10278);
nor U15415 (N_15415,N_14164,N_11405);
nor U15416 (N_15416,N_11511,N_14665);
nand U15417 (N_15417,N_14921,N_11153);
or U15418 (N_15418,N_13662,N_11689);
nand U15419 (N_15419,N_12171,N_11822);
nand U15420 (N_15420,N_10040,N_13075);
and U15421 (N_15421,N_14073,N_14553);
nor U15422 (N_15422,N_13570,N_10366);
nor U15423 (N_15423,N_11356,N_11458);
nor U15424 (N_15424,N_10280,N_11192);
and U15425 (N_15425,N_10303,N_14189);
nor U15426 (N_15426,N_13529,N_11535);
nor U15427 (N_15427,N_11117,N_13891);
or U15428 (N_15428,N_11572,N_12091);
or U15429 (N_15429,N_10494,N_13930);
and U15430 (N_15430,N_10937,N_10743);
xor U15431 (N_15431,N_13302,N_14929);
nand U15432 (N_15432,N_10609,N_10269);
or U15433 (N_15433,N_11944,N_11320);
nand U15434 (N_15434,N_14450,N_14817);
nor U15435 (N_15435,N_14834,N_12810);
or U15436 (N_15436,N_10420,N_14673);
nor U15437 (N_15437,N_12302,N_13937);
nor U15438 (N_15438,N_12905,N_14515);
xnor U15439 (N_15439,N_14851,N_12011);
xnor U15440 (N_15440,N_12110,N_10077);
and U15441 (N_15441,N_12288,N_11429);
and U15442 (N_15442,N_14327,N_13994);
or U15443 (N_15443,N_14566,N_13252);
nand U15444 (N_15444,N_12562,N_12195);
or U15445 (N_15445,N_10543,N_12962);
or U15446 (N_15446,N_13862,N_12006);
nor U15447 (N_15447,N_10279,N_12916);
or U15448 (N_15448,N_11054,N_10749);
nand U15449 (N_15449,N_11189,N_12637);
nor U15450 (N_15450,N_11901,N_12132);
nand U15451 (N_15451,N_13229,N_13808);
nand U15452 (N_15452,N_13143,N_12719);
or U15453 (N_15453,N_13118,N_11091);
and U15454 (N_15454,N_10282,N_14474);
nor U15455 (N_15455,N_13384,N_14154);
nor U15456 (N_15456,N_14113,N_14429);
and U15457 (N_15457,N_11080,N_10190);
nor U15458 (N_15458,N_12004,N_13593);
or U15459 (N_15459,N_14103,N_10338);
or U15460 (N_15460,N_11068,N_10918);
or U15461 (N_15461,N_11801,N_13000);
nor U15462 (N_15462,N_11145,N_14716);
or U15463 (N_15463,N_10555,N_14747);
xor U15464 (N_15464,N_10559,N_10098);
and U15465 (N_15465,N_13790,N_10713);
and U15466 (N_15466,N_12864,N_13511);
or U15467 (N_15467,N_14750,N_12429);
nor U15468 (N_15468,N_12218,N_14703);
nand U15469 (N_15469,N_10445,N_10095);
nand U15470 (N_15470,N_12948,N_12353);
and U15471 (N_15471,N_14922,N_14760);
nand U15472 (N_15472,N_14048,N_10192);
nor U15473 (N_15473,N_12813,N_13237);
nor U15474 (N_15474,N_10998,N_13172);
or U15475 (N_15475,N_14316,N_10263);
and U15476 (N_15476,N_13439,N_12760);
nor U15477 (N_15477,N_13573,N_10333);
xor U15478 (N_15478,N_11426,N_10909);
and U15479 (N_15479,N_10091,N_10828);
or U15480 (N_15480,N_10229,N_13974);
xor U15481 (N_15481,N_11787,N_14812);
and U15482 (N_15482,N_12816,N_12794);
nand U15483 (N_15483,N_10472,N_11367);
or U15484 (N_15484,N_11058,N_11712);
or U15485 (N_15485,N_14170,N_12903);
nor U15486 (N_15486,N_13491,N_11556);
nor U15487 (N_15487,N_10370,N_11342);
and U15488 (N_15488,N_11703,N_12678);
nand U15489 (N_15489,N_14243,N_12330);
and U15490 (N_15490,N_12706,N_10583);
nand U15491 (N_15491,N_12443,N_11628);
nand U15492 (N_15492,N_11690,N_14111);
nand U15493 (N_15493,N_10302,N_11364);
and U15494 (N_15494,N_11953,N_11600);
or U15495 (N_15495,N_11823,N_11508);
xnor U15496 (N_15496,N_12655,N_11821);
and U15497 (N_15497,N_12769,N_13803);
nor U15498 (N_15498,N_11624,N_10171);
nor U15499 (N_15499,N_12568,N_12336);
or U15500 (N_15500,N_13094,N_13463);
and U15501 (N_15501,N_12914,N_14104);
and U15502 (N_15502,N_14783,N_14919);
nor U15503 (N_15503,N_12125,N_10891);
nand U15504 (N_15504,N_12950,N_10039);
or U15505 (N_15505,N_14241,N_12873);
nand U15506 (N_15506,N_10122,N_14732);
or U15507 (N_15507,N_11397,N_14799);
and U15508 (N_15508,N_13886,N_14625);
or U15509 (N_15509,N_10938,N_11271);
nor U15510 (N_15510,N_11159,N_10389);
or U15511 (N_15511,N_13918,N_12584);
or U15512 (N_15512,N_10731,N_13047);
and U15513 (N_15513,N_12005,N_10885);
or U15514 (N_15514,N_14616,N_14976);
and U15515 (N_15515,N_11951,N_10975);
nand U15516 (N_15516,N_14421,N_10402);
and U15517 (N_15517,N_10884,N_14764);
or U15518 (N_15518,N_11740,N_11400);
nand U15519 (N_15519,N_14227,N_11392);
and U15520 (N_15520,N_11443,N_14045);
nor U15521 (N_15521,N_14757,N_14632);
and U15522 (N_15522,N_12550,N_10509);
and U15523 (N_15523,N_11891,N_14478);
nand U15524 (N_15524,N_13611,N_11521);
xnor U15525 (N_15525,N_14004,N_10151);
nor U15526 (N_15526,N_11503,N_14503);
nand U15527 (N_15527,N_13588,N_14668);
nand U15528 (N_15528,N_10427,N_13544);
nor U15529 (N_15529,N_13927,N_14219);
nor U15530 (N_15530,N_11693,N_12559);
nor U15531 (N_15531,N_10732,N_11843);
and U15532 (N_15532,N_13402,N_12861);
xor U15533 (N_15533,N_13429,N_14333);
or U15534 (N_15534,N_10625,N_11258);
or U15535 (N_15535,N_14292,N_14694);
nor U15536 (N_15536,N_10848,N_14717);
and U15537 (N_15537,N_14994,N_14131);
and U15538 (N_15538,N_13764,N_11865);
nand U15539 (N_15539,N_10469,N_14403);
or U15540 (N_15540,N_11409,N_10406);
nor U15541 (N_15541,N_10779,N_14749);
nand U15542 (N_15542,N_13201,N_13175);
or U15543 (N_15543,N_10951,N_10764);
and U15544 (N_15544,N_10173,N_14605);
and U15545 (N_15545,N_13663,N_11050);
and U15546 (N_15546,N_13103,N_14571);
xor U15547 (N_15547,N_13878,N_13989);
nor U15548 (N_15548,N_14078,N_14059);
nand U15549 (N_15549,N_10313,N_12220);
or U15550 (N_15550,N_10156,N_10023);
nor U15551 (N_15551,N_14128,N_11583);
nand U15552 (N_15552,N_14891,N_14397);
nor U15553 (N_15553,N_13104,N_11995);
and U15554 (N_15554,N_13951,N_13420);
and U15555 (N_15555,N_12904,N_11266);
or U15556 (N_15556,N_10318,N_13694);
xnor U15557 (N_15557,N_13601,N_14601);
nor U15558 (N_15558,N_12821,N_11365);
nor U15559 (N_15559,N_14305,N_13746);
nand U15560 (N_15560,N_10950,N_11137);
nand U15561 (N_15561,N_14721,N_14529);
and U15562 (N_15562,N_12844,N_14043);
xnor U15563 (N_15563,N_14123,N_11772);
or U15564 (N_15564,N_13860,N_13120);
nand U15565 (N_15565,N_11800,N_11464);
or U15566 (N_15566,N_14485,N_13203);
and U15567 (N_15567,N_13263,N_13939);
and U15568 (N_15568,N_10215,N_14461);
and U15569 (N_15569,N_10927,N_14985);
or U15570 (N_15570,N_13226,N_10357);
nand U15571 (N_15571,N_13411,N_13377);
or U15572 (N_15572,N_12370,N_12401);
xor U15573 (N_15573,N_13359,N_14543);
and U15574 (N_15574,N_13197,N_14466);
or U15575 (N_15575,N_14488,N_13795);
nand U15576 (N_15576,N_13220,N_10385);
nor U15577 (N_15577,N_11363,N_13382);
nand U15578 (N_15578,N_12164,N_13388);
nand U15579 (N_15579,N_13287,N_11826);
nand U15580 (N_15580,N_10778,N_13109);
nor U15581 (N_15581,N_13892,N_13395);
xnor U15582 (N_15582,N_13251,N_12452);
or U15583 (N_15583,N_11236,N_11872);
or U15584 (N_15584,N_11433,N_12516);
xor U15585 (N_15585,N_11473,N_10889);
or U15586 (N_15586,N_10193,N_12963);
xnor U15587 (N_15587,N_12457,N_12112);
nor U15588 (N_15588,N_11227,N_14785);
nor U15589 (N_15589,N_11928,N_10744);
nand U15590 (N_15590,N_14210,N_10869);
and U15591 (N_15591,N_13934,N_11873);
nand U15592 (N_15592,N_10719,N_14085);
nor U15593 (N_15593,N_11867,N_10425);
or U15594 (N_15594,N_11037,N_11638);
or U15595 (N_15595,N_11207,N_14857);
nand U15596 (N_15596,N_11734,N_14312);
and U15597 (N_15597,N_14708,N_12250);
nor U15598 (N_15598,N_11208,N_10925);
or U15599 (N_15599,N_10714,N_14674);
and U15600 (N_15600,N_12239,N_13861);
nand U15601 (N_15601,N_10348,N_10701);
nor U15602 (N_15602,N_10457,N_12988);
and U15603 (N_15603,N_10275,N_13633);
and U15604 (N_15604,N_13975,N_11333);
xor U15605 (N_15605,N_14822,N_12493);
or U15606 (N_15606,N_12297,N_14069);
nor U15607 (N_15607,N_12490,N_13240);
nand U15608 (N_15608,N_12304,N_14145);
xnor U15609 (N_15609,N_10688,N_14870);
nand U15610 (N_15610,N_14779,N_10068);
or U15611 (N_15611,N_11123,N_10364);
nand U15612 (N_15612,N_12393,N_12306);
and U15613 (N_15613,N_14562,N_12499);
xnor U15614 (N_15614,N_10307,N_11127);
and U15615 (N_15615,N_13840,N_14021);
or U15616 (N_15616,N_13696,N_12990);
xnor U15617 (N_15617,N_14497,N_13787);
and U15618 (N_15618,N_14672,N_12789);
nand U15619 (N_15619,N_12714,N_11135);
and U15620 (N_15620,N_11148,N_10600);
or U15621 (N_15621,N_13991,N_11957);
nor U15622 (N_15622,N_14400,N_12169);
or U15623 (N_15623,N_11056,N_13170);
and U15624 (N_15624,N_14140,N_14297);
and U15625 (N_15625,N_11188,N_12832);
and U15626 (N_15626,N_10462,N_11594);
or U15627 (N_15627,N_10514,N_10623);
or U15628 (N_15628,N_10994,N_14585);
and U15629 (N_15629,N_10393,N_10878);
and U15630 (N_15630,N_14392,N_10914);
nand U15631 (N_15631,N_11761,N_13483);
and U15632 (N_15632,N_11241,N_14776);
nand U15633 (N_15633,N_10671,N_12056);
nand U15634 (N_15634,N_12847,N_12155);
or U15635 (N_15635,N_11483,N_13775);
or U15636 (N_15636,N_10334,N_10970);
or U15637 (N_15637,N_14417,N_12042);
nor U15638 (N_15638,N_13216,N_12843);
xor U15639 (N_15639,N_10247,N_12147);
xor U15640 (N_15640,N_11278,N_11576);
xnor U15641 (N_15641,N_10409,N_14402);
or U15642 (N_15642,N_14731,N_14001);
and U15643 (N_15643,N_11131,N_11705);
nand U15644 (N_15644,N_10311,N_14805);
or U15645 (N_15645,N_10805,N_13198);
nor U15646 (N_15646,N_12135,N_14909);
nor U15647 (N_15647,N_12592,N_10290);
and U15648 (N_15648,N_13292,N_13299);
nand U15649 (N_15649,N_11834,N_11109);
and U15650 (N_15650,N_10223,N_14201);
nor U15651 (N_15651,N_11651,N_12889);
nand U15652 (N_15652,N_14293,N_13167);
and U15653 (N_15653,N_11482,N_13304);
and U15654 (N_15654,N_11981,N_12392);
nor U15655 (N_15655,N_14321,N_10523);
nand U15656 (N_15656,N_12126,N_14289);
or U15657 (N_15657,N_14284,N_14653);
and U15658 (N_15658,N_11407,N_10054);
nand U15659 (N_15659,N_14893,N_13389);
or U15660 (N_15660,N_14296,N_10407);
nand U15661 (N_15661,N_11292,N_13154);
nor U15662 (N_15662,N_11758,N_13548);
or U15663 (N_15663,N_12596,N_12368);
nor U15664 (N_15664,N_14607,N_11818);
xor U15665 (N_15665,N_11343,N_14931);
nand U15666 (N_15666,N_13277,N_11018);
nand U15667 (N_15667,N_13622,N_10770);
and U15668 (N_15668,N_10554,N_10396);
and U15669 (N_15669,N_14957,N_13947);
xor U15670 (N_15670,N_14455,N_14666);
nand U15671 (N_15671,N_10604,N_13644);
nor U15672 (N_15672,N_10112,N_12525);
nand U15673 (N_15673,N_13604,N_10960);
nor U15674 (N_15674,N_12822,N_12734);
nor U15675 (N_15675,N_14715,N_11937);
xor U15676 (N_15676,N_11013,N_10592);
or U15677 (N_15677,N_10658,N_10887);
or U15678 (N_15678,N_14500,N_13280);
nor U15679 (N_15679,N_13169,N_11664);
and U15680 (N_15680,N_10452,N_12901);
and U15681 (N_15681,N_13903,N_11530);
nor U15682 (N_15682,N_11332,N_10624);
or U15683 (N_15683,N_11554,N_12481);
nand U15684 (N_15684,N_11601,N_12815);
or U15685 (N_15685,N_11300,N_13316);
and U15686 (N_15686,N_12563,N_14682);
nor U15687 (N_15687,N_10710,N_12547);
or U15688 (N_15688,N_10941,N_13027);
nand U15689 (N_15689,N_13504,N_12325);
nor U15690 (N_15690,N_11825,N_10150);
nand U15691 (N_15691,N_10484,N_14551);
nor U15692 (N_15692,N_11280,N_12450);
nor U15693 (N_15693,N_10401,N_13676);
or U15694 (N_15694,N_12093,N_11128);
xor U15695 (N_15695,N_11675,N_13967);
xnor U15696 (N_15696,N_10754,N_14868);
or U15697 (N_15697,N_11379,N_13966);
or U15698 (N_15698,N_13004,N_14547);
nand U15699 (N_15699,N_14880,N_10249);
or U15700 (N_15700,N_13464,N_14641);
nand U15701 (N_15701,N_10288,N_13440);
nor U15702 (N_15702,N_13116,N_10777);
nor U15703 (N_15703,N_12165,N_12258);
nand U15704 (N_15704,N_11558,N_11835);
and U15705 (N_15705,N_10926,N_13121);
nand U15706 (N_15706,N_13954,N_14331);
nand U15707 (N_15707,N_14693,N_11692);
or U15708 (N_15708,N_10504,N_14956);
or U15709 (N_15709,N_11125,N_13437);
xor U15710 (N_15710,N_11178,N_14521);
and U15711 (N_15711,N_13952,N_12552);
nor U15712 (N_15712,N_14900,N_11183);
xnor U15713 (N_15713,N_13282,N_11450);
or U15714 (N_15714,N_10491,N_13265);
and U15715 (N_15715,N_12814,N_12464);
nand U15716 (N_15716,N_12482,N_10875);
nand U15717 (N_15717,N_10895,N_13376);
nor U15718 (N_15718,N_11413,N_10365);
xor U15719 (N_15719,N_13715,N_13176);
nand U15720 (N_15720,N_12066,N_12438);
and U15721 (N_15721,N_10563,N_12802);
nor U15722 (N_15722,N_10336,N_14705);
or U15723 (N_15723,N_11416,N_12357);
xor U15724 (N_15724,N_12600,N_13777);
xnor U15725 (N_15725,N_11751,N_14895);
or U15726 (N_15726,N_13457,N_12740);
xor U15727 (N_15727,N_10164,N_11448);
nor U15728 (N_15728,N_14802,N_10677);
nand U15729 (N_15729,N_10760,N_11753);
xor U15730 (N_15730,N_13505,N_14229);
or U15731 (N_15731,N_11531,N_10976);
or U15732 (N_15732,N_11459,N_10670);
and U15733 (N_15733,N_11808,N_14644);
nand U15734 (N_15734,N_11069,N_11452);
nand U15735 (N_15735,N_11308,N_11310);
nor U15736 (N_15736,N_10493,N_10440);
nand U15737 (N_15737,N_14563,N_11655);
xor U15738 (N_15738,N_10314,N_10446);
and U15739 (N_15739,N_13579,N_13159);
xor U15740 (N_15740,N_12222,N_12628);
nand U15741 (N_15741,N_10605,N_12884);
or U15742 (N_15742,N_13180,N_11688);
and U15743 (N_15743,N_11738,N_12458);
and U15744 (N_15744,N_11012,N_10272);
nand U15745 (N_15745,N_11175,N_10859);
and U15746 (N_15746,N_12504,N_11107);
nand U15747 (N_15747,N_12682,N_12020);
or U15748 (N_15748,N_11274,N_13735);
xnor U15749 (N_15749,N_12227,N_14695);
nor U15750 (N_15750,N_10296,N_13246);
nand U15751 (N_15751,N_11434,N_12090);
or U15752 (N_15752,N_10867,N_12415);
nand U15753 (N_15753,N_14807,N_14869);
and U15754 (N_15754,N_13023,N_14617);
xnor U15755 (N_15755,N_11839,N_12569);
nor U15756 (N_15756,N_13273,N_12406);
nand U15757 (N_15757,N_12599,N_10993);
and U15758 (N_15758,N_11929,N_12226);
or U15759 (N_15759,N_14094,N_12604);
nand U15760 (N_15760,N_11454,N_11828);
nand U15761 (N_15761,N_14438,N_11026);
nand U15762 (N_15762,N_11219,N_14158);
nand U15763 (N_15763,N_14663,N_14968);
nand U15764 (N_15764,N_14736,N_12783);
and U15765 (N_15765,N_13785,N_14575);
and U15766 (N_15766,N_11287,N_10900);
or U15767 (N_15767,N_10078,N_13747);
nand U15768 (N_15768,N_14072,N_12622);
nand U15769 (N_15769,N_10962,N_12386);
and U15770 (N_15770,N_12653,N_14102);
and U15771 (N_15771,N_12973,N_13125);
or U15772 (N_15772,N_12517,N_10408);
nand U15773 (N_15773,N_14756,N_12775);
and U15774 (N_15774,N_11742,N_13621);
nor U15775 (N_15775,N_14584,N_13845);
or U15776 (N_15776,N_13057,N_13066);
and U15777 (N_15777,N_14788,N_14148);
xnor U15778 (N_15778,N_14160,N_14178);
and U15779 (N_15779,N_12786,N_12223);
and U15780 (N_15780,N_12413,N_14960);
or U15781 (N_15781,N_11684,N_12649);
nor U15782 (N_15782,N_14649,N_13284);
or U15783 (N_15783,N_10179,N_12997);
nand U15784 (N_15784,N_10693,N_13731);
or U15785 (N_15785,N_13942,N_11745);
or U15786 (N_15786,N_13308,N_10662);
xnor U15787 (N_15787,N_14247,N_13629);
nand U15788 (N_15788,N_11602,N_10529);
nor U15789 (N_15789,N_11499,N_11152);
and U15790 (N_15790,N_11918,N_12369);
xnor U15791 (N_15791,N_11494,N_11071);
and U15792 (N_15792,N_13852,N_12548);
or U15793 (N_15793,N_13943,N_12846);
xor U15794 (N_15794,N_11305,N_12390);
xnor U15795 (N_15795,N_14533,N_10221);
and U15796 (N_15796,N_14179,N_11910);
xnor U15797 (N_15797,N_14713,N_14830);
and U15798 (N_15798,N_10800,N_10258);
and U15799 (N_15799,N_10207,N_11025);
and U15800 (N_15800,N_14054,N_12338);
nor U15801 (N_15801,N_10707,N_14955);
nor U15802 (N_15802,N_10430,N_14751);
xnor U15803 (N_15803,N_14537,N_10271);
nor U15804 (N_15804,N_10835,N_12937);
and U15805 (N_15805,N_11331,N_13824);
or U15806 (N_15806,N_12347,N_12692);
xor U15807 (N_15807,N_13354,N_11914);
and U15808 (N_15808,N_14885,N_14686);
nand U15809 (N_15809,N_13986,N_14412);
or U15810 (N_15810,N_13171,N_10847);
nor U15811 (N_15811,N_12561,N_13931);
and U15812 (N_15812,N_13294,N_11863);
nand U15813 (N_15813,N_11868,N_13070);
and U15814 (N_15814,N_13554,N_13837);
or U15815 (N_15815,N_10730,N_12921);
and U15816 (N_15816,N_11876,N_12284);
xor U15817 (N_15817,N_10668,N_10717);
nand U15818 (N_15818,N_10120,N_12329);
nand U15819 (N_15819,N_10978,N_10224);
nand U15820 (N_15820,N_10035,N_14637);
xor U15821 (N_15821,N_13691,N_10380);
nand U15822 (N_15822,N_11629,N_13615);
or U15823 (N_15823,N_11523,N_10211);
nand U15824 (N_15824,N_14849,N_10617);
nand U15825 (N_15825,N_13712,N_12729);
or U15826 (N_15826,N_12841,N_14090);
nand U15827 (N_15827,N_10027,N_11301);
and U15828 (N_15828,N_12735,N_14555);
and U15829 (N_15829,N_10345,N_10134);
nor U15830 (N_15830,N_10154,N_10036);
nor U15831 (N_15831,N_13088,N_12098);
nor U15832 (N_15832,N_13736,N_11652);
or U15833 (N_15833,N_13414,N_13829);
xnor U15834 (N_15834,N_11905,N_12652);
nor U15835 (N_15835,N_12546,N_13031);
and U15836 (N_15836,N_10005,N_10638);
nor U15837 (N_15837,N_14567,N_14506);
or U15838 (N_15838,N_12448,N_11341);
and U15839 (N_15839,N_11627,N_12811);
or U15840 (N_15840,N_11488,N_12445);
and U15841 (N_15841,N_12544,N_13028);
or U15842 (N_15842,N_12310,N_12922);
or U15843 (N_15843,N_13911,N_11831);
nand U15844 (N_15844,N_10079,N_14032);
or U15845 (N_15845,N_12268,N_13678);
nand U15846 (N_15846,N_11892,N_10839);
nand U15847 (N_15847,N_12793,N_12644);
nand U15848 (N_15848,N_11325,N_11377);
or U15849 (N_15849,N_12856,N_14525);
and U15850 (N_15850,N_13161,N_13489);
nand U15851 (N_15851,N_13026,N_14268);
or U15852 (N_15852,N_13857,N_13339);
nor U15853 (N_15853,N_14639,N_13938);
or U15854 (N_15854,N_14290,N_12049);
and U15855 (N_15855,N_10264,N_10116);
and U15856 (N_15856,N_12378,N_10752);
xnor U15857 (N_15857,N_14107,N_11283);
xnor U15858 (N_15858,N_13879,N_12248);
or U15859 (N_15859,N_12566,N_10421);
and U15860 (N_15860,N_14545,N_14602);
and U15861 (N_15861,N_11945,N_13064);
nor U15862 (N_15862,N_10810,N_12824);
or U15863 (N_15863,N_14132,N_11485);
xnor U15864 (N_15864,N_12778,N_14301);
and U15865 (N_15865,N_10437,N_14494);
nor U15866 (N_15866,N_10695,N_14723);
xnor U15867 (N_15867,N_10961,N_12128);
nand U15868 (N_15868,N_14238,N_11802);
and U15869 (N_15869,N_13488,N_13421);
nand U15870 (N_15870,N_12381,N_10085);
nand U15871 (N_15871,N_10968,N_13689);
and U15872 (N_15872,N_12398,N_13110);
or U15873 (N_15873,N_12739,N_14251);
nand U15874 (N_15874,N_13900,N_14827);
and U15875 (N_15875,N_13961,N_10813);
nand U15876 (N_15876,N_13758,N_12087);
nor U15877 (N_15877,N_13750,N_10363);
or U15878 (N_15878,N_11306,N_14821);
nand U15879 (N_15879,N_10273,N_14249);
nand U15880 (N_15880,N_10560,N_13821);
or U15881 (N_15881,N_10454,N_10773);
nor U15882 (N_15882,N_13503,N_10152);
and U15883 (N_15883,N_12255,N_13725);
or U15884 (N_15884,N_10629,N_12032);
or U15885 (N_15885,N_13034,N_11545);
and U15886 (N_15886,N_12487,N_13160);
nand U15887 (N_15887,N_10682,N_13217);
nor U15888 (N_15888,N_14196,N_13055);
nand U15889 (N_15889,N_13784,N_10447);
nor U15890 (N_15890,N_11948,N_13100);
or U15891 (N_15891,N_12358,N_11940);
and U15892 (N_15892,N_11378,N_12860);
xor U15893 (N_15893,N_14481,N_14942);
nor U15894 (N_15894,N_10404,N_10517);
nand U15895 (N_15895,N_10200,N_14388);
or U15896 (N_15896,N_12360,N_14444);
and U15897 (N_15897,N_13702,N_11567);
nor U15898 (N_15898,N_13560,N_14386);
nor U15899 (N_15899,N_11449,N_12497);
nor U15900 (N_15900,N_13754,N_12295);
xnor U15901 (N_15901,N_10608,N_11357);
and U15902 (N_15902,N_13578,N_12564);
nor U15903 (N_15903,N_12565,N_12671);
nand U15904 (N_15904,N_13185,N_10083);
nand U15905 (N_15905,N_10274,N_10020);
or U15906 (N_15906,N_10107,N_14358);
or U15907 (N_15907,N_10433,N_13541);
or U15908 (N_15908,N_13258,N_13468);
or U15909 (N_15909,N_12116,N_10432);
or U15910 (N_15910,N_11559,N_14161);
nand U15911 (N_15911,N_11549,N_13510);
nand U15912 (N_15912,N_13922,N_12100);
nor U15913 (N_15913,N_14133,N_13778);
nor U15914 (N_15914,N_14095,N_10341);
and U15915 (N_15915,N_13397,N_12251);
nand U15916 (N_15916,N_10099,N_14710);
nor U15917 (N_15917,N_10840,N_12594);
nand U15918 (N_15918,N_11595,N_14544);
xor U15919 (N_15919,N_11996,N_14353);
or U15920 (N_15920,N_13738,N_12666);
or U15921 (N_15921,N_14634,N_14472);
or U15922 (N_15922,N_11644,N_11729);
and U15923 (N_15923,N_11904,N_10822);
or U15924 (N_15924,N_10958,N_13124);
nand U15925 (N_15925,N_12648,N_10656);
nand U15926 (N_15926,N_13630,N_13446);
nand U15927 (N_15927,N_11903,N_13972);
or U15928 (N_15928,N_11146,N_11707);
nor U15929 (N_15929,N_13854,N_10512);
nand U15930 (N_15930,N_11218,N_12882);
nand U15931 (N_15931,N_14524,N_11103);
nor U15932 (N_15932,N_12010,N_14084);
nor U15933 (N_15933,N_14759,N_14624);
or U15934 (N_15934,N_14635,N_13233);
and U15935 (N_15935,N_12167,N_14896);
nor U15936 (N_15936,N_12511,N_12736);
nand U15937 (N_15937,N_13259,N_12555);
nand U15938 (N_15938,N_12528,N_13009);
or U15939 (N_15939,N_12143,N_14561);
nand U15940 (N_15940,N_12084,N_14042);
nand U15941 (N_15941,N_10359,N_10352);
or U15942 (N_15942,N_12588,N_13475);
nand U15943 (N_15943,N_14187,N_14911);
or U15944 (N_15944,N_12507,N_14855);
or U15945 (N_15945,N_10924,N_14097);
and U15946 (N_15946,N_13516,N_10992);
xnor U15947 (N_15947,N_11023,N_11971);
nand U15948 (N_15948,N_11330,N_10735);
and U15949 (N_15949,N_10952,N_10117);
and U15950 (N_15950,N_13737,N_12383);
nand U15951 (N_15951,N_13813,N_13239);
nand U15952 (N_15952,N_13971,N_12192);
nor U15953 (N_15953,N_10377,N_13914);
nand U15954 (N_15954,N_12553,N_12750);
nor U15955 (N_15955,N_11181,N_14475);
and U15956 (N_15956,N_13108,N_11987);
nand U15957 (N_15957,N_11898,N_10939);
and U15958 (N_15958,N_11949,N_14800);
or U15959 (N_15959,N_12435,N_14894);
and U15960 (N_15960,N_14765,N_12286);
nor U15961 (N_15961,N_12621,N_12003);
nand U15962 (N_15962,N_11555,N_13347);
xor U15963 (N_15963,N_10048,N_10921);
nand U15964 (N_15964,N_12261,N_13380);
and U15965 (N_15965,N_12718,N_13155);
nor U15966 (N_15966,N_11882,N_13782);
or U15967 (N_15967,N_11479,N_12068);
and U15968 (N_15968,N_12984,N_11896);
and U15969 (N_15969,N_14744,N_12388);
nor U15970 (N_15970,N_14887,N_12605);
nor U15971 (N_15971,N_12659,N_11842);
and U15972 (N_15972,N_13734,N_10681);
nor U15973 (N_15973,N_12679,N_11381);
or U15974 (N_15974,N_10097,N_10630);
or U15975 (N_15975,N_14987,N_12685);
nor U15976 (N_15976,N_10570,N_14075);
xnor U15977 (N_15977,N_14309,N_10418);
and U15978 (N_15978,N_12540,N_13062);
or U15979 (N_15979,N_12193,N_14137);
or U15980 (N_15980,N_12007,N_12927);
nand U15981 (N_15981,N_11014,N_11991);
nor U15982 (N_15982,N_12784,N_14135);
or U15983 (N_15983,N_13291,N_10284);
nor U15984 (N_15984,N_11066,N_12845);
nor U15985 (N_15985,N_13311,N_10988);
nand U15986 (N_15986,N_14062,N_13069);
and U15987 (N_15987,N_13005,N_14176);
or U15988 (N_15988,N_14267,N_14603);
nor U15989 (N_15989,N_11697,N_10483);
or U15990 (N_15990,N_12733,N_14029);
and U15991 (N_15991,N_10374,N_11619);
and U15992 (N_15992,N_14590,N_14594);
and U15993 (N_15993,N_11766,N_12875);
nor U15994 (N_15994,N_10757,N_11247);
and U15995 (N_15995,N_14018,N_14791);
nand U15996 (N_15996,N_13042,N_11269);
nor U15997 (N_15997,N_14300,N_14009);
xnor U15998 (N_15998,N_12342,N_13628);
nand U15999 (N_15999,N_13643,N_14356);
nor U16000 (N_16000,N_10610,N_13366);
or U16001 (N_16001,N_11253,N_12907);
nand U16002 (N_16002,N_12681,N_10326);
or U16003 (N_16003,N_13177,N_11672);
nand U16004 (N_16004,N_14056,N_14239);
nor U16005 (N_16005,N_11653,N_14700);
and U16006 (N_16006,N_13956,N_14262);
or U16007 (N_16007,N_12680,N_11374);
or U16008 (N_16008,N_11884,N_12518);
nand U16009 (N_16009,N_13751,N_13194);
and U16010 (N_16010,N_13236,N_10169);
and U16011 (N_16011,N_13533,N_13329);
nor U16012 (N_16012,N_12515,N_13234);
nor U16013 (N_16013,N_11246,N_11446);
and U16014 (N_16014,N_14707,N_14938);
and U16015 (N_16015,N_10115,N_14833);
and U16016 (N_16016,N_11517,N_11691);
or U16017 (N_16017,N_10191,N_12198);
nor U16018 (N_16018,N_10544,N_11584);
or U16019 (N_16019,N_14044,N_13481);
nor U16020 (N_16020,N_10003,N_10475);
nand U16021 (N_16021,N_13598,N_12809);
nor U16022 (N_16022,N_14369,N_10118);
or U16023 (N_16023,N_12075,N_11108);
nand U16024 (N_16024,N_11314,N_10977);
or U16025 (N_16025,N_12920,N_11935);
nand U16026 (N_16026,N_13126,N_14809);
nor U16027 (N_16027,N_14913,N_13798);
or U16028 (N_16028,N_13335,N_10834);
or U16029 (N_16029,N_12939,N_14655);
xor U16030 (N_16030,N_12346,N_12023);
and U16031 (N_16031,N_14967,N_12377);
or U16032 (N_16032,N_13363,N_13462);
and U16033 (N_16033,N_11880,N_12618);
nor U16034 (N_16034,N_14404,N_11350);
nor U16035 (N_16035,N_14359,N_13897);
or U16036 (N_16036,N_11480,N_12851);
and U16037 (N_16037,N_13493,N_12048);
or U16038 (N_16038,N_14557,N_11355);
and U16039 (N_16039,N_14587,N_14910);
nor U16040 (N_16040,N_12439,N_11793);
or U16041 (N_16041,N_10572,N_13594);
xor U16042 (N_16042,N_12945,N_14339);
or U16043 (N_16043,N_10786,N_11604);
or U16044 (N_16044,N_13313,N_13863);
or U16045 (N_16045,N_10400,N_14628);
nor U16046 (N_16046,N_14832,N_12237);
or U16047 (N_16047,N_14523,N_10070);
nor U16048 (N_16048,N_10213,N_11008);
and U16049 (N_16049,N_11956,N_12956);
nand U16050 (N_16050,N_12229,N_14795);
or U16051 (N_16051,N_13331,N_12301);
xnor U16052 (N_16052,N_14231,N_10037);
nand U16053 (N_16053,N_10185,N_10802);
nand U16054 (N_16054,N_12465,N_13648);
or U16055 (N_16055,N_12154,N_12343);
or U16056 (N_16056,N_11052,N_12298);
nor U16057 (N_16057,N_10212,N_14698);
and U16058 (N_16058,N_11104,N_10076);
nor U16059 (N_16059,N_14035,N_14996);
xnor U16060 (N_16060,N_14577,N_10612);
xnor U16061 (N_16061,N_10826,N_12433);
and U16062 (N_16062,N_12853,N_14039);
and U16063 (N_16063,N_13811,N_12660);
and U16064 (N_16064,N_11217,N_11858);
or U16065 (N_16065,N_12633,N_14516);
and U16066 (N_16066,N_11425,N_10379);
and U16067 (N_16067,N_10718,N_10471);
and U16068 (N_16068,N_11447,N_11771);
and U16069 (N_16069,N_14511,N_12277);
or U16070 (N_16070,N_11960,N_14990);
and U16071 (N_16071,N_13473,N_13298);
or U16072 (N_16072,N_13129,N_10022);
nand U16073 (N_16073,N_11256,N_13518);
or U16074 (N_16074,N_11760,N_12998);
xnor U16075 (N_16075,N_12541,N_11286);
nand U16076 (N_16076,N_12854,N_13305);
xor U16077 (N_16077,N_12543,N_11958);
nand U16078 (N_16078,N_13152,N_10546);
xnor U16079 (N_16079,N_10528,N_11992);
or U16080 (N_16080,N_11129,N_13684);
nand U16081 (N_16081,N_12807,N_12918);
xor U16082 (N_16082,N_10502,N_10585);
nand U16083 (N_16083,N_12712,N_13261);
nand U16084 (N_16084,N_12094,N_11603);
xnor U16085 (N_16085,N_14781,N_14986);
nand U16086 (N_16086,N_13016,N_13178);
nand U16087 (N_16087,N_12942,N_11106);
xor U16088 (N_16088,N_13249,N_13864);
and U16089 (N_16089,N_14023,N_13929);
or U16090 (N_16090,N_14924,N_12179);
and U16091 (N_16091,N_10367,N_11755);
or U16092 (N_16092,N_12989,N_10674);
nand U16093 (N_16093,N_13191,N_14499);
nor U16094 (N_16094,N_13209,N_12919);
or U16095 (N_16095,N_14174,N_10281);
nor U16096 (N_16096,N_12204,N_11318);
nand U16097 (N_16097,N_14906,N_12488);
or U16098 (N_16098,N_12715,N_10403);
nor U16099 (N_16099,N_12523,N_13707);
nand U16100 (N_16100,N_13033,N_14542);
and U16101 (N_16101,N_11430,N_14410);
and U16102 (N_16102,N_13571,N_14886);
nor U16103 (N_16103,N_14767,N_14433);
and U16104 (N_16104,N_10963,N_12314);
or U16105 (N_16105,N_10990,N_14409);
nor U16106 (N_16106,N_12421,N_13106);
or U16107 (N_16107,N_10460,N_10140);
xnor U16108 (N_16108,N_11670,N_14079);
and U16109 (N_16109,N_13836,N_12610);
or U16110 (N_16110,N_11820,N_10862);
or U16111 (N_16111,N_11284,N_13398);
xnor U16112 (N_16112,N_12819,N_10356);
nand U16113 (N_16113,N_13909,N_12158);
nor U16114 (N_16114,N_10545,N_11788);
or U16115 (N_16115,N_10890,N_14645);
nand U16116 (N_16116,N_11469,N_13297);
nand U16117 (N_16117,N_11795,N_11575);
and U16118 (N_16118,N_10294,N_14777);
nor U16119 (N_16119,N_10399,N_12000);
nor U16120 (N_16120,N_12946,N_10167);
and U16121 (N_16121,N_13761,N_13416);
and U16122 (N_16122,N_13225,N_13901);
or U16123 (N_16123,N_11396,N_13856);
nand U16124 (N_16124,N_13321,N_12432);
or U16125 (N_16125,N_12142,N_11179);
nor U16126 (N_16126,N_14454,N_12670);
or U16127 (N_16127,N_12966,N_11041);
nor U16128 (N_16128,N_14495,N_11092);
or U16129 (N_16129,N_10231,N_14933);
and U16130 (N_16130,N_14232,N_11295);
nand U16131 (N_16131,N_10907,N_12213);
or U16132 (N_16132,N_11156,N_13820);
nand U16133 (N_16133,N_14711,N_13501);
or U16134 (N_16134,N_12276,N_13855);
or U16135 (N_16135,N_14675,N_11936);
nand U16136 (N_16136,N_13039,N_10225);
xor U16137 (N_16137,N_10080,N_10496);
and U16138 (N_16138,N_14477,N_14143);
nand U16139 (N_16139,N_10153,N_10017);
nor U16140 (N_16140,N_10295,N_13566);
nand U16141 (N_16141,N_14928,N_14367);
or U16142 (N_16142,N_13616,N_10188);
nor U16143 (N_16143,N_10982,N_14277);
nand U16144 (N_16144,N_13221,N_14873);
xor U16145 (N_16145,N_14192,N_10690);
nand U16146 (N_16146,N_10727,N_12305);
nor U16147 (N_16147,N_13068,N_14633);
and U16148 (N_16148,N_13877,N_11859);
and U16149 (N_16149,N_10238,N_13638);
and U16150 (N_16150,N_12571,N_12603);
nor U16151 (N_16151,N_11022,N_10102);
nand U16152 (N_16152,N_10553,N_11387);
nand U16153 (N_16153,N_13285,N_10149);
and U16154 (N_16154,N_14735,N_12964);
nand U16155 (N_16155,N_10945,N_11886);
nor U16156 (N_16156,N_14264,N_12573);
or U16157 (N_16157,N_11925,N_13887);
nor U16158 (N_16158,N_10157,N_10860);
xor U16159 (N_16159,N_13576,N_13454);
nand U16160 (N_16160,N_13642,N_11451);
nor U16161 (N_16161,N_10756,N_14748);
nand U16162 (N_16162,N_14228,N_12623);
and U16163 (N_16163,N_11830,N_12410);
nor U16164 (N_16164,N_13685,N_14012);
and U16165 (N_16165,N_12199,N_13426);
nor U16166 (N_16166,N_10825,N_11252);
or U16167 (N_16167,N_10703,N_14874);
nor U16168 (N_16168,N_13276,N_14871);
xor U16169 (N_16169,N_10160,N_10721);
or U16170 (N_16170,N_13535,N_10722);
nand U16171 (N_16171,N_14630,N_12269);
nor U16172 (N_16172,N_14470,N_10763);
or U16173 (N_16173,N_14853,N_13772);
nand U16174 (N_16174,N_13067,N_10882);
or U16175 (N_16175,N_14722,N_14487);
and U16176 (N_16176,N_13520,N_13895);
nor U16177 (N_16177,N_11916,N_14431);
and U16178 (N_16178,N_10026,N_14741);
or U16179 (N_16179,N_13865,N_13040);
nor U16180 (N_16180,N_13584,N_14153);
nand U16181 (N_16181,N_12161,N_12852);
nor U16182 (N_16182,N_12911,N_12893);
nand U16183 (N_16183,N_13247,N_11028);
nor U16184 (N_16184,N_11136,N_14696);
and U16185 (N_16185,N_10780,N_14982);
and U16186 (N_16186,N_14340,N_14093);
or U16187 (N_16187,N_12028,N_11019);
nor U16188 (N_16188,N_10024,N_14168);
nand U16189 (N_16189,N_12619,N_13525);
nand U16190 (N_16190,N_12139,N_11248);
and U16191 (N_16191,N_13773,N_13568);
nor U16192 (N_16192,N_10587,N_12728);
nor U16193 (N_16193,N_12500,N_11965);
and U16194 (N_16194,N_14124,N_12440);
nand U16195 (N_16195,N_10482,N_13844);
nand U16196 (N_16196,N_13563,N_11607);
nand U16197 (N_16197,N_14743,N_10903);
and U16198 (N_16198,N_12501,N_12777);
nand U16199 (N_16199,N_13608,N_13998);
or U16200 (N_16200,N_10838,N_14540);
or U16201 (N_16201,N_14337,N_14884);
nor U16202 (N_16202,N_11348,N_14341);
nand U16203 (N_16203,N_10182,N_14350);
and U16204 (N_16204,N_11726,N_12716);
nor U16205 (N_16205,N_13983,N_14368);
nor U16206 (N_16206,N_10997,N_12486);
nor U16207 (N_16207,N_14269,N_12025);
nand U16208 (N_16208,N_12943,N_11002);
nand U16209 (N_16209,N_14803,N_13403);
nand U16210 (N_16210,N_13453,N_13567);
or U16211 (N_16211,N_12070,N_11616);
or U16212 (N_16212,N_14993,N_13499);
or U16213 (N_16213,N_13669,N_11921);
nor U16214 (N_16214,N_11763,N_13144);
or U16215 (N_16215,N_14375,N_10424);
and U16216 (N_16216,N_11962,N_12355);
nand U16217 (N_16217,N_12332,N_10183);
nor U16218 (N_16218,N_11111,N_10589);
xnor U16219 (N_16219,N_10306,N_12591);
nor U16220 (N_16220,N_14804,N_11090);
or U16221 (N_16221,N_14789,N_12535);
or U16222 (N_16222,N_13149,N_13728);
xnor U16223 (N_16223,N_14941,N_10508);
nor U16224 (N_16224,N_12146,N_14623);
nand U16225 (N_16225,N_11371,N_12118);
or U16226 (N_16226,N_12589,N_14801);
nor U16227 (N_16227,N_10738,N_12182);
and U16228 (N_16228,N_13517,N_10248);
nor U16229 (N_16229,N_10375,N_13322);
xnor U16230 (N_16230,N_10395,N_10979);
or U16231 (N_16231,N_11866,N_13370);
or U16232 (N_16232,N_12934,N_14464);
nand U16233 (N_16233,N_11003,N_11072);
and U16234 (N_16234,N_12790,N_11539);
and U16235 (N_16235,N_11676,N_12881);
xnor U16236 (N_16236,N_12908,N_14037);
xor U16237 (N_16237,N_10959,N_13577);
nand U16238 (N_16238,N_13153,N_10031);
nand U16239 (N_16239,N_13123,N_12088);
or U16240 (N_16240,N_14932,N_11526);
nand U16241 (N_16241,N_13551,N_10561);
nand U16242 (N_16242,N_14377,N_11162);
xor U16243 (N_16243,N_14077,N_10310);
xor U16244 (N_16244,N_10716,N_12354);
nor U16245 (N_16245,N_12322,N_13213);
and U16246 (N_16246,N_12551,N_13105);
nor U16247 (N_16247,N_11959,N_14948);
and U16248 (N_16248,N_14294,N_11727);
or U16249 (N_16249,N_10711,N_12316);
or U16250 (N_16250,N_12156,N_12583);
or U16251 (N_16251,N_14202,N_13327);
or U16252 (N_16252,N_13726,N_14038);
nand U16253 (N_16253,N_10346,N_11047);
or U16254 (N_16254,N_11060,N_10806);
and U16255 (N_16255,N_13241,N_11877);
nand U16256 (N_16256,N_13988,N_13809);
nand U16257 (N_16257,N_14794,N_14916);
nor U16258 (N_16258,N_13227,N_14216);
and U16259 (N_16259,N_12496,N_11394);
or U16260 (N_16260,N_13826,N_13330);
nor U16261 (N_16261,N_10983,N_14411);
or U16262 (N_16262,N_14773,N_10949);
or U16263 (N_16263,N_14435,N_11048);
nand U16264 (N_16264,N_10855,N_14049);
or U16265 (N_16265,N_13206,N_12124);
or U16266 (N_16266,N_10208,N_11743);
and U16267 (N_16267,N_10811,N_11319);
nand U16268 (N_16268,N_12216,N_14136);
and U16269 (N_16269,N_14583,N_11166);
and U16270 (N_16270,N_12249,N_13324);
nor U16271 (N_16271,N_13884,N_10226);
nor U16272 (N_16272,N_10342,N_11055);
and U16273 (N_16273,N_12642,N_10793);
nor U16274 (N_16274,N_10967,N_10055);
and U16275 (N_16275,N_14618,N_14858);
and U16276 (N_16276,N_13848,N_14146);
nor U16277 (N_16277,N_10197,N_12234);
or U16278 (N_16278,N_12917,N_12333);
or U16279 (N_16279,N_10378,N_10931);
xnor U16280 (N_16280,N_14599,N_12359);
and U16281 (N_16281,N_13542,N_14322);
or U16282 (N_16282,N_14546,N_12542);
and U16283 (N_16283,N_11848,N_14549);
nand U16284 (N_16284,N_12701,N_14977);
and U16285 (N_16285,N_12579,N_13238);
nand U16286 (N_16286,N_11582,N_13823);
and U16287 (N_16287,N_12224,N_10861);
nand U16288 (N_16288,N_12334,N_12188);
xnor U16289 (N_16289,N_11563,N_13459);
nand U16290 (N_16290,N_11706,N_10165);
or U16291 (N_16291,N_12096,N_13763);
or U16292 (N_16292,N_10148,N_10726);
or U16293 (N_16293,N_11061,N_11427);
and U16294 (N_16294,N_13513,N_11418);
nand U16295 (N_16295,N_10209,N_12871);
or U16296 (N_16296,N_10880,N_13352);
or U16297 (N_16297,N_11466,N_11122);
or U16298 (N_16298,N_10235,N_13435);
nand U16299 (N_16299,N_11774,N_13405);
and U16300 (N_16300,N_14596,N_13469);
or U16301 (N_16301,N_10245,N_13408);
nor U16302 (N_16302,N_12363,N_14390);
and U16303 (N_16303,N_12527,N_11908);
nor U16304 (N_16304,N_11245,N_11560);
and U16305 (N_16305,N_11210,N_10106);
nand U16306 (N_16306,N_13915,N_10046);
nor U16307 (N_16307,N_13358,N_13631);
or U16308 (N_16308,N_10981,N_11390);
and U16309 (N_16309,N_10206,N_14016);
or U16310 (N_16310,N_13456,N_14372);
or U16311 (N_16311,N_12071,N_14496);
xnor U16312 (N_16312,N_12521,N_12940);
nor U16313 (N_16313,N_12206,N_13211);
or U16314 (N_16314,N_10651,N_12266);
or U16315 (N_16315,N_14589,N_12315);
and U16316 (N_16316,N_12570,N_14307);
nor U16317 (N_16317,N_12677,N_14091);
or U16318 (N_16318,N_11372,N_12219);
and U16319 (N_16319,N_10014,N_10841);
xnor U16320 (N_16320,N_10911,N_10172);
nor U16321 (N_16321,N_10593,N_12503);
xor U16322 (N_16322,N_14425,N_11654);
nor U16323 (N_16323,N_13851,N_10577);
nor U16324 (N_16324,N_14983,N_11442);
and U16325 (N_16325,N_12133,N_12101);
nand U16326 (N_16326,N_13944,N_13965);
xnor U16327 (N_16327,N_12174,N_12483);
and U16328 (N_16328,N_11082,N_14257);
or U16329 (N_16329,N_10381,N_13272);
xnor U16330 (N_16330,N_13202,N_12683);
xnor U16331 (N_16331,N_12050,N_10506);
and U16332 (N_16332,N_14361,N_10291);
nand U16333 (N_16333,N_12166,N_13672);
and U16334 (N_16334,N_13112,N_11307);
nand U16335 (N_16335,N_12034,N_11327);
and U16336 (N_16336,N_12150,N_11035);
or U16337 (N_16337,N_11557,N_10660);
nor U16338 (N_16338,N_12044,N_14276);
nand U16339 (N_16339,N_10110,N_10038);
or U16340 (N_16340,N_11746,N_12138);
or U16341 (N_16341,N_11569,N_14570);
or U16342 (N_16342,N_14920,N_11847);
nand U16343 (N_16343,N_12387,N_14336);
nor U16344 (N_16344,N_13948,N_14859);
nor U16345 (N_16345,N_11259,N_13872);
or U16346 (N_16346,N_12560,N_10567);
nor U16347 (N_16347,N_10644,N_13797);
and U16348 (N_16348,N_11414,N_14966);
nand U16349 (N_16349,N_10390,N_13796);
nand U16350 (N_16350,N_13163,N_12141);
and U16351 (N_16351,N_11161,N_14762);
nand U16352 (N_16352,N_10933,N_11864);
and U16353 (N_16353,N_12799,N_10416);
nor U16354 (N_16354,N_12601,N_13286);
nand U16355 (N_16355,N_13080,N_14391);
and U16356 (N_16356,N_13679,N_12796);
or U16357 (N_16357,N_10143,N_13700);
or U16358 (N_16358,N_12173,N_10383);
nand U16359 (N_16359,N_13036,N_10327);
or U16360 (N_16360,N_14360,N_11754);
xor U16361 (N_16361,N_14598,N_14724);
xnor U16362 (N_16362,N_13935,N_14255);
nand U16363 (N_16363,N_13162,N_11285);
or U16364 (N_16364,N_13021,N_14671);
nor U16365 (N_16365,N_13507,N_12104);
or U16366 (N_16366,N_14183,N_10901);
xor U16367 (N_16367,N_10218,N_14287);
and U16368 (N_16368,N_10598,N_11942);
nand U16369 (N_16369,N_13107,N_13574);
or U16370 (N_16370,N_13675,N_11110);
or U16371 (N_16371,N_12757,N_13199);
nand U16372 (N_16372,N_13482,N_14437);
and U16373 (N_16373,N_11696,N_13232);
and U16374 (N_16374,N_13041,N_10648);
and U16375 (N_16375,N_13447,N_14426);
or U16376 (N_16376,N_11932,N_13906);
xor U16377 (N_16377,N_14027,N_10094);
nor U16378 (N_16378,N_10252,N_12980);
or U16379 (N_16379,N_10320,N_11923);
nand U16380 (N_16380,N_12259,N_13385);
nand U16381 (N_16381,N_12103,N_14690);
nor U16382 (N_16382,N_14286,N_10059);
or U16383 (N_16383,N_13079,N_11422);
nor U16384 (N_16384,N_11366,N_10679);
nor U16385 (N_16385,N_10620,N_14867);
and U16386 (N_16386,N_11577,N_11881);
or U16387 (N_16387,N_13074,N_13869);
nor U16388 (N_16388,N_12178,N_14423);
or U16389 (N_16389,N_14457,N_13933);
and U16390 (N_16390,N_10603,N_10527);
or U16391 (N_16391,N_13721,N_13443);
nor U16392 (N_16392,N_12602,N_14517);
and U16393 (N_16393,N_14092,N_10680);
nor U16394 (N_16394,N_14193,N_10029);
nor U16395 (N_16395,N_11986,N_10340);
xnor U16396 (N_16396,N_11985,N_14022);
nand U16397 (N_16397,N_12238,N_13733);
nor U16398 (N_16398,N_10292,N_14739);
nand U16399 (N_16399,N_11215,N_12955);
or U16400 (N_16400,N_14237,N_13050);
or U16401 (N_16401,N_11095,N_13290);
nand U16402 (N_16402,N_12379,N_11358);
nor U16403 (N_16403,N_10361,N_11140);
or U16404 (N_16404,N_14047,N_12773);
nor U16405 (N_16405,N_14825,N_11502);
xor U16406 (N_16406,N_14656,N_10797);
or U16407 (N_16407,N_13681,N_12041);
or U16408 (N_16408,N_13214,N_11338);
or U16409 (N_16409,N_14303,N_13135);
and U16410 (N_16410,N_12134,N_14820);
nor U16411 (N_16411,N_14622,N_13637);
or U16412 (N_16412,N_12800,N_10100);
xor U16413 (N_16413,N_10794,N_10692);
nand U16414 (N_16414,N_13244,N_12925);
and U16415 (N_16415,N_11202,N_10872);
nor U16416 (N_16416,N_12119,N_11270);
and U16417 (N_16417,N_13394,N_10818);
and U16418 (N_16418,N_10686,N_11875);
nor U16419 (N_16419,N_14040,N_10019);
nand U16420 (N_16420,N_14452,N_13653);
nand U16421 (N_16421,N_14513,N_11625);
and U16422 (N_16422,N_13924,N_13534);
nand U16423 (N_16423,N_10659,N_10808);
or U16424 (N_16424,N_12089,N_13357);
nor U16425 (N_16425,N_11201,N_12311);
or U16426 (N_16426,N_10614,N_14066);
and U16427 (N_16427,N_11335,N_12912);
or U16428 (N_16428,N_14007,N_10299);
nor U16429 (N_16429,N_10239,N_12935);
nor U16430 (N_16430,N_14484,N_12144);
nor U16431 (N_16431,N_10734,N_14011);
and U16432 (N_16432,N_14279,N_13973);
or U16433 (N_16433,N_13744,N_13046);
or U16434 (N_16434,N_11154,N_13583);
and U16435 (N_16435,N_13119,N_14197);
xor U16436 (N_16436,N_14502,N_13379);
nor U16437 (N_16437,N_10636,N_10991);
xnor U16438 (N_16438,N_10090,N_13010);
nand U16439 (N_16439,N_14326,N_12271);
nor U16440 (N_16440,N_11852,N_12233);
xnor U16441 (N_16441,N_13219,N_13096);
and U16442 (N_16442,N_12477,N_14507);
nand U16443 (N_16443,N_11861,N_13508);
and U16444 (N_16444,N_14020,N_14240);
xnor U16445 (N_16445,N_13060,N_10666);
or U16446 (N_16446,N_13677,N_13344);
nand U16447 (N_16447,N_12558,N_10473);
xnor U16448 (N_16448,N_11339,N_12744);
nand U16449 (N_16449,N_13314,N_10868);
nor U16450 (N_16450,N_10204,N_13687);
nor U16451 (N_16451,N_14220,N_12791);
or U16452 (N_16452,N_13765,N_11507);
nor U16453 (N_16453,N_13978,N_12242);
or U16454 (N_16454,N_14901,N_13591);
and U16455 (N_16455,N_10556,N_10684);
nor U16456 (N_16456,N_12848,N_10873);
and U16457 (N_16457,N_13614,N_14527);
and U16458 (N_16458,N_13650,N_14394);
and U16459 (N_16459,N_13928,N_13723);
nand U16460 (N_16460,N_14510,N_12194);
nor U16461 (N_16461,N_12615,N_12635);
nor U16462 (N_16462,N_11681,N_10723);
or U16463 (N_16463,N_11970,N_14453);
or U16464 (N_16464,N_13436,N_13945);
nand U16465 (N_16465,N_10758,N_12668);
nor U16466 (N_16466,N_12232,N_12212);
or U16467 (N_16467,N_13139,N_12513);
nor U16468 (N_16468,N_11185,N_13345);
nand U16469 (N_16469,N_13982,N_14230);
xnor U16470 (N_16470,N_12466,N_12285);
nor U16471 (N_16471,N_10824,N_11472);
nor U16472 (N_16472,N_12992,N_14875);
nand U16473 (N_16473,N_11496,N_11733);
xnor U16474 (N_16474,N_11211,N_12394);
or U16475 (N_16475,N_13818,N_14182);
nand U16476 (N_16476,N_10548,N_11832);
or U16477 (N_16477,N_14083,N_12640);
or U16478 (N_16478,N_14074,N_14905);
nand U16479 (N_16479,N_11133,N_10343);
nor U16480 (N_16480,N_11457,N_12713);
nor U16481 (N_16481,N_10673,N_11273);
or U16482 (N_16482,N_12062,N_13969);
and U16483 (N_16483,N_10266,N_10147);
xor U16484 (N_16484,N_12054,N_12746);
or U16485 (N_16485,N_12960,N_14185);
xor U16486 (N_16486,N_12281,N_13204);
and U16487 (N_16487,N_12866,N_11978);
nand U16488 (N_16488,N_11551,N_12631);
nand U16489 (N_16489,N_12556,N_10753);
nand U16490 (N_16490,N_13557,N_10534);
nor U16491 (N_16491,N_12382,N_13001);
nor U16492 (N_16492,N_10866,N_13866);
or U16493 (N_16493,N_11514,N_14548);
nor U16494 (N_16494,N_12046,N_12373);
nor U16495 (N_16495,N_10431,N_11177);
nor U16496 (N_16496,N_14476,N_12484);
or U16497 (N_16497,N_14769,N_11143);
and U16498 (N_16498,N_13753,N_12083);
nor U16499 (N_16499,N_10807,N_14304);
or U16500 (N_16500,N_13173,N_14917);
and U16501 (N_16501,N_12909,N_11345);
and U16502 (N_16502,N_10205,N_12549);
nor U16503 (N_16503,N_12290,N_11750);
nand U16504 (N_16504,N_10599,N_12774);
or U16505 (N_16505,N_12765,N_11509);
nor U16506 (N_16506,N_10109,N_10580);
and U16507 (N_16507,N_14687,N_12797);
nor U16508 (N_16508,N_12923,N_12024);
or U16509 (N_16509,N_14105,N_13910);
xor U16510 (N_16510,N_13053,N_13281);
nand U16511 (N_16511,N_10814,N_11516);
and U16512 (N_16512,N_11924,N_13476);
and U16513 (N_16513,N_14719,N_14127);
and U16514 (N_16514,N_11085,N_12779);
and U16515 (N_16515,N_14352,N_11701);
xnor U16516 (N_16516,N_14381,N_10220);
xor U16517 (N_16517,N_11679,N_10762);
nand U16518 (N_16518,N_13955,N_10595);
nor U16519 (N_16519,N_13883,N_12825);
and U16520 (N_16520,N_12446,N_10187);
and U16521 (N_16521,N_13387,N_13843);
or U16522 (N_16522,N_11309,N_10852);
and U16523 (N_16523,N_11941,N_14784);
and U16524 (N_16524,N_10384,N_13071);
nor U16525 (N_16525,N_11118,N_14125);
and U16526 (N_16526,N_11524,N_14771);
xor U16527 (N_16527,N_11671,N_12371);
and U16528 (N_16528,N_14141,N_13894);
or U16529 (N_16529,N_11370,N_12858);
nand U16530 (N_16530,N_13827,N_11816);
nor U16531 (N_16531,N_13318,N_10350);
or U16532 (N_16532,N_11541,N_12639);
xor U16533 (N_16533,N_11979,N_14385);
or U16534 (N_16534,N_14442,N_11169);
and U16535 (N_16535,N_14138,N_13320);
nor U16536 (N_16536,N_12838,N_12002);
nor U16537 (N_16537,N_10300,N_14647);
and U16538 (N_16538,N_13834,N_14233);
nand U16539 (N_16539,N_13812,N_10222);
and U16540 (N_16540,N_13430,N_14465);
or U16541 (N_16541,N_14888,N_13623);
nor U16542 (N_16542,N_14405,N_12981);
nand U16543 (N_16543,N_12183,N_12060);
or U16544 (N_16544,N_14738,N_12898);
xor U16545 (N_16545,N_11543,N_11453);
and U16546 (N_16546,N_13540,N_14349);
nand U16547 (N_16547,N_14063,N_14188);
or U16548 (N_16548,N_13506,N_11998);
nor U16549 (N_16549,N_10705,N_12035);
and U16550 (N_16550,N_13367,N_10531);
nand U16551 (N_16551,N_13779,N_13831);
or U16552 (N_16552,N_11420,N_12627);
nor U16553 (N_16553,N_10386,N_10428);
and U16554 (N_16554,N_10571,N_12574);
and U16555 (N_16555,N_12282,N_14854);
and U16556 (N_16556,N_12260,N_11561);
or U16557 (N_16557,N_10089,N_10564);
nand U16558 (N_16558,N_10650,N_14271);
nor U16559 (N_16559,N_10072,N_14399);
nand U16560 (N_16560,N_10507,N_14396);
nor U16561 (N_16561,N_11562,N_11182);
or U16562 (N_16562,N_13743,N_10073);
nor U16563 (N_16563,N_11157,N_11578);
and U16564 (N_16564,N_11815,N_12108);
and U16565 (N_16565,N_12959,N_10836);
nand U16566 (N_16566,N_12662,N_10877);
or U16567 (N_16567,N_11321,N_10270);
nand U16568 (N_16568,N_13756,N_12456);
nand U16569 (N_16569,N_10450,N_12176);
or U16570 (N_16570,N_13810,N_11408);
and U16571 (N_16571,N_14298,N_12741);
nor U16572 (N_16572,N_12145,N_13452);
nor U16573 (N_16573,N_14824,N_13635);
or U16574 (N_16574,N_12013,N_12872);
xor U16575 (N_16575,N_12630,N_12079);
nand U16576 (N_16576,N_14166,N_11708);
or U16577 (N_16577,N_10845,N_14416);
or U16578 (N_16578,N_12246,N_14329);
or U16579 (N_16579,N_12428,N_12175);
nand U16580 (N_16580,N_11279,N_11120);
or U16581 (N_16581,N_12272,N_13759);
or U16582 (N_16582,N_14661,N_11234);
xnor U16583 (N_16583,N_11659,N_12840);
nor U16584 (N_16584,N_11439,N_10126);
nand U16585 (N_16585,N_12426,N_10865);
and U16586 (N_16586,N_14415,N_11836);
or U16587 (N_16587,N_14946,N_13705);
and U16588 (N_16588,N_12471,N_10135);
xnor U16589 (N_16589,N_11931,N_10915);
nor U16590 (N_16590,N_11029,N_12407);
and U16591 (N_16591,N_13867,N_12289);
nand U16592 (N_16592,N_10198,N_13138);
nor U16593 (N_16593,N_10687,N_11384);
nor U16594 (N_16594,N_13921,N_12015);
nand U16595 (N_16595,N_10562,N_14734);
or U16596 (N_16596,N_11988,N_12663);
or U16597 (N_16597,N_12827,N_14670);
or U16598 (N_16598,N_11982,N_12781);
nand U16599 (N_16599,N_10557,N_13254);
and U16600 (N_16600,N_13325,N_12021);
nand U16601 (N_16601,N_10016,N_13661);
xor U16602 (N_16602,N_11435,N_11081);
or U16603 (N_16603,N_13151,N_10074);
or U16604 (N_16604,N_13303,N_10316);
nand U16605 (N_16605,N_12667,N_12265);
nand U16606 (N_16606,N_11724,N_13825);
xnor U16607 (N_16607,N_13407,N_13390);
nor U16608 (N_16608,N_11878,N_13553);
nand U16609 (N_16609,N_14890,N_14579);
and U16610 (N_16610,N_11168,N_10255);
or U16611 (N_16611,N_10057,N_11762);
nand U16612 (N_16612,N_12578,N_13655);
and U16613 (N_16613,N_12932,N_11596);
and U16614 (N_16614,N_14954,N_13306);
and U16615 (N_16615,N_11786,N_13266);
or U16616 (N_16616,N_10476,N_10293);
and U16617 (N_16617,N_13940,N_14492);
and U16618 (N_16618,N_10893,N_12085);
nand U16619 (N_16619,N_10894,N_14959);
and U16620 (N_16620,N_10236,N_10542);
xor U16621 (N_16621,N_11850,N_10304);
and U16622 (N_16622,N_13880,N_11683);
nor U16623 (N_16623,N_12951,N_11780);
or U16624 (N_16624,N_12294,N_13528);
and U16625 (N_16625,N_14469,N_13674);
nor U16626 (N_16626,N_11084,N_13458);
nor U16627 (N_16627,N_12976,N_13279);
xnor U16628 (N_16628,N_12442,N_10669);
or U16629 (N_16629,N_10104,N_10550);
nand U16630 (N_16630,N_10565,N_10536);
nor U16631 (N_16631,N_14973,N_10788);
nand U16632 (N_16632,N_10373,N_13569);
and U16633 (N_16633,N_14681,N_14775);
nand U16634 (N_16634,N_13846,N_14014);
nor U16635 (N_16635,N_10184,N_12425);
nand U16636 (N_16636,N_13415,N_11773);
or U16637 (N_16637,N_11010,N_10071);
and U16638 (N_16638,N_13373,N_12534);
nand U16639 (N_16639,N_13355,N_10129);
or U16640 (N_16640,N_13061,N_14774);
and U16641 (N_16641,N_14953,N_10616);
or U16642 (N_16642,N_10217,N_12768);
nand U16643 (N_16643,N_10001,N_12512);
nand U16644 (N_16644,N_13898,N_12587);
and U16645 (N_16645,N_12928,N_13800);
or U16646 (N_16646,N_13356,N_13187);
nand U16647 (N_16647,N_11200,N_10241);
or U16648 (N_16648,N_12077,N_10351);
and U16649 (N_16649,N_13701,N_12533);
nor U16650 (N_16650,N_13904,N_11977);
xnor U16651 (N_16651,N_12217,N_14033);
and U16652 (N_16652,N_12244,N_12361);
nor U16653 (N_16653,N_10201,N_11074);
or U16654 (N_16654,N_14057,N_14872);
or U16655 (N_16655,N_13839,N_14573);
and U16656 (N_16656,N_12828,N_11947);
nand U16657 (N_16657,N_12826,N_13195);
and U16658 (N_16658,N_13024,N_10199);
nand U16659 (N_16659,N_10464,N_10930);
or U16660 (N_16660,N_10954,N_14864);
or U16661 (N_16661,N_14281,N_14620);
or U16662 (N_16662,N_10820,N_10176);
nand U16663 (N_16663,N_12404,N_10216);
or U16664 (N_16664,N_10655,N_12626);
nor U16665 (N_16665,N_12078,N_11281);
or U16666 (N_16666,N_13137,N_13885);
nor U16667 (N_16667,N_12424,N_14541);
or U16668 (N_16668,N_13641,N_10922);
xor U16669 (N_16669,N_10372,N_14787);
or U16670 (N_16670,N_11412,N_11720);
nor U16671 (N_16671,N_11187,N_13134);
and U16672 (N_16672,N_11501,N_14036);
nor U16673 (N_16673,N_14981,N_14283);
nand U16674 (N_16674,N_12172,N_14539);
and U16675 (N_16675,N_12759,N_11767);
nor U16676 (N_16676,N_14699,N_13500);
nand U16677 (N_16677,N_10510,N_12296);
xor U16678 (N_16678,N_11471,N_11101);
nor U16679 (N_16679,N_12467,N_13714);
nor U16680 (N_16680,N_11571,N_13020);
or U16681 (N_16681,N_11897,N_11695);
xor U16682 (N_16682,N_14207,N_10459);
and U16683 (N_16683,N_14806,N_10804);
and U16684 (N_16684,N_14117,N_10795);
nor U16685 (N_16685,N_14489,N_12656);
nand U16686 (N_16686,N_14848,N_13375);
nand U16687 (N_16687,N_11765,N_11038);
nor U16688 (N_16688,N_13222,N_14393);
nand U16689 (N_16689,N_13300,N_12069);
nand U16690 (N_16690,N_12669,N_13460);
nor U16691 (N_16691,N_14878,N_13432);
xnor U16692 (N_16692,N_11461,N_12254);
or U16693 (N_16693,N_10261,N_14772);
or U16694 (N_16694,N_14308,N_11254);
nand U16695 (N_16695,N_12634,N_12751);
or U16696 (N_16696,N_12017,N_14768);
nand U16697 (N_16697,N_14988,N_14940);
nand U16698 (N_16698,N_12857,N_14152);
or U16699 (N_16699,N_11568,N_14162);
nand U16700 (N_16700,N_14319,N_12885);
nand U16701 (N_16701,N_11796,N_14642);
and U16702 (N_16702,N_14882,N_13555);
or U16703 (N_16703,N_13386,N_12263);
and U16704 (N_16704,N_11226,N_11717);
nand U16705 (N_16705,N_11804,N_10061);
or U16706 (N_16706,N_13657,N_13995);
nor U16707 (N_16707,N_14980,N_11840);
or U16708 (N_16708,N_13478,N_13147);
xor U16709 (N_16709,N_10329,N_13295);
and U16710 (N_16710,N_12723,N_13130);
or U16711 (N_16711,N_11141,N_13870);
and U16712 (N_16712,N_11076,N_14114);
or U16713 (N_16713,N_13451,N_14798);
nor U16714 (N_16714,N_11871,N_14816);
or U16715 (N_16715,N_10033,N_14291);
or U16716 (N_16716,N_11036,N_10330);
nor U16717 (N_16717,N_11265,N_12508);
nor U16718 (N_16718,N_11167,N_12539);
xnor U16719 (N_16719,N_14991,N_10790);
or U16720 (N_16720,N_14740,N_14518);
nand U16721 (N_16721,N_10004,N_14080);
nor U16722 (N_16722,N_14604,N_14149);
nor U16723 (N_16723,N_12495,N_11040);
and U16724 (N_16724,N_10526,N_13932);
nor U16725 (N_16725,N_11838,N_10056);
or U16726 (N_16726,N_13418,N_13065);
and U16727 (N_16727,N_12767,N_10417);
or U16728 (N_16728,N_10558,N_14151);
nor U16729 (N_16729,N_11782,N_11635);
nor U16730 (N_16730,N_11057,N_12896);
or U16731 (N_16731,N_11853,N_12650);
nand U16732 (N_16732,N_14949,N_11272);
nand U16733 (N_16733,N_13054,N_14184);
and U16734 (N_16734,N_13011,N_10649);
xnor U16735 (N_16735,N_11715,N_14943);
xnor U16736 (N_16736,N_13369,N_12480);
or U16737 (N_16737,N_14755,N_13908);
nor U16738 (N_16738,N_10495,N_12247);
nor U16739 (N_16739,N_10642,N_10344);
nand U16740 (N_16740,N_11612,N_12862);
and U16741 (N_16741,N_12965,N_14691);
or U16742 (N_16742,N_13413,N_11411);
or U16743 (N_16743,N_11512,N_14652);
or U16744 (N_16744,N_14205,N_12834);
nand U16745 (N_16745,N_14664,N_12280);
nand U16746 (N_16746,N_13871,N_13612);
and U16747 (N_16747,N_12324,N_13141);
xor U16748 (N_16748,N_14324,N_10766);
nand U16749 (N_16749,N_11805,N_14689);
nand U16750 (N_16750,N_12431,N_11585);
or U16751 (N_16751,N_11021,N_14320);
nand U16752 (N_16752,N_13873,N_12208);
and U16753 (N_16753,N_11650,N_10174);
nor U16754 (N_16754,N_12632,N_10262);
nand U16755 (N_16755,N_14199,N_14447);
xor U16756 (N_16756,N_11222,N_13275);
nand U16757 (N_16757,N_10538,N_11952);
and U16758 (N_16758,N_11657,N_14728);
xor U16759 (N_16759,N_10832,N_12537);
xor U16760 (N_16760,N_11326,N_10725);
nor U16761 (N_16761,N_12349,N_13699);
nand U16762 (N_16762,N_11460,N_12641);
nor U16763 (N_16763,N_10257,N_14462);
nor U16764 (N_16764,N_14568,N_12074);
or U16765 (N_16765,N_11116,N_11573);
xnor U16766 (N_16766,N_11334,N_12576);
nand U16767 (N_16767,N_11075,N_11220);
or U16768 (N_16768,N_11436,N_11546);
and U16769 (N_16769,N_12327,N_14850);
or U16770 (N_16770,N_13248,N_12163);
nor U16771 (N_16771,N_12878,N_13620);
xnor U16772 (N_16772,N_11889,N_10133);
or U16773 (N_16773,N_10876,N_12874);
xnor U16774 (N_16774,N_14401,N_13362);
and U16775 (N_16775,N_13383,N_14203);
and U16776 (N_16776,N_14814,N_13817);
nand U16777 (N_16777,N_11099,N_14274);
xnor U16778 (N_16778,N_14245,N_11172);
and U16779 (N_16779,N_14729,N_13752);
nor U16780 (N_16780,N_12120,N_11630);
and U16781 (N_16781,N_10964,N_10368);
xor U16782 (N_16782,N_12514,N_10145);
nand U16783 (N_16783,N_14157,N_11368);
or U16784 (N_16784,N_14246,N_11437);
or U16785 (N_16785,N_12749,N_14186);
nor U16786 (N_16786,N_11373,N_14427);
or U16787 (N_16787,N_14667,N_13582);
and U16788 (N_16788,N_10458,N_10741);
or U16789 (N_16789,N_13361,N_11070);
nor U16790 (N_16790,N_10809,N_14119);
nor U16791 (N_16791,N_12545,N_10339);
or U16792 (N_16792,N_10449,N_13441);
or U16793 (N_16793,N_13902,N_13364);
or U16794 (N_16794,N_14684,N_12585);
xnor U16795 (N_16795,N_12895,N_11351);
nand U16796 (N_16796,N_13063,N_10667);
and U16797 (N_16797,N_11972,N_11045);
nor U16798 (N_16798,N_13990,N_12225);
nor U16799 (N_16799,N_13757,N_14531);
and U16800 (N_16800,N_14212,N_14129);
and U16801 (N_16801,N_13013,N_12820);
or U16802 (N_16802,N_12798,N_12709);
and U16803 (N_16803,N_12027,N_11130);
nor U16804 (N_16804,N_14958,N_11618);
nor U16805 (N_16805,N_14338,N_11049);
xor U16806 (N_16806,N_12947,N_11934);
xor U16807 (N_16807,N_11424,N_12764);
nand U16808 (N_16808,N_11403,N_13115);
xnor U16809 (N_16809,N_10423,N_10028);
and U16810 (N_16810,N_10268,N_10639);
and U16811 (N_16811,N_10058,N_11983);
xor U16812 (N_16812,N_10888,N_10503);
and U16813 (N_16813,N_12412,N_14150);
nand U16814 (N_16814,N_12030,N_11230);
nand U16815 (N_16815,N_13338,N_11854);
and U16816 (N_16816,N_14797,N_11731);
nor U16817 (N_16817,N_13968,N_14588);
or U16818 (N_16818,N_11150,N_13896);
nand U16819 (N_16819,N_12187,N_11324);
nand U16820 (N_16820,N_14058,N_14904);
xnor U16821 (N_16821,N_13710,N_14581);
and U16822 (N_16822,N_11004,N_12472);
xnor U16823 (N_16823,N_12256,N_11752);
or U16824 (N_16824,N_11911,N_12913);
or U16825 (N_16825,N_11349,N_12308);
nand U16826 (N_16826,N_12257,N_11102);
nor U16827 (N_16827,N_11432,N_12397);
xor U16828 (N_16828,N_14702,N_12961);
nor U16829 (N_16829,N_12869,N_14204);
nand U16830 (N_16830,N_10729,N_11519);
or U16831 (N_16831,N_12231,N_13654);
nand U16832 (N_16832,N_14313,N_11062);
nand U16833 (N_16833,N_14252,N_13917);
or U16834 (N_16834,N_12364,N_14147);
nor U16835 (N_16835,N_12065,N_13301);
nor U16836 (N_16836,N_11817,N_12418);
and U16837 (N_16837,N_14536,N_13748);
or U16838 (N_16838,N_14134,N_10755);
xor U16839 (N_16839,N_10919,N_13950);
nor U16840 (N_16840,N_11574,N_10522);
or U16841 (N_16841,N_10652,N_13122);
and U16842 (N_16842,N_12673,N_14130);
or U16843 (N_16843,N_10082,N_14118);
nor U16844 (N_16844,N_10774,N_14939);
nor U16845 (N_16845,N_13378,N_13183);
nand U16846 (N_16846,N_10470,N_13783);
nor U16847 (N_16847,N_11922,N_10627);
or U16848 (N_16848,N_12703,N_14560);
and U16849 (N_16849,N_11073,N_14998);
and U16850 (N_16850,N_14214,N_13496);
and U16851 (N_16851,N_14490,N_14195);
and U16852 (N_16852,N_13521,N_11100);
xor U16853 (N_16853,N_14019,N_12273);
nand U16854 (N_16854,N_11315,N_10382);
nor U16855 (N_16855,N_14155,N_10746);
or U16856 (N_16856,N_10101,N_12968);
or U16857 (N_16857,N_10516,N_11165);
nand U16858 (N_16858,N_11522,N_13830);
or U16859 (N_16859,N_12121,N_14669);
nor U16860 (N_16860,N_11709,N_13076);
and U16861 (N_16861,N_10704,N_12986);
and U16862 (N_16862,N_10645,N_13853);
nand U16863 (N_16863,N_10874,N_13003);
nand U16864 (N_16864,N_12894,N_12982);
or U16865 (N_16865,N_10626,N_13835);
nor U16866 (N_16866,N_11078,N_11083);
nor U16867 (N_16867,N_10857,N_12929);
xor U16868 (N_16868,N_14840,N_10347);
or U16869 (N_16869,N_13959,N_12253);
nand U16870 (N_16870,N_13980,N_14480);
or U16871 (N_16871,N_12674,N_12350);
nor U16872 (N_16872,N_14742,N_12732);
and U16873 (N_16873,N_12738,N_11686);
nand U16874 (N_16874,N_11142,N_14089);
and U16875 (N_16875,N_14565,N_10349);
or U16876 (N_16876,N_12064,N_13312);
and U16877 (N_16877,N_12941,N_12510);
nor U16878 (N_16878,N_10905,N_12469);
xnor U16879 (N_16879,N_10588,N_12197);
xnor U16880 (N_16880,N_13838,N_13179);
nor U16881 (N_16881,N_11290,N_13760);
nand U16882 (N_16882,N_11098,N_13716);
nor U16883 (N_16883,N_14530,N_11328);
nor U16884 (N_16884,N_10849,N_13401);
xnor U16885 (N_16885,N_11553,N_11510);
or U16886 (N_16886,N_12267,N_10902);
and U16887 (N_16887,N_12762,N_12320);
nand U16888 (N_16888,N_10972,N_11257);
nor U16889 (N_16889,N_14701,N_10525);
nand U16890 (N_16890,N_13140,N_10267);
xor U16891 (N_16891,N_11615,N_13255);
or U16892 (N_16892,N_10579,N_11806);
and U16893 (N_16893,N_12328,N_11094);
and U16894 (N_16894,N_12954,N_11984);
and U16895 (N_16895,N_14819,N_14432);
xnor U16896 (N_16896,N_13882,N_12307);
and U16897 (N_16897,N_13522,N_13719);
or U16898 (N_16898,N_11431,N_11064);
or U16899 (N_16899,N_12177,N_14613);
nor U16900 (N_16900,N_10843,N_14813);
and U16901 (N_16901,N_10898,N_11728);
nor U16902 (N_16902,N_12189,N_12890);
nand U16903 (N_16903,N_14419,N_14071);
and U16904 (N_16904,N_13166,N_14334);
xnor U16905 (N_16905,N_13235,N_11608);
or U16906 (N_16906,N_10043,N_13051);
and U16907 (N_16907,N_12694,N_13196);
nand U16908 (N_16908,N_13717,N_14501);
nor U16909 (N_16909,N_14826,N_13564);
xnor U16910 (N_16910,N_11814,N_11685);
nor U16911 (N_16911,N_14384,N_11857);
or U16912 (N_16912,N_11739,N_12362);
xor U16913 (N_16913,N_11477,N_14101);
nor U16914 (N_16914,N_10635,N_11700);
and U16915 (N_16915,N_13193,N_13890);
xnor U16916 (N_16916,N_12771,N_11015);
nor U16917 (N_16917,N_12742,N_11647);
and U16918 (N_16918,N_14619,N_14165);
or U16919 (N_16919,N_12159,N_12726);
xor U16920 (N_16920,N_13342,N_12262);
or U16921 (N_16921,N_10928,N_14109);
nor U16922 (N_16922,N_14451,N_13495);
and U16923 (N_16923,N_13278,N_14408);
nand U16924 (N_16924,N_13997,N_13128);
or U16925 (N_16925,N_10539,N_12264);
nor U16926 (N_16926,N_14842,N_13832);
nor U16927 (N_16927,N_10309,N_10641);
nor U16928 (N_16928,N_10412,N_10009);
or U16929 (N_16929,N_10461,N_12944);
nand U16930 (N_16930,N_10596,N_11209);
nand U16931 (N_16931,N_14688,N_13461);
and U16932 (N_16932,N_13547,N_13186);
nor U16933 (N_16933,N_14837,N_10319);
nand U16934 (N_16934,N_14685,N_11946);
nor U16935 (N_16935,N_10955,N_14512);
nor U16936 (N_16936,N_12506,N_11809);
or U16937 (N_16937,N_13698,N_10488);
nor U16938 (N_16938,N_14024,N_10203);
or U16939 (N_16939,N_13791,N_13805);
nand U16940 (N_16940,N_13127,N_13624);
and U16941 (N_16941,N_12867,N_10566);
nor U16942 (N_16942,N_12366,N_14348);
or U16943 (N_16943,N_11033,N_13472);
xor U16944 (N_16944,N_10286,N_11869);
or U16945 (N_16945,N_12380,N_13876);
nand U16946 (N_16946,N_11807,N_14572);
xnor U16947 (N_16947,N_13333,N_11221);
or U16948 (N_16948,N_10830,N_10159);
nand U16949 (N_16949,N_12492,N_14061);
nand U16950 (N_16950,N_12113,N_10973);
nor U16951 (N_16951,N_13448,N_11621);
nor U16952 (N_16952,N_11065,N_12427);
xnor U16953 (N_16953,N_11119,N_14002);
nor U16954 (N_16954,N_13718,N_13984);
nor U16955 (N_16955,N_11275,N_10256);
nand U16956 (N_16956,N_10166,N_14030);
nor U16957 (N_16957,N_12389,N_14458);
nand U16958 (N_16958,N_10971,N_10010);
and U16959 (N_16959,N_12831,N_13532);
nor U16960 (N_16960,N_12972,N_14096);
nand U16961 (N_16961,N_14116,N_11296);
nor U16962 (N_16962,N_10044,N_13727);
nand U16963 (N_16963,N_12109,N_11710);
nand U16964 (N_16964,N_13018,N_10260);
nor U16965 (N_16965,N_14407,N_10590);
nor U16966 (N_16966,N_13979,N_14493);
and U16967 (N_16967,N_12837,N_12967);
nand U16968 (N_16968,N_14373,N_10740);
or U16969 (N_16969,N_14430,N_13595);
xnor U16970 (N_16970,N_11216,N_12441);
nand U16971 (N_16971,N_12312,N_14752);
xor U16972 (N_16972,N_11735,N_11611);
or U16973 (N_16973,N_14733,N_14413);
and U16974 (N_16974,N_14569,N_10619);
nor U16975 (N_16975,N_11044,N_10767);
and U16976 (N_16976,N_14031,N_13833);
and U16977 (N_16977,N_10466,N_10244);
nand U16978 (N_16978,N_13148,N_14288);
xor U16979 (N_16979,N_13059,N_13958);
nor U16980 (N_16980,N_13465,N_10138);
and U16981 (N_16981,N_11759,N_13487);
nand U16982 (N_16982,N_10250,N_14295);
nand U16983 (N_16983,N_13686,N_12745);
nor U16984 (N_16984,N_13941,N_13793);
or U16985 (N_16985,N_14678,N_10317);
nor U16986 (N_16986,N_10552,N_13600);
nor U16987 (N_16987,N_13842,N_13596);
nor U16988 (N_16988,N_11124,N_11147);
nor U16989 (N_16989,N_14876,N_10946);
nor U16990 (N_16990,N_10956,N_10720);
and U16991 (N_16991,N_10618,N_11566);
xor U16992 (N_16992,N_12416,N_13977);
xor U16993 (N_16993,N_11537,N_14509);
xnor U16994 (N_16994,N_12702,N_14597);
and U16995 (N_16995,N_10601,N_11176);
nand U16996 (N_16996,N_13695,N_13828);
nor U16997 (N_16997,N_11534,N_14659);
or U16998 (N_16998,N_11337,N_14253);
nor U16999 (N_16999,N_10879,N_11768);
xor U17000 (N_17000,N_13498,N_14250);
nor U17001 (N_17001,N_14640,N_14720);
nand U17002 (N_17002,N_13963,N_13058);
nor U17003 (N_17003,N_14414,N_12292);
or U17004 (N_17004,N_14260,N_12468);
or U17005 (N_17005,N_12170,N_13250);
nand U17006 (N_17006,N_14654,N_11195);
nand U17007 (N_17007,N_11620,N_13419);
nor U17008 (N_17008,N_11194,N_10113);
or U17009 (N_17009,N_10021,N_11529);
nand U17010 (N_17010,N_11232,N_10935);
nand U17011 (N_17011,N_14970,N_13692);
nor U17012 (N_17012,N_11385,N_11698);
xor U17013 (N_17013,N_10637,N_10665);
nand U17014 (N_17014,N_13215,N_11500);
xor U17015 (N_17015,N_11323,N_14448);
nand U17016 (N_17016,N_13703,N_12752);
nand U17017 (N_17017,N_11277,N_14311);
and U17018 (N_17018,N_14374,N_11239);
xnor U17019 (N_17019,N_11347,N_11598);
nand U17020 (N_17020,N_10487,N_13617);
nand U17021 (N_17021,N_14811,N_12067);
nor U17022 (N_17022,N_10259,N_14180);
nand U17023 (N_17023,N_12902,N_14763);
nor U17024 (N_17024,N_12106,N_14528);
and U17025 (N_17025,N_13433,N_12105);
or U17026 (N_17026,N_13083,N_12717);
or U17027 (N_17027,N_13730,N_13671);
nor U17028 (N_17028,N_14629,N_13086);
nand U17029 (N_17029,N_12696,N_12038);
and U17030 (N_17030,N_14558,N_11470);
nor U17031 (N_17031,N_11126,N_14144);
or U17032 (N_17032,N_14115,N_12235);
or U17033 (N_17033,N_10283,N_10549);
or U17034 (N_17034,N_11587,N_11391);
nand U17035 (N_17035,N_11313,N_14486);
nor U17036 (N_17036,N_11229,N_14810);
nand U17037 (N_17037,N_14355,N_11716);
nor U17038 (N_17038,N_10498,N_14861);
xnor U17039 (N_17039,N_14576,N_11846);
or U17040 (N_17040,N_11662,N_12061);
or U17041 (N_17041,N_13683,N_12293);
or U17042 (N_17042,N_10715,N_10551);
nand U17043 (N_17043,N_10739,N_10864);
and U17044 (N_17044,N_13771,N_14559);
and U17045 (N_17045,N_11344,N_10397);
or U17046 (N_17046,N_11900,N_14440);
and U17047 (N_17047,N_13526,N_11380);
nor U17048 (N_17048,N_10706,N_14258);
nor U17049 (N_17049,N_14218,N_10335);
and U17050 (N_17050,N_10434,N_13341);
nor U17051 (N_17051,N_12526,N_11845);
nand U17052 (N_17052,N_10791,N_14908);
or U17053 (N_17053,N_10142,N_12420);
xnor U17054 (N_17054,N_13328,N_11894);
or U17055 (N_17055,N_13315,N_13479);
and U17056 (N_17056,N_10130,N_11909);
and U17057 (N_17057,N_11260,N_11173);
nand U17058 (N_17058,N_12059,N_11719);
xor U17059 (N_17059,N_11288,N_10923);
xor U17060 (N_17060,N_12008,N_14346);
nand U17061 (N_17061,N_13091,N_13627);
nor U17062 (N_17062,N_13431,N_11811);
and U17063 (N_17063,N_12763,N_11096);
nand U17064 (N_17064,N_14342,N_11276);
or U17065 (N_17065,N_11158,N_10782);
or U17066 (N_17066,N_10500,N_11538);
or U17067 (N_17067,N_12122,N_11088);
or U17068 (N_17068,N_10784,N_13309);
nor U17069 (N_17069,N_10155,N_12019);
nand U17070 (N_17070,N_11819,N_13090);
or U17071 (N_17071,N_10948,N_12612);
nand U17072 (N_17072,N_11669,N_10521);
xor U17073 (N_17073,N_13048,N_14318);
and U17074 (N_17074,N_12279,N_11917);
nand U17075 (N_17075,N_11515,N_14275);
nor U17076 (N_17076,N_13270,N_11282);
or U17077 (N_17077,N_13340,N_14236);
nor U17078 (N_17078,N_10086,N_14974);
or U17079 (N_17079,N_14347,N_10492);
or U17080 (N_17080,N_11677,N_11233);
xnor U17081 (N_17081,N_11077,N_14866);
xor U17082 (N_17082,N_12129,N_10957);
nor U17083 (N_17083,N_13274,N_10006);
or U17084 (N_17084,N_12337,N_11267);
or U17085 (N_17085,N_11293,N_12808);
nand U17086 (N_17086,N_10065,N_13228);
nor U17087 (N_17087,N_13396,N_12883);
or U17088 (N_17088,N_14969,N_11730);
or U17089 (N_17089,N_12818,N_10640);
nor U17090 (N_17090,N_10067,N_11665);
nand U17091 (N_17091,N_14508,N_11623);
nand U17092 (N_17092,N_10358,N_13993);
or U17093 (N_17093,N_10537,N_10584);
xnor U17094 (N_17094,N_11588,N_10634);
xor U17095 (N_17095,N_12200,N_11639);
nor U17096 (N_17096,N_13688,N_13289);
nand U17097 (N_17097,N_13084,N_14766);
nor U17098 (N_17098,N_10353,N_11792);
or U17099 (N_17099,N_13946,N_13101);
nor U17100 (N_17100,N_13207,N_11043);
and U17101 (N_17101,N_10456,N_11299);
or U17102 (N_17102,N_13445,N_14892);
or U17103 (N_17103,N_12485,N_10441);
or U17104 (N_17104,N_12730,N_11622);
and U17105 (N_17105,N_10515,N_11833);
or U17106 (N_17106,N_13794,N_13212);
nand U17107 (N_17107,N_13740,N_10410);
nor U17108 (N_17108,N_11034,N_11649);
nor U17109 (N_17109,N_14591,N_10322);
nand U17110 (N_17110,N_10647,N_11086);
and U17111 (N_17111,N_11410,N_13697);
nand U17112 (N_17112,N_12131,N_11186);
nor U17113 (N_17113,N_10787,N_12252);
nand U17114 (N_17114,N_10415,N_12018);
or U17115 (N_17115,N_14142,N_13256);
and U17116 (N_17116,N_10093,N_12606);
and U17117 (N_17117,N_10892,N_13585);
nand U17118 (N_17118,N_14428,N_12203);
xnor U17119 (N_17119,N_13015,N_14026);
or U17120 (N_17120,N_11467,N_14221);
and U17121 (N_17121,N_10505,N_14200);
or U17122 (N_17122,N_14456,N_14100);
nor U17123 (N_17123,N_13858,N_14177);
nand U17124 (N_17124,N_11359,N_14903);
nand U17125 (N_17125,N_13607,N_14614);
nand U17126 (N_17126,N_11139,N_13769);
nand U17127 (N_17127,N_11678,N_12491);
nor U17128 (N_17128,N_11498,N_11190);
nor U17129 (N_17129,N_11723,N_12888);
or U17130 (N_17130,N_13960,N_11919);
xor U17131 (N_17131,N_12335,N_13804);
and U17132 (N_17132,N_10240,N_11404);
or U17133 (N_17133,N_13711,N_10047);
nor U17134 (N_17134,N_10748,N_12724);
nor U17135 (N_17135,N_13073,N_14790);
or U17136 (N_17136,N_12210,N_13647);
and U17137 (N_17137,N_14025,N_12114);
or U17138 (N_17138,N_14215,N_12720);
or U17139 (N_17139,N_14171,N_11870);
xnor U17140 (N_17140,N_12690,N_11132);
or U17141 (N_17141,N_12409,N_10995);
or U17142 (N_17142,N_14999,N_14365);
nand U17143 (N_17143,N_12859,N_13913);
and U17144 (N_17144,N_11463,N_12137);
nand U17145 (N_17145,N_12036,N_12437);
and U17146 (N_17146,N_11860,N_11398);
xnor U17147 (N_17147,N_12645,N_11741);
nor U17148 (N_17148,N_14424,N_12657);
nor U17149 (N_17149,N_11386,N_12076);
nor U17150 (N_17150,N_14997,N_14989);
and U17151 (N_17151,N_13749,N_12721);
xnor U17152 (N_17152,N_10751,N_11699);
and U17153 (N_17153,N_10965,N_11067);
or U17154 (N_17154,N_10087,N_11827);
nor U17155 (N_17155,N_12806,N_13181);
and U17156 (N_17156,N_10547,N_14758);
nand U17157 (N_17157,N_11495,N_13673);
nand U17158 (N_17158,N_12123,N_12676);
nand U17159 (N_17159,N_14190,N_14856);
and U17160 (N_17160,N_12029,N_10569);
xor U17161 (N_17161,N_11844,N_10728);
nor U17162 (N_17162,N_13490,N_10277);
nor U17163 (N_17163,N_14272,N_11362);
or U17164 (N_17164,N_10886,N_10242);
xor U17165 (N_17165,N_13720,N_13666);
xor U17166 (N_17166,N_12996,N_10000);
and U17167 (N_17167,N_10141,N_12475);
nand U17168 (N_17168,N_12855,N_10578);
xnor U17169 (N_17169,N_11484,N_12522);
nand U17170 (N_17170,N_10478,N_14082);
xor U17171 (N_17171,N_10041,N_13581);
xnor U17172 (N_17172,N_11354,N_10485);
or U17173 (N_17173,N_11660,N_10783);
xnor U17174 (N_17174,N_13704,N_12699);
nand U17175 (N_17175,N_12688,N_13146);
or U17176 (N_17176,N_11474,N_14877);
nor U17177 (N_17177,N_13442,N_14595);
nand U17178 (N_17178,N_11938,N_12529);
or U17179 (N_17179,N_12536,N_11527);
nand U17180 (N_17180,N_14934,N_12753);
nand U17181 (N_17181,N_13822,N_13562);
or U17182 (N_17182,N_10096,N_13645);
or U17183 (N_17183,N_12168,N_14680);
nor U17184 (N_17184,N_14606,N_11976);
xor U17185 (N_17185,N_10663,N_13022);
nor U17186 (N_17186,N_11444,N_13606);
and U17187 (N_17187,N_13670,N_13755);
nor U17188 (N_17188,N_13332,N_14979);
and U17189 (N_17189,N_11893,N_13561);
nor U17190 (N_17190,N_10497,N_13690);
nor U17191 (N_17191,N_12788,N_13444);
and U17192 (N_17192,N_12933,N_13243);
nor U17193 (N_17193,N_11063,N_13531);
and U17194 (N_17194,N_13925,N_11428);
nor U17195 (N_17195,N_10541,N_12664);
and U17196 (N_17196,N_14070,N_14709);
nor U17197 (N_17197,N_11163,N_14112);
and U17198 (N_17198,N_10163,N_13519);
and U17199 (N_17199,N_14961,N_10700);
nor U17200 (N_17200,N_12849,N_13613);
and U17201 (N_17201,N_12743,N_14780);
nor U17202 (N_17202,N_12608,N_11213);
nand U17203 (N_17203,N_10940,N_11506);
or U17204 (N_17204,N_13188,N_10468);
and U17205 (N_17205,N_14972,N_13786);
nand U17206 (N_17206,N_14046,N_12016);
and U17207 (N_17207,N_14611,N_14964);
nor U17208 (N_17208,N_11492,N_12865);
or U17209 (N_17209,N_14538,N_13815);
or U17210 (N_17210,N_14845,N_13636);
or U17211 (N_17211,N_13037,N_10934);
or U17212 (N_17212,N_14156,N_14554);
or U17213 (N_17213,N_11643,N_12953);
xor U17214 (N_17214,N_10829,N_14064);
nand U17215 (N_17215,N_12971,N_11375);
or U17216 (N_17216,N_10823,N_11415);
nor U17217 (N_17217,N_12520,N_12058);
xnor U17218 (N_17218,N_11570,N_14631);
nor U17219 (N_17219,N_11913,N_11565);
nand U17220 (N_17220,N_13283,N_11682);
and U17221 (N_17221,N_11749,N_13205);
or U17222 (N_17222,N_11964,N_12153);
and U17223 (N_17223,N_10785,N_11610);
nor U17224 (N_17224,N_10858,N_11829);
nand U17225 (N_17225,N_10568,N_14662);
or U17226 (N_17226,N_10996,N_13268);
and U17227 (N_17227,N_13082,N_11475);
or U17228 (N_17228,N_11243,N_10388);
nor U17229 (N_17229,N_13722,N_14351);
nor U17230 (N_17230,N_13158,N_11798);
or U17231 (N_17231,N_10354,N_11794);
nor U17232 (N_17232,N_11093,N_12494);
nor U17233 (N_17233,N_11856,N_12453);
or U17234 (N_17234,N_10691,N_10999);
nand U17235 (N_17235,N_12687,N_13558);
nand U17236 (N_17236,N_13350,N_14330);
and U17237 (N_17237,N_13422,N_14068);
nor U17238 (N_17238,N_12461,N_13552);
nor U17239 (N_17239,N_11933,N_14364);
and U17240 (N_17240,N_14899,N_14556);
xor U17241 (N_17241,N_12829,N_11614);
and U17242 (N_17242,N_10315,N_11799);
or U17243 (N_17243,N_13524,N_12614);
or U17244 (N_17244,N_13709,N_11989);
and U17245 (N_17245,N_11711,N_14067);
and U17246 (N_17246,N_12434,N_14266);
nor U17247 (N_17247,N_13546,N_13002);
nand U17248 (N_17248,N_11784,N_11419);
nand U17249 (N_17249,N_14863,N_13789);
nor U17250 (N_17250,N_12097,N_12977);
xor U17251 (N_17251,N_10285,N_10435);
and U17252 (N_17252,N_13572,N_11926);
nor U17253 (N_17253,N_12636,N_11781);
nor U17254 (N_17254,N_10108,N_13680);
and U17255 (N_17255,N_12665,N_13165);
nand U17256 (N_17256,N_12419,N_10771);
or U17257 (N_17257,N_10479,N_13539);
and U17258 (N_17258,N_10511,N_12402);
nand U17259 (N_17259,N_13423,N_10111);
or U17260 (N_17260,N_14060,N_13097);
nand U17261 (N_17261,N_11969,N_14120);
xor U17262 (N_17262,N_13847,N_12317);
and U17263 (N_17263,N_14839,N_10246);
nand U17264 (N_17264,N_13916,N_14357);
xnor U17265 (N_17265,N_10846,N_11954);
nor U17266 (N_17266,N_14532,N_11640);
xor U17267 (N_17267,N_14898,N_11016);
nand U17268 (N_17268,N_11997,N_10615);
nand U17269 (N_17269,N_10697,N_13334);
nand U17270 (N_17270,N_12451,N_10518);
nor U17271 (N_17271,N_11666,N_12877);
and U17272 (N_17272,N_12057,N_10831);
nor U17273 (N_17273,N_14473,N_13708);
xor U17274 (N_17274,N_12747,N_11191);
xor U17275 (N_17275,N_13792,N_11694);
nor U17276 (N_17276,N_10481,N_12755);
or U17277 (N_17277,N_12647,N_11747);
or U17278 (N_17278,N_11564,N_13527);
and U17279 (N_17279,N_10195,N_12340);
or U17280 (N_17280,N_13008,N_14099);
xnor U17281 (N_17281,N_13587,N_14006);
xnor U17282 (N_17282,N_12031,N_14041);
or U17283 (N_17283,N_11151,N_13610);
and U17284 (N_17284,N_10254,N_14285);
nor U17285 (N_17285,N_10121,N_14051);
nand U17286 (N_17286,N_12323,N_11237);
nand U17287 (N_17287,N_11393,N_14159);
nand U17288 (N_17288,N_14952,N_12400);
nor U17289 (N_17289,N_10321,N_11144);
nand U17290 (N_17290,N_13586,N_10489);
or U17291 (N_17291,N_14265,N_13260);
and U17292 (N_17292,N_11702,N_10501);
nand U17293 (N_17293,N_13639,N_13374);
nor U17294 (N_17294,N_14586,N_13538);
nor U17295 (N_17295,N_11255,N_12957);
and U17296 (N_17296,N_11663,N_13875);
nand U17297 (N_17297,N_13077,N_10816);
nand U17298 (N_17298,N_11950,N_10980);
xor U17299 (N_17299,N_14055,N_13919);
or U17300 (N_17300,N_13806,N_12479);
nand U17301 (N_17301,N_11294,N_12782);
nor U17302 (N_17302,N_12910,N_13609);
nand U17303 (N_17303,N_11196,N_13807);
or U17304 (N_17304,N_10661,N_10881);
and U17305 (N_17305,N_14389,N_12906);
xnor U17306 (N_17306,N_10985,N_10775);
nand U17307 (N_17307,N_14434,N_14468);
and U17308 (N_17308,N_11298,N_13486);
nor U17309 (N_17309,N_14660,N_11636);
xnor U17310 (N_17310,N_13087,N_11089);
nand U17311 (N_17311,N_10324,N_13781);
and U17312 (N_17312,N_13536,N_14902);
nand U17313 (N_17313,N_10429,N_12454);
nand U17314 (N_17314,N_13257,N_13849);
nor U17315 (N_17315,N_11641,N_11581);
nor U17316 (N_17316,N_11402,N_13599);
nor U17317 (N_17317,N_11605,N_13575);
nand U17318 (N_17318,N_12331,N_13245);
nand U17319 (N_17319,N_11490,N_10653);
xor U17320 (N_17320,N_11617,N_14714);
or U17321 (N_17321,N_14278,N_10986);
and U17322 (N_17322,N_11421,N_14003);
or U17323 (N_17323,N_10974,N_14912);
and U17324 (N_17324,N_12275,N_12081);
nor U17325 (N_17325,N_11855,N_13337);
xnor U17326 (N_17326,N_10105,N_10799);
or U17327 (N_17327,N_10916,N_13434);
and U17328 (N_17328,N_13117,N_10664);
and U17329 (N_17329,N_14730,N_13492);
and U17330 (N_17330,N_11406,N_12758);
nand U17331 (N_17331,N_12897,N_13427);
nor U17332 (N_17332,N_11505,N_11930);
nand U17333 (N_17333,N_12938,N_10772);
nor U17334 (N_17334,N_10136,N_11225);
or U17335 (N_17335,N_12748,N_11336);
or U17336 (N_17336,N_13466,N_11170);
nor U17337 (N_17337,N_11112,N_11810);
and U17338 (N_17338,N_12991,N_14883);
xnor U17339 (N_17339,N_11540,N_14770);
or U17340 (N_17340,N_10576,N_13509);
nor U17341 (N_17341,N_14950,N_11303);
or U17342 (N_17342,N_10178,N_10175);
nand U17343 (N_17343,N_12001,N_11389);
and U17344 (N_17344,N_10066,N_11240);
xnor U17345 (N_17345,N_13133,N_11592);
nand U17346 (N_17346,N_12411,N_12924);
nor U17347 (N_17347,N_14280,N_11441);
nand U17348 (N_17348,N_10081,N_14017);
nor U17349 (N_17349,N_13025,N_12620);
nor U17350 (N_17350,N_14314,N_11042);
nand U17351 (N_17351,N_13372,N_10181);
and U17352 (N_17352,N_13467,N_10530);
and U17353 (N_17353,N_12202,N_12374);
or U17354 (N_17354,N_13907,N_12463);
and U17355 (N_17355,N_12376,N_14181);
or U17356 (N_17356,N_13970,N_11249);
xnor U17357 (N_17357,N_13264,N_11533);
nor U17358 (N_17358,N_10733,N_13497);
nor U17359 (N_17359,N_13881,N_10853);
or U17360 (N_17360,N_11360,N_12162);
and U17361 (N_17361,N_12891,N_13007);
and U17362 (N_17362,N_14420,N_11783);
or U17363 (N_17363,N_10052,N_12509);
nor U17364 (N_17364,N_10844,N_11631);
or U17365 (N_17365,N_11489,N_12037);
nand U17366 (N_17366,N_13189,N_10827);
xor U17367 (N_17367,N_12396,N_12414);
nand U17368 (N_17368,N_10124,N_12812);
and U17369 (N_17369,N_14621,N_11242);
nand U17370 (N_17370,N_11548,N_14651);
or U17371 (N_17371,N_14211,N_10745);
and U17372 (N_17372,N_10899,N_11261);
and U17373 (N_17373,N_12695,N_13113);
and U17374 (N_17374,N_13494,N_12575);
nand U17375 (N_17375,N_13006,N_10520);
nor U17376 (N_17376,N_10709,N_13580);
and U17377 (N_17377,N_14439,N_11478);
nand U17378 (N_17378,N_14593,N_10103);
nand U17379 (N_17379,N_13926,N_12348);
nor U17380 (N_17380,N_13549,N_12318);
and U17381 (N_17381,N_14841,N_13184);
nor U17382 (N_17382,N_12152,N_11920);
nor U17383 (N_17383,N_14580,N_13724);
nor U17384 (N_17384,N_14110,N_11593);
nand U17385 (N_17385,N_12157,N_10486);
xor U17386 (N_17386,N_11465,N_13404);
and U17387 (N_17387,N_10643,N_13368);
or U17388 (N_17388,N_14163,N_14612);
nand U17389 (N_17389,N_13156,N_11268);
or U17390 (N_17390,N_13343,N_13072);
nor U17391 (N_17391,N_13814,N_14646);
and U17392 (N_17392,N_13543,N_10419);
or U17393 (N_17393,N_14534,N_11223);
nand U17394 (N_17394,N_12365,N_12300);
and U17395 (N_17395,N_10042,N_10532);
nand U17396 (N_17396,N_10084,N_11382);
nor U17397 (N_17397,N_14209,N_14962);
and U17398 (N_17398,N_12341,N_12180);
nor U17399 (N_17399,N_13200,N_14422);
nor U17400 (N_17400,N_11974,N_13455);
and U17401 (N_17401,N_13515,N_12970);
nor U17402 (N_17402,N_11369,N_11890);
and U17403 (N_17403,N_12698,N_12617);
xnor U17404 (N_17404,N_14087,N_14449);
and U17405 (N_17405,N_10586,N_13474);
or U17406 (N_17406,N_10422,N_12423);
nor U17407 (N_17407,N_13208,N_10851);
or U17408 (N_17408,N_14648,N_10051);
nand U17409 (N_17409,N_10332,N_10989);
and U17410 (N_17410,N_14808,N_12839);
nor U17411 (N_17411,N_11885,N_13346);
nand U17412 (N_17412,N_10289,N_10265);
nand U17413 (N_17413,N_11642,N_10837);
and U17414 (N_17414,N_13660,N_13044);
nor U17415 (N_17415,N_13530,N_11383);
or U17416 (N_17416,N_10675,N_13893);
and U17417 (N_17417,N_10597,N_14753);
or U17418 (N_17418,N_10438,N_11346);
xnor U17419 (N_17419,N_11203,N_11803);
nor U17420 (N_17420,N_12051,N_13999);
nand U17421 (N_17421,N_11525,N_10448);
or U17422 (N_17422,N_10312,N_10443);
and U17423 (N_17423,N_13912,N_11973);
nor U17424 (N_17424,N_11059,N_12823);
and U17425 (N_17425,N_11455,N_14737);
or U17426 (N_17426,N_11423,N_11597);
nor U17427 (N_17427,N_13136,N_12643);
or U17428 (N_17428,N_14923,N_13111);
or U17429 (N_17429,N_12609,N_11968);
nand U17430 (N_17430,N_14638,N_10442);
nor U17431 (N_17431,N_13190,N_12754);
and U17432 (N_17432,N_14519,N_14354);
and U17433 (N_17433,N_14235,N_14198);
nand U17434 (N_17434,N_10297,N_12356);
and U17435 (N_17435,N_10908,N_12422);
or U17436 (N_17436,N_12191,N_11673);
and U17437 (N_17437,N_10953,N_13590);
or U17438 (N_17438,N_10678,N_10702);
nor U17439 (N_17439,N_11532,N_10162);
nand U17440 (N_17440,N_13556,N_12243);
nor U17441 (N_17441,N_12772,N_13417);
nor U17442 (N_17442,N_11748,N_11401);
and U17443 (N_17443,N_14363,N_10850);
or U17444 (N_17444,N_10912,N_14010);
nor U17445 (N_17445,N_13649,N_11722);
xnor U17446 (N_17446,N_14835,N_10984);
nand U17447 (N_17447,N_14862,N_11497);
nor U17448 (N_17448,N_12658,N_10050);
nor U17449 (N_17449,N_13052,N_14383);
and U17450 (N_17450,N_11251,N_10870);
nand U17451 (N_17451,N_13038,N_12804);
nor U17452 (N_17452,N_10298,N_14467);
and U17453 (N_17453,N_10513,N_10092);
xor U17454 (N_17454,N_13962,N_12900);
nand U17455 (N_17455,N_13602,N_11250);
nand U17456 (N_17456,N_14995,N_12572);
nor U17457 (N_17457,N_12476,N_14076);
nor U17458 (N_17458,N_14657,N_12221);
nand U17459 (N_17459,N_13780,N_10943);
or U17460 (N_17460,N_14610,N_13056);
nand U17461 (N_17461,N_14459,N_14398);
nor U17462 (N_17462,N_12478,N_13450);
nand U17463 (N_17463,N_10287,N_12577);
and U17464 (N_17464,N_12770,N_12130);
nand U17465 (N_17465,N_14299,N_14106);
nor U17466 (N_17466,N_10842,N_12473);
or U17467 (N_17467,N_12780,N_13348);
nand U17468 (N_17468,N_12385,N_10053);
and U17469 (N_17469,N_12868,N_10606);
nand U17470 (N_17470,N_11212,N_12099);
nor U17471 (N_17471,N_10792,N_11789);
or U17472 (N_17472,N_11785,N_14362);
nand U17473 (N_17473,N_12593,N_12245);
nor U17474 (N_17474,N_10331,N_14992);
nand U17475 (N_17475,N_12375,N_12115);
and U17476 (N_17476,N_14086,N_13030);
and U17477 (N_17477,N_11206,N_14679);
nor U17478 (N_17478,N_14263,N_13742);
nand U17479 (N_17479,N_13625,N_12737);
nand U17480 (N_17480,N_10477,N_12870);
and U17481 (N_17481,N_12505,N_14984);
or U17482 (N_17482,N_11721,N_13597);
nor U17483 (N_17483,N_11027,N_11032);
or U17484 (N_17484,N_13410,N_11812);
and U17485 (N_17485,N_14259,N_12999);
nor U17486 (N_17486,N_11777,N_10196);
nor U17487 (N_17487,N_11813,N_10798);
nand U17488 (N_17488,N_11736,N_13399);
or U17489 (N_17489,N_11718,N_11668);
nor U17490 (N_17490,N_12842,N_11725);
nand U17491 (N_17491,N_13816,N_11197);
nand U17492 (N_17492,N_10821,N_12449);
or U17493 (N_17493,N_11121,N_12072);
or U17494 (N_17494,N_13145,N_12952);
nand U17495 (N_17495,N_13269,N_14222);
or U17496 (N_17496,N_13693,N_12460);
or U17497 (N_17497,N_13799,N_10177);
or U17498 (N_17498,N_11680,N_12403);
or U17499 (N_17499,N_12321,N_13899);
or U17500 (N_17500,N_14710,N_14110);
or U17501 (N_17501,N_11343,N_12698);
and U17502 (N_17502,N_11745,N_12873);
and U17503 (N_17503,N_14174,N_14487);
and U17504 (N_17504,N_11925,N_13521);
and U17505 (N_17505,N_14683,N_12802);
or U17506 (N_17506,N_10673,N_11559);
or U17507 (N_17507,N_13158,N_14106);
nor U17508 (N_17508,N_11198,N_10274);
or U17509 (N_17509,N_13374,N_12094);
nand U17510 (N_17510,N_13836,N_12204);
or U17511 (N_17511,N_11755,N_10971);
nand U17512 (N_17512,N_13059,N_14144);
or U17513 (N_17513,N_13060,N_14963);
and U17514 (N_17514,N_14622,N_13630);
nor U17515 (N_17515,N_10455,N_12928);
nor U17516 (N_17516,N_12477,N_14188);
and U17517 (N_17517,N_11855,N_11351);
nand U17518 (N_17518,N_13980,N_10390);
nor U17519 (N_17519,N_12573,N_11361);
xor U17520 (N_17520,N_10589,N_13301);
and U17521 (N_17521,N_11159,N_10750);
or U17522 (N_17522,N_12344,N_10464);
nand U17523 (N_17523,N_10553,N_12647);
or U17524 (N_17524,N_13797,N_13757);
nor U17525 (N_17525,N_10640,N_13956);
nand U17526 (N_17526,N_10876,N_12200);
xor U17527 (N_17527,N_14783,N_13965);
nor U17528 (N_17528,N_12236,N_13432);
nand U17529 (N_17529,N_14644,N_13731);
xnor U17530 (N_17530,N_14792,N_12979);
nor U17531 (N_17531,N_12403,N_12969);
nor U17532 (N_17532,N_13794,N_12339);
nor U17533 (N_17533,N_11206,N_10821);
xor U17534 (N_17534,N_13433,N_13478);
nor U17535 (N_17535,N_12015,N_14652);
nor U17536 (N_17536,N_11274,N_13124);
or U17537 (N_17537,N_12065,N_10353);
or U17538 (N_17538,N_12346,N_11259);
nand U17539 (N_17539,N_11691,N_14575);
or U17540 (N_17540,N_12459,N_11875);
xor U17541 (N_17541,N_14379,N_12221);
xnor U17542 (N_17542,N_13033,N_14835);
or U17543 (N_17543,N_14588,N_12221);
xor U17544 (N_17544,N_10085,N_11211);
and U17545 (N_17545,N_11702,N_11226);
and U17546 (N_17546,N_11274,N_13227);
or U17547 (N_17547,N_11277,N_11909);
and U17548 (N_17548,N_12616,N_13631);
and U17549 (N_17549,N_10122,N_10231);
and U17550 (N_17550,N_11197,N_14573);
xor U17551 (N_17551,N_14483,N_14505);
and U17552 (N_17552,N_10091,N_10451);
xor U17553 (N_17553,N_12746,N_10559);
nor U17554 (N_17554,N_12953,N_13332);
nand U17555 (N_17555,N_12405,N_11508);
nor U17556 (N_17556,N_14834,N_11016);
or U17557 (N_17557,N_14095,N_10719);
and U17558 (N_17558,N_13585,N_10357);
nand U17559 (N_17559,N_11118,N_13295);
and U17560 (N_17560,N_10532,N_10049);
nor U17561 (N_17561,N_14555,N_12842);
xnor U17562 (N_17562,N_12071,N_11453);
nand U17563 (N_17563,N_14107,N_13222);
xor U17564 (N_17564,N_12475,N_12980);
and U17565 (N_17565,N_10757,N_14333);
nand U17566 (N_17566,N_12184,N_12807);
and U17567 (N_17567,N_14916,N_12172);
or U17568 (N_17568,N_10518,N_13985);
nor U17569 (N_17569,N_12292,N_14555);
xnor U17570 (N_17570,N_11353,N_10711);
or U17571 (N_17571,N_11614,N_10228);
nor U17572 (N_17572,N_12841,N_10856);
and U17573 (N_17573,N_12898,N_10190);
nand U17574 (N_17574,N_12860,N_13114);
nor U17575 (N_17575,N_12761,N_12872);
or U17576 (N_17576,N_13628,N_11840);
and U17577 (N_17577,N_13820,N_14679);
nor U17578 (N_17578,N_12898,N_13172);
or U17579 (N_17579,N_14832,N_11753);
nand U17580 (N_17580,N_13623,N_12183);
nor U17581 (N_17581,N_13634,N_13890);
nand U17582 (N_17582,N_10455,N_13199);
or U17583 (N_17583,N_13872,N_14790);
nor U17584 (N_17584,N_13060,N_13255);
or U17585 (N_17585,N_10437,N_11590);
nor U17586 (N_17586,N_14579,N_14702);
and U17587 (N_17587,N_14769,N_14420);
and U17588 (N_17588,N_11460,N_13902);
or U17589 (N_17589,N_12268,N_10896);
nor U17590 (N_17590,N_11265,N_14218);
nor U17591 (N_17591,N_14967,N_13608);
nor U17592 (N_17592,N_13371,N_11997);
nand U17593 (N_17593,N_14137,N_14260);
and U17594 (N_17594,N_14614,N_11284);
nand U17595 (N_17595,N_11225,N_10656);
or U17596 (N_17596,N_12518,N_12523);
nor U17597 (N_17597,N_10115,N_13226);
nor U17598 (N_17598,N_12486,N_10881);
xnor U17599 (N_17599,N_10124,N_14600);
xor U17600 (N_17600,N_14704,N_12646);
and U17601 (N_17601,N_12740,N_12359);
nor U17602 (N_17602,N_10777,N_14047);
nor U17603 (N_17603,N_11533,N_14846);
xnor U17604 (N_17604,N_12595,N_11551);
and U17605 (N_17605,N_12326,N_12225);
or U17606 (N_17606,N_11090,N_14443);
nor U17607 (N_17607,N_11243,N_12351);
nand U17608 (N_17608,N_10468,N_12975);
or U17609 (N_17609,N_11674,N_11700);
nand U17610 (N_17610,N_11729,N_11663);
and U17611 (N_17611,N_14705,N_10355);
nor U17612 (N_17612,N_10996,N_12785);
and U17613 (N_17613,N_10689,N_14702);
nor U17614 (N_17614,N_10789,N_13324);
or U17615 (N_17615,N_10693,N_11757);
nor U17616 (N_17616,N_13196,N_14859);
xnor U17617 (N_17617,N_13505,N_11852);
or U17618 (N_17618,N_13317,N_10649);
or U17619 (N_17619,N_14690,N_10576);
xnor U17620 (N_17620,N_12329,N_10166);
nand U17621 (N_17621,N_13596,N_10709);
nor U17622 (N_17622,N_13910,N_10076);
or U17623 (N_17623,N_11694,N_10059);
nand U17624 (N_17624,N_11300,N_11581);
nand U17625 (N_17625,N_14946,N_12050);
nor U17626 (N_17626,N_13573,N_10935);
or U17627 (N_17627,N_14139,N_14495);
nor U17628 (N_17628,N_12395,N_12764);
nand U17629 (N_17629,N_12622,N_12816);
or U17630 (N_17630,N_12889,N_14104);
and U17631 (N_17631,N_13142,N_12153);
nand U17632 (N_17632,N_11740,N_14936);
xor U17633 (N_17633,N_14860,N_14255);
and U17634 (N_17634,N_10521,N_10171);
or U17635 (N_17635,N_11513,N_10137);
and U17636 (N_17636,N_12617,N_14892);
and U17637 (N_17637,N_10348,N_14990);
nor U17638 (N_17638,N_12958,N_14301);
nand U17639 (N_17639,N_14980,N_13641);
or U17640 (N_17640,N_10986,N_11540);
nor U17641 (N_17641,N_12707,N_13825);
and U17642 (N_17642,N_10489,N_14106);
and U17643 (N_17643,N_11816,N_14139);
or U17644 (N_17644,N_11256,N_10708);
and U17645 (N_17645,N_10629,N_12007);
or U17646 (N_17646,N_14543,N_14881);
nor U17647 (N_17647,N_14140,N_14570);
nor U17648 (N_17648,N_10967,N_13587);
or U17649 (N_17649,N_11428,N_13279);
or U17650 (N_17650,N_11300,N_10444);
or U17651 (N_17651,N_11923,N_12911);
nor U17652 (N_17652,N_12400,N_13069);
and U17653 (N_17653,N_12150,N_11452);
and U17654 (N_17654,N_13856,N_12294);
and U17655 (N_17655,N_12114,N_12909);
nor U17656 (N_17656,N_11650,N_14875);
nor U17657 (N_17657,N_10031,N_10173);
and U17658 (N_17658,N_10267,N_14781);
or U17659 (N_17659,N_13464,N_10871);
xnor U17660 (N_17660,N_13966,N_13174);
nor U17661 (N_17661,N_10411,N_12194);
xnor U17662 (N_17662,N_10849,N_14831);
or U17663 (N_17663,N_11710,N_12166);
or U17664 (N_17664,N_14877,N_13005);
or U17665 (N_17665,N_10884,N_12845);
and U17666 (N_17666,N_11540,N_13883);
or U17667 (N_17667,N_13698,N_10346);
nand U17668 (N_17668,N_11227,N_12804);
and U17669 (N_17669,N_12938,N_13059);
nor U17670 (N_17670,N_10166,N_13231);
or U17671 (N_17671,N_12510,N_11955);
nand U17672 (N_17672,N_13329,N_13766);
and U17673 (N_17673,N_12647,N_10112);
nand U17674 (N_17674,N_11564,N_14301);
nor U17675 (N_17675,N_11069,N_13623);
xor U17676 (N_17676,N_10710,N_10917);
or U17677 (N_17677,N_13719,N_10736);
and U17678 (N_17678,N_13347,N_12059);
xnor U17679 (N_17679,N_12130,N_10106);
or U17680 (N_17680,N_11929,N_14519);
nor U17681 (N_17681,N_12806,N_14086);
nand U17682 (N_17682,N_11564,N_10264);
nor U17683 (N_17683,N_11162,N_14587);
nor U17684 (N_17684,N_11868,N_13292);
nand U17685 (N_17685,N_10062,N_12405);
nor U17686 (N_17686,N_11354,N_12818);
nand U17687 (N_17687,N_13100,N_10949);
and U17688 (N_17688,N_12931,N_12316);
xor U17689 (N_17689,N_10697,N_12992);
or U17690 (N_17690,N_12067,N_13523);
and U17691 (N_17691,N_11087,N_11094);
nand U17692 (N_17692,N_13921,N_12062);
xnor U17693 (N_17693,N_12750,N_13987);
or U17694 (N_17694,N_12554,N_12810);
and U17695 (N_17695,N_11547,N_14382);
or U17696 (N_17696,N_10523,N_13539);
nand U17697 (N_17697,N_14534,N_11805);
or U17698 (N_17698,N_13181,N_10018);
and U17699 (N_17699,N_11743,N_11766);
nand U17700 (N_17700,N_10412,N_10809);
nand U17701 (N_17701,N_10558,N_12296);
nor U17702 (N_17702,N_11998,N_10886);
or U17703 (N_17703,N_10927,N_13858);
or U17704 (N_17704,N_12503,N_11126);
nand U17705 (N_17705,N_10177,N_14707);
or U17706 (N_17706,N_13798,N_13456);
nand U17707 (N_17707,N_10038,N_12704);
and U17708 (N_17708,N_13858,N_10125);
or U17709 (N_17709,N_14934,N_14185);
xor U17710 (N_17710,N_10791,N_10810);
and U17711 (N_17711,N_14446,N_12252);
and U17712 (N_17712,N_14028,N_11376);
nand U17713 (N_17713,N_10992,N_11424);
nor U17714 (N_17714,N_14904,N_11134);
or U17715 (N_17715,N_14940,N_12111);
nor U17716 (N_17716,N_13049,N_13403);
nand U17717 (N_17717,N_13335,N_11201);
nand U17718 (N_17718,N_14407,N_10979);
nor U17719 (N_17719,N_11448,N_12733);
and U17720 (N_17720,N_14712,N_11288);
and U17721 (N_17721,N_12577,N_13058);
nor U17722 (N_17722,N_12358,N_11656);
and U17723 (N_17723,N_11404,N_11129);
or U17724 (N_17724,N_14211,N_14695);
xnor U17725 (N_17725,N_12575,N_13749);
or U17726 (N_17726,N_13945,N_12164);
nand U17727 (N_17727,N_11294,N_12161);
xnor U17728 (N_17728,N_11179,N_12155);
and U17729 (N_17729,N_11825,N_13187);
nand U17730 (N_17730,N_12452,N_14873);
and U17731 (N_17731,N_14480,N_13347);
and U17732 (N_17732,N_14211,N_11653);
or U17733 (N_17733,N_14487,N_13669);
or U17734 (N_17734,N_12984,N_10746);
or U17735 (N_17735,N_13435,N_10065);
or U17736 (N_17736,N_10660,N_11886);
nor U17737 (N_17737,N_14380,N_13356);
xnor U17738 (N_17738,N_12335,N_10162);
xnor U17739 (N_17739,N_13025,N_10356);
or U17740 (N_17740,N_11669,N_12796);
or U17741 (N_17741,N_11184,N_10950);
and U17742 (N_17742,N_10911,N_12857);
and U17743 (N_17743,N_11942,N_13187);
nand U17744 (N_17744,N_10813,N_12493);
and U17745 (N_17745,N_14514,N_14310);
and U17746 (N_17746,N_14535,N_11615);
nand U17747 (N_17747,N_10460,N_14614);
or U17748 (N_17748,N_10283,N_11595);
nor U17749 (N_17749,N_14654,N_11058);
nand U17750 (N_17750,N_12305,N_11163);
nor U17751 (N_17751,N_12379,N_13887);
and U17752 (N_17752,N_13829,N_11363);
xnor U17753 (N_17753,N_14614,N_14822);
nor U17754 (N_17754,N_10441,N_13348);
nand U17755 (N_17755,N_14123,N_12092);
or U17756 (N_17756,N_13007,N_12509);
and U17757 (N_17757,N_12687,N_12829);
and U17758 (N_17758,N_12373,N_10691);
xor U17759 (N_17759,N_11360,N_12457);
nand U17760 (N_17760,N_14147,N_13901);
xnor U17761 (N_17761,N_13043,N_10747);
xor U17762 (N_17762,N_14856,N_12787);
and U17763 (N_17763,N_13841,N_14994);
nand U17764 (N_17764,N_10062,N_13185);
and U17765 (N_17765,N_12686,N_10792);
and U17766 (N_17766,N_13671,N_13697);
xnor U17767 (N_17767,N_11730,N_13868);
or U17768 (N_17768,N_14043,N_14778);
and U17769 (N_17769,N_11680,N_10631);
xor U17770 (N_17770,N_11502,N_12854);
or U17771 (N_17771,N_10982,N_14362);
nor U17772 (N_17772,N_11556,N_11371);
and U17773 (N_17773,N_11103,N_14655);
or U17774 (N_17774,N_11104,N_11939);
or U17775 (N_17775,N_14349,N_11665);
or U17776 (N_17776,N_13741,N_12331);
or U17777 (N_17777,N_13170,N_11896);
or U17778 (N_17778,N_13122,N_13945);
or U17779 (N_17779,N_14918,N_13642);
nand U17780 (N_17780,N_12001,N_11416);
nor U17781 (N_17781,N_12044,N_13607);
or U17782 (N_17782,N_13733,N_12811);
or U17783 (N_17783,N_12272,N_10071);
nand U17784 (N_17784,N_12987,N_14693);
nand U17785 (N_17785,N_13925,N_12472);
and U17786 (N_17786,N_10874,N_12699);
and U17787 (N_17787,N_10694,N_10391);
nand U17788 (N_17788,N_13639,N_10564);
xnor U17789 (N_17789,N_14345,N_14289);
or U17790 (N_17790,N_11008,N_11866);
and U17791 (N_17791,N_13262,N_12330);
and U17792 (N_17792,N_11889,N_11332);
or U17793 (N_17793,N_14916,N_12279);
and U17794 (N_17794,N_11112,N_10747);
and U17795 (N_17795,N_11479,N_11235);
or U17796 (N_17796,N_14720,N_13834);
and U17797 (N_17797,N_13218,N_14846);
nand U17798 (N_17798,N_10186,N_14996);
or U17799 (N_17799,N_12409,N_14605);
or U17800 (N_17800,N_10935,N_14035);
nand U17801 (N_17801,N_14002,N_10625);
xor U17802 (N_17802,N_10780,N_11681);
and U17803 (N_17803,N_14938,N_11041);
and U17804 (N_17804,N_10293,N_12392);
nand U17805 (N_17805,N_11498,N_13851);
nand U17806 (N_17806,N_11338,N_13781);
nand U17807 (N_17807,N_14392,N_14079);
xor U17808 (N_17808,N_14421,N_13779);
xor U17809 (N_17809,N_14108,N_14776);
nor U17810 (N_17810,N_14881,N_11704);
xor U17811 (N_17811,N_11357,N_10217);
nand U17812 (N_17812,N_11898,N_14774);
nor U17813 (N_17813,N_14358,N_10361);
and U17814 (N_17814,N_10218,N_14808);
xnor U17815 (N_17815,N_13956,N_13935);
nand U17816 (N_17816,N_10303,N_12632);
or U17817 (N_17817,N_14431,N_11381);
nand U17818 (N_17818,N_14038,N_12836);
nor U17819 (N_17819,N_10807,N_13218);
and U17820 (N_17820,N_12354,N_14337);
nand U17821 (N_17821,N_10840,N_10043);
nand U17822 (N_17822,N_13330,N_14715);
nor U17823 (N_17823,N_13097,N_10411);
and U17824 (N_17824,N_14319,N_10342);
nor U17825 (N_17825,N_11839,N_10307);
or U17826 (N_17826,N_10024,N_13612);
and U17827 (N_17827,N_14965,N_13745);
nor U17828 (N_17828,N_12822,N_12221);
nor U17829 (N_17829,N_10297,N_13643);
or U17830 (N_17830,N_12328,N_13861);
nor U17831 (N_17831,N_12595,N_13737);
nand U17832 (N_17832,N_14351,N_11921);
xnor U17833 (N_17833,N_10097,N_11298);
nor U17834 (N_17834,N_12857,N_13495);
and U17835 (N_17835,N_13461,N_14986);
nor U17836 (N_17836,N_11868,N_10928);
nor U17837 (N_17837,N_11164,N_12272);
nand U17838 (N_17838,N_12759,N_12632);
or U17839 (N_17839,N_13447,N_10140);
and U17840 (N_17840,N_11881,N_11603);
nand U17841 (N_17841,N_11549,N_10814);
nand U17842 (N_17842,N_13430,N_12824);
nand U17843 (N_17843,N_11184,N_14166);
and U17844 (N_17844,N_11963,N_11756);
or U17845 (N_17845,N_12228,N_12923);
and U17846 (N_17846,N_11398,N_11667);
nor U17847 (N_17847,N_13971,N_11141);
or U17848 (N_17848,N_12895,N_14647);
xor U17849 (N_17849,N_12798,N_12629);
nor U17850 (N_17850,N_13490,N_14220);
nand U17851 (N_17851,N_11558,N_10221);
nand U17852 (N_17852,N_14191,N_14230);
nand U17853 (N_17853,N_10706,N_12614);
or U17854 (N_17854,N_13503,N_13211);
and U17855 (N_17855,N_11252,N_14721);
or U17856 (N_17856,N_13544,N_11216);
xor U17857 (N_17857,N_11884,N_13423);
or U17858 (N_17858,N_11727,N_14318);
nor U17859 (N_17859,N_10864,N_11449);
nand U17860 (N_17860,N_11975,N_13311);
or U17861 (N_17861,N_10302,N_12409);
nor U17862 (N_17862,N_12539,N_11402);
or U17863 (N_17863,N_12300,N_11157);
nor U17864 (N_17864,N_11907,N_13217);
nor U17865 (N_17865,N_10066,N_14171);
nand U17866 (N_17866,N_13030,N_13910);
and U17867 (N_17867,N_11144,N_13006);
or U17868 (N_17868,N_12770,N_11469);
nor U17869 (N_17869,N_11033,N_13742);
nor U17870 (N_17870,N_10624,N_10729);
and U17871 (N_17871,N_12921,N_11395);
and U17872 (N_17872,N_12536,N_12056);
nand U17873 (N_17873,N_14503,N_10042);
or U17874 (N_17874,N_13837,N_12095);
or U17875 (N_17875,N_13487,N_12313);
nor U17876 (N_17876,N_11963,N_13542);
xnor U17877 (N_17877,N_13777,N_12112);
xor U17878 (N_17878,N_12071,N_13848);
and U17879 (N_17879,N_14989,N_13626);
and U17880 (N_17880,N_10020,N_10271);
or U17881 (N_17881,N_13259,N_14590);
or U17882 (N_17882,N_14370,N_14016);
nor U17883 (N_17883,N_10269,N_11258);
or U17884 (N_17884,N_10823,N_13156);
nand U17885 (N_17885,N_14126,N_12394);
nand U17886 (N_17886,N_13878,N_10195);
nor U17887 (N_17887,N_10912,N_12195);
nand U17888 (N_17888,N_12074,N_11369);
nand U17889 (N_17889,N_10849,N_10525);
nor U17890 (N_17890,N_14842,N_14593);
xnor U17891 (N_17891,N_13252,N_10414);
nor U17892 (N_17892,N_10118,N_13876);
or U17893 (N_17893,N_10230,N_11804);
nor U17894 (N_17894,N_13775,N_11036);
or U17895 (N_17895,N_12640,N_11312);
nor U17896 (N_17896,N_13387,N_11083);
nor U17897 (N_17897,N_10368,N_14971);
nand U17898 (N_17898,N_11758,N_12613);
or U17899 (N_17899,N_14890,N_10869);
nand U17900 (N_17900,N_12939,N_10780);
nor U17901 (N_17901,N_14875,N_10497);
nor U17902 (N_17902,N_11374,N_14275);
and U17903 (N_17903,N_11233,N_12584);
or U17904 (N_17904,N_14142,N_11854);
nor U17905 (N_17905,N_10819,N_13450);
nor U17906 (N_17906,N_10392,N_11972);
and U17907 (N_17907,N_12959,N_12503);
nor U17908 (N_17908,N_10160,N_12363);
xor U17909 (N_17909,N_11049,N_11521);
nand U17910 (N_17910,N_14253,N_13286);
and U17911 (N_17911,N_13697,N_12115);
or U17912 (N_17912,N_10836,N_12794);
and U17913 (N_17913,N_12409,N_13364);
and U17914 (N_17914,N_13458,N_11842);
or U17915 (N_17915,N_13237,N_10318);
xnor U17916 (N_17916,N_11952,N_14665);
or U17917 (N_17917,N_10122,N_12326);
and U17918 (N_17918,N_14428,N_10426);
nand U17919 (N_17919,N_12446,N_11956);
nor U17920 (N_17920,N_14935,N_13364);
and U17921 (N_17921,N_13399,N_14995);
or U17922 (N_17922,N_12347,N_13029);
xnor U17923 (N_17923,N_13932,N_14903);
and U17924 (N_17924,N_14880,N_10907);
and U17925 (N_17925,N_14569,N_12442);
and U17926 (N_17926,N_14094,N_13511);
or U17927 (N_17927,N_13231,N_10176);
nor U17928 (N_17928,N_11279,N_10503);
nor U17929 (N_17929,N_11292,N_12839);
or U17930 (N_17930,N_13062,N_13623);
nand U17931 (N_17931,N_10815,N_11821);
nor U17932 (N_17932,N_12432,N_14422);
nor U17933 (N_17933,N_14256,N_13413);
or U17934 (N_17934,N_11331,N_12885);
xor U17935 (N_17935,N_13205,N_11243);
nor U17936 (N_17936,N_12523,N_14956);
nor U17937 (N_17937,N_11026,N_14708);
nand U17938 (N_17938,N_12474,N_14465);
and U17939 (N_17939,N_11632,N_12168);
nand U17940 (N_17940,N_14170,N_10007);
and U17941 (N_17941,N_10229,N_13839);
nand U17942 (N_17942,N_14753,N_12111);
nor U17943 (N_17943,N_11634,N_11737);
nor U17944 (N_17944,N_10401,N_12508);
and U17945 (N_17945,N_10083,N_14318);
nand U17946 (N_17946,N_11188,N_11378);
nand U17947 (N_17947,N_10077,N_12245);
nor U17948 (N_17948,N_12797,N_14428);
nand U17949 (N_17949,N_11185,N_10294);
xor U17950 (N_17950,N_13884,N_11196);
nand U17951 (N_17951,N_13381,N_13432);
nand U17952 (N_17952,N_11589,N_11299);
or U17953 (N_17953,N_11633,N_13388);
nand U17954 (N_17954,N_10643,N_13453);
nand U17955 (N_17955,N_10984,N_10952);
or U17956 (N_17956,N_14687,N_10873);
nand U17957 (N_17957,N_13972,N_13362);
or U17958 (N_17958,N_11168,N_11775);
nor U17959 (N_17959,N_14468,N_13717);
nand U17960 (N_17960,N_11561,N_10378);
or U17961 (N_17961,N_14208,N_11104);
or U17962 (N_17962,N_13851,N_13504);
or U17963 (N_17963,N_11523,N_10277);
or U17964 (N_17964,N_11459,N_12423);
nor U17965 (N_17965,N_11793,N_11863);
or U17966 (N_17966,N_10278,N_13310);
xor U17967 (N_17967,N_12422,N_14655);
or U17968 (N_17968,N_11972,N_12829);
and U17969 (N_17969,N_14871,N_13883);
or U17970 (N_17970,N_14824,N_14108);
and U17971 (N_17971,N_13719,N_13479);
or U17972 (N_17972,N_14109,N_12415);
and U17973 (N_17973,N_11146,N_12766);
nor U17974 (N_17974,N_12022,N_10626);
or U17975 (N_17975,N_11118,N_11499);
xnor U17976 (N_17976,N_12817,N_11220);
nor U17977 (N_17977,N_14414,N_11955);
nor U17978 (N_17978,N_14551,N_13670);
nor U17979 (N_17979,N_11358,N_12016);
xor U17980 (N_17980,N_12811,N_13902);
or U17981 (N_17981,N_10622,N_10304);
nand U17982 (N_17982,N_13256,N_14686);
xnor U17983 (N_17983,N_11673,N_12447);
or U17984 (N_17984,N_14381,N_14245);
nor U17985 (N_17985,N_12579,N_13748);
and U17986 (N_17986,N_14229,N_10406);
xor U17987 (N_17987,N_11274,N_11107);
nand U17988 (N_17988,N_12571,N_13060);
or U17989 (N_17989,N_11085,N_10528);
nand U17990 (N_17990,N_11006,N_14275);
and U17991 (N_17991,N_13968,N_13264);
or U17992 (N_17992,N_12844,N_10307);
or U17993 (N_17993,N_10129,N_11723);
nor U17994 (N_17994,N_11075,N_14916);
xnor U17995 (N_17995,N_10579,N_12318);
nand U17996 (N_17996,N_11922,N_11727);
nand U17997 (N_17997,N_13570,N_11758);
and U17998 (N_17998,N_13542,N_13969);
and U17999 (N_17999,N_13215,N_11315);
nor U18000 (N_18000,N_12244,N_11668);
nand U18001 (N_18001,N_14320,N_12488);
and U18002 (N_18002,N_10755,N_11961);
or U18003 (N_18003,N_10563,N_10613);
or U18004 (N_18004,N_11695,N_12674);
xor U18005 (N_18005,N_13664,N_12767);
nand U18006 (N_18006,N_10368,N_12586);
and U18007 (N_18007,N_14224,N_13262);
or U18008 (N_18008,N_11306,N_11670);
or U18009 (N_18009,N_13473,N_10429);
and U18010 (N_18010,N_11642,N_14082);
nor U18011 (N_18011,N_10191,N_12974);
nand U18012 (N_18012,N_14184,N_12427);
and U18013 (N_18013,N_12352,N_14313);
or U18014 (N_18014,N_12481,N_14872);
and U18015 (N_18015,N_13179,N_11882);
nand U18016 (N_18016,N_11650,N_10387);
or U18017 (N_18017,N_11422,N_14521);
or U18018 (N_18018,N_10726,N_10101);
or U18019 (N_18019,N_12683,N_14457);
or U18020 (N_18020,N_13544,N_10707);
nor U18021 (N_18021,N_14278,N_14464);
and U18022 (N_18022,N_13349,N_12862);
and U18023 (N_18023,N_13780,N_11378);
nand U18024 (N_18024,N_14570,N_13398);
nand U18025 (N_18025,N_14121,N_10690);
and U18026 (N_18026,N_12353,N_12630);
or U18027 (N_18027,N_12371,N_12126);
and U18028 (N_18028,N_10909,N_11091);
and U18029 (N_18029,N_14058,N_11688);
nand U18030 (N_18030,N_13518,N_10866);
nand U18031 (N_18031,N_13311,N_11830);
or U18032 (N_18032,N_14985,N_13020);
and U18033 (N_18033,N_11454,N_14131);
and U18034 (N_18034,N_12738,N_14407);
or U18035 (N_18035,N_13829,N_13145);
nor U18036 (N_18036,N_12286,N_10044);
nand U18037 (N_18037,N_11024,N_12438);
and U18038 (N_18038,N_10548,N_10185);
or U18039 (N_18039,N_10475,N_11310);
xor U18040 (N_18040,N_13515,N_14700);
nor U18041 (N_18041,N_12932,N_12765);
and U18042 (N_18042,N_12069,N_10941);
or U18043 (N_18043,N_11984,N_12156);
or U18044 (N_18044,N_14401,N_13198);
or U18045 (N_18045,N_11323,N_11848);
nor U18046 (N_18046,N_10117,N_14446);
or U18047 (N_18047,N_12562,N_11162);
nor U18048 (N_18048,N_12921,N_12551);
nand U18049 (N_18049,N_14061,N_11965);
and U18050 (N_18050,N_12511,N_11919);
or U18051 (N_18051,N_10664,N_14923);
nand U18052 (N_18052,N_11750,N_13419);
nand U18053 (N_18053,N_14839,N_13676);
nor U18054 (N_18054,N_11883,N_14576);
or U18055 (N_18055,N_13342,N_12853);
nor U18056 (N_18056,N_12501,N_10717);
and U18057 (N_18057,N_14112,N_11302);
and U18058 (N_18058,N_11515,N_11114);
nor U18059 (N_18059,N_10221,N_12322);
nand U18060 (N_18060,N_13001,N_14052);
or U18061 (N_18061,N_14356,N_13903);
and U18062 (N_18062,N_10242,N_12984);
and U18063 (N_18063,N_13076,N_13442);
nor U18064 (N_18064,N_12257,N_14624);
xor U18065 (N_18065,N_14117,N_12404);
xnor U18066 (N_18066,N_10965,N_11166);
nand U18067 (N_18067,N_11230,N_12938);
xor U18068 (N_18068,N_13197,N_11035);
and U18069 (N_18069,N_13016,N_13858);
and U18070 (N_18070,N_13371,N_12962);
nor U18071 (N_18071,N_13050,N_13065);
nor U18072 (N_18072,N_13556,N_10388);
nand U18073 (N_18073,N_10164,N_14083);
and U18074 (N_18074,N_14867,N_11223);
or U18075 (N_18075,N_12096,N_12401);
and U18076 (N_18076,N_12826,N_13904);
or U18077 (N_18077,N_11896,N_14934);
nand U18078 (N_18078,N_11770,N_10290);
or U18079 (N_18079,N_11140,N_12201);
nor U18080 (N_18080,N_13452,N_12999);
xor U18081 (N_18081,N_12388,N_14504);
and U18082 (N_18082,N_10340,N_14875);
xnor U18083 (N_18083,N_12575,N_14957);
nor U18084 (N_18084,N_11623,N_11164);
xnor U18085 (N_18085,N_10228,N_12439);
or U18086 (N_18086,N_12069,N_13364);
nor U18087 (N_18087,N_14986,N_13539);
nand U18088 (N_18088,N_11242,N_14716);
and U18089 (N_18089,N_12052,N_14456);
nor U18090 (N_18090,N_14253,N_14243);
or U18091 (N_18091,N_14078,N_11309);
or U18092 (N_18092,N_13752,N_10683);
and U18093 (N_18093,N_11969,N_11632);
and U18094 (N_18094,N_11432,N_13350);
nand U18095 (N_18095,N_10819,N_10547);
and U18096 (N_18096,N_14004,N_14817);
nor U18097 (N_18097,N_11186,N_11190);
nand U18098 (N_18098,N_12628,N_10536);
or U18099 (N_18099,N_11151,N_11964);
nor U18100 (N_18100,N_14665,N_10052);
and U18101 (N_18101,N_13339,N_10793);
or U18102 (N_18102,N_13771,N_12375);
or U18103 (N_18103,N_13811,N_11353);
and U18104 (N_18104,N_12141,N_12237);
or U18105 (N_18105,N_12890,N_14259);
xor U18106 (N_18106,N_12425,N_12662);
nand U18107 (N_18107,N_10646,N_10401);
or U18108 (N_18108,N_11951,N_10672);
nor U18109 (N_18109,N_12709,N_11919);
or U18110 (N_18110,N_14692,N_11602);
nor U18111 (N_18111,N_11153,N_10942);
nand U18112 (N_18112,N_11384,N_14676);
or U18113 (N_18113,N_12794,N_11238);
nor U18114 (N_18114,N_10099,N_11816);
nor U18115 (N_18115,N_10502,N_11195);
or U18116 (N_18116,N_12321,N_13843);
xnor U18117 (N_18117,N_12082,N_12745);
and U18118 (N_18118,N_10204,N_14921);
nor U18119 (N_18119,N_12118,N_11472);
and U18120 (N_18120,N_12050,N_11234);
nand U18121 (N_18121,N_14443,N_14367);
nand U18122 (N_18122,N_14192,N_12025);
or U18123 (N_18123,N_12018,N_14390);
nand U18124 (N_18124,N_10787,N_11973);
nor U18125 (N_18125,N_12628,N_12203);
xnor U18126 (N_18126,N_10635,N_14044);
and U18127 (N_18127,N_13441,N_11200);
nand U18128 (N_18128,N_13189,N_14548);
nand U18129 (N_18129,N_13495,N_10745);
and U18130 (N_18130,N_14546,N_13411);
and U18131 (N_18131,N_14114,N_11382);
nor U18132 (N_18132,N_11982,N_14546);
or U18133 (N_18133,N_12320,N_12350);
nor U18134 (N_18134,N_12828,N_10762);
nor U18135 (N_18135,N_14489,N_13191);
xnor U18136 (N_18136,N_13973,N_12067);
or U18137 (N_18137,N_10714,N_13385);
or U18138 (N_18138,N_13981,N_14340);
xor U18139 (N_18139,N_11857,N_11541);
and U18140 (N_18140,N_12838,N_14691);
and U18141 (N_18141,N_13863,N_13690);
nand U18142 (N_18142,N_11670,N_12837);
nor U18143 (N_18143,N_12073,N_11328);
nand U18144 (N_18144,N_11009,N_14609);
nor U18145 (N_18145,N_13795,N_14100);
xnor U18146 (N_18146,N_14872,N_10203);
and U18147 (N_18147,N_11003,N_11902);
nand U18148 (N_18148,N_14089,N_14563);
nand U18149 (N_18149,N_10518,N_10080);
nand U18150 (N_18150,N_14758,N_12426);
xor U18151 (N_18151,N_10352,N_10800);
and U18152 (N_18152,N_13305,N_10546);
nor U18153 (N_18153,N_10020,N_11677);
and U18154 (N_18154,N_13935,N_14127);
nand U18155 (N_18155,N_12150,N_10554);
nor U18156 (N_18156,N_13402,N_14638);
nor U18157 (N_18157,N_11834,N_12122);
nand U18158 (N_18158,N_11761,N_12623);
xnor U18159 (N_18159,N_13910,N_14921);
nand U18160 (N_18160,N_14287,N_11770);
and U18161 (N_18161,N_13997,N_13030);
nor U18162 (N_18162,N_14282,N_10900);
nand U18163 (N_18163,N_10595,N_12304);
nor U18164 (N_18164,N_14908,N_11895);
nand U18165 (N_18165,N_10338,N_14389);
nor U18166 (N_18166,N_13463,N_11110);
nand U18167 (N_18167,N_13279,N_13432);
nor U18168 (N_18168,N_13148,N_14688);
nor U18169 (N_18169,N_14790,N_10687);
and U18170 (N_18170,N_13822,N_14035);
or U18171 (N_18171,N_14634,N_12068);
nand U18172 (N_18172,N_13345,N_10046);
or U18173 (N_18173,N_14406,N_14285);
nand U18174 (N_18174,N_12812,N_12206);
nand U18175 (N_18175,N_12854,N_11685);
nor U18176 (N_18176,N_12171,N_13121);
xnor U18177 (N_18177,N_11546,N_12755);
or U18178 (N_18178,N_14224,N_13387);
or U18179 (N_18179,N_14889,N_14243);
nor U18180 (N_18180,N_13513,N_14983);
nor U18181 (N_18181,N_11486,N_10892);
and U18182 (N_18182,N_13170,N_13067);
nor U18183 (N_18183,N_12112,N_14722);
and U18184 (N_18184,N_13802,N_12013);
xor U18185 (N_18185,N_11068,N_12098);
nand U18186 (N_18186,N_10938,N_11237);
or U18187 (N_18187,N_12273,N_12056);
or U18188 (N_18188,N_11045,N_10539);
nor U18189 (N_18189,N_10263,N_10917);
or U18190 (N_18190,N_10487,N_11822);
nor U18191 (N_18191,N_10497,N_13143);
nor U18192 (N_18192,N_13414,N_12847);
or U18193 (N_18193,N_12830,N_13732);
and U18194 (N_18194,N_10628,N_10866);
and U18195 (N_18195,N_14846,N_14507);
nor U18196 (N_18196,N_11979,N_10877);
or U18197 (N_18197,N_12410,N_11993);
and U18198 (N_18198,N_13655,N_11092);
or U18199 (N_18199,N_14920,N_12781);
or U18200 (N_18200,N_12986,N_14233);
xnor U18201 (N_18201,N_14386,N_12484);
or U18202 (N_18202,N_14602,N_14704);
or U18203 (N_18203,N_11127,N_13677);
or U18204 (N_18204,N_13824,N_13401);
xnor U18205 (N_18205,N_14786,N_14055);
or U18206 (N_18206,N_10576,N_10249);
or U18207 (N_18207,N_14801,N_12680);
nand U18208 (N_18208,N_12475,N_12062);
nand U18209 (N_18209,N_12556,N_10675);
nand U18210 (N_18210,N_11785,N_14350);
or U18211 (N_18211,N_13306,N_13023);
and U18212 (N_18212,N_14572,N_14786);
nor U18213 (N_18213,N_12559,N_13903);
nand U18214 (N_18214,N_14851,N_14902);
or U18215 (N_18215,N_11647,N_12735);
nand U18216 (N_18216,N_10483,N_12013);
nor U18217 (N_18217,N_11355,N_11998);
nor U18218 (N_18218,N_10756,N_14157);
xnor U18219 (N_18219,N_12993,N_11588);
nand U18220 (N_18220,N_10289,N_14357);
xor U18221 (N_18221,N_13818,N_11606);
nand U18222 (N_18222,N_13566,N_11989);
nand U18223 (N_18223,N_14351,N_10903);
nor U18224 (N_18224,N_11043,N_10816);
xnor U18225 (N_18225,N_12771,N_14678);
nor U18226 (N_18226,N_10559,N_11093);
or U18227 (N_18227,N_10515,N_13447);
xor U18228 (N_18228,N_10651,N_12620);
nor U18229 (N_18229,N_11019,N_12278);
or U18230 (N_18230,N_12496,N_12273);
or U18231 (N_18231,N_12679,N_14939);
nand U18232 (N_18232,N_14580,N_14511);
or U18233 (N_18233,N_12432,N_12003);
xor U18234 (N_18234,N_12947,N_13386);
or U18235 (N_18235,N_11205,N_14859);
and U18236 (N_18236,N_11234,N_12305);
or U18237 (N_18237,N_14895,N_12498);
and U18238 (N_18238,N_13683,N_10148);
and U18239 (N_18239,N_14986,N_12939);
nor U18240 (N_18240,N_11852,N_11317);
nand U18241 (N_18241,N_12827,N_14405);
and U18242 (N_18242,N_14807,N_10907);
and U18243 (N_18243,N_14254,N_12012);
nor U18244 (N_18244,N_12895,N_10531);
and U18245 (N_18245,N_11094,N_11563);
nor U18246 (N_18246,N_12695,N_13852);
and U18247 (N_18247,N_12849,N_10851);
nor U18248 (N_18248,N_11465,N_11694);
xor U18249 (N_18249,N_12326,N_11663);
and U18250 (N_18250,N_10714,N_12768);
and U18251 (N_18251,N_14191,N_14509);
nand U18252 (N_18252,N_10308,N_13058);
nand U18253 (N_18253,N_13141,N_14162);
nand U18254 (N_18254,N_12662,N_11612);
nand U18255 (N_18255,N_13847,N_14904);
and U18256 (N_18256,N_11532,N_12906);
nand U18257 (N_18257,N_12677,N_12859);
or U18258 (N_18258,N_11092,N_10937);
and U18259 (N_18259,N_11175,N_10300);
nor U18260 (N_18260,N_13196,N_11788);
or U18261 (N_18261,N_10110,N_12120);
and U18262 (N_18262,N_10829,N_11098);
or U18263 (N_18263,N_10618,N_11476);
nand U18264 (N_18264,N_11983,N_10374);
or U18265 (N_18265,N_11088,N_11465);
or U18266 (N_18266,N_12882,N_12845);
xor U18267 (N_18267,N_12335,N_12993);
or U18268 (N_18268,N_14507,N_13510);
xor U18269 (N_18269,N_10430,N_11696);
nand U18270 (N_18270,N_10628,N_13198);
or U18271 (N_18271,N_11799,N_10790);
and U18272 (N_18272,N_14660,N_14714);
or U18273 (N_18273,N_10566,N_10491);
nand U18274 (N_18274,N_12615,N_14854);
nand U18275 (N_18275,N_11076,N_10677);
nor U18276 (N_18276,N_12298,N_11611);
nand U18277 (N_18277,N_14367,N_11661);
or U18278 (N_18278,N_10602,N_11429);
or U18279 (N_18279,N_11897,N_12794);
and U18280 (N_18280,N_13753,N_12725);
nor U18281 (N_18281,N_13320,N_11683);
and U18282 (N_18282,N_12770,N_13071);
and U18283 (N_18283,N_12128,N_11949);
and U18284 (N_18284,N_14196,N_13574);
nor U18285 (N_18285,N_13616,N_12305);
or U18286 (N_18286,N_11555,N_11500);
nand U18287 (N_18287,N_10026,N_14023);
nor U18288 (N_18288,N_10644,N_10341);
xnor U18289 (N_18289,N_13141,N_11000);
and U18290 (N_18290,N_13813,N_12473);
nor U18291 (N_18291,N_12940,N_12552);
nand U18292 (N_18292,N_13443,N_11449);
and U18293 (N_18293,N_14142,N_10303);
nor U18294 (N_18294,N_11670,N_12302);
nand U18295 (N_18295,N_13616,N_10735);
and U18296 (N_18296,N_14471,N_10961);
nand U18297 (N_18297,N_12000,N_12451);
nand U18298 (N_18298,N_13815,N_10538);
or U18299 (N_18299,N_10103,N_11785);
nor U18300 (N_18300,N_12584,N_11044);
nor U18301 (N_18301,N_12178,N_13448);
nand U18302 (N_18302,N_11385,N_13261);
nand U18303 (N_18303,N_13022,N_12540);
xnor U18304 (N_18304,N_13499,N_12780);
xnor U18305 (N_18305,N_14632,N_11668);
or U18306 (N_18306,N_14210,N_11244);
or U18307 (N_18307,N_14043,N_13535);
nor U18308 (N_18308,N_10314,N_12694);
and U18309 (N_18309,N_10548,N_14252);
nor U18310 (N_18310,N_14823,N_12186);
or U18311 (N_18311,N_10323,N_11313);
or U18312 (N_18312,N_14748,N_10888);
and U18313 (N_18313,N_10032,N_14972);
and U18314 (N_18314,N_11846,N_11787);
and U18315 (N_18315,N_12076,N_10400);
and U18316 (N_18316,N_10256,N_10423);
xnor U18317 (N_18317,N_13893,N_12628);
xor U18318 (N_18318,N_14198,N_11573);
nand U18319 (N_18319,N_14332,N_13199);
xnor U18320 (N_18320,N_11125,N_10368);
nor U18321 (N_18321,N_11445,N_12121);
xor U18322 (N_18322,N_14977,N_12419);
and U18323 (N_18323,N_14173,N_13164);
nor U18324 (N_18324,N_12600,N_12450);
nand U18325 (N_18325,N_13541,N_13550);
and U18326 (N_18326,N_13882,N_13514);
nand U18327 (N_18327,N_10662,N_12648);
or U18328 (N_18328,N_10493,N_14322);
nor U18329 (N_18329,N_14202,N_12368);
and U18330 (N_18330,N_12991,N_10749);
and U18331 (N_18331,N_12772,N_11577);
and U18332 (N_18332,N_11820,N_11077);
and U18333 (N_18333,N_13577,N_10636);
or U18334 (N_18334,N_13875,N_12442);
nand U18335 (N_18335,N_11989,N_12899);
xor U18336 (N_18336,N_13307,N_10559);
or U18337 (N_18337,N_11759,N_10932);
nand U18338 (N_18338,N_10120,N_13049);
or U18339 (N_18339,N_10081,N_13122);
xnor U18340 (N_18340,N_12691,N_14013);
and U18341 (N_18341,N_12598,N_14837);
nor U18342 (N_18342,N_12328,N_10666);
and U18343 (N_18343,N_12365,N_12352);
and U18344 (N_18344,N_10073,N_14122);
and U18345 (N_18345,N_10266,N_12944);
and U18346 (N_18346,N_11461,N_12166);
or U18347 (N_18347,N_11249,N_13995);
nor U18348 (N_18348,N_13556,N_12515);
nor U18349 (N_18349,N_14121,N_12055);
nor U18350 (N_18350,N_12827,N_10316);
or U18351 (N_18351,N_13226,N_13372);
nor U18352 (N_18352,N_11092,N_12352);
nor U18353 (N_18353,N_14798,N_13544);
nand U18354 (N_18354,N_12561,N_10363);
nor U18355 (N_18355,N_10278,N_13856);
nor U18356 (N_18356,N_10111,N_14377);
nor U18357 (N_18357,N_14337,N_11782);
or U18358 (N_18358,N_12491,N_12776);
nand U18359 (N_18359,N_14260,N_14522);
and U18360 (N_18360,N_13065,N_11252);
nor U18361 (N_18361,N_13633,N_11920);
nor U18362 (N_18362,N_11066,N_13387);
nor U18363 (N_18363,N_12989,N_13719);
and U18364 (N_18364,N_13077,N_10974);
and U18365 (N_18365,N_14554,N_12888);
or U18366 (N_18366,N_12909,N_12566);
nor U18367 (N_18367,N_13538,N_14990);
nor U18368 (N_18368,N_10537,N_14788);
and U18369 (N_18369,N_10359,N_12546);
or U18370 (N_18370,N_11895,N_11069);
nor U18371 (N_18371,N_10228,N_10189);
or U18372 (N_18372,N_11176,N_10599);
or U18373 (N_18373,N_14222,N_13897);
and U18374 (N_18374,N_12249,N_14899);
and U18375 (N_18375,N_10592,N_12427);
or U18376 (N_18376,N_12685,N_11208);
nor U18377 (N_18377,N_13092,N_11324);
nand U18378 (N_18378,N_14137,N_13880);
nor U18379 (N_18379,N_11126,N_13422);
xnor U18380 (N_18380,N_13239,N_11097);
or U18381 (N_18381,N_12814,N_11221);
nand U18382 (N_18382,N_12828,N_11679);
nand U18383 (N_18383,N_12544,N_11861);
and U18384 (N_18384,N_11688,N_13575);
and U18385 (N_18385,N_14029,N_12925);
nand U18386 (N_18386,N_10111,N_14392);
and U18387 (N_18387,N_11088,N_13885);
nor U18388 (N_18388,N_14023,N_14993);
nand U18389 (N_18389,N_11045,N_13838);
or U18390 (N_18390,N_11096,N_10223);
or U18391 (N_18391,N_12353,N_14103);
or U18392 (N_18392,N_14556,N_12918);
and U18393 (N_18393,N_11498,N_12365);
and U18394 (N_18394,N_11010,N_10709);
nor U18395 (N_18395,N_12813,N_14396);
nor U18396 (N_18396,N_10199,N_12320);
and U18397 (N_18397,N_14929,N_11098);
and U18398 (N_18398,N_12737,N_14992);
and U18399 (N_18399,N_10305,N_14184);
nor U18400 (N_18400,N_14213,N_13012);
nor U18401 (N_18401,N_12991,N_14064);
and U18402 (N_18402,N_14486,N_10184);
nand U18403 (N_18403,N_10779,N_11942);
nand U18404 (N_18404,N_11339,N_11561);
nor U18405 (N_18405,N_13890,N_14707);
or U18406 (N_18406,N_13039,N_12685);
nor U18407 (N_18407,N_14312,N_10255);
and U18408 (N_18408,N_13384,N_13767);
nand U18409 (N_18409,N_12103,N_13221);
nor U18410 (N_18410,N_14495,N_11728);
nor U18411 (N_18411,N_10401,N_10879);
and U18412 (N_18412,N_11976,N_10388);
or U18413 (N_18413,N_13579,N_14193);
xnor U18414 (N_18414,N_11814,N_10443);
or U18415 (N_18415,N_14765,N_13098);
nor U18416 (N_18416,N_13060,N_10421);
xnor U18417 (N_18417,N_11229,N_14020);
nand U18418 (N_18418,N_14496,N_13349);
nor U18419 (N_18419,N_13645,N_13180);
xor U18420 (N_18420,N_10818,N_14781);
nor U18421 (N_18421,N_10197,N_12565);
and U18422 (N_18422,N_13917,N_14306);
and U18423 (N_18423,N_13638,N_10529);
and U18424 (N_18424,N_10229,N_10297);
and U18425 (N_18425,N_12645,N_10877);
or U18426 (N_18426,N_11552,N_13989);
nand U18427 (N_18427,N_14368,N_10247);
nor U18428 (N_18428,N_10147,N_12776);
or U18429 (N_18429,N_14389,N_11319);
nor U18430 (N_18430,N_14500,N_11183);
and U18431 (N_18431,N_10011,N_14256);
and U18432 (N_18432,N_11418,N_12330);
and U18433 (N_18433,N_10075,N_12753);
and U18434 (N_18434,N_14641,N_10884);
xor U18435 (N_18435,N_14838,N_13690);
xnor U18436 (N_18436,N_12218,N_11566);
nor U18437 (N_18437,N_13577,N_14295);
nand U18438 (N_18438,N_13382,N_13787);
nand U18439 (N_18439,N_12835,N_11248);
nor U18440 (N_18440,N_10882,N_10764);
nand U18441 (N_18441,N_11626,N_13213);
and U18442 (N_18442,N_11588,N_11811);
and U18443 (N_18443,N_13673,N_14487);
and U18444 (N_18444,N_14925,N_11373);
or U18445 (N_18445,N_12636,N_14607);
and U18446 (N_18446,N_10870,N_11417);
nand U18447 (N_18447,N_14297,N_10668);
xor U18448 (N_18448,N_14296,N_13314);
and U18449 (N_18449,N_12960,N_14330);
or U18450 (N_18450,N_10910,N_13497);
or U18451 (N_18451,N_10918,N_12677);
nor U18452 (N_18452,N_12892,N_14631);
or U18453 (N_18453,N_10178,N_13384);
nand U18454 (N_18454,N_12160,N_11089);
nand U18455 (N_18455,N_11024,N_11166);
nand U18456 (N_18456,N_13175,N_10872);
nand U18457 (N_18457,N_13947,N_12179);
nand U18458 (N_18458,N_11091,N_14281);
xnor U18459 (N_18459,N_12263,N_12804);
or U18460 (N_18460,N_14639,N_11425);
nor U18461 (N_18461,N_10015,N_12187);
nor U18462 (N_18462,N_12843,N_10990);
nand U18463 (N_18463,N_13331,N_14949);
xnor U18464 (N_18464,N_11351,N_11827);
and U18465 (N_18465,N_11899,N_10394);
and U18466 (N_18466,N_10985,N_10770);
xnor U18467 (N_18467,N_12298,N_12800);
nor U18468 (N_18468,N_14691,N_11866);
and U18469 (N_18469,N_13436,N_10475);
or U18470 (N_18470,N_11329,N_12449);
nand U18471 (N_18471,N_12138,N_13444);
and U18472 (N_18472,N_12474,N_12212);
nor U18473 (N_18473,N_11572,N_10217);
or U18474 (N_18474,N_13433,N_11355);
nand U18475 (N_18475,N_14981,N_13037);
nand U18476 (N_18476,N_11488,N_14236);
xor U18477 (N_18477,N_13654,N_11154);
and U18478 (N_18478,N_10592,N_10868);
xor U18479 (N_18479,N_14905,N_10227);
xnor U18480 (N_18480,N_12657,N_10181);
xor U18481 (N_18481,N_11085,N_10130);
and U18482 (N_18482,N_13076,N_12826);
nor U18483 (N_18483,N_11869,N_13309);
nand U18484 (N_18484,N_11528,N_12559);
nand U18485 (N_18485,N_11002,N_13149);
or U18486 (N_18486,N_12079,N_11720);
and U18487 (N_18487,N_14314,N_13926);
nor U18488 (N_18488,N_11093,N_10528);
nand U18489 (N_18489,N_10092,N_14247);
xnor U18490 (N_18490,N_11591,N_11496);
and U18491 (N_18491,N_13709,N_12003);
or U18492 (N_18492,N_14076,N_13169);
and U18493 (N_18493,N_13307,N_12155);
xnor U18494 (N_18494,N_12343,N_14378);
nor U18495 (N_18495,N_13969,N_10291);
nand U18496 (N_18496,N_12456,N_10317);
nor U18497 (N_18497,N_14701,N_12879);
and U18498 (N_18498,N_12782,N_12513);
and U18499 (N_18499,N_12398,N_14710);
or U18500 (N_18500,N_14042,N_13310);
nand U18501 (N_18501,N_11149,N_12671);
or U18502 (N_18502,N_11294,N_13320);
or U18503 (N_18503,N_12575,N_14851);
and U18504 (N_18504,N_12190,N_14970);
nand U18505 (N_18505,N_12768,N_14876);
nor U18506 (N_18506,N_13821,N_13201);
or U18507 (N_18507,N_12515,N_14056);
xor U18508 (N_18508,N_10820,N_14842);
or U18509 (N_18509,N_14542,N_10562);
nor U18510 (N_18510,N_12332,N_10565);
nor U18511 (N_18511,N_11967,N_10802);
nand U18512 (N_18512,N_13552,N_13238);
and U18513 (N_18513,N_11641,N_10939);
nand U18514 (N_18514,N_14726,N_14261);
xor U18515 (N_18515,N_12928,N_14625);
xor U18516 (N_18516,N_12468,N_14831);
or U18517 (N_18517,N_10243,N_14354);
nor U18518 (N_18518,N_12599,N_14023);
nand U18519 (N_18519,N_11952,N_11605);
nor U18520 (N_18520,N_12767,N_10807);
and U18521 (N_18521,N_12414,N_14623);
or U18522 (N_18522,N_14084,N_12687);
nand U18523 (N_18523,N_11980,N_11713);
or U18524 (N_18524,N_11730,N_10984);
and U18525 (N_18525,N_12762,N_14748);
and U18526 (N_18526,N_14175,N_12585);
nand U18527 (N_18527,N_10427,N_12451);
nand U18528 (N_18528,N_10074,N_13432);
or U18529 (N_18529,N_14534,N_13285);
and U18530 (N_18530,N_10228,N_11273);
nor U18531 (N_18531,N_14532,N_14887);
nor U18532 (N_18532,N_13833,N_11501);
nor U18533 (N_18533,N_11628,N_13835);
or U18534 (N_18534,N_11500,N_14113);
nor U18535 (N_18535,N_11559,N_12776);
or U18536 (N_18536,N_10160,N_12686);
nor U18537 (N_18537,N_12734,N_11503);
or U18538 (N_18538,N_10460,N_11579);
and U18539 (N_18539,N_14604,N_10844);
nor U18540 (N_18540,N_14633,N_11940);
or U18541 (N_18541,N_11244,N_14789);
nor U18542 (N_18542,N_11104,N_13465);
nor U18543 (N_18543,N_14338,N_12440);
nand U18544 (N_18544,N_14820,N_14310);
and U18545 (N_18545,N_10563,N_13055);
or U18546 (N_18546,N_12323,N_13567);
or U18547 (N_18547,N_14903,N_14173);
nand U18548 (N_18548,N_14564,N_10667);
nand U18549 (N_18549,N_11019,N_14288);
or U18550 (N_18550,N_12101,N_10436);
and U18551 (N_18551,N_10442,N_11986);
and U18552 (N_18552,N_10157,N_12632);
xor U18553 (N_18553,N_12894,N_11277);
and U18554 (N_18554,N_13305,N_11422);
and U18555 (N_18555,N_13332,N_14279);
or U18556 (N_18556,N_14053,N_11199);
and U18557 (N_18557,N_11573,N_14312);
and U18558 (N_18558,N_10323,N_10055);
and U18559 (N_18559,N_14337,N_13874);
xnor U18560 (N_18560,N_11822,N_13656);
and U18561 (N_18561,N_13192,N_14084);
nor U18562 (N_18562,N_10877,N_10118);
and U18563 (N_18563,N_10486,N_11179);
nand U18564 (N_18564,N_13826,N_14593);
nor U18565 (N_18565,N_12521,N_13626);
and U18566 (N_18566,N_10744,N_12182);
nor U18567 (N_18567,N_14611,N_12646);
and U18568 (N_18568,N_11538,N_11837);
xor U18569 (N_18569,N_14258,N_10399);
or U18570 (N_18570,N_14097,N_14533);
and U18571 (N_18571,N_12553,N_14258);
nor U18572 (N_18572,N_14638,N_13338);
nor U18573 (N_18573,N_11464,N_10650);
xor U18574 (N_18574,N_10877,N_13200);
nand U18575 (N_18575,N_14762,N_10947);
xor U18576 (N_18576,N_11419,N_11988);
and U18577 (N_18577,N_10884,N_10139);
or U18578 (N_18578,N_10252,N_13025);
or U18579 (N_18579,N_11928,N_14843);
xor U18580 (N_18580,N_10656,N_12559);
and U18581 (N_18581,N_11226,N_10530);
and U18582 (N_18582,N_10869,N_12328);
nor U18583 (N_18583,N_10670,N_13928);
or U18584 (N_18584,N_13775,N_12608);
xnor U18585 (N_18585,N_11256,N_11094);
and U18586 (N_18586,N_14479,N_11829);
and U18587 (N_18587,N_13619,N_13770);
or U18588 (N_18588,N_14723,N_11816);
nand U18589 (N_18589,N_10358,N_10968);
nand U18590 (N_18590,N_10388,N_13802);
or U18591 (N_18591,N_10683,N_14113);
nand U18592 (N_18592,N_13209,N_11711);
and U18593 (N_18593,N_13410,N_12952);
xor U18594 (N_18594,N_10592,N_13547);
or U18595 (N_18595,N_10260,N_11019);
and U18596 (N_18596,N_11665,N_11580);
nand U18597 (N_18597,N_13988,N_13804);
nor U18598 (N_18598,N_14907,N_10909);
nand U18599 (N_18599,N_11636,N_13130);
nor U18600 (N_18600,N_12102,N_12590);
nor U18601 (N_18601,N_10840,N_10826);
or U18602 (N_18602,N_12194,N_14551);
nand U18603 (N_18603,N_13862,N_12447);
or U18604 (N_18604,N_12583,N_14434);
nor U18605 (N_18605,N_11869,N_10339);
or U18606 (N_18606,N_14113,N_13224);
nor U18607 (N_18607,N_10591,N_14348);
nand U18608 (N_18608,N_13907,N_14376);
nor U18609 (N_18609,N_12848,N_11195);
and U18610 (N_18610,N_12785,N_12741);
or U18611 (N_18611,N_11988,N_10455);
xor U18612 (N_18612,N_14909,N_14237);
nor U18613 (N_18613,N_13391,N_14472);
nor U18614 (N_18614,N_14568,N_12354);
nand U18615 (N_18615,N_13518,N_11076);
nor U18616 (N_18616,N_12871,N_12665);
or U18617 (N_18617,N_14795,N_13472);
nor U18618 (N_18618,N_11909,N_11152);
and U18619 (N_18619,N_11334,N_12870);
and U18620 (N_18620,N_11920,N_10272);
nand U18621 (N_18621,N_13034,N_10881);
and U18622 (N_18622,N_13959,N_11905);
nand U18623 (N_18623,N_12787,N_14793);
nor U18624 (N_18624,N_14032,N_13639);
or U18625 (N_18625,N_12733,N_10363);
xnor U18626 (N_18626,N_12942,N_13480);
nand U18627 (N_18627,N_12565,N_12457);
nor U18628 (N_18628,N_14957,N_13999);
and U18629 (N_18629,N_14399,N_11340);
or U18630 (N_18630,N_12707,N_12415);
nor U18631 (N_18631,N_14792,N_12512);
or U18632 (N_18632,N_11381,N_10045);
and U18633 (N_18633,N_13700,N_12933);
nor U18634 (N_18634,N_13374,N_12363);
or U18635 (N_18635,N_12567,N_12263);
or U18636 (N_18636,N_14079,N_10533);
and U18637 (N_18637,N_14034,N_12624);
nand U18638 (N_18638,N_11880,N_10081);
nand U18639 (N_18639,N_10852,N_12588);
and U18640 (N_18640,N_10632,N_10049);
or U18641 (N_18641,N_12938,N_11716);
nand U18642 (N_18642,N_12156,N_10924);
nor U18643 (N_18643,N_14036,N_14012);
or U18644 (N_18644,N_13708,N_11945);
or U18645 (N_18645,N_12125,N_12043);
xor U18646 (N_18646,N_13309,N_13460);
and U18647 (N_18647,N_13555,N_10253);
xnor U18648 (N_18648,N_10120,N_12224);
or U18649 (N_18649,N_10830,N_13901);
or U18650 (N_18650,N_14528,N_14668);
nor U18651 (N_18651,N_12801,N_14528);
nor U18652 (N_18652,N_11629,N_14083);
nor U18653 (N_18653,N_14146,N_12315);
nor U18654 (N_18654,N_14258,N_12729);
nand U18655 (N_18655,N_11620,N_14164);
and U18656 (N_18656,N_12683,N_12930);
and U18657 (N_18657,N_13945,N_10148);
and U18658 (N_18658,N_12859,N_10268);
nand U18659 (N_18659,N_12483,N_14808);
or U18660 (N_18660,N_10096,N_11895);
or U18661 (N_18661,N_11159,N_11771);
or U18662 (N_18662,N_13094,N_10071);
nor U18663 (N_18663,N_12279,N_14529);
nor U18664 (N_18664,N_12718,N_12415);
nor U18665 (N_18665,N_12702,N_11333);
nand U18666 (N_18666,N_11448,N_14986);
nor U18667 (N_18667,N_14444,N_12724);
nand U18668 (N_18668,N_13846,N_14187);
nand U18669 (N_18669,N_12431,N_13599);
nand U18670 (N_18670,N_14268,N_10425);
and U18671 (N_18671,N_12491,N_13934);
nor U18672 (N_18672,N_13334,N_12549);
nor U18673 (N_18673,N_11465,N_14396);
nand U18674 (N_18674,N_14336,N_13448);
xnor U18675 (N_18675,N_13994,N_14402);
and U18676 (N_18676,N_10377,N_12867);
nand U18677 (N_18677,N_14914,N_10127);
xor U18678 (N_18678,N_11696,N_14491);
nor U18679 (N_18679,N_14767,N_13137);
xnor U18680 (N_18680,N_14882,N_14499);
nand U18681 (N_18681,N_10299,N_13540);
or U18682 (N_18682,N_12978,N_14132);
xor U18683 (N_18683,N_13967,N_10355);
nor U18684 (N_18684,N_12803,N_12116);
nor U18685 (N_18685,N_10590,N_14372);
or U18686 (N_18686,N_13073,N_11417);
or U18687 (N_18687,N_14511,N_10785);
and U18688 (N_18688,N_13570,N_10384);
and U18689 (N_18689,N_13094,N_10144);
xnor U18690 (N_18690,N_14349,N_11369);
or U18691 (N_18691,N_13287,N_10260);
nand U18692 (N_18692,N_12321,N_14844);
xor U18693 (N_18693,N_11998,N_14065);
or U18694 (N_18694,N_12104,N_10250);
nor U18695 (N_18695,N_12293,N_10995);
nor U18696 (N_18696,N_10011,N_10271);
xor U18697 (N_18697,N_12175,N_11393);
nand U18698 (N_18698,N_11365,N_12194);
or U18699 (N_18699,N_12350,N_13607);
or U18700 (N_18700,N_13210,N_12521);
and U18701 (N_18701,N_13138,N_12726);
nor U18702 (N_18702,N_13570,N_13737);
and U18703 (N_18703,N_12451,N_14374);
nor U18704 (N_18704,N_10885,N_13158);
nor U18705 (N_18705,N_12753,N_12483);
nand U18706 (N_18706,N_14882,N_12082);
and U18707 (N_18707,N_10126,N_14417);
nor U18708 (N_18708,N_11206,N_12525);
nand U18709 (N_18709,N_11051,N_14419);
or U18710 (N_18710,N_14281,N_10100);
nand U18711 (N_18711,N_14342,N_11156);
nor U18712 (N_18712,N_13465,N_10237);
nand U18713 (N_18713,N_12209,N_13973);
nor U18714 (N_18714,N_14504,N_11716);
nand U18715 (N_18715,N_12773,N_11328);
and U18716 (N_18716,N_10024,N_14918);
and U18717 (N_18717,N_12801,N_13247);
and U18718 (N_18718,N_11476,N_13973);
or U18719 (N_18719,N_10875,N_13269);
and U18720 (N_18720,N_11532,N_11985);
nand U18721 (N_18721,N_10547,N_13365);
xnor U18722 (N_18722,N_11022,N_10030);
and U18723 (N_18723,N_12006,N_10245);
or U18724 (N_18724,N_10810,N_12661);
xor U18725 (N_18725,N_10824,N_12852);
and U18726 (N_18726,N_14040,N_14770);
and U18727 (N_18727,N_14141,N_12186);
nor U18728 (N_18728,N_14782,N_14387);
nand U18729 (N_18729,N_11715,N_13652);
or U18730 (N_18730,N_10646,N_11452);
nor U18731 (N_18731,N_11281,N_11097);
or U18732 (N_18732,N_11966,N_14188);
or U18733 (N_18733,N_11378,N_11956);
and U18734 (N_18734,N_12419,N_12410);
nor U18735 (N_18735,N_13669,N_12581);
and U18736 (N_18736,N_10222,N_10790);
and U18737 (N_18737,N_12057,N_10747);
nor U18738 (N_18738,N_12145,N_10637);
nor U18739 (N_18739,N_12485,N_11923);
nor U18740 (N_18740,N_12974,N_13872);
xnor U18741 (N_18741,N_13409,N_12431);
nand U18742 (N_18742,N_12129,N_12993);
xnor U18743 (N_18743,N_13684,N_12906);
or U18744 (N_18744,N_10170,N_11744);
or U18745 (N_18745,N_12463,N_10133);
or U18746 (N_18746,N_11788,N_12504);
nor U18747 (N_18747,N_11995,N_14836);
xnor U18748 (N_18748,N_12525,N_10091);
nand U18749 (N_18749,N_10880,N_12771);
and U18750 (N_18750,N_12721,N_14289);
or U18751 (N_18751,N_12380,N_13140);
nand U18752 (N_18752,N_11456,N_11290);
or U18753 (N_18753,N_12287,N_10865);
and U18754 (N_18754,N_11998,N_12645);
nor U18755 (N_18755,N_11086,N_13096);
nand U18756 (N_18756,N_13433,N_10812);
or U18757 (N_18757,N_10322,N_11597);
nand U18758 (N_18758,N_14286,N_13945);
or U18759 (N_18759,N_11793,N_10404);
nand U18760 (N_18760,N_10033,N_14796);
xor U18761 (N_18761,N_10842,N_13796);
and U18762 (N_18762,N_13870,N_12015);
or U18763 (N_18763,N_13825,N_14319);
or U18764 (N_18764,N_14682,N_13930);
xor U18765 (N_18765,N_10831,N_14262);
nor U18766 (N_18766,N_14914,N_10064);
nor U18767 (N_18767,N_12385,N_10564);
and U18768 (N_18768,N_10082,N_11699);
nor U18769 (N_18769,N_13229,N_14185);
or U18770 (N_18770,N_10992,N_14419);
and U18771 (N_18771,N_10438,N_12630);
nor U18772 (N_18772,N_12555,N_13651);
nor U18773 (N_18773,N_10017,N_11782);
xor U18774 (N_18774,N_10621,N_12291);
nor U18775 (N_18775,N_11816,N_11689);
or U18776 (N_18776,N_10025,N_11240);
xnor U18777 (N_18777,N_10617,N_10696);
nor U18778 (N_18778,N_14697,N_14515);
and U18779 (N_18779,N_13240,N_13565);
nor U18780 (N_18780,N_13815,N_12596);
nor U18781 (N_18781,N_12842,N_12548);
or U18782 (N_18782,N_12129,N_14484);
and U18783 (N_18783,N_11869,N_12430);
xor U18784 (N_18784,N_14352,N_10631);
and U18785 (N_18785,N_11869,N_12414);
nand U18786 (N_18786,N_14741,N_11140);
and U18787 (N_18787,N_14755,N_10922);
nor U18788 (N_18788,N_10658,N_13784);
nand U18789 (N_18789,N_10884,N_14276);
nand U18790 (N_18790,N_14288,N_13910);
and U18791 (N_18791,N_13681,N_13296);
xor U18792 (N_18792,N_11374,N_13825);
nand U18793 (N_18793,N_10964,N_14942);
or U18794 (N_18794,N_14434,N_10317);
nand U18795 (N_18795,N_13313,N_12293);
nor U18796 (N_18796,N_13372,N_12534);
xor U18797 (N_18797,N_11939,N_14581);
or U18798 (N_18798,N_12361,N_11527);
nand U18799 (N_18799,N_14506,N_12262);
or U18800 (N_18800,N_14044,N_13753);
nor U18801 (N_18801,N_10379,N_13019);
or U18802 (N_18802,N_12220,N_10753);
or U18803 (N_18803,N_13177,N_11591);
nor U18804 (N_18804,N_14589,N_14749);
or U18805 (N_18805,N_12182,N_11684);
nor U18806 (N_18806,N_11333,N_12670);
and U18807 (N_18807,N_11555,N_12319);
or U18808 (N_18808,N_10260,N_12805);
nor U18809 (N_18809,N_14253,N_11954);
xnor U18810 (N_18810,N_10746,N_13630);
and U18811 (N_18811,N_12721,N_13747);
nor U18812 (N_18812,N_14200,N_10756);
and U18813 (N_18813,N_12130,N_10998);
or U18814 (N_18814,N_13252,N_10111);
and U18815 (N_18815,N_10385,N_11789);
or U18816 (N_18816,N_14821,N_13025);
nor U18817 (N_18817,N_13756,N_14778);
or U18818 (N_18818,N_13133,N_12651);
xnor U18819 (N_18819,N_10126,N_11800);
or U18820 (N_18820,N_12796,N_13729);
or U18821 (N_18821,N_11543,N_12973);
and U18822 (N_18822,N_14522,N_13346);
nor U18823 (N_18823,N_10111,N_10350);
or U18824 (N_18824,N_10594,N_12991);
or U18825 (N_18825,N_13553,N_10184);
and U18826 (N_18826,N_14224,N_13412);
nor U18827 (N_18827,N_11484,N_11463);
nor U18828 (N_18828,N_10020,N_12576);
nor U18829 (N_18829,N_12859,N_13397);
and U18830 (N_18830,N_14729,N_10907);
xnor U18831 (N_18831,N_13154,N_12408);
nand U18832 (N_18832,N_11722,N_13398);
or U18833 (N_18833,N_10995,N_12597);
nor U18834 (N_18834,N_11636,N_13639);
and U18835 (N_18835,N_12001,N_13967);
nand U18836 (N_18836,N_11073,N_12352);
and U18837 (N_18837,N_10198,N_13897);
and U18838 (N_18838,N_13471,N_14222);
nor U18839 (N_18839,N_12313,N_12737);
and U18840 (N_18840,N_12152,N_10484);
nand U18841 (N_18841,N_12161,N_11118);
and U18842 (N_18842,N_11771,N_10000);
and U18843 (N_18843,N_11095,N_10021);
or U18844 (N_18844,N_10460,N_14354);
and U18845 (N_18845,N_12734,N_14685);
nor U18846 (N_18846,N_11901,N_14682);
and U18847 (N_18847,N_10309,N_11824);
nor U18848 (N_18848,N_10252,N_11953);
nor U18849 (N_18849,N_12032,N_13989);
nor U18850 (N_18850,N_12662,N_13884);
nor U18851 (N_18851,N_14218,N_12466);
and U18852 (N_18852,N_13576,N_12389);
nor U18853 (N_18853,N_14099,N_12973);
nand U18854 (N_18854,N_10784,N_13224);
nor U18855 (N_18855,N_14853,N_11847);
or U18856 (N_18856,N_12776,N_13330);
and U18857 (N_18857,N_13599,N_12779);
nor U18858 (N_18858,N_12878,N_12982);
nand U18859 (N_18859,N_12676,N_10469);
and U18860 (N_18860,N_11489,N_14084);
and U18861 (N_18861,N_14788,N_12918);
nand U18862 (N_18862,N_14466,N_14763);
or U18863 (N_18863,N_11997,N_11976);
or U18864 (N_18864,N_12567,N_13369);
nor U18865 (N_18865,N_13989,N_14700);
or U18866 (N_18866,N_13938,N_12865);
or U18867 (N_18867,N_14388,N_14701);
nand U18868 (N_18868,N_14096,N_12741);
or U18869 (N_18869,N_11671,N_13337);
nand U18870 (N_18870,N_12925,N_14555);
nand U18871 (N_18871,N_14972,N_13427);
and U18872 (N_18872,N_11458,N_10474);
nor U18873 (N_18873,N_11678,N_14827);
and U18874 (N_18874,N_14100,N_14318);
nand U18875 (N_18875,N_13026,N_11289);
or U18876 (N_18876,N_10915,N_10897);
and U18877 (N_18877,N_12239,N_13155);
nand U18878 (N_18878,N_13356,N_12272);
nand U18879 (N_18879,N_10110,N_14127);
and U18880 (N_18880,N_11578,N_11927);
or U18881 (N_18881,N_14231,N_10407);
nand U18882 (N_18882,N_10576,N_10385);
nor U18883 (N_18883,N_11246,N_14251);
or U18884 (N_18884,N_14558,N_12834);
xnor U18885 (N_18885,N_11068,N_12348);
or U18886 (N_18886,N_11365,N_14509);
and U18887 (N_18887,N_10030,N_10514);
nor U18888 (N_18888,N_13455,N_14587);
nand U18889 (N_18889,N_14054,N_14005);
nor U18890 (N_18890,N_14114,N_12680);
nor U18891 (N_18891,N_10004,N_14927);
and U18892 (N_18892,N_14802,N_12908);
or U18893 (N_18893,N_12769,N_11227);
nor U18894 (N_18894,N_10951,N_13564);
or U18895 (N_18895,N_12435,N_14963);
or U18896 (N_18896,N_14234,N_13404);
or U18897 (N_18897,N_10686,N_13825);
nor U18898 (N_18898,N_12168,N_13000);
and U18899 (N_18899,N_13000,N_12826);
or U18900 (N_18900,N_13251,N_12417);
nand U18901 (N_18901,N_14146,N_12154);
xnor U18902 (N_18902,N_10610,N_14992);
nand U18903 (N_18903,N_11995,N_12860);
nor U18904 (N_18904,N_10531,N_11123);
nor U18905 (N_18905,N_10742,N_14534);
nor U18906 (N_18906,N_11456,N_14662);
nand U18907 (N_18907,N_14933,N_11820);
nor U18908 (N_18908,N_12743,N_14469);
nor U18909 (N_18909,N_11365,N_13208);
nand U18910 (N_18910,N_12560,N_10020);
or U18911 (N_18911,N_10927,N_13119);
and U18912 (N_18912,N_13895,N_12350);
nor U18913 (N_18913,N_10970,N_12892);
nand U18914 (N_18914,N_13119,N_10049);
nor U18915 (N_18915,N_14363,N_13036);
nor U18916 (N_18916,N_14328,N_11300);
nor U18917 (N_18917,N_11376,N_14095);
and U18918 (N_18918,N_12807,N_10992);
and U18919 (N_18919,N_14545,N_14532);
nor U18920 (N_18920,N_12780,N_13899);
xnor U18921 (N_18921,N_12993,N_14857);
nor U18922 (N_18922,N_14366,N_12111);
nor U18923 (N_18923,N_12129,N_13799);
nand U18924 (N_18924,N_14840,N_14759);
nand U18925 (N_18925,N_10077,N_11201);
nand U18926 (N_18926,N_10982,N_12631);
xor U18927 (N_18927,N_12890,N_14731);
and U18928 (N_18928,N_12462,N_11833);
and U18929 (N_18929,N_10564,N_12207);
or U18930 (N_18930,N_13507,N_10453);
or U18931 (N_18931,N_13388,N_10782);
and U18932 (N_18932,N_14397,N_11433);
or U18933 (N_18933,N_11327,N_13370);
xnor U18934 (N_18934,N_13047,N_11571);
and U18935 (N_18935,N_11108,N_12419);
nand U18936 (N_18936,N_13028,N_10503);
or U18937 (N_18937,N_13526,N_14565);
and U18938 (N_18938,N_11823,N_11307);
and U18939 (N_18939,N_12507,N_10976);
nand U18940 (N_18940,N_13843,N_12127);
and U18941 (N_18941,N_12655,N_12360);
nor U18942 (N_18942,N_10360,N_14128);
and U18943 (N_18943,N_12576,N_13304);
and U18944 (N_18944,N_12362,N_10345);
nor U18945 (N_18945,N_10679,N_12122);
nand U18946 (N_18946,N_14550,N_12475);
and U18947 (N_18947,N_12725,N_14795);
or U18948 (N_18948,N_12748,N_13886);
nor U18949 (N_18949,N_14527,N_11839);
nand U18950 (N_18950,N_12255,N_13532);
nand U18951 (N_18951,N_10853,N_14250);
xor U18952 (N_18952,N_12823,N_12895);
nor U18953 (N_18953,N_12953,N_14181);
or U18954 (N_18954,N_10259,N_14616);
and U18955 (N_18955,N_13537,N_14228);
and U18956 (N_18956,N_10687,N_11318);
nand U18957 (N_18957,N_14429,N_10039);
and U18958 (N_18958,N_11990,N_13946);
nand U18959 (N_18959,N_11487,N_11886);
nor U18960 (N_18960,N_13429,N_11009);
or U18961 (N_18961,N_12269,N_12419);
or U18962 (N_18962,N_12255,N_11420);
and U18963 (N_18963,N_11508,N_11570);
nor U18964 (N_18964,N_11721,N_13924);
nand U18965 (N_18965,N_10960,N_10128);
nand U18966 (N_18966,N_14606,N_12559);
nand U18967 (N_18967,N_12447,N_13519);
nand U18968 (N_18968,N_12343,N_12221);
nor U18969 (N_18969,N_10529,N_11910);
and U18970 (N_18970,N_10613,N_14658);
nor U18971 (N_18971,N_12839,N_13277);
xor U18972 (N_18972,N_10103,N_12910);
nor U18973 (N_18973,N_11101,N_13541);
nand U18974 (N_18974,N_10601,N_12412);
nor U18975 (N_18975,N_13299,N_14172);
nor U18976 (N_18976,N_12912,N_10388);
and U18977 (N_18977,N_14022,N_11368);
nand U18978 (N_18978,N_11138,N_13212);
nor U18979 (N_18979,N_14616,N_14019);
nand U18980 (N_18980,N_14558,N_14372);
or U18981 (N_18981,N_14380,N_10595);
nor U18982 (N_18982,N_11797,N_13637);
nor U18983 (N_18983,N_14193,N_14595);
nor U18984 (N_18984,N_13862,N_13014);
or U18985 (N_18985,N_12409,N_12604);
and U18986 (N_18986,N_14123,N_14057);
and U18987 (N_18987,N_14587,N_12585);
nor U18988 (N_18988,N_14651,N_11161);
nor U18989 (N_18989,N_12259,N_12830);
nand U18990 (N_18990,N_12283,N_14533);
and U18991 (N_18991,N_11064,N_14045);
nor U18992 (N_18992,N_10320,N_13196);
or U18993 (N_18993,N_10238,N_11018);
or U18994 (N_18994,N_14779,N_10040);
nand U18995 (N_18995,N_12280,N_13566);
nor U18996 (N_18996,N_13979,N_13829);
or U18997 (N_18997,N_13684,N_10828);
xor U18998 (N_18998,N_10869,N_10863);
or U18999 (N_18999,N_10471,N_13095);
or U19000 (N_19000,N_14905,N_10396);
nand U19001 (N_19001,N_11420,N_14640);
and U19002 (N_19002,N_13529,N_14966);
or U19003 (N_19003,N_11382,N_14912);
nor U19004 (N_19004,N_12252,N_10922);
and U19005 (N_19005,N_10478,N_12953);
or U19006 (N_19006,N_13175,N_10472);
nand U19007 (N_19007,N_14600,N_14361);
and U19008 (N_19008,N_12154,N_14084);
or U19009 (N_19009,N_12001,N_11226);
nand U19010 (N_19010,N_10390,N_12845);
nor U19011 (N_19011,N_14911,N_14549);
nand U19012 (N_19012,N_13945,N_11658);
and U19013 (N_19013,N_13933,N_10248);
and U19014 (N_19014,N_10485,N_10478);
xor U19015 (N_19015,N_13201,N_11127);
or U19016 (N_19016,N_12835,N_13188);
or U19017 (N_19017,N_11225,N_14941);
and U19018 (N_19018,N_11329,N_12974);
xnor U19019 (N_19019,N_12603,N_13741);
and U19020 (N_19020,N_13785,N_14758);
nor U19021 (N_19021,N_13967,N_14082);
or U19022 (N_19022,N_12911,N_13159);
or U19023 (N_19023,N_10646,N_10041);
nand U19024 (N_19024,N_12367,N_14099);
nor U19025 (N_19025,N_12520,N_13408);
nand U19026 (N_19026,N_13462,N_11875);
and U19027 (N_19027,N_13979,N_12683);
or U19028 (N_19028,N_11450,N_10848);
and U19029 (N_19029,N_13229,N_14514);
and U19030 (N_19030,N_11109,N_11384);
or U19031 (N_19031,N_12119,N_11677);
nand U19032 (N_19032,N_10684,N_12359);
and U19033 (N_19033,N_13945,N_14461);
nor U19034 (N_19034,N_14303,N_11394);
nor U19035 (N_19035,N_11387,N_14998);
nor U19036 (N_19036,N_13211,N_13792);
nor U19037 (N_19037,N_13200,N_11490);
and U19038 (N_19038,N_14581,N_12199);
and U19039 (N_19039,N_12474,N_12044);
nor U19040 (N_19040,N_13159,N_14435);
nor U19041 (N_19041,N_11064,N_10315);
nor U19042 (N_19042,N_11193,N_14017);
nor U19043 (N_19043,N_10067,N_12114);
and U19044 (N_19044,N_14842,N_12477);
and U19045 (N_19045,N_14264,N_14041);
and U19046 (N_19046,N_14583,N_14727);
or U19047 (N_19047,N_10511,N_13393);
and U19048 (N_19048,N_10391,N_11847);
nor U19049 (N_19049,N_14162,N_12498);
or U19050 (N_19050,N_10010,N_12644);
or U19051 (N_19051,N_13322,N_10237);
and U19052 (N_19052,N_11657,N_12762);
and U19053 (N_19053,N_12917,N_14806);
xnor U19054 (N_19054,N_13494,N_12861);
nor U19055 (N_19055,N_14577,N_13830);
nand U19056 (N_19056,N_10784,N_12501);
or U19057 (N_19057,N_14087,N_10516);
or U19058 (N_19058,N_13367,N_13077);
or U19059 (N_19059,N_11812,N_11951);
nor U19060 (N_19060,N_11590,N_13661);
or U19061 (N_19061,N_12217,N_14726);
and U19062 (N_19062,N_10557,N_13824);
nand U19063 (N_19063,N_12776,N_10355);
nor U19064 (N_19064,N_13783,N_12824);
and U19065 (N_19065,N_13183,N_11353);
or U19066 (N_19066,N_10205,N_10059);
nand U19067 (N_19067,N_14799,N_10147);
nand U19068 (N_19068,N_11628,N_14627);
nand U19069 (N_19069,N_14019,N_13374);
nand U19070 (N_19070,N_13478,N_11986);
and U19071 (N_19071,N_10994,N_11653);
or U19072 (N_19072,N_10047,N_11948);
and U19073 (N_19073,N_13783,N_12244);
nand U19074 (N_19074,N_10327,N_14236);
or U19075 (N_19075,N_11700,N_11326);
or U19076 (N_19076,N_12082,N_10773);
and U19077 (N_19077,N_11140,N_11942);
and U19078 (N_19078,N_14377,N_10433);
nand U19079 (N_19079,N_10305,N_10269);
nor U19080 (N_19080,N_13476,N_14216);
or U19081 (N_19081,N_12887,N_10652);
nand U19082 (N_19082,N_11665,N_13979);
nand U19083 (N_19083,N_13539,N_13853);
nand U19084 (N_19084,N_13358,N_12868);
nand U19085 (N_19085,N_10205,N_12168);
and U19086 (N_19086,N_10530,N_12952);
or U19087 (N_19087,N_14970,N_11979);
or U19088 (N_19088,N_10304,N_10237);
and U19089 (N_19089,N_10092,N_10435);
or U19090 (N_19090,N_11746,N_13930);
nand U19091 (N_19091,N_12572,N_13285);
nor U19092 (N_19092,N_14317,N_12141);
xnor U19093 (N_19093,N_12220,N_13524);
or U19094 (N_19094,N_13476,N_12896);
nor U19095 (N_19095,N_14058,N_14112);
nor U19096 (N_19096,N_10803,N_13936);
nand U19097 (N_19097,N_11441,N_13691);
or U19098 (N_19098,N_14791,N_13545);
nor U19099 (N_19099,N_12686,N_11113);
xnor U19100 (N_19100,N_10070,N_12428);
or U19101 (N_19101,N_10291,N_12879);
nor U19102 (N_19102,N_11604,N_12988);
or U19103 (N_19103,N_14846,N_10955);
or U19104 (N_19104,N_14231,N_11211);
or U19105 (N_19105,N_14669,N_14048);
nand U19106 (N_19106,N_14168,N_14341);
nor U19107 (N_19107,N_13015,N_10029);
and U19108 (N_19108,N_12957,N_14560);
nand U19109 (N_19109,N_13863,N_13231);
nand U19110 (N_19110,N_10815,N_14950);
nor U19111 (N_19111,N_13819,N_13032);
nor U19112 (N_19112,N_14879,N_14594);
nand U19113 (N_19113,N_14590,N_10545);
or U19114 (N_19114,N_14651,N_12476);
xor U19115 (N_19115,N_14429,N_10435);
nor U19116 (N_19116,N_11745,N_14132);
nor U19117 (N_19117,N_11758,N_13408);
nand U19118 (N_19118,N_13910,N_11005);
or U19119 (N_19119,N_11399,N_13961);
nor U19120 (N_19120,N_10148,N_11809);
nand U19121 (N_19121,N_12164,N_11001);
or U19122 (N_19122,N_13737,N_12171);
nand U19123 (N_19123,N_12421,N_12648);
and U19124 (N_19124,N_12494,N_10894);
or U19125 (N_19125,N_14455,N_13931);
nor U19126 (N_19126,N_12290,N_11888);
nand U19127 (N_19127,N_12077,N_12080);
xor U19128 (N_19128,N_11144,N_11901);
nor U19129 (N_19129,N_12971,N_12541);
or U19130 (N_19130,N_10950,N_14926);
nand U19131 (N_19131,N_14787,N_13172);
nor U19132 (N_19132,N_14695,N_11402);
and U19133 (N_19133,N_14708,N_14844);
nor U19134 (N_19134,N_11778,N_13146);
or U19135 (N_19135,N_10258,N_12058);
or U19136 (N_19136,N_12387,N_10430);
nand U19137 (N_19137,N_11619,N_11756);
or U19138 (N_19138,N_11865,N_10652);
or U19139 (N_19139,N_12506,N_12675);
and U19140 (N_19140,N_11054,N_14023);
and U19141 (N_19141,N_12807,N_14230);
xor U19142 (N_19142,N_10405,N_13368);
nand U19143 (N_19143,N_14178,N_11560);
nand U19144 (N_19144,N_11214,N_12007);
or U19145 (N_19145,N_10428,N_11234);
or U19146 (N_19146,N_13498,N_14407);
and U19147 (N_19147,N_12713,N_12858);
nor U19148 (N_19148,N_12422,N_13765);
nand U19149 (N_19149,N_10587,N_10126);
and U19150 (N_19150,N_12573,N_12284);
or U19151 (N_19151,N_10623,N_11637);
xor U19152 (N_19152,N_10092,N_14036);
or U19153 (N_19153,N_10487,N_10415);
nor U19154 (N_19154,N_13433,N_11840);
or U19155 (N_19155,N_10054,N_11086);
nand U19156 (N_19156,N_12213,N_13955);
or U19157 (N_19157,N_11618,N_14192);
and U19158 (N_19158,N_12921,N_10582);
nor U19159 (N_19159,N_12085,N_12336);
nor U19160 (N_19160,N_14784,N_13875);
or U19161 (N_19161,N_11836,N_12983);
or U19162 (N_19162,N_12054,N_13398);
and U19163 (N_19163,N_13405,N_11705);
xnor U19164 (N_19164,N_14760,N_12428);
nor U19165 (N_19165,N_14723,N_13656);
or U19166 (N_19166,N_14927,N_11808);
and U19167 (N_19167,N_11868,N_12510);
or U19168 (N_19168,N_12243,N_14592);
and U19169 (N_19169,N_11027,N_14314);
nor U19170 (N_19170,N_14411,N_10607);
or U19171 (N_19171,N_10628,N_13524);
and U19172 (N_19172,N_12577,N_14595);
nand U19173 (N_19173,N_10352,N_10517);
or U19174 (N_19174,N_13875,N_10020);
nor U19175 (N_19175,N_12742,N_14748);
nor U19176 (N_19176,N_10594,N_12097);
nor U19177 (N_19177,N_13952,N_12666);
and U19178 (N_19178,N_12306,N_13220);
xor U19179 (N_19179,N_14987,N_12633);
nand U19180 (N_19180,N_12064,N_11991);
nor U19181 (N_19181,N_14580,N_14066);
nand U19182 (N_19182,N_11678,N_11704);
nor U19183 (N_19183,N_13964,N_11421);
nand U19184 (N_19184,N_14281,N_10181);
or U19185 (N_19185,N_10229,N_10330);
nor U19186 (N_19186,N_13378,N_13834);
nor U19187 (N_19187,N_11387,N_11214);
or U19188 (N_19188,N_10399,N_12833);
nand U19189 (N_19189,N_13740,N_11140);
or U19190 (N_19190,N_14274,N_13777);
nand U19191 (N_19191,N_14274,N_12633);
xnor U19192 (N_19192,N_14839,N_11630);
nand U19193 (N_19193,N_10304,N_13899);
nor U19194 (N_19194,N_14248,N_13707);
nand U19195 (N_19195,N_14149,N_13955);
nand U19196 (N_19196,N_11357,N_10327);
or U19197 (N_19197,N_12101,N_14938);
and U19198 (N_19198,N_11257,N_11317);
and U19199 (N_19199,N_12333,N_12406);
nor U19200 (N_19200,N_12833,N_11924);
or U19201 (N_19201,N_10668,N_10878);
or U19202 (N_19202,N_12757,N_11472);
and U19203 (N_19203,N_13846,N_14802);
and U19204 (N_19204,N_13874,N_13870);
nand U19205 (N_19205,N_12889,N_13262);
nand U19206 (N_19206,N_10348,N_13402);
nand U19207 (N_19207,N_10109,N_10176);
or U19208 (N_19208,N_11258,N_11593);
nand U19209 (N_19209,N_14556,N_12527);
nor U19210 (N_19210,N_14506,N_11279);
and U19211 (N_19211,N_11374,N_11653);
and U19212 (N_19212,N_11073,N_11817);
or U19213 (N_19213,N_14308,N_14815);
or U19214 (N_19214,N_10958,N_11170);
or U19215 (N_19215,N_14801,N_10958);
and U19216 (N_19216,N_11846,N_10919);
nand U19217 (N_19217,N_10434,N_10491);
or U19218 (N_19218,N_10375,N_12098);
nor U19219 (N_19219,N_11366,N_13818);
or U19220 (N_19220,N_12898,N_11789);
nand U19221 (N_19221,N_14844,N_12984);
nand U19222 (N_19222,N_10059,N_10731);
and U19223 (N_19223,N_11075,N_13891);
nor U19224 (N_19224,N_11106,N_12066);
xnor U19225 (N_19225,N_12346,N_10772);
or U19226 (N_19226,N_10109,N_11615);
nor U19227 (N_19227,N_11193,N_12619);
or U19228 (N_19228,N_10985,N_13287);
and U19229 (N_19229,N_14715,N_13226);
or U19230 (N_19230,N_13124,N_13149);
xnor U19231 (N_19231,N_11411,N_13239);
nor U19232 (N_19232,N_10424,N_14981);
nand U19233 (N_19233,N_10770,N_12678);
nor U19234 (N_19234,N_12967,N_14627);
nand U19235 (N_19235,N_14399,N_11114);
and U19236 (N_19236,N_14807,N_11757);
xor U19237 (N_19237,N_10447,N_11400);
nand U19238 (N_19238,N_10186,N_11027);
nand U19239 (N_19239,N_13534,N_12678);
nor U19240 (N_19240,N_12727,N_11158);
nor U19241 (N_19241,N_11859,N_12431);
or U19242 (N_19242,N_12780,N_11784);
and U19243 (N_19243,N_13449,N_12495);
nand U19244 (N_19244,N_11656,N_14319);
and U19245 (N_19245,N_10973,N_14052);
or U19246 (N_19246,N_14867,N_14356);
nand U19247 (N_19247,N_12581,N_11024);
nor U19248 (N_19248,N_10249,N_11521);
or U19249 (N_19249,N_10677,N_10652);
and U19250 (N_19250,N_11208,N_13358);
xor U19251 (N_19251,N_10457,N_13718);
nand U19252 (N_19252,N_11661,N_12573);
and U19253 (N_19253,N_12513,N_10224);
and U19254 (N_19254,N_14952,N_10373);
nand U19255 (N_19255,N_11672,N_11797);
and U19256 (N_19256,N_14657,N_11432);
nor U19257 (N_19257,N_12987,N_11287);
or U19258 (N_19258,N_14772,N_10385);
or U19259 (N_19259,N_13000,N_10241);
or U19260 (N_19260,N_11895,N_13552);
nand U19261 (N_19261,N_10283,N_10815);
nor U19262 (N_19262,N_10823,N_12839);
or U19263 (N_19263,N_12424,N_14027);
nor U19264 (N_19264,N_11718,N_11739);
and U19265 (N_19265,N_12520,N_13613);
and U19266 (N_19266,N_14129,N_10373);
xnor U19267 (N_19267,N_11684,N_10955);
nand U19268 (N_19268,N_12991,N_14203);
nor U19269 (N_19269,N_12421,N_11147);
or U19270 (N_19270,N_11049,N_12182);
nor U19271 (N_19271,N_14580,N_10154);
nor U19272 (N_19272,N_12564,N_10395);
nand U19273 (N_19273,N_13160,N_14826);
and U19274 (N_19274,N_11837,N_10343);
and U19275 (N_19275,N_12329,N_11677);
nand U19276 (N_19276,N_14299,N_12624);
nor U19277 (N_19277,N_13074,N_12829);
xnor U19278 (N_19278,N_13811,N_10129);
nand U19279 (N_19279,N_12905,N_12027);
nand U19280 (N_19280,N_14515,N_14973);
or U19281 (N_19281,N_10070,N_14988);
nor U19282 (N_19282,N_13390,N_10585);
nand U19283 (N_19283,N_11503,N_12493);
nand U19284 (N_19284,N_11339,N_13202);
nor U19285 (N_19285,N_12795,N_14128);
and U19286 (N_19286,N_14704,N_14372);
and U19287 (N_19287,N_13540,N_14181);
nand U19288 (N_19288,N_11340,N_12953);
or U19289 (N_19289,N_10923,N_10767);
nand U19290 (N_19290,N_12822,N_10835);
and U19291 (N_19291,N_10067,N_12280);
nor U19292 (N_19292,N_10834,N_12215);
or U19293 (N_19293,N_14605,N_10459);
and U19294 (N_19294,N_12455,N_12749);
and U19295 (N_19295,N_11126,N_14628);
nand U19296 (N_19296,N_14933,N_11977);
and U19297 (N_19297,N_13754,N_12977);
or U19298 (N_19298,N_12243,N_12426);
nor U19299 (N_19299,N_14434,N_10845);
or U19300 (N_19300,N_14357,N_11940);
xor U19301 (N_19301,N_13696,N_11573);
and U19302 (N_19302,N_11484,N_11038);
and U19303 (N_19303,N_12501,N_14129);
and U19304 (N_19304,N_13743,N_11105);
or U19305 (N_19305,N_14831,N_11431);
nand U19306 (N_19306,N_11340,N_11261);
nor U19307 (N_19307,N_10070,N_13618);
nor U19308 (N_19308,N_12172,N_13692);
and U19309 (N_19309,N_12684,N_11384);
nor U19310 (N_19310,N_11231,N_14017);
nand U19311 (N_19311,N_13983,N_10734);
and U19312 (N_19312,N_12201,N_11422);
and U19313 (N_19313,N_11443,N_12962);
nand U19314 (N_19314,N_11863,N_13827);
nand U19315 (N_19315,N_12129,N_13532);
nand U19316 (N_19316,N_14759,N_12363);
nor U19317 (N_19317,N_14984,N_14952);
or U19318 (N_19318,N_11157,N_14388);
nand U19319 (N_19319,N_13188,N_12251);
and U19320 (N_19320,N_12901,N_10701);
or U19321 (N_19321,N_14197,N_10303);
or U19322 (N_19322,N_14718,N_14652);
and U19323 (N_19323,N_11125,N_12427);
and U19324 (N_19324,N_13211,N_13131);
and U19325 (N_19325,N_12549,N_10903);
or U19326 (N_19326,N_11355,N_11049);
xnor U19327 (N_19327,N_13184,N_12220);
xnor U19328 (N_19328,N_14646,N_11159);
or U19329 (N_19329,N_11204,N_14826);
nor U19330 (N_19330,N_12952,N_14429);
nor U19331 (N_19331,N_11837,N_14052);
nor U19332 (N_19332,N_10914,N_12454);
nor U19333 (N_19333,N_13390,N_14252);
or U19334 (N_19334,N_10020,N_13530);
xor U19335 (N_19335,N_14066,N_13917);
or U19336 (N_19336,N_14698,N_11008);
xnor U19337 (N_19337,N_11836,N_11190);
xnor U19338 (N_19338,N_13777,N_10301);
nand U19339 (N_19339,N_13609,N_11703);
nor U19340 (N_19340,N_12837,N_11578);
and U19341 (N_19341,N_12508,N_11707);
xor U19342 (N_19342,N_12157,N_14045);
xor U19343 (N_19343,N_10459,N_14878);
nand U19344 (N_19344,N_12104,N_13339);
or U19345 (N_19345,N_10588,N_13788);
or U19346 (N_19346,N_11212,N_13826);
nand U19347 (N_19347,N_13575,N_13745);
nor U19348 (N_19348,N_12176,N_10097);
or U19349 (N_19349,N_11353,N_13103);
and U19350 (N_19350,N_13458,N_10096);
nor U19351 (N_19351,N_12509,N_11037);
and U19352 (N_19352,N_13656,N_13557);
nor U19353 (N_19353,N_10407,N_12639);
and U19354 (N_19354,N_10710,N_10461);
or U19355 (N_19355,N_14645,N_11874);
xnor U19356 (N_19356,N_10053,N_14620);
or U19357 (N_19357,N_10346,N_11285);
nand U19358 (N_19358,N_10222,N_14450);
and U19359 (N_19359,N_10445,N_12595);
or U19360 (N_19360,N_12224,N_12748);
and U19361 (N_19361,N_10174,N_10658);
nor U19362 (N_19362,N_12048,N_11069);
and U19363 (N_19363,N_10934,N_10952);
nand U19364 (N_19364,N_11242,N_10119);
or U19365 (N_19365,N_14402,N_12595);
nand U19366 (N_19366,N_12803,N_11943);
nand U19367 (N_19367,N_10297,N_10725);
or U19368 (N_19368,N_10089,N_10310);
or U19369 (N_19369,N_10239,N_11396);
and U19370 (N_19370,N_10611,N_13295);
nor U19371 (N_19371,N_12155,N_12710);
or U19372 (N_19372,N_13834,N_11200);
or U19373 (N_19373,N_13838,N_12101);
and U19374 (N_19374,N_10917,N_11802);
and U19375 (N_19375,N_10674,N_13463);
nor U19376 (N_19376,N_13935,N_13908);
nand U19377 (N_19377,N_10963,N_11831);
nand U19378 (N_19378,N_14991,N_14375);
nor U19379 (N_19379,N_11829,N_13382);
nor U19380 (N_19380,N_12093,N_10357);
and U19381 (N_19381,N_14336,N_14198);
xor U19382 (N_19382,N_10312,N_10960);
nand U19383 (N_19383,N_13356,N_12793);
or U19384 (N_19384,N_12124,N_11303);
nor U19385 (N_19385,N_11574,N_13745);
nor U19386 (N_19386,N_10902,N_12122);
nand U19387 (N_19387,N_10130,N_12599);
nor U19388 (N_19388,N_12518,N_10453);
and U19389 (N_19389,N_10889,N_14033);
or U19390 (N_19390,N_12982,N_10571);
or U19391 (N_19391,N_12763,N_12188);
nor U19392 (N_19392,N_11333,N_12749);
nand U19393 (N_19393,N_11952,N_14004);
nand U19394 (N_19394,N_14176,N_11325);
nand U19395 (N_19395,N_14422,N_14002);
nand U19396 (N_19396,N_14307,N_12133);
nor U19397 (N_19397,N_11597,N_13080);
and U19398 (N_19398,N_14176,N_10375);
nor U19399 (N_19399,N_10482,N_13936);
nor U19400 (N_19400,N_14766,N_14238);
and U19401 (N_19401,N_10116,N_11553);
nand U19402 (N_19402,N_14327,N_12183);
or U19403 (N_19403,N_12180,N_10843);
nor U19404 (N_19404,N_10010,N_11207);
and U19405 (N_19405,N_13251,N_10548);
nor U19406 (N_19406,N_14428,N_12746);
and U19407 (N_19407,N_13595,N_14760);
xor U19408 (N_19408,N_14233,N_11256);
nor U19409 (N_19409,N_11140,N_10030);
and U19410 (N_19410,N_14538,N_14326);
and U19411 (N_19411,N_11484,N_13811);
xor U19412 (N_19412,N_13081,N_11028);
and U19413 (N_19413,N_10052,N_11481);
nand U19414 (N_19414,N_14283,N_10137);
or U19415 (N_19415,N_11835,N_13691);
nand U19416 (N_19416,N_14584,N_11570);
nor U19417 (N_19417,N_14846,N_13618);
and U19418 (N_19418,N_12175,N_10544);
and U19419 (N_19419,N_11715,N_12943);
or U19420 (N_19420,N_10430,N_14208);
nor U19421 (N_19421,N_12814,N_13885);
nand U19422 (N_19422,N_13756,N_10437);
nor U19423 (N_19423,N_14183,N_14756);
nand U19424 (N_19424,N_14350,N_12795);
or U19425 (N_19425,N_13698,N_13226);
or U19426 (N_19426,N_10015,N_14928);
xor U19427 (N_19427,N_11983,N_14501);
nor U19428 (N_19428,N_10451,N_11576);
and U19429 (N_19429,N_12146,N_14347);
xor U19430 (N_19430,N_13290,N_12585);
or U19431 (N_19431,N_10388,N_13690);
xor U19432 (N_19432,N_12242,N_12877);
xnor U19433 (N_19433,N_12038,N_12562);
or U19434 (N_19434,N_13322,N_13478);
and U19435 (N_19435,N_12504,N_11692);
nor U19436 (N_19436,N_13785,N_13295);
xnor U19437 (N_19437,N_11320,N_14024);
xor U19438 (N_19438,N_11646,N_11339);
or U19439 (N_19439,N_11086,N_14178);
xnor U19440 (N_19440,N_10942,N_14940);
or U19441 (N_19441,N_10345,N_12505);
nand U19442 (N_19442,N_12358,N_11725);
nor U19443 (N_19443,N_13241,N_13118);
nor U19444 (N_19444,N_14796,N_12051);
and U19445 (N_19445,N_13343,N_11282);
nand U19446 (N_19446,N_13039,N_11870);
or U19447 (N_19447,N_14810,N_12483);
and U19448 (N_19448,N_10862,N_10365);
and U19449 (N_19449,N_11912,N_14053);
nor U19450 (N_19450,N_12457,N_10213);
nand U19451 (N_19451,N_11099,N_12722);
or U19452 (N_19452,N_14142,N_12108);
or U19453 (N_19453,N_11243,N_12420);
xor U19454 (N_19454,N_13464,N_14118);
or U19455 (N_19455,N_13489,N_11869);
and U19456 (N_19456,N_11723,N_11112);
or U19457 (N_19457,N_10388,N_14973);
or U19458 (N_19458,N_14908,N_12321);
nand U19459 (N_19459,N_11550,N_12371);
nand U19460 (N_19460,N_12642,N_12346);
or U19461 (N_19461,N_14647,N_13140);
nand U19462 (N_19462,N_10249,N_13192);
nor U19463 (N_19463,N_11307,N_11054);
nand U19464 (N_19464,N_12750,N_10668);
or U19465 (N_19465,N_13540,N_12235);
or U19466 (N_19466,N_13817,N_14110);
or U19467 (N_19467,N_10442,N_14441);
nand U19468 (N_19468,N_11454,N_10835);
nor U19469 (N_19469,N_11981,N_10475);
or U19470 (N_19470,N_11440,N_10687);
nand U19471 (N_19471,N_11208,N_10496);
or U19472 (N_19472,N_11568,N_13367);
nand U19473 (N_19473,N_12656,N_12234);
nor U19474 (N_19474,N_14149,N_14369);
xor U19475 (N_19475,N_13351,N_10780);
nand U19476 (N_19476,N_14551,N_14123);
and U19477 (N_19477,N_11751,N_11384);
nor U19478 (N_19478,N_11365,N_12186);
and U19479 (N_19479,N_10923,N_12676);
and U19480 (N_19480,N_13429,N_12329);
nor U19481 (N_19481,N_12877,N_12845);
nand U19482 (N_19482,N_13016,N_12463);
or U19483 (N_19483,N_12323,N_14193);
or U19484 (N_19484,N_14457,N_12892);
and U19485 (N_19485,N_13651,N_14778);
nand U19486 (N_19486,N_11903,N_11878);
nand U19487 (N_19487,N_11382,N_13971);
nor U19488 (N_19488,N_11046,N_14136);
or U19489 (N_19489,N_14234,N_13088);
nand U19490 (N_19490,N_14108,N_12084);
and U19491 (N_19491,N_13327,N_11478);
nand U19492 (N_19492,N_13768,N_12750);
and U19493 (N_19493,N_10487,N_10176);
nand U19494 (N_19494,N_14727,N_10325);
or U19495 (N_19495,N_11405,N_10070);
nor U19496 (N_19496,N_10031,N_13007);
and U19497 (N_19497,N_12851,N_14376);
and U19498 (N_19498,N_10459,N_10167);
nand U19499 (N_19499,N_11952,N_12521);
and U19500 (N_19500,N_10708,N_12556);
xor U19501 (N_19501,N_14755,N_11603);
nor U19502 (N_19502,N_13706,N_10244);
nor U19503 (N_19503,N_13381,N_10112);
nand U19504 (N_19504,N_11388,N_12414);
nand U19505 (N_19505,N_13402,N_14258);
and U19506 (N_19506,N_11655,N_10242);
and U19507 (N_19507,N_14550,N_11699);
or U19508 (N_19508,N_12401,N_10130);
and U19509 (N_19509,N_14914,N_10114);
nand U19510 (N_19510,N_12238,N_12107);
nand U19511 (N_19511,N_12849,N_14912);
and U19512 (N_19512,N_10203,N_12361);
or U19513 (N_19513,N_12915,N_10567);
or U19514 (N_19514,N_14967,N_14910);
xnor U19515 (N_19515,N_12297,N_12982);
or U19516 (N_19516,N_10314,N_13688);
nor U19517 (N_19517,N_14412,N_13253);
or U19518 (N_19518,N_11809,N_12666);
nor U19519 (N_19519,N_11169,N_12014);
and U19520 (N_19520,N_10631,N_14182);
or U19521 (N_19521,N_10811,N_11482);
or U19522 (N_19522,N_12546,N_14152);
and U19523 (N_19523,N_10051,N_11756);
xor U19524 (N_19524,N_13411,N_14247);
nand U19525 (N_19525,N_10173,N_12469);
and U19526 (N_19526,N_10321,N_14329);
and U19527 (N_19527,N_12199,N_11414);
xor U19528 (N_19528,N_14106,N_13103);
xor U19529 (N_19529,N_10068,N_14819);
and U19530 (N_19530,N_13406,N_13169);
nor U19531 (N_19531,N_14233,N_12152);
and U19532 (N_19532,N_12354,N_12822);
nor U19533 (N_19533,N_10929,N_14883);
nand U19534 (N_19534,N_14246,N_12085);
xnor U19535 (N_19535,N_12321,N_10607);
and U19536 (N_19536,N_14831,N_11652);
or U19537 (N_19537,N_12648,N_14775);
or U19538 (N_19538,N_13130,N_11953);
nand U19539 (N_19539,N_13328,N_13511);
nor U19540 (N_19540,N_14374,N_13210);
nand U19541 (N_19541,N_14059,N_14139);
and U19542 (N_19542,N_11007,N_13467);
nor U19543 (N_19543,N_12929,N_13438);
nand U19544 (N_19544,N_11047,N_10926);
and U19545 (N_19545,N_13019,N_10851);
or U19546 (N_19546,N_13394,N_12004);
nand U19547 (N_19547,N_14021,N_12746);
and U19548 (N_19548,N_10126,N_14447);
and U19549 (N_19549,N_11153,N_14165);
or U19550 (N_19550,N_10988,N_13001);
or U19551 (N_19551,N_11335,N_14222);
nor U19552 (N_19552,N_14572,N_11643);
nor U19553 (N_19553,N_14516,N_10585);
nor U19554 (N_19554,N_14327,N_14105);
and U19555 (N_19555,N_13135,N_13957);
nand U19556 (N_19556,N_10178,N_13507);
and U19557 (N_19557,N_11583,N_13708);
and U19558 (N_19558,N_13309,N_14089);
or U19559 (N_19559,N_13908,N_14742);
or U19560 (N_19560,N_14763,N_11894);
nand U19561 (N_19561,N_11097,N_13546);
or U19562 (N_19562,N_11854,N_12847);
or U19563 (N_19563,N_14069,N_14163);
nor U19564 (N_19564,N_11468,N_14123);
or U19565 (N_19565,N_13201,N_12955);
nor U19566 (N_19566,N_12956,N_12759);
nor U19567 (N_19567,N_13496,N_14483);
nand U19568 (N_19568,N_14229,N_14447);
nor U19569 (N_19569,N_11570,N_12507);
nand U19570 (N_19570,N_10256,N_11980);
nand U19571 (N_19571,N_10595,N_12850);
nand U19572 (N_19572,N_13306,N_12105);
and U19573 (N_19573,N_14002,N_13567);
nor U19574 (N_19574,N_12458,N_10081);
nor U19575 (N_19575,N_14075,N_10527);
nand U19576 (N_19576,N_10442,N_12653);
and U19577 (N_19577,N_14874,N_12322);
or U19578 (N_19578,N_10199,N_11928);
and U19579 (N_19579,N_10198,N_12116);
xor U19580 (N_19580,N_13755,N_12178);
or U19581 (N_19581,N_14735,N_14947);
and U19582 (N_19582,N_11026,N_12201);
and U19583 (N_19583,N_10056,N_14648);
nor U19584 (N_19584,N_12432,N_11349);
and U19585 (N_19585,N_10365,N_11893);
nand U19586 (N_19586,N_12132,N_14759);
xor U19587 (N_19587,N_14394,N_14033);
or U19588 (N_19588,N_13259,N_14802);
nor U19589 (N_19589,N_14964,N_12596);
or U19590 (N_19590,N_13671,N_12003);
and U19591 (N_19591,N_11586,N_11843);
nand U19592 (N_19592,N_10673,N_13508);
nor U19593 (N_19593,N_13517,N_10785);
and U19594 (N_19594,N_13466,N_10047);
and U19595 (N_19595,N_13381,N_12660);
nand U19596 (N_19596,N_11119,N_10113);
nand U19597 (N_19597,N_11419,N_12379);
nand U19598 (N_19598,N_13013,N_11882);
nor U19599 (N_19599,N_11951,N_12182);
and U19600 (N_19600,N_14408,N_13786);
nor U19601 (N_19601,N_11608,N_14853);
nand U19602 (N_19602,N_10970,N_10063);
nor U19603 (N_19603,N_12704,N_14684);
nor U19604 (N_19604,N_10533,N_13841);
nor U19605 (N_19605,N_14393,N_13643);
nand U19606 (N_19606,N_10136,N_10397);
or U19607 (N_19607,N_11590,N_11552);
nor U19608 (N_19608,N_11525,N_14372);
or U19609 (N_19609,N_13328,N_13390);
or U19610 (N_19610,N_13265,N_13660);
or U19611 (N_19611,N_12816,N_10813);
nor U19612 (N_19612,N_12404,N_10913);
or U19613 (N_19613,N_13692,N_13300);
and U19614 (N_19614,N_12450,N_13409);
or U19615 (N_19615,N_11975,N_12114);
and U19616 (N_19616,N_12906,N_11075);
nand U19617 (N_19617,N_13167,N_14820);
nor U19618 (N_19618,N_11388,N_11853);
nand U19619 (N_19619,N_11532,N_12414);
and U19620 (N_19620,N_13030,N_11229);
xnor U19621 (N_19621,N_12415,N_10555);
or U19622 (N_19622,N_11180,N_13101);
or U19623 (N_19623,N_13148,N_14666);
nand U19624 (N_19624,N_11243,N_11267);
or U19625 (N_19625,N_14137,N_11355);
nor U19626 (N_19626,N_12879,N_12957);
or U19627 (N_19627,N_12837,N_12783);
nand U19628 (N_19628,N_13134,N_10718);
nand U19629 (N_19629,N_10415,N_11810);
or U19630 (N_19630,N_10830,N_13977);
nor U19631 (N_19631,N_11612,N_13725);
nor U19632 (N_19632,N_11533,N_13124);
nor U19633 (N_19633,N_12970,N_10820);
and U19634 (N_19634,N_10148,N_13659);
nand U19635 (N_19635,N_11062,N_12501);
xor U19636 (N_19636,N_13708,N_12953);
nand U19637 (N_19637,N_14521,N_11109);
nand U19638 (N_19638,N_13922,N_14520);
and U19639 (N_19639,N_12041,N_11653);
or U19640 (N_19640,N_14798,N_10896);
and U19641 (N_19641,N_13740,N_13196);
and U19642 (N_19642,N_12400,N_14371);
xor U19643 (N_19643,N_13178,N_13855);
or U19644 (N_19644,N_14666,N_11112);
and U19645 (N_19645,N_11778,N_14573);
nor U19646 (N_19646,N_13029,N_12030);
nand U19647 (N_19647,N_12920,N_13849);
nor U19648 (N_19648,N_13637,N_10921);
nor U19649 (N_19649,N_10515,N_10715);
nand U19650 (N_19650,N_14053,N_12710);
nor U19651 (N_19651,N_10023,N_10994);
nor U19652 (N_19652,N_13842,N_14366);
and U19653 (N_19653,N_10366,N_10516);
or U19654 (N_19654,N_12505,N_10760);
xor U19655 (N_19655,N_12534,N_14393);
xnor U19656 (N_19656,N_12773,N_10627);
nor U19657 (N_19657,N_10831,N_11987);
nor U19658 (N_19658,N_11032,N_10697);
nor U19659 (N_19659,N_13034,N_11734);
or U19660 (N_19660,N_11796,N_10359);
or U19661 (N_19661,N_10754,N_14552);
and U19662 (N_19662,N_12728,N_12200);
xnor U19663 (N_19663,N_14561,N_12152);
nor U19664 (N_19664,N_13255,N_12216);
xor U19665 (N_19665,N_12644,N_10970);
xnor U19666 (N_19666,N_10514,N_11694);
or U19667 (N_19667,N_12562,N_12718);
nor U19668 (N_19668,N_12986,N_10232);
nand U19669 (N_19669,N_14682,N_12745);
or U19670 (N_19670,N_12297,N_10281);
nor U19671 (N_19671,N_10058,N_13161);
or U19672 (N_19672,N_11883,N_10361);
nor U19673 (N_19673,N_14485,N_10930);
and U19674 (N_19674,N_12117,N_10579);
or U19675 (N_19675,N_12467,N_11128);
nand U19676 (N_19676,N_10006,N_12397);
nand U19677 (N_19677,N_10932,N_14220);
or U19678 (N_19678,N_12586,N_12520);
nand U19679 (N_19679,N_14678,N_13361);
or U19680 (N_19680,N_14517,N_11217);
or U19681 (N_19681,N_10638,N_13327);
nor U19682 (N_19682,N_11216,N_11763);
nand U19683 (N_19683,N_13101,N_11758);
nand U19684 (N_19684,N_10367,N_14525);
xnor U19685 (N_19685,N_12920,N_12603);
nand U19686 (N_19686,N_11229,N_12425);
and U19687 (N_19687,N_10184,N_12323);
or U19688 (N_19688,N_14409,N_14283);
or U19689 (N_19689,N_13535,N_11814);
nor U19690 (N_19690,N_14737,N_14042);
or U19691 (N_19691,N_11833,N_10050);
nor U19692 (N_19692,N_13384,N_13261);
xnor U19693 (N_19693,N_10365,N_14577);
and U19694 (N_19694,N_11622,N_13943);
nor U19695 (N_19695,N_13954,N_14028);
and U19696 (N_19696,N_12222,N_13235);
and U19697 (N_19697,N_10749,N_12133);
or U19698 (N_19698,N_11295,N_14540);
or U19699 (N_19699,N_10159,N_12396);
nand U19700 (N_19700,N_13271,N_10983);
and U19701 (N_19701,N_14188,N_11586);
and U19702 (N_19702,N_14266,N_14024);
and U19703 (N_19703,N_14759,N_14279);
or U19704 (N_19704,N_11091,N_11840);
xor U19705 (N_19705,N_13784,N_12870);
nand U19706 (N_19706,N_12671,N_12601);
nor U19707 (N_19707,N_12240,N_13206);
and U19708 (N_19708,N_13424,N_13639);
nand U19709 (N_19709,N_11042,N_11102);
nand U19710 (N_19710,N_12687,N_14292);
or U19711 (N_19711,N_10609,N_14012);
xor U19712 (N_19712,N_14476,N_13489);
nand U19713 (N_19713,N_14998,N_11984);
nor U19714 (N_19714,N_11825,N_11338);
nand U19715 (N_19715,N_14650,N_10033);
or U19716 (N_19716,N_12472,N_10982);
nand U19717 (N_19717,N_13529,N_10907);
nor U19718 (N_19718,N_13771,N_12341);
nor U19719 (N_19719,N_12974,N_14467);
nor U19720 (N_19720,N_11883,N_11205);
or U19721 (N_19721,N_13801,N_14338);
xor U19722 (N_19722,N_11843,N_14530);
or U19723 (N_19723,N_13752,N_11745);
nand U19724 (N_19724,N_11293,N_11423);
xor U19725 (N_19725,N_12489,N_14363);
nand U19726 (N_19726,N_10730,N_11787);
or U19727 (N_19727,N_13675,N_14837);
nor U19728 (N_19728,N_14043,N_14384);
or U19729 (N_19729,N_12888,N_10510);
nand U19730 (N_19730,N_12032,N_10072);
xnor U19731 (N_19731,N_13071,N_13724);
nor U19732 (N_19732,N_13227,N_11113);
nor U19733 (N_19733,N_11205,N_10795);
nor U19734 (N_19734,N_14133,N_13289);
and U19735 (N_19735,N_14493,N_10358);
or U19736 (N_19736,N_11515,N_10579);
nor U19737 (N_19737,N_10833,N_13426);
xor U19738 (N_19738,N_10122,N_12501);
and U19739 (N_19739,N_10397,N_11731);
nand U19740 (N_19740,N_13933,N_14569);
and U19741 (N_19741,N_11243,N_13830);
and U19742 (N_19742,N_12883,N_11604);
or U19743 (N_19743,N_13633,N_13783);
nor U19744 (N_19744,N_14743,N_12156);
and U19745 (N_19745,N_12804,N_12192);
or U19746 (N_19746,N_14151,N_10784);
or U19747 (N_19747,N_11660,N_11420);
xor U19748 (N_19748,N_14656,N_11984);
nor U19749 (N_19749,N_11882,N_10053);
nor U19750 (N_19750,N_12693,N_11002);
nand U19751 (N_19751,N_12801,N_11513);
nor U19752 (N_19752,N_12658,N_12058);
nand U19753 (N_19753,N_12173,N_11285);
xor U19754 (N_19754,N_14263,N_10487);
and U19755 (N_19755,N_10317,N_10098);
and U19756 (N_19756,N_11487,N_12801);
nand U19757 (N_19757,N_11890,N_10461);
nand U19758 (N_19758,N_11786,N_14203);
nand U19759 (N_19759,N_11550,N_11925);
nand U19760 (N_19760,N_12107,N_13054);
nand U19761 (N_19761,N_12683,N_11271);
and U19762 (N_19762,N_12867,N_14028);
or U19763 (N_19763,N_13867,N_13826);
nand U19764 (N_19764,N_10060,N_11510);
and U19765 (N_19765,N_14490,N_10990);
and U19766 (N_19766,N_13908,N_14383);
or U19767 (N_19767,N_10967,N_14419);
nor U19768 (N_19768,N_14947,N_14270);
and U19769 (N_19769,N_14651,N_10944);
and U19770 (N_19770,N_14824,N_13155);
and U19771 (N_19771,N_10275,N_10889);
and U19772 (N_19772,N_14755,N_10730);
nand U19773 (N_19773,N_14147,N_12358);
xnor U19774 (N_19774,N_13050,N_13257);
and U19775 (N_19775,N_11622,N_14082);
and U19776 (N_19776,N_13627,N_10475);
xor U19777 (N_19777,N_10687,N_13133);
nand U19778 (N_19778,N_10839,N_13908);
nor U19779 (N_19779,N_13223,N_11823);
nor U19780 (N_19780,N_10067,N_12642);
or U19781 (N_19781,N_10872,N_13133);
or U19782 (N_19782,N_10720,N_13856);
nand U19783 (N_19783,N_13504,N_14241);
xor U19784 (N_19784,N_13223,N_13384);
nor U19785 (N_19785,N_10751,N_12678);
nand U19786 (N_19786,N_14371,N_11705);
nand U19787 (N_19787,N_10011,N_12073);
or U19788 (N_19788,N_14740,N_14705);
nor U19789 (N_19789,N_11714,N_11672);
nor U19790 (N_19790,N_13005,N_11557);
or U19791 (N_19791,N_10060,N_14006);
nor U19792 (N_19792,N_11578,N_13270);
or U19793 (N_19793,N_10493,N_12445);
or U19794 (N_19794,N_14839,N_10213);
nor U19795 (N_19795,N_10192,N_10330);
or U19796 (N_19796,N_12771,N_12667);
and U19797 (N_19797,N_10831,N_11596);
or U19798 (N_19798,N_14544,N_14548);
nor U19799 (N_19799,N_13799,N_10411);
xnor U19800 (N_19800,N_13802,N_14148);
or U19801 (N_19801,N_13170,N_14484);
or U19802 (N_19802,N_11495,N_14566);
and U19803 (N_19803,N_13039,N_10018);
nand U19804 (N_19804,N_11666,N_14189);
nand U19805 (N_19805,N_10855,N_12783);
or U19806 (N_19806,N_10826,N_14047);
xnor U19807 (N_19807,N_14579,N_13258);
and U19808 (N_19808,N_12584,N_14252);
nor U19809 (N_19809,N_12771,N_13766);
nand U19810 (N_19810,N_10965,N_14461);
and U19811 (N_19811,N_10771,N_14382);
xor U19812 (N_19812,N_14604,N_14965);
or U19813 (N_19813,N_12813,N_14994);
or U19814 (N_19814,N_12078,N_11097);
nand U19815 (N_19815,N_11468,N_12699);
or U19816 (N_19816,N_10935,N_14028);
nand U19817 (N_19817,N_14156,N_10476);
nor U19818 (N_19818,N_10013,N_14871);
or U19819 (N_19819,N_13834,N_12131);
xor U19820 (N_19820,N_10089,N_14367);
nor U19821 (N_19821,N_10010,N_13954);
xor U19822 (N_19822,N_11203,N_13114);
nor U19823 (N_19823,N_13433,N_10873);
xor U19824 (N_19824,N_11656,N_11618);
or U19825 (N_19825,N_13217,N_10853);
or U19826 (N_19826,N_14308,N_12514);
and U19827 (N_19827,N_13511,N_12081);
or U19828 (N_19828,N_14647,N_12799);
nor U19829 (N_19829,N_11534,N_12304);
and U19830 (N_19830,N_10012,N_13693);
xor U19831 (N_19831,N_14458,N_10357);
and U19832 (N_19832,N_14242,N_14435);
and U19833 (N_19833,N_12461,N_14203);
or U19834 (N_19834,N_13937,N_10678);
nor U19835 (N_19835,N_11693,N_13695);
and U19836 (N_19836,N_11697,N_14253);
and U19837 (N_19837,N_13660,N_11654);
nand U19838 (N_19838,N_14221,N_14950);
and U19839 (N_19839,N_11433,N_11945);
nor U19840 (N_19840,N_14439,N_10875);
and U19841 (N_19841,N_13499,N_14844);
and U19842 (N_19842,N_13804,N_11621);
or U19843 (N_19843,N_13797,N_11134);
or U19844 (N_19844,N_14847,N_14285);
xnor U19845 (N_19845,N_11736,N_13326);
xor U19846 (N_19846,N_13650,N_14680);
nand U19847 (N_19847,N_11437,N_11585);
nand U19848 (N_19848,N_13452,N_12332);
nor U19849 (N_19849,N_14049,N_14447);
nor U19850 (N_19850,N_10571,N_13621);
nand U19851 (N_19851,N_12782,N_11505);
and U19852 (N_19852,N_12648,N_12546);
xnor U19853 (N_19853,N_14182,N_11332);
nand U19854 (N_19854,N_12621,N_10489);
nor U19855 (N_19855,N_10846,N_13421);
nand U19856 (N_19856,N_11850,N_14075);
or U19857 (N_19857,N_11963,N_13928);
or U19858 (N_19858,N_11758,N_14212);
and U19859 (N_19859,N_13556,N_11370);
xor U19860 (N_19860,N_14155,N_13258);
or U19861 (N_19861,N_12617,N_14353);
or U19862 (N_19862,N_13604,N_11580);
xor U19863 (N_19863,N_11930,N_11508);
nand U19864 (N_19864,N_11961,N_11200);
or U19865 (N_19865,N_10091,N_11147);
and U19866 (N_19866,N_14577,N_10835);
xor U19867 (N_19867,N_10188,N_11087);
and U19868 (N_19868,N_14692,N_11133);
or U19869 (N_19869,N_10080,N_14648);
or U19870 (N_19870,N_10266,N_13956);
or U19871 (N_19871,N_14356,N_13492);
nor U19872 (N_19872,N_13762,N_11487);
nor U19873 (N_19873,N_13052,N_14120);
and U19874 (N_19874,N_13241,N_10387);
nor U19875 (N_19875,N_10009,N_14258);
or U19876 (N_19876,N_14275,N_12818);
or U19877 (N_19877,N_14901,N_11432);
or U19878 (N_19878,N_11952,N_12190);
nand U19879 (N_19879,N_12697,N_12341);
and U19880 (N_19880,N_10912,N_10735);
or U19881 (N_19881,N_10964,N_10841);
and U19882 (N_19882,N_14288,N_10924);
and U19883 (N_19883,N_13877,N_10949);
nor U19884 (N_19884,N_13114,N_14656);
or U19885 (N_19885,N_14450,N_12584);
xor U19886 (N_19886,N_12811,N_11024);
or U19887 (N_19887,N_11191,N_10073);
xnor U19888 (N_19888,N_10428,N_14673);
or U19889 (N_19889,N_12930,N_14492);
or U19890 (N_19890,N_12714,N_10668);
or U19891 (N_19891,N_14811,N_13636);
xnor U19892 (N_19892,N_12961,N_13179);
nand U19893 (N_19893,N_14339,N_12790);
nand U19894 (N_19894,N_14592,N_13445);
nor U19895 (N_19895,N_14402,N_14572);
nand U19896 (N_19896,N_13657,N_14109);
or U19897 (N_19897,N_11456,N_12168);
and U19898 (N_19898,N_13859,N_11299);
nand U19899 (N_19899,N_13480,N_13022);
or U19900 (N_19900,N_12087,N_11136);
and U19901 (N_19901,N_13755,N_11528);
nand U19902 (N_19902,N_13720,N_14614);
and U19903 (N_19903,N_12816,N_12667);
nand U19904 (N_19904,N_10397,N_11567);
or U19905 (N_19905,N_13408,N_13126);
and U19906 (N_19906,N_11556,N_10580);
or U19907 (N_19907,N_12902,N_12522);
nor U19908 (N_19908,N_13113,N_13102);
nor U19909 (N_19909,N_14617,N_13007);
nand U19910 (N_19910,N_13795,N_13091);
and U19911 (N_19911,N_13064,N_13753);
and U19912 (N_19912,N_10967,N_11283);
or U19913 (N_19913,N_12077,N_14030);
nor U19914 (N_19914,N_13420,N_12960);
or U19915 (N_19915,N_11834,N_11116);
xnor U19916 (N_19916,N_13520,N_14071);
and U19917 (N_19917,N_13652,N_12274);
nand U19918 (N_19918,N_10121,N_11416);
nand U19919 (N_19919,N_14232,N_13792);
xor U19920 (N_19920,N_10677,N_12558);
and U19921 (N_19921,N_14730,N_10304);
nor U19922 (N_19922,N_12144,N_12229);
or U19923 (N_19923,N_14616,N_12764);
and U19924 (N_19924,N_12523,N_10733);
nor U19925 (N_19925,N_12754,N_12346);
nor U19926 (N_19926,N_12126,N_13407);
nand U19927 (N_19927,N_11386,N_13953);
xor U19928 (N_19928,N_13833,N_10808);
nor U19929 (N_19929,N_13693,N_11952);
nor U19930 (N_19930,N_14646,N_13593);
or U19931 (N_19931,N_12122,N_10618);
or U19932 (N_19932,N_11374,N_11444);
nor U19933 (N_19933,N_14855,N_10671);
or U19934 (N_19934,N_11293,N_13817);
nor U19935 (N_19935,N_12883,N_12092);
xor U19936 (N_19936,N_11302,N_12161);
and U19937 (N_19937,N_13176,N_14135);
nor U19938 (N_19938,N_12789,N_12477);
xnor U19939 (N_19939,N_12767,N_12382);
and U19940 (N_19940,N_12215,N_11499);
nor U19941 (N_19941,N_10758,N_12466);
nand U19942 (N_19942,N_13062,N_12001);
nor U19943 (N_19943,N_12689,N_11687);
and U19944 (N_19944,N_12955,N_10471);
nor U19945 (N_19945,N_12577,N_10641);
or U19946 (N_19946,N_12425,N_10312);
nor U19947 (N_19947,N_12536,N_14231);
xnor U19948 (N_19948,N_14458,N_10836);
nor U19949 (N_19949,N_12598,N_13027);
and U19950 (N_19950,N_10626,N_10956);
nor U19951 (N_19951,N_13580,N_10126);
nor U19952 (N_19952,N_12681,N_11580);
or U19953 (N_19953,N_11457,N_14651);
and U19954 (N_19954,N_11300,N_11949);
and U19955 (N_19955,N_10994,N_11168);
and U19956 (N_19956,N_10461,N_12246);
and U19957 (N_19957,N_13202,N_13745);
or U19958 (N_19958,N_10336,N_13967);
nor U19959 (N_19959,N_10233,N_12093);
and U19960 (N_19960,N_13887,N_13776);
xor U19961 (N_19961,N_11864,N_13293);
nor U19962 (N_19962,N_12057,N_13060);
nand U19963 (N_19963,N_12979,N_12840);
and U19964 (N_19964,N_13748,N_10767);
nor U19965 (N_19965,N_13503,N_12887);
and U19966 (N_19966,N_10161,N_13496);
and U19967 (N_19967,N_13447,N_10263);
nor U19968 (N_19968,N_11935,N_11928);
nand U19969 (N_19969,N_11622,N_11649);
or U19970 (N_19970,N_12150,N_11825);
and U19971 (N_19971,N_10484,N_11363);
nand U19972 (N_19972,N_13399,N_13979);
and U19973 (N_19973,N_13638,N_14201);
nor U19974 (N_19974,N_13787,N_10811);
or U19975 (N_19975,N_11582,N_13133);
or U19976 (N_19976,N_10089,N_14745);
nor U19977 (N_19977,N_14168,N_10862);
and U19978 (N_19978,N_10249,N_10910);
and U19979 (N_19979,N_13069,N_13278);
nand U19980 (N_19980,N_12785,N_14012);
xor U19981 (N_19981,N_11414,N_11648);
nand U19982 (N_19982,N_13862,N_14141);
nand U19983 (N_19983,N_14237,N_13841);
or U19984 (N_19984,N_12664,N_10246);
and U19985 (N_19985,N_12515,N_14263);
or U19986 (N_19986,N_13844,N_13516);
and U19987 (N_19987,N_14385,N_12063);
nand U19988 (N_19988,N_13755,N_14502);
nor U19989 (N_19989,N_14913,N_11271);
nand U19990 (N_19990,N_14158,N_10830);
xor U19991 (N_19991,N_14329,N_11215);
xnor U19992 (N_19992,N_10178,N_12703);
nor U19993 (N_19993,N_12115,N_12655);
xnor U19994 (N_19994,N_13666,N_11728);
nand U19995 (N_19995,N_10025,N_14548);
nor U19996 (N_19996,N_12407,N_13282);
or U19997 (N_19997,N_11760,N_11012);
nand U19998 (N_19998,N_11921,N_10574);
or U19999 (N_19999,N_12367,N_13909);
nor U20000 (N_20000,N_16721,N_16060);
nor U20001 (N_20001,N_15003,N_15781);
nand U20002 (N_20002,N_17529,N_17517);
nand U20003 (N_20003,N_16324,N_15844);
or U20004 (N_20004,N_15870,N_19966);
nor U20005 (N_20005,N_16710,N_18611);
nand U20006 (N_20006,N_19247,N_15409);
nor U20007 (N_20007,N_16343,N_18831);
nor U20008 (N_20008,N_17575,N_19904);
or U20009 (N_20009,N_19537,N_17512);
nand U20010 (N_20010,N_17294,N_19182);
and U20011 (N_20011,N_15453,N_18185);
nor U20012 (N_20012,N_18087,N_16177);
and U20013 (N_20013,N_17227,N_16755);
or U20014 (N_20014,N_17859,N_19984);
nor U20015 (N_20015,N_19750,N_15364);
or U20016 (N_20016,N_15464,N_17785);
nand U20017 (N_20017,N_17135,N_19001);
nor U20018 (N_20018,N_19049,N_17425);
or U20019 (N_20019,N_16229,N_18782);
and U20020 (N_20020,N_15360,N_17649);
nor U20021 (N_20021,N_18534,N_17933);
nand U20022 (N_20022,N_19032,N_15495);
and U20023 (N_20023,N_17774,N_16331);
nand U20024 (N_20024,N_15880,N_19878);
or U20025 (N_20025,N_18771,N_18430);
or U20026 (N_20026,N_19948,N_16114);
and U20027 (N_20027,N_18973,N_16724);
nand U20028 (N_20028,N_15092,N_19592);
nor U20029 (N_20029,N_17751,N_16938);
nor U20030 (N_20030,N_17349,N_16901);
or U20031 (N_20031,N_17805,N_16923);
and U20032 (N_20032,N_16147,N_18914);
and U20033 (N_20033,N_19362,N_18815);
and U20034 (N_20034,N_19832,N_19691);
or U20035 (N_20035,N_18727,N_18979);
nor U20036 (N_20036,N_18106,N_19371);
nand U20037 (N_20037,N_19411,N_17794);
xnor U20038 (N_20038,N_15770,N_18671);
nor U20039 (N_20039,N_16879,N_18770);
nand U20040 (N_20040,N_19193,N_15219);
nor U20041 (N_20041,N_17252,N_19671);
and U20042 (N_20042,N_19215,N_15919);
nand U20043 (N_20043,N_18830,N_19583);
nor U20044 (N_20044,N_18392,N_16824);
nand U20045 (N_20045,N_17544,N_18472);
and U20046 (N_20046,N_15735,N_16756);
and U20047 (N_20047,N_15191,N_19239);
and U20048 (N_20048,N_15637,N_19559);
nand U20049 (N_20049,N_19316,N_18555);
and U20050 (N_20050,N_18048,N_18860);
or U20051 (N_20051,N_15171,N_15481);
nand U20052 (N_20052,N_18105,N_16789);
nor U20053 (N_20053,N_18221,N_15228);
nor U20054 (N_20054,N_15660,N_15862);
and U20055 (N_20055,N_19956,N_19120);
or U20056 (N_20056,N_15006,N_18981);
nand U20057 (N_20057,N_17118,N_17417);
or U20058 (N_20058,N_16822,N_16663);
nand U20059 (N_20059,N_16792,N_15542);
nand U20060 (N_20060,N_18485,N_18751);
nor U20061 (N_20061,N_16747,N_19159);
nor U20062 (N_20062,N_19970,N_16280);
nor U20063 (N_20063,N_15855,N_18900);
nor U20064 (N_20064,N_17664,N_16816);
xor U20065 (N_20065,N_17813,N_16194);
or U20066 (N_20066,N_18655,N_15716);
or U20067 (N_20067,N_17139,N_19479);
nand U20068 (N_20068,N_15966,N_17941);
nor U20069 (N_20069,N_18712,N_17490);
nand U20070 (N_20070,N_15188,N_16875);
or U20071 (N_20071,N_19125,N_19503);
xor U20072 (N_20072,N_15907,N_15877);
nor U20073 (N_20073,N_15462,N_15945);
nand U20074 (N_20074,N_19825,N_17606);
nor U20075 (N_20075,N_18670,N_17148);
nor U20076 (N_20076,N_16368,N_18019);
nand U20077 (N_20077,N_15471,N_18188);
xor U20078 (N_20078,N_15552,N_19968);
nor U20079 (N_20079,N_15725,N_19488);
nor U20080 (N_20080,N_17388,N_15574);
and U20081 (N_20081,N_15281,N_16381);
nor U20082 (N_20082,N_17103,N_15043);
xor U20083 (N_20083,N_15227,N_19643);
and U20084 (N_20084,N_15445,N_16803);
nand U20085 (N_20085,N_16785,N_18663);
and U20086 (N_20086,N_18078,N_15489);
xnor U20087 (N_20087,N_18255,N_16825);
or U20088 (N_20088,N_17494,N_18891);
nand U20089 (N_20089,N_18437,N_16205);
xor U20090 (N_20090,N_19084,N_15909);
nor U20091 (N_20091,N_18232,N_15347);
nand U20092 (N_20092,N_17170,N_15494);
and U20093 (N_20093,N_17625,N_18031);
nor U20094 (N_20094,N_16476,N_18781);
nand U20095 (N_20095,N_16491,N_18634);
nand U20096 (N_20096,N_18417,N_18546);
and U20097 (N_20097,N_19278,N_15582);
xnor U20098 (N_20098,N_18396,N_19368);
nor U20099 (N_20099,N_18451,N_19208);
nor U20100 (N_20100,N_16408,N_15968);
and U20101 (N_20101,N_16388,N_16187);
nor U20102 (N_20102,N_19821,N_19017);
or U20103 (N_20103,N_15602,N_15804);
and U20104 (N_20104,N_18657,N_18077);
nand U20105 (N_20105,N_17432,N_19581);
and U20106 (N_20106,N_18370,N_18146);
or U20107 (N_20107,N_18998,N_15189);
and U20108 (N_20108,N_18717,N_15833);
or U20109 (N_20109,N_16505,N_15013);
nand U20110 (N_20110,N_16083,N_17579);
xnor U20111 (N_20111,N_16518,N_17448);
and U20112 (N_20112,N_19720,N_16732);
nand U20113 (N_20113,N_19609,N_18277);
or U20114 (N_20114,N_19301,N_17855);
nand U20115 (N_20115,N_18354,N_17078);
nor U20116 (N_20116,N_16726,N_15728);
or U20117 (N_20117,N_15402,N_15841);
and U20118 (N_20118,N_17823,N_19109);
and U20119 (N_20119,N_18173,N_15882);
and U20120 (N_20120,N_16941,N_19858);
or U20121 (N_20121,N_15195,N_15576);
nor U20122 (N_20122,N_16853,N_16902);
and U20123 (N_20123,N_17628,N_15067);
or U20124 (N_20124,N_15640,N_19596);
nand U20125 (N_20125,N_16530,N_18487);
nor U20126 (N_20126,N_15001,N_16492);
or U20127 (N_20127,N_18114,N_17197);
and U20128 (N_20128,N_17931,N_18044);
or U20129 (N_20129,N_17314,N_19519);
nand U20130 (N_20130,N_19378,N_17532);
and U20131 (N_20131,N_17927,N_17757);
or U20132 (N_20132,N_19299,N_15987);
and U20133 (N_20133,N_17706,N_16386);
nor U20134 (N_20134,N_18462,N_16691);
or U20135 (N_20135,N_19327,N_15650);
nor U20136 (N_20136,N_15478,N_19726);
and U20137 (N_20137,N_16156,N_19361);
nor U20138 (N_20138,N_19561,N_19990);
or U20139 (N_20139,N_18647,N_19211);
nor U20140 (N_20140,N_15981,N_15423);
xnor U20141 (N_20141,N_17275,N_17693);
nor U20142 (N_20142,N_16043,N_16731);
nand U20143 (N_20143,N_19422,N_17109);
nor U20144 (N_20144,N_15399,N_18756);
nor U20145 (N_20145,N_19920,N_15962);
nand U20146 (N_20146,N_15821,N_19744);
and U20147 (N_20147,N_15524,N_19704);
nand U20148 (N_20148,N_19692,N_18536);
nor U20149 (N_20149,N_16576,N_17348);
nand U20150 (N_20150,N_18303,N_16104);
nor U20151 (N_20151,N_18151,N_15739);
or U20152 (N_20152,N_15479,N_18873);
nor U20153 (N_20153,N_15359,N_15801);
xnor U20154 (N_20154,N_17089,N_19283);
nand U20155 (N_20155,N_19250,N_17872);
nor U20156 (N_20156,N_19660,N_15289);
nor U20157 (N_20157,N_17120,N_15624);
or U20158 (N_20158,N_17746,N_16071);
or U20159 (N_20159,N_18264,N_18950);
and U20160 (N_20160,N_19797,N_15349);
or U20161 (N_20161,N_15087,N_15599);
or U20162 (N_20162,N_17374,N_15810);
or U20163 (N_20163,N_17600,N_15208);
or U20164 (N_20164,N_19908,N_15580);
xnor U20165 (N_20165,N_19253,N_16804);
nor U20166 (N_20166,N_17861,N_15727);
nor U20167 (N_20167,N_15717,N_19937);
nor U20168 (N_20168,N_18202,N_16794);
and U20169 (N_20169,N_17779,N_18788);
xnor U20170 (N_20170,N_16089,N_16238);
nor U20171 (N_20171,N_18501,N_18636);
nor U20172 (N_20172,N_16348,N_19779);
nand U20173 (N_20173,N_15572,N_15374);
nor U20174 (N_20174,N_17962,N_17955);
nand U20175 (N_20175,N_17057,N_16657);
nand U20176 (N_20176,N_16428,N_19381);
nand U20177 (N_20177,N_18988,N_19505);
nand U20178 (N_20178,N_18267,N_15772);
and U20179 (N_20179,N_17787,N_17145);
or U20180 (N_20180,N_17949,N_15839);
or U20181 (N_20181,N_17789,N_17034);
nand U20182 (N_20182,N_15285,N_17590);
or U20183 (N_20183,N_18650,N_18116);
or U20184 (N_20184,N_18424,N_19334);
or U20185 (N_20185,N_17504,N_19881);
nor U20186 (N_20186,N_17844,N_16859);
or U20187 (N_20187,N_16488,N_18579);
nor U20188 (N_20188,N_15142,N_19897);
xnor U20189 (N_20189,N_15361,N_15345);
xor U20190 (N_20190,N_17800,N_17188);
nand U20191 (N_20191,N_16351,N_19077);
or U20192 (N_20192,N_17418,N_15775);
or U20193 (N_20193,N_18644,N_16671);
and U20194 (N_20194,N_15262,N_15103);
xor U20195 (N_20195,N_18660,N_19845);
and U20196 (N_20196,N_18390,N_15504);
and U20197 (N_20197,N_15747,N_18183);
or U20198 (N_20198,N_18737,N_17480);
nor U20199 (N_20199,N_16556,N_19550);
xnor U20200 (N_20200,N_16734,N_18174);
nand U20201 (N_20201,N_19339,N_17905);
nand U20202 (N_20202,N_19453,N_17077);
and U20203 (N_20203,N_15267,N_16416);
and U20204 (N_20204,N_15999,N_16067);
or U20205 (N_20205,N_17142,N_17611);
nand U20206 (N_20206,N_17442,N_15398);
or U20207 (N_20207,N_17690,N_18394);
or U20208 (N_20208,N_18736,N_19628);
nand U20209 (N_20209,N_18672,N_18235);
nor U20210 (N_20210,N_18231,N_19147);
or U20211 (N_20211,N_18250,N_17887);
and U20212 (N_20212,N_17341,N_16797);
nand U20213 (N_20213,N_15199,N_17129);
nand U20214 (N_20214,N_15928,N_16338);
nand U20215 (N_20215,N_16310,N_18310);
or U20216 (N_20216,N_19263,N_18856);
nor U20217 (N_20217,N_16024,N_15930);
or U20218 (N_20218,N_17873,N_16312);
nor U20219 (N_20219,N_19444,N_18641);
and U20220 (N_20220,N_15150,N_17092);
or U20221 (N_20221,N_16033,N_18777);
or U20222 (N_20222,N_16969,N_17685);
nor U20223 (N_20223,N_17826,N_17242);
and U20224 (N_20224,N_16066,N_15136);
or U20225 (N_20225,N_17194,N_18679);
or U20226 (N_20226,N_17229,N_17498);
nand U20227 (N_20227,N_17760,N_15785);
xnor U20228 (N_20228,N_19407,N_18999);
or U20229 (N_20229,N_17722,N_16955);
nand U20230 (N_20230,N_16943,N_16693);
nand U20231 (N_20231,N_16313,N_17731);
nor U20232 (N_20232,N_18735,N_18119);
xor U20233 (N_20233,N_16904,N_19814);
nor U20234 (N_20234,N_18564,N_18141);
xnor U20235 (N_20235,N_19457,N_15522);
nand U20236 (N_20236,N_16744,N_17668);
and U20237 (N_20237,N_19261,N_16526);
and U20238 (N_20238,N_19273,N_17978);
xor U20239 (N_20239,N_17713,N_15330);
and U20240 (N_20240,N_16222,N_15221);
and U20241 (N_20241,N_16615,N_19560);
or U20242 (N_20242,N_15961,N_18924);
nand U20243 (N_20243,N_18402,N_15498);
nor U20244 (N_20244,N_16757,N_19372);
xnor U20245 (N_20245,N_17430,N_19186);
nor U20246 (N_20246,N_16144,N_18347);
nor U20247 (N_20247,N_15560,N_17121);
and U20248 (N_20248,N_19585,N_15419);
nand U20249 (N_20249,N_18653,N_19356);
nand U20250 (N_20250,N_16165,N_16515);
nor U20251 (N_20251,N_18866,N_16942);
or U20252 (N_20252,N_18126,N_16405);
nand U20253 (N_20253,N_16149,N_17535);
and U20254 (N_20254,N_15625,N_16051);
or U20255 (N_20255,N_15031,N_16211);
or U20256 (N_20256,N_16344,N_16117);
nor U20257 (N_20257,N_19673,N_16133);
and U20258 (N_20258,N_17870,N_17750);
nor U20259 (N_20259,N_15411,N_18335);
or U20260 (N_20260,N_19196,N_16329);
or U20261 (N_20261,N_18586,N_17093);
or U20262 (N_20262,N_19375,N_15109);
xor U20263 (N_20263,N_19954,N_18947);
and U20264 (N_20264,N_16784,N_16746);
nor U20265 (N_20265,N_17330,N_19936);
nor U20266 (N_20266,N_15593,N_16267);
and U20267 (N_20267,N_17683,N_18263);
nor U20268 (N_20268,N_17908,N_17133);
or U20269 (N_20269,N_17288,N_16143);
nor U20270 (N_20270,N_19003,N_16684);
and U20271 (N_20271,N_19044,N_18740);
nand U20272 (N_20272,N_19083,N_15940);
and U20273 (N_20273,N_19896,N_19168);
or U20274 (N_20274,N_17391,N_17096);
or U20275 (N_20275,N_18957,N_19341);
and U20276 (N_20276,N_15678,N_15714);
nand U20277 (N_20277,N_18904,N_18554);
and U20278 (N_20278,N_18509,N_16443);
nor U20279 (N_20279,N_17106,N_19798);
nand U20280 (N_20280,N_17111,N_16524);
nor U20281 (N_20281,N_17607,N_18387);
nand U20282 (N_20282,N_18172,N_17963);
nand U20283 (N_20283,N_17627,N_19235);
xor U20284 (N_20284,N_16619,N_18715);
or U20285 (N_20285,N_18014,N_19194);
and U20286 (N_20286,N_19487,N_18137);
nor U20287 (N_20287,N_15960,N_17682);
or U20288 (N_20288,N_16375,N_16290);
or U20289 (N_20289,N_15338,N_15311);
nor U20290 (N_20290,N_19342,N_16704);
xnor U20291 (N_20291,N_16586,N_17201);
xor U20292 (N_20292,N_17723,N_15258);
and U20293 (N_20293,N_19843,N_17198);
and U20294 (N_20294,N_17609,N_18313);
and U20295 (N_20295,N_19650,N_16537);
nand U20296 (N_20296,N_19626,N_19376);
or U20297 (N_20297,N_19013,N_17204);
nor U20298 (N_20298,N_17755,N_15197);
nand U20299 (N_20299,N_17210,N_19112);
nand U20300 (N_20300,N_19094,N_17810);
or U20301 (N_20301,N_17839,N_18719);
or U20302 (N_20302,N_16855,N_16627);
nand U20303 (N_20303,N_18571,N_15000);
and U20304 (N_20304,N_18694,N_17646);
nor U20305 (N_20305,N_15416,N_17333);
xnor U20306 (N_20306,N_16864,N_15662);
nand U20307 (N_20307,N_19326,N_15731);
and U20308 (N_20308,N_15809,N_17350);
or U20309 (N_20309,N_16644,N_16272);
nor U20310 (N_20310,N_18187,N_15892);
nor U20311 (N_20311,N_16982,N_19141);
nor U20312 (N_20312,N_15314,N_15965);
nor U20313 (N_20313,N_18055,N_18937);
nand U20314 (N_20314,N_18320,N_18018);
xnor U20315 (N_20315,N_17320,N_19288);
or U20316 (N_20316,N_15248,N_16101);
or U20317 (N_20317,N_15115,N_16018);
and U20318 (N_20318,N_15759,N_19806);
nor U20319 (N_20319,N_16300,N_19218);
nor U20320 (N_20320,N_18400,N_19739);
nand U20321 (N_20321,N_16134,N_18799);
xor U20322 (N_20322,N_19202,N_17977);
and U20323 (N_20323,N_16577,N_18618);
or U20324 (N_20324,N_17302,N_15851);
and U20325 (N_20325,N_18812,N_17586);
and U20326 (N_20326,N_19160,N_15861);
and U20327 (N_20327,N_16553,N_16285);
or U20328 (N_20328,N_19982,N_16517);
nor U20329 (N_20329,N_16400,N_19213);
and U20330 (N_20330,N_17122,N_19575);
and U20331 (N_20331,N_15754,N_16335);
or U20332 (N_20332,N_16620,N_16600);
nor U20333 (N_20333,N_15647,N_19976);
nor U20334 (N_20334,N_19593,N_15694);
and U20335 (N_20335,N_18810,N_15561);
and U20336 (N_20336,N_15200,N_19514);
nand U20337 (N_20337,N_16202,N_17205);
and U20338 (N_20338,N_16899,N_15057);
nor U20339 (N_20339,N_16493,N_16738);
nand U20340 (N_20340,N_18862,N_19469);
and U20341 (N_20341,N_18104,N_19981);
xor U20342 (N_20342,N_19354,N_15487);
nor U20343 (N_20343,N_16812,N_15070);
and U20344 (N_20344,N_18590,N_16836);
nor U20345 (N_20345,N_15286,N_18177);
or U20346 (N_20346,N_18423,N_15021);
or U20347 (N_20347,N_15900,N_18120);
and U20348 (N_20348,N_16543,N_15540);
and U20349 (N_20349,N_19577,N_18569);
nor U20350 (N_20350,N_16447,N_15808);
or U20351 (N_20351,N_18338,N_15519);
nor U20352 (N_20352,N_19258,N_19403);
nor U20353 (N_20353,N_19297,N_17837);
and U20354 (N_20354,N_17782,N_17191);
nor U20355 (N_20355,N_17564,N_16781);
xor U20356 (N_20356,N_18787,N_19226);
and U20357 (N_20357,N_17441,N_16076);
nor U20358 (N_20358,N_19494,N_18466);
and U20359 (N_20359,N_17484,N_18742);
nor U20360 (N_20360,N_15920,N_15817);
or U20361 (N_20361,N_17824,N_15350);
and U20362 (N_20362,N_18206,N_18438);
or U20363 (N_20363,N_16643,N_17486);
nor U20364 (N_20364,N_15768,N_19031);
nor U20365 (N_20365,N_18377,N_17551);
nand U20366 (N_20366,N_16799,N_19364);
or U20367 (N_20367,N_18455,N_19818);
nor U20368 (N_20368,N_15659,N_15098);
and U20369 (N_20369,N_15045,N_17657);
and U20370 (N_20370,N_18794,N_18955);
nor U20371 (N_20371,N_16362,N_18245);
nand U20372 (N_20372,N_18932,N_16891);
xnor U20373 (N_20373,N_16289,N_15414);
xnor U20374 (N_20374,N_17331,N_17738);
xor U20375 (N_20375,N_15904,N_16056);
and U20376 (N_20376,N_16714,N_18364);
and U20377 (N_20377,N_17289,N_19060);
and U20378 (N_20378,N_18021,N_19839);
or U20379 (N_20379,N_18213,N_15667);
or U20380 (N_20380,N_15060,N_19498);
and U20381 (N_20381,N_15251,N_18272);
xor U20382 (N_20382,N_18702,N_17406);
and U20383 (N_20383,N_18916,N_15569);
nand U20384 (N_20384,N_15065,N_17412);
nor U20385 (N_20385,N_17240,N_19582);
or U20386 (N_20386,N_16481,N_17354);
nand U20387 (N_20387,N_15636,N_18337);
nand U20388 (N_20388,N_15905,N_15866);
or U20389 (N_20389,N_18163,N_19370);
and U20390 (N_20390,N_15134,N_16345);
nor U20391 (N_20391,N_15293,N_15229);
or U20392 (N_20392,N_19713,N_16429);
nor U20393 (N_20393,N_19723,N_17334);
nor U20394 (N_20394,N_16639,N_19344);
nand U20395 (N_20395,N_17665,N_16469);
and U20396 (N_20396,N_19760,N_18314);
or U20397 (N_20397,N_16501,N_19535);
or U20398 (N_20398,N_17613,N_19078);
and U20399 (N_20399,N_16768,N_15310);
or U20400 (N_20400,N_17137,N_17904);
or U20401 (N_20401,N_16183,N_16733);
xnor U20402 (N_20402,N_17439,N_16094);
and U20403 (N_20403,N_15052,N_15983);
nor U20404 (N_20404,N_19601,N_15538);
and U20405 (N_20405,N_17042,N_15100);
and U20406 (N_20406,N_15680,N_15779);
and U20407 (N_20407,N_18557,N_18158);
or U20408 (N_20408,N_19868,N_17891);
and U20409 (N_20409,N_15784,N_17394);
nor U20410 (N_20410,N_16573,N_16878);
or U20411 (N_20411,N_16241,N_16540);
xnor U20412 (N_20412,N_17729,N_16893);
or U20413 (N_20413,N_15135,N_15544);
or U20414 (N_20414,N_15510,N_15496);
nand U20415 (N_20415,N_18881,N_16778);
and U20416 (N_20416,N_18203,N_15891);
or U20417 (N_20417,N_18409,N_18161);
or U20418 (N_20418,N_19985,N_17603);
nand U20419 (N_20419,N_15170,N_18459);
nand U20420 (N_20420,N_16158,N_15884);
or U20421 (N_20421,N_19799,N_16762);
nand U20422 (N_20422,N_17297,N_16178);
or U20423 (N_20423,N_17743,N_19068);
nor U20424 (N_20424,N_17992,N_19969);
and U20425 (N_20425,N_16887,N_18017);
nand U20426 (N_20426,N_17836,N_16589);
and U20427 (N_20427,N_18397,N_17518);
nor U20428 (N_20428,N_18926,N_19886);
or U20429 (N_20429,N_16145,N_16995);
xor U20430 (N_20430,N_17368,N_19611);
nand U20431 (N_20431,N_18069,N_15047);
nand U20432 (N_20432,N_16279,N_19617);
xor U20433 (N_20433,N_19678,N_16295);
nor U20434 (N_20434,N_18257,N_18271);
nand U20435 (N_20435,N_18329,N_18179);
or U20436 (N_20436,N_16990,N_18222);
xor U20437 (N_20437,N_19999,N_16499);
or U20438 (N_20438,N_16616,N_17361);
or U20439 (N_20439,N_19658,N_16379);
and U20440 (N_20440,N_19621,N_19396);
and U20441 (N_20441,N_16602,N_17593);
xnor U20442 (N_20442,N_19192,N_15936);
nor U20443 (N_20443,N_18075,N_17392);
and U20444 (N_20444,N_16707,N_16139);
and U20445 (N_20445,N_16508,N_16209);
and U20446 (N_20446,N_16422,N_19055);
and U20447 (N_20447,N_18109,N_16450);
or U20448 (N_20448,N_18906,N_16008);
or U20449 (N_20449,N_16782,N_19104);
or U20450 (N_20450,N_18654,N_18561);
or U20451 (N_20451,N_18797,N_15700);
xor U20452 (N_20452,N_17793,N_17671);
or U20453 (N_20453,N_17076,N_18913);
and U20454 (N_20454,N_17231,N_16017);
or U20455 (N_20455,N_18925,N_15849);
or U20456 (N_20456,N_17910,N_18285);
or U20457 (N_20457,N_19777,N_18391);
and U20458 (N_20458,N_17470,N_15268);
and U20459 (N_20459,N_19360,N_18268);
or U20460 (N_20460,N_15566,N_16698);
and U20461 (N_20461,N_18821,N_15749);
nand U20462 (N_20462,N_16949,N_19511);
nand U20463 (N_20463,N_17270,N_17832);
and U20464 (N_20464,N_15107,N_15664);
or U20465 (N_20465,N_19891,N_18418);
and U20466 (N_20466,N_15748,N_16580);
and U20467 (N_20467,N_16059,N_17301);
nor U20468 (N_20468,N_16411,N_19207);
nand U20469 (N_20469,N_18677,N_18484);
nand U20470 (N_20470,N_16695,N_19011);
nor U20471 (N_20471,N_19994,N_19964);
and U20472 (N_20472,N_16365,N_16182);
nor U20473 (N_20473,N_17276,N_18816);
or U20474 (N_20474,N_17986,N_16217);
and U20475 (N_20475,N_16304,N_16314);
nand U20476 (N_20476,N_15383,N_15832);
xor U20477 (N_20477,N_16281,N_15746);
or U20478 (N_20478,N_15492,N_18820);
nor U20479 (N_20479,N_18622,N_19106);
or U20480 (N_20480,N_17929,N_15812);
nor U20481 (N_20481,N_16937,N_19103);
and U20482 (N_20482,N_16532,N_17259);
xor U20483 (N_20483,N_17852,N_15715);
and U20484 (N_20484,N_19063,N_18166);
or U20485 (N_20485,N_18674,N_17655);
and U20486 (N_20486,N_18503,N_16519);
nand U20487 (N_20487,N_18627,N_18288);
and U20488 (N_20488,N_18351,N_19766);
nand U20489 (N_20489,N_17150,N_16819);
and U20490 (N_20490,N_16363,N_16545);
xnor U20491 (N_20491,N_19652,N_18454);
and U20492 (N_20492,N_18295,N_17193);
and U20493 (N_20493,N_18333,N_16699);
nor U20494 (N_20494,N_18444,N_16503);
xor U20495 (N_20495,N_15823,N_18518);
nor U20496 (N_20496,N_19882,N_15058);
and U20497 (N_20497,N_17695,N_16559);
nor U20498 (N_20498,N_19566,N_15484);
nor U20499 (N_20499,N_16884,N_17475);
and U20500 (N_20500,N_17857,N_18275);
nand U20501 (N_20501,N_17011,N_18698);
nor U20502 (N_20502,N_16903,N_15249);
nand U20503 (N_20503,N_16767,N_18208);
xor U20504 (N_20504,N_19402,N_15245);
or U20505 (N_20505,N_17635,N_18649);
nor U20506 (N_20506,N_15250,N_17526);
or U20507 (N_20507,N_17730,N_19705);
xor U20508 (N_20508,N_18992,N_19808);
nor U20509 (N_20509,N_15253,N_18869);
and U20510 (N_20510,N_18646,N_19312);
and U20511 (N_20511,N_15408,N_16035);
or U20512 (N_20512,N_15154,N_17572);
and U20513 (N_20513,N_17450,N_15686);
nor U20514 (N_20514,N_17890,N_17206);
xor U20515 (N_20515,N_19648,N_17726);
nor U20516 (N_20516,N_18365,N_19082);
or U20517 (N_20517,N_18958,N_15061);
or U20518 (N_20518,N_16701,N_19786);
nor U20519 (N_20519,N_18130,N_18690);
and U20520 (N_20520,N_16246,N_18847);
nor U20521 (N_20521,N_17402,N_19038);
xnor U20522 (N_20522,N_17939,N_19824);
and U20523 (N_20523,N_16783,N_17059);
nor U20524 (N_20524,N_15993,N_16849);
nand U20525 (N_20525,N_17262,N_19507);
or U20526 (N_20526,N_18884,N_15139);
and U20527 (N_20527,N_19431,N_15302);
nand U20528 (N_20528,N_15385,N_15159);
and U20529 (N_20529,N_17217,N_15737);
xor U20530 (N_20530,N_17553,N_18152);
and U20531 (N_20531,N_19623,N_17942);
nand U20532 (N_20532,N_16082,N_19244);
xnor U20533 (N_20533,N_16420,N_17436);
nand U20534 (N_20534,N_16474,N_17124);
or U20535 (N_20535,N_19091,N_16833);
xnor U20536 (N_20536,N_17419,N_15137);
nand U20537 (N_20537,N_18028,N_18039);
nand U20538 (N_20538,N_18239,N_19745);
nand U20539 (N_20539,N_19931,N_16265);
and U20540 (N_20540,N_19093,N_19852);
nor U20541 (N_20541,N_16821,N_19119);
and U20542 (N_20542,N_15722,N_15676);
nand U20543 (N_20543,N_19409,N_19815);
and U20544 (N_20544,N_18410,N_19796);
and U20545 (N_20545,N_18378,N_18469);
and U20546 (N_20546,N_15956,N_16844);
nor U20547 (N_20547,N_18291,N_18342);
nand U20548 (N_20548,N_16963,N_16337);
nand U20549 (N_20549,N_17786,N_15670);
nor U20550 (N_20550,N_17640,N_17525);
or U20551 (N_20551,N_18298,N_15015);
nor U20552 (N_20552,N_16448,N_18997);
or U20553 (N_20553,N_15284,N_19893);
nor U20554 (N_20554,N_17183,N_16658);
nand U20555 (N_20555,N_18020,N_19699);
or U20556 (N_20556,N_18135,N_15648);
nor U20557 (N_20557,N_15701,N_15413);
nand U20558 (N_20558,N_15366,N_16584);
nand U20559 (N_20559,N_15192,N_16213);
nor U20560 (N_20560,N_15308,N_19790);
xor U20561 (N_20561,N_19903,N_16551);
xnor U20562 (N_20562,N_17085,N_19480);
xor U20563 (N_20563,N_15220,N_16826);
nor U20564 (N_20564,N_17167,N_15842);
nor U20565 (N_20565,N_15549,N_19269);
and U20566 (N_20566,N_19458,N_17648);
and U20567 (N_20567,N_19940,N_18350);
nor U20568 (N_20568,N_19087,N_19268);
nor U20569 (N_20569,N_18718,N_17620);
nand U20570 (N_20570,N_19419,N_17728);
nor U20571 (N_20571,N_15089,N_18837);
nor U20572 (N_20572,N_19670,N_17060);
or U20573 (N_20573,N_19081,N_18949);
or U20574 (N_20574,N_16967,N_19146);
nand U20575 (N_20575,N_17783,N_18850);
nor U20576 (N_20576,N_16110,N_16687);
or U20577 (N_20577,N_18316,N_18961);
nor U20578 (N_20578,N_17666,N_19317);
or U20579 (N_20579,N_16052,N_17951);
or U20580 (N_20580,N_19659,N_15982);
and U20581 (N_20581,N_16357,N_16451);
or U20582 (N_20582,N_17151,N_19313);
nor U20583 (N_20583,N_17408,N_19006);
xor U20584 (N_20584,N_17416,N_19241);
nand U20585 (N_20585,N_19460,N_17458);
nand U20586 (N_20586,N_17375,N_18952);
nor U20587 (N_20587,N_15834,N_16549);
nand U20588 (N_20588,N_18595,N_19154);
nand U20589 (N_20589,N_16404,N_16055);
nor U20590 (N_20590,N_18261,N_16888);
nor U20591 (N_20591,N_19130,N_15603);
xor U20592 (N_20592,N_18624,N_17980);
or U20593 (N_20593,N_15019,N_19600);
or U20594 (N_20594,N_17952,N_17692);
nor U20595 (N_20595,N_19649,N_19425);
xor U20596 (N_20596,N_16471,N_19547);
or U20597 (N_20597,N_17537,N_18969);
and U20598 (N_20598,N_15455,N_19837);
nand U20599 (N_20599,N_15183,N_15953);
or U20600 (N_20600,N_16924,N_17843);
nor U20601 (N_20601,N_18845,N_19849);
or U20602 (N_20602,N_17175,N_19180);
or U20603 (N_20603,N_18253,N_17703);
nor U20604 (N_20604,N_18097,N_18523);
and U20605 (N_20605,N_15923,N_19545);
and U20606 (N_20606,N_15971,N_15023);
or U20607 (N_20607,N_17007,N_18854);
and U20608 (N_20608,N_15029,N_15612);
nand U20609 (N_20609,N_18994,N_16392);
and U20610 (N_20610,N_17009,N_16210);
xnor U20611 (N_20611,N_15073,N_15016);
xnor U20612 (N_20612,N_19683,N_15326);
nor U20613 (N_20613,N_19171,N_15879);
and U20614 (N_20614,N_19729,N_17223);
nor U20615 (N_20615,N_18504,N_16058);
nor U20616 (N_20616,N_19176,N_17047);
nor U20617 (N_20617,N_16261,N_19775);
or U20618 (N_20618,N_15578,N_17497);
nand U20619 (N_20619,N_16396,N_19747);
nand U20620 (N_20620,N_17756,N_15329);
and U20621 (N_20621,N_16814,N_19754);
and U20622 (N_20622,N_19382,N_18975);
and U20623 (N_20623,N_15468,N_15427);
nor U20624 (N_20624,N_18131,N_18897);
nand U20625 (N_20625,N_17686,N_15819);
nand U20626 (N_20626,N_16203,N_16557);
nand U20627 (N_20627,N_16457,N_18773);
nand U20628 (N_20628,N_17926,N_17975);
nand U20629 (N_20629,N_16542,N_18825);
xnor U20630 (N_20630,N_16236,N_18578);
or U20631 (N_20631,N_17364,N_18544);
nor U20632 (N_20632,N_19579,N_17894);
or U20633 (N_20633,N_16061,N_18107);
nand U20634 (N_20634,N_15184,N_19455);
or U20635 (N_20635,N_15247,N_18665);
nand U20636 (N_20636,N_18764,N_18058);
nor U20637 (N_20637,N_19025,N_16248);
and U20638 (N_20638,N_18893,N_17702);
nand U20639 (N_20639,N_15541,N_15179);
and U20640 (N_20640,N_19987,N_17560);
nor U20641 (N_20641,N_18332,N_17892);
or U20642 (N_20642,N_18465,N_15025);
nor U20643 (N_20643,N_19653,N_18761);
or U20644 (N_20644,N_16989,N_16087);
nand U20645 (N_20645,N_16424,N_15318);
or U20646 (N_20646,N_19132,N_18868);
xor U20647 (N_20647,N_19465,N_16005);
or U20648 (N_20648,N_16948,N_16108);
nor U20649 (N_20649,N_19447,N_16015);
and U20650 (N_20650,N_19838,N_17169);
and U20651 (N_20651,N_18818,N_19497);
nand U20652 (N_20652,N_17667,N_16098);
or U20653 (N_20653,N_18970,N_19847);
nand U20654 (N_20654,N_17046,N_18246);
xor U20655 (N_20655,N_19558,N_15325);
xnor U20656 (N_20656,N_18201,N_17511);
and U20657 (N_20657,N_17357,N_18522);
or U20658 (N_20658,N_15619,N_15932);
and U20659 (N_20659,N_18008,N_17616);
nand U20660 (N_20660,N_15649,N_16831);
nand U20661 (N_20661,N_19138,N_19406);
and U20662 (N_20662,N_15681,N_16996);
nor U20663 (N_20663,N_16111,N_18005);
or U20664 (N_20664,N_19466,N_16328);
nor U20665 (N_20665,N_19870,N_16851);
and U20666 (N_20666,N_15404,N_16900);
or U20667 (N_20667,N_15762,N_16307);
or U20668 (N_20668,N_18311,N_18813);
nand U20669 (N_20669,N_19439,N_16249);
nor U20670 (N_20670,N_18938,N_16601);
nand U20671 (N_20671,N_19432,N_16195);
and U20672 (N_20672,N_19385,N_17026);
and U20673 (N_20673,N_16006,N_19927);
and U20674 (N_20674,N_15825,N_19756);
or U20675 (N_20675,N_18903,N_19115);
or U20676 (N_20676,N_19199,N_19369);
nor U20677 (N_20677,N_16839,N_19733);
and U20678 (N_20678,N_16538,N_15127);
xnor U20679 (N_20679,N_16637,N_15244);
and U20680 (N_20680,N_16766,N_18468);
and U20681 (N_20681,N_17777,N_19532);
and U20682 (N_20682,N_15690,N_19963);
and U20683 (N_20683,N_17050,N_19635);
nand U20684 (N_20684,N_18507,N_17717);
nor U20685 (N_20685,N_16237,N_19928);
nand U20686 (N_20686,N_17817,N_19397);
nand U20687 (N_20687,N_16976,N_19462);
and U20688 (N_20688,N_18062,N_17192);
or U20689 (N_20689,N_17144,N_16497);
nand U20690 (N_20690,N_19228,N_16876);
xnor U20691 (N_20691,N_19538,N_18905);
nand U20692 (N_20692,N_16200,N_15653);
xnor U20693 (N_20693,N_16527,N_16048);
nand U20694 (N_20694,N_18894,N_19076);
and U20695 (N_20695,N_15274,N_18936);
nand U20696 (N_20696,N_19647,N_18695);
nand U20697 (N_20697,N_17835,N_19061);
nor U20698 (N_20698,N_18247,N_17338);
or U20699 (N_20699,N_18760,N_15548);
or U20700 (N_20700,N_17679,N_19096);
and U20701 (N_20701,N_19805,N_16273);
and U20702 (N_20702,N_16494,N_15559);
and U20703 (N_20703,N_18553,N_19501);
nor U20704 (N_20704,N_19026,N_15486);
nor U20705 (N_20705,N_19787,N_16962);
nor U20706 (N_20706,N_17538,N_16862);
nand U20707 (N_20707,N_16278,N_15467);
or U20708 (N_20708,N_16309,N_17546);
nand U20709 (N_20709,N_16513,N_17174);
and U20710 (N_20710,N_15642,N_18643);
xor U20711 (N_20711,N_18326,N_17523);
or U20712 (N_20712,N_17776,N_19276);
xor U20713 (N_20713,N_16449,N_19090);
nand U20714 (N_20714,N_19393,N_18068);
or U20715 (N_20715,N_18429,N_19349);
or U20716 (N_20716,N_15926,N_16649);
or U20717 (N_20717,N_19978,N_16169);
or U20718 (N_20718,N_19230,N_16652);
and U20719 (N_20719,N_19126,N_19571);
nand U20720 (N_20720,N_18061,N_15234);
nor U20721 (N_20721,N_19291,N_15611);
and U20722 (N_20722,N_18081,N_17922);
nor U20723 (N_20723,N_18072,N_18604);
nand U20724 (N_20724,N_19884,N_17195);
nand U20725 (N_20725,N_16742,N_15646);
and U20726 (N_20726,N_16847,N_18279);
and U20727 (N_20727,N_19315,N_18610);
nor U20728 (N_20728,N_19694,N_18360);
and U20729 (N_20729,N_17973,N_16977);
and U20730 (N_20730,N_15130,N_19175);
or U20731 (N_20731,N_16146,N_17687);
or U20732 (N_20732,N_15658,N_19546);
nand U20733 (N_20733,N_16907,N_15209);
or U20734 (N_20734,N_18315,N_16407);
and U20735 (N_20735,N_15094,N_18098);
or U20736 (N_20736,N_18852,N_15177);
xor U20737 (N_20737,N_19274,N_19792);
and U20738 (N_20738,N_17112,N_18965);
and U20739 (N_20739,N_15201,N_19092);
nand U20740 (N_20740,N_17116,N_15679);
nand U20741 (N_20741,N_15056,N_18563);
nor U20742 (N_20742,N_15654,N_19944);
or U20743 (N_20743,N_15205,N_19167);
nor U20744 (N_20744,N_15692,N_16679);
xnor U20745 (N_20745,N_15534,N_15925);
nor U20746 (N_20746,N_17225,N_17090);
nor U20747 (N_20747,N_18216,N_17984);
nand U20748 (N_20748,N_17156,N_17811);
and U20749 (N_20749,N_17024,N_16199);
or U20750 (N_20750,N_19300,N_17647);
nand U20751 (N_20751,N_19980,N_15908);
and U20752 (N_20752,N_18739,N_16818);
nand U20753 (N_20753,N_18870,N_15336);
nand U20754 (N_20754,N_18776,N_17916);
xor U20755 (N_20755,N_15613,N_17365);
nand U20756 (N_20756,N_19311,N_16670);
nand U20757 (N_20757,N_18506,N_16669);
nand U20758 (N_20758,N_15256,N_17732);
nor U20759 (N_20759,N_17882,N_15764);
nor U20760 (N_20760,N_17267,N_18796);
nand U20761 (N_20761,N_17736,N_17960);
or U20762 (N_20762,N_19735,N_17999);
nand U20763 (N_20763,N_18480,N_16242);
and U20764 (N_20764,N_17040,N_16102);
and U20765 (N_20765,N_17389,N_18099);
nand U20766 (N_20766,N_16034,N_16093);
and U20767 (N_20767,N_17382,N_19005);
xor U20768 (N_20768,N_16536,N_17554);
and U20769 (N_20769,N_16998,N_17282);
or U20770 (N_20770,N_18328,N_17213);
and U20771 (N_20771,N_17502,N_16456);
and U20772 (N_20772,N_19024,N_16592);
or U20773 (N_20773,N_16383,N_16713);
xor U20774 (N_20774,N_18642,N_19785);
nand U20775 (N_20775,N_18419,N_15622);
nor U20776 (N_20776,N_15763,N_16788);
xor U20777 (N_20777,N_18252,N_18804);
nor U20778 (N_20778,N_15948,N_16394);
nand U20779 (N_20779,N_15435,N_17164);
nor U20780 (N_20780,N_16629,N_15595);
nor U20781 (N_20781,N_16226,N_16820);
nand U20782 (N_20782,N_19145,N_18381);
nand U20783 (N_20783,N_17337,N_16945);
xor U20784 (N_20784,N_18157,N_18368);
and U20785 (N_20785,N_17626,N_19846);
nand U20786 (N_20786,N_16896,N_15601);
nor U20787 (N_20787,N_16906,N_17281);
xor U20788 (N_20788,N_16410,N_16270);
nand U20789 (N_20789,N_16239,N_19266);
or U20790 (N_20790,N_19391,N_15316);
xnor U20791 (N_20791,N_17715,N_15463);
nor U20792 (N_20792,N_15372,N_15111);
xnor U20793 (N_20793,N_15963,N_17202);
and U20794 (N_20794,N_15931,N_17309);
and U20795 (N_20795,N_19067,N_16320);
and U20796 (N_20796,N_16359,N_19850);
nor U20797 (N_20797,N_17815,N_16414);
nand U20798 (N_20798,N_17700,N_15674);
xor U20799 (N_20799,N_17994,N_17642);
nor U20800 (N_20800,N_19959,N_18223);
nand U20801 (N_20801,N_16939,N_18457);
xor U20802 (N_20802,N_18896,N_15598);
and U20803 (N_20803,N_17101,N_17264);
nand U20804 (N_20804,N_18525,N_18408);
or U20805 (N_20805,N_16672,N_15807);
nand U20806 (N_20806,N_17362,N_15906);
nor U20807 (N_20807,N_15859,N_19442);
xnor U20808 (N_20808,N_17663,N_18182);
and U20809 (N_20809,N_16935,N_16252);
nand U20810 (N_20810,N_15472,N_16268);
or U20811 (N_20811,N_15243,N_15126);
nor U20812 (N_20812,N_19638,N_16550);
nand U20813 (N_20813,N_15106,N_15511);
nand U20814 (N_20814,N_19758,N_16037);
or U20815 (N_20815,N_18538,N_16841);
or U20816 (N_20816,N_18389,N_18805);
nand U20817 (N_20817,N_19468,N_19553);
or U20818 (N_20818,N_16728,N_15610);
nand U20819 (N_20819,N_15752,N_16417);
xor U20820 (N_20820,N_15586,N_16306);
or U20821 (N_20821,N_15401,N_17923);
and U20822 (N_20822,N_18625,N_18361);
and U20823 (N_20823,N_16718,N_19184);
nor U20824 (N_20824,N_19252,N_16053);
nand U20825 (N_20825,N_16914,N_18091);
or U20826 (N_20826,N_15755,N_16830);
xor U20827 (N_20827,N_17907,N_16882);
or U20828 (N_20828,N_15490,N_17930);
and U20829 (N_20829,N_15352,N_15048);
nand U20830 (N_20830,N_18617,N_17998);
and U20831 (N_20831,N_16294,N_15026);
xor U20832 (N_20832,N_17015,N_18898);
nand U20833 (N_20833,N_15273,N_19696);
and U20834 (N_20834,N_17481,N_17107);
and U20835 (N_20835,N_17950,N_18224);
xor U20836 (N_20836,N_17804,N_15055);
nor U20837 (N_20837,N_16688,N_17125);
or U20838 (N_20838,N_15114,N_16872);
xnor U20839 (N_20839,N_15776,N_19906);
nor U20840 (N_20840,N_19088,N_19549);
nand U20841 (N_20841,N_18471,N_16617);
or U20842 (N_20842,N_17200,N_15915);
and U20843 (N_20843,N_15133,N_17398);
and U20844 (N_20844,N_16927,N_19198);
nand U20845 (N_20845,N_15080,N_17272);
nand U20846 (N_20846,N_17797,N_19045);
or U20847 (N_20847,N_19856,N_19187);
or U20848 (N_20848,N_17190,N_17018);
or U20849 (N_20849,N_17283,N_18631);
and U20850 (N_20850,N_19279,N_19221);
and U20851 (N_20851,N_19888,N_19737);
nor U20852 (N_20852,N_17074,N_18877);
nand U20853 (N_20853,N_18596,N_16026);
nand U20854 (N_20854,N_15477,N_18322);
and U20855 (N_20855,N_16735,N_19965);
and U20856 (N_20856,N_16574,N_17896);
and U20857 (N_20857,N_19421,N_16770);
nand U20858 (N_20858,N_15148,N_19347);
nor U20859 (N_20859,N_16594,N_19835);
nor U20860 (N_20860,N_18601,N_19495);
nor U20861 (N_20861,N_18100,N_16552);
xnor U20862 (N_20862,N_16869,N_18713);
or U20863 (N_20863,N_16356,N_19725);
and U20864 (N_20864,N_19027,N_19394);
or U20865 (N_20865,N_19086,N_17806);
and U20866 (N_20866,N_19163,N_19599);
nand U20867 (N_20867,N_17387,N_15750);
nor U20868 (N_20868,N_15131,N_15627);
or U20869 (N_20869,N_19639,N_16997);
and U20870 (N_20870,N_19173,N_15878);
or U20871 (N_20871,N_16193,N_17311);
and U20872 (N_20872,N_18366,N_16189);
nand U20873 (N_20873,N_18066,N_18102);
xnor U20874 (N_20874,N_18780,N_19489);
nor U20875 (N_20875,N_18412,N_15163);
or U20876 (N_20876,N_16634,N_16190);
nor U20877 (N_20877,N_19932,N_19050);
nand U20878 (N_20878,N_17029,N_15149);
or U20879 (N_20879,N_15334,N_18659);
or U20880 (N_20880,N_15696,N_15631);
nand U20881 (N_20881,N_19350,N_15447);
xnor U20882 (N_20882,N_18475,N_16922);
or U20883 (N_20883,N_17720,N_19028);
nand U20884 (N_20884,N_18880,N_16608);
nor U20885 (N_20885,N_17016,N_18530);
nand U20886 (N_20886,N_15998,N_18855);
and U20887 (N_20887,N_17110,N_15941);
and U20888 (N_20888,N_15488,N_15687);
and U20889 (N_20889,N_16212,N_16832);
xnor U20890 (N_20890,N_17754,N_17672);
or U20891 (N_20891,N_17796,N_18339);
and U20892 (N_20892,N_15480,N_15354);
nand U20893 (N_20893,N_17744,N_17299);
nor U20894 (N_20894,N_17239,N_18449);
and U20895 (N_20895,N_16012,N_15788);
and U20896 (N_20896,N_19657,N_15942);
nand U20897 (N_20897,N_16244,N_19452);
nor U20898 (N_20898,N_18899,N_16225);
xnor U20899 (N_20899,N_16486,N_19441);
xor U20900 (N_20900,N_16419,N_16905);
and U20901 (N_20901,N_19512,N_17141);
and U20902 (N_20902,N_17917,N_16341);
xnor U20903 (N_20903,N_15363,N_15943);
or U20904 (N_20904,N_15977,N_19724);
or U20905 (N_20905,N_16745,N_19543);
xor U20906 (N_20906,N_15793,N_18628);
nor U20907 (N_20907,N_15324,N_18473);
nor U20908 (N_20908,N_18945,N_17555);
nand U20909 (N_20909,N_19864,N_17065);
and U20910 (N_20910,N_16881,N_18282);
and U20911 (N_20911,N_19046,N_15012);
nand U20912 (N_20912,N_16224,N_17265);
and U20913 (N_20913,N_16890,N_18828);
nand U20914 (N_20914,N_15805,N_18321);
nand U20915 (N_20915,N_16593,N_15724);
or U20916 (N_20916,N_19333,N_17083);
and U20917 (N_20917,N_16609,N_19551);
and U20918 (N_20918,N_17318,N_17711);
and U20919 (N_20919,N_18714,N_17315);
nand U20920 (N_20920,N_18589,N_19121);
nand U20921 (N_20921,N_15704,N_19484);
nand U20922 (N_20922,N_19768,N_18138);
or U20923 (N_20923,N_17396,N_17261);
and U20924 (N_20924,N_16605,N_16013);
and U20925 (N_20925,N_15921,N_18848);
xnor U20926 (N_20926,N_19486,N_19128);
nor U20927 (N_20927,N_19539,N_16920);
or U20928 (N_20928,N_16460,N_17514);
nand U20929 (N_20929,N_17182,N_19129);
and U20930 (N_20930,N_16512,N_16126);
or U20931 (N_20931,N_17747,N_15896);
and U20932 (N_20932,N_18709,N_19408);
or U20933 (N_20933,N_19776,N_15225);
nor U20934 (N_20934,N_18720,N_15632);
and U20935 (N_20935,N_19445,N_18775);
nand U20936 (N_20936,N_16109,N_15180);
and U20937 (N_20937,N_17433,N_16854);
nor U20938 (N_20938,N_16489,N_16023);
and U20939 (N_20939,N_17454,N_18237);
or U20940 (N_20940,N_19450,N_19842);
nor U20941 (N_20941,N_18258,N_16283);
nand U20942 (N_20942,N_15840,N_15914);
xor U20943 (N_20943,N_17982,N_16260);
xor U20944 (N_20944,N_15265,N_18276);
or U20945 (N_20945,N_18605,N_19751);
and U20946 (N_20946,N_15837,N_19924);
nor U20947 (N_20947,N_16719,N_19533);
nand U20948 (N_20948,N_15307,N_17457);
nor U20949 (N_20949,N_19586,N_19749);
nand U20950 (N_20950,N_19329,N_18656);
or U20951 (N_20951,N_17765,N_17467);
or U20952 (N_20952,N_18550,N_15235);
nor U20953 (N_20953,N_17868,N_18294);
xnor U20954 (N_20954,N_16297,N_19042);
or U20955 (N_20955,N_16291,N_16112);
nor U20956 (N_20956,N_19022,N_17149);
or U20957 (N_20957,N_19015,N_18769);
nor U20958 (N_20958,N_19669,N_18919);
nor U20959 (N_20959,N_15152,N_17147);
nor U20960 (N_20960,N_15167,N_15518);
nand U20961 (N_20961,N_15796,N_15732);
nor U20962 (N_20962,N_18162,N_17644);
nor U20963 (N_20963,N_15269,N_16292);
nor U20964 (N_20964,N_17636,N_17208);
and U20965 (N_20965,N_16583,N_17650);
or U20966 (N_20966,N_16858,N_18090);
and U20967 (N_20967,N_15068,N_19500);
or U20968 (N_20968,N_19204,N_16039);
or U20969 (N_20969,N_19456,N_16399);
or U20970 (N_20970,N_16645,N_16323);
or U20971 (N_20971,N_16142,N_17513);
or U20972 (N_20972,N_19618,N_15778);
or U20973 (N_20973,N_16823,N_15387);
nand U20974 (N_20974,N_18933,N_15994);
or U20975 (N_20975,N_17324,N_19716);
nand U20976 (N_20976,N_16092,N_15008);
or U20977 (N_20977,N_16498,N_18346);
and U20978 (N_20978,N_19688,N_17269);
nor U20979 (N_20979,N_19052,N_17459);
or U20980 (N_20980,N_16681,N_16181);
or U20981 (N_20981,N_18708,N_15168);
or U20982 (N_20982,N_18023,N_16032);
and U20983 (N_20983,N_19957,N_15194);
and U20984 (N_20984,N_17601,N_16510);
nand U20985 (N_20985,N_18744,N_17017);
nand U20986 (N_20986,N_19883,N_18269);
nor U20987 (N_20987,N_17001,N_16740);
nor U20988 (N_20988,N_15430,N_19338);
nand U20989 (N_20989,N_19018,N_19428);
and U20990 (N_20990,N_18716,N_17566);
and U20991 (N_20991,N_18440,N_15426);
or U20992 (N_20992,N_16175,N_17071);
or U20993 (N_20993,N_15947,N_15836);
nand U20994 (N_20994,N_19155,N_18254);
nand U20995 (N_20995,N_16436,N_15800);
xor U20996 (N_20996,N_16259,N_19404);
or U20997 (N_20997,N_18452,N_18878);
nand U20998 (N_20998,N_15037,N_17641);
or U20999 (N_20999,N_19007,N_17897);
xor U21000 (N_21000,N_16483,N_18535);
xnor U21001 (N_21001,N_17733,N_17678);
nor U21002 (N_21002,N_19961,N_19153);
and U21003 (N_21003,N_17508,N_15757);
xnor U21004 (N_21004,N_15564,N_16739);
xnor U21005 (N_21005,N_16931,N_18178);
and U21006 (N_21006,N_19471,N_18363);
nand U21007 (N_21007,N_16020,N_17413);
and U21008 (N_21008,N_18591,N_15856);
nor U21009 (N_21009,N_15617,N_17559);
and U21010 (N_21010,N_17420,N_19708);
nand U21011 (N_21011,N_16316,N_17696);
or U21012 (N_21012,N_16484,N_16315);
and U21013 (N_21013,N_18567,N_15457);
or U21014 (N_21014,N_16829,N_16970);
and U21015 (N_21015,N_17162,N_17991);
nand U21016 (N_21016,N_19555,N_15989);
nor U21017 (N_21017,N_18865,N_16215);
nor U21018 (N_21018,N_16567,N_16885);
nor U21019 (N_21019,N_18700,N_16372);
nand U21020 (N_21020,N_15589,N_15271);
and U21021 (N_21021,N_18244,N_15449);
and U21022 (N_21022,N_17163,N_18745);
nand U21023 (N_21023,N_15382,N_18552);
nor U21024 (N_21024,N_15507,N_17689);
nor U21025 (N_21025,N_19988,N_18447);
nand U21026 (N_21026,N_19150,N_19216);
nand U21027 (N_21027,N_15438,N_15203);
or U21028 (N_21028,N_19188,N_17203);
and U21029 (N_21029,N_18696,N_18551);
and U21030 (N_21030,N_18549,N_17189);
nand U21031 (N_21031,N_15389,N_17263);
nor U21032 (N_21032,N_16848,N_17165);
nor U21033 (N_21033,N_18108,N_16384);
or U21034 (N_21034,N_19443,N_18917);
or U21035 (N_21035,N_15415,N_16800);
nor U21036 (N_21036,N_16912,N_17158);
nand U21037 (N_21037,N_16079,N_19183);
and U21038 (N_21038,N_16148,N_16651);
or U21039 (N_21039,N_18791,N_17426);
or U21040 (N_21040,N_15018,N_17014);
or U21041 (N_21041,N_17725,N_17912);
or U21042 (N_21042,N_15132,N_16004);
xnor U21043 (N_21043,N_15151,N_15321);
and U21044 (N_21044,N_17753,N_17943);
nor U21045 (N_21045,N_15525,N_17293);
or U21046 (N_21046,N_19860,N_15587);
and U21047 (N_21047,N_19828,N_16431);
and U21048 (N_21048,N_15938,N_15466);
or U21049 (N_21049,N_18143,N_16520);
nand U21050 (N_21050,N_17006,N_19414);
and U21051 (N_21051,N_15036,N_18879);
nand U21052 (N_21052,N_18920,N_15535);
nand U21053 (N_21053,N_19689,N_17506);
nor U21054 (N_21054,N_17515,N_15384);
or U21055 (N_21055,N_17997,N_16330);
nor U21056 (N_21056,N_15096,N_18059);
or U21057 (N_21057,N_18733,N_19384);
or U21058 (N_21058,N_19222,N_15157);
nand U21059 (N_21059,N_16680,N_17995);
or U21060 (N_21060,N_17360,N_15875);
or U21061 (N_21061,N_15034,N_16683);
or U21062 (N_21062,N_16137,N_19962);
and U21063 (N_21063,N_15911,N_15996);
or U21064 (N_21064,N_16123,N_15894);
or U21065 (N_21065,N_17431,N_16535);
nand U21066 (N_21066,N_16069,N_18514);
nand U21067 (N_21067,N_18249,N_17545);
nand U21068 (N_21068,N_16972,N_16690);
xnor U21069 (N_21069,N_17598,N_19014);
nand U21070 (N_21070,N_18007,N_19831);
or U21071 (N_21071,N_18491,N_17624);
xnor U21072 (N_21072,N_17134,N_19358);
xor U21073 (N_21073,N_17944,N_19251);
nor U21074 (N_21074,N_17035,N_15027);
nand U21075 (N_21075,N_19021,N_15712);
nand U21076 (N_21076,N_19946,N_17656);
nand U21077 (N_21077,N_16044,N_17914);
or U21078 (N_21078,N_19424,N_15473);
xor U21079 (N_21079,N_17632,N_18371);
and U21080 (N_21080,N_15461,N_16548);
nor U21081 (N_21081,N_18448,N_19314);
or U21082 (N_21082,N_19064,N_16132);
and U21083 (N_21083,N_15357,N_19826);
nand U21084 (N_21084,N_19795,N_19225);
nand U21085 (N_21085,N_17427,N_18149);
or U21086 (N_21086,N_16214,N_19178);
or U21087 (N_21087,N_16257,N_17479);
and U21088 (N_21088,N_18599,N_15729);
or U21089 (N_21089,N_18080,N_17902);
and U21090 (N_21090,N_16009,N_19714);
xnor U21091 (N_21091,N_17880,N_18836);
or U21092 (N_21092,N_16846,N_16461);
nand U21093 (N_21093,N_15218,N_15600);
or U21094 (N_21094,N_18142,N_18033);
or U21095 (N_21095,N_19080,N_18433);
nand U21096 (N_21096,N_19576,N_15420);
nand U21097 (N_21097,N_16642,N_17449);
nor U21098 (N_21098,N_18015,N_17915);
and U21099 (N_21099,N_19899,N_15829);
and U21100 (N_21100,N_19608,N_15575);
or U21101 (N_21101,N_16604,N_18259);
nor U21102 (N_21102,N_17965,N_16636);
nand U21103 (N_21103,N_19663,N_18526);
nand U21104 (N_21104,N_17557,N_15918);
and U21105 (N_21105,N_16221,N_15614);
nand U21106 (N_21106,N_19292,N_15083);
and U21107 (N_21107,N_16694,N_18580);
nand U21108 (N_21108,N_16958,N_18626);
and U21109 (N_21109,N_15356,N_19440);
nand U21110 (N_21110,N_17127,N_15091);
and U21111 (N_21111,N_19614,N_19803);
and U21112 (N_21112,N_15418,N_16442);
xnor U21113 (N_21113,N_15581,N_18047);
and U21114 (N_21114,N_16302,N_18616);
or U21115 (N_21115,N_18054,N_18425);
xnor U21116 (N_21116,N_18844,N_17326);
nand U21117 (N_21117,N_15075,N_17232);
or U21118 (N_21118,N_19973,N_17565);
and U21119 (N_21119,N_17858,N_17347);
xor U21120 (N_21120,N_18343,N_18428);
and U21121 (N_21121,N_17901,N_17058);
xnor U21122 (N_21122,N_18191,N_19874);
or U21123 (N_21123,N_16036,N_17591);
or U21124 (N_21124,N_19793,N_18548);
or U21125 (N_21125,N_18974,N_19770);
nand U21126 (N_21126,N_15118,N_19454);
and U21127 (N_21127,N_17247,N_18721);
nand U21128 (N_21128,N_15405,N_16014);
nor U21129 (N_21129,N_18755,N_16176);
nor U21130 (N_21130,N_15910,N_18562);
or U21131 (N_21131,N_17356,N_18823);
nor U21132 (N_21132,N_17780,N_16808);
nand U21133 (N_21133,N_15232,N_16752);
or U21134 (N_21134,N_17582,N_19727);
nand U21135 (N_21135,N_18833,N_16186);
and U21136 (N_21136,N_17157,N_16709);
and U21137 (N_21137,N_18895,N_19034);
or U21138 (N_21138,N_18688,N_15282);
nor U21139 (N_21139,N_19656,N_19029);
or U21140 (N_21140,N_15465,N_15433);
and U21141 (N_21141,N_15122,N_19020);
or U21142 (N_21142,N_15555,N_19470);
nor U21143 (N_21143,N_17166,N_17669);
nand U21144 (N_21144,N_16325,N_16534);
or U21145 (N_21145,N_18289,N_17547);
or U21146 (N_21146,N_18382,N_16564);
nand U21147 (N_21147,N_19912,N_15215);
nor U21148 (N_21148,N_19662,N_17358);
xor U21149 (N_21149,N_15570,N_18016);
or U21150 (N_21150,N_19661,N_16992);
or U21151 (N_21151,N_18667,N_15365);
nor U21152 (N_21152,N_15140,N_19114);
xor U21153 (N_21153,N_19876,N_16802);
or U21154 (N_21154,N_16434,N_18000);
nor U21155 (N_21155,N_17863,N_19930);
and U21156 (N_21156,N_16334,N_18405);
and U21157 (N_21157,N_17440,N_18645);
nor U21158 (N_21158,N_18542,N_19767);
nor U21159 (N_21159,N_16827,N_18401);
or U21160 (N_21160,N_18052,N_19271);
xnor U21161 (N_21161,N_19743,N_19958);
or U21162 (N_21162,N_15101,N_17469);
and U21163 (N_21163,N_16737,N_16445);
nor U21164 (N_21164,N_18724,N_15644);
and U21165 (N_21165,N_18730,N_16678);
and U21166 (N_21166,N_16458,N_19655);
nor U21167 (N_21167,N_19149,N_15119);
nand U21168 (N_21168,N_18808,N_15826);
and U21169 (N_21169,N_15095,N_18147);
and U21170 (N_21170,N_19938,N_17266);
and U21171 (N_21171,N_17493,N_17697);
nor U21172 (N_21172,N_16172,N_19203);
and U21173 (N_21173,N_19695,N_18991);
nand U21174 (N_21174,N_16528,N_19434);
nand U21175 (N_21175,N_18057,N_15410);
and U21176 (N_21176,N_17768,N_18705);
or U21177 (N_21177,N_19784,N_19270);
nor U21178 (N_21178,N_18959,N_17028);
nor U21179 (N_21179,N_16883,N_16353);
and U21180 (N_21180,N_18664,N_15024);
nand U21181 (N_21181,N_19232,N_18889);
and U21182 (N_21182,N_19634,N_15802);
nor U21183 (N_21183,N_19629,N_16595);
or U21184 (N_21184,N_19298,N_15072);
or U21185 (N_21185,N_16630,N_16702);
and U21186 (N_21186,N_16459,N_19430);
nor U21187 (N_21187,N_15064,N_17251);
or U21188 (N_21188,N_18757,N_15899);
nor U21189 (N_21189,N_18117,N_15469);
and U21190 (N_21190,N_16926,N_16703);
or U21191 (N_21191,N_17906,N_16668);
nor U21192 (N_21192,N_15207,N_15434);
nand U21193 (N_21193,N_17115,N_17987);
nor U21194 (N_21194,N_17934,N_16100);
nor U21195 (N_21195,N_15665,N_16790);
nand U21196 (N_21196,N_15799,N_18155);
nor U21197 (N_21197,N_16162,N_17808);
or U21198 (N_21198,N_15153,N_15604);
nand U21199 (N_21199,N_15517,N_16507);
nand U21200 (N_21200,N_17759,N_18956);
nor U21201 (N_21201,N_18603,N_19569);
and U21202 (N_21202,N_19179,N_17990);
or U21203 (N_21203,N_16954,N_16991);
nor U21204 (N_21204,N_18978,N_19504);
or U21205 (N_21205,N_15155,N_16606);
nor U21206 (N_21206,N_15375,N_16985);
nor U21207 (N_21207,N_17381,N_15677);
nand U21208 (N_21208,N_19399,N_18413);
nand U21209 (N_21209,N_19556,N_16258);
nor U21210 (N_21210,N_17244,N_17130);
nor U21211 (N_21211,N_19606,N_18883);
and U21212 (N_21212,N_16758,N_15508);
nand U21213 (N_21213,N_19667,N_18512);
xor U21214 (N_21214,N_17820,N_19822);
nor U21215 (N_21215,N_19437,N_19841);
xor U21216 (N_21216,N_18832,N_15066);
and U21217 (N_21217,N_18349,N_16207);
nand U21218 (N_21218,N_16361,N_17548);
nor U21219 (N_21219,N_15125,N_18299);
nor U21220 (N_21220,N_19165,N_15076);
or U21221 (N_21221,N_18948,N_19200);
or U21222 (N_21222,N_18909,N_15051);
nand U21223 (N_21223,N_19869,N_19058);
and U21224 (N_21224,N_17010,N_17983);
nand U21225 (N_21225,N_15745,N_16393);
or U21226 (N_21226,N_17707,N_19578);
and U21227 (N_21227,N_16895,N_18527);
or U21228 (N_21228,N_17181,N_19588);
nor U21229 (N_21229,N_16435,N_18439);
or U21230 (N_21230,N_17954,N_16174);
and U21231 (N_21231,N_19491,N_18939);
and U21232 (N_21232,N_19909,N_15751);
or U21233 (N_21233,N_19645,N_16866);
nand U21234 (N_21234,N_19426,N_15017);
and U21235 (N_21235,N_17862,N_17946);
and U21236 (N_21236,N_18801,N_16509);
or U21237 (N_21237,N_16730,N_15630);
or U21238 (N_21238,N_16613,N_15226);
or U21239 (N_21239,N_15997,N_15531);
and U21240 (N_21240,N_19780,N_16347);
and U21241 (N_21241,N_18307,N_19951);
or U21242 (N_21242,N_15571,N_15718);
xnor U21243 (N_21243,N_15585,N_18217);
and U21244 (N_21244,N_19474,N_16198);
nor U21245 (N_21245,N_17988,N_18505);
nor U21246 (N_21246,N_17869,N_18749);
xnor U21247 (N_21247,N_19820,N_17153);
xnor U21248 (N_21248,N_19907,N_18726);
and U21249 (N_21249,N_18481,N_17539);
nand U21250 (N_21250,N_18205,N_18632);
and U21251 (N_21251,N_15684,N_18792);
or U21252 (N_21252,N_16624,N_17680);
or U21253 (N_21253,N_17373,N_18284);
nor U21254 (N_21254,N_18331,N_18902);
nand U21255 (N_21255,N_17013,N_18464);
or U21256 (N_21256,N_18009,N_19254);
and U21257 (N_21257,N_16953,N_16463);
nor U21258 (N_21258,N_19925,N_16433);
nor U21259 (N_21259,N_16994,N_17438);
and U21260 (N_21260,N_18722,N_18297);
nor U21261 (N_21261,N_18483,N_18490);
nand U21262 (N_21262,N_18826,N_18934);
or U21263 (N_21263,N_16523,N_19711);
or U21264 (N_21264,N_19190,N_16633);
or U21265 (N_21265,N_15797,N_19387);
nor U21266 (N_21266,N_16340,N_15672);
or U21267 (N_21267,N_19782,N_18043);
or U21268 (N_21268,N_18543,N_16467);
and U21269 (N_21269,N_16843,N_17881);
xnor U21270 (N_21270,N_19351,N_18446);
and U21271 (N_21271,N_19591,N_18118);
and U21272 (N_21272,N_19541,N_16062);
nand U21273 (N_21273,N_15212,N_18461);
or U21274 (N_21274,N_16753,N_15628);
nand U21275 (N_21275,N_16692,N_16128);
nand U21276 (N_21276,N_19357,N_16596);
nand U21277 (N_21277,N_17925,N_19759);
and U21278 (N_21278,N_16590,N_17741);
or U21279 (N_21279,N_15697,N_15439);
and U21280 (N_21280,N_19008,N_15707);
and U21281 (N_21281,N_16930,N_19644);
nor U21282 (N_21282,N_16255,N_17002);
nor U21283 (N_21283,N_19584,N_19156);
or U21284 (N_21284,N_18195,N_19236);
nand U21285 (N_21285,N_18890,N_19637);
nor U21286 (N_21286,N_15533,N_15378);
nor U21287 (N_21287,N_18980,N_16160);
xnor U21288 (N_21288,N_18594,N_19955);
nor U21289 (N_21289,N_18513,N_17380);
nand U21290 (N_21290,N_19282,N_18960);
nand U21291 (N_21291,N_15085,N_15765);
and U21292 (N_21292,N_19844,N_19911);
and U21293 (N_21293,N_19885,N_17676);
xnor U21294 (N_21294,N_19877,N_16326);
xnor U21295 (N_21295,N_18026,N_18593);
nand U21296 (N_21296,N_16075,N_15795);
nor U21297 (N_21297,N_18436,N_18887);
and U21298 (N_21298,N_16437,N_18809);
nand U21299 (N_21299,N_17505,N_18309);
and U21300 (N_21300,N_18083,N_16786);
or U21301 (N_21301,N_18496,N_16027);
nor U21302 (N_21302,N_16563,N_18581);
and U21303 (N_21303,N_18256,N_18411);
and U21304 (N_21304,N_16284,N_16993);
or U21305 (N_21305,N_17045,N_15233);
and U21306 (N_21306,N_16271,N_17913);
or U21307 (N_21307,N_19654,N_17271);
xnor U21308 (N_21308,N_15263,N_15633);
nor U21309 (N_21309,N_18003,N_19863);
and U21310 (N_21310,N_16423,N_19875);
nand U21311 (N_21311,N_15456,N_18494);
or U21312 (N_21312,N_15988,N_19249);
and U21313 (N_21313,N_18537,N_16837);
or U21314 (N_21314,N_19325,N_16185);
and U21315 (N_21315,N_19490,N_18167);
or U21316 (N_21316,N_19374,N_18012);
nor U21317 (N_21317,N_17752,N_19161);
nand U21318 (N_21318,N_18278,N_15520);
or U21319 (N_21319,N_15460,N_19712);
nor U21320 (N_21320,N_16979,N_19336);
nor U21321 (N_21321,N_17662,N_17384);
nand U21322 (N_21322,N_15693,N_16163);
or U21323 (N_21323,N_16120,N_19122);
and U21324 (N_21324,N_19641,N_19295);
and U21325 (N_21325,N_19942,N_15020);
and U21326 (N_21326,N_19706,N_18668);
or U21327 (N_21327,N_17317,N_15705);
and U21328 (N_21328,N_16003,N_15629);
nor U21329 (N_21329,N_19703,N_17066);
nand U21330 (N_21330,N_18652,N_15590);
and U21331 (N_21331,N_18707,N_16978);
or U21332 (N_21332,N_18133,N_18327);
and U21333 (N_21333,N_17878,N_15615);
nand U21334 (N_21334,N_16299,N_18317);
nor U21335 (N_21335,N_17044,N_18558);
nand U21336 (N_21336,N_15206,N_19224);
nor U21337 (N_21337,N_15081,N_15290);
nand U21338 (N_21338,N_15721,N_16250);
nand U21339 (N_21339,N_15213,N_18038);
nor U21340 (N_21340,N_16095,N_15176);
nand U21341 (N_21341,N_18927,N_18115);
or U21342 (N_21342,N_19865,N_18993);
nand U21343 (N_21343,N_15973,N_16813);
nor U21344 (N_21344,N_15703,N_17437);
xnor U21345 (N_21345,N_18817,N_17841);
and U21346 (N_21346,N_15260,N_15331);
or U21347 (N_21347,N_18723,N_19185);
or U21348 (N_21348,N_17236,N_18750);
and U21349 (N_21349,N_15893,N_17631);
xor U21350 (N_21350,N_18575,N_17766);
and U21351 (N_21351,N_17030,N_19773);
or U21352 (N_21352,N_18829,N_15777);
nor U21353 (N_21353,N_17846,N_17543);
nand U21354 (N_21354,N_18943,N_15441);
or U21355 (N_21355,N_15482,N_19624);
xnor U21356 (N_21356,N_17608,N_15499);
nand U21357 (N_21357,N_15432,N_16852);
or U21358 (N_21358,N_18064,N_18403);
nand U21359 (N_21359,N_17528,N_17834);
nor U21360 (N_21360,N_19836,N_19979);
and U21361 (N_21361,N_17527,N_15547);
xor U21362 (N_21362,N_19380,N_16772);
or U21363 (N_21363,N_15088,N_19231);
or U21364 (N_21364,N_19700,N_17483);
and U21365 (N_21365,N_15039,N_15175);
or U21366 (N_21366,N_16610,N_19921);
or U21367 (N_21367,N_17761,N_15038);
or U21368 (N_21368,N_17556,N_18583);
nor U21369 (N_21369,N_15291,N_17886);
and U21370 (N_21370,N_19413,N_17928);
and U21371 (N_21371,N_19365,N_19718);
or U21372 (N_21372,N_16712,N_15874);
nand U21373 (N_21373,N_16029,N_16444);
and U21374 (N_21374,N_17428,N_15353);
nand U21375 (N_21375,N_17876,N_15315);
and U21376 (N_21376,N_19615,N_19675);
nor U21377 (N_21377,N_15429,N_17969);
or U21378 (N_21378,N_17698,N_16230);
or U21379 (N_21379,N_16247,N_17277);
nand U21380 (N_21380,N_16173,N_15579);
and U21381 (N_21381,N_17274,N_16339);
nor U21382 (N_21382,N_19554,N_19383);
nand U21383 (N_21383,N_18281,N_16472);
nand U21384 (N_21384,N_16166,N_16045);
nand U21385 (N_21385,N_19807,N_19340);
xnor U21386 (N_21386,N_18340,N_17250);
nand U21387 (N_21387,N_16479,N_16466);
or U21388 (N_21388,N_16022,N_15853);
xor U21389 (N_21389,N_15991,N_17818);
nor U21390 (N_21390,N_19783,N_17143);
nor U21391 (N_21391,N_19686,N_15688);
nand U21392 (N_21392,N_19905,N_18888);
nand U21393 (N_21393,N_17241,N_16231);
and U21394 (N_21394,N_15857,N_18691);
nor U21395 (N_21395,N_18983,N_16350);
xnor U21396 (N_21396,N_17569,N_18758);
or U21397 (N_21397,N_18234,N_16016);
nand U21398 (N_21398,N_16398,N_19810);
or U21399 (N_21399,N_18706,N_16801);
nand U21400 (N_21400,N_18684,N_16266);
nand U21401 (N_21401,N_15858,N_15475);
and U21402 (N_21402,N_17336,N_18807);
and U21403 (N_21403,N_19219,N_18565);
and U21404 (N_21404,N_15004,N_15264);
and U21405 (N_21405,N_18767,N_17771);
nand U21406 (N_21406,N_18103,N_16425);
or U21407 (N_21407,N_19223,N_16452);
or U21408 (N_21408,N_17020,N_15502);
and U21409 (N_21409,N_18225,N_19627);
or U21410 (N_21410,N_17114,N_19284);
or U21411 (N_21411,N_15355,N_18128);
nand U21412 (N_21412,N_18393,N_19580);
or U21413 (N_21413,N_18074,N_17856);
and U21414 (N_21414,N_18911,N_19043);
and U21415 (N_21415,N_18136,N_18602);
nand U21416 (N_21416,N_19960,N_17562);
or U21417 (N_21417,N_15706,N_15254);
and U21418 (N_21418,N_19328,N_19862);
xor U21419 (N_21419,N_17589,N_17445);
nor U21420 (N_21420,N_19722,N_16354);
and U21421 (N_21421,N_17874,N_17465);
nor U21422 (N_21422,N_19492,N_19085);
or U21423 (N_21423,N_17405,N_17477);
nand U21424 (N_21424,N_18262,N_19265);
nand U21425 (N_21425,N_17867,N_19528);
or U21426 (N_21426,N_19625,N_16725);
and U21427 (N_21427,N_17948,N_19151);
nor U21428 (N_21428,N_16791,N_16073);
nor U21429 (N_21429,N_15417,N_17864);
xnor U21430 (N_21430,N_16127,N_18923);
nand U21431 (N_21431,N_15806,N_15608);
and U21432 (N_21432,N_19913,N_15123);
nand U21433 (N_21433,N_18260,N_15902);
nor U21434 (N_21434,N_17871,N_15110);
or U21435 (N_21435,N_16751,N_15885);
and U21436 (N_21436,N_15259,N_19478);
and U21437 (N_21437,N_19594,N_16360);
nor U21438 (N_21438,N_15964,N_18470);
and U21439 (N_21439,N_17536,N_19481);
and U21440 (N_21440,N_17772,N_18515);
nor U21441 (N_21441,N_16940,N_16125);
nor U21442 (N_21442,N_18073,N_19433);
and U21443 (N_21443,N_17712,N_18359);
nand U21444 (N_21444,N_19170,N_16981);
or U21445 (N_21445,N_18002,N_15128);
or U21446 (N_21446,N_16919,N_15816);
and U21447 (N_21447,N_16065,N_15760);
xor U21448 (N_21448,N_16966,N_16478);
or U21449 (N_21449,N_16562,N_16611);
or U21450 (N_21450,N_16641,N_15532);
and U21451 (N_21451,N_16441,N_18241);
and U21452 (N_21452,N_16566,N_18037);
or U21453 (N_21453,N_18150,N_17745);
and U21454 (N_21454,N_16475,N_15500);
nand U21455 (N_21455,N_17084,N_16749);
nor U21456 (N_21456,N_18651,N_15386);
or U21457 (N_21457,N_17541,N_16845);
or U21458 (N_21458,N_18233,N_15231);
nand U21459 (N_21459,N_17290,N_18519);
and U21460 (N_21460,N_16454,N_18964);
xnor U21461 (N_21461,N_17246,N_18334);
nand U21462 (N_21462,N_16277,N_17850);
nor U21463 (N_21463,N_15074,N_18639);
or U21464 (N_21464,N_19933,N_19229);
and U21465 (N_21465,N_16421,N_16287);
nand U21466 (N_21466,N_15181,N_15377);
nand U21467 (N_21467,N_19287,N_15121);
or U21468 (N_21468,N_15391,N_15283);
and U21469 (N_21469,N_16286,N_19079);
nor U21470 (N_21470,N_18318,N_17840);
and U21471 (N_21471,N_16743,N_19306);
and U21472 (N_21472,N_15108,N_18215);
nand U21473 (N_21473,N_17146,N_18374);
or U21474 (N_21474,N_17764,N_19630);
and U21475 (N_21475,N_16925,N_18372);
and U21476 (N_21476,N_17615,N_18111);
xor U21477 (N_21477,N_16971,N_19095);
nor U21478 (N_21478,N_17588,N_16319);
xor U21479 (N_21479,N_16072,N_16950);
nand U21480 (N_21480,N_15854,N_19565);
and U21481 (N_21481,N_18274,N_17653);
and U21482 (N_21482,N_17443,N_15974);
and U21483 (N_21483,N_15340,N_19245);
nor U21484 (N_21484,N_19322,N_18729);
or U21485 (N_21485,N_19366,N_16780);
xor U21486 (N_21486,N_17964,N_17604);
and U21487 (N_21487,N_19684,N_17638);
or U21488 (N_21488,N_18189,N_18227);
nor U21489 (N_21489,N_16440,N_17221);
and U21490 (N_21490,N_17673,N_16391);
nor U21491 (N_21491,N_16750,N_17968);
or U21492 (N_21492,N_18200,N_17435);
nand U21493 (N_21493,N_15675,N_18517);
nor U21494 (N_21494,N_17619,N_18835);
or U21495 (N_21495,N_17621,N_17885);
and U21496 (N_21496,N_17173,N_15639);
nor U21497 (N_21497,N_17784,N_17884);
nand U21498 (N_21498,N_19423,N_18265);
and U21499 (N_21499,N_16038,N_16656);
or U21500 (N_21500,N_16874,N_17567);
and U21501 (N_21501,N_19152,N_17849);
nand U21502 (N_21502,N_19390,N_17054);
and U21503 (N_21503,N_18946,N_16377);
and U21504 (N_21504,N_18822,N_17633);
or U21505 (N_21505,N_16355,N_17019);
or U21506 (N_21506,N_18573,N_16046);
nor U21507 (N_21507,N_15141,N_17462);
nand U21508 (N_21508,N_15863,N_19873);
and U21509 (N_21509,N_19568,N_15202);
nand U21510 (N_21510,N_19070,N_19294);
and U21511 (N_21511,N_18966,N_15516);
and U21512 (N_21512,N_15761,N_18858);
nor U21513 (N_21513,N_18082,N_17404);
nor U21514 (N_21514,N_17037,N_16349);
nand U21515 (N_21515,N_18540,N_18145);
and U21516 (N_21516,N_15010,N_17491);
xnor U21517 (N_21517,N_19914,N_18467);
or U21518 (N_21518,N_19054,N_18910);
or U21519 (N_21519,N_19257,N_18140);
nor U21520 (N_21520,N_16119,N_15975);
and U21521 (N_21521,N_15824,N_15972);
and U21522 (N_21522,N_15236,N_16086);
or U21523 (N_21523,N_16655,N_15657);
or U21524 (N_21524,N_17699,N_16465);
and U21525 (N_21525,N_15343,N_15623);
nand U21526 (N_21526,N_19619,N_17935);
or U21527 (N_21527,N_17827,N_16157);
xor U21528 (N_21528,N_18319,N_18682);
or U21529 (N_21529,N_16975,N_17492);
nand U21530 (N_21530,N_19748,N_16769);
and U21531 (N_21531,N_17287,N_17531);
xor U21532 (N_21532,N_16897,N_18030);
or U21533 (N_21533,N_15313,N_18236);
or U21534 (N_21534,N_16091,N_19548);
nor U21535 (N_21535,N_19827,N_16380);
or U21536 (N_21536,N_15030,N_19308);
or U21537 (N_21537,N_18989,N_19573);
and U21538 (N_21538,N_17342,N_19685);
and U21539 (N_21539,N_19730,N_17967);
or U21540 (N_21540,N_17307,N_16107);
and U21541 (N_21541,N_18132,N_17482);
nor U21542 (N_21542,N_19293,N_18341);
or U21543 (N_21543,N_17177,N_15158);
and U21544 (N_21544,N_15606,N_17099);
or U21545 (N_21545,N_17719,N_15813);
nor U21546 (N_21546,N_18511,N_16909);
or U21547 (N_21547,N_19975,N_19389);
nor U21548 (N_21548,N_18577,N_19267);
or U21549 (N_21549,N_16856,N_15305);
nor U21550 (N_21550,N_18434,N_19039);
and U21551 (N_21551,N_19040,N_19892);
nor U21552 (N_21552,N_15515,N_18547);
nand U21553 (N_21553,N_16317,N_17086);
nand U21554 (N_21554,N_17451,N_17352);
xor U21555 (N_21555,N_19467,N_17825);
nor U21556 (N_21556,N_17522,N_16251);
and U21557 (N_21557,N_17094,N_16298);
xnor U21558 (N_21558,N_15689,N_18785);
nand U21559 (N_21559,N_18041,N_16318);
nor U21560 (N_21560,N_18982,N_18824);
and U21561 (N_21561,N_19681,N_17742);
nand U21562 (N_21562,N_15954,N_18477);
or U21563 (N_21563,N_19065,N_19952);
and U21564 (N_21564,N_19646,N_19734);
nor U21565 (N_21565,N_19324,N_16984);
nand U21566 (N_21566,N_17452,N_16121);
nor U21567 (N_21567,N_16216,N_17583);
nand U21568 (N_21568,N_17854,N_16081);
or U21569 (N_21569,N_19834,N_16603);
nor U21570 (N_21570,N_18853,N_15246);
xor U21571 (N_21571,N_17705,N_17296);
nor U21572 (N_21572,N_19062,N_17224);
nor U21573 (N_21573,N_15645,N_18693);
and U21574 (N_21574,N_17739,N_18598);
or U21575 (N_21575,N_18025,N_15339);
and U21576 (N_21576,N_18095,N_17594);
nor U21577 (N_21577,N_18686,N_19761);
nor U21578 (N_21578,N_16409,N_17207);
and U21579 (N_21579,N_15470,N_18210);
nor U21580 (N_21580,N_16068,N_19405);
or U21581 (N_21581,N_15145,N_15241);
or U21582 (N_21582,N_17674,N_19331);
xor U21583 (N_21583,N_16096,N_15820);
or U21584 (N_21584,N_15393,N_18089);
or U21585 (N_21585,N_15166,N_18270);
nor U21586 (N_21586,N_18197,N_18524);
or U21587 (N_21587,N_16151,N_19346);
or U21588 (N_21588,N_16892,N_17095);
and U21589 (N_21589,N_19935,N_17829);
nor U21590 (N_21590,N_16911,N_15933);
and U21591 (N_21591,N_17280,N_18325);
nand U21592 (N_21592,N_19567,N_19260);
nand U21593 (N_21593,N_18704,N_19513);
and U21594 (N_21594,N_19765,N_15514);
nand U21595 (N_21595,N_16179,N_15451);
nand U21596 (N_21596,N_18421,N_15897);
or U21597 (N_21597,N_16000,N_18585);
or U21598 (N_21598,N_18406,N_17429);
and U21599 (N_21599,N_18035,N_19506);
nor U21600 (N_21600,N_16765,N_15078);
nand U21601 (N_21601,N_16946,N_19056);
nor U21602 (N_21602,N_17051,N_17651);
and U21603 (N_21603,N_18772,N_17749);
nor U21604 (N_21604,N_18230,N_19926);
and U21605 (N_21605,N_17321,N_15944);
nand U21606 (N_21606,N_17610,N_17088);
nand U21607 (N_21607,N_17081,N_16311);
or U21608 (N_21608,N_19212,N_19164);
nand U21609 (N_21609,N_19037,N_18500);
and U21610 (N_21610,N_19923,N_17027);
or U21611 (N_21611,N_18112,N_19135);
nand U21612 (N_21612,N_15959,N_17570);
nor U21613 (N_21613,N_16676,N_15929);
xor U21614 (N_21614,N_19941,N_19947);
and U21615 (N_21615,N_18790,N_16432);
and U21616 (N_21616,N_17386,N_16579);
or U21617 (N_21617,N_15295,N_17938);
nor U21618 (N_21618,N_15117,N_16654);
nand U21619 (N_21619,N_16988,N_17407);
nor U21620 (N_21620,N_18286,N_16514);
nor U21621 (N_21621,N_19916,N_18678);
and U21622 (N_21622,N_17721,N_18204);
or U21623 (N_21623,N_15272,N_18876);
nand U21624 (N_21624,N_19731,N_17075);
and U21625 (N_21625,N_19610,N_15557);
xor U21626 (N_21626,N_16446,N_19752);
nand U21627 (N_21627,N_16571,N_18171);
or U21628 (N_21628,N_15831,N_15656);
nor U21629 (N_21629,N_17708,N_15239);
nand U21630 (N_21630,N_17346,N_19323);
xor U21631 (N_21631,N_15257,N_17102);
xor U21632 (N_21632,N_18305,N_16122);
and U21633 (N_21633,N_18928,N_16597);
nor U21634 (N_21634,N_19742,N_17370);
or U21635 (N_21635,N_19256,N_17091);
or U21636 (N_21636,N_17171,N_17119);
xor U21637 (N_21637,N_18607,N_19448);
nor U21638 (N_21638,N_19998,N_15577);
or U21639 (N_21639,N_19880,N_15952);
nor U21640 (N_21640,N_16544,N_19233);
nand U21641 (N_21641,N_17209,N_15710);
and U21642 (N_21642,N_17587,N_17233);
nor U21643 (N_21643,N_19004,N_19986);
nand U21644 (N_21644,N_16254,N_15161);
and U21645 (N_21645,N_19971,N_17300);
xor U21646 (N_21646,N_19530,N_18560);
xor U21647 (N_21647,N_18778,N_15007);
or U21648 (N_21648,N_19321,N_19597);
nand U21649 (N_21649,N_18375,N_18996);
xnor U21650 (N_21650,N_19526,N_16761);
nand U21651 (N_21651,N_19209,N_17285);
nor U21652 (N_21652,N_17773,N_18931);
or U21653 (N_21653,N_15425,N_18990);
nand U21654 (N_21654,N_16074,N_18053);
and U21655 (N_21655,N_16196,N_15436);
and U21656 (N_21656,N_15422,N_16233);
and U21657 (N_21657,N_15766,N_17478);
nor U21658 (N_21658,N_18592,N_16607);
nor U21659 (N_21659,N_17025,N_19557);
or U21660 (N_21660,N_17652,N_17000);
and U21661 (N_21661,N_18498,N_16253);
or U21662 (N_21662,N_15255,N_18872);
nor U21663 (N_21663,N_17473,N_15917);
or U21664 (N_21664,N_17612,N_19116);
xnor U21665 (N_21665,N_15651,N_18587);
or U21666 (N_21666,N_18545,N_17257);
and U21667 (N_21667,N_16376,N_18814);
nand U21668 (N_21668,N_15371,N_16352);
and U21669 (N_21669,N_15193,N_19804);
xnor U21670 (N_21670,N_16263,N_18148);
nor U21671 (N_21671,N_15172,N_18427);
nand U21672 (N_21672,N_19632,N_18711);
nor U21673 (N_21673,N_16674,N_16276);
and U21674 (N_21674,N_16980,N_18811);
nand U21675 (N_21675,N_17339,N_19134);
and U21676 (N_21676,N_18779,N_15671);
and U21677 (N_21677,N_16516,N_15683);
nor U21678 (N_21678,N_15079,N_18838);
or U21679 (N_21679,N_19520,N_17959);
and U21680 (N_21680,N_18458,N_18942);
xor U21681 (N_21681,N_17395,N_19697);
nor U21682 (N_21682,N_16587,N_17126);
or U21683 (N_21683,N_19320,N_19690);
and U21684 (N_21684,N_16558,N_17578);
nor U21685 (N_21685,N_17041,N_18915);
nor U21686 (N_21686,N_15738,N_18582);
and U21687 (N_21687,N_18300,N_18834);
and U21688 (N_21688,N_19977,N_19993);
and U21689 (N_21689,N_19201,N_19636);
and U21690 (N_21690,N_15216,N_19246);
or U21691 (N_21691,N_16957,N_15898);
and U21692 (N_21692,N_18386,N_18330);
nand U21693 (N_21693,N_16180,N_15444);
and U21694 (N_21694,N_15771,N_17453);
or U21695 (N_21695,N_19373,N_17803);
or U21696 (N_21696,N_19420,N_19137);
nor U21697 (N_21697,N_17468,N_15883);
nor U21698 (N_21698,N_19522,N_15210);
or U21699 (N_21699,N_15124,N_15702);
nor U21700 (N_21700,N_16001,N_18388);
nor U21701 (N_21701,N_17359,N_15144);
nor U21702 (N_21702,N_17248,N_15028);
nor U21703 (N_21703,N_16116,N_18747);
nor U21704 (N_21704,N_15828,N_18584);
nand U21705 (N_21705,N_17466,N_17184);
nor U21706 (N_21706,N_16860,N_15513);
nand U21707 (N_21707,N_18929,N_19510);
or U21708 (N_21708,N_16412,N_16373);
nand U21709 (N_21709,N_17053,N_18180);
and U21710 (N_21710,N_17677,N_18597);
nor U21711 (N_21711,N_16531,N_17561);
and U21712 (N_21712,N_17634,N_19781);
nand U21713 (N_21713,N_17372,N_15980);
and U21714 (N_21714,N_15506,N_18908);
or U21715 (N_21715,N_15077,N_17180);
or U21716 (N_21716,N_19436,N_15476);
and U21717 (N_21717,N_18376,N_19967);
nand U21718 (N_21718,N_19379,N_15044);
nand U21719 (N_21719,N_16932,N_18160);
and U21720 (N_21720,N_17838,N_19010);
or U21721 (N_21721,N_15638,N_17371);
or U21722 (N_21722,N_18209,N_16934);
or U21723 (N_21723,N_19764,N_19097);
nor U21724 (N_21724,N_16168,N_18683);
nor U21725 (N_21725,N_15635,N_18092);
and U21726 (N_21726,N_17310,N_17821);
and U21727 (N_21727,N_18242,N_19642);
and U21728 (N_21728,N_15102,N_16947);
or U21729 (N_21729,N_19939,N_16647);
or U21730 (N_21730,N_16124,N_15530);
nor U21731 (N_21731,N_18042,N_16031);
nor U21732 (N_21732,N_15033,N_15459);
xor U21733 (N_21733,N_19162,N_19895);
nor U21734 (N_21734,N_15850,N_17781);
nor U21735 (N_21735,N_18086,N_15887);
nor U21736 (N_21736,N_18441,N_15002);
or U21737 (N_21737,N_17082,N_19890);
and U21738 (N_21738,N_19259,N_16321);
nand U21739 (N_21739,N_19483,N_15937);
or U21740 (N_21740,N_18385,N_15505);
nor U21741 (N_21741,N_15984,N_19707);
nor U21742 (N_21742,N_19286,N_15868);
nor U21743 (N_21743,N_17298,N_16468);
nand U21744 (N_21744,N_15780,N_18783);
nor U21745 (N_21745,N_15888,N_15733);
or U21746 (N_21746,N_17893,N_15616);
nor U21747 (N_21747,N_19540,N_18731);
and U21748 (N_21748,N_15277,N_15187);
nor U21749 (N_21749,N_19887,N_15164);
nor U21750 (N_21750,N_15069,N_16150);
nand U21751 (N_21751,N_15421,N_15713);
or U21752 (N_21752,N_17540,N_16582);
or U21753 (N_21753,N_18169,N_17446);
nand U21754 (N_21754,N_19829,N_15655);
nand U21755 (N_21755,N_16569,N_15303);
nand U21756 (N_21756,N_16840,N_16700);
and U21757 (N_21757,N_18445,N_17291);
or U21758 (N_21758,N_16464,N_18024);
nand U21759 (N_21759,N_17168,N_16987);
or U21760 (N_21760,N_19143,N_18011);
and U21761 (N_21761,N_15323,N_15528);
and U21762 (N_21762,N_15605,N_17108);
nor U21763 (N_21763,N_19305,N_18497);
or U21764 (N_21764,N_19677,N_18912);
and U21765 (N_21765,N_17008,N_17552);
and U21766 (N_21766,N_15287,N_16282);
nor U21767 (N_21767,N_18859,N_17883);
and U21768 (N_21768,N_19100,N_16736);
and U21769 (N_21769,N_16480,N_17316);
nand U21770 (N_21770,N_19395,N_19801);
nand U21771 (N_21771,N_18976,N_17185);
and U21772 (N_21772,N_17716,N_18987);
nor U21773 (N_21773,N_17363,N_19997);
nor U21774 (N_21774,N_15546,N_17199);
or U21775 (N_21775,N_18986,N_17414);
nand U21776 (N_21776,N_15266,N_17012);
nand U21777 (N_21777,N_15536,N_17292);
nor U21778 (N_21778,N_18967,N_17812);
and U21779 (N_21779,N_16342,N_17802);
or U21780 (N_21780,N_17461,N_18559);
and U21781 (N_21781,N_15093,N_16541);
xnor U21782 (N_21782,N_18004,N_18367);
and U21783 (N_21783,N_16857,N_16113);
nand U21784 (N_21784,N_16723,N_16131);
nor U21785 (N_21785,N_17132,N_18312);
or U21786 (N_21786,N_17617,N_17421);
and U21787 (N_21787,N_15120,N_17376);
and U21788 (N_21788,N_15978,N_19023);
nand U21789 (N_21789,N_18675,N_18676);
nand U21790 (N_21790,N_17585,N_18689);
xnor U21791 (N_21791,N_17516,N_18290);
and U21792 (N_21792,N_15995,N_19515);
nor U21793 (N_21793,N_18687,N_15949);
nor U21794 (N_21794,N_16218,N_16870);
and U21795 (N_21795,N_15165,N_16490);
nor U21796 (N_21796,N_16366,N_18212);
and U21797 (N_21797,N_16397,N_18034);
and U21798 (N_21798,N_16387,N_15558);
or U21799 (N_21799,N_19552,N_18006);
nor U21800 (N_21800,N_17979,N_15967);
nor U21801 (N_21801,N_17597,N_19721);
nand U21802 (N_21802,N_15362,N_18892);
xor U21803 (N_21803,N_19900,N_19523);
and U21804 (N_21804,N_16243,N_15886);
and U21805 (N_21805,N_18192,N_17228);
nor U21806 (N_21806,N_16555,N_15053);
nand U21807 (N_21807,N_15912,N_15440);
and U21808 (N_21808,N_15240,N_15529);
nand U21809 (N_21809,N_19771,N_19359);
or U21810 (N_21810,N_17936,N_16760);
and U21811 (N_21811,N_19949,N_16141);
or U21812 (N_21812,N_18572,N_19345);
or U21813 (N_21813,N_19800,N_16099);
nand U21814 (N_21814,N_19009,N_17214);
nor U21815 (N_21815,N_17159,N_15348);
nor U21816 (N_21816,N_17900,N_17278);
nand U21817 (N_21817,N_18529,N_16164);
and U21818 (N_21818,N_17681,N_19992);
nor U21819 (N_21819,N_15406,N_16402);
and U21820 (N_21820,N_17932,N_18101);
nand U21821 (N_21821,N_18637,N_16256);
or U21822 (N_21822,N_17385,N_19590);
nand U21823 (N_21823,N_17503,N_18630);
nor U21824 (N_21824,N_15390,N_16064);
nor U21825 (N_21825,N_15871,N_17888);
and U21826 (N_21826,N_19762,N_19701);
and U21827 (N_21827,N_17104,N_16806);
or U21828 (N_21828,N_16097,N_15214);
nand U21829 (N_21829,N_16332,N_17256);
and U21830 (N_21830,N_17788,N_17098);
and U21831 (N_21831,N_16648,N_17970);
and U21832 (N_21832,N_16504,N_15951);
or U21833 (N_21833,N_19889,N_16077);
nand U21834 (N_21834,N_16685,N_19693);
or U21835 (N_21835,N_19353,N_17684);
xor U21836 (N_21836,N_19463,N_17622);
and U21837 (N_21837,N_15032,N_19746);
or U21838 (N_21838,N_18453,N_16201);
xnor U21839 (N_21839,N_18638,N_16913);
and U21840 (N_21840,N_16019,N_18766);
or U21841 (N_21841,N_19871,N_19983);
and U21842 (N_21842,N_18301,N_17581);
nor U21843 (N_21843,N_16561,N_17643);
nor U21844 (N_21844,N_15173,N_17063);
nor U21845 (N_21845,N_15726,N_16974);
nor U21846 (N_21846,N_16085,N_16296);
and U21847 (N_21847,N_19872,N_16626);
and U21848 (N_21848,N_16511,N_16775);
nor U21849 (N_21849,N_19461,N_15835);
nor U21850 (N_21850,N_18144,N_17295);
and U21851 (N_21851,N_16426,N_15105);
nor U21852 (N_21852,N_17637,N_17830);
xnor U21853 (N_21853,N_19485,N_19310);
nor U21854 (N_21854,N_15474,N_15872);
or U21855 (N_21855,N_17630,N_18324);
or U21856 (N_21856,N_17021,N_16227);
or U21857 (N_21857,N_15403,N_19598);
nand U21858 (N_21858,N_17956,N_19189);
xor U21859 (N_21859,N_18292,N_15969);
or U21860 (N_21860,N_18786,N_19166);
and U21861 (N_21861,N_15698,N_17434);
nor U21862 (N_21862,N_16834,N_17629);
or U21863 (N_21863,N_17989,N_18369);
nor U21864 (N_21864,N_17161,N_15822);
and U21865 (N_21865,N_15652,N_15054);
nor U21866 (N_21866,N_18701,N_16057);
and U21867 (N_21867,N_19732,N_15442);
and U21868 (N_21868,N_18482,N_15211);
and U21869 (N_21869,N_19000,N_17351);
nand U21870 (N_21870,N_18431,N_17899);
nand U21871 (N_21871,N_15458,N_15730);
xor U21872 (N_21872,N_16274,N_15881);
nand U21873 (N_21873,N_19595,N_17499);
or U21874 (N_21874,N_18619,N_16047);
and U21875 (N_21875,N_18358,N_16115);
nor U21876 (N_21876,N_16959,N_19616);
nand U21877 (N_21877,N_17488,N_19417);
xnor U21878 (N_21878,N_16364,N_17792);
or U21879 (N_21879,N_15381,N_17322);
nor U21880 (N_21880,N_15129,N_18532);
nand U21881 (N_21881,N_19449,N_15022);
and U21882 (N_21882,N_17568,N_18251);
or U21883 (N_21883,N_16720,N_19794);
nor U21884 (N_21884,N_16167,N_19255);
nand U21885 (N_21885,N_19464,N_15512);
and U21886 (N_21886,N_17485,N_15005);
and U21887 (N_21887,N_15395,N_16090);
or U21888 (N_21888,N_17329,N_16470);
nand U21889 (N_21889,N_15424,N_19791);
or U21890 (N_21890,N_19197,N_18738);
nand U21891 (N_21891,N_15450,N_16533);
or U21892 (N_21892,N_16689,N_15924);
or U21893 (N_21893,N_15443,N_16908);
xor U21894 (N_21894,N_18426,N_17056);
nor U21895 (N_21895,N_19934,N_18753);
nor U21896 (N_21896,N_16264,N_19277);
and U21897 (N_21897,N_19352,N_18165);
nor U21898 (N_21898,N_18944,N_15838);
nor U21899 (N_21899,N_16028,N_15562);
or U21900 (N_21900,N_16653,N_17043);
xnor U21901 (N_21901,N_17410,N_16522);
or U21902 (N_21902,N_18492,N_18198);
xor U21903 (N_21903,N_17152,N_16951);
nand U21904 (N_21904,N_18849,N_18851);
or U21905 (N_21905,N_18079,N_19867);
or U21906 (N_21906,N_19071,N_19281);
or U21907 (N_21907,N_17661,N_16631);
or U21908 (N_21908,N_19717,N_16219);
nor U21909 (N_21909,N_17791,N_17070);
nor U21910 (N_21910,N_15509,N_18306);
nor U21911 (N_21911,N_18442,N_19107);
and U21912 (N_21912,N_16614,N_17062);
xor U21913 (N_21913,N_19953,N_19753);
nor U21914 (N_21914,N_19131,N_17775);
and U21915 (N_21915,N_18795,N_19665);
and U21916 (N_21916,N_17004,N_19680);
nor U21917 (N_21917,N_19702,N_17521);
xnor U21918 (N_21918,N_16136,N_15297);
and U21919 (N_21919,N_18864,N_15556);
nand U21920 (N_21920,N_17123,N_18159);
nor U21921 (N_21921,N_15394,N_17069);
or U21922 (N_21922,N_17128,N_17769);
nor U21923 (N_21923,N_15237,N_15843);
nor U21924 (N_21924,N_19142,N_16933);
nand U21925 (N_21925,N_19136,N_17501);
nand U21926 (N_21926,N_16638,N_18875);
nand U21927 (N_21927,N_15830,N_19217);
or U21928 (N_21928,N_15437,N_18355);
nand U21929 (N_21929,N_17972,N_19518);
and U21930 (N_21930,N_15368,N_16635);
and U21931 (N_21931,N_17230,N_17623);
or U21932 (N_21932,N_15869,N_15059);
xor U21933 (N_21933,N_16088,N_18398);
nor U21934 (N_21934,N_18669,N_17958);
and U21935 (N_21935,N_17379,N_16506);
nor U21936 (N_21936,N_19303,N_19047);
or U21937 (N_21937,N_16049,N_15641);
and U21938 (N_21938,N_15876,N_18186);
xnor U21939 (N_21939,N_17460,N_16560);
nor U21940 (N_21940,N_16968,N_19473);
nand U21941 (N_21941,N_17801,N_18456);
or U21942 (N_21942,N_15583,N_15742);
nor U21943 (N_21943,N_19123,N_17155);
or U21944 (N_21944,N_16191,N_15097);
and U21945 (N_21945,N_17966,N_18615);
nand U21946 (N_21946,N_15634,N_19631);
nand U21947 (N_21947,N_17220,N_18193);
or U21948 (N_21948,N_16661,N_18840);
nand U21949 (N_21949,N_18608,N_17718);
and U21950 (N_21950,N_16161,N_18566);
and U21951 (N_21951,N_18027,N_16711);
nor U21952 (N_21952,N_17268,N_17378);
nand U21953 (N_21953,N_18539,N_17367);
nand U21954 (N_21954,N_15553,N_18085);
or U21955 (N_21955,N_16650,N_17500);
or U21956 (N_21956,N_18623,N_19830);
nand U21957 (N_21957,N_17117,N_16696);
and U21958 (N_21958,N_15138,N_17187);
or U21959 (N_21959,N_18857,N_19757);
and U21960 (N_21960,N_17399,N_17957);
and U21961 (N_21961,N_16129,N_16403);
nor U21962 (N_21962,N_17584,N_19234);
nor U21963 (N_21963,N_19769,N_19089);
nor U21964 (N_21964,N_19995,N_17534);
xnor U21965 (N_21965,N_18874,N_17758);
xnor U21966 (N_21966,N_16697,N_18499);
nand U21967 (N_21967,N_19041,N_15178);
and U21968 (N_21968,N_18741,N_19855);
or U21969 (N_21969,N_16581,N_16773);
or U21970 (N_21970,N_19861,N_15491);
or U21971 (N_21971,N_16002,N_17790);
or U21972 (N_21972,N_19392,N_15741);
or U21973 (N_21973,N_17472,N_19451);
or U21974 (N_21974,N_19174,N_18063);
or U21975 (N_21975,N_15774,N_17487);
xor U21976 (N_21976,N_16204,N_15786);
nor U21977 (N_21977,N_19817,N_18032);
nor U21978 (N_21978,N_19534,N_16138);
or U21979 (N_21979,N_18907,N_17489);
xor U21980 (N_21980,N_18614,N_16999);
xnor U21981 (N_21981,N_16815,N_15668);
xor U21982 (N_21982,N_18521,N_15699);
and U21983 (N_21983,N_19823,N_19710);
and U21984 (N_21984,N_17172,N_15261);
nand U21985 (N_21985,N_16305,N_15367);
nor U21986 (N_21986,N_17327,N_15798);
or U21987 (N_21987,N_18629,N_19521);
nor U21988 (N_21988,N_19833,N_18219);
nor U21989 (N_21989,N_18071,N_15815);
and U21990 (N_21990,N_19237,N_18843);
or U21991 (N_21991,N_17464,N_16764);
or U21992 (N_21992,N_15050,N_16153);
or U21993 (N_21993,N_16050,N_18725);
or U21994 (N_21994,N_19572,N_17654);
or U21995 (N_21995,N_16708,N_17895);
and U21996 (N_21996,N_17226,N_17325);
nor U21997 (N_21997,N_15301,N_17875);
nor U21998 (N_21998,N_16208,N_15573);
nor U21999 (N_21999,N_17286,N_17369);
nor U22000 (N_22000,N_15756,N_19280);
and U22001 (N_22001,N_17542,N_16741);
and U22002 (N_22002,N_16220,N_16546);
and U22003 (N_22003,N_18127,N_16415);
nor U22004 (N_22004,N_17596,N_16722);
or U22005 (N_22005,N_19416,N_18046);
and U22006 (N_22006,N_17496,N_15501);
nand U22007 (N_22007,N_16206,N_19674);
xnor U22008 (N_22008,N_16382,N_17455);
or U22009 (N_22009,N_17770,N_17237);
nor U22010 (N_22010,N_19475,N_17533);
and U22011 (N_22011,N_15063,N_15753);
or U22012 (N_22012,N_17312,N_17853);
and U22013 (N_22013,N_16105,N_18612);
or U22014 (N_22014,N_16439,N_18789);
and U22015 (N_22015,N_19177,N_15169);
nand U22016 (N_22016,N_19048,N_19740);
and U22017 (N_22017,N_19811,N_18520);
nor U22018 (N_22018,N_16640,N_16262);
nor U22019 (N_22019,N_19427,N_18170);
nor U22020 (N_22020,N_15889,N_19666);
or U22021 (N_22021,N_15782,N_16346);
nand U22022 (N_22022,N_15865,N_18648);
or U22023 (N_22023,N_15903,N_18416);
nand U22024 (N_22024,N_18125,N_15400);
and U22025 (N_22025,N_18703,N_19111);
or U22026 (N_22026,N_19238,N_18613);
nor U22027 (N_22027,N_19110,N_17573);
nor U22028 (N_22028,N_19438,N_17737);
nor U22029 (N_22029,N_15970,N_15049);
nor U22030 (N_22030,N_18861,N_19036);
nand U22031 (N_22031,N_15174,N_15682);
and U22032 (N_22032,N_15673,N_15827);
nand U22033 (N_22033,N_17179,N_19651);
and U22034 (N_22034,N_17176,N_18533);
nand U22035 (N_22035,N_16578,N_18362);
nand U22036 (N_22036,N_15112,N_18029);
or U22037 (N_22037,N_17724,N_19929);
or U22038 (N_22038,N_19335,N_18373);
or U22039 (N_22039,N_19840,N_16418);
and U22040 (N_22040,N_15190,N_17366);
nor U22041 (N_22041,N_16010,N_19272);
and U22042 (N_22042,N_15986,N_18621);
nor U22043 (N_22043,N_19412,N_16159);
nand U22044 (N_22044,N_15597,N_18356);
nand U22045 (N_22045,N_17061,N_17848);
nand U22046 (N_22046,N_18803,N_15147);
xnor U22047 (N_22047,N_15116,N_16171);
or U22048 (N_22048,N_15927,N_16727);
xnor U22049 (N_22049,N_18110,N_15312);
nand U22050 (N_22050,N_16809,N_17710);
nand U22051 (N_22051,N_16358,N_17714);
and U22052 (N_22052,N_15661,N_17456);
or U22053 (N_22053,N_16659,N_16406);
nor U22054 (N_22054,N_19172,N_16395);
and U22055 (N_22055,N_17080,N_17659);
nand U22056 (N_22056,N_19687,N_19772);
nor U22057 (N_22057,N_16042,N_15740);
nand U22058 (N_22058,N_17474,N_18001);
and U22059 (N_22059,N_17393,N_17073);
nand U22060 (N_22060,N_15335,N_19738);
nor U22061 (N_22061,N_18380,N_18752);
nor U22062 (N_22062,N_19715,N_19108);
nand U22063 (N_22063,N_19918,N_15913);
nand U22064 (N_22064,N_19059,N_16621);
and U22065 (N_22065,N_16054,N_17186);
and U22066 (N_22066,N_19525,N_15497);
nor U22067 (N_22067,N_19264,N_18474);
or U22068 (N_22068,N_18134,N_17131);
nand U22069 (N_22069,N_19248,N_16763);
nor U22070 (N_22070,N_15791,N_17799);
nand U22071 (N_22071,N_17323,N_17704);
nor U22072 (N_22072,N_19813,N_15042);
xor U22073 (N_22073,N_17903,N_18352);
nand U22074 (N_22074,N_17520,N_19227);
or U22075 (N_22075,N_16944,N_18067);
and U22076 (N_22076,N_18214,N_15332);
xnor U22077 (N_22077,N_15280,N_17463);
nand U22078 (N_22078,N_16598,N_18930);
xnor U22079 (N_22079,N_18762,N_18296);
or U22080 (N_22080,N_15223,N_18871);
or U22081 (N_22081,N_15568,N_15369);
and U22082 (N_22082,N_16664,N_19069);
nand U22083 (N_22083,N_15818,N_18443);
nand U22084 (N_22084,N_19012,N_17898);
xnor U22085 (N_22085,N_16983,N_15523);
and U22086 (N_22086,N_18218,N_15327);
xnor U22087 (N_22087,N_16130,N_19051);
nand U22088 (N_22088,N_17319,N_15976);
xnor U22089 (N_22089,N_17422,N_19972);
or U22090 (N_22090,N_17974,N_15379);
xor U22091 (N_22091,N_19719,N_17550);
nand U22092 (N_22092,N_19242,N_17100);
nand U22093 (N_22093,N_17831,N_19319);
nor U22094 (N_22094,N_19682,N_16135);
nand U22095 (N_22095,N_18666,N_19318);
xnor U22096 (N_22096,N_18407,N_18404);
nand U22097 (N_22097,N_17595,N_18435);
nor U22098 (N_22098,N_18065,N_19307);
xnor U22099 (N_22099,N_18516,N_17865);
nor U22100 (N_22100,N_19057,N_19158);
nand U22101 (N_22101,N_15596,N_17701);
or U22102 (N_22102,N_15565,N_18600);
or U22103 (N_22103,N_19072,N_15860);
nor U22104 (N_22104,N_19330,N_15814);
nor U22105 (N_22105,N_19563,N_16568);
nand U22106 (N_22106,N_17423,N_17216);
or U22107 (N_22107,N_17762,N_15563);
or U22108 (N_22108,N_16293,N_17340);
nor U22109 (N_22109,N_19517,N_18839);
or U22110 (N_22110,N_17549,N_16430);
and U22111 (N_22111,N_16835,N_15204);
nand U22112 (N_22112,N_18754,N_18680);
nor U22113 (N_22113,N_18123,N_19622);
xnor U22114 (N_22114,N_15304,N_16080);
nor U22115 (N_22115,N_15773,N_17087);
and U22116 (N_22116,N_19789,N_15146);
nor U22117 (N_22117,N_16103,N_17254);
nor U22118 (N_22118,N_19819,N_17238);
or U22119 (N_22119,N_18588,N_18743);
and U22120 (N_22120,N_15845,N_15990);
or U22121 (N_22121,N_17592,N_16776);
nor U22122 (N_22122,N_15319,N_15767);
nor U22123 (N_22123,N_16041,N_18885);
or U22124 (N_22124,N_15446,N_15333);
nand U22125 (N_22125,N_15607,N_18175);
nand U22126 (N_22126,N_19472,N_19996);
nand U22127 (N_22127,N_18570,N_18129);
nor U22128 (N_22128,N_16565,N_15275);
or U22129 (N_22129,N_17409,N_19139);
nand U22130 (N_22130,N_17235,N_17924);
nand U22131 (N_22131,N_19206,N_15099);
nor U22132 (N_22132,N_19157,N_17332);
nor U22133 (N_22133,N_17814,N_19205);
and U22134 (N_22134,N_17571,N_18793);
or U22135 (N_22135,N_16921,N_18228);
nor U22136 (N_22136,N_17985,N_17767);
nor U22137 (N_22137,N_16660,N_19337);
nor U22138 (N_22138,N_17937,N_15113);
nor U22139 (N_22139,N_18531,N_17911);
xor U22140 (N_22140,N_17136,N_19191);
nand U22141 (N_22141,N_19367,N_17851);
nand U22142 (N_22142,N_16715,N_15709);
or U22143 (N_22143,N_19502,N_16473);
xnor U22144 (N_22144,N_18827,N_18882);
and U22145 (N_22145,N_15230,N_16106);
nor U22146 (N_22146,N_18010,N_18420);
or U22147 (N_22147,N_19002,N_15895);
nand U22148 (N_22148,N_17519,N_17919);
or U22149 (N_22149,N_16570,N_15320);
nand U22150 (N_22150,N_19943,N_18460);
xor U22151 (N_22151,N_19446,N_16371);
and U22152 (N_22152,N_15852,N_15309);
nor U22153 (N_22153,N_19802,N_19974);
nand U22154 (N_22154,N_18124,N_16401);
and U22155 (N_22155,N_19075,N_19066);
xnor U22156 (N_22156,N_17335,N_19053);
nand U22157 (N_22157,N_15743,N_19496);
and U22158 (N_22158,N_18323,N_19989);
nor U22159 (N_22159,N_17510,N_18953);
nor U22160 (N_22160,N_19388,N_17049);
nor U22161 (N_22161,N_15337,N_15992);
nor U22162 (N_22162,N_16748,N_17602);
nor U22163 (N_22163,N_17558,N_16686);
nand U22164 (N_22164,N_16496,N_15720);
and U22165 (N_22165,N_16677,N_16591);
nor U22166 (N_22166,N_15736,N_17798);
nor U22167 (N_22167,N_15014,N_17809);
nand U22168 (N_22168,N_17691,N_15789);
nor U22169 (N_22169,N_16588,N_18121);
nand U22170 (N_22170,N_18802,N_18345);
nand U22171 (N_22171,N_16910,N_16389);
or U22172 (N_22172,N_18867,N_17645);
or U22173 (N_22173,N_17079,N_19210);
nor U22174 (N_22174,N_19476,N_18963);
nand U22175 (N_22175,N_18951,N_18336);
or U22176 (N_22176,N_15341,N_15543);
xor U22177 (N_22177,N_16487,N_17306);
nor U22178 (N_22178,N_15454,N_16873);
and U22179 (N_22179,N_18685,N_18798);
xnor U22180 (N_22180,N_17996,N_15143);
nand U22181 (N_22181,N_15537,N_18732);
and U22182 (N_22182,N_17889,N_19127);
xor U22183 (N_22183,N_16525,N_18486);
nand U22184 (N_22184,N_17476,N_15592);
xor U22185 (N_22185,N_19945,N_17154);
and U22186 (N_22186,N_18658,N_15270);
nand U22187 (N_22187,N_17828,N_17688);
nand U22188 (N_22188,N_15186,N_18308);
or U22189 (N_22189,N_17670,N_18640);
and U22190 (N_22190,N_19133,N_18574);
and U22191 (N_22191,N_19602,N_19275);
and U22192 (N_22192,N_15090,N_18240);
or U22193 (N_22193,N_18863,N_16777);
nor U22194 (N_22194,N_19418,N_16917);
or U22195 (N_22195,N_18774,N_17580);
and U22196 (N_22196,N_18800,N_19901);
nor U22197 (N_22197,N_16192,N_17211);
nor U22198 (N_22198,N_16807,N_18606);
or U22199 (N_22199,N_15539,N_16453);
or U22200 (N_22200,N_15621,N_17344);
and U22201 (N_22201,N_17945,N_18036);
and U22202 (N_22202,N_17215,N_17748);
or U22203 (N_22203,N_15626,N_15934);
or U22204 (N_22204,N_19493,N_19398);
and U22205 (N_22205,N_16850,N_18977);
or U22206 (N_22206,N_17599,N_15278);
nor U22207 (N_22207,N_17447,N_17605);
xnor U22208 (N_22208,N_16070,N_16675);
or U22209 (N_22209,N_15322,N_17694);
nand U22210 (N_22210,N_15071,N_19285);
nor U22211 (N_22211,N_19144,N_16779);
and U22212 (N_22212,N_18383,N_19917);
nor U22213 (N_22213,N_18962,N_16828);
nand U22214 (N_22214,N_17509,N_15708);
and U22215 (N_22215,N_15196,N_18918);
nor U22216 (N_22216,N_17218,N_16554);
xnor U22217 (N_22217,N_15198,N_16880);
and U22218 (N_22218,N_16811,N_15620);
and U22219 (N_22219,N_18609,N_19848);
or U22220 (N_22220,N_19289,N_15376);
nand U22221 (N_22221,N_16898,N_17795);
nand U22222 (N_22222,N_16063,N_19074);
nor U22223 (N_22223,N_17258,N_15618);
or U22224 (N_22224,N_15803,N_17842);
or U22225 (N_22225,N_16798,N_18229);
and U22226 (N_22226,N_18985,N_16154);
nand U22227 (N_22227,N_18084,N_16771);
and U22228 (N_22228,N_18122,N_19728);
and U22229 (N_22229,N_19101,N_16868);
nor U22230 (N_22230,N_16301,N_16228);
or U22231 (N_22231,N_18450,N_17971);
or U22232 (N_22232,N_17245,N_15792);
nor U22233 (N_22233,N_15663,N_17033);
nor U22234 (N_22234,N_16986,N_17067);
and U22235 (N_22235,N_19240,N_15811);
or U22236 (N_22236,N_15182,N_16632);
or U22237 (N_22237,N_18765,N_17709);
and U22238 (N_22238,N_15922,N_16232);
nor U22239 (N_22239,N_18168,N_16787);
and U22240 (N_22240,N_17574,N_17530);
nand U22241 (N_22241,N_15358,N_15939);
xnor U22242 (N_22242,N_18556,N_16385);
nor U22243 (N_22243,N_16889,N_19574);
nor U22244 (N_22244,N_16521,N_18842);
nor U22245 (N_22245,N_17032,N_18784);
and U22246 (N_22246,N_16390,N_18886);
nor U22247 (N_22247,N_19812,N_15380);
nand U22248 (N_22248,N_16245,N_16477);
and U22249 (N_22249,N_17981,N_17921);
nor U22250 (N_22250,N_18207,N_18283);
or U22251 (N_22251,N_16547,N_15901);
nand U22252 (N_22252,N_16795,N_17052);
and U22253 (N_22253,N_19664,N_15317);
nor U22254 (N_22254,N_18051,N_19309);
nor U22255 (N_22255,N_17105,N_16871);
nand U22256 (N_22256,N_15156,N_16118);
or U22257 (N_22257,N_17816,N_19148);
nand U22258 (N_22258,N_17212,N_16774);
nand U22259 (N_22259,N_18156,N_17113);
nor U22260 (N_22260,N_18710,N_15397);
or U22261 (N_22261,N_17304,N_15503);
or U22262 (N_22262,N_16333,N_18040);
nand U22263 (N_22263,N_15550,N_19030);
nand U22264 (N_22264,N_15342,N_19736);
nand U22265 (N_22265,N_17048,N_16964);
nand U22266 (N_22266,N_18576,N_16140);
nand U22267 (N_22267,N_16529,N_15790);
and U22268 (N_22268,N_17495,N_18154);
nand U22269 (N_22269,N_19073,N_16717);
nand U22270 (N_22270,N_19508,N_17313);
nand U22271 (N_22271,N_17308,N_19544);
nor U22272 (N_22272,N_15979,N_19531);
or U22273 (N_22273,N_16413,N_19410);
nor U22274 (N_22274,N_19102,N_17390);
nand U22275 (N_22275,N_19589,N_19668);
and U22276 (N_22276,N_15691,N_16682);
nand U22277 (N_22277,N_19709,N_19564);
and U22278 (N_22278,N_16502,N_18968);
nor U22279 (N_22279,N_15431,N_17383);
or U22280 (N_22280,N_16084,N_18302);
and U22281 (N_22281,N_16863,N_18995);
xor U22282 (N_22282,N_18190,N_16462);
or U22283 (N_22283,N_18113,N_19035);
or U22284 (N_22284,N_15062,N_16928);
and U22285 (N_22285,N_15734,N_17219);
nor U22286 (N_22286,N_18164,N_15084);
nor U22287 (N_22287,N_15252,N_15396);
or U22288 (N_22288,N_15695,N_18568);
nor U22289 (N_22289,N_15217,N_18076);
xnor U22290 (N_22290,N_17303,N_18050);
or U22291 (N_22291,N_17072,N_19302);
or U22292 (N_22292,N_18673,N_15666);
or U22293 (N_22293,N_19603,N_18476);
nor U22294 (N_22294,N_16793,N_19348);
nor U22295 (N_22295,N_19640,N_18819);
or U22296 (N_22296,N_17400,N_16894);
nand U22297 (N_22297,N_17918,N_15483);
nor U22298 (N_22298,N_17036,N_16370);
and U22299 (N_22299,N_18049,N_19809);
xnor U22300 (N_22300,N_19698,N_17866);
nand U22301 (N_22301,N_17353,N_18415);
or U22302 (N_22302,N_16705,N_16152);
nor U22303 (N_22303,N_17734,N_15292);
nand U22304 (N_22304,N_17763,N_18681);
xor U22305 (N_22305,N_19477,N_18348);
or U22306 (N_22306,N_17577,N_16223);
nand U22307 (N_22307,N_19482,N_18841);
and U22308 (N_22308,N_15758,N_16599);
or U22309 (N_22309,N_15035,N_15009);
xnor U22310 (N_22310,N_19676,N_16021);
or U22311 (N_22311,N_19019,N_16322);
or U22312 (N_22312,N_16805,N_19016);
nor U22313 (N_22313,N_15935,N_19296);
or U22314 (N_22314,N_19633,N_19915);
xor U22315 (N_22315,N_19343,N_17807);
and U22316 (N_22316,N_16025,N_19755);
or U22317 (N_22317,N_18088,N_19113);
nand U22318 (N_22318,N_19620,N_18941);
and U22319 (N_22319,N_16915,N_16539);
xnor U22320 (N_22320,N_18528,N_15104);
and U22321 (N_22321,N_16269,N_17735);
or U22322 (N_22322,N_19778,N_19613);
or U22323 (N_22323,N_19922,N_18984);
nand U22324 (N_22324,N_19763,N_15864);
and U22325 (N_22325,N_17345,N_18488);
nor U22326 (N_22326,N_18510,N_16155);
nand U22327 (N_22327,N_15279,N_19181);
and U22328 (N_22328,N_16378,N_16759);
nor U22329 (N_22329,N_19118,N_18238);
nand U22330 (N_22330,N_15594,N_15162);
and U22331 (N_22331,N_17055,N_17284);
nor U22332 (N_22332,N_16575,N_15185);
nor U22333 (N_22333,N_17940,N_15160);
and U22334 (N_22334,N_18060,N_16867);
or U22335 (N_22335,N_16170,N_18901);
nand U22336 (N_22336,N_18293,N_17845);
nand U22337 (N_22337,N_17524,N_18045);
nand U22338 (N_22338,N_15328,N_16623);
and U22339 (N_22339,N_16197,N_15373);
and U22340 (N_22340,N_15783,N_17401);
or U22341 (N_22341,N_15609,N_16184);
and U22342 (N_22342,N_19562,N_16817);
and U22343 (N_22343,N_17328,N_19105);
nand U22344 (N_22344,N_17023,N_15744);
and U22345 (N_22345,N_15847,N_17660);
nand U22346 (N_22346,N_19672,N_18266);
or U22347 (N_22347,N_16572,N_15588);
and U22348 (N_22348,N_15916,N_17411);
nor U22349 (N_22349,N_15890,N_17860);
and U22350 (N_22350,N_18399,N_17415);
nand U22351 (N_22351,N_16646,N_16078);
nor U22352 (N_22352,N_19612,N_16367);
nand U22353 (N_22353,N_19587,N_19499);
or U22354 (N_22354,N_15867,N_18384);
and U22355 (N_22355,N_15955,N_18196);
nand U22356 (N_22356,N_17196,N_19788);
nand U22357 (N_22357,N_19435,N_15046);
and U22358 (N_22358,N_17005,N_18940);
nor U22359 (N_22359,N_16796,N_15794);
nand U22360 (N_22360,N_15527,N_16665);
or U22361 (N_22361,N_19363,N_18422);
nand U22362 (N_22362,N_17397,N_17377);
and U22363 (N_22363,N_17675,N_17563);
and U22364 (N_22364,N_17403,N_15485);
and U22365 (N_22365,N_18304,N_18344);
or U22366 (N_22366,N_19243,N_15306);
nand U22367 (N_22367,N_15370,N_15787);
and U22368 (N_22368,N_16427,N_17355);
or U22369 (N_22369,N_15946,N_16952);
nand U22370 (N_22370,N_19386,N_19902);
and U22371 (N_22371,N_17993,N_19605);
or U22372 (N_22372,N_19910,N_19290);
or U22373 (N_22373,N_17255,N_17279);
xnor U22374 (N_22374,N_17507,N_15584);
xor U22375 (N_22375,N_15344,N_17576);
or U22376 (N_22376,N_19898,N_16585);
and U22377 (N_22377,N_17253,N_18728);
nor U22378 (N_22378,N_17022,N_17822);
or U22379 (N_22379,N_16754,N_16916);
xor U22380 (N_22380,N_18211,N_19524);
nand U22381 (N_22381,N_19117,N_15719);
and U22382 (N_22382,N_16716,N_18972);
nand U22383 (N_22383,N_16455,N_18746);
nor U22384 (N_22384,N_18357,N_18479);
nor U22385 (N_22385,N_17064,N_15294);
nand U22386 (N_22386,N_17305,N_15407);
and U22387 (N_22387,N_19332,N_19529);
and U22388 (N_22388,N_18395,N_17819);
nor U22389 (N_22389,N_16495,N_15521);
and U22390 (N_22390,N_15452,N_17471);
nor U22391 (N_22391,N_18692,N_19774);
nand U22392 (N_22392,N_18199,N_16240);
and U22393 (N_22393,N_15545,N_17920);
or U22394 (N_22394,N_17003,N_15526);
nand U22395 (N_22395,N_19741,N_18495);
or U22396 (N_22396,N_19033,N_18635);
nand U22397 (N_22397,N_15846,N_15873);
or U22398 (N_22398,N_18379,N_15493);
nor U22399 (N_22399,N_17178,N_15296);
xor U22400 (N_22400,N_19570,N_16673);
or U22401 (N_22401,N_16485,N_18493);
and U22402 (N_22402,N_15298,N_18220);
nor U22403 (N_22403,N_16234,N_16622);
and U22404 (N_22404,N_15723,N_19459);
and U22405 (N_22405,N_15591,N_17138);
and U22406 (N_22406,N_19220,N_16973);
nand U22407 (N_22407,N_16960,N_17031);
nor U22408 (N_22408,N_16929,N_17343);
nor U22409 (N_22409,N_19950,N_19169);
nor U22410 (N_22410,N_19859,N_15011);
xor U22411 (N_22411,N_19853,N_18273);
and U22412 (N_22412,N_19816,N_15957);
nand U22413 (N_22413,N_17877,N_18181);
or U22414 (N_22414,N_16918,N_18806);
nand U22415 (N_22415,N_18194,N_16007);
or U22416 (N_22416,N_15950,N_15428);
and U22417 (N_22417,N_17833,N_17097);
or U22418 (N_22418,N_18846,N_16961);
nor U22419 (N_22419,N_16886,N_19401);
and U22420 (N_22420,N_19604,N_15351);
nand U22421 (N_22421,N_16011,N_18489);
or U22422 (N_22422,N_15242,N_17961);
nand U22423 (N_22423,N_17909,N_18013);
nor U22424 (N_22424,N_19214,N_16336);
nor U22425 (N_22425,N_17249,N_15041);
and U22426 (N_22426,N_18541,N_18662);
nor U22427 (N_22427,N_15769,N_18280);
nand U22428 (N_22428,N_15412,N_18153);
xor U22429 (N_22429,N_18748,N_18463);
or U22430 (N_22430,N_18734,N_18478);
or U22431 (N_22431,N_19607,N_18139);
nand U22432 (N_22432,N_15711,N_16438);
or U22433 (N_22433,N_18971,N_19195);
nand U22434 (N_22434,N_18921,N_17847);
nand U22435 (N_22435,N_18759,N_19536);
nand U22436 (N_22436,N_18922,N_15238);
or U22437 (N_22437,N_16288,N_17444);
or U22438 (N_22438,N_19124,N_17140);
nor U22439 (N_22439,N_16865,N_18243);
xnor U22440 (N_22440,N_17879,N_18022);
and U22441 (N_22441,N_15222,N_16729);
and U22442 (N_22442,N_17953,N_18697);
and U22443 (N_22443,N_15224,N_15567);
xor U22444 (N_22444,N_19866,N_16842);
nor U22445 (N_22445,N_18620,N_16662);
and U22446 (N_22446,N_16936,N_17234);
nor U22447 (N_22447,N_17639,N_17778);
nor U22448 (N_22448,N_16303,N_18763);
or U22449 (N_22449,N_19509,N_15985);
or U22450 (N_22450,N_19304,N_18248);
xor U22451 (N_22451,N_15276,N_18935);
or U22452 (N_22452,N_18184,N_17614);
or U22453 (N_22453,N_19140,N_16838);
and U22454 (N_22454,N_16308,N_19679);
nor U22455 (N_22455,N_15082,N_16667);
nor U22456 (N_22456,N_15388,N_17260);
or U22457 (N_22457,N_18226,N_19851);
xor U22458 (N_22458,N_16877,N_15392);
or U22459 (N_22459,N_16482,N_19894);
nor U22460 (N_22460,N_17222,N_15299);
nor U22461 (N_22461,N_18432,N_16235);
or U22462 (N_22462,N_18096,N_19377);
or U22463 (N_22463,N_19262,N_18176);
and U22464 (N_22464,N_18056,N_18661);
or U22465 (N_22465,N_16706,N_16327);
and U22466 (N_22466,N_16861,N_16275);
nor U22467 (N_22467,N_15958,N_15685);
nand U22468 (N_22468,N_16628,N_18699);
nand U22469 (N_22469,N_15448,N_16956);
nor U22470 (N_22470,N_16618,N_16612);
nor U22471 (N_22471,N_19400,N_18633);
nor U22472 (N_22472,N_19415,N_17243);
nand U22473 (N_22473,N_16625,N_18954);
or U22474 (N_22474,N_17740,N_19098);
xnor U22475 (N_22475,N_19527,N_17038);
or U22476 (N_22476,N_17424,N_19854);
and U22477 (N_22477,N_18287,N_15040);
nand U22478 (N_22478,N_17273,N_16040);
or U22479 (N_22479,N_19355,N_18508);
nand U22480 (N_22480,N_16369,N_17039);
or U22481 (N_22481,N_16188,N_17976);
nand U22482 (N_22482,N_16374,N_17727);
xnor U22483 (N_22483,N_16666,N_19991);
and U22484 (N_22484,N_16965,N_15643);
and U22485 (N_22485,N_16810,N_16030);
and U22486 (N_22486,N_19542,N_15086);
and U22487 (N_22487,N_19099,N_19429);
nor U22488 (N_22488,N_15288,N_17068);
or U22489 (N_22489,N_15551,N_18094);
and U22490 (N_22490,N_19879,N_18070);
nor U22491 (N_22491,N_15848,N_18502);
or U22492 (N_22492,N_15300,N_17658);
and U22493 (N_22493,N_18414,N_15554);
nor U22494 (N_22494,N_18768,N_18353);
nand U22495 (N_22495,N_19516,N_17947);
nor U22496 (N_22496,N_15346,N_19919);
or U22497 (N_22497,N_19857,N_18093);
nor U22498 (N_22498,N_15669,N_17618);
xnor U22499 (N_22499,N_17160,N_16500);
or U22500 (N_22500,N_18922,N_18792);
nand U22501 (N_22501,N_19262,N_17656);
nor U22502 (N_22502,N_18371,N_15406);
and U22503 (N_22503,N_15536,N_18325);
or U22504 (N_22504,N_19837,N_16720);
and U22505 (N_22505,N_16544,N_18470);
xor U22506 (N_22506,N_19313,N_15351);
nor U22507 (N_22507,N_16982,N_16604);
and U22508 (N_22508,N_17416,N_18778);
nor U22509 (N_22509,N_18891,N_17152);
nor U22510 (N_22510,N_18660,N_16947);
or U22511 (N_22511,N_19838,N_15272);
nand U22512 (N_22512,N_18729,N_15241);
xnor U22513 (N_22513,N_16032,N_18811);
nor U22514 (N_22514,N_17474,N_18023);
nand U22515 (N_22515,N_17609,N_15779);
nand U22516 (N_22516,N_17511,N_16762);
and U22517 (N_22517,N_17970,N_19084);
nand U22518 (N_22518,N_18371,N_19577);
nor U22519 (N_22519,N_15727,N_19378);
nor U22520 (N_22520,N_19702,N_18159);
and U22521 (N_22521,N_15223,N_19761);
or U22522 (N_22522,N_15027,N_18841);
nand U22523 (N_22523,N_16852,N_15659);
and U22524 (N_22524,N_19355,N_15717);
nand U22525 (N_22525,N_19990,N_19445);
nand U22526 (N_22526,N_18473,N_19109);
xnor U22527 (N_22527,N_18426,N_17636);
nand U22528 (N_22528,N_18355,N_15522);
or U22529 (N_22529,N_15565,N_17270);
and U22530 (N_22530,N_18145,N_18761);
or U22531 (N_22531,N_15343,N_19488);
or U22532 (N_22532,N_19915,N_15981);
nand U22533 (N_22533,N_16937,N_19760);
nor U22534 (N_22534,N_19226,N_17025);
or U22535 (N_22535,N_18896,N_16646);
or U22536 (N_22536,N_15067,N_16112);
nor U22537 (N_22537,N_17380,N_17951);
nor U22538 (N_22538,N_18027,N_18126);
and U22539 (N_22539,N_15666,N_15172);
nand U22540 (N_22540,N_15914,N_17705);
or U22541 (N_22541,N_15838,N_16541);
nor U22542 (N_22542,N_16967,N_16810);
nor U22543 (N_22543,N_16834,N_19363);
nand U22544 (N_22544,N_19141,N_15893);
nand U22545 (N_22545,N_15508,N_19508);
or U22546 (N_22546,N_19407,N_18494);
nand U22547 (N_22547,N_15219,N_16580);
nor U22548 (N_22548,N_17710,N_17519);
and U22549 (N_22549,N_18232,N_19591);
and U22550 (N_22550,N_19111,N_19987);
or U22551 (N_22551,N_17111,N_15464);
xor U22552 (N_22552,N_19645,N_17150);
nand U22553 (N_22553,N_19387,N_15125);
and U22554 (N_22554,N_16696,N_15185);
nor U22555 (N_22555,N_16284,N_19206);
and U22556 (N_22556,N_15609,N_19641);
nor U22557 (N_22557,N_17417,N_19471);
nor U22558 (N_22558,N_19402,N_19793);
and U22559 (N_22559,N_19228,N_15607);
or U22560 (N_22560,N_17661,N_16274);
nand U22561 (N_22561,N_18324,N_18105);
nand U22562 (N_22562,N_18258,N_19581);
nand U22563 (N_22563,N_18008,N_16312);
and U22564 (N_22564,N_16225,N_16668);
xnor U22565 (N_22565,N_19837,N_15974);
or U22566 (N_22566,N_18548,N_17731);
and U22567 (N_22567,N_19083,N_16368);
and U22568 (N_22568,N_15401,N_16499);
or U22569 (N_22569,N_19709,N_17403);
and U22570 (N_22570,N_17725,N_15407);
xor U22571 (N_22571,N_19502,N_17754);
nand U22572 (N_22572,N_16709,N_19282);
or U22573 (N_22573,N_15864,N_18069);
nor U22574 (N_22574,N_15422,N_19159);
or U22575 (N_22575,N_17310,N_18141);
nand U22576 (N_22576,N_17360,N_15660);
xor U22577 (N_22577,N_19743,N_16975);
and U22578 (N_22578,N_17080,N_15160);
nor U22579 (N_22579,N_16802,N_16117);
and U22580 (N_22580,N_17682,N_15590);
and U22581 (N_22581,N_16045,N_18992);
nand U22582 (N_22582,N_17126,N_17976);
nor U22583 (N_22583,N_19851,N_19446);
or U22584 (N_22584,N_17391,N_17229);
or U22585 (N_22585,N_18173,N_16156);
or U22586 (N_22586,N_17366,N_18965);
nand U22587 (N_22587,N_19258,N_19808);
nand U22588 (N_22588,N_18967,N_15734);
nand U22589 (N_22589,N_15525,N_15716);
or U22590 (N_22590,N_16221,N_17651);
or U22591 (N_22591,N_15888,N_15266);
or U22592 (N_22592,N_18025,N_16121);
nor U22593 (N_22593,N_19719,N_18946);
and U22594 (N_22594,N_16743,N_18120);
nor U22595 (N_22595,N_18684,N_19735);
and U22596 (N_22596,N_15550,N_19106);
or U22597 (N_22597,N_18202,N_18162);
nand U22598 (N_22598,N_16509,N_17960);
or U22599 (N_22599,N_16894,N_15101);
nand U22600 (N_22600,N_15126,N_19037);
or U22601 (N_22601,N_18450,N_19450);
nor U22602 (N_22602,N_19545,N_18486);
nand U22603 (N_22603,N_16080,N_17018);
nor U22604 (N_22604,N_16215,N_18126);
or U22605 (N_22605,N_15784,N_16150);
xnor U22606 (N_22606,N_17465,N_17827);
and U22607 (N_22607,N_18833,N_17158);
nand U22608 (N_22608,N_15648,N_15970);
and U22609 (N_22609,N_16865,N_16796);
and U22610 (N_22610,N_19752,N_16392);
nand U22611 (N_22611,N_15609,N_18945);
nor U22612 (N_22612,N_17613,N_16223);
xnor U22613 (N_22613,N_16185,N_17527);
nor U22614 (N_22614,N_15349,N_19445);
xor U22615 (N_22615,N_17416,N_17675);
nand U22616 (N_22616,N_16140,N_15125);
nand U22617 (N_22617,N_19854,N_17320);
nor U22618 (N_22618,N_17338,N_15175);
xnor U22619 (N_22619,N_16732,N_18999);
xnor U22620 (N_22620,N_16952,N_19133);
nor U22621 (N_22621,N_19213,N_16428);
nor U22622 (N_22622,N_18138,N_19550);
nor U22623 (N_22623,N_16424,N_17661);
and U22624 (N_22624,N_17910,N_19673);
nand U22625 (N_22625,N_19643,N_18188);
nor U22626 (N_22626,N_19171,N_15299);
nand U22627 (N_22627,N_19231,N_16379);
nor U22628 (N_22628,N_19575,N_15096);
xor U22629 (N_22629,N_15829,N_19100);
and U22630 (N_22630,N_18026,N_18869);
nand U22631 (N_22631,N_19107,N_19366);
and U22632 (N_22632,N_17934,N_15387);
and U22633 (N_22633,N_18119,N_19539);
nor U22634 (N_22634,N_16066,N_16345);
nand U22635 (N_22635,N_19020,N_15444);
or U22636 (N_22636,N_15568,N_17770);
and U22637 (N_22637,N_17770,N_19023);
nor U22638 (N_22638,N_18835,N_17712);
nand U22639 (N_22639,N_17448,N_17867);
nor U22640 (N_22640,N_19795,N_15774);
nand U22641 (N_22641,N_15659,N_18572);
or U22642 (N_22642,N_16130,N_17069);
nor U22643 (N_22643,N_16250,N_16227);
nand U22644 (N_22644,N_16027,N_15140);
nor U22645 (N_22645,N_15653,N_17016);
nand U22646 (N_22646,N_17189,N_18704);
nor U22647 (N_22647,N_19225,N_15113);
or U22648 (N_22648,N_19772,N_16320);
nor U22649 (N_22649,N_18016,N_16413);
nor U22650 (N_22650,N_17926,N_16714);
or U22651 (N_22651,N_16199,N_17010);
or U22652 (N_22652,N_19063,N_18984);
and U22653 (N_22653,N_19944,N_19889);
and U22654 (N_22654,N_19879,N_18477);
and U22655 (N_22655,N_18899,N_16463);
and U22656 (N_22656,N_18859,N_16567);
and U22657 (N_22657,N_18324,N_18556);
xor U22658 (N_22658,N_15669,N_19866);
or U22659 (N_22659,N_18281,N_19964);
nand U22660 (N_22660,N_15240,N_17180);
or U22661 (N_22661,N_19017,N_15997);
or U22662 (N_22662,N_19256,N_19791);
or U22663 (N_22663,N_18224,N_16611);
and U22664 (N_22664,N_18443,N_19487);
nand U22665 (N_22665,N_19206,N_17814);
or U22666 (N_22666,N_19362,N_16313);
nor U22667 (N_22667,N_16650,N_19473);
or U22668 (N_22668,N_18047,N_19782);
and U22669 (N_22669,N_15924,N_16607);
and U22670 (N_22670,N_18325,N_18656);
or U22671 (N_22671,N_15021,N_15529);
nor U22672 (N_22672,N_17926,N_19885);
nor U22673 (N_22673,N_17250,N_18316);
nand U22674 (N_22674,N_18819,N_15533);
nand U22675 (N_22675,N_19477,N_16882);
nand U22676 (N_22676,N_15281,N_17973);
and U22677 (N_22677,N_17577,N_17160);
nor U22678 (N_22678,N_19591,N_18662);
or U22679 (N_22679,N_18353,N_18002);
nor U22680 (N_22680,N_15704,N_16898);
and U22681 (N_22681,N_19159,N_17466);
nor U22682 (N_22682,N_16435,N_18874);
or U22683 (N_22683,N_18015,N_18136);
nand U22684 (N_22684,N_18515,N_16083);
nor U22685 (N_22685,N_15488,N_18290);
nor U22686 (N_22686,N_17651,N_17752);
and U22687 (N_22687,N_17939,N_18841);
nor U22688 (N_22688,N_15206,N_17467);
nor U22689 (N_22689,N_17683,N_17055);
nand U22690 (N_22690,N_15779,N_16983);
nand U22691 (N_22691,N_17989,N_16389);
or U22692 (N_22692,N_15855,N_17427);
nor U22693 (N_22693,N_16503,N_17308);
or U22694 (N_22694,N_19445,N_15820);
or U22695 (N_22695,N_19789,N_19029);
nor U22696 (N_22696,N_18922,N_19977);
nor U22697 (N_22697,N_17954,N_19199);
and U22698 (N_22698,N_19973,N_17754);
nand U22699 (N_22699,N_16146,N_15729);
and U22700 (N_22700,N_17896,N_16023);
and U22701 (N_22701,N_15228,N_15878);
and U22702 (N_22702,N_15752,N_18685);
and U22703 (N_22703,N_18017,N_17814);
or U22704 (N_22704,N_19260,N_17878);
or U22705 (N_22705,N_19426,N_15812);
nor U22706 (N_22706,N_17145,N_18386);
nor U22707 (N_22707,N_19571,N_19543);
xor U22708 (N_22708,N_16097,N_16782);
nor U22709 (N_22709,N_19974,N_19519);
and U22710 (N_22710,N_17981,N_17747);
nor U22711 (N_22711,N_15503,N_18904);
xnor U22712 (N_22712,N_15731,N_15910);
and U22713 (N_22713,N_17193,N_18030);
nand U22714 (N_22714,N_17243,N_16330);
or U22715 (N_22715,N_15403,N_17647);
and U22716 (N_22716,N_16431,N_19835);
nor U22717 (N_22717,N_18516,N_18228);
nand U22718 (N_22718,N_19540,N_17910);
or U22719 (N_22719,N_16294,N_17099);
xor U22720 (N_22720,N_18200,N_16711);
nor U22721 (N_22721,N_17184,N_18246);
nand U22722 (N_22722,N_19082,N_16259);
or U22723 (N_22723,N_18561,N_15630);
xnor U22724 (N_22724,N_18991,N_19113);
or U22725 (N_22725,N_16732,N_18351);
nor U22726 (N_22726,N_16257,N_19763);
nand U22727 (N_22727,N_15919,N_19653);
and U22728 (N_22728,N_17581,N_15303);
nand U22729 (N_22729,N_16068,N_18481);
or U22730 (N_22730,N_15339,N_16651);
nand U22731 (N_22731,N_19783,N_18885);
or U22732 (N_22732,N_17073,N_17967);
or U22733 (N_22733,N_16673,N_17278);
and U22734 (N_22734,N_18213,N_19523);
and U22735 (N_22735,N_16147,N_16014);
and U22736 (N_22736,N_16084,N_15896);
xnor U22737 (N_22737,N_15737,N_17692);
or U22738 (N_22738,N_19819,N_18451);
and U22739 (N_22739,N_16662,N_15104);
nor U22740 (N_22740,N_16634,N_19074);
or U22741 (N_22741,N_18211,N_15100);
or U22742 (N_22742,N_19844,N_19999);
and U22743 (N_22743,N_17023,N_16931);
or U22744 (N_22744,N_18072,N_17245);
nand U22745 (N_22745,N_16712,N_16318);
xor U22746 (N_22746,N_18550,N_19079);
nor U22747 (N_22747,N_15179,N_17262);
and U22748 (N_22748,N_18366,N_15985);
or U22749 (N_22749,N_17063,N_15997);
nor U22750 (N_22750,N_15643,N_19044);
nor U22751 (N_22751,N_16501,N_17114);
nor U22752 (N_22752,N_19243,N_19866);
nor U22753 (N_22753,N_19814,N_17401);
or U22754 (N_22754,N_18622,N_17339);
and U22755 (N_22755,N_19300,N_15192);
nand U22756 (N_22756,N_17335,N_19529);
nor U22757 (N_22757,N_15266,N_15853);
nand U22758 (N_22758,N_17028,N_19207);
nor U22759 (N_22759,N_17220,N_18407);
nor U22760 (N_22760,N_16256,N_16541);
xor U22761 (N_22761,N_19626,N_16798);
and U22762 (N_22762,N_18898,N_19740);
and U22763 (N_22763,N_15684,N_16599);
nor U22764 (N_22764,N_19943,N_16037);
and U22765 (N_22765,N_16935,N_16195);
and U22766 (N_22766,N_15573,N_15479);
and U22767 (N_22767,N_18064,N_16767);
and U22768 (N_22768,N_15063,N_16621);
xor U22769 (N_22769,N_16738,N_15032);
nor U22770 (N_22770,N_18884,N_17610);
and U22771 (N_22771,N_15074,N_17563);
nor U22772 (N_22772,N_15977,N_17981);
nor U22773 (N_22773,N_19634,N_19702);
nand U22774 (N_22774,N_16016,N_17791);
xnor U22775 (N_22775,N_17619,N_16710);
xnor U22776 (N_22776,N_15476,N_16631);
or U22777 (N_22777,N_18032,N_19639);
and U22778 (N_22778,N_15873,N_17188);
or U22779 (N_22779,N_18725,N_15532);
nor U22780 (N_22780,N_19327,N_15192);
nor U22781 (N_22781,N_18142,N_19142);
nor U22782 (N_22782,N_17884,N_17461);
and U22783 (N_22783,N_18251,N_16481);
nor U22784 (N_22784,N_19465,N_19597);
or U22785 (N_22785,N_17210,N_15294);
nor U22786 (N_22786,N_19374,N_15626);
and U22787 (N_22787,N_16076,N_18772);
nand U22788 (N_22788,N_15682,N_16656);
and U22789 (N_22789,N_17644,N_17601);
and U22790 (N_22790,N_17813,N_16819);
nor U22791 (N_22791,N_15541,N_18425);
nand U22792 (N_22792,N_18453,N_19004);
nor U22793 (N_22793,N_18045,N_16647);
nand U22794 (N_22794,N_15053,N_15630);
nand U22795 (N_22795,N_18906,N_18504);
nor U22796 (N_22796,N_16582,N_17737);
nor U22797 (N_22797,N_16519,N_16196);
nor U22798 (N_22798,N_16284,N_18550);
nor U22799 (N_22799,N_15681,N_18944);
or U22800 (N_22800,N_18786,N_18123);
and U22801 (N_22801,N_19584,N_16548);
nand U22802 (N_22802,N_17711,N_19767);
or U22803 (N_22803,N_17118,N_19405);
nor U22804 (N_22804,N_16661,N_15976);
nor U22805 (N_22805,N_19619,N_19894);
xnor U22806 (N_22806,N_19982,N_18459);
and U22807 (N_22807,N_18385,N_18932);
and U22808 (N_22808,N_16976,N_15971);
and U22809 (N_22809,N_18538,N_17446);
nor U22810 (N_22810,N_16832,N_15225);
nor U22811 (N_22811,N_19824,N_17713);
nand U22812 (N_22812,N_19093,N_16642);
nand U22813 (N_22813,N_15073,N_17294);
or U22814 (N_22814,N_16338,N_18709);
nor U22815 (N_22815,N_19801,N_15465);
nand U22816 (N_22816,N_16983,N_19935);
and U22817 (N_22817,N_15056,N_19011);
and U22818 (N_22818,N_17360,N_16313);
or U22819 (N_22819,N_15664,N_17516);
xor U22820 (N_22820,N_17788,N_16156);
xor U22821 (N_22821,N_15949,N_15529);
or U22822 (N_22822,N_19610,N_17194);
and U22823 (N_22823,N_16672,N_17807);
nand U22824 (N_22824,N_16066,N_19692);
and U22825 (N_22825,N_15708,N_19931);
and U22826 (N_22826,N_18377,N_17052);
nand U22827 (N_22827,N_15754,N_15601);
nand U22828 (N_22828,N_16765,N_19621);
and U22829 (N_22829,N_19794,N_18267);
or U22830 (N_22830,N_17853,N_15678);
or U22831 (N_22831,N_18263,N_15488);
nor U22832 (N_22832,N_16145,N_15199);
nor U22833 (N_22833,N_19878,N_18221);
nor U22834 (N_22834,N_17797,N_17761);
nand U22835 (N_22835,N_15354,N_17293);
nor U22836 (N_22836,N_19889,N_18901);
nor U22837 (N_22837,N_16076,N_18427);
or U22838 (N_22838,N_17236,N_19336);
nor U22839 (N_22839,N_16724,N_17835);
xnor U22840 (N_22840,N_16562,N_15856);
or U22841 (N_22841,N_17885,N_16611);
xnor U22842 (N_22842,N_19283,N_19731);
nand U22843 (N_22843,N_15195,N_19670);
xor U22844 (N_22844,N_17178,N_15276);
xor U22845 (N_22845,N_19372,N_17771);
nor U22846 (N_22846,N_18411,N_15360);
and U22847 (N_22847,N_16939,N_18961);
nor U22848 (N_22848,N_15816,N_16079);
or U22849 (N_22849,N_19417,N_18434);
and U22850 (N_22850,N_18494,N_19324);
and U22851 (N_22851,N_15910,N_17729);
and U22852 (N_22852,N_16403,N_16895);
and U22853 (N_22853,N_18702,N_18920);
xnor U22854 (N_22854,N_19115,N_15070);
nor U22855 (N_22855,N_17076,N_16795);
xor U22856 (N_22856,N_19858,N_15404);
nand U22857 (N_22857,N_19975,N_16519);
nor U22858 (N_22858,N_16250,N_19526);
xor U22859 (N_22859,N_15238,N_19061);
nor U22860 (N_22860,N_16521,N_15667);
or U22861 (N_22861,N_15103,N_15241);
or U22862 (N_22862,N_15405,N_18523);
nor U22863 (N_22863,N_15992,N_17571);
or U22864 (N_22864,N_18999,N_19731);
and U22865 (N_22865,N_18103,N_16986);
nor U22866 (N_22866,N_16509,N_17861);
or U22867 (N_22867,N_16562,N_18354);
or U22868 (N_22868,N_17642,N_17491);
and U22869 (N_22869,N_17137,N_18193);
nand U22870 (N_22870,N_15837,N_16913);
nor U22871 (N_22871,N_17874,N_18590);
nor U22872 (N_22872,N_19443,N_17317);
nor U22873 (N_22873,N_18402,N_16146);
nand U22874 (N_22874,N_16027,N_15862);
and U22875 (N_22875,N_17561,N_18475);
and U22876 (N_22876,N_16046,N_18882);
xor U22877 (N_22877,N_17563,N_18607);
xnor U22878 (N_22878,N_18287,N_17417);
nand U22879 (N_22879,N_17120,N_15644);
or U22880 (N_22880,N_15636,N_18663);
nor U22881 (N_22881,N_18996,N_17843);
or U22882 (N_22882,N_19518,N_15467);
nand U22883 (N_22883,N_18959,N_15105);
and U22884 (N_22884,N_15449,N_16181);
or U22885 (N_22885,N_19434,N_15112);
xor U22886 (N_22886,N_17927,N_17731);
nor U22887 (N_22887,N_16247,N_15791);
or U22888 (N_22888,N_15833,N_16336);
or U22889 (N_22889,N_19193,N_15509);
nor U22890 (N_22890,N_18105,N_16692);
or U22891 (N_22891,N_18130,N_19969);
nor U22892 (N_22892,N_18631,N_18756);
nand U22893 (N_22893,N_18798,N_18372);
and U22894 (N_22894,N_16024,N_16226);
and U22895 (N_22895,N_18902,N_16460);
or U22896 (N_22896,N_17060,N_18160);
and U22897 (N_22897,N_19520,N_17819);
xnor U22898 (N_22898,N_16401,N_18691);
nor U22899 (N_22899,N_16818,N_15921);
and U22900 (N_22900,N_16579,N_18512);
nand U22901 (N_22901,N_15608,N_19403);
nor U22902 (N_22902,N_17305,N_19666);
nor U22903 (N_22903,N_16031,N_15676);
nand U22904 (N_22904,N_17952,N_15419);
nor U22905 (N_22905,N_19119,N_19890);
or U22906 (N_22906,N_17048,N_18046);
or U22907 (N_22907,N_16087,N_18521);
nor U22908 (N_22908,N_17298,N_15418);
and U22909 (N_22909,N_17509,N_17212);
nand U22910 (N_22910,N_17143,N_17944);
nor U22911 (N_22911,N_17529,N_19292);
nand U22912 (N_22912,N_15492,N_15485);
nor U22913 (N_22913,N_18034,N_17057);
and U22914 (N_22914,N_15429,N_17785);
xor U22915 (N_22915,N_17477,N_16025);
or U22916 (N_22916,N_17384,N_18126);
nor U22917 (N_22917,N_16504,N_17107);
xor U22918 (N_22918,N_18286,N_18251);
or U22919 (N_22919,N_19438,N_15358);
nand U22920 (N_22920,N_19832,N_19979);
or U22921 (N_22921,N_18904,N_18862);
and U22922 (N_22922,N_16543,N_16742);
nor U22923 (N_22923,N_16167,N_15900);
nor U22924 (N_22924,N_19728,N_15079);
and U22925 (N_22925,N_17365,N_16499);
or U22926 (N_22926,N_18939,N_15715);
nand U22927 (N_22927,N_17441,N_19966);
nand U22928 (N_22928,N_17703,N_17964);
nor U22929 (N_22929,N_16515,N_19704);
nand U22930 (N_22930,N_18893,N_19926);
nand U22931 (N_22931,N_19896,N_15092);
nor U22932 (N_22932,N_17572,N_15940);
nor U22933 (N_22933,N_17806,N_16805);
and U22934 (N_22934,N_16683,N_15618);
nand U22935 (N_22935,N_19335,N_16351);
nor U22936 (N_22936,N_19304,N_16041);
xor U22937 (N_22937,N_18999,N_15232);
or U22938 (N_22938,N_15110,N_15543);
xnor U22939 (N_22939,N_15195,N_19834);
and U22940 (N_22940,N_18164,N_17114);
nor U22941 (N_22941,N_19583,N_15486);
xnor U22942 (N_22942,N_18511,N_17497);
nand U22943 (N_22943,N_18155,N_19258);
or U22944 (N_22944,N_17996,N_15104);
nor U22945 (N_22945,N_18445,N_17261);
or U22946 (N_22946,N_16173,N_17672);
and U22947 (N_22947,N_17066,N_16103);
nor U22948 (N_22948,N_16700,N_17743);
nand U22949 (N_22949,N_19453,N_19697);
nand U22950 (N_22950,N_19682,N_19232);
nor U22951 (N_22951,N_19123,N_19427);
and U22952 (N_22952,N_16335,N_17359);
xnor U22953 (N_22953,N_19100,N_19516);
nor U22954 (N_22954,N_17211,N_19446);
nand U22955 (N_22955,N_19002,N_15294);
nand U22956 (N_22956,N_18369,N_17084);
or U22957 (N_22957,N_18842,N_19439);
nand U22958 (N_22958,N_16272,N_16472);
nand U22959 (N_22959,N_16509,N_19620);
and U22960 (N_22960,N_17703,N_17305);
xor U22961 (N_22961,N_15162,N_17487);
nand U22962 (N_22962,N_19736,N_15417);
or U22963 (N_22963,N_16785,N_17052);
and U22964 (N_22964,N_16937,N_16533);
and U22965 (N_22965,N_18019,N_19462);
or U22966 (N_22966,N_18111,N_17924);
nor U22967 (N_22967,N_18991,N_19745);
or U22968 (N_22968,N_18764,N_15844);
nand U22969 (N_22969,N_16580,N_17093);
nand U22970 (N_22970,N_17335,N_18911);
nor U22971 (N_22971,N_17225,N_19635);
or U22972 (N_22972,N_18476,N_15603);
nor U22973 (N_22973,N_16896,N_15404);
or U22974 (N_22974,N_19270,N_18192);
and U22975 (N_22975,N_18867,N_19205);
and U22976 (N_22976,N_19275,N_19848);
or U22977 (N_22977,N_15967,N_16705);
nand U22978 (N_22978,N_19217,N_16745);
and U22979 (N_22979,N_15415,N_17817);
or U22980 (N_22980,N_18694,N_16346);
nand U22981 (N_22981,N_16534,N_15102);
nor U22982 (N_22982,N_16012,N_17834);
xnor U22983 (N_22983,N_15390,N_18519);
nand U22984 (N_22984,N_19417,N_17958);
nor U22985 (N_22985,N_17564,N_15251);
nand U22986 (N_22986,N_15141,N_16557);
xor U22987 (N_22987,N_18929,N_16070);
and U22988 (N_22988,N_17277,N_18390);
and U22989 (N_22989,N_17853,N_15917);
nor U22990 (N_22990,N_19212,N_19005);
and U22991 (N_22991,N_19778,N_18900);
nand U22992 (N_22992,N_17055,N_18654);
and U22993 (N_22993,N_19064,N_15682);
or U22994 (N_22994,N_16737,N_18550);
nor U22995 (N_22995,N_17903,N_15565);
or U22996 (N_22996,N_16718,N_18206);
nand U22997 (N_22997,N_16486,N_15235);
or U22998 (N_22998,N_17737,N_18752);
or U22999 (N_22999,N_16843,N_18452);
xnor U23000 (N_23000,N_19685,N_16758);
nor U23001 (N_23001,N_18407,N_18567);
and U23002 (N_23002,N_19164,N_17316);
and U23003 (N_23003,N_18378,N_18256);
nand U23004 (N_23004,N_19670,N_16041);
and U23005 (N_23005,N_19902,N_15008);
nand U23006 (N_23006,N_18140,N_19488);
and U23007 (N_23007,N_15299,N_18885);
and U23008 (N_23008,N_19385,N_17106);
and U23009 (N_23009,N_17493,N_18895);
nand U23010 (N_23010,N_19752,N_17816);
nor U23011 (N_23011,N_19161,N_18475);
or U23012 (N_23012,N_16112,N_15905);
nor U23013 (N_23013,N_18796,N_19730);
or U23014 (N_23014,N_15490,N_18719);
xnor U23015 (N_23015,N_17580,N_16956);
nor U23016 (N_23016,N_18003,N_17916);
or U23017 (N_23017,N_15741,N_18682);
nand U23018 (N_23018,N_17768,N_19496);
and U23019 (N_23019,N_19749,N_17489);
or U23020 (N_23020,N_16370,N_19653);
and U23021 (N_23021,N_17212,N_17583);
nor U23022 (N_23022,N_17753,N_18953);
and U23023 (N_23023,N_17399,N_17347);
and U23024 (N_23024,N_15741,N_18379);
and U23025 (N_23025,N_18330,N_18454);
nand U23026 (N_23026,N_18158,N_19378);
nand U23027 (N_23027,N_17508,N_18361);
and U23028 (N_23028,N_16025,N_16688);
and U23029 (N_23029,N_17285,N_17199);
and U23030 (N_23030,N_19530,N_19029);
nor U23031 (N_23031,N_15549,N_17624);
nor U23032 (N_23032,N_17866,N_19858);
nand U23033 (N_23033,N_15136,N_18148);
nor U23034 (N_23034,N_17307,N_16629);
xnor U23035 (N_23035,N_19231,N_18108);
nand U23036 (N_23036,N_16914,N_18060);
or U23037 (N_23037,N_17669,N_17501);
or U23038 (N_23038,N_18342,N_18083);
nand U23039 (N_23039,N_19052,N_15172);
nor U23040 (N_23040,N_19950,N_17799);
or U23041 (N_23041,N_19557,N_16571);
or U23042 (N_23042,N_15592,N_19091);
nor U23043 (N_23043,N_16211,N_16239);
nor U23044 (N_23044,N_19862,N_18783);
and U23045 (N_23045,N_17832,N_17617);
nor U23046 (N_23046,N_15476,N_19561);
nand U23047 (N_23047,N_16484,N_16127);
nor U23048 (N_23048,N_17494,N_16153);
or U23049 (N_23049,N_17190,N_15784);
and U23050 (N_23050,N_16086,N_16905);
nand U23051 (N_23051,N_18604,N_15320);
or U23052 (N_23052,N_18836,N_17358);
xor U23053 (N_23053,N_18257,N_19833);
nand U23054 (N_23054,N_16361,N_15685);
nor U23055 (N_23055,N_17416,N_17190);
or U23056 (N_23056,N_17345,N_16517);
and U23057 (N_23057,N_16678,N_18353);
or U23058 (N_23058,N_17254,N_18639);
nor U23059 (N_23059,N_19132,N_18568);
nand U23060 (N_23060,N_15318,N_15691);
nand U23061 (N_23061,N_19341,N_16030);
and U23062 (N_23062,N_16859,N_19822);
nand U23063 (N_23063,N_16739,N_17658);
and U23064 (N_23064,N_18226,N_16376);
nor U23065 (N_23065,N_18084,N_18069);
or U23066 (N_23066,N_16990,N_19933);
nand U23067 (N_23067,N_19757,N_19872);
nand U23068 (N_23068,N_17965,N_15693);
and U23069 (N_23069,N_17701,N_16493);
nor U23070 (N_23070,N_15168,N_17585);
xnor U23071 (N_23071,N_19224,N_15203);
nand U23072 (N_23072,N_19276,N_15294);
and U23073 (N_23073,N_17308,N_15379);
and U23074 (N_23074,N_16983,N_15469);
nand U23075 (N_23075,N_15839,N_17693);
or U23076 (N_23076,N_18284,N_18692);
and U23077 (N_23077,N_15300,N_15321);
nor U23078 (N_23078,N_17705,N_19211);
nand U23079 (N_23079,N_16224,N_18510);
xor U23080 (N_23080,N_15441,N_18724);
and U23081 (N_23081,N_19919,N_19995);
nor U23082 (N_23082,N_19602,N_17453);
nand U23083 (N_23083,N_19982,N_17144);
and U23084 (N_23084,N_19699,N_16925);
nor U23085 (N_23085,N_15525,N_16701);
and U23086 (N_23086,N_18753,N_17934);
nor U23087 (N_23087,N_15193,N_19849);
or U23088 (N_23088,N_16938,N_18862);
or U23089 (N_23089,N_17598,N_17037);
nor U23090 (N_23090,N_16964,N_17865);
nand U23091 (N_23091,N_18420,N_15162);
or U23092 (N_23092,N_15591,N_16736);
or U23093 (N_23093,N_18195,N_17046);
or U23094 (N_23094,N_17450,N_15274);
nand U23095 (N_23095,N_19046,N_18476);
nor U23096 (N_23096,N_19881,N_17356);
nand U23097 (N_23097,N_15970,N_17756);
nand U23098 (N_23098,N_15086,N_19544);
or U23099 (N_23099,N_18211,N_16375);
nor U23100 (N_23100,N_17471,N_17021);
or U23101 (N_23101,N_17132,N_17358);
nor U23102 (N_23102,N_15809,N_15225);
nor U23103 (N_23103,N_19346,N_17372);
nand U23104 (N_23104,N_17539,N_18840);
or U23105 (N_23105,N_19159,N_18284);
or U23106 (N_23106,N_19947,N_16308);
nor U23107 (N_23107,N_17933,N_17799);
or U23108 (N_23108,N_19012,N_16749);
nor U23109 (N_23109,N_17491,N_18146);
nor U23110 (N_23110,N_15724,N_19702);
xnor U23111 (N_23111,N_16906,N_15976);
or U23112 (N_23112,N_17396,N_19798);
or U23113 (N_23113,N_18670,N_18069);
nand U23114 (N_23114,N_17087,N_15481);
xnor U23115 (N_23115,N_17766,N_15099);
nand U23116 (N_23116,N_19114,N_16846);
or U23117 (N_23117,N_19574,N_17622);
or U23118 (N_23118,N_19169,N_16316);
xor U23119 (N_23119,N_16228,N_15374);
nand U23120 (N_23120,N_19058,N_19255);
nand U23121 (N_23121,N_19130,N_18324);
or U23122 (N_23122,N_19250,N_18002);
nor U23123 (N_23123,N_16613,N_19125);
and U23124 (N_23124,N_18600,N_18828);
nor U23125 (N_23125,N_18882,N_16816);
and U23126 (N_23126,N_18822,N_15132);
nor U23127 (N_23127,N_16167,N_16923);
nor U23128 (N_23128,N_19623,N_17728);
nor U23129 (N_23129,N_17891,N_17596);
nand U23130 (N_23130,N_19548,N_19589);
nand U23131 (N_23131,N_19893,N_15863);
or U23132 (N_23132,N_19778,N_15026);
or U23133 (N_23133,N_18157,N_17722);
or U23134 (N_23134,N_16222,N_19613);
nand U23135 (N_23135,N_17184,N_15153);
or U23136 (N_23136,N_18762,N_18568);
and U23137 (N_23137,N_19053,N_18351);
nand U23138 (N_23138,N_17684,N_16653);
and U23139 (N_23139,N_17148,N_16814);
nor U23140 (N_23140,N_17009,N_17359);
xor U23141 (N_23141,N_17030,N_16513);
and U23142 (N_23142,N_18720,N_15908);
nand U23143 (N_23143,N_19387,N_19190);
nand U23144 (N_23144,N_18059,N_19081);
nand U23145 (N_23145,N_19611,N_18690);
nand U23146 (N_23146,N_18371,N_19433);
nand U23147 (N_23147,N_18314,N_16358);
nand U23148 (N_23148,N_17105,N_18855);
nor U23149 (N_23149,N_16837,N_19605);
or U23150 (N_23150,N_15613,N_16037);
xor U23151 (N_23151,N_18146,N_17952);
xnor U23152 (N_23152,N_16226,N_18991);
or U23153 (N_23153,N_17419,N_17528);
and U23154 (N_23154,N_16208,N_18242);
and U23155 (N_23155,N_15194,N_19019);
nor U23156 (N_23156,N_15465,N_16458);
nand U23157 (N_23157,N_18353,N_16745);
or U23158 (N_23158,N_17061,N_18638);
nor U23159 (N_23159,N_18809,N_19958);
and U23160 (N_23160,N_18241,N_15883);
or U23161 (N_23161,N_16767,N_18747);
or U23162 (N_23162,N_15109,N_18229);
and U23163 (N_23163,N_17661,N_17360);
nand U23164 (N_23164,N_15637,N_17465);
and U23165 (N_23165,N_15369,N_16013);
and U23166 (N_23166,N_19747,N_19796);
or U23167 (N_23167,N_19438,N_19897);
or U23168 (N_23168,N_18844,N_18170);
nor U23169 (N_23169,N_18799,N_17817);
or U23170 (N_23170,N_17054,N_18451);
or U23171 (N_23171,N_17923,N_18032);
or U23172 (N_23172,N_15322,N_19750);
nor U23173 (N_23173,N_16389,N_19631);
or U23174 (N_23174,N_17447,N_17743);
and U23175 (N_23175,N_17393,N_16960);
or U23176 (N_23176,N_17205,N_15818);
nor U23177 (N_23177,N_19273,N_16969);
nor U23178 (N_23178,N_19771,N_17003);
or U23179 (N_23179,N_18744,N_15602);
and U23180 (N_23180,N_18923,N_19405);
nor U23181 (N_23181,N_19625,N_19419);
nand U23182 (N_23182,N_18771,N_17484);
and U23183 (N_23183,N_16620,N_17629);
or U23184 (N_23184,N_19157,N_19564);
and U23185 (N_23185,N_18658,N_18089);
nand U23186 (N_23186,N_17100,N_19404);
nand U23187 (N_23187,N_18739,N_18953);
nand U23188 (N_23188,N_16081,N_19500);
and U23189 (N_23189,N_15110,N_19148);
nor U23190 (N_23190,N_16672,N_15427);
or U23191 (N_23191,N_15179,N_16694);
nand U23192 (N_23192,N_16020,N_17350);
and U23193 (N_23193,N_19043,N_18267);
or U23194 (N_23194,N_17769,N_16678);
nand U23195 (N_23195,N_18650,N_17965);
nand U23196 (N_23196,N_19673,N_17247);
xnor U23197 (N_23197,N_18980,N_18057);
and U23198 (N_23198,N_15212,N_15119);
nand U23199 (N_23199,N_18962,N_16231);
and U23200 (N_23200,N_15525,N_17049);
and U23201 (N_23201,N_19963,N_15847);
nor U23202 (N_23202,N_16692,N_18898);
nand U23203 (N_23203,N_15613,N_17903);
or U23204 (N_23204,N_18133,N_17368);
xor U23205 (N_23205,N_17761,N_17624);
nand U23206 (N_23206,N_16373,N_19846);
nor U23207 (N_23207,N_19307,N_18590);
xnor U23208 (N_23208,N_15270,N_19226);
nand U23209 (N_23209,N_18016,N_19252);
and U23210 (N_23210,N_15609,N_16942);
or U23211 (N_23211,N_19893,N_17162);
and U23212 (N_23212,N_19822,N_18903);
or U23213 (N_23213,N_15597,N_15194);
nand U23214 (N_23214,N_19574,N_19141);
nand U23215 (N_23215,N_18731,N_17932);
and U23216 (N_23216,N_18978,N_16528);
nor U23217 (N_23217,N_18628,N_19551);
xnor U23218 (N_23218,N_15582,N_15315);
nand U23219 (N_23219,N_15026,N_17905);
nand U23220 (N_23220,N_16022,N_16389);
and U23221 (N_23221,N_18308,N_19035);
or U23222 (N_23222,N_18703,N_18701);
nor U23223 (N_23223,N_18773,N_19447);
nand U23224 (N_23224,N_19407,N_19512);
xnor U23225 (N_23225,N_15693,N_17989);
and U23226 (N_23226,N_16123,N_17930);
or U23227 (N_23227,N_18419,N_19301);
or U23228 (N_23228,N_19972,N_17643);
and U23229 (N_23229,N_18144,N_18870);
nand U23230 (N_23230,N_15765,N_19614);
nor U23231 (N_23231,N_19967,N_18157);
nand U23232 (N_23232,N_17117,N_15746);
or U23233 (N_23233,N_16448,N_19861);
and U23234 (N_23234,N_19579,N_18453);
and U23235 (N_23235,N_16906,N_17080);
nand U23236 (N_23236,N_17974,N_18624);
and U23237 (N_23237,N_16967,N_17697);
or U23238 (N_23238,N_16357,N_15463);
nor U23239 (N_23239,N_19629,N_19399);
or U23240 (N_23240,N_15172,N_17078);
or U23241 (N_23241,N_19632,N_19168);
or U23242 (N_23242,N_19431,N_19978);
nor U23243 (N_23243,N_19928,N_17077);
nand U23244 (N_23244,N_15963,N_15954);
xor U23245 (N_23245,N_19825,N_19943);
nand U23246 (N_23246,N_16248,N_17576);
and U23247 (N_23247,N_15690,N_16516);
nand U23248 (N_23248,N_16746,N_15666);
and U23249 (N_23249,N_17639,N_18917);
and U23250 (N_23250,N_16004,N_17739);
and U23251 (N_23251,N_17119,N_15232);
nand U23252 (N_23252,N_15428,N_19317);
nor U23253 (N_23253,N_16656,N_18034);
xnor U23254 (N_23254,N_15172,N_17401);
and U23255 (N_23255,N_18663,N_15774);
nor U23256 (N_23256,N_15273,N_15467);
or U23257 (N_23257,N_15923,N_15255);
or U23258 (N_23258,N_18752,N_19873);
nor U23259 (N_23259,N_16529,N_17327);
nor U23260 (N_23260,N_16289,N_19508);
xnor U23261 (N_23261,N_18674,N_15617);
and U23262 (N_23262,N_15018,N_15957);
or U23263 (N_23263,N_15593,N_15898);
xor U23264 (N_23264,N_16589,N_17514);
nor U23265 (N_23265,N_17565,N_15766);
nor U23266 (N_23266,N_17657,N_17554);
or U23267 (N_23267,N_17180,N_15025);
nor U23268 (N_23268,N_19178,N_18727);
and U23269 (N_23269,N_15327,N_19733);
nor U23270 (N_23270,N_18413,N_17052);
and U23271 (N_23271,N_16784,N_15915);
or U23272 (N_23272,N_19731,N_16086);
nor U23273 (N_23273,N_15469,N_19244);
nand U23274 (N_23274,N_19414,N_15217);
nor U23275 (N_23275,N_17578,N_19778);
and U23276 (N_23276,N_18153,N_15024);
or U23277 (N_23277,N_18298,N_17202);
and U23278 (N_23278,N_17780,N_17839);
or U23279 (N_23279,N_18156,N_17110);
nor U23280 (N_23280,N_17113,N_15397);
nand U23281 (N_23281,N_18361,N_15851);
xnor U23282 (N_23282,N_15035,N_16308);
or U23283 (N_23283,N_16738,N_15592);
nor U23284 (N_23284,N_17668,N_16313);
xor U23285 (N_23285,N_16831,N_17734);
or U23286 (N_23286,N_19227,N_15460);
and U23287 (N_23287,N_15456,N_17548);
nor U23288 (N_23288,N_17246,N_18617);
nand U23289 (N_23289,N_18622,N_16046);
and U23290 (N_23290,N_15232,N_18323);
xnor U23291 (N_23291,N_16666,N_15346);
or U23292 (N_23292,N_19910,N_16091);
nor U23293 (N_23293,N_16840,N_16343);
nand U23294 (N_23294,N_19426,N_17671);
and U23295 (N_23295,N_19578,N_18331);
nand U23296 (N_23296,N_18439,N_15416);
or U23297 (N_23297,N_17533,N_18308);
nand U23298 (N_23298,N_15073,N_19703);
nor U23299 (N_23299,N_18108,N_18332);
nand U23300 (N_23300,N_18456,N_17035);
xnor U23301 (N_23301,N_17635,N_18611);
nand U23302 (N_23302,N_18891,N_16216);
nor U23303 (N_23303,N_18007,N_15470);
nor U23304 (N_23304,N_16429,N_19109);
xnor U23305 (N_23305,N_18524,N_17728);
nand U23306 (N_23306,N_16647,N_16431);
nor U23307 (N_23307,N_17916,N_19305);
and U23308 (N_23308,N_17681,N_17026);
and U23309 (N_23309,N_18219,N_18370);
xnor U23310 (N_23310,N_17075,N_19622);
nand U23311 (N_23311,N_18559,N_15253);
nor U23312 (N_23312,N_15764,N_16161);
and U23313 (N_23313,N_15572,N_18525);
nand U23314 (N_23314,N_15880,N_18400);
or U23315 (N_23315,N_18678,N_18229);
nand U23316 (N_23316,N_17010,N_16018);
and U23317 (N_23317,N_17704,N_19152);
nand U23318 (N_23318,N_17995,N_19941);
or U23319 (N_23319,N_18295,N_19488);
nand U23320 (N_23320,N_17254,N_18429);
nor U23321 (N_23321,N_15631,N_17110);
or U23322 (N_23322,N_16181,N_17459);
and U23323 (N_23323,N_17925,N_16433);
and U23324 (N_23324,N_19847,N_18942);
nor U23325 (N_23325,N_17451,N_18734);
and U23326 (N_23326,N_17248,N_19638);
nand U23327 (N_23327,N_15682,N_17891);
nor U23328 (N_23328,N_17874,N_17601);
and U23329 (N_23329,N_16766,N_18071);
nor U23330 (N_23330,N_17277,N_17544);
nor U23331 (N_23331,N_18836,N_16820);
nor U23332 (N_23332,N_17400,N_15049);
nor U23333 (N_23333,N_18068,N_17422);
nor U23334 (N_23334,N_17279,N_15335);
nor U23335 (N_23335,N_17949,N_16719);
and U23336 (N_23336,N_15959,N_15691);
nor U23337 (N_23337,N_19414,N_15533);
and U23338 (N_23338,N_16405,N_19389);
and U23339 (N_23339,N_17318,N_15841);
or U23340 (N_23340,N_18897,N_17488);
nor U23341 (N_23341,N_19350,N_19701);
or U23342 (N_23342,N_19614,N_19252);
or U23343 (N_23343,N_15198,N_17487);
or U23344 (N_23344,N_15152,N_17142);
or U23345 (N_23345,N_16699,N_17728);
and U23346 (N_23346,N_16468,N_18637);
nand U23347 (N_23347,N_19843,N_15352);
and U23348 (N_23348,N_19788,N_17863);
and U23349 (N_23349,N_16026,N_19513);
nor U23350 (N_23350,N_15041,N_18756);
or U23351 (N_23351,N_18807,N_17754);
nand U23352 (N_23352,N_17001,N_18095);
xnor U23353 (N_23353,N_18659,N_19815);
and U23354 (N_23354,N_16649,N_19297);
xnor U23355 (N_23355,N_15581,N_19064);
nor U23356 (N_23356,N_17032,N_17938);
nor U23357 (N_23357,N_18190,N_16870);
nor U23358 (N_23358,N_16670,N_17115);
nand U23359 (N_23359,N_19767,N_15572);
xor U23360 (N_23360,N_16184,N_15854);
nand U23361 (N_23361,N_15107,N_17842);
and U23362 (N_23362,N_17456,N_16171);
nand U23363 (N_23363,N_16055,N_15173);
nor U23364 (N_23364,N_16980,N_18799);
nor U23365 (N_23365,N_17298,N_17313);
or U23366 (N_23366,N_17085,N_18036);
and U23367 (N_23367,N_15013,N_17643);
and U23368 (N_23368,N_15482,N_16029);
or U23369 (N_23369,N_15998,N_18978);
nand U23370 (N_23370,N_16925,N_18386);
xor U23371 (N_23371,N_16406,N_19847);
nand U23372 (N_23372,N_19771,N_17510);
nor U23373 (N_23373,N_18517,N_15066);
or U23374 (N_23374,N_18856,N_16415);
nor U23375 (N_23375,N_15585,N_19160);
or U23376 (N_23376,N_16215,N_17329);
xor U23377 (N_23377,N_17356,N_18028);
nor U23378 (N_23378,N_15061,N_19180);
nand U23379 (N_23379,N_17752,N_19154);
nor U23380 (N_23380,N_16046,N_15124);
and U23381 (N_23381,N_19578,N_17235);
nor U23382 (N_23382,N_17871,N_19632);
nand U23383 (N_23383,N_19604,N_19982);
or U23384 (N_23384,N_16272,N_18726);
and U23385 (N_23385,N_18376,N_18215);
nand U23386 (N_23386,N_18424,N_18479);
or U23387 (N_23387,N_18034,N_18194);
nand U23388 (N_23388,N_15987,N_17348);
and U23389 (N_23389,N_16239,N_17936);
nand U23390 (N_23390,N_18883,N_15575);
nand U23391 (N_23391,N_17478,N_15509);
nor U23392 (N_23392,N_16705,N_19712);
nand U23393 (N_23393,N_17278,N_15776);
or U23394 (N_23394,N_17945,N_15827);
and U23395 (N_23395,N_18175,N_15621);
nor U23396 (N_23396,N_15642,N_19891);
and U23397 (N_23397,N_18884,N_15520);
and U23398 (N_23398,N_16441,N_19316);
nand U23399 (N_23399,N_16539,N_15717);
and U23400 (N_23400,N_16093,N_19538);
nor U23401 (N_23401,N_19427,N_18152);
nand U23402 (N_23402,N_18066,N_16213);
nor U23403 (N_23403,N_17018,N_16883);
nand U23404 (N_23404,N_15220,N_18269);
xor U23405 (N_23405,N_17442,N_19201);
nor U23406 (N_23406,N_18261,N_19232);
nor U23407 (N_23407,N_18074,N_15006);
nor U23408 (N_23408,N_18092,N_18619);
nor U23409 (N_23409,N_19535,N_18847);
or U23410 (N_23410,N_15258,N_18765);
and U23411 (N_23411,N_16453,N_16145);
and U23412 (N_23412,N_18191,N_15091);
or U23413 (N_23413,N_19637,N_18171);
and U23414 (N_23414,N_17642,N_17121);
nor U23415 (N_23415,N_17033,N_16722);
nor U23416 (N_23416,N_17622,N_17731);
xnor U23417 (N_23417,N_19931,N_17011);
or U23418 (N_23418,N_15859,N_19393);
or U23419 (N_23419,N_17892,N_19575);
nand U23420 (N_23420,N_16266,N_19583);
and U23421 (N_23421,N_15030,N_19597);
nor U23422 (N_23422,N_18393,N_15395);
xnor U23423 (N_23423,N_15548,N_18702);
nand U23424 (N_23424,N_19882,N_16465);
or U23425 (N_23425,N_18463,N_16215);
nor U23426 (N_23426,N_19739,N_18551);
nand U23427 (N_23427,N_15155,N_15945);
nor U23428 (N_23428,N_19947,N_16625);
nor U23429 (N_23429,N_19467,N_18686);
nand U23430 (N_23430,N_17588,N_16401);
nand U23431 (N_23431,N_15260,N_16668);
nor U23432 (N_23432,N_17054,N_15349);
nor U23433 (N_23433,N_16887,N_16737);
nor U23434 (N_23434,N_15134,N_17783);
or U23435 (N_23435,N_18342,N_15627);
nor U23436 (N_23436,N_18068,N_18838);
nor U23437 (N_23437,N_19244,N_17748);
xor U23438 (N_23438,N_19142,N_16014);
nand U23439 (N_23439,N_15120,N_19926);
nand U23440 (N_23440,N_19583,N_15383);
or U23441 (N_23441,N_17993,N_16491);
or U23442 (N_23442,N_17733,N_17634);
and U23443 (N_23443,N_16524,N_16509);
or U23444 (N_23444,N_17305,N_18924);
and U23445 (N_23445,N_18390,N_18009);
nor U23446 (N_23446,N_17137,N_19880);
or U23447 (N_23447,N_17741,N_19596);
or U23448 (N_23448,N_19607,N_16953);
and U23449 (N_23449,N_16042,N_15344);
nor U23450 (N_23450,N_19965,N_17014);
and U23451 (N_23451,N_17242,N_18127);
or U23452 (N_23452,N_19767,N_15839);
xor U23453 (N_23453,N_18823,N_19331);
and U23454 (N_23454,N_17851,N_16145);
nor U23455 (N_23455,N_19917,N_18352);
nor U23456 (N_23456,N_18848,N_15339);
nand U23457 (N_23457,N_15544,N_19523);
or U23458 (N_23458,N_19806,N_15311);
nor U23459 (N_23459,N_18516,N_18572);
or U23460 (N_23460,N_18890,N_19840);
nand U23461 (N_23461,N_16747,N_16847);
nor U23462 (N_23462,N_15009,N_19328);
and U23463 (N_23463,N_15869,N_18596);
or U23464 (N_23464,N_19326,N_18578);
or U23465 (N_23465,N_18564,N_16895);
nor U23466 (N_23466,N_15545,N_19900);
nor U23467 (N_23467,N_19699,N_18113);
and U23468 (N_23468,N_17911,N_15612);
nor U23469 (N_23469,N_19083,N_19746);
nor U23470 (N_23470,N_18268,N_15854);
xnor U23471 (N_23471,N_15688,N_17065);
nor U23472 (N_23472,N_19844,N_15368);
and U23473 (N_23473,N_18306,N_19336);
or U23474 (N_23474,N_18123,N_17830);
nor U23475 (N_23475,N_15832,N_18452);
nor U23476 (N_23476,N_18647,N_18419);
nor U23477 (N_23477,N_15695,N_16736);
nand U23478 (N_23478,N_18918,N_16020);
and U23479 (N_23479,N_16948,N_18507);
and U23480 (N_23480,N_18103,N_17736);
xor U23481 (N_23481,N_19108,N_18536);
and U23482 (N_23482,N_15126,N_19929);
xor U23483 (N_23483,N_16623,N_16512);
nor U23484 (N_23484,N_15977,N_17844);
nand U23485 (N_23485,N_16999,N_17161);
nand U23486 (N_23486,N_15445,N_15260);
xor U23487 (N_23487,N_16676,N_19922);
nor U23488 (N_23488,N_18161,N_15403);
nand U23489 (N_23489,N_17467,N_19268);
or U23490 (N_23490,N_15143,N_16408);
nand U23491 (N_23491,N_18619,N_19074);
and U23492 (N_23492,N_16215,N_18471);
nand U23493 (N_23493,N_15045,N_18277);
or U23494 (N_23494,N_15102,N_19023);
nor U23495 (N_23495,N_15328,N_17544);
xor U23496 (N_23496,N_15350,N_16347);
nand U23497 (N_23497,N_17596,N_15316);
nand U23498 (N_23498,N_19211,N_19361);
and U23499 (N_23499,N_15389,N_19134);
nor U23500 (N_23500,N_17652,N_19791);
and U23501 (N_23501,N_16531,N_16880);
or U23502 (N_23502,N_17755,N_16237);
and U23503 (N_23503,N_17943,N_18287);
nor U23504 (N_23504,N_17323,N_18446);
nand U23505 (N_23505,N_19838,N_19835);
or U23506 (N_23506,N_17734,N_16315);
or U23507 (N_23507,N_17189,N_18404);
or U23508 (N_23508,N_15759,N_15768);
or U23509 (N_23509,N_18290,N_17017);
or U23510 (N_23510,N_15690,N_15296);
nand U23511 (N_23511,N_19300,N_17713);
nand U23512 (N_23512,N_18816,N_17141);
xor U23513 (N_23513,N_19519,N_18173);
xnor U23514 (N_23514,N_18853,N_18528);
nand U23515 (N_23515,N_19804,N_16517);
and U23516 (N_23516,N_15541,N_15380);
nand U23517 (N_23517,N_15631,N_18493);
nand U23518 (N_23518,N_16002,N_17468);
or U23519 (N_23519,N_16380,N_19441);
or U23520 (N_23520,N_16764,N_17100);
nand U23521 (N_23521,N_19101,N_16072);
nand U23522 (N_23522,N_15756,N_19681);
nor U23523 (N_23523,N_18094,N_19469);
nor U23524 (N_23524,N_16132,N_15281);
xnor U23525 (N_23525,N_18553,N_19023);
or U23526 (N_23526,N_19505,N_15669);
nor U23527 (N_23527,N_16577,N_16062);
and U23528 (N_23528,N_19134,N_18241);
and U23529 (N_23529,N_19769,N_16487);
or U23530 (N_23530,N_18419,N_17779);
and U23531 (N_23531,N_19092,N_18645);
nand U23532 (N_23532,N_16421,N_17922);
or U23533 (N_23533,N_19498,N_19584);
nor U23534 (N_23534,N_18996,N_16148);
and U23535 (N_23535,N_18147,N_16484);
xor U23536 (N_23536,N_15323,N_17645);
nor U23537 (N_23537,N_17984,N_17456);
nand U23538 (N_23538,N_16219,N_16020);
or U23539 (N_23539,N_15813,N_19377);
nor U23540 (N_23540,N_16324,N_15986);
nor U23541 (N_23541,N_19775,N_16978);
nor U23542 (N_23542,N_16895,N_19802);
nand U23543 (N_23543,N_16492,N_15591);
nand U23544 (N_23544,N_16738,N_15113);
and U23545 (N_23545,N_16637,N_19406);
nor U23546 (N_23546,N_17853,N_17333);
xnor U23547 (N_23547,N_17691,N_15594);
nor U23548 (N_23548,N_15031,N_16840);
and U23549 (N_23549,N_18332,N_19661);
and U23550 (N_23550,N_18958,N_19298);
xor U23551 (N_23551,N_19984,N_15566);
nor U23552 (N_23552,N_15564,N_15856);
or U23553 (N_23553,N_19999,N_15217);
nand U23554 (N_23554,N_19431,N_18541);
nand U23555 (N_23555,N_18541,N_17301);
or U23556 (N_23556,N_17786,N_18507);
nand U23557 (N_23557,N_19212,N_16167);
and U23558 (N_23558,N_17194,N_19445);
nand U23559 (N_23559,N_17431,N_16981);
nor U23560 (N_23560,N_17921,N_18776);
nor U23561 (N_23561,N_15727,N_18701);
nand U23562 (N_23562,N_19274,N_18890);
and U23563 (N_23563,N_16873,N_17822);
nor U23564 (N_23564,N_17468,N_17249);
nor U23565 (N_23565,N_18164,N_19219);
xnor U23566 (N_23566,N_16810,N_18458);
or U23567 (N_23567,N_15926,N_17685);
nand U23568 (N_23568,N_16012,N_17724);
nor U23569 (N_23569,N_16566,N_19519);
nor U23570 (N_23570,N_16446,N_16521);
nor U23571 (N_23571,N_16877,N_19157);
xor U23572 (N_23572,N_17319,N_17562);
nor U23573 (N_23573,N_19695,N_19798);
nand U23574 (N_23574,N_17273,N_16112);
and U23575 (N_23575,N_18236,N_19804);
nor U23576 (N_23576,N_16395,N_16477);
or U23577 (N_23577,N_19579,N_17956);
and U23578 (N_23578,N_15344,N_19402);
and U23579 (N_23579,N_19429,N_18148);
or U23580 (N_23580,N_19865,N_15938);
or U23581 (N_23581,N_16429,N_15626);
and U23582 (N_23582,N_16642,N_15881);
or U23583 (N_23583,N_19827,N_18894);
nor U23584 (N_23584,N_15614,N_17667);
nand U23585 (N_23585,N_16608,N_15977);
xor U23586 (N_23586,N_18072,N_18672);
xor U23587 (N_23587,N_15594,N_16732);
or U23588 (N_23588,N_18371,N_15369);
nand U23589 (N_23589,N_19249,N_17166);
and U23590 (N_23590,N_18819,N_17798);
xor U23591 (N_23591,N_15115,N_16963);
or U23592 (N_23592,N_18224,N_17900);
nand U23593 (N_23593,N_19916,N_16916);
and U23594 (N_23594,N_18798,N_17034);
or U23595 (N_23595,N_15467,N_18086);
nand U23596 (N_23596,N_18553,N_15485);
and U23597 (N_23597,N_17382,N_19633);
or U23598 (N_23598,N_19804,N_19628);
nor U23599 (N_23599,N_17304,N_18121);
or U23600 (N_23600,N_19716,N_19175);
nand U23601 (N_23601,N_17980,N_19073);
and U23602 (N_23602,N_15439,N_19630);
xnor U23603 (N_23603,N_18244,N_15725);
nor U23604 (N_23604,N_18044,N_17759);
xor U23605 (N_23605,N_16544,N_17770);
and U23606 (N_23606,N_17074,N_15882);
nor U23607 (N_23607,N_19928,N_18885);
nand U23608 (N_23608,N_19538,N_18660);
or U23609 (N_23609,N_15872,N_16155);
or U23610 (N_23610,N_19467,N_15457);
or U23611 (N_23611,N_18184,N_19321);
nor U23612 (N_23612,N_15084,N_18232);
nor U23613 (N_23613,N_16058,N_16524);
xor U23614 (N_23614,N_15091,N_17291);
and U23615 (N_23615,N_17386,N_16871);
and U23616 (N_23616,N_17387,N_15221);
nor U23617 (N_23617,N_18370,N_19859);
nor U23618 (N_23618,N_16145,N_16775);
or U23619 (N_23619,N_19165,N_18152);
nor U23620 (N_23620,N_15381,N_17662);
and U23621 (N_23621,N_16862,N_18131);
nand U23622 (N_23622,N_15893,N_17882);
and U23623 (N_23623,N_18007,N_19214);
nand U23624 (N_23624,N_17294,N_15921);
nor U23625 (N_23625,N_15877,N_15236);
xnor U23626 (N_23626,N_19899,N_16474);
nand U23627 (N_23627,N_18802,N_17480);
nor U23628 (N_23628,N_17230,N_15037);
xnor U23629 (N_23629,N_17582,N_17123);
nand U23630 (N_23630,N_18119,N_17455);
or U23631 (N_23631,N_16830,N_19892);
nor U23632 (N_23632,N_17010,N_19153);
nand U23633 (N_23633,N_19890,N_19381);
nand U23634 (N_23634,N_15626,N_16642);
nand U23635 (N_23635,N_19161,N_16704);
nand U23636 (N_23636,N_19338,N_15651);
nor U23637 (N_23637,N_16341,N_18411);
nor U23638 (N_23638,N_16423,N_17005);
and U23639 (N_23639,N_19248,N_19316);
and U23640 (N_23640,N_17101,N_15134);
nand U23641 (N_23641,N_18901,N_17881);
nor U23642 (N_23642,N_15921,N_19403);
and U23643 (N_23643,N_19173,N_19919);
nor U23644 (N_23644,N_17773,N_17182);
and U23645 (N_23645,N_19904,N_16906);
and U23646 (N_23646,N_18390,N_18950);
and U23647 (N_23647,N_17898,N_18955);
nor U23648 (N_23648,N_17639,N_19784);
nand U23649 (N_23649,N_16794,N_19046);
and U23650 (N_23650,N_15509,N_16970);
nor U23651 (N_23651,N_17244,N_19295);
nand U23652 (N_23652,N_19879,N_16551);
or U23653 (N_23653,N_15406,N_19535);
and U23654 (N_23654,N_15645,N_19222);
or U23655 (N_23655,N_17689,N_16513);
and U23656 (N_23656,N_16901,N_17405);
xor U23657 (N_23657,N_18280,N_15226);
and U23658 (N_23658,N_17855,N_18287);
and U23659 (N_23659,N_17137,N_15533);
nand U23660 (N_23660,N_18055,N_16742);
and U23661 (N_23661,N_16600,N_15952);
nand U23662 (N_23662,N_18114,N_19011);
nor U23663 (N_23663,N_16723,N_16571);
nor U23664 (N_23664,N_17515,N_17079);
nand U23665 (N_23665,N_15141,N_17745);
or U23666 (N_23666,N_18688,N_18026);
or U23667 (N_23667,N_15915,N_19801);
or U23668 (N_23668,N_19512,N_16901);
or U23669 (N_23669,N_17852,N_15842);
and U23670 (N_23670,N_16772,N_16863);
or U23671 (N_23671,N_19021,N_18041);
nand U23672 (N_23672,N_19175,N_16062);
xor U23673 (N_23673,N_15965,N_15530);
nand U23674 (N_23674,N_15534,N_15951);
or U23675 (N_23675,N_16318,N_15678);
or U23676 (N_23676,N_17971,N_15811);
or U23677 (N_23677,N_16201,N_17222);
and U23678 (N_23678,N_15225,N_16488);
and U23679 (N_23679,N_16307,N_18091);
xor U23680 (N_23680,N_16867,N_16489);
and U23681 (N_23681,N_15892,N_18605);
nor U23682 (N_23682,N_17271,N_17233);
nand U23683 (N_23683,N_17163,N_16948);
xor U23684 (N_23684,N_16247,N_17978);
nand U23685 (N_23685,N_15833,N_15157);
or U23686 (N_23686,N_17247,N_19342);
nand U23687 (N_23687,N_15631,N_18623);
nor U23688 (N_23688,N_19578,N_19778);
or U23689 (N_23689,N_17490,N_19138);
and U23690 (N_23690,N_16887,N_19775);
nand U23691 (N_23691,N_19176,N_18846);
and U23692 (N_23692,N_17740,N_15618);
and U23693 (N_23693,N_19466,N_17725);
and U23694 (N_23694,N_16269,N_17068);
or U23695 (N_23695,N_18566,N_19876);
and U23696 (N_23696,N_17942,N_17757);
or U23697 (N_23697,N_17666,N_16677);
nor U23698 (N_23698,N_17055,N_19946);
and U23699 (N_23699,N_18985,N_16946);
or U23700 (N_23700,N_19973,N_16959);
nand U23701 (N_23701,N_18748,N_18263);
nor U23702 (N_23702,N_18506,N_17517);
nor U23703 (N_23703,N_15131,N_19873);
xor U23704 (N_23704,N_16062,N_17338);
or U23705 (N_23705,N_15753,N_16096);
nand U23706 (N_23706,N_16897,N_16668);
xnor U23707 (N_23707,N_18425,N_15642);
or U23708 (N_23708,N_15853,N_18616);
nor U23709 (N_23709,N_19136,N_19464);
and U23710 (N_23710,N_16658,N_16979);
nand U23711 (N_23711,N_19609,N_17755);
or U23712 (N_23712,N_16246,N_16365);
or U23713 (N_23713,N_19158,N_19723);
nor U23714 (N_23714,N_16223,N_17640);
xor U23715 (N_23715,N_18642,N_18585);
nor U23716 (N_23716,N_18454,N_19035);
or U23717 (N_23717,N_15984,N_16105);
or U23718 (N_23718,N_15198,N_15681);
and U23719 (N_23719,N_16147,N_19916);
nand U23720 (N_23720,N_15997,N_18289);
and U23721 (N_23721,N_15694,N_16864);
nor U23722 (N_23722,N_19902,N_15380);
or U23723 (N_23723,N_17709,N_17251);
or U23724 (N_23724,N_15864,N_18241);
nor U23725 (N_23725,N_18836,N_16633);
nor U23726 (N_23726,N_15539,N_17156);
and U23727 (N_23727,N_19329,N_17971);
or U23728 (N_23728,N_18558,N_17478);
nor U23729 (N_23729,N_15565,N_15439);
nor U23730 (N_23730,N_17488,N_19364);
xor U23731 (N_23731,N_17396,N_15077);
and U23732 (N_23732,N_15635,N_18884);
or U23733 (N_23733,N_19897,N_18948);
xor U23734 (N_23734,N_17501,N_15309);
nand U23735 (N_23735,N_15975,N_16836);
and U23736 (N_23736,N_19280,N_19157);
or U23737 (N_23737,N_16240,N_15933);
and U23738 (N_23738,N_19103,N_18595);
nor U23739 (N_23739,N_18688,N_17734);
nor U23740 (N_23740,N_17015,N_19553);
or U23741 (N_23741,N_19228,N_19221);
or U23742 (N_23742,N_19466,N_15228);
and U23743 (N_23743,N_19456,N_15404);
xnor U23744 (N_23744,N_18722,N_16106);
xnor U23745 (N_23745,N_17752,N_19709);
and U23746 (N_23746,N_18184,N_18487);
and U23747 (N_23747,N_18368,N_19936);
nor U23748 (N_23748,N_15051,N_16442);
nor U23749 (N_23749,N_18243,N_16385);
nor U23750 (N_23750,N_19378,N_18506);
and U23751 (N_23751,N_17035,N_15581);
xnor U23752 (N_23752,N_16262,N_15087);
nand U23753 (N_23753,N_17489,N_18712);
nor U23754 (N_23754,N_16912,N_16611);
and U23755 (N_23755,N_19807,N_16909);
nand U23756 (N_23756,N_18812,N_19884);
nand U23757 (N_23757,N_15103,N_18215);
and U23758 (N_23758,N_16180,N_16334);
xnor U23759 (N_23759,N_15503,N_18531);
xnor U23760 (N_23760,N_16801,N_15552);
or U23761 (N_23761,N_18030,N_18362);
or U23762 (N_23762,N_17440,N_17888);
nand U23763 (N_23763,N_19591,N_18599);
and U23764 (N_23764,N_18879,N_15748);
nor U23765 (N_23765,N_16499,N_19480);
nor U23766 (N_23766,N_16685,N_17090);
xnor U23767 (N_23767,N_19833,N_17457);
nor U23768 (N_23768,N_19999,N_15904);
and U23769 (N_23769,N_17785,N_16675);
nand U23770 (N_23770,N_16286,N_18781);
or U23771 (N_23771,N_17441,N_18480);
nand U23772 (N_23772,N_16090,N_18725);
nand U23773 (N_23773,N_17859,N_19408);
and U23774 (N_23774,N_17500,N_19994);
xnor U23775 (N_23775,N_18192,N_17980);
nand U23776 (N_23776,N_18485,N_16526);
or U23777 (N_23777,N_15417,N_15819);
nand U23778 (N_23778,N_17897,N_18650);
and U23779 (N_23779,N_19851,N_15619);
nand U23780 (N_23780,N_18337,N_19317);
and U23781 (N_23781,N_18668,N_18911);
or U23782 (N_23782,N_19512,N_15802);
and U23783 (N_23783,N_18422,N_18089);
nand U23784 (N_23784,N_16677,N_17905);
and U23785 (N_23785,N_15617,N_19677);
nor U23786 (N_23786,N_18698,N_17731);
nand U23787 (N_23787,N_17156,N_17107);
xor U23788 (N_23788,N_19962,N_18168);
or U23789 (N_23789,N_19968,N_16671);
nor U23790 (N_23790,N_19502,N_18907);
and U23791 (N_23791,N_18103,N_15877);
xnor U23792 (N_23792,N_18361,N_19592);
nor U23793 (N_23793,N_17145,N_19965);
nand U23794 (N_23794,N_16985,N_18698);
nand U23795 (N_23795,N_16493,N_18587);
and U23796 (N_23796,N_18129,N_19571);
or U23797 (N_23797,N_16029,N_16792);
xor U23798 (N_23798,N_15971,N_18415);
nor U23799 (N_23799,N_18589,N_16043);
or U23800 (N_23800,N_18709,N_19519);
and U23801 (N_23801,N_19515,N_16366);
nor U23802 (N_23802,N_18179,N_15572);
and U23803 (N_23803,N_18164,N_15893);
nor U23804 (N_23804,N_16693,N_19523);
and U23805 (N_23805,N_16142,N_18279);
nand U23806 (N_23806,N_16666,N_16919);
and U23807 (N_23807,N_19367,N_15736);
nand U23808 (N_23808,N_15902,N_17306);
nand U23809 (N_23809,N_15156,N_15733);
xnor U23810 (N_23810,N_18245,N_19213);
and U23811 (N_23811,N_17065,N_19481);
or U23812 (N_23812,N_16985,N_15271);
or U23813 (N_23813,N_16302,N_15406);
nand U23814 (N_23814,N_17728,N_15320);
nor U23815 (N_23815,N_17982,N_16361);
and U23816 (N_23816,N_17291,N_17770);
or U23817 (N_23817,N_16170,N_19065);
nand U23818 (N_23818,N_18698,N_16113);
nor U23819 (N_23819,N_15957,N_19981);
nand U23820 (N_23820,N_19671,N_17022);
nand U23821 (N_23821,N_19031,N_16501);
nor U23822 (N_23822,N_16334,N_19310);
and U23823 (N_23823,N_19238,N_19748);
or U23824 (N_23824,N_19212,N_19839);
or U23825 (N_23825,N_18343,N_18583);
and U23826 (N_23826,N_15886,N_15040);
or U23827 (N_23827,N_19053,N_15300);
nand U23828 (N_23828,N_17410,N_16848);
nor U23829 (N_23829,N_15075,N_15179);
nor U23830 (N_23830,N_19988,N_18678);
and U23831 (N_23831,N_19176,N_16264);
nand U23832 (N_23832,N_19585,N_15309);
nand U23833 (N_23833,N_18495,N_19673);
nand U23834 (N_23834,N_19748,N_18775);
and U23835 (N_23835,N_16473,N_18143);
xnor U23836 (N_23836,N_17747,N_19236);
xnor U23837 (N_23837,N_15477,N_17956);
nor U23838 (N_23838,N_18321,N_17477);
or U23839 (N_23839,N_16549,N_18899);
and U23840 (N_23840,N_19293,N_19054);
nand U23841 (N_23841,N_16612,N_18824);
and U23842 (N_23842,N_19444,N_16809);
and U23843 (N_23843,N_15733,N_18846);
nand U23844 (N_23844,N_17583,N_19708);
and U23845 (N_23845,N_15432,N_18147);
and U23846 (N_23846,N_17145,N_15727);
or U23847 (N_23847,N_18849,N_16301);
or U23848 (N_23848,N_15745,N_19199);
and U23849 (N_23849,N_15750,N_16064);
or U23850 (N_23850,N_17423,N_16680);
and U23851 (N_23851,N_19838,N_19050);
and U23852 (N_23852,N_18347,N_18820);
and U23853 (N_23853,N_19188,N_15243);
nand U23854 (N_23854,N_16968,N_18857);
or U23855 (N_23855,N_17810,N_16313);
nor U23856 (N_23856,N_16911,N_16633);
or U23857 (N_23857,N_19008,N_15638);
and U23858 (N_23858,N_15599,N_19141);
nand U23859 (N_23859,N_18290,N_15624);
nand U23860 (N_23860,N_16704,N_15143);
nor U23861 (N_23861,N_19775,N_15028);
nor U23862 (N_23862,N_17402,N_19120);
nor U23863 (N_23863,N_18776,N_19742);
nand U23864 (N_23864,N_17535,N_16278);
nor U23865 (N_23865,N_16511,N_18021);
xor U23866 (N_23866,N_18462,N_18379);
nand U23867 (N_23867,N_19231,N_19167);
nand U23868 (N_23868,N_15651,N_15064);
nand U23869 (N_23869,N_16155,N_15494);
nand U23870 (N_23870,N_18192,N_18066);
xor U23871 (N_23871,N_16113,N_15433);
nor U23872 (N_23872,N_18452,N_17341);
nand U23873 (N_23873,N_17193,N_15723);
and U23874 (N_23874,N_19543,N_19045);
nand U23875 (N_23875,N_18118,N_15133);
and U23876 (N_23876,N_16664,N_18013);
nor U23877 (N_23877,N_17715,N_19175);
nand U23878 (N_23878,N_15901,N_15696);
and U23879 (N_23879,N_15725,N_19988);
or U23880 (N_23880,N_15833,N_16405);
or U23881 (N_23881,N_17531,N_17782);
or U23882 (N_23882,N_15725,N_16994);
xnor U23883 (N_23883,N_19732,N_17140);
or U23884 (N_23884,N_18215,N_16071);
nand U23885 (N_23885,N_16833,N_15452);
nand U23886 (N_23886,N_16685,N_15649);
and U23887 (N_23887,N_15418,N_19040);
and U23888 (N_23888,N_19687,N_16711);
nand U23889 (N_23889,N_18569,N_17927);
or U23890 (N_23890,N_19869,N_18499);
or U23891 (N_23891,N_19014,N_19827);
nor U23892 (N_23892,N_17458,N_18406);
nor U23893 (N_23893,N_18554,N_17837);
nor U23894 (N_23894,N_15607,N_15690);
or U23895 (N_23895,N_16562,N_15577);
and U23896 (N_23896,N_19637,N_19822);
or U23897 (N_23897,N_16352,N_18883);
nand U23898 (N_23898,N_17823,N_18993);
and U23899 (N_23899,N_19923,N_18674);
and U23900 (N_23900,N_17728,N_16102);
nand U23901 (N_23901,N_17825,N_16222);
nor U23902 (N_23902,N_19363,N_17894);
nor U23903 (N_23903,N_15282,N_18748);
and U23904 (N_23904,N_17458,N_18176);
nor U23905 (N_23905,N_15616,N_19323);
and U23906 (N_23906,N_15550,N_17689);
nand U23907 (N_23907,N_19278,N_17328);
nand U23908 (N_23908,N_18157,N_17102);
or U23909 (N_23909,N_15423,N_19072);
or U23910 (N_23910,N_16398,N_16958);
nor U23911 (N_23911,N_19777,N_16629);
or U23912 (N_23912,N_19887,N_17763);
or U23913 (N_23913,N_17557,N_18460);
nor U23914 (N_23914,N_17774,N_16399);
or U23915 (N_23915,N_16382,N_16793);
nor U23916 (N_23916,N_18709,N_17675);
and U23917 (N_23917,N_15762,N_16950);
nor U23918 (N_23918,N_18691,N_17827);
and U23919 (N_23919,N_16572,N_18134);
nor U23920 (N_23920,N_18500,N_16865);
or U23921 (N_23921,N_15531,N_19337);
xor U23922 (N_23922,N_15781,N_17040);
and U23923 (N_23923,N_19514,N_15231);
nand U23924 (N_23924,N_15875,N_16900);
xnor U23925 (N_23925,N_15920,N_18545);
nor U23926 (N_23926,N_18855,N_16491);
nor U23927 (N_23927,N_17089,N_18502);
nor U23928 (N_23928,N_18540,N_18968);
and U23929 (N_23929,N_15800,N_16353);
nor U23930 (N_23930,N_15580,N_17351);
nor U23931 (N_23931,N_17268,N_18955);
nor U23932 (N_23932,N_19099,N_18990);
or U23933 (N_23933,N_15553,N_17257);
nor U23934 (N_23934,N_16163,N_15234);
or U23935 (N_23935,N_16246,N_19970);
and U23936 (N_23936,N_16874,N_18472);
nor U23937 (N_23937,N_17587,N_17053);
nand U23938 (N_23938,N_19180,N_15765);
or U23939 (N_23939,N_16552,N_19604);
nand U23940 (N_23940,N_18642,N_15987);
nand U23941 (N_23941,N_16570,N_18637);
nand U23942 (N_23942,N_19256,N_19871);
nor U23943 (N_23943,N_17483,N_16562);
nor U23944 (N_23944,N_17205,N_19564);
nor U23945 (N_23945,N_18162,N_16379);
nand U23946 (N_23946,N_16318,N_16209);
and U23947 (N_23947,N_17897,N_18937);
nand U23948 (N_23948,N_16041,N_16743);
nor U23949 (N_23949,N_17934,N_18062);
and U23950 (N_23950,N_17651,N_16345);
or U23951 (N_23951,N_15844,N_16561);
nand U23952 (N_23952,N_17280,N_16048);
nand U23953 (N_23953,N_18422,N_19772);
and U23954 (N_23954,N_16107,N_17383);
nand U23955 (N_23955,N_15291,N_15743);
and U23956 (N_23956,N_16378,N_18188);
xnor U23957 (N_23957,N_17169,N_18475);
nor U23958 (N_23958,N_17597,N_15320);
xor U23959 (N_23959,N_17014,N_15931);
and U23960 (N_23960,N_19404,N_15864);
nand U23961 (N_23961,N_17042,N_17263);
or U23962 (N_23962,N_16550,N_16937);
or U23963 (N_23963,N_15334,N_15538);
nand U23964 (N_23964,N_19665,N_19922);
nor U23965 (N_23965,N_18443,N_16722);
or U23966 (N_23966,N_15976,N_17663);
or U23967 (N_23967,N_17283,N_18925);
or U23968 (N_23968,N_15726,N_15256);
nand U23969 (N_23969,N_16585,N_15035);
and U23970 (N_23970,N_15481,N_16191);
nand U23971 (N_23971,N_16668,N_17150);
nor U23972 (N_23972,N_19497,N_17337);
nand U23973 (N_23973,N_16147,N_19264);
nor U23974 (N_23974,N_15853,N_17164);
and U23975 (N_23975,N_15510,N_15772);
or U23976 (N_23976,N_16466,N_16243);
or U23977 (N_23977,N_17438,N_18565);
or U23978 (N_23978,N_16870,N_16131);
or U23979 (N_23979,N_15192,N_19801);
or U23980 (N_23980,N_15157,N_18905);
or U23981 (N_23981,N_19004,N_19231);
and U23982 (N_23982,N_19352,N_16888);
xnor U23983 (N_23983,N_17503,N_19299);
and U23984 (N_23984,N_15942,N_17573);
xnor U23985 (N_23985,N_17986,N_15211);
or U23986 (N_23986,N_18167,N_16432);
or U23987 (N_23987,N_15998,N_19760);
nand U23988 (N_23988,N_17389,N_16527);
xnor U23989 (N_23989,N_19781,N_18990);
nor U23990 (N_23990,N_17149,N_16519);
nor U23991 (N_23991,N_15940,N_17092);
nand U23992 (N_23992,N_17244,N_17408);
and U23993 (N_23993,N_19946,N_17755);
or U23994 (N_23994,N_16580,N_19245);
nand U23995 (N_23995,N_15015,N_15777);
nor U23996 (N_23996,N_15511,N_19880);
or U23997 (N_23997,N_15993,N_16318);
or U23998 (N_23998,N_17152,N_18580);
nor U23999 (N_23999,N_16165,N_15277);
or U24000 (N_24000,N_18673,N_19108);
nand U24001 (N_24001,N_16138,N_17451);
xor U24002 (N_24002,N_16052,N_16899);
nand U24003 (N_24003,N_18328,N_17779);
nand U24004 (N_24004,N_16153,N_18494);
xnor U24005 (N_24005,N_16740,N_15317);
nor U24006 (N_24006,N_19087,N_15730);
nand U24007 (N_24007,N_17493,N_15291);
or U24008 (N_24008,N_16251,N_15790);
xor U24009 (N_24009,N_16115,N_17769);
nor U24010 (N_24010,N_17245,N_15578);
nand U24011 (N_24011,N_19192,N_19886);
nor U24012 (N_24012,N_17235,N_17361);
xor U24013 (N_24013,N_19056,N_15113);
and U24014 (N_24014,N_19119,N_15757);
and U24015 (N_24015,N_18455,N_15900);
and U24016 (N_24016,N_19335,N_15338);
nand U24017 (N_24017,N_18663,N_17616);
nor U24018 (N_24018,N_19836,N_19551);
or U24019 (N_24019,N_16010,N_18161);
xor U24020 (N_24020,N_15060,N_17074);
or U24021 (N_24021,N_15929,N_19204);
and U24022 (N_24022,N_15496,N_18363);
or U24023 (N_24023,N_15539,N_17222);
nor U24024 (N_24024,N_15554,N_17328);
or U24025 (N_24025,N_17877,N_19847);
nor U24026 (N_24026,N_19693,N_19880);
and U24027 (N_24027,N_18746,N_17844);
nand U24028 (N_24028,N_18454,N_19496);
and U24029 (N_24029,N_17077,N_15954);
or U24030 (N_24030,N_19004,N_17940);
nor U24031 (N_24031,N_16324,N_18017);
and U24032 (N_24032,N_16945,N_15865);
or U24033 (N_24033,N_16372,N_16053);
and U24034 (N_24034,N_17875,N_19250);
nand U24035 (N_24035,N_15161,N_16441);
or U24036 (N_24036,N_16726,N_15197);
or U24037 (N_24037,N_15545,N_17765);
nand U24038 (N_24038,N_17878,N_15266);
and U24039 (N_24039,N_16247,N_16903);
xnor U24040 (N_24040,N_16152,N_18262);
or U24041 (N_24041,N_16238,N_18384);
or U24042 (N_24042,N_16809,N_18495);
and U24043 (N_24043,N_16190,N_19974);
nor U24044 (N_24044,N_17865,N_17307);
nor U24045 (N_24045,N_18967,N_18552);
or U24046 (N_24046,N_15967,N_16521);
and U24047 (N_24047,N_18601,N_19959);
or U24048 (N_24048,N_16254,N_15819);
nand U24049 (N_24049,N_15675,N_17959);
and U24050 (N_24050,N_15385,N_19275);
nand U24051 (N_24051,N_16126,N_18318);
nand U24052 (N_24052,N_17181,N_18017);
and U24053 (N_24053,N_17942,N_16188);
nand U24054 (N_24054,N_17009,N_18013);
nand U24055 (N_24055,N_19808,N_15651);
nand U24056 (N_24056,N_17211,N_16386);
nand U24057 (N_24057,N_18190,N_15171);
nor U24058 (N_24058,N_16202,N_15081);
nand U24059 (N_24059,N_16746,N_15059);
or U24060 (N_24060,N_16932,N_17600);
nand U24061 (N_24061,N_15890,N_16015);
or U24062 (N_24062,N_17642,N_15427);
nor U24063 (N_24063,N_17204,N_19928);
nand U24064 (N_24064,N_17160,N_16707);
and U24065 (N_24065,N_17947,N_19193);
nor U24066 (N_24066,N_17576,N_17618);
nor U24067 (N_24067,N_19928,N_18516);
nand U24068 (N_24068,N_19377,N_16063);
nor U24069 (N_24069,N_16825,N_19083);
nor U24070 (N_24070,N_15380,N_15621);
or U24071 (N_24071,N_15467,N_19263);
nand U24072 (N_24072,N_19118,N_19490);
xor U24073 (N_24073,N_18895,N_16914);
and U24074 (N_24074,N_19668,N_19689);
or U24075 (N_24075,N_19986,N_17833);
nor U24076 (N_24076,N_19675,N_16864);
nor U24077 (N_24077,N_15027,N_15981);
nor U24078 (N_24078,N_17118,N_19866);
and U24079 (N_24079,N_17946,N_18060);
nor U24080 (N_24080,N_16521,N_16805);
or U24081 (N_24081,N_17376,N_17890);
nor U24082 (N_24082,N_19948,N_16518);
xor U24083 (N_24083,N_16980,N_15836);
or U24084 (N_24084,N_16975,N_18252);
or U24085 (N_24085,N_16988,N_15865);
xnor U24086 (N_24086,N_17912,N_19471);
or U24087 (N_24087,N_18850,N_19281);
or U24088 (N_24088,N_16262,N_19215);
nor U24089 (N_24089,N_19396,N_17726);
or U24090 (N_24090,N_15061,N_19073);
and U24091 (N_24091,N_16807,N_18368);
nand U24092 (N_24092,N_17949,N_16184);
nor U24093 (N_24093,N_16499,N_16966);
and U24094 (N_24094,N_15893,N_19582);
nand U24095 (N_24095,N_15352,N_15005);
nand U24096 (N_24096,N_18676,N_17540);
xnor U24097 (N_24097,N_15214,N_17307);
nor U24098 (N_24098,N_15369,N_19482);
nor U24099 (N_24099,N_19186,N_16755);
nand U24100 (N_24100,N_15699,N_17091);
nand U24101 (N_24101,N_18851,N_17178);
nor U24102 (N_24102,N_16081,N_15757);
nand U24103 (N_24103,N_19029,N_16892);
and U24104 (N_24104,N_17834,N_18015);
xor U24105 (N_24105,N_16435,N_19144);
nand U24106 (N_24106,N_19481,N_16511);
or U24107 (N_24107,N_16560,N_18234);
or U24108 (N_24108,N_18338,N_19884);
or U24109 (N_24109,N_19152,N_17803);
nand U24110 (N_24110,N_16395,N_15355);
or U24111 (N_24111,N_17101,N_15276);
or U24112 (N_24112,N_15398,N_15760);
and U24113 (N_24113,N_18698,N_18871);
and U24114 (N_24114,N_17706,N_18276);
or U24115 (N_24115,N_18170,N_16934);
or U24116 (N_24116,N_19008,N_15327);
or U24117 (N_24117,N_17110,N_16514);
or U24118 (N_24118,N_18761,N_17135);
or U24119 (N_24119,N_17427,N_19895);
or U24120 (N_24120,N_18425,N_16455);
nor U24121 (N_24121,N_17850,N_18745);
and U24122 (N_24122,N_18056,N_19268);
nor U24123 (N_24123,N_15036,N_17660);
or U24124 (N_24124,N_17097,N_15967);
or U24125 (N_24125,N_18324,N_16647);
or U24126 (N_24126,N_18126,N_17992);
or U24127 (N_24127,N_19410,N_16538);
or U24128 (N_24128,N_17835,N_18060);
xnor U24129 (N_24129,N_17952,N_15995);
nor U24130 (N_24130,N_16707,N_15474);
nand U24131 (N_24131,N_19375,N_17643);
or U24132 (N_24132,N_18792,N_17749);
or U24133 (N_24133,N_18502,N_18474);
or U24134 (N_24134,N_15664,N_17866);
nor U24135 (N_24135,N_15460,N_19729);
nand U24136 (N_24136,N_15133,N_15426);
nor U24137 (N_24137,N_16541,N_17161);
nand U24138 (N_24138,N_15060,N_15208);
or U24139 (N_24139,N_18208,N_15331);
xor U24140 (N_24140,N_16118,N_17289);
nand U24141 (N_24141,N_15101,N_19555);
nand U24142 (N_24142,N_15282,N_16843);
and U24143 (N_24143,N_16576,N_16929);
or U24144 (N_24144,N_19215,N_17372);
and U24145 (N_24145,N_15361,N_17104);
nand U24146 (N_24146,N_16667,N_17057);
nor U24147 (N_24147,N_15080,N_15114);
nand U24148 (N_24148,N_18816,N_19632);
or U24149 (N_24149,N_18033,N_15900);
nand U24150 (N_24150,N_19554,N_18331);
or U24151 (N_24151,N_16320,N_16240);
or U24152 (N_24152,N_16673,N_19761);
nand U24153 (N_24153,N_16635,N_17285);
nor U24154 (N_24154,N_18853,N_17345);
nor U24155 (N_24155,N_15321,N_19360);
nand U24156 (N_24156,N_15003,N_18501);
nand U24157 (N_24157,N_16737,N_16062);
or U24158 (N_24158,N_17806,N_15867);
and U24159 (N_24159,N_18391,N_18778);
or U24160 (N_24160,N_19123,N_16011);
or U24161 (N_24161,N_19781,N_18019);
and U24162 (N_24162,N_16107,N_15107);
nand U24163 (N_24163,N_16604,N_17736);
nor U24164 (N_24164,N_16438,N_15951);
nand U24165 (N_24165,N_19398,N_16984);
nor U24166 (N_24166,N_19352,N_17396);
or U24167 (N_24167,N_15809,N_19615);
xnor U24168 (N_24168,N_19489,N_19536);
nand U24169 (N_24169,N_15420,N_17238);
xnor U24170 (N_24170,N_15166,N_19858);
and U24171 (N_24171,N_16940,N_16004);
and U24172 (N_24172,N_17021,N_17246);
nor U24173 (N_24173,N_17622,N_16382);
or U24174 (N_24174,N_17983,N_19414);
or U24175 (N_24175,N_19643,N_15524);
nor U24176 (N_24176,N_16866,N_17066);
nor U24177 (N_24177,N_17482,N_19847);
nand U24178 (N_24178,N_19918,N_15794);
nand U24179 (N_24179,N_18258,N_17266);
and U24180 (N_24180,N_17718,N_19954);
nand U24181 (N_24181,N_17720,N_16182);
nor U24182 (N_24182,N_17065,N_17498);
nand U24183 (N_24183,N_16314,N_15775);
nand U24184 (N_24184,N_15055,N_16339);
nor U24185 (N_24185,N_15236,N_15214);
nor U24186 (N_24186,N_18279,N_16405);
nand U24187 (N_24187,N_17142,N_17391);
and U24188 (N_24188,N_17995,N_19068);
or U24189 (N_24189,N_17693,N_16238);
nand U24190 (N_24190,N_17892,N_18409);
or U24191 (N_24191,N_15618,N_15198);
or U24192 (N_24192,N_18878,N_17509);
and U24193 (N_24193,N_16757,N_16597);
nand U24194 (N_24194,N_17638,N_18882);
nor U24195 (N_24195,N_15034,N_16276);
and U24196 (N_24196,N_17076,N_17004);
nand U24197 (N_24197,N_18041,N_19736);
and U24198 (N_24198,N_18894,N_15827);
nor U24199 (N_24199,N_18981,N_15280);
and U24200 (N_24200,N_19005,N_19040);
and U24201 (N_24201,N_19810,N_16628);
xor U24202 (N_24202,N_18581,N_18733);
nor U24203 (N_24203,N_16492,N_17586);
nand U24204 (N_24204,N_15268,N_18333);
xor U24205 (N_24205,N_17869,N_15502);
or U24206 (N_24206,N_18387,N_19913);
or U24207 (N_24207,N_17376,N_18187);
or U24208 (N_24208,N_18852,N_16947);
and U24209 (N_24209,N_17790,N_17659);
or U24210 (N_24210,N_19787,N_16438);
nand U24211 (N_24211,N_15816,N_19897);
and U24212 (N_24212,N_17432,N_18136);
nand U24213 (N_24213,N_15849,N_18355);
xnor U24214 (N_24214,N_18757,N_15547);
nor U24215 (N_24215,N_16738,N_15623);
nor U24216 (N_24216,N_17978,N_19201);
nor U24217 (N_24217,N_18595,N_16702);
nor U24218 (N_24218,N_15729,N_18988);
nand U24219 (N_24219,N_16818,N_19628);
xor U24220 (N_24220,N_18774,N_19381);
nor U24221 (N_24221,N_19444,N_19769);
nand U24222 (N_24222,N_15227,N_16129);
or U24223 (N_24223,N_19841,N_19675);
and U24224 (N_24224,N_19349,N_16624);
and U24225 (N_24225,N_18969,N_17128);
or U24226 (N_24226,N_15735,N_19751);
or U24227 (N_24227,N_18515,N_19570);
or U24228 (N_24228,N_19917,N_19053);
xnor U24229 (N_24229,N_17532,N_15129);
xnor U24230 (N_24230,N_16702,N_16044);
or U24231 (N_24231,N_15154,N_15110);
or U24232 (N_24232,N_18087,N_18188);
nand U24233 (N_24233,N_18121,N_19771);
or U24234 (N_24234,N_17620,N_16410);
nor U24235 (N_24235,N_17233,N_18645);
or U24236 (N_24236,N_15595,N_19578);
nor U24237 (N_24237,N_15244,N_17100);
and U24238 (N_24238,N_16249,N_18950);
or U24239 (N_24239,N_18252,N_16597);
nand U24240 (N_24240,N_16246,N_17418);
and U24241 (N_24241,N_18418,N_15039);
and U24242 (N_24242,N_15707,N_15918);
and U24243 (N_24243,N_17717,N_19056);
nand U24244 (N_24244,N_17924,N_18135);
nand U24245 (N_24245,N_18265,N_19536);
nor U24246 (N_24246,N_15658,N_15642);
and U24247 (N_24247,N_19803,N_17975);
or U24248 (N_24248,N_16858,N_15883);
or U24249 (N_24249,N_17963,N_19164);
nand U24250 (N_24250,N_17773,N_18113);
and U24251 (N_24251,N_15070,N_17726);
nor U24252 (N_24252,N_17802,N_17576);
nor U24253 (N_24253,N_18592,N_18606);
nand U24254 (N_24254,N_15398,N_15355);
and U24255 (N_24255,N_17427,N_18411);
nand U24256 (N_24256,N_15250,N_19615);
or U24257 (N_24257,N_19406,N_15163);
or U24258 (N_24258,N_15729,N_19448);
xnor U24259 (N_24259,N_16095,N_17660);
or U24260 (N_24260,N_19003,N_17989);
nand U24261 (N_24261,N_16418,N_19800);
and U24262 (N_24262,N_16388,N_15389);
nand U24263 (N_24263,N_19070,N_18829);
or U24264 (N_24264,N_15639,N_16751);
xor U24265 (N_24265,N_17489,N_15785);
or U24266 (N_24266,N_15406,N_17051);
xnor U24267 (N_24267,N_19379,N_15174);
nand U24268 (N_24268,N_18273,N_19375);
nor U24269 (N_24269,N_16645,N_16606);
or U24270 (N_24270,N_19022,N_17751);
nor U24271 (N_24271,N_17732,N_17990);
nand U24272 (N_24272,N_18637,N_19796);
xor U24273 (N_24273,N_15861,N_17666);
or U24274 (N_24274,N_15474,N_18428);
nor U24275 (N_24275,N_16735,N_16017);
xnor U24276 (N_24276,N_15159,N_18197);
and U24277 (N_24277,N_17862,N_19538);
nand U24278 (N_24278,N_17468,N_19330);
or U24279 (N_24279,N_15013,N_15469);
and U24280 (N_24280,N_17772,N_16806);
or U24281 (N_24281,N_19197,N_18876);
or U24282 (N_24282,N_18646,N_17045);
and U24283 (N_24283,N_19279,N_17876);
nor U24284 (N_24284,N_16910,N_15467);
and U24285 (N_24285,N_16426,N_15039);
and U24286 (N_24286,N_15284,N_16825);
and U24287 (N_24287,N_17550,N_15617);
nor U24288 (N_24288,N_19804,N_17787);
nor U24289 (N_24289,N_16800,N_16365);
nand U24290 (N_24290,N_18506,N_17443);
xor U24291 (N_24291,N_19366,N_18484);
or U24292 (N_24292,N_16372,N_17105);
or U24293 (N_24293,N_18451,N_15528);
or U24294 (N_24294,N_19845,N_17866);
nor U24295 (N_24295,N_17504,N_15412);
nand U24296 (N_24296,N_16240,N_17121);
xor U24297 (N_24297,N_17390,N_15464);
nand U24298 (N_24298,N_15840,N_19007);
or U24299 (N_24299,N_16583,N_19673);
nand U24300 (N_24300,N_17885,N_17031);
and U24301 (N_24301,N_18539,N_19964);
nand U24302 (N_24302,N_16436,N_17795);
xnor U24303 (N_24303,N_15083,N_18887);
nor U24304 (N_24304,N_17045,N_17674);
and U24305 (N_24305,N_19137,N_15906);
and U24306 (N_24306,N_17272,N_15376);
nor U24307 (N_24307,N_16332,N_16079);
xor U24308 (N_24308,N_17874,N_19351);
nand U24309 (N_24309,N_18103,N_17279);
nand U24310 (N_24310,N_19966,N_16063);
and U24311 (N_24311,N_15773,N_16358);
nand U24312 (N_24312,N_15120,N_17747);
and U24313 (N_24313,N_18441,N_18534);
xnor U24314 (N_24314,N_16195,N_16430);
nand U24315 (N_24315,N_18540,N_15960);
or U24316 (N_24316,N_19850,N_17691);
nand U24317 (N_24317,N_15128,N_16345);
nand U24318 (N_24318,N_17675,N_17030);
and U24319 (N_24319,N_17905,N_19804);
or U24320 (N_24320,N_17402,N_17423);
nor U24321 (N_24321,N_15424,N_15890);
nand U24322 (N_24322,N_15508,N_16500);
or U24323 (N_24323,N_17990,N_17100);
or U24324 (N_24324,N_19709,N_18413);
nor U24325 (N_24325,N_15744,N_19568);
nand U24326 (N_24326,N_15115,N_18053);
nor U24327 (N_24327,N_15578,N_17596);
and U24328 (N_24328,N_19709,N_19777);
nand U24329 (N_24329,N_19353,N_19509);
or U24330 (N_24330,N_19241,N_19663);
and U24331 (N_24331,N_17478,N_16853);
and U24332 (N_24332,N_15043,N_18057);
or U24333 (N_24333,N_17073,N_17046);
nand U24334 (N_24334,N_16382,N_15501);
and U24335 (N_24335,N_15019,N_16929);
xnor U24336 (N_24336,N_19874,N_18498);
nor U24337 (N_24337,N_18351,N_17438);
nor U24338 (N_24338,N_19534,N_15764);
nor U24339 (N_24339,N_16180,N_15954);
nand U24340 (N_24340,N_15484,N_15287);
nand U24341 (N_24341,N_17011,N_16388);
nor U24342 (N_24342,N_15298,N_19177);
nor U24343 (N_24343,N_17963,N_19358);
and U24344 (N_24344,N_17702,N_18282);
or U24345 (N_24345,N_16480,N_15437);
and U24346 (N_24346,N_17636,N_18166);
or U24347 (N_24347,N_19244,N_16990);
or U24348 (N_24348,N_19841,N_16004);
or U24349 (N_24349,N_17413,N_16427);
nor U24350 (N_24350,N_19680,N_16168);
or U24351 (N_24351,N_17447,N_15472);
nand U24352 (N_24352,N_16936,N_16335);
or U24353 (N_24353,N_17033,N_15195);
and U24354 (N_24354,N_16669,N_18770);
nand U24355 (N_24355,N_17124,N_18616);
nand U24356 (N_24356,N_15674,N_17798);
nor U24357 (N_24357,N_16187,N_17740);
or U24358 (N_24358,N_19312,N_18502);
or U24359 (N_24359,N_19773,N_16512);
xnor U24360 (N_24360,N_16368,N_17073);
or U24361 (N_24361,N_17136,N_18263);
nand U24362 (N_24362,N_16145,N_19308);
nand U24363 (N_24363,N_17728,N_16327);
and U24364 (N_24364,N_16339,N_18673);
nand U24365 (N_24365,N_18052,N_18725);
nand U24366 (N_24366,N_17394,N_19179);
and U24367 (N_24367,N_16655,N_19771);
or U24368 (N_24368,N_15753,N_19271);
nand U24369 (N_24369,N_19246,N_15239);
nand U24370 (N_24370,N_15991,N_18889);
or U24371 (N_24371,N_16955,N_19077);
nor U24372 (N_24372,N_19405,N_16928);
xor U24373 (N_24373,N_19290,N_15042);
and U24374 (N_24374,N_17989,N_18157);
or U24375 (N_24375,N_15643,N_15335);
or U24376 (N_24376,N_15601,N_15588);
nor U24377 (N_24377,N_15937,N_17378);
xor U24378 (N_24378,N_17916,N_19088);
and U24379 (N_24379,N_16143,N_17118);
and U24380 (N_24380,N_16668,N_18948);
and U24381 (N_24381,N_17883,N_17768);
xnor U24382 (N_24382,N_18092,N_19820);
nor U24383 (N_24383,N_18085,N_17713);
and U24384 (N_24384,N_15394,N_17491);
nor U24385 (N_24385,N_15939,N_16305);
or U24386 (N_24386,N_19173,N_15739);
nor U24387 (N_24387,N_17635,N_18348);
and U24388 (N_24388,N_17996,N_16119);
or U24389 (N_24389,N_16086,N_17578);
nor U24390 (N_24390,N_19780,N_19819);
and U24391 (N_24391,N_18395,N_17154);
or U24392 (N_24392,N_19554,N_15274);
and U24393 (N_24393,N_16700,N_19534);
nand U24394 (N_24394,N_15258,N_17479);
nor U24395 (N_24395,N_19080,N_18907);
and U24396 (N_24396,N_18713,N_17679);
and U24397 (N_24397,N_16674,N_16201);
and U24398 (N_24398,N_16150,N_15023);
nand U24399 (N_24399,N_19495,N_15705);
nor U24400 (N_24400,N_18908,N_18151);
or U24401 (N_24401,N_17153,N_17681);
nand U24402 (N_24402,N_16578,N_17090);
or U24403 (N_24403,N_17153,N_17829);
and U24404 (N_24404,N_19966,N_17172);
xor U24405 (N_24405,N_17102,N_19683);
or U24406 (N_24406,N_18974,N_17550);
and U24407 (N_24407,N_17955,N_16635);
xor U24408 (N_24408,N_19321,N_15397);
xnor U24409 (N_24409,N_15099,N_17562);
and U24410 (N_24410,N_16117,N_17499);
nor U24411 (N_24411,N_18442,N_19458);
xnor U24412 (N_24412,N_16510,N_19251);
nand U24413 (N_24413,N_16217,N_16343);
and U24414 (N_24414,N_17499,N_19091);
and U24415 (N_24415,N_18824,N_19683);
and U24416 (N_24416,N_17109,N_16696);
nand U24417 (N_24417,N_17131,N_16989);
and U24418 (N_24418,N_19896,N_19716);
nand U24419 (N_24419,N_19289,N_18646);
nand U24420 (N_24420,N_17696,N_17931);
and U24421 (N_24421,N_19554,N_19350);
nor U24422 (N_24422,N_16838,N_16095);
and U24423 (N_24423,N_18325,N_18662);
nand U24424 (N_24424,N_19684,N_15218);
nand U24425 (N_24425,N_17755,N_16523);
and U24426 (N_24426,N_16212,N_18917);
xnor U24427 (N_24427,N_18765,N_15897);
nor U24428 (N_24428,N_19064,N_18498);
and U24429 (N_24429,N_18264,N_19267);
nand U24430 (N_24430,N_17256,N_16583);
nor U24431 (N_24431,N_17839,N_18835);
xnor U24432 (N_24432,N_15423,N_17580);
and U24433 (N_24433,N_17262,N_19131);
and U24434 (N_24434,N_15510,N_18898);
nor U24435 (N_24435,N_18799,N_16298);
and U24436 (N_24436,N_18404,N_17897);
or U24437 (N_24437,N_16851,N_17511);
xor U24438 (N_24438,N_15690,N_16667);
xor U24439 (N_24439,N_17088,N_19902);
nor U24440 (N_24440,N_19736,N_16277);
or U24441 (N_24441,N_18527,N_15099);
and U24442 (N_24442,N_15468,N_15049);
and U24443 (N_24443,N_19512,N_19343);
or U24444 (N_24444,N_17134,N_18680);
and U24445 (N_24445,N_16614,N_19672);
nand U24446 (N_24446,N_18503,N_16115);
or U24447 (N_24447,N_16316,N_15165);
nor U24448 (N_24448,N_15836,N_18191);
or U24449 (N_24449,N_19941,N_19668);
xnor U24450 (N_24450,N_18488,N_16068);
nor U24451 (N_24451,N_19007,N_15945);
nand U24452 (N_24452,N_19931,N_19667);
and U24453 (N_24453,N_18729,N_19731);
nand U24454 (N_24454,N_15558,N_15079);
or U24455 (N_24455,N_18080,N_16108);
nand U24456 (N_24456,N_16259,N_17202);
xnor U24457 (N_24457,N_19970,N_19945);
nand U24458 (N_24458,N_16819,N_16761);
nand U24459 (N_24459,N_19267,N_16868);
nor U24460 (N_24460,N_17032,N_18612);
nor U24461 (N_24461,N_15430,N_15307);
and U24462 (N_24462,N_17899,N_16932);
and U24463 (N_24463,N_17030,N_18689);
or U24464 (N_24464,N_18662,N_17183);
or U24465 (N_24465,N_17707,N_15483);
nor U24466 (N_24466,N_19470,N_16412);
nor U24467 (N_24467,N_16200,N_17042);
or U24468 (N_24468,N_18357,N_19108);
nand U24469 (N_24469,N_15793,N_15957);
nand U24470 (N_24470,N_16720,N_15622);
nor U24471 (N_24471,N_16682,N_19490);
and U24472 (N_24472,N_19335,N_19173);
nand U24473 (N_24473,N_15501,N_19387);
nor U24474 (N_24474,N_15910,N_15219);
nand U24475 (N_24475,N_17666,N_19263);
or U24476 (N_24476,N_16516,N_19508);
nand U24477 (N_24477,N_16956,N_17284);
nand U24478 (N_24478,N_19752,N_17716);
or U24479 (N_24479,N_15334,N_19728);
and U24480 (N_24480,N_18041,N_15435);
xor U24481 (N_24481,N_17019,N_18740);
xor U24482 (N_24482,N_19312,N_16476);
xor U24483 (N_24483,N_15774,N_18597);
nand U24484 (N_24484,N_17613,N_18866);
nand U24485 (N_24485,N_19059,N_15316);
nand U24486 (N_24486,N_17585,N_18717);
nand U24487 (N_24487,N_18171,N_18460);
and U24488 (N_24488,N_16541,N_15105);
or U24489 (N_24489,N_19617,N_15556);
or U24490 (N_24490,N_16684,N_18183);
xnor U24491 (N_24491,N_19894,N_17781);
nand U24492 (N_24492,N_15450,N_19481);
nor U24493 (N_24493,N_15021,N_19384);
nand U24494 (N_24494,N_18247,N_17670);
nand U24495 (N_24495,N_19172,N_18809);
nor U24496 (N_24496,N_17318,N_15851);
nor U24497 (N_24497,N_17935,N_17361);
nand U24498 (N_24498,N_17078,N_15754);
or U24499 (N_24499,N_19928,N_19017);
or U24500 (N_24500,N_16758,N_19704);
nor U24501 (N_24501,N_19388,N_19856);
or U24502 (N_24502,N_19189,N_19356);
and U24503 (N_24503,N_17729,N_17254);
or U24504 (N_24504,N_18271,N_18196);
nor U24505 (N_24505,N_18979,N_17022);
and U24506 (N_24506,N_17973,N_15092);
xor U24507 (N_24507,N_18868,N_19312);
or U24508 (N_24508,N_16473,N_18851);
nand U24509 (N_24509,N_19802,N_18553);
and U24510 (N_24510,N_19315,N_16182);
or U24511 (N_24511,N_16396,N_18817);
or U24512 (N_24512,N_19979,N_15062);
or U24513 (N_24513,N_19136,N_16802);
and U24514 (N_24514,N_19130,N_15394);
or U24515 (N_24515,N_16664,N_18899);
or U24516 (N_24516,N_19487,N_17021);
nor U24517 (N_24517,N_16955,N_17886);
and U24518 (N_24518,N_15281,N_19170);
or U24519 (N_24519,N_19688,N_16820);
and U24520 (N_24520,N_17790,N_16494);
nand U24521 (N_24521,N_19556,N_19070);
and U24522 (N_24522,N_17272,N_19276);
and U24523 (N_24523,N_15044,N_15985);
or U24524 (N_24524,N_19821,N_16746);
nand U24525 (N_24525,N_16380,N_17866);
nand U24526 (N_24526,N_16834,N_15480);
nor U24527 (N_24527,N_19318,N_15592);
nand U24528 (N_24528,N_18111,N_16435);
nor U24529 (N_24529,N_15434,N_19939);
xor U24530 (N_24530,N_19232,N_17384);
and U24531 (N_24531,N_17448,N_16429);
and U24532 (N_24532,N_18307,N_19231);
xor U24533 (N_24533,N_19978,N_18834);
nor U24534 (N_24534,N_18841,N_17266);
nor U24535 (N_24535,N_17622,N_19864);
and U24536 (N_24536,N_15640,N_16545);
nand U24537 (N_24537,N_18809,N_17426);
nor U24538 (N_24538,N_16461,N_17393);
nand U24539 (N_24539,N_17021,N_16901);
nand U24540 (N_24540,N_15051,N_15263);
and U24541 (N_24541,N_17554,N_19467);
nand U24542 (N_24542,N_15511,N_17314);
and U24543 (N_24543,N_19621,N_19532);
and U24544 (N_24544,N_15048,N_16890);
nor U24545 (N_24545,N_17246,N_17673);
xor U24546 (N_24546,N_16006,N_18526);
or U24547 (N_24547,N_18035,N_16072);
nor U24548 (N_24548,N_19437,N_16673);
nor U24549 (N_24549,N_15433,N_18065);
nand U24550 (N_24550,N_18263,N_17133);
nor U24551 (N_24551,N_19569,N_15323);
and U24552 (N_24552,N_15012,N_19842);
or U24553 (N_24553,N_17874,N_16039);
nand U24554 (N_24554,N_16546,N_18446);
and U24555 (N_24555,N_18195,N_16197);
nand U24556 (N_24556,N_15077,N_15859);
nand U24557 (N_24557,N_17985,N_17353);
and U24558 (N_24558,N_19180,N_17762);
or U24559 (N_24559,N_18065,N_15970);
nand U24560 (N_24560,N_18414,N_19909);
nand U24561 (N_24561,N_19544,N_17640);
nand U24562 (N_24562,N_16559,N_17541);
or U24563 (N_24563,N_17552,N_18965);
xnor U24564 (N_24564,N_19501,N_15717);
nor U24565 (N_24565,N_16732,N_17295);
or U24566 (N_24566,N_15509,N_17936);
and U24567 (N_24567,N_18102,N_17457);
nand U24568 (N_24568,N_15412,N_15291);
or U24569 (N_24569,N_18726,N_17236);
nor U24570 (N_24570,N_16873,N_17700);
and U24571 (N_24571,N_19335,N_15522);
or U24572 (N_24572,N_15035,N_15811);
and U24573 (N_24573,N_15965,N_18343);
nor U24574 (N_24574,N_16329,N_17314);
or U24575 (N_24575,N_19709,N_15312);
and U24576 (N_24576,N_18318,N_17331);
or U24577 (N_24577,N_18868,N_16467);
nor U24578 (N_24578,N_16825,N_15663);
and U24579 (N_24579,N_16619,N_17387);
nor U24580 (N_24580,N_19572,N_17966);
and U24581 (N_24581,N_19292,N_18713);
and U24582 (N_24582,N_15528,N_17532);
and U24583 (N_24583,N_19405,N_16248);
nor U24584 (N_24584,N_19731,N_19736);
nand U24585 (N_24585,N_15327,N_18395);
nor U24586 (N_24586,N_16038,N_16923);
xor U24587 (N_24587,N_19936,N_19100);
nand U24588 (N_24588,N_19595,N_18536);
or U24589 (N_24589,N_15617,N_15917);
and U24590 (N_24590,N_16233,N_18467);
or U24591 (N_24591,N_15889,N_19905);
nand U24592 (N_24592,N_18808,N_18460);
or U24593 (N_24593,N_16046,N_15540);
nor U24594 (N_24594,N_16800,N_19364);
nor U24595 (N_24595,N_15672,N_19061);
nand U24596 (N_24596,N_16890,N_15688);
and U24597 (N_24597,N_19612,N_16923);
xor U24598 (N_24598,N_18219,N_16207);
and U24599 (N_24599,N_15452,N_17008);
nand U24600 (N_24600,N_16379,N_19652);
nand U24601 (N_24601,N_16810,N_19567);
nor U24602 (N_24602,N_17466,N_17567);
or U24603 (N_24603,N_16681,N_16528);
or U24604 (N_24604,N_16948,N_16411);
nor U24605 (N_24605,N_18025,N_19791);
nor U24606 (N_24606,N_15474,N_17810);
nand U24607 (N_24607,N_16607,N_18624);
nand U24608 (N_24608,N_16935,N_19694);
xor U24609 (N_24609,N_16798,N_15156);
nand U24610 (N_24610,N_19152,N_17617);
or U24611 (N_24611,N_16643,N_15665);
nor U24612 (N_24612,N_18669,N_16467);
or U24613 (N_24613,N_15121,N_18165);
or U24614 (N_24614,N_18999,N_16465);
or U24615 (N_24615,N_19433,N_17113);
nor U24616 (N_24616,N_18409,N_15278);
nand U24617 (N_24617,N_15162,N_16115);
nor U24618 (N_24618,N_17136,N_16364);
nor U24619 (N_24619,N_18863,N_16500);
nor U24620 (N_24620,N_18674,N_19292);
or U24621 (N_24621,N_18479,N_16328);
or U24622 (N_24622,N_18018,N_19421);
nand U24623 (N_24623,N_16393,N_16169);
xnor U24624 (N_24624,N_19710,N_18066);
xnor U24625 (N_24625,N_18552,N_18211);
nand U24626 (N_24626,N_17899,N_18651);
and U24627 (N_24627,N_16990,N_15391);
nand U24628 (N_24628,N_19911,N_18635);
nand U24629 (N_24629,N_16100,N_15614);
xnor U24630 (N_24630,N_15538,N_17888);
or U24631 (N_24631,N_17042,N_16250);
xor U24632 (N_24632,N_17941,N_19264);
nor U24633 (N_24633,N_15036,N_17522);
nor U24634 (N_24634,N_19090,N_15240);
nand U24635 (N_24635,N_18283,N_19591);
nor U24636 (N_24636,N_19346,N_17645);
nor U24637 (N_24637,N_17689,N_18936);
or U24638 (N_24638,N_18190,N_17548);
and U24639 (N_24639,N_16249,N_15906);
nand U24640 (N_24640,N_18044,N_17055);
or U24641 (N_24641,N_15564,N_19816);
or U24642 (N_24642,N_18716,N_18125);
nor U24643 (N_24643,N_19302,N_15120);
nand U24644 (N_24644,N_16464,N_15813);
and U24645 (N_24645,N_16190,N_15797);
nor U24646 (N_24646,N_18096,N_16012);
nor U24647 (N_24647,N_16360,N_19747);
or U24648 (N_24648,N_18318,N_15675);
nor U24649 (N_24649,N_15062,N_19663);
nand U24650 (N_24650,N_17559,N_17926);
nor U24651 (N_24651,N_16086,N_16018);
nor U24652 (N_24652,N_17688,N_15186);
and U24653 (N_24653,N_16969,N_16108);
xor U24654 (N_24654,N_17234,N_18757);
nand U24655 (N_24655,N_16270,N_16294);
and U24656 (N_24656,N_15728,N_15137);
xnor U24657 (N_24657,N_15932,N_18298);
and U24658 (N_24658,N_15592,N_17050);
and U24659 (N_24659,N_17539,N_16843);
nor U24660 (N_24660,N_17053,N_19916);
and U24661 (N_24661,N_16840,N_18602);
or U24662 (N_24662,N_16416,N_15145);
and U24663 (N_24663,N_19488,N_19138);
nor U24664 (N_24664,N_17014,N_17283);
or U24665 (N_24665,N_18293,N_18755);
nand U24666 (N_24666,N_17408,N_18493);
nand U24667 (N_24667,N_18634,N_18119);
nand U24668 (N_24668,N_17478,N_18705);
nor U24669 (N_24669,N_17805,N_15366);
or U24670 (N_24670,N_16682,N_16727);
nand U24671 (N_24671,N_17549,N_17264);
or U24672 (N_24672,N_16818,N_19459);
xnor U24673 (N_24673,N_18559,N_17442);
and U24674 (N_24674,N_15991,N_18768);
and U24675 (N_24675,N_17092,N_18156);
nor U24676 (N_24676,N_19655,N_16879);
nor U24677 (N_24677,N_19061,N_17896);
and U24678 (N_24678,N_15181,N_15948);
and U24679 (N_24679,N_16121,N_16099);
nand U24680 (N_24680,N_16690,N_18035);
and U24681 (N_24681,N_19721,N_18817);
and U24682 (N_24682,N_15060,N_19357);
and U24683 (N_24683,N_19980,N_15812);
xnor U24684 (N_24684,N_16188,N_15268);
nand U24685 (N_24685,N_19182,N_18332);
or U24686 (N_24686,N_19716,N_17064);
nand U24687 (N_24687,N_18494,N_19169);
nand U24688 (N_24688,N_19779,N_17147);
and U24689 (N_24689,N_19571,N_16194);
nor U24690 (N_24690,N_18887,N_18781);
nor U24691 (N_24691,N_18152,N_16057);
and U24692 (N_24692,N_19636,N_16644);
or U24693 (N_24693,N_15872,N_15527);
xnor U24694 (N_24694,N_16187,N_17849);
and U24695 (N_24695,N_18118,N_15505);
nor U24696 (N_24696,N_18536,N_19520);
xor U24697 (N_24697,N_18963,N_18800);
nor U24698 (N_24698,N_16466,N_16714);
nor U24699 (N_24699,N_17790,N_18932);
or U24700 (N_24700,N_19500,N_18683);
and U24701 (N_24701,N_19754,N_18208);
and U24702 (N_24702,N_17305,N_18443);
or U24703 (N_24703,N_17591,N_16943);
xor U24704 (N_24704,N_15576,N_17786);
nor U24705 (N_24705,N_17469,N_15625);
nand U24706 (N_24706,N_18195,N_15230);
nor U24707 (N_24707,N_15909,N_17359);
nand U24708 (N_24708,N_17227,N_19466);
and U24709 (N_24709,N_15362,N_15153);
nor U24710 (N_24710,N_17029,N_15743);
or U24711 (N_24711,N_19967,N_17589);
nand U24712 (N_24712,N_19382,N_18487);
and U24713 (N_24713,N_16189,N_15617);
and U24714 (N_24714,N_17356,N_17691);
and U24715 (N_24715,N_15495,N_17053);
nor U24716 (N_24716,N_18056,N_18617);
nor U24717 (N_24717,N_18560,N_16180);
nor U24718 (N_24718,N_18433,N_17496);
nor U24719 (N_24719,N_19873,N_15642);
and U24720 (N_24720,N_16044,N_16273);
and U24721 (N_24721,N_16767,N_15570);
and U24722 (N_24722,N_16076,N_19715);
xor U24723 (N_24723,N_18969,N_17047);
or U24724 (N_24724,N_17864,N_18241);
or U24725 (N_24725,N_18304,N_19967);
and U24726 (N_24726,N_18968,N_17669);
nor U24727 (N_24727,N_15555,N_15309);
or U24728 (N_24728,N_16523,N_15277);
xor U24729 (N_24729,N_17776,N_16975);
and U24730 (N_24730,N_15975,N_16536);
nand U24731 (N_24731,N_16095,N_19879);
and U24732 (N_24732,N_18015,N_19350);
nand U24733 (N_24733,N_17827,N_17666);
xor U24734 (N_24734,N_18023,N_18142);
nor U24735 (N_24735,N_16404,N_19080);
and U24736 (N_24736,N_19253,N_19379);
and U24737 (N_24737,N_18419,N_18356);
and U24738 (N_24738,N_15652,N_17629);
nor U24739 (N_24739,N_18093,N_19558);
and U24740 (N_24740,N_15559,N_15161);
xnor U24741 (N_24741,N_15007,N_16221);
nor U24742 (N_24742,N_17786,N_19111);
nor U24743 (N_24743,N_16956,N_19547);
and U24744 (N_24744,N_19606,N_19601);
or U24745 (N_24745,N_15494,N_16380);
and U24746 (N_24746,N_15049,N_15773);
nand U24747 (N_24747,N_15433,N_19815);
and U24748 (N_24748,N_18996,N_18878);
nor U24749 (N_24749,N_15335,N_15851);
or U24750 (N_24750,N_15710,N_18544);
nor U24751 (N_24751,N_16131,N_17007);
nor U24752 (N_24752,N_17131,N_18534);
and U24753 (N_24753,N_17031,N_16182);
and U24754 (N_24754,N_18443,N_15275);
and U24755 (N_24755,N_16758,N_16916);
and U24756 (N_24756,N_17828,N_15138);
nand U24757 (N_24757,N_16729,N_17668);
nand U24758 (N_24758,N_19084,N_16802);
nand U24759 (N_24759,N_17032,N_19695);
and U24760 (N_24760,N_18169,N_19195);
nand U24761 (N_24761,N_16866,N_17854);
nand U24762 (N_24762,N_15467,N_19802);
nand U24763 (N_24763,N_19078,N_19851);
nand U24764 (N_24764,N_18144,N_16632);
nand U24765 (N_24765,N_17793,N_19324);
xor U24766 (N_24766,N_16111,N_18023);
nand U24767 (N_24767,N_18325,N_17428);
or U24768 (N_24768,N_15843,N_19284);
nand U24769 (N_24769,N_19147,N_16597);
or U24770 (N_24770,N_18127,N_16237);
and U24771 (N_24771,N_15029,N_17708);
nand U24772 (N_24772,N_15314,N_18215);
and U24773 (N_24773,N_16546,N_19348);
nor U24774 (N_24774,N_15052,N_18165);
nor U24775 (N_24775,N_19286,N_15632);
and U24776 (N_24776,N_15285,N_18570);
nand U24777 (N_24777,N_15863,N_16145);
xnor U24778 (N_24778,N_16236,N_18694);
and U24779 (N_24779,N_15306,N_16782);
xnor U24780 (N_24780,N_15641,N_15448);
and U24781 (N_24781,N_15985,N_15845);
and U24782 (N_24782,N_19311,N_17871);
and U24783 (N_24783,N_19749,N_16476);
nand U24784 (N_24784,N_17807,N_15403);
or U24785 (N_24785,N_19790,N_17023);
or U24786 (N_24786,N_16760,N_17076);
nand U24787 (N_24787,N_17296,N_15313);
or U24788 (N_24788,N_19864,N_19845);
nand U24789 (N_24789,N_17676,N_17527);
and U24790 (N_24790,N_16571,N_16587);
nand U24791 (N_24791,N_16942,N_15276);
nor U24792 (N_24792,N_19064,N_19289);
nor U24793 (N_24793,N_15858,N_17659);
or U24794 (N_24794,N_16529,N_16523);
nor U24795 (N_24795,N_15755,N_15884);
or U24796 (N_24796,N_18884,N_18915);
or U24797 (N_24797,N_18405,N_16227);
and U24798 (N_24798,N_16295,N_16990);
and U24799 (N_24799,N_16856,N_18606);
or U24800 (N_24800,N_17410,N_15341);
xor U24801 (N_24801,N_19127,N_17439);
nor U24802 (N_24802,N_19777,N_16606);
xnor U24803 (N_24803,N_17889,N_15413);
nor U24804 (N_24804,N_18874,N_17583);
nand U24805 (N_24805,N_19462,N_19968);
xnor U24806 (N_24806,N_18882,N_19944);
or U24807 (N_24807,N_16756,N_19409);
nor U24808 (N_24808,N_15146,N_19730);
nand U24809 (N_24809,N_15110,N_17069);
or U24810 (N_24810,N_19429,N_15738);
nor U24811 (N_24811,N_16458,N_16196);
or U24812 (N_24812,N_15436,N_17188);
and U24813 (N_24813,N_15591,N_18605);
nand U24814 (N_24814,N_16149,N_15460);
nand U24815 (N_24815,N_18795,N_16116);
nand U24816 (N_24816,N_16995,N_19743);
and U24817 (N_24817,N_19139,N_16132);
nand U24818 (N_24818,N_15603,N_17797);
nand U24819 (N_24819,N_17955,N_15714);
nand U24820 (N_24820,N_15024,N_17419);
and U24821 (N_24821,N_15233,N_18765);
xnor U24822 (N_24822,N_17954,N_16770);
nand U24823 (N_24823,N_19493,N_15140);
nor U24824 (N_24824,N_17996,N_17420);
or U24825 (N_24825,N_19169,N_17452);
and U24826 (N_24826,N_17829,N_19411);
or U24827 (N_24827,N_17157,N_17416);
or U24828 (N_24828,N_15704,N_18278);
and U24829 (N_24829,N_17704,N_16148);
nor U24830 (N_24830,N_17182,N_15629);
nand U24831 (N_24831,N_17636,N_16790);
nor U24832 (N_24832,N_19887,N_19757);
or U24833 (N_24833,N_18158,N_19938);
and U24834 (N_24834,N_19614,N_19459);
nand U24835 (N_24835,N_15908,N_15246);
nor U24836 (N_24836,N_19150,N_17005);
and U24837 (N_24837,N_16375,N_19220);
nand U24838 (N_24838,N_19878,N_17744);
or U24839 (N_24839,N_17443,N_19804);
and U24840 (N_24840,N_18012,N_18794);
nand U24841 (N_24841,N_19341,N_16085);
nand U24842 (N_24842,N_17352,N_18559);
or U24843 (N_24843,N_16036,N_17500);
or U24844 (N_24844,N_15473,N_18565);
nor U24845 (N_24845,N_17186,N_17371);
xor U24846 (N_24846,N_15832,N_15451);
nor U24847 (N_24847,N_18247,N_15960);
nand U24848 (N_24848,N_18060,N_19320);
nor U24849 (N_24849,N_19371,N_16039);
nor U24850 (N_24850,N_16537,N_16329);
or U24851 (N_24851,N_18318,N_15952);
nand U24852 (N_24852,N_18584,N_18316);
nor U24853 (N_24853,N_19507,N_19413);
or U24854 (N_24854,N_18417,N_16760);
nand U24855 (N_24855,N_15378,N_16090);
nor U24856 (N_24856,N_19593,N_16856);
and U24857 (N_24857,N_17419,N_19365);
or U24858 (N_24858,N_18714,N_15964);
nand U24859 (N_24859,N_16321,N_19370);
or U24860 (N_24860,N_18280,N_15378);
and U24861 (N_24861,N_16055,N_19097);
or U24862 (N_24862,N_16313,N_16140);
xor U24863 (N_24863,N_15037,N_17059);
nand U24864 (N_24864,N_18450,N_15831);
nand U24865 (N_24865,N_18435,N_18246);
xnor U24866 (N_24866,N_19485,N_17415);
and U24867 (N_24867,N_19909,N_19933);
nand U24868 (N_24868,N_15916,N_19912);
nand U24869 (N_24869,N_16974,N_15921);
nand U24870 (N_24870,N_17722,N_19978);
or U24871 (N_24871,N_18137,N_15436);
nand U24872 (N_24872,N_19994,N_19018);
nor U24873 (N_24873,N_18799,N_18002);
nand U24874 (N_24874,N_17257,N_16484);
nor U24875 (N_24875,N_18040,N_16901);
nor U24876 (N_24876,N_18049,N_16171);
and U24877 (N_24877,N_15955,N_19056);
and U24878 (N_24878,N_17528,N_16915);
and U24879 (N_24879,N_18210,N_15121);
nand U24880 (N_24880,N_19258,N_17431);
nand U24881 (N_24881,N_16295,N_16455);
and U24882 (N_24882,N_17256,N_16398);
xor U24883 (N_24883,N_16975,N_19247);
and U24884 (N_24884,N_17530,N_19188);
nor U24885 (N_24885,N_17915,N_18581);
and U24886 (N_24886,N_16495,N_15137);
or U24887 (N_24887,N_16383,N_19354);
and U24888 (N_24888,N_18969,N_19547);
nor U24889 (N_24889,N_15820,N_16671);
or U24890 (N_24890,N_15397,N_19455);
and U24891 (N_24891,N_16528,N_17321);
nand U24892 (N_24892,N_18820,N_17206);
and U24893 (N_24893,N_19087,N_17274);
nand U24894 (N_24894,N_17650,N_15937);
nand U24895 (N_24895,N_17849,N_19459);
nor U24896 (N_24896,N_19976,N_17866);
nor U24897 (N_24897,N_15613,N_18120);
nor U24898 (N_24898,N_16104,N_18314);
and U24899 (N_24899,N_17294,N_15312);
nor U24900 (N_24900,N_17624,N_18636);
nand U24901 (N_24901,N_16504,N_19554);
nor U24902 (N_24902,N_15833,N_15418);
nor U24903 (N_24903,N_15070,N_15783);
or U24904 (N_24904,N_19539,N_16672);
and U24905 (N_24905,N_18742,N_18800);
nand U24906 (N_24906,N_17183,N_18481);
and U24907 (N_24907,N_16713,N_15559);
and U24908 (N_24908,N_17317,N_16325);
and U24909 (N_24909,N_17057,N_16300);
nor U24910 (N_24910,N_18647,N_16505);
and U24911 (N_24911,N_16346,N_19578);
or U24912 (N_24912,N_16591,N_17369);
and U24913 (N_24913,N_19519,N_18802);
nor U24914 (N_24914,N_17277,N_19610);
or U24915 (N_24915,N_16120,N_18295);
or U24916 (N_24916,N_17658,N_19025);
nor U24917 (N_24917,N_19041,N_16490);
or U24918 (N_24918,N_15270,N_18766);
nand U24919 (N_24919,N_18630,N_17805);
nor U24920 (N_24920,N_19798,N_17115);
or U24921 (N_24921,N_17989,N_18895);
nor U24922 (N_24922,N_19767,N_17613);
or U24923 (N_24923,N_18869,N_18372);
nand U24924 (N_24924,N_19180,N_18251);
or U24925 (N_24925,N_18340,N_18120);
or U24926 (N_24926,N_16286,N_15019);
or U24927 (N_24927,N_18258,N_16744);
nor U24928 (N_24928,N_15039,N_16163);
nor U24929 (N_24929,N_16132,N_18818);
and U24930 (N_24930,N_18483,N_17316);
and U24931 (N_24931,N_18563,N_15696);
or U24932 (N_24932,N_19495,N_16059);
and U24933 (N_24933,N_15780,N_17744);
nor U24934 (N_24934,N_18527,N_18585);
nor U24935 (N_24935,N_19064,N_16616);
xor U24936 (N_24936,N_19353,N_17741);
or U24937 (N_24937,N_18484,N_15735);
or U24938 (N_24938,N_17257,N_17216);
nor U24939 (N_24939,N_18655,N_18150);
nand U24940 (N_24940,N_16558,N_16957);
xor U24941 (N_24941,N_15228,N_18426);
and U24942 (N_24942,N_15025,N_17102);
or U24943 (N_24943,N_19257,N_18024);
and U24944 (N_24944,N_17349,N_15927);
nand U24945 (N_24945,N_15615,N_17712);
nor U24946 (N_24946,N_16171,N_17915);
nand U24947 (N_24947,N_18606,N_19786);
nor U24948 (N_24948,N_15072,N_17783);
nor U24949 (N_24949,N_17391,N_19722);
or U24950 (N_24950,N_19146,N_16477);
nand U24951 (N_24951,N_18655,N_16944);
and U24952 (N_24952,N_19751,N_17542);
nor U24953 (N_24953,N_16888,N_16798);
xnor U24954 (N_24954,N_18177,N_19050);
nor U24955 (N_24955,N_16359,N_19976);
nand U24956 (N_24956,N_18599,N_16488);
xnor U24957 (N_24957,N_17555,N_19287);
nor U24958 (N_24958,N_17839,N_16454);
nand U24959 (N_24959,N_15853,N_17689);
nand U24960 (N_24960,N_16519,N_18133);
nor U24961 (N_24961,N_16129,N_17516);
nor U24962 (N_24962,N_17120,N_17386);
nor U24963 (N_24963,N_18181,N_16483);
nor U24964 (N_24964,N_19060,N_17332);
and U24965 (N_24965,N_16593,N_19142);
and U24966 (N_24966,N_17949,N_18801);
xor U24967 (N_24967,N_19358,N_18423);
or U24968 (N_24968,N_19477,N_18930);
nand U24969 (N_24969,N_19289,N_19641);
nand U24970 (N_24970,N_18695,N_15127);
and U24971 (N_24971,N_15166,N_18703);
nand U24972 (N_24972,N_16967,N_15279);
nand U24973 (N_24973,N_17753,N_18883);
nor U24974 (N_24974,N_17978,N_19154);
nor U24975 (N_24975,N_17074,N_19263);
and U24976 (N_24976,N_19815,N_17056);
nand U24977 (N_24977,N_15153,N_17165);
nand U24978 (N_24978,N_15493,N_17787);
nand U24979 (N_24979,N_18492,N_19011);
nor U24980 (N_24980,N_18785,N_18307);
or U24981 (N_24981,N_18176,N_17344);
xnor U24982 (N_24982,N_16748,N_15416);
or U24983 (N_24983,N_17561,N_16458);
and U24984 (N_24984,N_17886,N_17922);
nor U24985 (N_24985,N_19097,N_15116);
nand U24986 (N_24986,N_16598,N_16078);
nor U24987 (N_24987,N_18261,N_18295);
and U24988 (N_24988,N_17470,N_19163);
xor U24989 (N_24989,N_16701,N_15455);
or U24990 (N_24990,N_19801,N_17407);
nor U24991 (N_24991,N_16033,N_18701);
nor U24992 (N_24992,N_19186,N_18972);
nand U24993 (N_24993,N_18244,N_17582);
nand U24994 (N_24994,N_19948,N_19083);
nand U24995 (N_24995,N_17399,N_15311);
xnor U24996 (N_24996,N_17508,N_18784);
or U24997 (N_24997,N_19074,N_19291);
or U24998 (N_24998,N_15978,N_19558);
nor U24999 (N_24999,N_19270,N_17009);
nor U25000 (N_25000,N_22645,N_20490);
nor U25001 (N_25001,N_21240,N_23647);
nor U25002 (N_25002,N_24856,N_22691);
or U25003 (N_25003,N_24277,N_22769);
and U25004 (N_25004,N_22113,N_22754);
or U25005 (N_25005,N_22631,N_22501);
nor U25006 (N_25006,N_22097,N_21399);
nand U25007 (N_25007,N_24103,N_20969);
nor U25008 (N_25008,N_20405,N_24032);
nor U25009 (N_25009,N_20571,N_23805);
nor U25010 (N_25010,N_20799,N_23782);
and U25011 (N_25011,N_20046,N_23347);
and U25012 (N_25012,N_22298,N_22863);
nand U25013 (N_25013,N_21865,N_24173);
and U25014 (N_25014,N_24185,N_24026);
or U25015 (N_25015,N_24944,N_20999);
or U25016 (N_25016,N_24101,N_21824);
and U25017 (N_25017,N_20621,N_20473);
and U25018 (N_25018,N_20005,N_20390);
or U25019 (N_25019,N_23915,N_23322);
or U25020 (N_25020,N_22433,N_21985);
and U25021 (N_25021,N_21683,N_20185);
and U25022 (N_25022,N_20223,N_23662);
nor U25023 (N_25023,N_21339,N_22713);
or U25024 (N_25024,N_23914,N_21484);
nor U25025 (N_25025,N_22219,N_23889);
nor U25026 (N_25026,N_23818,N_21634);
nand U25027 (N_25027,N_21598,N_21546);
xnor U25028 (N_25028,N_23502,N_21156);
and U25029 (N_25029,N_23195,N_24138);
xnor U25030 (N_25030,N_23918,N_22104);
nor U25031 (N_25031,N_22218,N_20182);
nand U25032 (N_25032,N_21224,N_21489);
and U25033 (N_25033,N_23724,N_20441);
nand U25034 (N_25034,N_21932,N_24407);
and U25035 (N_25035,N_20610,N_21565);
nor U25036 (N_25036,N_24079,N_23944);
or U25037 (N_25037,N_22276,N_21609);
nand U25038 (N_25038,N_23119,N_23768);
or U25039 (N_25039,N_23019,N_24510);
nand U25040 (N_25040,N_23552,N_20931);
and U25041 (N_25041,N_23631,N_24442);
xnor U25042 (N_25042,N_20471,N_24557);
nor U25043 (N_25043,N_23152,N_21508);
or U25044 (N_25044,N_20312,N_21409);
and U25045 (N_25045,N_24848,N_21052);
nor U25046 (N_25046,N_21148,N_22616);
and U25047 (N_25047,N_21806,N_22838);
or U25048 (N_25048,N_20128,N_24934);
nor U25049 (N_25049,N_23381,N_24445);
nor U25050 (N_25050,N_20144,N_22361);
and U25051 (N_25051,N_22239,N_22170);
nor U25052 (N_25052,N_23190,N_20674);
nand U25053 (N_25053,N_23695,N_23710);
nand U25054 (N_25054,N_21811,N_20180);
or U25055 (N_25055,N_22382,N_24212);
nand U25056 (N_25056,N_21213,N_22423);
nor U25057 (N_25057,N_21757,N_23830);
or U25058 (N_25058,N_22799,N_21397);
xor U25059 (N_25059,N_20380,N_23547);
xnor U25060 (N_25060,N_24807,N_20825);
nand U25061 (N_25061,N_21365,N_23900);
nand U25062 (N_25062,N_20332,N_24721);
xnor U25063 (N_25063,N_21143,N_23241);
nor U25064 (N_25064,N_22485,N_22374);
xnor U25065 (N_25065,N_20749,N_20083);
or U25066 (N_25066,N_21228,N_20225);
nand U25067 (N_25067,N_21058,N_21694);
xnor U25068 (N_25068,N_20634,N_22269);
and U25069 (N_25069,N_24907,N_23472);
and U25070 (N_25070,N_23635,N_22355);
nor U25071 (N_25071,N_22638,N_23079);
and U25072 (N_25072,N_23581,N_23361);
nor U25073 (N_25073,N_21647,N_23038);
and U25074 (N_25074,N_24868,N_24652);
or U25075 (N_25075,N_21251,N_21466);
nand U25076 (N_25076,N_23794,N_24544);
nand U25077 (N_25077,N_24403,N_24877);
or U25078 (N_25078,N_24792,N_23941);
and U25079 (N_25079,N_24260,N_23184);
nand U25080 (N_25080,N_20461,N_24859);
or U25081 (N_25081,N_20142,N_20813);
and U25082 (N_25082,N_24874,N_23682);
nor U25083 (N_25083,N_21208,N_22100);
or U25084 (N_25084,N_23855,N_23133);
nand U25085 (N_25085,N_20566,N_24521);
nor U25086 (N_25086,N_21418,N_22749);
or U25087 (N_25087,N_21169,N_23189);
nor U25088 (N_25088,N_22917,N_22342);
xor U25089 (N_25089,N_20288,N_22284);
and U25090 (N_25090,N_21073,N_20482);
nand U25091 (N_25091,N_22384,N_22392);
xor U25092 (N_25092,N_24554,N_23793);
nand U25093 (N_25093,N_23601,N_20488);
nand U25094 (N_25094,N_22233,N_23899);
or U25095 (N_25095,N_20311,N_23626);
or U25096 (N_25096,N_21098,N_24064);
nand U25097 (N_25097,N_20994,N_24775);
nand U25098 (N_25098,N_21205,N_22800);
and U25099 (N_25099,N_23965,N_23265);
xor U25100 (N_25100,N_23122,N_24805);
or U25101 (N_25101,N_22983,N_20743);
xor U25102 (N_25102,N_20370,N_20844);
nand U25103 (N_25103,N_22312,N_24146);
nor U25104 (N_25104,N_20788,N_22866);
or U25105 (N_25105,N_22425,N_23978);
or U25106 (N_25106,N_24106,N_20369);
nand U25107 (N_25107,N_23962,N_22347);
xnor U25108 (N_25108,N_22172,N_21914);
nor U25109 (N_25109,N_24712,N_24120);
or U25110 (N_25110,N_24595,N_23881);
and U25111 (N_25111,N_21117,N_24522);
nand U25112 (N_25112,N_20885,N_24741);
and U25113 (N_25113,N_23450,N_22770);
nand U25114 (N_25114,N_22292,N_22237);
or U25115 (N_25115,N_21087,N_24958);
nand U25116 (N_25116,N_23592,N_22553);
xnor U25117 (N_25117,N_21133,N_22011);
or U25118 (N_25118,N_24147,N_21509);
nor U25119 (N_25119,N_20608,N_22280);
or U25120 (N_25120,N_24576,N_23104);
nor U25121 (N_25121,N_20345,N_21572);
or U25122 (N_25122,N_22459,N_20734);
or U25123 (N_25123,N_20922,N_24885);
nand U25124 (N_25124,N_20156,N_20964);
nand U25125 (N_25125,N_24084,N_20555);
nor U25126 (N_25126,N_22061,N_23884);
nor U25127 (N_25127,N_22891,N_20572);
or U25128 (N_25128,N_22614,N_21235);
nand U25129 (N_25129,N_23760,N_20830);
nor U25130 (N_25130,N_20248,N_23051);
and U25131 (N_25131,N_22213,N_24936);
or U25132 (N_25132,N_20918,N_21522);
nand U25133 (N_25133,N_24745,N_21836);
or U25134 (N_25134,N_23239,N_22108);
or U25135 (N_25135,N_23575,N_22448);
and U25136 (N_25136,N_22796,N_21167);
nor U25137 (N_25137,N_22340,N_21216);
nor U25138 (N_25138,N_22144,N_21407);
xnor U25139 (N_25139,N_24425,N_24221);
and U25140 (N_25140,N_22181,N_23542);
or U25141 (N_25141,N_22438,N_21255);
and U25142 (N_25142,N_23062,N_23233);
nand U25143 (N_25143,N_24402,N_22489);
xnor U25144 (N_25144,N_22856,N_20512);
xnor U25145 (N_25145,N_20138,N_23072);
nor U25146 (N_25146,N_21613,N_23728);
and U25147 (N_25147,N_21866,N_24399);
or U25148 (N_25148,N_22937,N_24621);
or U25149 (N_25149,N_22165,N_23549);
or U25150 (N_25150,N_23288,N_22212);
nor U25151 (N_25151,N_23652,N_24112);
or U25152 (N_25152,N_23819,N_24482);
nor U25153 (N_25153,N_24584,N_24426);
or U25154 (N_25154,N_21280,N_24520);
and U25155 (N_25155,N_23888,N_22632);
xor U25156 (N_25156,N_24016,N_23012);
nand U25157 (N_25157,N_24880,N_21467);
or U25158 (N_25158,N_21942,N_22069);
and U25159 (N_25159,N_21913,N_21666);
nand U25160 (N_25160,N_23902,N_20363);
or U25161 (N_25161,N_23734,N_24606);
xnor U25162 (N_25162,N_22506,N_20262);
nand U25163 (N_25163,N_24704,N_23524);
nand U25164 (N_25164,N_21154,N_23546);
or U25165 (N_25165,N_22319,N_20597);
nor U25166 (N_25166,N_20212,N_22858);
and U25167 (N_25167,N_23188,N_22888);
nand U25168 (N_25168,N_23130,N_24428);
and U25169 (N_25169,N_23317,N_23298);
and U25170 (N_25170,N_22180,N_23800);
or U25171 (N_25171,N_21031,N_23833);
or U25172 (N_25172,N_20333,N_20159);
nor U25173 (N_25173,N_23954,N_23314);
or U25174 (N_25174,N_22153,N_22791);
and U25175 (N_25175,N_21144,N_22855);
nor U25176 (N_25176,N_21193,N_22872);
or U25177 (N_25177,N_21475,N_22998);
or U25178 (N_25178,N_22480,N_21113);
and U25179 (N_25179,N_23931,N_22018);
nand U25180 (N_25180,N_21338,N_21881);
or U25181 (N_25181,N_21192,N_23209);
nand U25182 (N_25182,N_23260,N_23453);
nor U25183 (N_25183,N_22474,N_22297);
nand U25184 (N_25184,N_20792,N_23413);
nand U25185 (N_25185,N_22341,N_21272);
or U25186 (N_25186,N_21402,N_22223);
nand U25187 (N_25187,N_20705,N_23766);
and U25188 (N_25188,N_24686,N_23562);
xnor U25189 (N_25189,N_23625,N_23779);
or U25190 (N_25190,N_24396,N_20733);
or U25191 (N_25191,N_24730,N_21783);
nor U25192 (N_25192,N_24242,N_21054);
nor U25193 (N_25193,N_21422,N_21009);
nand U25194 (N_25194,N_22941,N_22934);
nor U25195 (N_25195,N_23258,N_21555);
and U25196 (N_25196,N_21545,N_23333);
nor U25197 (N_25197,N_23909,N_22593);
xor U25198 (N_25198,N_23560,N_21086);
xnor U25199 (N_25199,N_20872,N_21254);
xor U25200 (N_25200,N_22327,N_23481);
nor U25201 (N_25201,N_24314,N_23840);
nand U25202 (N_25202,N_24136,N_22129);
xor U25203 (N_25203,N_23252,N_23335);
and U25204 (N_25204,N_23667,N_21763);
and U25205 (N_25205,N_21896,N_20320);
nor U25206 (N_25206,N_21525,N_21573);
or U25207 (N_25207,N_22288,N_20754);
or U25208 (N_25208,N_24491,N_22469);
and U25209 (N_25209,N_23434,N_23423);
or U25210 (N_25210,N_24200,N_21848);
and U25211 (N_25211,N_23616,N_21905);
or U25212 (N_25212,N_21071,N_24224);
and U25213 (N_25213,N_20874,N_22668);
and U25214 (N_25214,N_21306,N_23674);
and U25215 (N_25215,N_21158,N_21954);
nor U25216 (N_25216,N_23798,N_22383);
nor U25217 (N_25217,N_21882,N_23593);
nand U25218 (N_25218,N_22176,N_23221);
or U25219 (N_25219,N_20219,N_20745);
or U25220 (N_25220,N_24273,N_23679);
nor U25221 (N_25221,N_20949,N_23113);
xor U25222 (N_25222,N_23653,N_21273);
or U25223 (N_25223,N_22294,N_21206);
nor U25224 (N_25224,N_24619,N_20859);
nand U25225 (N_25225,N_22889,N_23222);
or U25226 (N_25226,N_23808,N_20140);
or U25227 (N_25227,N_22993,N_24793);
xor U25228 (N_25228,N_23214,N_24981);
nand U25229 (N_25229,N_23493,N_24891);
and U25230 (N_25230,N_21926,N_21602);
nor U25231 (N_25231,N_20860,N_24896);
nand U25232 (N_25232,N_23420,N_24168);
nor U25233 (N_25233,N_21720,N_24909);
nand U25234 (N_25234,N_23429,N_23312);
xor U25235 (N_25235,N_21662,N_21685);
nor U25236 (N_25236,N_20588,N_21129);
or U25237 (N_25237,N_24693,N_20015);
or U25238 (N_25238,N_23082,N_24542);
nor U25239 (N_25239,N_23203,N_21064);
or U25240 (N_25240,N_22461,N_20064);
or U25241 (N_25241,N_23947,N_23256);
and U25242 (N_25242,N_21699,N_21379);
or U25243 (N_25243,N_21390,N_23530);
xor U25244 (N_25244,N_24455,N_20116);
nand U25245 (N_25245,N_24748,N_24561);
nand U25246 (N_25246,N_20952,N_24598);
and U25247 (N_25247,N_23811,N_21155);
or U25248 (N_25248,N_23860,N_23338);
nor U25249 (N_25249,N_21004,N_24247);
or U25250 (N_25250,N_20718,N_20656);
nor U25251 (N_25251,N_24430,N_21210);
nor U25252 (N_25252,N_23852,N_24747);
nand U25253 (N_25253,N_24804,N_21925);
nand U25254 (N_25254,N_24568,N_21289);
xor U25255 (N_25255,N_24135,N_22723);
nand U25256 (N_25256,N_22894,N_20750);
nand U25257 (N_25257,N_24148,N_20677);
xnor U25258 (N_25258,N_23357,N_23398);
and U25259 (N_25259,N_24964,N_22070);
and U25260 (N_25260,N_23110,N_21577);
or U25261 (N_25261,N_24263,N_24073);
nor U25262 (N_25262,N_21329,N_20496);
nor U25263 (N_25263,N_21775,N_24011);
and U25264 (N_25264,N_22596,N_20030);
and U25265 (N_25265,N_22503,N_23358);
and U25266 (N_25266,N_22162,N_20125);
or U25267 (N_25267,N_24875,N_24065);
xor U25268 (N_25268,N_22865,N_23966);
nor U25269 (N_25269,N_22844,N_21533);
nand U25270 (N_25270,N_22360,N_20620);
or U25271 (N_25271,N_24341,N_24955);
nor U25272 (N_25272,N_20661,N_24512);
or U25273 (N_25273,N_21060,N_20547);
xnor U25274 (N_25274,N_21336,N_20599);
and U25275 (N_25275,N_23092,N_21599);
and U25276 (N_25276,N_24800,N_21414);
nor U25277 (N_25277,N_22078,N_22756);
nand U25278 (N_25278,N_23248,N_20829);
nor U25279 (N_25279,N_23597,N_24657);
and U25280 (N_25280,N_24708,N_20143);
xor U25281 (N_25281,N_24631,N_24329);
xor U25282 (N_25282,N_24272,N_22063);
xor U25283 (N_25283,N_24029,N_23293);
or U25284 (N_25284,N_24806,N_20044);
nand U25285 (N_25285,N_23689,N_20777);
nand U25286 (N_25286,N_20124,N_23269);
nand U25287 (N_25287,N_21604,N_21966);
nor U25288 (N_25288,N_22258,N_21716);
or U25289 (N_25289,N_22470,N_20183);
or U25290 (N_25290,N_24849,N_23956);
and U25291 (N_25291,N_22546,N_21723);
or U25292 (N_25292,N_20462,N_24753);
or U25293 (N_25293,N_22033,N_21114);
and U25294 (N_25294,N_23864,N_23587);
nor U25295 (N_25295,N_24304,N_21945);
nor U25296 (N_25296,N_23834,N_23661);
nand U25297 (N_25297,N_21356,N_24483);
and U25298 (N_25298,N_21179,N_24563);
nor U25299 (N_25299,N_22516,N_20973);
or U25300 (N_25300,N_24600,N_20649);
nor U25301 (N_25301,N_20652,N_20385);
nor U25302 (N_25302,N_20020,N_22378);
nor U25303 (N_25303,N_21267,N_22232);
nor U25304 (N_25304,N_23250,N_24904);
xnor U25305 (N_25305,N_24646,N_21698);
nand U25306 (N_25306,N_23576,N_24344);
and U25307 (N_25307,N_21752,N_20121);
nand U25308 (N_25308,N_20321,N_23080);
or U25309 (N_25309,N_20475,N_21534);
nor U25310 (N_25310,N_20536,N_21519);
or U25311 (N_25311,N_22709,N_21068);
xnor U25312 (N_25312,N_20856,N_22807);
nor U25313 (N_25313,N_21851,N_24833);
nand U25314 (N_25314,N_24181,N_21184);
or U25315 (N_25315,N_20072,N_21987);
and U25316 (N_25316,N_22116,N_21044);
nand U25317 (N_25317,N_20575,N_21963);
nor U25318 (N_25318,N_22651,N_24627);
nand U25319 (N_25319,N_22529,N_24530);
or U25320 (N_25320,N_20979,N_22436);
nand U25321 (N_25321,N_22817,N_23162);
and U25322 (N_25322,N_22979,N_21819);
nand U25323 (N_25323,N_20346,N_23433);
nor U25324 (N_25324,N_23046,N_24952);
xor U25325 (N_25325,N_21130,N_20455);
nor U25326 (N_25326,N_24443,N_22608);
nor U25327 (N_25327,N_22710,N_24256);
or U25328 (N_25328,N_24691,N_20631);
or U25329 (N_25329,N_20444,N_23309);
or U25330 (N_25330,N_24565,N_22833);
and U25331 (N_25331,N_21258,N_22085);
or U25332 (N_25332,N_20006,N_21436);
nor U25333 (N_25333,N_20474,N_24917);
nor U25334 (N_25334,N_22882,N_23343);
or U25335 (N_25335,N_20676,N_23109);
or U25336 (N_25336,N_22657,N_23174);
and U25337 (N_25337,N_20974,N_20366);
nand U25338 (N_25338,N_22569,N_24743);
nand U25339 (N_25339,N_22274,N_24054);
nand U25340 (N_25340,N_21047,N_22444);
nor U25341 (N_25341,N_24682,N_20200);
or U25342 (N_25342,N_24332,N_20744);
or U25343 (N_25343,N_20177,N_20360);
nand U25344 (N_25344,N_23255,N_22938);
nor U25345 (N_25345,N_20145,N_21089);
nor U25346 (N_25346,N_21299,N_23476);
and U25347 (N_25347,N_24170,N_20246);
or U25348 (N_25348,N_24724,N_20304);
nor U25349 (N_25349,N_22059,N_23839);
and U25350 (N_25350,N_20472,N_22183);
and U25351 (N_25351,N_23972,N_24469);
nor U25352 (N_25352,N_21287,N_21998);
nand U25353 (N_25353,N_21850,N_21642);
and U25354 (N_25354,N_24191,N_24262);
or U25355 (N_25355,N_23197,N_20950);
nand U25356 (N_25356,N_24988,N_21878);
and U25357 (N_25357,N_21332,N_22602);
nand U25358 (N_25358,N_23712,N_24668);
nor U25359 (N_25359,N_22397,N_23973);
or U25360 (N_25360,N_24725,N_23693);
nor U25361 (N_25361,N_20741,N_23348);
nor U25362 (N_25362,N_22262,N_22279);
nor U25363 (N_25363,N_20167,N_20569);
nand U25364 (N_25364,N_24642,N_22377);
or U25365 (N_25365,N_24369,N_22661);
xnor U25366 (N_25366,N_23711,N_23611);
and U25367 (N_25367,N_21428,N_20076);
nand U25368 (N_25368,N_20197,N_24705);
and U25369 (N_25369,N_23351,N_22561);
nand U25370 (N_25370,N_24791,N_20139);
nand U25371 (N_25371,N_23690,N_22247);
nor U25372 (N_25372,N_20094,N_20134);
nand U25373 (N_25373,N_22605,N_22852);
nor U25374 (N_25374,N_20552,N_20172);
and U25375 (N_25375,N_20570,N_23128);
xnor U25376 (N_25376,N_20663,N_24549);
nor U25377 (N_25377,N_20232,N_22477);
and U25378 (N_25378,N_20340,N_20082);
and U25379 (N_25379,N_23304,N_21246);
nor U25380 (N_25380,N_24843,N_21293);
xnor U25381 (N_25381,N_24149,N_23061);
xnor U25382 (N_25382,N_24995,N_20255);
or U25383 (N_25383,N_21371,N_20839);
and U25384 (N_25384,N_24975,N_22483);
or U25385 (N_25385,N_23186,N_24673);
and U25386 (N_25386,N_21984,N_23218);
or U25387 (N_25387,N_22222,N_23262);
and U25388 (N_25388,N_24845,N_20236);
nor U25389 (N_25389,N_20237,N_24354);
nand U25390 (N_25390,N_20221,N_20654);
nor U25391 (N_25391,N_22096,N_23791);
nor U25392 (N_25392,N_24312,N_22492);
and U25393 (N_25393,N_22025,N_22389);
and U25394 (N_25394,N_20896,N_20239);
or U25395 (N_25395,N_23686,N_20836);
and U25396 (N_25396,N_20463,N_24915);
or U25397 (N_25397,N_22135,N_22495);
nor U25398 (N_25398,N_22077,N_22324);
and U25399 (N_25399,N_20001,N_22620);
nand U25400 (N_25400,N_21679,N_23028);
or U25401 (N_25401,N_21632,N_21396);
or U25402 (N_25402,N_20514,N_20268);
nor U25403 (N_25403,N_20178,N_23731);
or U25404 (N_25404,N_20504,N_23774);
nor U25405 (N_25405,N_22793,N_22350);
and U25406 (N_25406,N_21784,N_23564);
and U25407 (N_25407,N_20402,N_20506);
nand U25408 (N_25408,N_21075,N_20133);
nor U25409 (N_25409,N_24411,N_20722);
and U25410 (N_25410,N_23848,N_21768);
or U25411 (N_25411,N_22160,N_23844);
or U25412 (N_25412,N_21550,N_22060);
and U25413 (N_25413,N_23063,N_22512);
and U25414 (N_25414,N_23415,N_23105);
or U25415 (N_25415,N_21949,N_21145);
nor U25416 (N_25416,N_21080,N_23383);
or U25417 (N_25417,N_24470,N_23905);
and U25418 (N_25418,N_22745,N_21430);
nor U25419 (N_25419,N_23267,N_23571);
or U25420 (N_25420,N_22301,N_21105);
nor U25421 (N_25421,N_20598,N_20120);
xnor U25422 (N_25422,N_23360,N_24355);
and U25423 (N_25423,N_24220,N_21975);
nor U25424 (N_25424,N_24675,N_21808);
nand U25425 (N_25425,N_23488,N_24838);
nor U25426 (N_25426,N_24062,N_22246);
and U25427 (N_25427,N_21681,N_22446);
nor U25428 (N_25428,N_20645,N_22803);
and U25429 (N_25429,N_22066,N_24940);
and U25430 (N_25430,N_22974,N_20330);
nor U25431 (N_25431,N_23574,N_24339);
nor U25432 (N_25432,N_23446,N_24444);
nor U25433 (N_25433,N_24986,N_20841);
nor U25434 (N_25434,N_23173,N_23388);
nor U25435 (N_25435,N_21626,N_20748);
xor U25436 (N_25436,N_20034,N_22261);
xor U25437 (N_25437,N_23163,N_24816);
or U25438 (N_25438,N_24229,N_23949);
nand U25439 (N_25439,N_23595,N_21275);
nand U25440 (N_25440,N_23033,N_20119);
nand U25441 (N_25441,N_20410,N_21186);
and U25442 (N_25442,N_22878,N_23404);
nor U25443 (N_25443,N_21168,N_21579);
or U25444 (N_25444,N_22640,N_21199);
or U25445 (N_25445,N_21491,N_22772);
nand U25446 (N_25446,N_21278,N_20636);
nor U25447 (N_25447,N_23518,N_22747);
and U25448 (N_25448,N_21551,N_24882);
and U25449 (N_25449,N_21279,N_20938);
xnor U25450 (N_25450,N_20558,N_22435);
or U25451 (N_25451,N_21030,N_24920);
nand U25452 (N_25452,N_21753,N_23158);
nand U25453 (N_25453,N_24335,N_21459);
or U25454 (N_25454,N_24334,N_20935);
or U25455 (N_25455,N_22753,N_22410);
nor U25456 (N_25456,N_20227,N_22650);
nor U25457 (N_25457,N_21005,N_24254);
or U25458 (N_25458,N_22226,N_22551);
and U25459 (N_25459,N_22945,N_20553);
xnor U25460 (N_25460,N_22079,N_21857);
and U25461 (N_25461,N_24346,N_21868);
xnor U25462 (N_25462,N_22320,N_21268);
xnor U25463 (N_25463,N_21286,N_24954);
and U25464 (N_25464,N_21797,N_24033);
or U25465 (N_25465,N_24360,N_22789);
or U25466 (N_25466,N_20580,N_24143);
xor U25467 (N_25467,N_24299,N_22944);
and U25468 (N_25468,N_21476,N_24710);
or U25469 (N_25469,N_23193,N_24573);
or U25470 (N_25470,N_20240,N_22317);
nor U25471 (N_25471,N_24440,N_20493);
nand U25472 (N_25472,N_24685,N_20639);
nor U25473 (N_25473,N_24420,N_23192);
nand U25474 (N_25474,N_21479,N_22128);
nand U25475 (N_25475,N_21653,N_24830);
or U25476 (N_25476,N_22071,N_20155);
or U25477 (N_25477,N_23023,N_23268);
xnor U25478 (N_25478,N_24580,N_22766);
or U25479 (N_25479,N_22271,N_24773);
or U25480 (N_25480,N_21063,N_20694);
xnor U25481 (N_25481,N_22310,N_22131);
or U25482 (N_25482,N_23443,N_21944);
nor U25483 (N_25483,N_24860,N_23447);
nor U25484 (N_25484,N_22388,N_20698);
xor U25485 (N_25485,N_20202,N_24599);
or U25486 (N_25486,N_22566,N_24067);
nor U25487 (N_25487,N_24210,N_21712);
nand U25488 (N_25488,N_21357,N_20365);
xnor U25489 (N_25489,N_24236,N_22394);
or U25490 (N_25490,N_21084,N_24715);
and U25491 (N_25491,N_20800,N_20867);
nor U25492 (N_25492,N_24169,N_21081);
nand U25493 (N_25493,N_22671,N_21701);
nor U25494 (N_25494,N_21016,N_22193);
nand U25495 (N_25495,N_23098,N_20100);
and U25496 (N_25496,N_21842,N_23912);
nor U25497 (N_25497,N_23796,N_20446);
xor U25498 (N_25498,N_24572,N_20301);
nand U25499 (N_25499,N_22381,N_24189);
or U25500 (N_25500,N_21025,N_24723);
nand U25501 (N_25501,N_22267,N_24498);
and U25502 (N_25502,N_20768,N_21812);
and U25503 (N_25503,N_21673,N_24996);
or U25504 (N_25504,N_22748,N_24095);
nand U25505 (N_25505,N_21368,N_23814);
nor U25506 (N_25506,N_22065,N_23328);
xnor U25507 (N_25507,N_24553,N_21314);
nor U25508 (N_25508,N_23726,N_20175);
and U25509 (N_25509,N_22798,N_21474);
nor U25510 (N_25510,N_22903,N_20894);
xor U25511 (N_25511,N_24605,N_23910);
and U25512 (N_25512,N_24662,N_22430);
nand U25513 (N_25513,N_22613,N_22263);
xor U25514 (N_25514,N_24000,N_20003);
nor U25515 (N_25515,N_20525,N_23424);
nor U25516 (N_25516,N_22963,N_24384);
nand U25517 (N_25517,N_23648,N_24292);
nand U25518 (N_25518,N_22952,N_22041);
or U25519 (N_25519,N_22291,N_21628);
or U25520 (N_25520,N_21049,N_23005);
and U25521 (N_25521,N_20928,N_21022);
or U25522 (N_25522,N_22089,N_24091);
nand U25523 (N_25523,N_24731,N_21324);
nand U25524 (N_25524,N_23922,N_24234);
and U25525 (N_25525,N_20650,N_24233);
xnor U25526 (N_25526,N_22151,N_24861);
and U25527 (N_25527,N_23286,N_23789);
or U25528 (N_25528,N_22019,N_22904);
and U25529 (N_25529,N_21782,N_24979);
nand U25530 (N_25530,N_23134,N_23555);
nor U25531 (N_25531,N_20022,N_21302);
or U25532 (N_25532,N_21695,N_22149);
or U25533 (N_25533,N_22224,N_23874);
and U25534 (N_25534,N_23963,N_21469);
and U25535 (N_25535,N_20560,N_24752);
and U25536 (N_25536,N_22890,N_21636);
nor U25537 (N_25537,N_21420,N_23159);
nor U25538 (N_25538,N_23401,N_24388);
nor U25539 (N_25539,N_22850,N_23083);
xnor U25540 (N_25540,N_23350,N_20840);
or U25541 (N_25541,N_20616,N_21334);
nand U25542 (N_25542,N_24110,N_20398);
or U25543 (N_25543,N_21408,N_22035);
or U25544 (N_25544,N_24331,N_20888);
or U25545 (N_25545,N_20215,N_23979);
nand U25546 (N_25546,N_20282,N_21729);
and U25547 (N_25547,N_23906,N_24457);
nor U25548 (N_25548,N_21471,N_23125);
and U25549 (N_25549,N_23621,N_22848);
nand U25550 (N_25550,N_22414,N_24279);
or U25551 (N_25551,N_23890,N_21090);
and U25552 (N_25552,N_24495,N_24918);
nor U25553 (N_25553,N_23499,N_22623);
nor U25554 (N_25554,N_24467,N_20310);
nand U25555 (N_25555,N_22921,N_21814);
nor U25556 (N_25556,N_20089,N_21326);
nor U25557 (N_25557,N_21252,N_24130);
nor U25558 (N_25558,N_24528,N_24991);
nor U25559 (N_25559,N_22259,N_22510);
nand U25560 (N_25560,N_22765,N_22926);
nor U25561 (N_25561,N_22366,N_23753);
or U25562 (N_25562,N_24552,N_22680);
nand U25563 (N_25563,N_23373,N_21921);
nor U25564 (N_25564,N_21977,N_24265);
nor U25565 (N_25565,N_22426,N_21037);
or U25566 (N_25566,N_22139,N_23723);
nor U25567 (N_25567,N_23206,N_24985);
or U25568 (N_25568,N_21443,N_21523);
or U25569 (N_25569,N_23633,N_22992);
xnor U25570 (N_25570,N_23013,N_23067);
xor U25571 (N_25571,N_21520,N_21557);
or U25572 (N_25572,N_24007,N_23925);
and U25573 (N_25573,N_21751,N_22051);
nand U25574 (N_25574,N_20457,N_21686);
nand U25575 (N_25575,N_20880,N_22639);
nand U25576 (N_25576,N_22664,N_24799);
nor U25577 (N_25577,N_24362,N_21655);
nor U25578 (N_25578,N_20562,N_24921);
nand U25579 (N_25579,N_22622,N_23389);
nand U25580 (N_25580,N_21091,N_22244);
and U25581 (N_25581,N_23020,N_24754);
nand U25582 (N_25582,N_20152,N_20104);
xor U25583 (N_25583,N_23449,N_24374);
xnor U25584 (N_25584,N_20737,N_24161);
nand U25585 (N_25585,N_24379,N_23516);
or U25586 (N_25586,N_22462,N_22556);
or U25587 (N_25587,N_24156,N_20921);
nor U25588 (N_25588,N_21585,N_20900);
and U25589 (N_25589,N_24010,N_24577);
nor U25590 (N_25590,N_23435,N_22105);
or U25591 (N_25591,N_24121,N_21488);
nor U25592 (N_25592,N_21237,N_20438);
nand U25593 (N_25593,N_22346,N_22257);
nand U25594 (N_25594,N_20238,N_22666);
and U25595 (N_25595,N_22243,N_23330);
or U25596 (N_25596,N_20413,N_20662);
nand U25597 (N_25597,N_20218,N_20528);
xor U25598 (N_25598,N_23452,N_24543);
and U25599 (N_25599,N_20179,N_23714);
and U25600 (N_25600,N_21503,N_23971);
and U25601 (N_25601,N_23573,N_21664);
or U25602 (N_25602,N_23369,N_23319);
nand U25603 (N_25603,N_20584,N_20758);
or U25604 (N_25604,N_23980,N_22202);
and U25605 (N_25605,N_24583,N_20685);
nand U25606 (N_25606,N_22829,N_23820);
nand U25607 (N_25607,N_20554,N_20158);
nor U25608 (N_25608,N_24513,N_21317);
xor U25609 (N_25609,N_24041,N_23933);
and U25610 (N_25610,N_20804,N_24751);
nand U25611 (N_25611,N_24216,N_20926);
xor U25612 (N_25612,N_22467,N_21377);
nand U25613 (N_25613,N_23300,N_22764);
and U25614 (N_25614,N_24898,N_23074);
nand U25615 (N_25615,N_24591,N_20408);
nand U25616 (N_25616,N_23660,N_23836);
xor U25617 (N_25617,N_23213,N_20527);
nor U25618 (N_25618,N_22416,N_22635);
and U25619 (N_25619,N_22174,N_22603);
nor U25620 (N_25620,N_20068,N_21386);
and U25621 (N_25621,N_22665,N_20538);
nand U25622 (N_25622,N_22229,N_21162);
xnor U25623 (N_25623,N_21359,N_24968);
nor U25624 (N_25624,N_20546,N_21918);
nand U25625 (N_25625,N_20613,N_21319);
xnor U25626 (N_25626,N_24432,N_20932);
or U25627 (N_25627,N_23187,N_22456);
and U25628 (N_25628,N_22252,N_22812);
or U25629 (N_25629,N_21384,N_24894);
and U25630 (N_25630,N_20352,N_21959);
and U25631 (N_25631,N_23022,N_20923);
nand U25632 (N_25632,N_22082,N_21643);
and U25633 (N_25633,N_24261,N_24461);
nor U25634 (N_25634,N_20899,N_21660);
nand U25635 (N_25635,N_20087,N_24757);
or U25636 (N_25636,N_20978,N_24046);
or U25637 (N_25637,N_20765,N_24966);
and U25638 (N_25638,N_23039,N_24145);
or U25639 (N_25639,N_24177,N_23536);
or U25640 (N_25640,N_21810,N_20819);
or U25641 (N_25641,N_22695,N_23868);
nand U25642 (N_25642,N_21730,N_20298);
and U25643 (N_25643,N_21248,N_23111);
nor U25644 (N_25644,N_21126,N_24421);
nor U25645 (N_25645,N_20760,N_24307);
nor U25646 (N_25646,N_20803,N_20358);
nand U25647 (N_25647,N_22804,N_21873);
nor U25648 (N_25648,N_23002,N_23034);
nor U25649 (N_25649,N_24912,N_24139);
nor U25650 (N_25650,N_21305,N_23064);
nor U25651 (N_25651,N_23229,N_20578);
nor U25652 (N_25652,N_20959,N_22732);
nand U25653 (N_25653,N_23170,N_21136);
nand U25654 (N_25654,N_20037,N_22173);
nand U25655 (N_25655,N_24298,N_21906);
or U25656 (N_25656,N_23837,N_24288);
or U25657 (N_25657,N_24831,N_21558);
nor U25658 (N_25658,N_23253,N_22737);
and U25659 (N_25659,N_23341,N_22576);
or U25660 (N_25660,N_23588,N_21612);
nand U25661 (N_25661,N_21256,N_23483);
xor U25662 (N_25662,N_20081,N_22148);
and U25663 (N_25663,N_23777,N_20724);
and U25664 (N_25664,N_20386,N_24460);
and U25665 (N_25665,N_21138,N_23851);
nor U25666 (N_25666,N_22114,N_20216);
nor U25667 (N_25667,N_22086,N_24020);
nand U25668 (N_25668,N_22859,N_24654);
and U25669 (N_25669,N_23327,N_21625);
or U25670 (N_25670,N_21736,N_20230);
nor U25671 (N_25671,N_22092,N_20141);
nand U25672 (N_25672,N_22995,N_23232);
xnor U25673 (N_25673,N_24687,N_21521);
nand U25674 (N_25674,N_23418,N_21748);
or U25675 (N_25675,N_21790,N_22642);
nor U25676 (N_25676,N_22359,N_23437);
xnor U25677 (N_25677,N_22724,N_21744);
or U25678 (N_25678,N_23372,N_20495);
or U25679 (N_25679,N_24375,N_23175);
nor U25680 (N_25680,N_21311,N_21161);
or U25681 (N_25681,N_21756,N_24784);
nand U25682 (N_25682,N_20207,N_21600);
nand U25683 (N_25683,N_21627,N_22731);
nand U25684 (N_25684,N_21956,N_21127);
nor U25685 (N_25685,N_23746,N_23469);
or U25686 (N_25686,N_21217,N_23997);
nor U25687 (N_25687,N_23526,N_23377);
or U25688 (N_25688,N_20818,N_24957);
nor U25689 (N_25689,N_20071,N_21595);
or U25690 (N_25690,N_21735,N_24165);
nand U25691 (N_25691,N_22368,N_22827);
nor U25692 (N_25692,N_24586,N_21387);
and U25693 (N_25693,N_24325,N_24309);
nor U25694 (N_25694,N_20245,N_24639);
or U25695 (N_25695,N_23586,N_24082);
nor U25696 (N_25696,N_20032,N_21174);
nor U25697 (N_25697,N_23606,N_20399);
nand U25698 (N_25698,N_22419,N_23259);
nor U25699 (N_25699,N_24303,N_23094);
nor U25700 (N_25700,N_24953,N_21363);
nor U25701 (N_25701,N_22098,N_21835);
and U25702 (N_25702,N_21492,N_22658);
nor U25703 (N_25703,N_23112,N_21920);
or U25704 (N_25704,N_23295,N_23102);
or U25705 (N_25705,N_22867,N_20335);
and U25706 (N_25706,N_24154,N_22951);
nand U25707 (N_25707,N_23145,N_23417);
xor U25708 (N_25708,N_23930,N_23946);
xor U25709 (N_25709,N_20679,N_24287);
and U25710 (N_25710,N_22486,N_21487);
and U25711 (N_25711,N_21137,N_22519);
or U25712 (N_25712,N_24398,N_21528);
nor U25713 (N_25713,N_23321,N_22336);
nand U25714 (N_25714,N_22836,N_21958);
nor U25715 (N_25715,N_22124,N_23540);
or U25716 (N_25716,N_20590,N_20367);
nor U25717 (N_25717,N_24815,N_24187);
nand U25718 (N_25718,N_23095,N_22358);
nor U25719 (N_25719,N_20283,N_21470);
or U25720 (N_25720,N_21564,N_20286);
nor U25721 (N_25721,N_22725,N_23479);
and U25722 (N_25722,N_23928,N_23178);
and U25723 (N_25723,N_23756,N_20466);
nand U25724 (N_25724,N_24706,N_24835);
nor U25725 (N_25725,N_24560,N_21884);
nand U25726 (N_25726,N_20431,N_22329);
nand U25727 (N_25727,N_20516,N_22006);
nor U25728 (N_25728,N_22959,N_23151);
nand U25729 (N_25729,N_20354,N_22190);
nor U25730 (N_25730,N_22038,N_24243);
xnor U25731 (N_25731,N_20975,N_23807);
and U25732 (N_25732,N_23289,N_22647);
nor U25733 (N_25733,N_21142,N_21473);
nor U25734 (N_25734,N_22221,N_22729);
nor U25735 (N_25735,N_24756,N_22530);
or U25736 (N_25736,N_21445,N_22058);
nand U25737 (N_25737,N_20510,N_23056);
xor U25738 (N_25738,N_23441,N_23088);
and U25739 (N_25739,N_22048,N_24180);
or U25740 (N_25740,N_24186,N_24204);
and U25741 (N_25741,N_24625,N_20543);
nor U25742 (N_25742,N_21103,N_23826);
nor U25743 (N_25743,N_24094,N_23371);
nand U25744 (N_25744,N_21298,N_20868);
nor U25745 (N_25745,N_20933,N_20626);
nor U25746 (N_25746,N_21821,N_24496);
nor U25747 (N_25747,N_23583,N_20864);
and U25748 (N_25748,N_24057,N_23994);
or U25749 (N_25749,N_24133,N_20789);
nor U25750 (N_25750,N_23367,N_21490);
xor U25751 (N_25751,N_23283,N_24195);
and U25752 (N_25752,N_20297,N_20026);
or U25753 (N_25753,N_24152,N_21742);
nor U25754 (N_25754,N_22076,N_20680);
xnor U25755 (N_25755,N_20033,N_23409);
and U25756 (N_25756,N_23582,N_24906);
nand U25757 (N_25757,N_21308,N_21739);
xor U25758 (N_25758,N_20151,N_21777);
nor U25759 (N_25759,N_23827,N_24707);
and U25760 (N_25760,N_20257,N_20492);
nand U25761 (N_25761,N_24230,N_23430);
and U25762 (N_25762,N_23938,N_24418);
nor U25763 (N_25763,N_21743,N_21423);
nor U25764 (N_25764,N_21755,N_21309);
nand U25765 (N_25765,N_22245,N_24477);
nand U25766 (N_25766,N_24383,N_20469);
and U25767 (N_25767,N_23943,N_22217);
or U25768 (N_25768,N_22655,N_24787);
or U25769 (N_25769,N_20292,N_21234);
and U25770 (N_25770,N_24617,N_24232);
nor U25771 (N_25771,N_22195,N_21046);
xor U25772 (N_25772,N_23656,N_21991);
nand U25773 (N_25773,N_21391,N_20039);
nand U25774 (N_25774,N_23871,N_24658);
nor U25775 (N_25775,N_23984,N_24059);
or U25776 (N_25776,N_24039,N_21780);
or U25777 (N_25777,N_20853,N_20250);
and U25778 (N_25778,N_22004,N_21907);
nand U25779 (N_25779,N_23663,N_21079);
xnor U25780 (N_25780,N_20794,N_24297);
nor U25781 (N_25781,N_24078,N_20837);
or U25782 (N_25782,N_24028,N_20927);
or U25783 (N_25783,N_22468,N_24419);
nor U25784 (N_25784,N_22841,N_24789);
nand U25785 (N_25785,N_20548,N_23440);
nand U25786 (N_25786,N_22656,N_21680);
nand U25787 (N_25787,N_24300,N_20574);
or U25788 (N_25788,N_22242,N_21971);
and U25789 (N_25789,N_24870,N_23510);
or U25790 (N_25790,N_23870,N_22654);
nor U25791 (N_25791,N_20252,N_24994);
nand U25792 (N_25792,N_23296,N_23610);
and U25793 (N_25793,N_20582,N_21362);
or U25794 (N_25794,N_23495,N_21547);
xnor U25795 (N_25795,N_23215,N_23847);
and U25796 (N_25796,N_24679,N_22907);
nor U25797 (N_25797,N_20669,N_22847);
and U25798 (N_25798,N_22568,N_20643);
nand U25799 (N_25799,N_22824,N_23865);
and U25800 (N_25800,N_20735,N_24689);
nor U25801 (N_25801,N_23744,N_22107);
nand U25802 (N_25802,N_21191,N_23568);
or U25803 (N_25803,N_21218,N_23687);
nand U25804 (N_25804,N_23942,N_20194);
or U25805 (N_25805,N_23216,N_20721);
or U25806 (N_25806,N_22371,N_22906);
nand U25807 (N_25807,N_24251,N_23604);
xnor U25808 (N_25808,N_20336,N_23788);
nor U25809 (N_25809,N_22481,N_22552);
or U25810 (N_25810,N_23736,N_21325);
or U25811 (N_25811,N_24492,N_23684);
nor U25812 (N_25812,N_23903,N_22750);
or U25813 (N_25813,N_23993,N_23272);
nand U25814 (N_25814,N_21171,N_22207);
or U25815 (N_25815,N_21580,N_23866);
nand U25816 (N_25816,N_21629,N_22960);
nand U25817 (N_25817,N_24289,N_22424);
or U25818 (N_25818,N_23026,N_24650);
and U25819 (N_25819,N_23557,N_22667);
or U25820 (N_25820,N_24801,N_23786);
nor U25821 (N_25821,N_21043,N_23374);
or U25822 (N_25822,N_24134,N_22618);
xor U25823 (N_25823,N_23853,N_20397);
nand U25824 (N_25824,N_24127,N_23815);
nand U25825 (N_25825,N_20787,N_20762);
and U25826 (N_25826,N_22591,N_24632);
or U25827 (N_25827,N_22509,N_24140);
nor U25828 (N_25828,N_23748,N_21781);
xor U25829 (N_25829,N_22930,N_21870);
or U25830 (N_25830,N_22412,N_22117);
nor U25831 (N_25831,N_21581,N_23701);
or U25832 (N_25832,N_21203,N_22285);
or U25833 (N_25833,N_21266,N_24910);
nor U25834 (N_25834,N_24950,N_23230);
xor U25835 (N_25835,N_23344,N_24248);
or U25836 (N_25836,N_20485,N_23605);
xor U25837 (N_25837,N_21141,N_21960);
nor U25838 (N_25838,N_24726,N_22774);
and U25839 (N_25839,N_24391,N_21654);
nand U25840 (N_25840,N_24956,N_21465);
nor U25841 (N_25841,N_20858,N_21726);
or U25842 (N_25842,N_21901,N_21854);
nand U25843 (N_25843,N_21056,N_20449);
or U25844 (N_25844,N_20757,N_20113);
or U25845 (N_25845,N_23001,N_23349);
nand U25846 (N_25846,N_22589,N_21766);
and U25847 (N_25847,N_20682,N_24515);
nand U25848 (N_25848,N_23114,N_20817);
xor U25849 (N_25849,N_21513,N_20112);
nand U25850 (N_25850,N_22682,N_22626);
nand U25851 (N_25851,N_23913,N_22201);
xnor U25852 (N_25852,N_20617,N_23846);
or U25853 (N_25853,N_22099,N_20781);
nand U25854 (N_25854,N_22379,N_20080);
nand U25855 (N_25855,N_20387,N_24651);
or U25856 (N_25856,N_22819,N_23543);
or U25857 (N_25857,N_23131,N_23566);
and U25858 (N_25858,N_24338,N_23108);
xor U25859 (N_25859,N_20135,N_23060);
xnor U25860 (N_25860,N_22199,N_21721);
nor U25861 (N_25861,N_23136,N_20376);
or U25862 (N_25862,N_23952,N_20334);
and U25863 (N_25863,N_22711,N_24817);
nor U25864 (N_25864,N_24048,N_21454);
and U25865 (N_25865,N_20118,N_21164);
nand U25866 (N_25866,N_23934,N_24526);
nand U25867 (N_25867,N_21693,N_21198);
nor U25868 (N_25868,N_21432,N_20937);
or U25869 (N_25869,N_21890,N_24961);
nor U25870 (N_25870,N_20233,N_22741);
and U25871 (N_25871,N_20425,N_22964);
nor U25872 (N_25872,N_24014,N_21276);
nand U25873 (N_25873,N_22164,N_20035);
nor U25874 (N_25874,N_20851,N_20291);
nand U25875 (N_25875,N_21318,N_20041);
nor U25876 (N_25876,N_22472,N_24100);
xnor U25877 (N_25877,N_22376,N_22525);
or U25878 (N_25878,N_21434,N_22455);
or U25879 (N_25879,N_24739,N_23670);
and U25880 (N_25880,N_21750,N_23363);
nand U25881 (N_25881,N_22056,N_20623);
and U25882 (N_25882,N_20778,N_20767);
xnor U25883 (N_25883,N_20454,N_22323);
nand U25884 (N_25884,N_24601,N_20747);
or U25885 (N_25885,N_24164,N_21859);
and U25886 (N_25886,N_20326,N_24376);
or U25887 (N_25887,N_22528,N_22592);
xnor U25888 (N_25888,N_23691,N_23523);
or U25889 (N_25889,N_20289,N_23044);
xor U25890 (N_25890,N_21707,N_21222);
nor U25891 (N_25891,N_22830,N_20199);
and U25892 (N_25892,N_23897,N_24881);
nor U25893 (N_25893,N_21804,N_24162);
xnor U25894 (N_25894,N_23795,N_20861);
nor U25895 (N_25895,N_21011,N_24851);
nand U25896 (N_25896,N_22152,N_24174);
and U25897 (N_25897,N_23442,N_23725);
xor U25898 (N_25898,N_21691,N_21233);
and U25899 (N_25899,N_21493,N_24244);
and U25900 (N_25900,N_24319,N_22028);
nand U25901 (N_25901,N_20137,N_20092);
nor U25902 (N_25902,N_20168,N_21328);
nand U25903 (N_25903,N_21085,N_20515);
and U25904 (N_25904,N_24814,N_22020);
nand U25905 (N_25905,N_22735,N_24562);
xnor U25906 (N_25906,N_23146,N_20074);
and U25907 (N_25907,N_23480,N_24222);
nand U25908 (N_25908,N_22478,N_21979);
and U25909 (N_25909,N_23612,N_24400);
nand U25910 (N_25910,N_22797,N_22899);
nand U25911 (N_25911,N_21074,N_22954);
or U25912 (N_25912,N_23685,N_20166);
nand U25913 (N_25913,N_21134,N_21355);
or U25914 (N_25914,N_20213,N_20117);
nand U25915 (N_25915,N_23008,N_21860);
or U25916 (N_25916,N_20911,N_21822);
and U25917 (N_25917,N_23396,N_22454);
nor U25918 (N_25918,N_20946,N_20392);
xnor U25919 (N_25919,N_23445,N_20647);
or U25920 (N_25920,N_23740,N_23985);
or U25921 (N_25921,N_24770,N_22869);
nand U25922 (N_25922,N_22784,N_20146);
nand U25923 (N_25923,N_22885,N_20666);
nand U25924 (N_25924,N_20920,N_23556);
nand U25925 (N_25925,N_20323,N_22008);
nor U25926 (N_25926,N_21997,N_24765);
nor U25927 (N_25927,N_24660,N_20675);
nand U25928 (N_25928,N_24749,N_24937);
nor U25929 (N_25929,N_21669,N_24983);
or U25930 (N_25930,N_21661,N_21367);
xor U25931 (N_25931,N_21505,N_21110);
nand U25932 (N_25932,N_20619,N_20173);
or U25933 (N_25933,N_22513,N_20189);
nor U25934 (N_25934,N_21530,N_23027);
nand U25935 (N_25935,N_20802,N_20388);
and U25936 (N_25936,N_20419,N_22123);
nor U25937 (N_25937,N_21895,N_22929);
nand U25938 (N_25938,N_22777,N_23273);
or U25939 (N_25939,N_22767,N_24372);
nor U25940 (N_25940,N_24570,N_24356);
nor U25941 (N_25941,N_21543,N_21758);
nand U25942 (N_25942,N_23261,N_20790);
or U25943 (N_25943,N_22036,N_21996);
or U25944 (N_25944,N_24141,N_20912);
nand U25945 (N_25945,N_20337,N_22978);
and U25946 (N_25946,N_21532,N_24060);
and U25947 (N_25947,N_22864,N_22922);
or U25948 (N_25948,N_23885,N_20256);
or U25949 (N_25949,N_20491,N_20281);
nor U25950 (N_25950,N_24821,N_24427);
nor U25951 (N_25951,N_21096,N_22815);
nor U25952 (N_25952,N_22254,N_24893);
xnor U25953 (N_25953,N_24392,N_21215);
nand U25954 (N_25954,N_22234,N_20883);
and U25955 (N_25955,N_24524,N_24716);
or U25956 (N_25956,N_21274,N_21879);
nor U25957 (N_25957,N_23511,N_20850);
nor U25958 (N_25958,N_22887,N_24285);
or U25959 (N_25959,N_24090,N_20556);
nor U25960 (N_25960,N_21951,N_21893);
nor U25961 (N_25961,N_22783,N_22400);
nand U25962 (N_25962,N_20436,N_24925);
and U25963 (N_25963,N_22133,N_22950);
nand U25964 (N_25964,N_22574,N_22648);
nor U25965 (N_25965,N_24235,N_20537);
xnor U25966 (N_25966,N_20414,N_23164);
nand U25967 (N_25967,N_23591,N_20807);
and U25968 (N_25968,N_21500,N_22849);
or U25969 (N_25969,N_23031,N_22734);
or U25970 (N_25970,N_23759,N_24390);
nand U25971 (N_25971,N_22633,N_22475);
nand U25972 (N_25972,N_20625,N_20214);
nor U25973 (N_25973,N_20513,N_20418);
and U25974 (N_25974,N_22005,N_20458);
nand U25975 (N_25975,N_20328,N_24439);
nand U25976 (N_25976,N_22704,N_24750);
and U25977 (N_25977,N_22787,N_20075);
nand U25978 (N_25978,N_21100,N_23454);
nor U25979 (N_25979,N_22730,N_24719);
nor U25980 (N_25980,N_20095,N_21147);
and U25981 (N_25981,N_21259,N_22604);
or U25982 (N_25982,N_24674,N_23375);
and U25983 (N_25983,N_20632,N_22441);
xnor U25984 (N_25984,N_24633,N_22701);
nand U25985 (N_25985,N_24182,N_22508);
and U25986 (N_25986,N_23990,N_22987);
or U25987 (N_25987,N_21713,N_21950);
nor U25988 (N_25988,N_21066,N_23140);
and U25989 (N_25989,N_23353,N_23916);
and U25990 (N_25990,N_20795,N_21962);
or U25991 (N_25991,N_24585,N_24231);
xor U25992 (N_25992,N_22338,N_21917);
nor U25993 (N_25993,N_24947,N_22806);
nor U25994 (N_25994,N_24245,N_23142);
nand U25995 (N_25995,N_21630,N_22505);
nor U25996 (N_25996,N_24306,N_21271);
nor U25997 (N_25997,N_21904,N_21212);
and U25998 (N_25998,N_24107,N_23882);
nand U25999 (N_25999,N_22169,N_20877);
nor U26000 (N_26000,N_21157,N_20925);
nand U26001 (N_26001,N_22809,N_22049);
nand U26002 (N_26002,N_21463,N_23249);
and U26003 (N_26003,N_24343,N_21722);
and U26004 (N_26004,N_20742,N_22928);
nor U26005 (N_26005,N_21864,N_24834);
and U26006 (N_26006,N_20186,N_23713);
xnor U26007 (N_26007,N_24846,N_23719);
and U26008 (N_26008,N_23803,N_23704);
xnor U26009 (N_26009,N_23761,N_20191);
and U26010 (N_26010,N_23720,N_24615);
and U26011 (N_26011,N_24463,N_23421);
nor U26012 (N_26012,N_21173,N_21152);
nor U26013 (N_26013,N_24665,N_23049);
nand U26014 (N_26014,N_24634,N_21511);
and U26015 (N_26015,N_22473,N_21957);
or U26016 (N_26016,N_21741,N_22281);
and U26017 (N_26017,N_21514,N_21934);
or U26018 (N_26018,N_20866,N_23519);
nor U26019 (N_26019,N_22641,N_21415);
and U26020 (N_26020,N_24364,N_21121);
or U26021 (N_26021,N_24124,N_20708);
nor U26022 (N_26022,N_21082,N_20423);
and U26023 (N_26023,N_23506,N_22192);
or U26024 (N_26024,N_21392,N_24813);
nand U26025 (N_26025,N_21594,N_22565);
xnor U26026 (N_26026,N_21799,N_20561);
or U26027 (N_26027,N_24559,N_20589);
nor U26028 (N_26028,N_22870,N_21591);
and U26029 (N_26029,N_21740,N_20264);
nor U26030 (N_26030,N_23737,N_24620);
nand U26031 (N_26031,N_22915,N_22306);
and U26032 (N_26032,N_21583,N_24865);
nand U26033 (N_26033,N_24209,N_23379);
nand U26034 (N_26034,N_20247,N_23477);
nor U26035 (N_26035,N_20791,N_20091);
and U26036 (N_26036,N_21510,N_23368);
nand U26037 (N_26037,N_23182,N_22688);
and U26038 (N_26038,N_22428,N_21702);
nand U26039 (N_26039,N_24386,N_23311);
or U26040 (N_26040,N_20389,N_22391);
or U26041 (N_26041,N_21115,N_22411);
nor U26042 (N_26042,N_24729,N_23354);
nand U26043 (N_26043,N_22062,N_21903);
nor U26044 (N_26044,N_22064,N_22443);
nand U26045 (N_26045,N_23004,N_22445);
nor U26046 (N_26046,N_24777,N_22628);
nor U26047 (N_26047,N_21874,N_23554);
nand U26048 (N_26048,N_21832,N_23775);
nand U26049 (N_26049,N_23224,N_22722);
and U26050 (N_26050,N_24490,N_23638);
and U26051 (N_26051,N_23394,N_23287);
or U26052 (N_26052,N_21566,N_20531);
xnor U26053 (N_26053,N_23970,N_20271);
nand U26054 (N_26054,N_24313,N_24878);
nand U26055 (N_26055,N_24201,N_24422);
nand U26056 (N_26056,N_21180,N_24217);
nand U26057 (N_26057,N_20261,N_20593);
xor U26058 (N_26058,N_22146,N_20344);
nand U26059 (N_26059,N_21282,N_22331);
or U26060 (N_26060,N_21732,N_22045);
and U26061 (N_26061,N_21265,N_23313);
and U26062 (N_26062,N_20870,N_21540);
or U26063 (N_26063,N_21119,N_20690);
or U26064 (N_26064,N_24333,N_24879);
and U26065 (N_26065,N_22610,N_21961);
and U26066 (N_26066,N_21575,N_21623);
xnor U26067 (N_26067,N_24034,N_23727);
nand U26068 (N_26068,N_20919,N_22823);
nand U26069 (N_26069,N_20755,N_22740);
nor U26070 (N_26070,N_23356,N_23520);
nand U26071 (N_26071,N_23829,N_24280);
or U26072 (N_26072,N_21029,N_21793);
or U26073 (N_26073,N_21809,N_22716);
or U26074 (N_26074,N_22080,N_20967);
and U26075 (N_26075,N_21244,N_23512);
or U26076 (N_26076,N_21370,N_24590);
xor U26077 (N_26077,N_23590,N_21335);
nor U26078 (N_26078,N_21340,N_24984);
nor U26079 (N_26079,N_21765,N_20318);
or U26080 (N_26080,N_21862,N_21831);
nand U26081 (N_26081,N_20309,N_20521);
or U26082 (N_26082,N_21537,N_23243);
or U26083 (N_26083,N_22555,N_23733);
and U26084 (N_26084,N_23747,N_21095);
nor U26085 (N_26085,N_22502,N_24602);
nand U26086 (N_26086,N_22687,N_21458);
nor U26087 (N_26087,N_23901,N_23127);
or U26088 (N_26088,N_22103,N_20822);
nand U26089 (N_26089,N_22211,N_20231);
nor U26090 (N_26090,N_20732,N_24895);
and U26091 (N_26091,N_22991,N_24172);
xnor U26092 (N_26092,N_24047,N_22832);
and U26093 (N_26093,N_20109,N_24096);
or U26094 (N_26094,N_24608,N_20591);
and U26095 (N_26095,N_22465,N_20042);
nor U26096 (N_26096,N_20009,N_20210);
or U26097 (N_26097,N_20209,N_23758);
nand U26098 (N_26098,N_23935,N_20008);
xnor U26099 (N_26099,N_22575,N_22494);
nand U26100 (N_26100,N_22779,N_21501);
and U26101 (N_26101,N_24157,N_21820);
nand U26102 (N_26102,N_24199,N_22043);
nor U26103 (N_26103,N_23129,N_23570);
nor U26104 (N_26104,N_23923,N_20898);
nand U26105 (N_26105,N_22989,N_22464);
and U26106 (N_26106,N_21648,N_23563);
nand U26107 (N_26107,N_20417,N_21441);
xor U26108 (N_26108,N_22678,N_22590);
nor U26109 (N_26109,N_24926,N_21687);
and U26110 (N_26110,N_22299,N_21670);
or U26111 (N_26111,N_20222,N_20459);
or U26112 (N_26112,N_21437,N_24558);
xor U26113 (N_26113,N_22594,N_20391);
and U26114 (N_26114,N_23559,N_22652);
and U26115 (N_26115,N_20343,N_23507);
or U26116 (N_26116,N_21773,N_22236);
or U26117 (N_26117,N_20305,N_22304);
xor U26118 (N_26118,N_24914,N_24582);
nand U26119 (N_26119,N_23065,N_21894);
nor U26120 (N_26120,N_21239,N_22788);
nand U26121 (N_26121,N_22268,N_21953);
and U26122 (N_26122,N_23580,N_23271);
xnor U26123 (N_26123,N_21974,N_21406);
nand U26124 (N_26124,N_23976,N_22000);
and U26125 (N_26125,N_21160,N_20050);
or U26126 (N_26126,N_24810,N_23041);
xor U26127 (N_26127,N_21348,N_24015);
nor U26128 (N_26128,N_23832,N_20486);
nand U26129 (N_26129,N_24545,N_20824);
and U26130 (N_26130,N_22188,N_23729);
or U26131 (N_26131,N_20293,N_20736);
and U26132 (N_26132,N_21816,N_21946);
or U26133 (N_26133,N_23282,N_22612);
xor U26134 (N_26134,N_21062,N_22497);
or U26135 (N_26135,N_24128,N_22265);
nand U26136 (N_26136,N_24676,N_22283);
and U26137 (N_26137,N_21875,N_22395);
nand U26138 (N_26138,N_20422,N_21446);
nor U26139 (N_26139,N_24167,N_20347);
or U26140 (N_26140,N_24575,N_21794);
nand U26141 (N_26141,N_24647,N_20697);
or U26142 (N_26142,N_24017,N_24732);
nor U26143 (N_26143,N_21107,N_21584);
and U26144 (N_26144,N_24353,N_23675);
nor U26145 (N_26145,N_20810,N_24395);
and U26146 (N_26146,N_20306,N_21759);
or U26147 (N_26147,N_20940,N_20400);
nor U26148 (N_26148,N_24922,N_20057);
nand U26149 (N_26149,N_22572,N_24890);
or U26150 (N_26150,N_21065,N_20769);
nor U26151 (N_26151,N_20518,N_20559);
or U26152 (N_26152,N_23075,N_23534);
and U26153 (N_26153,N_23664,N_22685);
or U26154 (N_26154,N_23336,N_20351);
nand U26155 (N_26155,N_22184,N_23517);
xor U26156 (N_26156,N_22785,N_20869);
and U26157 (N_26157,N_22690,N_22083);
xnor U26158 (N_26158,N_20706,N_23639);
and U26159 (N_26159,N_23156,N_22825);
or U26160 (N_26160,N_24385,N_20443);
nor U26161 (N_26161,N_21749,N_20909);
or U26162 (N_26162,N_23974,N_21924);
and U26163 (N_26163,N_22142,N_22571);
and U26164 (N_26164,N_23773,N_22260);
nor U26165 (N_26165,N_22256,N_22681);
and U26166 (N_26166,N_21676,N_21448);
or U26167 (N_26167,N_23010,N_20224);
and U26168 (N_26168,N_22034,N_21845);
nor U26169 (N_26169,N_20110,N_23967);
or U26170 (N_26170,N_22037,N_23455);
or U26171 (N_26171,N_24417,N_21313);
nor U26172 (N_26172,N_22578,N_22039);
nand U26173 (N_26173,N_21855,N_23100);
xnor U26174 (N_26174,N_21341,N_21754);
or U26175 (N_26175,N_22003,N_22322);
and U26176 (N_26176,N_23071,N_24340);
nand U26177 (N_26177,N_22200,N_20097);
xor U26178 (N_26178,N_20642,N_24780);
nand U26179 (N_26179,N_22241,N_24667);
and U26180 (N_26180,N_21710,N_20295);
nor U26181 (N_26181,N_23843,N_24892);
nand U26182 (N_26182,N_21178,N_23077);
or U26183 (N_26183,N_24628,N_24454);
nand U26184 (N_26184,N_21916,N_21315);
and U26185 (N_26185,N_23054,N_22499);
nor U26186 (N_26186,N_21175,N_22965);
or U26187 (N_26187,N_24250,N_20059);
nand U26188 (N_26188,N_20269,N_20357);
nor U26189 (N_26189,N_24268,N_22422);
or U26190 (N_26190,N_21041,N_20947);
nor U26191 (N_26191,N_22914,N_24493);
nor U26192 (N_26192,N_23378,N_22696);
xnor U26193 (N_26193,N_21369,N_24872);
nand U26194 (N_26194,N_22762,N_24258);
nor U26195 (N_26195,N_23153,N_23823);
nand U26196 (N_26196,N_22539,N_24607);
or U26197 (N_26197,N_21719,N_23887);
or U26198 (N_26198,N_22325,N_20456);
and U26199 (N_26199,N_23579,N_24031);
xor U26200 (N_26200,N_23799,N_22988);
nor U26201 (N_26201,N_21040,N_20696);
nand U26202 (N_26202,N_20382,N_23244);
and U26203 (N_26203,N_23732,N_21188);
nand U26204 (N_26204,N_23176,N_20953);
xnor U26205 (N_26205,N_24246,N_22662);
and U26206 (N_26206,N_22248,N_23609);
and U26207 (N_26207,N_24899,N_24760);
nor U26208 (N_26208,N_23755,N_20601);
xnor U26209 (N_26209,N_22898,N_23456);
xnor U26210 (N_26210,N_24858,N_20498);
or U26211 (N_26211,N_23411,N_20668);
nor U26212 (N_26212,N_20464,N_23785);
nor U26213 (N_26213,N_21531,N_21183);
or U26214 (N_26214,N_23646,N_20707);
nor U26215 (N_26215,N_20192,N_23299);
nor U26216 (N_26216,N_22924,N_23919);
or U26217 (N_26217,N_21885,N_20372);
or U26218 (N_26218,N_24270,N_21012);
nand U26219 (N_26219,N_21568,N_24755);
nor U26220 (N_26220,N_21570,N_23324);
nand U26221 (N_26221,N_21843,N_20070);
nor U26222 (N_26222,N_20426,N_22584);
and U26223 (N_26223,N_24196,N_22720);
nand U26224 (N_26224,N_24844,N_23490);
or U26225 (N_26225,N_20624,N_21798);
nand U26226 (N_26226,N_24252,N_23245);
xnor U26227 (N_26227,N_20157,N_21076);
or U26228 (N_26228,N_20618,N_20628);
xnor U26229 (N_26229,N_21517,N_20489);
or U26230 (N_26230,N_20439,N_24761);
and U26231 (N_26231,N_22386,N_22496);
and U26232 (N_26232,N_20451,N_23138);
nor U26233 (N_26233,N_20784,N_21805);
or U26234 (N_26234,N_20835,N_20341);
and U26235 (N_26235,N_23867,N_20079);
nand U26236 (N_26236,N_24864,N_23204);
nand U26237 (N_26237,N_22997,N_20375);
or U26238 (N_26238,N_21563,N_21659);
nor U26239 (N_26239,N_24122,N_21504);
nand U26240 (N_26240,N_24278,N_22763);
xnor U26241 (N_26241,N_23845,N_23886);
nor U26242 (N_26242,N_20445,N_20077);
and U26243 (N_26243,N_21109,N_24008);
or U26244 (N_26244,N_24581,N_23598);
xor U26245 (N_26245,N_23135,N_22874);
and U26246 (N_26246,N_22781,N_22549);
and U26247 (N_26247,N_22328,N_21374);
nor U26248 (N_26248,N_20043,N_21108);
xnor U26249 (N_26249,N_23091,N_23961);
nor U26250 (N_26250,N_24535,N_24822);
or U26251 (N_26251,N_20229,N_21734);
and U26252 (N_26252,N_22611,N_20651);
and U26253 (N_26253,N_21700,N_20401);
nand U26254 (N_26254,N_22837,N_22345);
and U26255 (N_26255,N_20198,N_20296);
and U26256 (N_26256,N_24114,N_22457);
or U26257 (N_26257,N_22161,N_22409);
or U26258 (N_26258,N_22822,N_24699);
nand U26259 (N_26259,N_22178,N_22790);
nand U26260 (N_26260,N_24847,N_22369);
or U26261 (N_26261,N_20751,N_24735);
nand U26262 (N_26262,N_20424,N_23821);
xnor U26263 (N_26263,N_24703,N_23926);
and U26264 (N_26264,N_21976,N_20901);
nand U26265 (N_26265,N_20673,N_21980);
or U26266 (N_26266,N_24267,N_22880);
and U26267 (N_26267,N_22860,N_21002);
or U26268 (N_26268,N_24451,N_23059);
or U26269 (N_26269,N_24850,N_20361);
and U26270 (N_26270,N_22542,N_24929);
xor U26271 (N_26271,N_20982,N_22540);
and U26272 (N_26272,N_22524,N_24973);
and U26273 (N_26273,N_22387,N_21597);
and U26274 (N_26274,N_20303,N_24505);
xor U26275 (N_26275,N_21512,N_22517);
or U26276 (N_26276,N_23382,N_22821);
xor U26277 (N_26277,N_20826,N_22831);
nand U26278 (N_26278,N_20205,N_24286);
nand U26279 (N_26279,N_20184,N_24175);
or U26280 (N_26280,N_22440,N_24214);
and U26281 (N_26281,N_20557,N_22700);
nor U26282 (N_26282,N_24450,N_23577);
xor U26283 (N_26283,N_24967,N_22318);
or U26284 (N_26284,N_20873,N_24030);
or U26285 (N_26285,N_21770,N_20983);
and U26286 (N_26286,N_20823,N_24155);
or U26287 (N_26287,N_23717,N_24321);
nand U26288 (N_26288,N_22932,N_24476);
nor U26289 (N_26289,N_23144,N_21631);
nor U26290 (N_26290,N_24836,N_23955);
and U26291 (N_26291,N_20437,N_22759);
and U26292 (N_26292,N_22853,N_24255);
nor U26293 (N_26293,N_20939,N_22702);
nand U26294 (N_26294,N_22778,N_22794);
and U26295 (N_26295,N_23572,N_21795);
or U26296 (N_26296,N_23730,N_21846);
nand U26297 (N_26297,N_21639,N_24429);
nor U26298 (N_26298,N_20242,N_22857);
nor U26299 (N_26299,N_24342,N_21211);
nor U26300 (N_26300,N_24311,N_21871);
or U26301 (N_26301,N_21967,N_24993);
or U26302 (N_26302,N_24166,N_24382);
nand U26303 (N_26303,N_24992,N_23765);
nand U26304 (N_26304,N_20395,N_21442);
or U26305 (N_26305,N_21185,N_22973);
nor U26306 (N_26306,N_24924,N_23052);
and U26307 (N_26307,N_20160,N_23920);
or U26308 (N_26308,N_21172,N_23438);
nand U26309 (N_26309,N_24862,N_24105);
or U26310 (N_26310,N_23671,N_22040);
nand U26311 (N_26311,N_24219,N_22296);
nand U26312 (N_26312,N_24109,N_24629);
or U26313 (N_26313,N_22027,N_20355);
and U26314 (N_26314,N_24215,N_21982);
or U26315 (N_26315,N_24855,N_21292);
nor U26316 (N_26316,N_23011,N_24796);
and U26317 (N_26317,N_22087,N_24742);
nand U26318 (N_26318,N_22214,N_20981);
and U26319 (N_26319,N_20396,N_24911);
and U26320 (N_26320,N_20048,N_22015);
xnor U26321 (N_26321,N_23068,N_21696);
nor U26322 (N_26322,N_20406,N_21455);
and U26323 (N_26323,N_24663,N_20373);
and U26324 (N_26324,N_22600,N_20078);
and U26325 (N_26325,N_23619,N_21652);
nand U26326 (N_26326,N_23809,N_20957);
or U26327 (N_26327,N_22068,N_22044);
xor U26328 (N_26328,N_23550,N_23911);
or U26329 (N_26329,N_21457,N_24499);
nor U26330 (N_26330,N_21048,N_21731);
nor U26331 (N_26331,N_23387,N_23048);
and U26332 (N_26332,N_22653,N_22805);
or U26333 (N_26333,N_21665,N_23069);
nor U26334 (N_26334,N_21197,N_24794);
or U26335 (N_26335,N_20606,N_23376);
and U26336 (N_26336,N_24027,N_21684);
or U26337 (N_26337,N_21883,N_20307);
nand U26338 (N_26338,N_23366,N_23600);
nand U26339 (N_26339,N_21578,N_23822);
or U26340 (N_26340,N_20052,N_20924);
and U26341 (N_26341,N_20067,N_24409);
nand U26342 (N_26342,N_24132,N_22834);
or U26343 (N_26343,N_22500,N_21576);
nand U26344 (N_26344,N_22541,N_22111);
and U26345 (N_26345,N_24198,N_20519);
or U26346 (N_26346,N_23090,N_24465);
xor U26347 (N_26347,N_23117,N_21919);
or U26348 (N_26348,N_24464,N_20258);
nor U26349 (N_26349,N_24960,N_22673);
nand U26350 (N_26350,N_23147,N_22399);
and U26351 (N_26351,N_20470,N_22595);
and U26352 (N_26352,N_23270,N_22876);
nand U26353 (N_26353,N_20833,N_24508);
or U26354 (N_26354,N_23463,N_23672);
or U26355 (N_26355,N_24459,N_21416);
and U26356 (N_26356,N_22093,N_20726);
and U26357 (N_26357,N_20993,N_22913);
or U26358 (N_26358,N_22240,N_20943);
nand U26359 (N_26359,N_22933,N_20773);
nand U26360 (N_26360,N_22923,N_24348);
or U26361 (N_26361,N_20153,N_23650);
nand U26362 (N_26362,N_22585,N_22187);
and U26363 (N_26363,N_21181,N_23485);
nand U26364 (N_26364,N_22277,N_24604);
nor U26365 (N_26365,N_21717,N_23482);
and U26366 (N_26366,N_24190,N_24211);
nor U26367 (N_26367,N_20266,N_20713);
nand U26368 (N_26368,N_20681,N_21346);
or U26369 (N_26369,N_21219,N_24179);
xor U26370 (N_26370,N_22676,N_23154);
nor U26371 (N_26371,N_21964,N_22939);
or U26372 (N_26372,N_22482,N_22046);
nand U26373 (N_26373,N_21791,N_20704);
or U26374 (N_26374,N_23776,N_24447);
xnor U26375 (N_26375,N_20154,N_21027);
nor U26376 (N_26376,N_21833,N_22736);
xor U26377 (N_26377,N_21616,N_22873);
xnor U26378 (N_26378,N_21093,N_20204);
nor U26379 (N_26379,N_24024,N_22196);
and U26380 (N_26380,N_23416,N_21364);
and U26381 (N_26381,N_24987,N_21159);
and U26382 (N_26382,N_24240,N_21312);
xnor U26383 (N_26383,N_24871,N_23842);
and U26384 (N_26384,N_22871,N_20544);
and U26385 (N_26385,N_21801,N_23532);
nor U26386 (N_26386,N_21620,N_24086);
nor U26387 (N_26387,N_24001,N_22073);
nand U26388 (N_26388,N_24823,N_23099);
and U26389 (N_26389,N_23365,N_20339);
nor U26390 (N_26390,N_24963,N_22311);
nor U26391 (N_26391,N_23739,N_23657);
nor U26392 (N_26392,N_21619,N_20432);
nor U26393 (N_26393,N_24423,N_24012);
or U26394 (N_26394,N_20629,N_22543);
xor U26395 (N_26395,N_21485,N_24655);
nand U26396 (N_26396,N_23608,N_22157);
nand U26397 (N_26397,N_20517,N_22977);
nand U26398 (N_26398,N_24717,N_24795);
and U26399 (N_26399,N_20812,N_21667);
nor U26400 (N_26400,N_20381,N_23895);
and U26401 (N_26401,N_22215,N_21036);
nand U26402 (N_26402,N_20098,N_24637);
or U26403 (N_26403,N_21923,N_22090);
nand U26404 (N_26404,N_23466,N_21936);
xor U26405 (N_26405,N_20852,N_24630);
or U26406 (N_26406,N_21986,N_23677);
and U26407 (N_26407,N_20480,N_21571);
and U26408 (N_26408,N_21050,N_22868);
and U26409 (N_26409,N_20942,N_21366);
or U26410 (N_26410,N_20587,N_24446);
nand U26411 (N_26411,N_23932,N_22694);
and U26412 (N_26412,N_22877,N_24322);
and U26413 (N_26413,N_21010,N_22644);
xnor U26414 (N_26414,N_24116,N_22795);
or U26415 (N_26415,N_20220,N_22780);
or U26416 (N_26416,N_20700,N_21034);
nor U26417 (N_26417,N_22693,N_24802);
nor U26418 (N_26418,N_23066,N_23665);
and U26419 (N_26419,N_20727,N_20887);
xnor U26420 (N_26420,N_23702,N_20053);
nand U26421 (N_26421,N_22684,N_20522);
nor U26422 (N_26422,N_23742,N_21376);
or U26423 (N_26423,N_24564,N_23310);
or U26424 (N_26424,N_23471,N_21718);
or U26425 (N_26425,N_21900,N_20875);
nor U26426 (N_26426,N_21083,N_20805);
nand U26427 (N_26427,N_24820,N_21381);
nor U26428 (N_26428,N_24044,N_22270);
nor U26429 (N_26429,N_21516,N_23316);
or U26430 (N_26430,N_21242,N_23470);
nor U26431 (N_26431,N_22175,N_24588);
nand U26432 (N_26432,N_21912,N_21711);
and U26433 (N_26433,N_20715,N_22646);
and U26434 (N_26434,N_20181,N_24774);
xnor U26435 (N_26435,N_20892,N_20995);
xnor U26436 (N_26436,N_20526,N_21640);
nand U26437 (N_26437,N_23645,N_23410);
xnor U26438 (N_26438,N_22966,N_23073);
nor U26439 (N_26439,N_20379,N_20693);
xnor U26440 (N_26440,N_23462,N_23180);
nand U26441 (N_26441,N_20793,N_20740);
nand U26442 (N_26442,N_24316,N_23749);
or U26443 (N_26443,N_23017,N_22118);
or U26444 (N_26444,N_23030,N_24373);
or U26445 (N_26445,N_20468,N_20066);
or U26446 (N_26446,N_23810,N_24959);
nor U26447 (N_26447,N_23681,N_22074);
or U26448 (N_26448,N_24239,N_23617);
nor U26449 (N_26449,N_24085,N_24293);
xor U26450 (N_26450,N_21995,N_21725);
nor U26451 (N_26451,N_23084,N_21772);
nor U26452 (N_26452,N_24759,N_21728);
or U26453 (N_26453,N_20130,N_23334);
or U26454 (N_26454,N_20783,N_23735);
and U26455 (N_26455,N_22629,N_23628);
nor U26456 (N_26456,N_24183,N_21856);
nand U26457 (N_26457,N_21561,N_23620);
and U26458 (N_26458,N_20646,N_22390);
and U26459 (N_26459,N_23143,N_21608);
nor U26460 (N_26460,N_20090,N_22919);
nand U26461 (N_26461,N_24282,N_20884);
and U26462 (N_26462,N_23160,N_21170);
nor U26463 (N_26463,N_21017,N_24203);
xor U26464 (N_26464,N_22980,N_22630);
and U26465 (N_26465,N_21250,N_24718);
nor U26466 (N_26466,N_21556,N_23858);
xnor U26467 (N_26467,N_20500,N_20435);
or U26468 (N_26468,N_20478,N_20099);
and U26469 (N_26469,N_21858,N_22697);
nand U26470 (N_26470,N_21788,N_21554);
or U26471 (N_26471,N_22002,N_23484);
or U26472 (N_26472,N_22544,N_24645);
nand U26473 (N_26473,N_22367,N_22303);
or U26474 (N_26474,N_23680,N_20985);
and U26475 (N_26475,N_21419,N_21658);
or U26476 (N_26476,N_23649,N_23167);
xnor U26477 (N_26477,N_21388,N_20782);
nand U26478 (N_26478,N_20038,N_22659);
and U26479 (N_26479,N_22032,N_21281);
nor U26480 (N_26480,N_24819,N_24700);
nand U26481 (N_26481,N_24763,N_20383);
xnor U26482 (N_26482,N_23318,N_21106);
nor U26483 (N_26483,N_22198,N_21241);
and U26484 (N_26484,N_20404,N_24635);
nand U26485 (N_26485,N_22249,N_21182);
nand U26486 (N_26486,N_24709,N_22460);
and U26487 (N_26487,N_20963,N_22166);
nor U26488 (N_26488,N_24501,N_20004);
nor U26489 (N_26489,N_20671,N_24518);
nand U26490 (N_26490,N_23303,N_20832);
and U26491 (N_26491,N_20612,N_24803);
nand U26492 (N_26492,N_24345,N_22171);
nor U26493 (N_26493,N_22273,N_21383);
nor U26494 (N_26494,N_21637,N_24045);
and U26495 (N_26495,N_23236,N_20058);
nand U26496 (N_26496,N_23362,N_24271);
or U26497 (N_26497,N_24525,N_23959);
nor U26498 (N_26498,N_23936,N_22567);
and U26499 (N_26499,N_20107,N_23089);
nand U26500 (N_26500,N_22637,N_21515);
nor U26501 (N_26501,N_22708,N_21544);
nand U26502 (N_26502,N_24126,N_20359);
nor U26503 (N_26503,N_22452,N_20615);
or U26504 (N_26504,N_20479,N_21838);
nor U26505 (N_26505,N_24058,N_23274);
nand U26506 (N_26506,N_20069,N_22115);
xnor U26507 (N_26507,N_21385,N_20274);
nor U26508 (N_26508,N_20956,N_22875);
nor U26509 (N_26509,N_21394,N_22401);
and U26510 (N_26510,N_23277,N_23623);
and U26511 (N_26511,N_22972,N_23016);
nand U26512 (N_26512,N_21796,N_23872);
nor U26513 (N_26513,N_22334,N_21502);
and U26514 (N_26514,N_23467,N_24514);
or U26515 (N_26515,N_20941,N_21221);
or U26516 (N_26516,N_23533,N_21834);
nor U26517 (N_26517,N_24367,N_21296);
nand U26518 (N_26518,N_20915,N_20796);
nor U26519 (N_26519,N_23355,N_20665);
nor U26520 (N_26520,N_20831,N_24009);
or U26521 (N_26521,N_23996,N_21952);
and U26522 (N_26522,N_21094,N_24827);
and U26523 (N_26523,N_24358,N_22293);
nor U26524 (N_26524,N_20808,N_21483);
or U26525 (N_26525,N_23986,N_20019);
or U26526 (N_26526,N_24453,N_23315);
and U26527 (N_26527,N_23769,N_21227);
nand U26528 (N_26528,N_20944,N_24643);
or U26529 (N_26529,N_21261,N_22286);
nand U26530 (N_26530,N_23225,N_22121);
nand U26531 (N_26531,N_21638,N_21078);
or U26532 (N_26532,N_24672,N_21033);
nor U26533 (N_26533,N_24649,N_22599);
nand U26534 (N_26534,N_20672,N_23457);
nor U26535 (N_26535,N_21097,N_24531);
nor U26536 (N_26536,N_21606,N_20416);
or U26537 (N_26537,N_20893,N_23201);
and U26538 (N_26538,N_20433,N_21549);
or U26539 (N_26539,N_21452,N_23181);
nand U26540 (N_26540,N_22862,N_20827);
or U26541 (N_26541,N_20958,N_20955);
or U26542 (N_26542,N_20148,N_21358);
and U26543 (N_26543,N_22615,N_23781);
nor U26544 (N_26544,N_23908,N_20093);
and U26545 (N_26545,N_21269,N_23326);
and U26546 (N_26546,N_21284,N_24962);
nand U26547 (N_26547,N_22141,N_20730);
nor U26548 (N_26548,N_20951,N_21204);
nand U26549 (N_26549,N_20254,N_23541);
nand U26550 (N_26550,N_20450,N_20889);
nand U26551 (N_26551,N_24022,N_22580);
or U26552 (N_26552,N_21536,N_20085);
xnor U26553 (N_26553,N_23929,N_20534);
nand U26554 (N_26554,N_22816,N_24040);
nor U26555 (N_26555,N_20602,N_20609);
nor U26556 (N_26556,N_23183,N_21277);
and U26557 (N_26557,N_20904,N_24061);
or U26558 (N_26558,N_21023,N_24736);
nor U26559 (N_26559,N_23279,N_21938);
or U26560 (N_26560,N_23716,N_24226);
nor U26561 (N_26561,N_20630,N_22413);
nor U26562 (N_26562,N_20011,N_22352);
nor U26563 (N_26563,N_23364,N_24974);
and U26564 (N_26564,N_24004,N_22001);
and U26565 (N_26565,N_21935,N_20966);
nor U26566 (N_26566,N_21948,N_21323);
or U26567 (N_26567,N_22362,N_23505);
xnor U26568 (N_26568,N_23045,N_23501);
nor U26569 (N_26569,N_24746,N_24284);
xor U26570 (N_26570,N_21337,N_20913);
or U26571 (N_26571,N_23537,N_24113);
xor U26572 (N_26572,N_23459,N_24769);
and U26573 (N_26573,N_24473,N_23521);
or U26574 (N_26574,N_21343,N_24178);
nor U26575 (N_26575,N_21291,N_24659);
nor U26576 (N_26576,N_21380,N_24692);
and U26577 (N_26577,N_24593,N_22984);
nor U26578 (N_26578,N_22953,N_20596);
or U26579 (N_26579,N_22278,N_24551);
nand U26580 (N_26580,N_20541,N_23790);
nand U26581 (N_26581,N_24866,N_22900);
or U26582 (N_26582,N_23042,N_22021);
or U26583 (N_26583,N_20524,N_24069);
nor U26584 (N_26584,N_22617,N_21908);
nor U26585 (N_26585,N_24075,N_23655);
xor U26586 (N_26586,N_22417,N_21290);
xor U26587 (N_26587,N_24768,N_24828);
nand U26588 (N_26588,N_23529,N_23640);
or U26589 (N_26589,N_24118,N_23958);
nor U26590 (N_26590,N_24171,N_23806);
or U26591 (N_26591,N_24035,N_23070);
or U26592 (N_26592,N_21972,N_21927);
xor U26593 (N_26593,N_20460,N_24697);
nor U26594 (N_26594,N_23264,N_23280);
nand U26595 (N_26595,N_23448,N_24253);
and U26596 (N_26596,N_20976,N_24666);
nor U26597 (N_26597,N_20467,N_23745);
or U26598 (N_26598,N_20054,N_21417);
nand U26599 (N_26599,N_22289,N_20226);
nor U26600 (N_26600,N_22137,N_20086);
nor U26601 (N_26601,N_23325,N_23053);
or U26602 (N_26602,N_20683,N_21863);
and U26603 (N_26603,N_20771,N_23783);
xor U26604 (N_26604,N_24502,N_22253);
or U26605 (N_26605,N_24529,N_22942);
and U26606 (N_26606,N_21787,N_24609);
or U26607 (N_26607,N_22609,N_23627);
nand U26608 (N_26608,N_23854,N_20627);
nor U26609 (N_26609,N_21300,N_22427);
and U26610 (N_26610,N_21983,N_22775);
or U26611 (N_26611,N_24387,N_23339);
and U26612 (N_26612,N_24566,N_24684);
xnor U26613 (N_26613,N_24976,N_21818);
xnor U26614 (N_26614,N_24310,N_23393);
and U26615 (N_26615,N_22986,N_23323);
nand U26616 (N_26616,N_23427,N_22109);
or U26617 (N_26617,N_23718,N_21539);
and U26618 (N_26618,N_24616,N_23509);
or U26619 (N_26619,N_24404,N_21304);
or U26620 (N_26620,N_20581,N_20161);
nor U26621 (N_26621,N_22282,N_21553);
nand U26622 (N_26622,N_20062,N_22905);
nor U26623 (N_26623,N_23850,N_23006);
nand U26624 (N_26624,N_22067,N_22538);
or U26625 (N_26625,N_21902,N_22537);
or U26626 (N_26626,N_24160,N_20244);
and U26627 (N_26627,N_23078,N_24337);
and U26628 (N_26628,N_21677,N_20905);
nor U26629 (N_26629,N_23503,N_20217);
xor U26630 (N_26630,N_22703,N_22698);
and U26631 (N_26631,N_20916,N_22266);
and U26632 (N_26632,N_24965,N_22408);
or U26633 (N_26633,N_21605,N_23743);
and U26634 (N_26634,N_24003,N_24811);
nor U26635 (N_26635,N_23722,N_23055);
and U26636 (N_26636,N_24111,N_21928);
or U26637 (N_26637,N_24808,N_21481);
and U26638 (N_26638,N_21429,N_22167);
nor U26639 (N_26639,N_20476,N_24125);
nor U26640 (N_26640,N_21413,N_24611);
nand U26641 (N_26641,N_21123,N_21593);
and U26642 (N_26642,N_21826,N_20411);
or U26643 (N_26643,N_21070,N_20655);
or U26644 (N_26644,N_22026,N_24998);
or U26645 (N_26645,N_24474,N_22909);
nor U26646 (N_26646,N_20989,N_21592);
or U26647 (N_26647,N_24897,N_22031);
and U26648 (N_26648,N_24023,N_21807);
nor U26649 (N_26649,N_24664,N_21615);
or U26650 (N_26650,N_21897,N_21727);
nor U26651 (N_26651,N_23750,N_21354);
nand U26652 (N_26652,N_23439,N_24948);
and U26653 (N_26653,N_21245,N_24488);
and U26654 (N_26654,N_23115,N_24481);
nor U26655 (N_26655,N_23496,N_24475);
nor U26656 (N_26656,N_21150,N_21970);
nor U26657 (N_26657,N_23939,N_21214);
and U26658 (N_26658,N_23771,N_20287);
nor U26659 (N_26659,N_20327,N_21891);
or U26660 (N_26660,N_20638,N_21941);
or U26661 (N_26661,N_24257,N_22712);
xor U26662 (N_26662,N_23003,N_24083);
nand U26663 (N_26663,N_22562,N_24176);
and U26664 (N_26664,N_22920,N_21650);
and U26665 (N_26665,N_22373,N_23015);
or U26666 (N_26666,N_21747,N_20353);
and U26667 (N_26667,N_23763,N_21829);
and U26668 (N_26668,N_22643,N_20280);
or U26669 (N_26669,N_24677,N_20136);
nor U26670 (N_26670,N_22030,N_23629);
nand U26671 (N_26671,N_21038,N_20028);
or U26672 (N_26672,N_22893,N_24587);
and U26673 (N_26673,N_20393,N_21061);
or U26674 (N_26674,N_23263,N_21345);
and U26675 (N_26675,N_22177,N_24497);
nand U26676 (N_26676,N_24097,N_21477);
nand U26677 (N_26677,N_20577,N_20891);
or U26678 (N_26678,N_21641,N_21177);
and U26679 (N_26679,N_23132,N_24541);
nand U26680 (N_26680,N_21389,N_21724);
nand U26681 (N_26681,N_22808,N_22163);
nand U26682 (N_26682,N_21830,N_22370);
nand U26683 (N_26683,N_20565,N_23879);
nor U26684 (N_26684,N_24393,N_24824);
xnor U26685 (N_26685,N_22431,N_24873);
nand U26686 (N_26686,N_22520,N_24613);
xor U26687 (N_26687,N_20821,N_23177);
or U26688 (N_26688,N_24517,N_20481);
nor U26689 (N_26689,N_21360,N_23697);
and U26690 (N_26690,N_23226,N_22886);
or U26691 (N_26691,N_23508,N_21294);
or U26692 (N_26692,N_24555,N_20319);
and U26693 (N_26693,N_20284,N_20187);
or U26694 (N_26694,N_24516,N_23242);
nand U26695 (N_26695,N_24088,N_23386);
nor U26696 (N_26696,N_23539,N_21877);
or U26697 (N_26697,N_24104,N_22895);
xor U26698 (N_26698,N_24361,N_24678);
nand U26699 (N_26699,N_23345,N_24927);
nor U26700 (N_26700,N_20507,N_22943);
and U26701 (N_26701,N_21400,N_22743);
and U26702 (N_26702,N_23873,N_24698);
and U26703 (N_26703,N_20881,N_21451);
or U26704 (N_26704,N_24762,N_21678);
or U26705 (N_26705,N_23880,N_23487);
nor U26706 (N_26706,N_20126,N_20549);
nor U26707 (N_26707,N_21869,N_22235);
and U26708 (N_26708,N_24972,N_23018);
nand U26709 (N_26709,N_20122,N_24913);
nand U26710 (N_26710,N_22168,N_24546);
or U26711 (N_26711,N_23121,N_24537);
nand U26712 (N_26712,N_21929,N_21940);
and U26713 (N_26713,N_21586,N_20169);
xor U26714 (N_26714,N_24092,N_20051);
nor U26715 (N_26715,N_21295,N_23085);
nor U26716 (N_26716,N_23157,N_23599);
xnor U26717 (N_26717,N_22140,N_23528);
nor U26718 (N_26718,N_22403,N_20325);
or U26719 (N_26719,N_20105,N_22490);
nand U26720 (N_26720,N_24695,N_20149);
nor U26721 (N_26721,N_23991,N_21425);
nand U26722 (N_26722,N_24448,N_20717);
and U26723 (N_26723,N_20906,N_24938);
nor U26724 (N_26724,N_24197,N_23878);
nor U26725 (N_26725,N_24053,N_23291);
and U26726 (N_26726,N_21861,N_23715);
nand U26727 (N_26727,N_22091,N_21464);
nor U26728 (N_26728,N_23869,N_21887);
xor U26729 (N_26729,N_23498,N_21440);
and U26730 (N_26730,N_20766,N_20992);
or U26731 (N_26731,N_20908,N_20403);
nand U26732 (N_26732,N_20917,N_22675);
nor U26733 (N_26733,N_24205,N_24788);
nor U26734 (N_26734,N_24042,N_20234);
nand U26735 (N_26735,N_23141,N_24485);
nor U26736 (N_26736,N_21395,N_24733);
nand U26737 (N_26737,N_24291,N_22179);
and U26738 (N_26738,N_23370,N_20196);
xor U26739 (N_26739,N_21844,N_21663);
nand U26740 (N_26740,N_22670,N_20622);
nor U26741 (N_26741,N_24347,N_22016);
xnor U26742 (N_26742,N_21426,N_23391);
nor U26743 (N_26743,N_23254,N_22726);
nand U26744 (N_26744,N_21931,N_20529);
or U26745 (N_26745,N_22660,N_22156);
and U26746 (N_26746,N_22315,N_21373);
nand U26747 (N_26747,N_24826,N_24326);
or U26748 (N_26748,N_20322,N_22439);
or U26749 (N_26749,N_23861,N_21055);
nor U26750 (N_26750,N_24863,N_24478);
or U26751 (N_26751,N_22818,N_23812);
nand U26752 (N_26752,N_24223,N_24052);
or U26753 (N_26753,N_21231,N_20586);
xnor U26754 (N_26754,N_22047,N_21943);
xnor U26755 (N_26755,N_20550,N_21349);
nor U26756 (N_26756,N_24424,N_20686);
nand U26757 (N_26757,N_24068,N_22122);
nand U26758 (N_26758,N_24738,N_20930);
nand U26759 (N_26759,N_21603,N_20016);
and U26760 (N_26760,N_23802,N_24302);
and U26761 (N_26761,N_23632,N_23235);
or U26762 (N_26762,N_20394,N_23465);
nor U26763 (N_26763,N_20374,N_24056);
and U26764 (N_26764,N_20592,N_20025);
xnor U26765 (N_26765,N_23461,N_21542);
nor U26766 (N_26766,N_22287,N_22625);
and U26767 (N_26767,N_24416,N_22627);
nand U26768 (N_26768,N_24905,N_21410);
nor U26769 (N_26769,N_23924,N_24365);
or U26770 (N_26770,N_20265,N_23669);
and U26771 (N_26771,N_20285,N_20452);
or U26772 (N_26772,N_21527,N_21131);
and U26773 (N_26773,N_22757,N_24318);
and U26774 (N_26774,N_22476,N_21120);
or U26775 (N_26775,N_20228,N_22981);
or U26776 (N_26776,N_23211,N_23960);
xnor U26777 (N_26777,N_20371,N_21910);
or U26778 (N_26778,N_22204,N_24005);
nor U26779 (N_26779,N_24072,N_22861);
or U26780 (N_26780,N_24989,N_24051);
nor U26781 (N_26781,N_22935,N_22110);
and U26782 (N_26782,N_23953,N_22990);
or U26783 (N_26783,N_21852,N_21552);
nand U26784 (N_26784,N_22839,N_23859);
or U26785 (N_26785,N_21202,N_22719);
nor U26786 (N_26786,N_21088,N_21853);
nor U26787 (N_26787,N_22357,N_20820);
nand U26788 (N_26788,N_24612,N_24487);
nor U26789 (N_26789,N_22208,N_21051);
and U26790 (N_26790,N_24489,N_22010);
nand U26791 (N_26791,N_22084,N_22669);
nor U26792 (N_26792,N_22739,N_22398);
or U26793 (N_26793,N_22883,N_21303);
or U26794 (N_26794,N_20338,N_24077);
nor U26795 (N_26795,N_22471,N_20914);
or U26796 (N_26796,N_22802,N_21288);
nor U26797 (N_26797,N_21243,N_22372);
nor U26798 (N_26798,N_23678,N_24484);
nand U26799 (N_26799,N_20876,N_22351);
and U26800 (N_26800,N_20711,N_23097);
and U26801 (N_26801,N_23999,N_21745);
or U26802 (N_26802,N_20123,N_21715);
nand U26803 (N_26803,N_22349,N_24982);
nand U26804 (N_26804,N_20447,N_21001);
and U26805 (N_26805,N_21111,N_22479);
or U26806 (N_26806,N_24225,N_20731);
and U26807 (N_26807,N_23414,N_23384);
nand U26808 (N_26808,N_20719,N_22225);
and U26809 (N_26809,N_21771,N_22811);
nand U26810 (N_26810,N_24415,N_20968);
or U26811 (N_26811,N_23297,N_22820);
xor U26812 (N_26812,N_20483,N_20031);
nand U26813 (N_26813,N_21350,N_20049);
nand U26814 (N_26814,N_22017,N_22782);
or U26815 (N_26815,N_20302,N_23831);
or U26816 (N_26816,N_23863,N_22969);
nand U26817 (N_26817,N_22896,N_23544);
or U26818 (N_26818,N_22746,N_23359);
xor U26819 (N_26819,N_22955,N_21310);
nand U26820 (N_26820,N_24359,N_23337);
and U26821 (N_26821,N_24472,N_23150);
or U26822 (N_26822,N_22484,N_20096);
nor U26823 (N_26823,N_23118,N_21621);
and U26824 (N_26824,N_24720,N_22488);
xnor U26825 (N_26825,N_22550,N_22112);
or U26826 (N_26826,N_20998,N_20816);
and U26827 (N_26827,N_22940,N_20660);
nand U26828 (N_26828,N_21196,N_23780);
nor U26829 (N_26829,N_21020,N_22216);
or U26830 (N_26830,N_22182,N_22587);
and U26831 (N_26831,N_21307,N_20678);
or U26832 (N_26832,N_23828,N_20174);
or U26833 (N_26833,N_22205,N_23087);
or U26834 (N_26834,N_24357,N_24503);
and U26835 (N_26835,N_24117,N_24099);
or U26836 (N_26836,N_24837,N_24980);
xor U26837 (N_26837,N_20102,N_23412);
nand U26838 (N_26838,N_20350,N_22407);
and U26839 (N_26839,N_21496,N_21688);
and U26840 (N_26840,N_24767,N_24089);
and U26841 (N_26841,N_22573,N_23801);
nand U26842 (N_26842,N_22466,N_22843);
and U26843 (N_26843,N_20573,N_24301);
nor U26844 (N_26844,N_23120,N_24536);
nor U26845 (N_26845,N_23982,N_21965);
nor U26846 (N_26846,N_23169,N_21922);
nor U26847 (N_26847,N_20862,N_20772);
or U26848 (N_26848,N_24349,N_22094);
nor U26849 (N_26849,N_20997,N_21013);
or U26850 (N_26850,N_22560,N_21968);
xor U26851 (N_26851,N_20688,N_23569);
nor U26852 (N_26852,N_23565,N_24527);
nor U26853 (N_26853,N_20600,N_21746);
nand U26854 (N_26854,N_22210,N_21769);
nand U26855 (N_26855,N_21092,N_22014);
nor U26856 (N_26856,N_24889,N_24764);
nor U26857 (N_26857,N_23340,N_24533);
and U26858 (N_26858,N_23764,N_20845);
or U26859 (N_26859,N_24999,N_21590);
and U26860 (N_26860,N_23940,N_20907);
or U26861 (N_26861,N_21344,N_21270);
nor U26862 (N_26862,N_20753,N_21840);
nand U26863 (N_26863,N_22851,N_20977);
nor U26864 (N_26864,N_24908,N_22956);
or U26865 (N_26865,N_21176,N_22072);
xnor U26866 (N_26866,N_23257,N_24188);
nor U26867 (N_26867,N_24623,N_23251);
nand U26868 (N_26868,N_24037,N_22343);
nor U26869 (N_26869,N_22194,N_21057);
or U26870 (N_26870,N_20317,N_24977);
or U26871 (N_26871,N_24315,N_24449);
and U26872 (N_26872,N_20484,N_21738);
nor U26873 (N_26873,N_23698,N_20934);
or U26874 (N_26874,N_24638,N_20163);
nor U26875 (N_26875,N_20448,N_24825);
and U26876 (N_26876,N_20540,N_22996);
xnor U26877 (N_26877,N_22143,N_21301);
or U26878 (N_26878,N_20409,N_24413);
nand U26879 (N_26879,N_24540,N_23904);
nand U26880 (N_26880,N_20775,N_23585);
and U26881 (N_26881,N_22564,N_22533);
and U26882 (N_26882,N_21817,N_21462);
and U26883 (N_26883,N_23666,N_21548);
nor U26884 (N_26884,N_23238,N_20961);
nand U26885 (N_26885,N_24013,N_23494);
nor U26886 (N_26886,N_22007,N_21933);
nor U26887 (N_26887,N_23589,N_21468);
nor U26888 (N_26888,N_22751,N_21035);
nand U26889 (N_26889,N_23614,N_24098);
nor U26890 (N_26890,N_24018,N_20106);
and U26891 (N_26891,N_20243,N_22534);
and U26892 (N_26892,N_24151,N_24019);
and U26893 (N_26893,N_22119,N_20501);
and U26894 (N_26894,N_23392,N_23497);
and U26895 (N_26895,N_21767,N_22522);
nand U26896 (N_26896,N_21032,N_22925);
nor U26897 (N_26897,N_24930,N_24320);
nor U26898 (N_26898,N_23284,N_20814);
nor U26899 (N_26899,N_20604,N_21994);
nand U26900 (N_26900,N_23431,N_20324);
or U26901 (N_26901,N_22364,N_22053);
or U26902 (N_26902,N_22699,N_20407);
nand U26903 (N_26903,N_20551,N_21847);
nand U26904 (N_26904,N_23228,N_20251);
nand U26905 (N_26905,N_23762,N_24412);
nor U26906 (N_26906,N_23618,N_23651);
and U26907 (N_26907,N_23643,N_24437);
nor U26908 (N_26908,N_23917,N_23199);
or U26909 (N_26909,N_24901,N_21657);
nand U26910 (N_26910,N_23352,N_20882);
nand U26911 (N_26911,N_24237,N_20428);
nor U26912 (N_26912,N_20739,N_21993);
and U26913 (N_26913,N_22231,N_23514);
nand U26914 (N_26914,N_21132,N_22892);
nand U26915 (N_26915,N_24548,N_24150);
and U26916 (N_26916,N_20579,N_23751);
or U26917 (N_26917,N_24569,N_22758);
nand U26918 (N_26918,N_21672,N_20114);
nor U26919 (N_26919,N_23202,N_20962);
nor U26920 (N_26920,N_22348,N_22840);
nand U26921 (N_26921,N_21999,N_20040);
xnor U26922 (N_26922,N_24818,N_22994);
or U26923 (N_26923,N_24080,N_20879);
and U26924 (N_26924,N_22406,N_23696);
or U26925 (N_26925,N_20785,N_24504);
nand U26926 (N_26926,N_23278,N_20725);
and U26927 (N_26927,N_20108,N_22786);
or U26928 (N_26928,N_20848,N_20348);
or U26929 (N_26929,N_22554,N_22309);
nor U26930 (N_26930,N_24714,N_21524);
nand U26931 (N_26931,N_22912,N_20171);
nand U26932 (N_26932,N_23500,N_22531);
xor U26933 (N_26933,N_24669,N_21825);
and U26934 (N_26934,N_22752,N_20176);
and U26935 (N_26935,N_20023,N_20583);
xnor U26936 (N_26936,N_20331,N_21472);
and U26937 (N_26937,N_23124,N_22683);
and U26938 (N_26938,N_20027,N_23992);
or U26939 (N_26939,N_20545,N_20368);
nor U26940 (N_26940,N_20865,N_23172);
nor U26941 (N_26941,N_22674,N_22487);
or U26942 (N_26942,N_24656,N_23699);
or U26943 (N_26943,N_22429,N_24592);
nand U26944 (N_26944,N_24269,N_24074);
nand U26945 (N_26945,N_24547,N_23937);
or U26946 (N_26946,N_20300,N_23468);
and U26947 (N_26947,N_23436,N_21003);
xor U26948 (N_26948,N_24308,N_24931);
nor U26949 (N_26949,N_21507,N_22948);
and U26950 (N_26950,N_23492,N_24969);
nor U26951 (N_26951,N_22744,N_21112);
xnor U26952 (N_26952,N_21187,N_20712);
or U26953 (N_26953,N_22536,N_23998);
and U26954 (N_26954,N_20002,N_22705);
nor U26955 (N_26955,N_21973,N_22102);
nand U26956 (N_26956,N_21102,N_21737);
or U26957 (N_26957,N_21320,N_24534);
xnor U26958 (N_26958,N_22075,N_22826);
and U26959 (N_26959,N_21480,N_20530);
nor U26960 (N_26960,N_24076,N_23464);
or U26961 (N_26961,N_23531,N_20728);
nand U26962 (N_26962,N_21153,N_20828);
xor U26963 (N_26963,N_23191,N_20315);
and U26964 (N_26964,N_23000,N_20509);
xnor U26965 (N_26965,N_23767,N_24266);
and U26966 (N_26966,N_23862,N_23995);
nand U26967 (N_26967,N_20203,N_23050);
nor U26968 (N_26968,N_24971,N_21411);
or U26969 (N_26969,N_21802,N_24290);
nand U26970 (N_26970,N_24264,N_22380);
and U26971 (N_26971,N_22559,N_24366);
and U26972 (N_26972,N_23856,N_22326);
nor U26973 (N_26973,N_23246,N_24511);
or U26974 (N_26974,N_21618,N_24238);
nor U26975 (N_26975,N_20871,N_20235);
and U26976 (N_26976,N_24614,N_23302);
nand U26977 (N_26977,N_20948,N_24928);
and U26978 (N_26978,N_24624,N_23285);
xnor U26979 (N_26979,N_24812,N_23668);
and U26980 (N_26980,N_23706,N_24227);
and U26981 (N_26981,N_20855,N_24785);
nor U26982 (N_26982,N_21645,N_23407);
nor U26983 (N_26983,N_20421,N_23857);
and U26984 (N_26984,N_22101,N_22518);
nand U26985 (N_26985,N_24941,N_24327);
and U26986 (N_26986,N_21898,N_22586);
xor U26987 (N_26987,N_20420,N_22911);
xor U26988 (N_26988,N_23968,N_20886);
or U26989 (N_26989,N_21264,N_21849);
nor U26990 (N_26990,N_21911,N_21789);
or U26991 (N_26991,N_21225,N_22828);
nand U26992 (N_26992,N_22197,N_21689);
nor U26993 (N_26993,N_21342,N_23292);
or U26994 (N_26994,N_21122,N_20563);
and U26995 (N_26995,N_20763,N_22527);
or U26996 (N_26996,N_22545,N_24441);
nor U26997 (N_26997,N_22396,N_23772);
and U26998 (N_26998,N_21008,N_22437);
or U26999 (N_26999,N_22022,N_20729);
or U27000 (N_27000,N_22052,N_23329);
nor U27001 (N_27001,N_22760,N_24970);
or U27002 (N_27002,N_23460,N_20505);
nor U27003 (N_27003,N_24438,N_21668);
and U27004 (N_27004,N_20267,N_22801);
and U27005 (N_27005,N_24523,N_23898);
or U27006 (N_27006,N_23567,N_23787);
nor U27007 (N_27007,N_21435,N_24778);
or U27008 (N_27008,N_24202,N_23168);
xnor U27009 (N_27009,N_21053,N_20063);
and U27010 (N_27010,N_23346,N_21779);
or U27011 (N_27011,N_23804,N_23196);
nor U27012 (N_27012,N_23676,N_23977);
nor U27013 (N_27013,N_22275,N_23123);
and U27014 (N_27014,N_23281,N_24330);
nor U27015 (N_27015,N_24782,N_23161);
or U27016 (N_27016,N_24567,N_21412);
nor U27017 (N_27017,N_20585,N_21101);
nor U27018 (N_27018,N_23155,N_22127);
xnor U27019 (N_27019,N_21889,N_24038);
nand U27020 (N_27020,N_23921,N_23594);
nor U27021 (N_27021,N_21226,N_21567);
nand U27022 (N_27022,N_24618,N_24867);
or U27023 (N_27023,N_23212,N_21498);
nand U27024 (N_27024,N_21876,N_23849);
or U27025 (N_27025,N_23551,N_20356);
and U27026 (N_27026,N_20648,N_21582);
nand U27027 (N_27027,N_24842,N_23473);
nand U27028 (N_27028,N_22967,N_23171);
nor U27029 (N_27029,N_20260,N_21257);
nor U27030 (N_27030,N_21778,N_21190);
nand U27031 (N_27031,N_22493,N_23237);
nor U27032 (N_27032,N_22420,N_22689);
nor U27033 (N_27033,N_24766,N_21026);
and U27034 (N_27034,N_24414,N_22191);
nor U27035 (N_27035,N_23106,N_24435);
and U27036 (N_27036,N_20201,N_23877);
xnor U27037 (N_27037,N_23927,N_23636);
or U27038 (N_27038,N_21460,N_22846);
or U27039 (N_27039,N_20494,N_24781);
or U27040 (N_27040,N_21827,N_20259);
xor U27041 (N_27041,N_24888,N_21128);
and U27042 (N_27042,N_24405,N_24840);
and U27043 (N_27043,N_22845,N_20637);
and U27044 (N_27044,N_23223,N_21450);
nand U27045 (N_27045,N_20061,N_24610);
nand U27046 (N_27046,N_24661,N_24696);
nand U27047 (N_27047,N_23578,N_24550);
nor U27048 (N_27048,N_24946,N_24538);
nor U27049 (N_27049,N_22910,N_23892);
or U27050 (N_27050,N_23989,N_23290);
xor U27051 (N_27051,N_21587,N_23615);
or U27052 (N_27052,N_20430,N_21124);
or U27053 (N_27053,N_21014,N_22447);
and U27054 (N_27054,N_24500,N_24305);
and U27055 (N_27055,N_20659,N_23525);
and U27056 (N_27056,N_21760,N_24671);
and U27057 (N_27057,N_22185,N_24887);
and U27058 (N_27058,N_21989,N_20746);
nand U27059 (N_27059,N_22728,N_21042);
nand U27060 (N_27060,N_23040,N_21433);
nand U27061 (N_27061,N_23101,N_20811);
nand U27062 (N_27062,N_21526,N_21560);
nor U27063 (N_27063,N_24102,N_24352);
or U27064 (N_27064,N_24323,N_22095);
nor U27065 (N_27065,N_22421,N_23425);
nor U27066 (N_27066,N_23703,N_22353);
or U27067 (N_27067,N_22582,N_22663);
and U27068 (N_27068,N_22055,N_24949);
or U27069 (N_27069,N_21709,N_20605);
nor U27070 (N_27070,N_20607,N_24933);
or U27071 (N_27071,N_22330,N_20290);
nand U27072 (N_27072,N_23240,N_21059);
and U27073 (N_27073,N_24194,N_24653);
nand U27074 (N_27074,N_23835,N_22621);
nor U27075 (N_27075,N_21886,N_23007);
and U27076 (N_27076,N_22718,N_22088);
xnor U27077 (N_27077,N_23596,N_21238);
or U27078 (N_27078,N_21461,N_20710);
nor U27079 (N_27079,N_20774,N_24737);
nand U27080 (N_27080,N_21447,N_20695);
and U27081 (N_27081,N_24509,N_23705);
and U27082 (N_27082,N_21045,N_23116);
nand U27083 (N_27083,N_23047,N_22238);
nand U27084 (N_27084,N_24579,N_22931);
nand U27085 (N_27085,N_21880,N_20611);
xor U27086 (N_27086,N_20716,N_23948);
and U27087 (N_27087,N_24479,N_20313);
nor U27088 (N_27088,N_21118,N_22738);
and U27089 (N_27089,N_22916,N_21486);
nand U27090 (N_27090,N_21899,N_20007);
nand U27091 (N_27091,N_21135,N_20190);
nor U27092 (N_27092,N_22814,N_22491);
and U27093 (N_27093,N_20564,N_24681);
and U27094 (N_27094,N_22453,N_22404);
and U27095 (N_27095,N_23951,N_20684);
nor U27096 (N_27096,N_22365,N_21230);
or U27097 (N_27097,N_23385,N_24869);
and U27098 (N_27098,N_23219,N_20701);
and U27099 (N_27099,N_22971,N_24218);
nand U27100 (N_27100,N_20111,N_21776);
or U27101 (N_27101,N_21589,N_22228);
nand U27102 (N_27102,N_22333,N_22363);
xnor U27103 (N_27103,N_21194,N_22557);
or U27104 (N_27104,N_23893,N_20614);
or U27105 (N_27105,N_21028,N_22250);
or U27106 (N_27106,N_20275,N_23402);
nor U27107 (N_27107,N_23637,N_22813);
and U27108 (N_27108,N_20702,N_22220);
or U27109 (N_27109,N_21283,N_20378);
nand U27110 (N_27110,N_23166,N_21099);
and U27111 (N_27111,N_22251,N_21021);
or U27112 (N_27112,N_24589,N_20465);
and U27113 (N_27113,N_22154,N_23491);
nor U27114 (N_27114,N_24744,N_20047);
and U27115 (N_27115,N_21353,N_24480);
nand U27116 (N_27116,N_20806,N_22206);
and U27117 (N_27117,N_23400,N_24108);
nor U27118 (N_27118,N_21990,N_22526);
and U27119 (N_27119,N_22308,N_24380);
nand U27120 (N_27120,N_24350,N_21347);
nor U27121 (N_27121,N_22649,N_23700);
or U27122 (N_27122,N_22985,N_20088);
xnor U27123 (N_27123,N_24050,N_21969);
nand U27124 (N_27124,N_22962,N_20206);
nand U27125 (N_27125,N_20477,N_20276);
nand U27126 (N_27126,N_22393,N_24184);
xor U27127 (N_27127,N_23778,N_24853);
and U27128 (N_27128,N_22451,N_23964);
and U27129 (N_27129,N_21937,N_24431);
or U27130 (N_27130,N_20147,N_20029);
nand U27131 (N_27131,N_22449,N_24532);
and U27132 (N_27132,N_24758,N_23210);
or U27133 (N_27133,N_20170,N_20415);
and U27134 (N_27134,N_21644,N_22264);
and U27135 (N_27135,N_23301,N_24713);
nor U27136 (N_27136,N_23057,N_21535);
nor U27137 (N_27137,N_21562,N_22458);
nand U27138 (N_27138,N_24294,N_24797);
or U27139 (N_27139,N_20965,N_20000);
nor U27140 (N_27140,N_23988,N_20842);
nor U27141 (N_27141,N_20752,N_24603);
nor U27142 (N_27142,N_23813,N_20703);
xnor U27143 (N_27143,N_23561,N_23545);
xor U27144 (N_27144,N_20972,N_22405);
or U27145 (N_27145,N_22186,N_21456);
nand U27146 (N_27146,N_20910,N_21405);
nor U27147 (N_27147,N_24935,N_21529);
nor U27148 (N_27148,N_20539,N_21704);
nor U27149 (N_27149,N_20084,N_20687);
xnor U27150 (N_27150,N_22511,N_20013);
and U27151 (N_27151,N_20497,N_24990);
or U27152 (N_27152,N_23896,N_20644);
or U27153 (N_27153,N_20012,N_23451);
and U27154 (N_27154,N_23603,N_20764);
nor U27155 (N_27155,N_20036,N_22970);
nand U27156 (N_27156,N_24295,N_21220);
xnor U27157 (N_27157,N_21067,N_22054);
nand U27158 (N_27158,N_23305,N_20060);
nor U27159 (N_27159,N_24644,N_21444);
and U27160 (N_27160,N_21541,N_20714);
xnor U27161 (N_27161,N_24119,N_23137);
nand U27162 (N_27162,N_22947,N_22012);
nor U27163 (N_27163,N_23025,N_23797);
or U27164 (N_27164,N_24153,N_21149);
nand U27165 (N_27165,N_20195,N_22854);
or U27166 (N_27166,N_22332,N_23194);
or U27167 (N_27167,N_22272,N_21909);
nand U27168 (N_27168,N_20897,N_22434);
or U27169 (N_27169,N_23658,N_21892);
or U27170 (N_27170,N_24622,N_23683);
and U27171 (N_27171,N_23630,N_22450);
nand U27172 (N_27172,N_24494,N_24462);
nand U27173 (N_27173,N_20362,N_22042);
and U27174 (N_27174,N_20567,N_23907);
or U27175 (N_27175,N_20653,N_24368);
nor U27176 (N_27176,N_20249,N_24900);
xnor U27177 (N_27177,N_20857,N_20756);
and U27178 (N_27178,N_23380,N_23139);
nand U27179 (N_27179,N_22961,N_22521);
xnor U27180 (N_27180,N_21559,N_23504);
or U27181 (N_27181,N_21189,N_24556);
or U27182 (N_27182,N_21682,N_23390);
nor U27183 (N_27183,N_22583,N_22624);
and U27184 (N_27184,N_24208,N_20045);
nand U27185 (N_27185,N_22957,N_24945);
and U27186 (N_27186,N_22013,N_24771);
nand U27187 (N_27187,N_23981,N_24137);
nor U27188 (N_27188,N_24506,N_22290);
and U27189 (N_27189,N_22120,N_24241);
nand U27190 (N_27190,N_22936,N_21588);
and U27191 (N_27191,N_23816,N_20308);
nor U27192 (N_27192,N_21453,N_22727);
nor U27193 (N_27193,N_20532,N_24902);
xor U27194 (N_27194,N_24274,N_20129);
nor U27195 (N_27195,N_23478,N_21260);
nor U27196 (N_27196,N_23096,N_21375);
nor U27197 (N_27197,N_22316,N_21166);
and U27198 (N_27198,N_20377,N_24213);
nor U27199 (N_27199,N_24043,N_21774);
or U27200 (N_27200,N_22597,N_23987);
nand U27201 (N_27201,N_20520,N_23406);
nand U27202 (N_27202,N_21930,N_22792);
and U27203 (N_27203,N_21656,N_21146);
nor U27204 (N_27204,N_22134,N_21232);
xnor U27205 (N_27205,N_22607,N_20502);
nor U27206 (N_27206,N_20838,N_20576);
nand U27207 (N_27207,N_20759,N_23522);
or U27208 (N_27208,N_23673,N_22949);
xor U27209 (N_27209,N_21209,N_21939);
or U27210 (N_27210,N_22677,N_23217);
xnor U27211 (N_27211,N_24123,N_23688);
nand U27212 (N_27212,N_22768,N_20895);
and U27213 (N_27213,N_20635,N_24594);
nor U27214 (N_27214,N_21988,N_20709);
nand U27215 (N_27215,N_21607,N_22442);
xor U27216 (N_27216,N_24436,N_24507);
or U27217 (N_27217,N_23426,N_21785);
or U27218 (N_27218,N_22057,N_21764);
or U27219 (N_27219,N_20073,N_21708);
xor U27220 (N_27220,N_22158,N_24055);
and U27221 (N_27221,N_20987,N_21733);
or U27222 (N_27222,N_22810,N_20903);
nor U27223 (N_27223,N_24401,N_24539);
xor U27224 (N_27224,N_24683,N_24249);
or U27225 (N_27225,N_22601,N_24434);
nor U27226 (N_27226,N_24378,N_22145);
xnor U27227 (N_27227,N_24690,N_21125);
or U27228 (N_27228,N_20797,N_20991);
nand U27229 (N_27229,N_21116,N_24734);
nor U27230 (N_27230,N_23694,N_24854);
xnor U27231 (N_27231,N_21614,N_22209);
and U27232 (N_27232,N_21104,N_22776);
or U27233 (N_27233,N_20017,N_23227);
nor U27234 (N_27234,N_22432,N_20633);
nand U27235 (N_27235,N_23875,N_24883);
xnor U27236 (N_27236,N_22375,N_24371);
xor U27237 (N_27237,N_24351,N_22968);
nand U27238 (N_27238,N_20014,N_21427);
or U27239 (N_27239,N_21761,N_23103);
nor U27240 (N_27240,N_24389,N_23622);
and U27241 (N_27241,N_20945,N_22227);
and U27242 (N_27242,N_20277,N_21690);
or U27243 (N_27243,N_23306,N_23838);
nor U27244 (N_27244,N_22147,N_24578);
nand U27245 (N_27245,N_21352,N_23331);
and U27246 (N_27246,N_21867,N_21378);
and U27247 (N_27247,N_21163,N_23198);
nor U27248 (N_27248,N_20664,N_23024);
or U27249 (N_27249,N_24839,N_20273);
and U27250 (N_27250,N_20779,N_24142);
or U27251 (N_27251,N_24324,N_20801);
xor U27252 (N_27252,N_21236,N_22761);
nor U27253 (N_27253,N_22463,N_24841);
or U27254 (N_27254,N_20815,N_24932);
or U27255 (N_27255,N_22707,N_24471);
and U27256 (N_27256,N_21635,N_23607);
nor U27257 (N_27257,N_23602,N_23548);
nor U27258 (N_27258,N_21786,N_24021);
or U27259 (N_27259,N_23513,N_21803);
xnor U27260 (N_27260,N_23876,N_24919);
nand U27261 (N_27261,N_20984,N_20878);
and U27262 (N_27262,N_20208,N_20487);
or U27263 (N_27263,N_24740,N_24049);
xnor U27264 (N_27264,N_21611,N_24722);
xor U27265 (N_27265,N_22515,N_20412);
xor U27266 (N_27266,N_22155,N_23043);
xnor U27267 (N_27267,N_23824,N_23817);
nor U27268 (N_27268,N_20384,N_21823);
nand U27269 (N_27269,N_24680,N_24943);
nand U27270 (N_27270,N_22189,N_20349);
nor U27271 (N_27271,N_22203,N_20640);
xor U27272 (N_27272,N_22159,N_24923);
xnor U27273 (N_27273,N_21247,N_21633);
nand U27274 (N_27274,N_20761,N_20132);
or U27275 (N_27275,N_21675,N_20843);
nand U27276 (N_27276,N_22679,N_22773);
or U27277 (N_27277,N_22976,N_22927);
nand U27278 (N_27278,N_22385,N_24410);
and U27279 (N_27279,N_24648,N_22548);
or U27280 (N_27280,N_23945,N_24727);
xor U27281 (N_27281,N_20798,N_23770);
and U27282 (N_27282,N_24093,N_24452);
nand U27283 (N_27283,N_22024,N_20523);
and U27284 (N_27284,N_20508,N_21139);
and U27285 (N_27285,N_20720,N_24786);
nor U27286 (N_27286,N_24978,N_21223);
xor U27287 (N_27287,N_21714,N_23489);
xnor U27288 (N_27288,N_23983,N_22982);
xor U27289 (N_27289,N_20846,N_21495);
nor U27290 (N_27290,N_23200,N_20699);
or U27291 (N_27291,N_20890,N_23558);
nor U27292 (N_27292,N_22563,N_20434);
and U27293 (N_27293,N_24903,N_21165);
and U27294 (N_27294,N_22918,N_20270);
nand U27295 (N_27295,N_24025,N_23035);
or U27296 (N_27296,N_20056,N_23553);
or U27297 (N_27297,N_21263,N_24370);
and U27298 (N_27298,N_22619,N_20986);
and U27299 (N_27299,N_22686,N_23784);
nand U27300 (N_27300,N_23422,N_24798);
nor U27301 (N_27301,N_23266,N_23231);
xor U27302 (N_27302,N_21449,N_22714);
or U27303 (N_27303,N_23475,N_21200);
nor U27304 (N_27304,N_23642,N_20150);
or U27305 (N_27305,N_20427,N_23014);
or U27306 (N_27306,N_21482,N_20990);
nor U27307 (N_27307,N_24317,N_21601);
nor U27308 (N_27308,N_21403,N_24597);
nor U27309 (N_27309,N_24071,N_23634);
and U27310 (N_27310,N_22307,N_21674);
nor U27311 (N_27311,N_21000,N_20294);
nor U27312 (N_27312,N_24328,N_21841);
nand U27313 (N_27313,N_24192,N_22498);
or U27314 (N_27314,N_21331,N_24466);
xor U27315 (N_27315,N_20849,N_22884);
or U27316 (N_27316,N_20568,N_23428);
nor U27317 (N_27317,N_21506,N_23613);
nor U27318 (N_27318,N_22050,N_21072);
xnor U27319 (N_27319,N_21229,N_22106);
nor U27320 (N_27320,N_24688,N_22999);
or U27321 (N_27321,N_23708,N_21646);
xor U27322 (N_27322,N_24951,N_20193);
and U27323 (N_27323,N_23641,N_23408);
and U27324 (N_27324,N_20603,N_24783);
nand U27325 (N_27325,N_20960,N_24206);
and U27326 (N_27326,N_24884,N_22946);
and U27327 (N_27327,N_23584,N_22570);
nor U27328 (N_27328,N_21201,N_20162);
or U27329 (N_27329,N_24036,N_23757);
or U27330 (N_27330,N_24163,N_22029);
nor U27331 (N_27331,N_21792,N_24876);
or U27332 (N_27332,N_24468,N_22009);
and U27333 (N_27333,N_21478,N_20936);
nor U27334 (N_27334,N_23205,N_21649);
nor U27335 (N_27335,N_20776,N_22634);
and U27336 (N_27336,N_23624,N_21888);
nand U27337 (N_27337,N_24519,N_20533);
nand U27338 (N_27338,N_24626,N_21574);
or U27339 (N_27339,N_23399,N_23957);
xor U27340 (N_27340,N_21624,N_23276);
and U27341 (N_27341,N_24276,N_22507);
xnor U27342 (N_27342,N_23220,N_20065);
nor U27343 (N_27343,N_24916,N_21992);
and U27344 (N_27344,N_21069,N_22126);
and U27345 (N_27345,N_23021,N_20263);
or U27346 (N_27346,N_21947,N_23738);
nand U27347 (N_27347,N_22577,N_21006);
nor U27348 (N_27348,N_20018,N_20101);
nor U27349 (N_27349,N_20786,N_23037);
or U27350 (N_27350,N_23841,N_21494);
xnor U27351 (N_27351,N_22581,N_22415);
or U27352 (N_27352,N_21019,N_20542);
or U27353 (N_27353,N_20641,N_22721);
nand U27354 (N_27354,N_23741,N_23032);
and U27355 (N_27355,N_20780,N_24081);
nand U27356 (N_27356,N_22138,N_20024);
and U27357 (N_27357,N_21322,N_24670);
nand U27358 (N_27358,N_21151,N_21297);
nor U27359 (N_27359,N_20595,N_22402);
nor U27360 (N_27360,N_21610,N_21316);
nand U27361 (N_27361,N_20055,N_20127);
xnor U27362 (N_27362,N_20440,N_20854);
or U27363 (N_27363,N_21195,N_22588);
and U27364 (N_27364,N_24711,N_22547);
xnor U27365 (N_27365,N_21382,N_21697);
and U27366 (N_27366,N_23058,N_24857);
nand U27367 (N_27367,N_22717,N_24776);
and U27368 (N_27368,N_20329,N_23076);
nor U27369 (N_27369,N_20691,N_20738);
nand U27370 (N_27370,N_23403,N_23538);
or U27371 (N_27371,N_24193,N_23535);
and U27372 (N_27372,N_22344,N_24228);
xnor U27373 (N_27373,N_22150,N_23752);
or U27374 (N_27374,N_22958,N_21617);
nand U27375 (N_27375,N_20658,N_20241);
and U27376 (N_27376,N_24809,N_23207);
nand U27377 (N_27377,N_23081,N_21815);
nand U27378 (N_27378,N_20010,N_22130);
or U27379 (N_27379,N_21361,N_24640);
nand U27380 (N_27380,N_21015,N_22305);
nand U27381 (N_27381,N_24131,N_22579);
nor U27382 (N_27382,N_24377,N_21327);
or U27383 (N_27383,N_22535,N_24939);
and U27384 (N_27384,N_21140,N_24641);
and U27385 (N_27385,N_22255,N_21018);
and U27386 (N_27386,N_21706,N_24406);
nor U27387 (N_27387,N_21351,N_24296);
nor U27388 (N_27388,N_20929,N_20503);
and U27389 (N_27389,N_23659,N_20980);
nor U27390 (N_27390,N_24207,N_22313);
xor U27391 (N_27391,N_20847,N_20988);
nand U27392 (N_27392,N_24144,N_23444);
nand U27393 (N_27393,N_24159,N_21499);
and U27394 (N_27394,N_23308,N_24574);
nor U27395 (N_27395,N_22901,N_21837);
and U27396 (N_27396,N_23185,N_24772);
nor U27397 (N_27397,N_24694,N_21596);
or U27398 (N_27398,N_21249,N_23432);
or U27399 (N_27399,N_22125,N_20279);
and U27400 (N_27400,N_21424,N_24397);
nor U27401 (N_27401,N_24281,N_22132);
or U27402 (N_27402,N_22908,N_20253);
or U27403 (N_27403,N_21253,N_23969);
and U27404 (N_27404,N_23709,N_20278);
and U27405 (N_27405,N_20834,N_20442);
or U27406 (N_27406,N_22558,N_23148);
nor U27407 (N_27407,N_24728,N_23036);
nor U27408 (N_27408,N_24063,N_21439);
nor U27409 (N_27409,N_23644,N_20272);
and U27410 (N_27410,N_21024,N_23086);
nand U27411 (N_27411,N_22523,N_22842);
xor U27412 (N_27412,N_22755,N_21039);
nor U27413 (N_27413,N_23692,N_22606);
nor U27414 (N_27414,N_23179,N_24002);
and U27415 (N_27415,N_22230,N_21321);
nor U27416 (N_27416,N_23894,N_21333);
nand U27417 (N_27417,N_20970,N_20364);
and U27418 (N_27418,N_20299,N_20429);
nand U27419 (N_27419,N_22504,N_20453);
and U27420 (N_27420,N_22706,N_22715);
nor U27421 (N_27421,N_24596,N_21692);
nor U27422 (N_27422,N_20971,N_20314);
and U27423 (N_27423,N_21872,N_24832);
nand U27424 (N_27424,N_21401,N_21705);
or U27425 (N_27425,N_21651,N_22337);
and U27426 (N_27426,N_23950,N_24070);
or U27427 (N_27427,N_24408,N_20188);
or U27428 (N_27428,N_22636,N_20689);
and U27429 (N_27429,N_23009,N_20499);
nand U27430 (N_27430,N_23654,N_20164);
xor U27431 (N_27431,N_24115,N_23975);
nand U27432 (N_27432,N_23883,N_20021);
and U27433 (N_27433,N_21398,N_20809);
or U27434 (N_27434,N_23419,N_23165);
or U27435 (N_27435,N_22902,N_24259);
nand U27436 (N_27436,N_24636,N_22881);
and U27437 (N_27437,N_23721,N_24129);
and U27438 (N_27438,N_21518,N_21828);
nor U27439 (N_27439,N_24336,N_23332);
or U27440 (N_27440,N_23792,N_24158);
and U27441 (N_27441,N_24394,N_22532);
and U27442 (N_27442,N_24852,N_21569);
nand U27443 (N_27443,N_22733,N_21077);
or U27444 (N_27444,N_22356,N_23515);
xnor U27445 (N_27445,N_22742,N_22975);
and U27446 (N_27446,N_24829,N_21438);
nand U27447 (N_27447,N_21285,N_23707);
nor U27448 (N_27448,N_20594,N_24997);
nand U27449 (N_27449,N_22354,N_23825);
or U27450 (N_27450,N_22879,N_22339);
or U27451 (N_27451,N_21622,N_20103);
or U27452 (N_27452,N_24701,N_23126);
or U27453 (N_27453,N_23107,N_22136);
nor U27454 (N_27454,N_23458,N_21421);
nand U27455 (N_27455,N_24087,N_20692);
or U27456 (N_27456,N_24790,N_21262);
nor U27457 (N_27457,N_22418,N_22897);
nand U27458 (N_27458,N_20657,N_22023);
xnor U27459 (N_27459,N_22835,N_20211);
and U27460 (N_27460,N_24571,N_20131);
nand U27461 (N_27461,N_20863,N_21839);
nand U27462 (N_27462,N_23294,N_20723);
nand U27463 (N_27463,N_23486,N_21762);
xor U27464 (N_27464,N_21813,N_21703);
nor U27465 (N_27465,N_20511,N_24066);
nor U27466 (N_27466,N_24486,N_20902);
xor U27467 (N_27467,N_24381,N_20342);
nand U27468 (N_27468,N_21372,N_23149);
or U27469 (N_27469,N_23029,N_22771);
nand U27470 (N_27470,N_20770,N_24283);
or U27471 (N_27471,N_20667,N_22672);
xor U27472 (N_27472,N_21497,N_24779);
nor U27473 (N_27473,N_20954,N_20115);
nand U27474 (N_27474,N_22302,N_22321);
or U27475 (N_27475,N_21431,N_21955);
or U27476 (N_27476,N_23474,N_21981);
nor U27477 (N_27477,N_24275,N_22314);
nand U27478 (N_27478,N_24363,N_21393);
nand U27479 (N_27479,N_24458,N_21007);
or U27480 (N_27480,N_23527,N_20535);
nor U27481 (N_27481,N_22692,N_21404);
nand U27482 (N_27482,N_22081,N_22598);
nand U27483 (N_27483,N_22295,N_21671);
or U27484 (N_27484,N_23234,N_24702);
xor U27485 (N_27485,N_22514,N_23320);
nor U27486 (N_27486,N_24433,N_21538);
or U27487 (N_27487,N_22335,N_20165);
nor U27488 (N_27488,N_23405,N_20316);
nor U27489 (N_27489,N_24006,N_21207);
nor U27490 (N_27490,N_21330,N_24942);
and U27491 (N_27491,N_23395,N_23342);
and U27492 (N_27492,N_23247,N_23891);
or U27493 (N_27493,N_23208,N_23093);
nand U27494 (N_27494,N_24886,N_24456);
or U27495 (N_27495,N_20996,N_23754);
nand U27496 (N_27496,N_22300,N_21800);
nor U27497 (N_27497,N_23275,N_21915);
nand U27498 (N_27498,N_23307,N_20670);
and U27499 (N_27499,N_23397,N_21978);
nand U27500 (N_27500,N_23902,N_21104);
nand U27501 (N_27501,N_20508,N_24109);
and U27502 (N_27502,N_21039,N_21705);
and U27503 (N_27503,N_24192,N_20613);
nor U27504 (N_27504,N_23419,N_22959);
nand U27505 (N_27505,N_23145,N_22197);
nand U27506 (N_27506,N_23288,N_24055);
and U27507 (N_27507,N_24557,N_21960);
and U27508 (N_27508,N_22734,N_21500);
nor U27509 (N_27509,N_24533,N_23124);
and U27510 (N_27510,N_24125,N_20510);
nand U27511 (N_27511,N_23055,N_23293);
nor U27512 (N_27512,N_20308,N_20902);
nand U27513 (N_27513,N_22567,N_21816);
nor U27514 (N_27514,N_22523,N_23810);
or U27515 (N_27515,N_20413,N_23202);
nor U27516 (N_27516,N_22269,N_22012);
nor U27517 (N_27517,N_21100,N_21012);
and U27518 (N_27518,N_22489,N_23363);
and U27519 (N_27519,N_23652,N_22146);
nand U27520 (N_27520,N_20018,N_22100);
nor U27521 (N_27521,N_22487,N_23833);
xnor U27522 (N_27522,N_22724,N_23874);
or U27523 (N_27523,N_20291,N_24877);
and U27524 (N_27524,N_23303,N_21069);
nor U27525 (N_27525,N_21915,N_24951);
or U27526 (N_27526,N_20108,N_24638);
nor U27527 (N_27527,N_22968,N_24802);
nand U27528 (N_27528,N_22885,N_23990);
xor U27529 (N_27529,N_21862,N_24215);
and U27530 (N_27530,N_20540,N_24829);
and U27531 (N_27531,N_22695,N_23578);
xor U27532 (N_27532,N_21936,N_23824);
nand U27533 (N_27533,N_21415,N_21153);
nand U27534 (N_27534,N_24717,N_20117);
and U27535 (N_27535,N_20205,N_21573);
or U27536 (N_27536,N_20783,N_22848);
and U27537 (N_27537,N_23992,N_21714);
or U27538 (N_27538,N_20171,N_22891);
nand U27539 (N_27539,N_22883,N_23529);
or U27540 (N_27540,N_23968,N_24939);
and U27541 (N_27541,N_22350,N_21366);
nand U27542 (N_27542,N_22869,N_23164);
nor U27543 (N_27543,N_22659,N_24886);
xor U27544 (N_27544,N_20713,N_22604);
nor U27545 (N_27545,N_22670,N_24959);
and U27546 (N_27546,N_20192,N_20378);
nand U27547 (N_27547,N_24610,N_21214);
nand U27548 (N_27548,N_20515,N_24346);
nor U27549 (N_27549,N_22856,N_24229);
nand U27550 (N_27550,N_24024,N_24712);
xor U27551 (N_27551,N_20190,N_21573);
or U27552 (N_27552,N_24096,N_21927);
or U27553 (N_27553,N_22496,N_24159);
nand U27554 (N_27554,N_23262,N_20832);
nand U27555 (N_27555,N_21447,N_20833);
and U27556 (N_27556,N_22688,N_20060);
nor U27557 (N_27557,N_23751,N_24943);
and U27558 (N_27558,N_24885,N_21604);
and U27559 (N_27559,N_22462,N_21513);
nor U27560 (N_27560,N_20300,N_21928);
nand U27561 (N_27561,N_21690,N_22284);
nand U27562 (N_27562,N_22449,N_23326);
nand U27563 (N_27563,N_21331,N_21185);
nor U27564 (N_27564,N_23414,N_20868);
nand U27565 (N_27565,N_22515,N_24136);
or U27566 (N_27566,N_20637,N_22462);
and U27567 (N_27567,N_22772,N_20534);
and U27568 (N_27568,N_23440,N_21848);
and U27569 (N_27569,N_24576,N_21604);
nand U27570 (N_27570,N_21538,N_23061);
xnor U27571 (N_27571,N_21056,N_21231);
and U27572 (N_27572,N_22007,N_21988);
and U27573 (N_27573,N_22299,N_20540);
nand U27574 (N_27574,N_20966,N_24505);
nor U27575 (N_27575,N_23663,N_20983);
or U27576 (N_27576,N_21459,N_23455);
nand U27577 (N_27577,N_24639,N_20860);
nor U27578 (N_27578,N_20268,N_22661);
nand U27579 (N_27579,N_21432,N_20813);
nor U27580 (N_27580,N_22774,N_20543);
nor U27581 (N_27581,N_21133,N_24234);
and U27582 (N_27582,N_21808,N_24865);
or U27583 (N_27583,N_21303,N_22389);
or U27584 (N_27584,N_20135,N_20351);
and U27585 (N_27585,N_24377,N_23279);
xor U27586 (N_27586,N_22513,N_24731);
nand U27587 (N_27587,N_24707,N_20092);
xnor U27588 (N_27588,N_24117,N_21235);
or U27589 (N_27589,N_21705,N_22117);
or U27590 (N_27590,N_23418,N_24836);
or U27591 (N_27591,N_23603,N_23006);
nand U27592 (N_27592,N_24768,N_24484);
or U27593 (N_27593,N_20096,N_23472);
and U27594 (N_27594,N_24695,N_20060);
nor U27595 (N_27595,N_24792,N_20296);
nand U27596 (N_27596,N_24420,N_23948);
or U27597 (N_27597,N_22771,N_21464);
nand U27598 (N_27598,N_22634,N_23965);
and U27599 (N_27599,N_22011,N_23836);
and U27600 (N_27600,N_21433,N_20176);
and U27601 (N_27601,N_23542,N_22114);
xnor U27602 (N_27602,N_21994,N_24474);
or U27603 (N_27603,N_22667,N_22692);
or U27604 (N_27604,N_20053,N_23687);
and U27605 (N_27605,N_20300,N_22971);
nand U27606 (N_27606,N_20424,N_24218);
and U27607 (N_27607,N_20384,N_21919);
or U27608 (N_27608,N_21094,N_23019);
nand U27609 (N_27609,N_20528,N_21296);
or U27610 (N_27610,N_21529,N_21371);
xnor U27611 (N_27611,N_21433,N_21983);
and U27612 (N_27612,N_21532,N_21802);
and U27613 (N_27613,N_20203,N_20985);
and U27614 (N_27614,N_23475,N_22690);
nand U27615 (N_27615,N_20442,N_23934);
and U27616 (N_27616,N_21460,N_21387);
nand U27617 (N_27617,N_20195,N_22132);
or U27618 (N_27618,N_20328,N_20146);
and U27619 (N_27619,N_22901,N_24795);
and U27620 (N_27620,N_23278,N_22091);
and U27621 (N_27621,N_22361,N_20085);
and U27622 (N_27622,N_24940,N_21007);
nor U27623 (N_27623,N_24518,N_22188);
or U27624 (N_27624,N_21214,N_22605);
xnor U27625 (N_27625,N_21398,N_22638);
or U27626 (N_27626,N_20138,N_21574);
and U27627 (N_27627,N_21771,N_22593);
nor U27628 (N_27628,N_21849,N_22416);
nand U27629 (N_27629,N_24026,N_21087);
and U27630 (N_27630,N_20030,N_20715);
and U27631 (N_27631,N_20872,N_24341);
nor U27632 (N_27632,N_22994,N_20922);
and U27633 (N_27633,N_24745,N_23937);
xnor U27634 (N_27634,N_24512,N_23168);
xnor U27635 (N_27635,N_20892,N_21568);
nor U27636 (N_27636,N_20990,N_22378);
or U27637 (N_27637,N_24184,N_23695);
nor U27638 (N_27638,N_22394,N_23715);
nand U27639 (N_27639,N_24810,N_23377);
nand U27640 (N_27640,N_22036,N_20744);
and U27641 (N_27641,N_22721,N_24571);
and U27642 (N_27642,N_20473,N_22058);
xnor U27643 (N_27643,N_21737,N_22858);
nor U27644 (N_27644,N_24958,N_20832);
and U27645 (N_27645,N_22546,N_23656);
or U27646 (N_27646,N_24600,N_24571);
nor U27647 (N_27647,N_21183,N_20730);
nand U27648 (N_27648,N_24558,N_22981);
nor U27649 (N_27649,N_20325,N_23032);
nand U27650 (N_27650,N_22466,N_24220);
and U27651 (N_27651,N_20868,N_20490);
and U27652 (N_27652,N_22205,N_22725);
nand U27653 (N_27653,N_24025,N_20576);
and U27654 (N_27654,N_23276,N_21751);
nor U27655 (N_27655,N_21446,N_21595);
and U27656 (N_27656,N_22785,N_23462);
xnor U27657 (N_27657,N_21135,N_22595);
xnor U27658 (N_27658,N_22199,N_22827);
nand U27659 (N_27659,N_20268,N_20498);
and U27660 (N_27660,N_21535,N_24808);
nand U27661 (N_27661,N_23808,N_24481);
nor U27662 (N_27662,N_22597,N_23424);
nor U27663 (N_27663,N_22993,N_20872);
or U27664 (N_27664,N_20448,N_23956);
or U27665 (N_27665,N_23672,N_24040);
nor U27666 (N_27666,N_22413,N_24428);
or U27667 (N_27667,N_23782,N_21070);
nand U27668 (N_27668,N_22363,N_24310);
or U27669 (N_27669,N_22270,N_21159);
and U27670 (N_27670,N_23733,N_21679);
and U27671 (N_27671,N_22120,N_21013);
or U27672 (N_27672,N_24393,N_23818);
xnor U27673 (N_27673,N_21986,N_22459);
nand U27674 (N_27674,N_21207,N_22070);
nand U27675 (N_27675,N_22597,N_22760);
nand U27676 (N_27676,N_24466,N_22807);
nor U27677 (N_27677,N_24686,N_21576);
and U27678 (N_27678,N_23345,N_23619);
or U27679 (N_27679,N_24791,N_21271);
or U27680 (N_27680,N_20553,N_24554);
nand U27681 (N_27681,N_24181,N_22089);
or U27682 (N_27682,N_22589,N_22860);
nor U27683 (N_27683,N_23263,N_20409);
xnor U27684 (N_27684,N_23486,N_22666);
or U27685 (N_27685,N_21398,N_23065);
xor U27686 (N_27686,N_22667,N_22572);
or U27687 (N_27687,N_22231,N_20633);
nor U27688 (N_27688,N_20628,N_22749);
or U27689 (N_27689,N_23701,N_23744);
or U27690 (N_27690,N_22789,N_21686);
or U27691 (N_27691,N_23935,N_24170);
or U27692 (N_27692,N_23723,N_21725);
and U27693 (N_27693,N_21577,N_20197);
nand U27694 (N_27694,N_23662,N_24172);
or U27695 (N_27695,N_20010,N_23333);
and U27696 (N_27696,N_22784,N_22417);
or U27697 (N_27697,N_21396,N_20029);
nand U27698 (N_27698,N_24569,N_22597);
or U27699 (N_27699,N_23432,N_24421);
and U27700 (N_27700,N_20149,N_20493);
nor U27701 (N_27701,N_24489,N_23728);
or U27702 (N_27702,N_20494,N_22239);
or U27703 (N_27703,N_20609,N_21039);
or U27704 (N_27704,N_23040,N_24979);
xnor U27705 (N_27705,N_22839,N_21444);
xor U27706 (N_27706,N_20648,N_21382);
or U27707 (N_27707,N_24297,N_23965);
nand U27708 (N_27708,N_20868,N_20458);
nand U27709 (N_27709,N_24073,N_24751);
and U27710 (N_27710,N_21004,N_24798);
or U27711 (N_27711,N_20125,N_22480);
nand U27712 (N_27712,N_22533,N_23990);
or U27713 (N_27713,N_21811,N_24652);
nor U27714 (N_27714,N_21749,N_22925);
and U27715 (N_27715,N_22836,N_21619);
nand U27716 (N_27716,N_22676,N_22272);
or U27717 (N_27717,N_24753,N_23722);
and U27718 (N_27718,N_24026,N_20922);
nor U27719 (N_27719,N_24275,N_24419);
or U27720 (N_27720,N_23078,N_22541);
and U27721 (N_27721,N_23167,N_23432);
nor U27722 (N_27722,N_23498,N_23061);
or U27723 (N_27723,N_21611,N_22324);
and U27724 (N_27724,N_22372,N_20838);
or U27725 (N_27725,N_24540,N_24837);
xnor U27726 (N_27726,N_22627,N_23834);
or U27727 (N_27727,N_21072,N_22693);
or U27728 (N_27728,N_20942,N_24711);
and U27729 (N_27729,N_20770,N_21957);
or U27730 (N_27730,N_21971,N_23197);
xor U27731 (N_27731,N_22208,N_22177);
xnor U27732 (N_27732,N_20420,N_22242);
or U27733 (N_27733,N_23389,N_20824);
nand U27734 (N_27734,N_23458,N_21109);
nor U27735 (N_27735,N_24049,N_23066);
nand U27736 (N_27736,N_22473,N_21142);
xnor U27737 (N_27737,N_20504,N_24753);
or U27738 (N_27738,N_20308,N_21066);
xor U27739 (N_27739,N_23757,N_21506);
nand U27740 (N_27740,N_22496,N_23187);
and U27741 (N_27741,N_23899,N_21662);
nor U27742 (N_27742,N_23740,N_22390);
nand U27743 (N_27743,N_22677,N_23887);
and U27744 (N_27744,N_21677,N_23868);
nand U27745 (N_27745,N_24962,N_23265);
and U27746 (N_27746,N_20691,N_20797);
nand U27747 (N_27747,N_20854,N_20375);
or U27748 (N_27748,N_21374,N_22421);
and U27749 (N_27749,N_24310,N_21218);
xor U27750 (N_27750,N_22937,N_20775);
nand U27751 (N_27751,N_24471,N_22992);
nand U27752 (N_27752,N_21311,N_23019);
and U27753 (N_27753,N_24179,N_22688);
nor U27754 (N_27754,N_20180,N_23541);
or U27755 (N_27755,N_24304,N_23396);
nand U27756 (N_27756,N_21626,N_22903);
and U27757 (N_27757,N_23541,N_21373);
and U27758 (N_27758,N_24237,N_20895);
or U27759 (N_27759,N_23063,N_22869);
xnor U27760 (N_27760,N_24927,N_24245);
nor U27761 (N_27761,N_20220,N_24474);
nand U27762 (N_27762,N_22947,N_20966);
xnor U27763 (N_27763,N_22457,N_20945);
xnor U27764 (N_27764,N_22942,N_20511);
nand U27765 (N_27765,N_23792,N_22902);
nor U27766 (N_27766,N_20970,N_20955);
and U27767 (N_27767,N_20793,N_20291);
and U27768 (N_27768,N_24421,N_24688);
nand U27769 (N_27769,N_22778,N_20717);
xnor U27770 (N_27770,N_24258,N_23723);
or U27771 (N_27771,N_22278,N_20283);
nand U27772 (N_27772,N_23254,N_22612);
nand U27773 (N_27773,N_23355,N_20597);
and U27774 (N_27774,N_22959,N_24684);
nor U27775 (N_27775,N_21767,N_21221);
xnor U27776 (N_27776,N_21370,N_23695);
nor U27777 (N_27777,N_21045,N_21442);
or U27778 (N_27778,N_24999,N_23157);
nor U27779 (N_27779,N_23551,N_22423);
or U27780 (N_27780,N_23018,N_23956);
or U27781 (N_27781,N_24502,N_22288);
and U27782 (N_27782,N_24363,N_22168);
or U27783 (N_27783,N_22824,N_24681);
nor U27784 (N_27784,N_24156,N_21538);
nor U27785 (N_27785,N_20439,N_20239);
or U27786 (N_27786,N_24679,N_23324);
nor U27787 (N_27787,N_21018,N_23576);
nor U27788 (N_27788,N_23042,N_24682);
nor U27789 (N_27789,N_21561,N_21451);
nor U27790 (N_27790,N_24368,N_23945);
nor U27791 (N_27791,N_22087,N_22338);
and U27792 (N_27792,N_20689,N_20813);
xor U27793 (N_27793,N_23071,N_20249);
xor U27794 (N_27794,N_22498,N_21940);
nor U27795 (N_27795,N_21788,N_23246);
or U27796 (N_27796,N_20110,N_20431);
and U27797 (N_27797,N_24160,N_24631);
nand U27798 (N_27798,N_23588,N_20331);
or U27799 (N_27799,N_22721,N_23195);
and U27800 (N_27800,N_24914,N_22340);
nand U27801 (N_27801,N_24614,N_24991);
nand U27802 (N_27802,N_23400,N_23503);
nand U27803 (N_27803,N_23194,N_20431);
nand U27804 (N_27804,N_21590,N_22955);
xor U27805 (N_27805,N_24079,N_23305);
and U27806 (N_27806,N_22083,N_21479);
nand U27807 (N_27807,N_20980,N_21647);
or U27808 (N_27808,N_24820,N_21948);
or U27809 (N_27809,N_20096,N_24680);
or U27810 (N_27810,N_21083,N_22920);
and U27811 (N_27811,N_20688,N_23112);
nand U27812 (N_27812,N_21798,N_24204);
nor U27813 (N_27813,N_24690,N_24396);
nand U27814 (N_27814,N_22993,N_22086);
and U27815 (N_27815,N_23456,N_21327);
nand U27816 (N_27816,N_24669,N_24017);
and U27817 (N_27817,N_22096,N_21204);
and U27818 (N_27818,N_21650,N_23206);
nor U27819 (N_27819,N_20062,N_24588);
and U27820 (N_27820,N_20088,N_23073);
nor U27821 (N_27821,N_24985,N_22283);
and U27822 (N_27822,N_24491,N_21143);
nor U27823 (N_27823,N_24789,N_22855);
nand U27824 (N_27824,N_24069,N_21590);
xor U27825 (N_27825,N_24484,N_21235);
nor U27826 (N_27826,N_22153,N_23748);
nor U27827 (N_27827,N_23409,N_23461);
and U27828 (N_27828,N_21300,N_23080);
and U27829 (N_27829,N_21851,N_24426);
and U27830 (N_27830,N_20510,N_20560);
xor U27831 (N_27831,N_23728,N_21009);
or U27832 (N_27832,N_24891,N_21900);
nor U27833 (N_27833,N_20432,N_22594);
xor U27834 (N_27834,N_22257,N_23212);
and U27835 (N_27835,N_20859,N_20313);
nor U27836 (N_27836,N_21461,N_24376);
and U27837 (N_27837,N_21750,N_24736);
nand U27838 (N_27838,N_23034,N_22386);
and U27839 (N_27839,N_24372,N_21699);
nor U27840 (N_27840,N_21291,N_21805);
nor U27841 (N_27841,N_24983,N_20220);
or U27842 (N_27842,N_22995,N_20248);
nand U27843 (N_27843,N_22947,N_22650);
and U27844 (N_27844,N_21773,N_24699);
or U27845 (N_27845,N_20647,N_24615);
nor U27846 (N_27846,N_22170,N_23713);
nor U27847 (N_27847,N_23597,N_23085);
and U27848 (N_27848,N_21151,N_23727);
or U27849 (N_27849,N_20714,N_20295);
or U27850 (N_27850,N_20961,N_24938);
nor U27851 (N_27851,N_23776,N_21832);
xor U27852 (N_27852,N_20664,N_24750);
nand U27853 (N_27853,N_24607,N_23121);
nor U27854 (N_27854,N_23350,N_22113);
and U27855 (N_27855,N_24626,N_23515);
xor U27856 (N_27856,N_24301,N_24857);
xor U27857 (N_27857,N_21092,N_22982);
and U27858 (N_27858,N_23532,N_22390);
nor U27859 (N_27859,N_20746,N_20504);
and U27860 (N_27860,N_22292,N_23669);
nor U27861 (N_27861,N_22969,N_23049);
or U27862 (N_27862,N_24422,N_21103);
or U27863 (N_27863,N_23407,N_23479);
and U27864 (N_27864,N_22338,N_21682);
or U27865 (N_27865,N_23109,N_22237);
nand U27866 (N_27866,N_23592,N_20143);
and U27867 (N_27867,N_20451,N_24388);
nor U27868 (N_27868,N_23652,N_23512);
nand U27869 (N_27869,N_21653,N_20629);
and U27870 (N_27870,N_23075,N_22411);
nand U27871 (N_27871,N_21436,N_21486);
nand U27872 (N_27872,N_20908,N_23968);
nand U27873 (N_27873,N_22235,N_23153);
and U27874 (N_27874,N_21884,N_21683);
nand U27875 (N_27875,N_21203,N_21680);
and U27876 (N_27876,N_22632,N_20393);
nor U27877 (N_27877,N_24482,N_21075);
xor U27878 (N_27878,N_22939,N_21488);
nand U27879 (N_27879,N_24709,N_20010);
or U27880 (N_27880,N_20985,N_20969);
xnor U27881 (N_27881,N_20991,N_20062);
or U27882 (N_27882,N_20093,N_22917);
or U27883 (N_27883,N_21062,N_21006);
and U27884 (N_27884,N_24692,N_21504);
nand U27885 (N_27885,N_23055,N_22205);
nor U27886 (N_27886,N_22108,N_24397);
nor U27887 (N_27887,N_21606,N_21392);
xor U27888 (N_27888,N_23618,N_20330);
nor U27889 (N_27889,N_20034,N_20759);
and U27890 (N_27890,N_22603,N_21861);
nor U27891 (N_27891,N_22929,N_21707);
nor U27892 (N_27892,N_20531,N_21690);
xor U27893 (N_27893,N_23378,N_22041);
or U27894 (N_27894,N_24685,N_24968);
or U27895 (N_27895,N_24901,N_24869);
nand U27896 (N_27896,N_21952,N_21992);
nand U27897 (N_27897,N_24401,N_20464);
nand U27898 (N_27898,N_21766,N_23694);
and U27899 (N_27899,N_20427,N_21547);
and U27900 (N_27900,N_23509,N_21264);
and U27901 (N_27901,N_24972,N_22839);
nand U27902 (N_27902,N_20163,N_23878);
and U27903 (N_27903,N_20974,N_22682);
nand U27904 (N_27904,N_24315,N_21391);
nand U27905 (N_27905,N_23627,N_20306);
nor U27906 (N_27906,N_24449,N_20457);
nand U27907 (N_27907,N_22173,N_24948);
and U27908 (N_27908,N_20638,N_21477);
and U27909 (N_27909,N_21261,N_23692);
or U27910 (N_27910,N_20613,N_23923);
or U27911 (N_27911,N_23911,N_20839);
nor U27912 (N_27912,N_23982,N_24671);
xnor U27913 (N_27913,N_22529,N_22597);
nand U27914 (N_27914,N_24705,N_24866);
xor U27915 (N_27915,N_23232,N_23774);
or U27916 (N_27916,N_21970,N_21666);
nand U27917 (N_27917,N_24105,N_20514);
nor U27918 (N_27918,N_20224,N_21694);
nor U27919 (N_27919,N_22626,N_22566);
nor U27920 (N_27920,N_22484,N_20039);
xor U27921 (N_27921,N_24346,N_22269);
and U27922 (N_27922,N_23409,N_24380);
or U27923 (N_27923,N_21745,N_21342);
nand U27924 (N_27924,N_21694,N_20229);
and U27925 (N_27925,N_23759,N_22056);
nor U27926 (N_27926,N_22462,N_21006);
nand U27927 (N_27927,N_24491,N_20638);
and U27928 (N_27928,N_20472,N_20513);
nand U27929 (N_27929,N_20052,N_20715);
and U27930 (N_27930,N_23553,N_22735);
or U27931 (N_27931,N_24120,N_23956);
or U27932 (N_27932,N_21842,N_21311);
nor U27933 (N_27933,N_20410,N_22272);
xnor U27934 (N_27934,N_24797,N_22425);
or U27935 (N_27935,N_21130,N_24921);
nand U27936 (N_27936,N_22461,N_21886);
and U27937 (N_27937,N_22529,N_20048);
or U27938 (N_27938,N_24714,N_21571);
nor U27939 (N_27939,N_22538,N_20918);
nor U27940 (N_27940,N_22685,N_22560);
nand U27941 (N_27941,N_23265,N_21359);
nand U27942 (N_27942,N_22277,N_24482);
and U27943 (N_27943,N_21265,N_22416);
nor U27944 (N_27944,N_23381,N_22310);
or U27945 (N_27945,N_23957,N_20070);
or U27946 (N_27946,N_22240,N_24985);
and U27947 (N_27947,N_20070,N_22045);
nand U27948 (N_27948,N_20339,N_23066);
and U27949 (N_27949,N_21414,N_24809);
and U27950 (N_27950,N_24778,N_23865);
or U27951 (N_27951,N_20316,N_20752);
nand U27952 (N_27952,N_24731,N_21054);
xnor U27953 (N_27953,N_20784,N_20463);
and U27954 (N_27954,N_23926,N_22262);
and U27955 (N_27955,N_21632,N_20023);
nand U27956 (N_27956,N_20246,N_21013);
and U27957 (N_27957,N_20823,N_24463);
nand U27958 (N_27958,N_21030,N_23517);
or U27959 (N_27959,N_23031,N_24898);
and U27960 (N_27960,N_22976,N_24300);
nor U27961 (N_27961,N_22538,N_23743);
xnor U27962 (N_27962,N_24615,N_20661);
nor U27963 (N_27963,N_21981,N_21240);
nor U27964 (N_27964,N_21132,N_22409);
nand U27965 (N_27965,N_22986,N_24622);
or U27966 (N_27966,N_24133,N_23237);
or U27967 (N_27967,N_21145,N_20166);
and U27968 (N_27968,N_23601,N_20745);
nand U27969 (N_27969,N_21374,N_21182);
or U27970 (N_27970,N_20597,N_24137);
or U27971 (N_27971,N_20447,N_24354);
nor U27972 (N_27972,N_21047,N_22889);
xnor U27973 (N_27973,N_22148,N_21562);
nor U27974 (N_27974,N_24417,N_20896);
nand U27975 (N_27975,N_22246,N_20346);
and U27976 (N_27976,N_24461,N_22720);
nor U27977 (N_27977,N_20413,N_23451);
and U27978 (N_27978,N_23253,N_24204);
and U27979 (N_27979,N_23850,N_24759);
and U27980 (N_27980,N_24030,N_21416);
or U27981 (N_27981,N_22655,N_24101);
nor U27982 (N_27982,N_21361,N_20936);
xnor U27983 (N_27983,N_23135,N_24057);
or U27984 (N_27984,N_21690,N_20912);
nand U27985 (N_27985,N_21497,N_20042);
xor U27986 (N_27986,N_21521,N_22390);
nand U27987 (N_27987,N_23876,N_22305);
and U27988 (N_27988,N_20716,N_22344);
nor U27989 (N_27989,N_24963,N_21465);
or U27990 (N_27990,N_20837,N_22717);
or U27991 (N_27991,N_21206,N_22700);
or U27992 (N_27992,N_22562,N_22939);
or U27993 (N_27993,N_21455,N_20038);
and U27994 (N_27994,N_23203,N_21771);
and U27995 (N_27995,N_21482,N_20848);
or U27996 (N_27996,N_23230,N_24571);
nand U27997 (N_27997,N_23683,N_20667);
nor U27998 (N_27998,N_24297,N_23307);
or U27999 (N_27999,N_24123,N_21133);
nor U28000 (N_28000,N_20049,N_20684);
xnor U28001 (N_28001,N_21066,N_23968);
nand U28002 (N_28002,N_24455,N_22475);
or U28003 (N_28003,N_23685,N_20881);
xnor U28004 (N_28004,N_24540,N_20901);
and U28005 (N_28005,N_22281,N_23463);
nor U28006 (N_28006,N_20449,N_22489);
xor U28007 (N_28007,N_24000,N_21135);
nor U28008 (N_28008,N_24140,N_24173);
and U28009 (N_28009,N_20246,N_23812);
nor U28010 (N_28010,N_21260,N_20342);
nand U28011 (N_28011,N_20932,N_23836);
or U28012 (N_28012,N_21732,N_24420);
xnor U28013 (N_28013,N_21348,N_23623);
and U28014 (N_28014,N_21347,N_24569);
nor U28015 (N_28015,N_24183,N_24771);
or U28016 (N_28016,N_22883,N_22479);
nor U28017 (N_28017,N_22237,N_23781);
nand U28018 (N_28018,N_22393,N_24087);
and U28019 (N_28019,N_23009,N_23780);
and U28020 (N_28020,N_22962,N_20695);
and U28021 (N_28021,N_23266,N_24935);
nor U28022 (N_28022,N_23390,N_24907);
xor U28023 (N_28023,N_21417,N_21776);
nor U28024 (N_28024,N_24726,N_23268);
xnor U28025 (N_28025,N_23036,N_23478);
nor U28026 (N_28026,N_22736,N_21195);
nor U28027 (N_28027,N_24956,N_24145);
nor U28028 (N_28028,N_23134,N_23833);
nor U28029 (N_28029,N_22845,N_20862);
nand U28030 (N_28030,N_24795,N_24004);
nor U28031 (N_28031,N_23580,N_22490);
nand U28032 (N_28032,N_20885,N_24342);
nand U28033 (N_28033,N_23832,N_24188);
and U28034 (N_28034,N_23871,N_20414);
nand U28035 (N_28035,N_21430,N_21556);
nor U28036 (N_28036,N_23180,N_24827);
nor U28037 (N_28037,N_23283,N_23855);
and U28038 (N_28038,N_20171,N_21875);
and U28039 (N_28039,N_20471,N_24430);
nand U28040 (N_28040,N_21700,N_22047);
or U28041 (N_28041,N_21828,N_24477);
or U28042 (N_28042,N_23331,N_20326);
nor U28043 (N_28043,N_22142,N_21157);
nand U28044 (N_28044,N_21288,N_24636);
and U28045 (N_28045,N_20691,N_20688);
nand U28046 (N_28046,N_23585,N_21754);
or U28047 (N_28047,N_24190,N_23400);
and U28048 (N_28048,N_21763,N_21145);
and U28049 (N_28049,N_22373,N_22655);
and U28050 (N_28050,N_21002,N_24840);
nand U28051 (N_28051,N_22678,N_20409);
and U28052 (N_28052,N_22450,N_21637);
nand U28053 (N_28053,N_21598,N_22523);
nand U28054 (N_28054,N_22838,N_20313);
and U28055 (N_28055,N_21850,N_22991);
xnor U28056 (N_28056,N_23522,N_24890);
nand U28057 (N_28057,N_24721,N_23925);
nor U28058 (N_28058,N_24944,N_24069);
and U28059 (N_28059,N_22941,N_20905);
nor U28060 (N_28060,N_21433,N_23370);
or U28061 (N_28061,N_22749,N_23595);
nor U28062 (N_28062,N_23102,N_21187);
nand U28063 (N_28063,N_23060,N_21255);
nor U28064 (N_28064,N_23282,N_20232);
nor U28065 (N_28065,N_24359,N_22087);
and U28066 (N_28066,N_23856,N_24688);
nand U28067 (N_28067,N_21450,N_23728);
nor U28068 (N_28068,N_23677,N_21968);
nor U28069 (N_28069,N_23590,N_23133);
and U28070 (N_28070,N_23073,N_22133);
nand U28071 (N_28071,N_20119,N_22256);
nand U28072 (N_28072,N_23746,N_20817);
or U28073 (N_28073,N_20363,N_20729);
nand U28074 (N_28074,N_24969,N_22049);
nor U28075 (N_28075,N_24109,N_24471);
nand U28076 (N_28076,N_20245,N_22430);
nand U28077 (N_28077,N_24119,N_23564);
or U28078 (N_28078,N_21833,N_23564);
nor U28079 (N_28079,N_22219,N_20898);
nor U28080 (N_28080,N_20427,N_20731);
nor U28081 (N_28081,N_21471,N_22790);
nand U28082 (N_28082,N_24258,N_21985);
nor U28083 (N_28083,N_22061,N_21366);
nand U28084 (N_28084,N_20426,N_20564);
nor U28085 (N_28085,N_23644,N_24815);
or U28086 (N_28086,N_22576,N_20690);
nand U28087 (N_28087,N_24181,N_23610);
nand U28088 (N_28088,N_24230,N_24821);
or U28089 (N_28089,N_22565,N_24045);
or U28090 (N_28090,N_24877,N_24619);
nor U28091 (N_28091,N_22340,N_20532);
nand U28092 (N_28092,N_22407,N_20242);
and U28093 (N_28093,N_24388,N_20596);
or U28094 (N_28094,N_20068,N_23633);
or U28095 (N_28095,N_21342,N_21999);
and U28096 (N_28096,N_21073,N_23787);
and U28097 (N_28097,N_22112,N_21761);
and U28098 (N_28098,N_20559,N_20644);
nand U28099 (N_28099,N_20218,N_24427);
and U28100 (N_28100,N_24150,N_21436);
and U28101 (N_28101,N_22179,N_21494);
and U28102 (N_28102,N_20683,N_23494);
and U28103 (N_28103,N_23127,N_23742);
and U28104 (N_28104,N_21626,N_23505);
nor U28105 (N_28105,N_24021,N_24790);
nor U28106 (N_28106,N_23415,N_21245);
nor U28107 (N_28107,N_23477,N_21633);
nor U28108 (N_28108,N_24734,N_22213);
nor U28109 (N_28109,N_20876,N_24816);
xnor U28110 (N_28110,N_22815,N_20793);
and U28111 (N_28111,N_21745,N_22404);
nor U28112 (N_28112,N_21226,N_22285);
nor U28113 (N_28113,N_22748,N_20500);
or U28114 (N_28114,N_24360,N_23739);
nand U28115 (N_28115,N_23943,N_24313);
nand U28116 (N_28116,N_24065,N_23957);
nand U28117 (N_28117,N_24817,N_22562);
nor U28118 (N_28118,N_23131,N_20436);
and U28119 (N_28119,N_24255,N_24041);
nand U28120 (N_28120,N_23698,N_24598);
nor U28121 (N_28121,N_24748,N_21798);
xnor U28122 (N_28122,N_23756,N_23331);
and U28123 (N_28123,N_21525,N_24332);
or U28124 (N_28124,N_20885,N_23772);
xor U28125 (N_28125,N_24398,N_22518);
nor U28126 (N_28126,N_22450,N_22207);
and U28127 (N_28127,N_23449,N_23862);
nand U28128 (N_28128,N_24169,N_21874);
nand U28129 (N_28129,N_20362,N_24507);
nand U28130 (N_28130,N_24494,N_20774);
and U28131 (N_28131,N_24406,N_22870);
nand U28132 (N_28132,N_24040,N_24395);
or U28133 (N_28133,N_21876,N_23139);
xor U28134 (N_28134,N_24327,N_24190);
nor U28135 (N_28135,N_22952,N_22869);
nor U28136 (N_28136,N_23832,N_21353);
nor U28137 (N_28137,N_24799,N_23392);
and U28138 (N_28138,N_24950,N_20896);
nor U28139 (N_28139,N_22103,N_22206);
or U28140 (N_28140,N_23538,N_20229);
nor U28141 (N_28141,N_20715,N_22770);
nand U28142 (N_28142,N_21198,N_23024);
and U28143 (N_28143,N_21587,N_22201);
nor U28144 (N_28144,N_22546,N_24863);
and U28145 (N_28145,N_24404,N_22468);
nor U28146 (N_28146,N_23030,N_22416);
and U28147 (N_28147,N_22056,N_20048);
nor U28148 (N_28148,N_23714,N_23884);
nor U28149 (N_28149,N_22404,N_24498);
nand U28150 (N_28150,N_22877,N_20851);
or U28151 (N_28151,N_24736,N_22648);
nand U28152 (N_28152,N_20149,N_22738);
nor U28153 (N_28153,N_21344,N_21983);
nor U28154 (N_28154,N_20041,N_24524);
nand U28155 (N_28155,N_23318,N_22801);
or U28156 (N_28156,N_20969,N_22465);
nand U28157 (N_28157,N_22288,N_24501);
or U28158 (N_28158,N_22688,N_24404);
nand U28159 (N_28159,N_20483,N_21566);
and U28160 (N_28160,N_20794,N_22997);
nand U28161 (N_28161,N_24126,N_20740);
nor U28162 (N_28162,N_23533,N_20052);
or U28163 (N_28163,N_22221,N_24796);
or U28164 (N_28164,N_23986,N_24235);
xnor U28165 (N_28165,N_21887,N_24410);
or U28166 (N_28166,N_20703,N_20226);
or U28167 (N_28167,N_22939,N_22883);
or U28168 (N_28168,N_20973,N_22584);
nand U28169 (N_28169,N_20269,N_23213);
and U28170 (N_28170,N_20517,N_23225);
nand U28171 (N_28171,N_23352,N_23670);
nor U28172 (N_28172,N_22703,N_22513);
nand U28173 (N_28173,N_21125,N_23906);
or U28174 (N_28174,N_21208,N_21062);
nand U28175 (N_28175,N_23948,N_23898);
or U28176 (N_28176,N_22620,N_20661);
nor U28177 (N_28177,N_24696,N_20068);
or U28178 (N_28178,N_24404,N_24288);
and U28179 (N_28179,N_21471,N_23680);
xor U28180 (N_28180,N_21612,N_21402);
nand U28181 (N_28181,N_20002,N_20593);
and U28182 (N_28182,N_20167,N_20040);
and U28183 (N_28183,N_20588,N_21845);
and U28184 (N_28184,N_21729,N_23446);
or U28185 (N_28185,N_20133,N_22835);
nor U28186 (N_28186,N_22510,N_21977);
and U28187 (N_28187,N_24188,N_21886);
or U28188 (N_28188,N_20187,N_23585);
nor U28189 (N_28189,N_21259,N_23581);
nor U28190 (N_28190,N_20776,N_21726);
nand U28191 (N_28191,N_24604,N_20247);
or U28192 (N_28192,N_24494,N_20502);
or U28193 (N_28193,N_22524,N_20317);
nand U28194 (N_28194,N_24573,N_24472);
and U28195 (N_28195,N_22748,N_23167);
xnor U28196 (N_28196,N_24572,N_22904);
nand U28197 (N_28197,N_21959,N_24515);
and U28198 (N_28198,N_21594,N_20585);
and U28199 (N_28199,N_20398,N_24985);
nand U28200 (N_28200,N_21147,N_22555);
nor U28201 (N_28201,N_24378,N_22811);
and U28202 (N_28202,N_21540,N_24764);
or U28203 (N_28203,N_20948,N_24362);
xnor U28204 (N_28204,N_21402,N_22995);
and U28205 (N_28205,N_20683,N_21829);
nor U28206 (N_28206,N_23598,N_20277);
nor U28207 (N_28207,N_22659,N_23042);
or U28208 (N_28208,N_22583,N_23851);
xor U28209 (N_28209,N_23436,N_24863);
or U28210 (N_28210,N_24580,N_23898);
and U28211 (N_28211,N_21524,N_22891);
or U28212 (N_28212,N_22027,N_20725);
xnor U28213 (N_28213,N_21409,N_21535);
xnor U28214 (N_28214,N_21901,N_23640);
nand U28215 (N_28215,N_22265,N_20847);
or U28216 (N_28216,N_24112,N_24825);
nor U28217 (N_28217,N_20046,N_20610);
nor U28218 (N_28218,N_24188,N_23328);
xnor U28219 (N_28219,N_20837,N_20353);
nand U28220 (N_28220,N_20483,N_24724);
nor U28221 (N_28221,N_20852,N_23033);
nand U28222 (N_28222,N_23202,N_23287);
nand U28223 (N_28223,N_23174,N_20609);
xor U28224 (N_28224,N_23397,N_23898);
or U28225 (N_28225,N_21050,N_21670);
or U28226 (N_28226,N_22204,N_20970);
and U28227 (N_28227,N_20930,N_22535);
or U28228 (N_28228,N_22920,N_23977);
nand U28229 (N_28229,N_23794,N_20423);
nor U28230 (N_28230,N_23373,N_24157);
or U28231 (N_28231,N_20503,N_23739);
nand U28232 (N_28232,N_24725,N_21812);
nor U28233 (N_28233,N_22482,N_23806);
nand U28234 (N_28234,N_24452,N_24979);
nor U28235 (N_28235,N_24293,N_23609);
nand U28236 (N_28236,N_23250,N_24591);
nand U28237 (N_28237,N_21039,N_24227);
or U28238 (N_28238,N_21792,N_21644);
and U28239 (N_28239,N_22515,N_21050);
nand U28240 (N_28240,N_22010,N_21099);
or U28241 (N_28241,N_20179,N_20494);
and U28242 (N_28242,N_22632,N_24475);
or U28243 (N_28243,N_24879,N_23050);
nor U28244 (N_28244,N_20643,N_24559);
nor U28245 (N_28245,N_23200,N_22589);
or U28246 (N_28246,N_21970,N_24018);
nand U28247 (N_28247,N_21699,N_22056);
xnor U28248 (N_28248,N_22122,N_20755);
and U28249 (N_28249,N_24412,N_22651);
nand U28250 (N_28250,N_24984,N_24126);
nor U28251 (N_28251,N_22351,N_24484);
nand U28252 (N_28252,N_20637,N_24353);
or U28253 (N_28253,N_21502,N_20249);
nor U28254 (N_28254,N_21016,N_23410);
nor U28255 (N_28255,N_23451,N_22936);
or U28256 (N_28256,N_23819,N_22630);
or U28257 (N_28257,N_20035,N_20760);
and U28258 (N_28258,N_23137,N_21753);
nand U28259 (N_28259,N_22547,N_23578);
nor U28260 (N_28260,N_23206,N_22031);
nand U28261 (N_28261,N_22777,N_20648);
nand U28262 (N_28262,N_24652,N_22746);
xnor U28263 (N_28263,N_21938,N_22222);
nand U28264 (N_28264,N_20758,N_21666);
and U28265 (N_28265,N_20721,N_23494);
nor U28266 (N_28266,N_24146,N_21236);
nand U28267 (N_28267,N_21755,N_23724);
nor U28268 (N_28268,N_21371,N_24372);
nand U28269 (N_28269,N_20682,N_24566);
nor U28270 (N_28270,N_20292,N_22877);
nor U28271 (N_28271,N_21211,N_23057);
and U28272 (N_28272,N_23896,N_23793);
nor U28273 (N_28273,N_22238,N_20381);
nor U28274 (N_28274,N_20357,N_24740);
or U28275 (N_28275,N_20840,N_21726);
nor U28276 (N_28276,N_20817,N_20571);
nor U28277 (N_28277,N_23283,N_23140);
nand U28278 (N_28278,N_21683,N_24899);
and U28279 (N_28279,N_24221,N_21705);
nor U28280 (N_28280,N_23224,N_22597);
nand U28281 (N_28281,N_23485,N_20011);
nand U28282 (N_28282,N_24657,N_21155);
and U28283 (N_28283,N_21350,N_23382);
and U28284 (N_28284,N_22076,N_24148);
and U28285 (N_28285,N_21369,N_20546);
or U28286 (N_28286,N_24492,N_21011);
or U28287 (N_28287,N_23576,N_23987);
and U28288 (N_28288,N_21043,N_20489);
xnor U28289 (N_28289,N_21604,N_21280);
and U28290 (N_28290,N_21396,N_24728);
and U28291 (N_28291,N_24712,N_22693);
nor U28292 (N_28292,N_23004,N_24916);
nor U28293 (N_28293,N_20744,N_20607);
and U28294 (N_28294,N_22671,N_24229);
nor U28295 (N_28295,N_24144,N_24917);
nand U28296 (N_28296,N_21737,N_23893);
xor U28297 (N_28297,N_22132,N_21935);
nor U28298 (N_28298,N_23002,N_23599);
or U28299 (N_28299,N_23630,N_22449);
nor U28300 (N_28300,N_24898,N_23270);
xnor U28301 (N_28301,N_21560,N_21998);
nor U28302 (N_28302,N_21175,N_24914);
nand U28303 (N_28303,N_22255,N_21027);
and U28304 (N_28304,N_23731,N_22175);
xnor U28305 (N_28305,N_20259,N_21152);
or U28306 (N_28306,N_22120,N_22415);
or U28307 (N_28307,N_20365,N_23380);
or U28308 (N_28308,N_20740,N_21701);
nor U28309 (N_28309,N_23308,N_20442);
nor U28310 (N_28310,N_23186,N_20809);
or U28311 (N_28311,N_24582,N_21618);
nand U28312 (N_28312,N_20522,N_21856);
nor U28313 (N_28313,N_21155,N_20649);
nand U28314 (N_28314,N_23555,N_21462);
nor U28315 (N_28315,N_21772,N_24395);
nor U28316 (N_28316,N_20061,N_21862);
nand U28317 (N_28317,N_23030,N_24777);
and U28318 (N_28318,N_23385,N_24251);
xor U28319 (N_28319,N_20713,N_23894);
and U28320 (N_28320,N_20522,N_23630);
and U28321 (N_28321,N_20503,N_20687);
nand U28322 (N_28322,N_22980,N_22054);
nand U28323 (N_28323,N_23909,N_21640);
nand U28324 (N_28324,N_24532,N_23960);
and U28325 (N_28325,N_20382,N_22679);
xor U28326 (N_28326,N_23381,N_24164);
and U28327 (N_28327,N_22841,N_23655);
nand U28328 (N_28328,N_23582,N_23702);
or U28329 (N_28329,N_21362,N_24610);
and U28330 (N_28330,N_24590,N_23436);
nor U28331 (N_28331,N_23308,N_20170);
nand U28332 (N_28332,N_24942,N_24538);
xor U28333 (N_28333,N_23896,N_22603);
nor U28334 (N_28334,N_24048,N_20290);
nand U28335 (N_28335,N_24158,N_21520);
or U28336 (N_28336,N_20916,N_22876);
or U28337 (N_28337,N_22648,N_24725);
or U28338 (N_28338,N_20079,N_20956);
or U28339 (N_28339,N_23399,N_20843);
nand U28340 (N_28340,N_24973,N_20331);
nand U28341 (N_28341,N_22124,N_22434);
nand U28342 (N_28342,N_20468,N_22636);
xor U28343 (N_28343,N_21879,N_22025);
nor U28344 (N_28344,N_22537,N_24004);
nor U28345 (N_28345,N_23349,N_22042);
nand U28346 (N_28346,N_23548,N_20937);
xnor U28347 (N_28347,N_24980,N_22908);
and U28348 (N_28348,N_22983,N_24218);
and U28349 (N_28349,N_21096,N_24063);
nand U28350 (N_28350,N_24403,N_20574);
nor U28351 (N_28351,N_21949,N_20988);
nor U28352 (N_28352,N_20191,N_22064);
nand U28353 (N_28353,N_23372,N_23645);
or U28354 (N_28354,N_23281,N_20007);
nand U28355 (N_28355,N_20940,N_21737);
nand U28356 (N_28356,N_21347,N_20363);
and U28357 (N_28357,N_22532,N_23475);
and U28358 (N_28358,N_20582,N_22102);
nand U28359 (N_28359,N_22583,N_21817);
nor U28360 (N_28360,N_23886,N_23753);
xnor U28361 (N_28361,N_21630,N_24697);
nand U28362 (N_28362,N_23049,N_21264);
nand U28363 (N_28363,N_22482,N_23764);
and U28364 (N_28364,N_20105,N_22691);
and U28365 (N_28365,N_24424,N_23963);
or U28366 (N_28366,N_20486,N_24142);
or U28367 (N_28367,N_22298,N_23593);
and U28368 (N_28368,N_21117,N_24281);
and U28369 (N_28369,N_22863,N_21771);
nand U28370 (N_28370,N_23988,N_21032);
or U28371 (N_28371,N_23119,N_22801);
and U28372 (N_28372,N_20117,N_24167);
and U28373 (N_28373,N_23327,N_22025);
or U28374 (N_28374,N_24041,N_22564);
or U28375 (N_28375,N_22289,N_24920);
and U28376 (N_28376,N_22709,N_22312);
nor U28377 (N_28377,N_20033,N_23245);
or U28378 (N_28378,N_23305,N_22746);
nand U28379 (N_28379,N_24198,N_20407);
nand U28380 (N_28380,N_24177,N_22502);
or U28381 (N_28381,N_20586,N_21899);
and U28382 (N_28382,N_23586,N_21775);
and U28383 (N_28383,N_23741,N_22312);
nor U28384 (N_28384,N_22110,N_20770);
nand U28385 (N_28385,N_22476,N_21286);
or U28386 (N_28386,N_23836,N_22395);
nor U28387 (N_28387,N_21000,N_23918);
or U28388 (N_28388,N_21577,N_22136);
or U28389 (N_28389,N_22103,N_21269);
xnor U28390 (N_28390,N_24968,N_20424);
nor U28391 (N_28391,N_22843,N_21181);
and U28392 (N_28392,N_24370,N_23209);
nand U28393 (N_28393,N_20554,N_20220);
xnor U28394 (N_28394,N_21420,N_22654);
and U28395 (N_28395,N_22688,N_24133);
and U28396 (N_28396,N_21497,N_20605);
or U28397 (N_28397,N_22249,N_21070);
nor U28398 (N_28398,N_20419,N_21074);
xnor U28399 (N_28399,N_24910,N_21830);
or U28400 (N_28400,N_22495,N_22909);
or U28401 (N_28401,N_24532,N_21101);
and U28402 (N_28402,N_22188,N_24204);
nand U28403 (N_28403,N_23039,N_20322);
nor U28404 (N_28404,N_21526,N_24647);
nand U28405 (N_28405,N_22595,N_22472);
xnor U28406 (N_28406,N_21251,N_24187);
nand U28407 (N_28407,N_21898,N_23663);
nand U28408 (N_28408,N_21944,N_23228);
or U28409 (N_28409,N_22614,N_20628);
or U28410 (N_28410,N_20810,N_22157);
nor U28411 (N_28411,N_24975,N_24400);
xnor U28412 (N_28412,N_23244,N_24201);
nor U28413 (N_28413,N_20047,N_20945);
nand U28414 (N_28414,N_20951,N_20445);
xnor U28415 (N_28415,N_23259,N_23997);
nand U28416 (N_28416,N_21576,N_21015);
nand U28417 (N_28417,N_23993,N_23831);
or U28418 (N_28418,N_22707,N_22468);
nand U28419 (N_28419,N_20511,N_20534);
nand U28420 (N_28420,N_20508,N_24099);
or U28421 (N_28421,N_21111,N_22665);
and U28422 (N_28422,N_24192,N_21002);
nand U28423 (N_28423,N_21324,N_20200);
and U28424 (N_28424,N_20303,N_21787);
or U28425 (N_28425,N_23440,N_23275);
and U28426 (N_28426,N_24032,N_21061);
nand U28427 (N_28427,N_22140,N_22723);
or U28428 (N_28428,N_20362,N_21714);
or U28429 (N_28429,N_23011,N_22250);
nand U28430 (N_28430,N_22160,N_20181);
and U28431 (N_28431,N_22110,N_21243);
nand U28432 (N_28432,N_22320,N_20651);
nand U28433 (N_28433,N_23424,N_24459);
nor U28434 (N_28434,N_21863,N_22142);
or U28435 (N_28435,N_20447,N_21868);
and U28436 (N_28436,N_21665,N_23821);
nor U28437 (N_28437,N_24469,N_22659);
or U28438 (N_28438,N_20488,N_21942);
nor U28439 (N_28439,N_21592,N_21395);
nor U28440 (N_28440,N_23938,N_22136);
nand U28441 (N_28441,N_24094,N_23812);
xor U28442 (N_28442,N_24854,N_21437);
nand U28443 (N_28443,N_23498,N_20308);
xnor U28444 (N_28444,N_20638,N_23174);
nor U28445 (N_28445,N_23526,N_21629);
nand U28446 (N_28446,N_21131,N_21562);
and U28447 (N_28447,N_21464,N_24698);
and U28448 (N_28448,N_20753,N_23010);
nand U28449 (N_28449,N_20259,N_24041);
or U28450 (N_28450,N_23926,N_21377);
or U28451 (N_28451,N_21577,N_22216);
nor U28452 (N_28452,N_20392,N_20011);
nor U28453 (N_28453,N_20903,N_22113);
nand U28454 (N_28454,N_23172,N_24716);
and U28455 (N_28455,N_23673,N_20850);
nand U28456 (N_28456,N_20561,N_22367);
nand U28457 (N_28457,N_23954,N_24059);
and U28458 (N_28458,N_23230,N_22707);
nand U28459 (N_28459,N_22781,N_21535);
and U28460 (N_28460,N_21304,N_21891);
and U28461 (N_28461,N_21478,N_24934);
or U28462 (N_28462,N_23447,N_20497);
nor U28463 (N_28463,N_23559,N_21266);
nor U28464 (N_28464,N_22117,N_24528);
xnor U28465 (N_28465,N_20219,N_24053);
xor U28466 (N_28466,N_20552,N_20413);
nand U28467 (N_28467,N_21283,N_22188);
nor U28468 (N_28468,N_23311,N_22611);
nor U28469 (N_28469,N_23827,N_24883);
and U28470 (N_28470,N_24982,N_21810);
nand U28471 (N_28471,N_22444,N_21894);
nand U28472 (N_28472,N_21985,N_22985);
and U28473 (N_28473,N_24578,N_20496);
xnor U28474 (N_28474,N_23003,N_21750);
nand U28475 (N_28475,N_24236,N_21207);
or U28476 (N_28476,N_20989,N_23270);
and U28477 (N_28477,N_24742,N_24466);
nor U28478 (N_28478,N_23517,N_24109);
or U28479 (N_28479,N_20724,N_23125);
or U28480 (N_28480,N_22867,N_20845);
nand U28481 (N_28481,N_24785,N_24121);
and U28482 (N_28482,N_24261,N_21663);
or U28483 (N_28483,N_23773,N_22072);
nor U28484 (N_28484,N_24415,N_24398);
nand U28485 (N_28485,N_24863,N_21170);
and U28486 (N_28486,N_21044,N_21631);
nor U28487 (N_28487,N_23233,N_20567);
nor U28488 (N_28488,N_20579,N_21607);
or U28489 (N_28489,N_24743,N_20855);
and U28490 (N_28490,N_24869,N_22403);
nand U28491 (N_28491,N_22342,N_22629);
or U28492 (N_28492,N_23601,N_23287);
and U28493 (N_28493,N_21230,N_20144);
nor U28494 (N_28494,N_23860,N_22764);
xnor U28495 (N_28495,N_22912,N_22560);
nand U28496 (N_28496,N_21678,N_20934);
xor U28497 (N_28497,N_21171,N_24459);
xnor U28498 (N_28498,N_23657,N_22138);
xnor U28499 (N_28499,N_24093,N_20197);
or U28500 (N_28500,N_20607,N_22691);
nor U28501 (N_28501,N_20652,N_20671);
nor U28502 (N_28502,N_23977,N_23985);
nand U28503 (N_28503,N_21848,N_21802);
or U28504 (N_28504,N_23211,N_22326);
nand U28505 (N_28505,N_22691,N_21694);
nor U28506 (N_28506,N_22059,N_23628);
or U28507 (N_28507,N_22403,N_24965);
xnor U28508 (N_28508,N_20772,N_23429);
xnor U28509 (N_28509,N_22642,N_23926);
nand U28510 (N_28510,N_23842,N_20044);
nand U28511 (N_28511,N_24861,N_22898);
nand U28512 (N_28512,N_21941,N_22500);
nor U28513 (N_28513,N_23476,N_21698);
or U28514 (N_28514,N_21757,N_22598);
nand U28515 (N_28515,N_20382,N_20977);
nor U28516 (N_28516,N_23960,N_24015);
nor U28517 (N_28517,N_21146,N_21077);
nor U28518 (N_28518,N_23120,N_23952);
nor U28519 (N_28519,N_21614,N_21848);
nand U28520 (N_28520,N_23937,N_20526);
or U28521 (N_28521,N_24651,N_22070);
nor U28522 (N_28522,N_23688,N_22803);
xor U28523 (N_28523,N_20706,N_20963);
nor U28524 (N_28524,N_21115,N_23737);
nand U28525 (N_28525,N_22118,N_22232);
nand U28526 (N_28526,N_23566,N_20315);
and U28527 (N_28527,N_24656,N_22763);
and U28528 (N_28528,N_23813,N_20492);
or U28529 (N_28529,N_21121,N_21950);
or U28530 (N_28530,N_22352,N_23386);
nand U28531 (N_28531,N_24283,N_22152);
xnor U28532 (N_28532,N_23805,N_23788);
nor U28533 (N_28533,N_22090,N_23964);
and U28534 (N_28534,N_23448,N_22002);
nor U28535 (N_28535,N_23902,N_24692);
nor U28536 (N_28536,N_20183,N_22686);
nor U28537 (N_28537,N_23831,N_23779);
nor U28538 (N_28538,N_22761,N_24531);
nand U28539 (N_28539,N_20346,N_24899);
and U28540 (N_28540,N_21708,N_23119);
nand U28541 (N_28541,N_23307,N_22103);
and U28542 (N_28542,N_22664,N_20083);
or U28543 (N_28543,N_24950,N_22344);
nand U28544 (N_28544,N_23529,N_24749);
or U28545 (N_28545,N_22550,N_22600);
nor U28546 (N_28546,N_22977,N_24444);
or U28547 (N_28547,N_24355,N_22699);
or U28548 (N_28548,N_21893,N_21863);
or U28549 (N_28549,N_22798,N_20499);
or U28550 (N_28550,N_20713,N_23926);
xnor U28551 (N_28551,N_21527,N_21295);
nor U28552 (N_28552,N_23517,N_22534);
and U28553 (N_28553,N_22965,N_24365);
xnor U28554 (N_28554,N_24214,N_24837);
or U28555 (N_28555,N_23421,N_20996);
and U28556 (N_28556,N_21061,N_20273);
nand U28557 (N_28557,N_21655,N_24965);
nor U28558 (N_28558,N_21750,N_22487);
and U28559 (N_28559,N_24106,N_22953);
nor U28560 (N_28560,N_21051,N_24838);
nor U28561 (N_28561,N_21800,N_22075);
nor U28562 (N_28562,N_21901,N_22894);
nor U28563 (N_28563,N_23175,N_21646);
nor U28564 (N_28564,N_24502,N_20064);
nor U28565 (N_28565,N_21099,N_20679);
nor U28566 (N_28566,N_22177,N_22866);
and U28567 (N_28567,N_24742,N_24814);
and U28568 (N_28568,N_22753,N_22617);
nor U28569 (N_28569,N_22682,N_20256);
nor U28570 (N_28570,N_24813,N_20648);
nor U28571 (N_28571,N_23765,N_21383);
nand U28572 (N_28572,N_21105,N_23120);
or U28573 (N_28573,N_20074,N_23948);
and U28574 (N_28574,N_22906,N_22377);
nand U28575 (N_28575,N_24679,N_24063);
nor U28576 (N_28576,N_20882,N_22548);
xor U28577 (N_28577,N_24628,N_23325);
or U28578 (N_28578,N_23835,N_21220);
nand U28579 (N_28579,N_22181,N_23150);
and U28580 (N_28580,N_24965,N_23247);
nor U28581 (N_28581,N_24825,N_22090);
nand U28582 (N_28582,N_20983,N_22724);
or U28583 (N_28583,N_20683,N_22305);
and U28584 (N_28584,N_23277,N_24535);
nand U28585 (N_28585,N_24021,N_24625);
or U28586 (N_28586,N_21652,N_23429);
or U28587 (N_28587,N_23847,N_20125);
nand U28588 (N_28588,N_23986,N_21439);
nand U28589 (N_28589,N_22615,N_20172);
nand U28590 (N_28590,N_20117,N_22327);
and U28591 (N_28591,N_22715,N_20061);
nand U28592 (N_28592,N_21372,N_24107);
and U28593 (N_28593,N_23973,N_23574);
nor U28594 (N_28594,N_20991,N_22735);
nor U28595 (N_28595,N_23769,N_20178);
nand U28596 (N_28596,N_24070,N_21405);
or U28597 (N_28597,N_21084,N_22229);
nand U28598 (N_28598,N_23558,N_22474);
xor U28599 (N_28599,N_21849,N_24260);
nor U28600 (N_28600,N_21624,N_24111);
nor U28601 (N_28601,N_21905,N_24811);
xnor U28602 (N_28602,N_22868,N_22987);
nand U28603 (N_28603,N_23172,N_20137);
and U28604 (N_28604,N_23201,N_21185);
or U28605 (N_28605,N_22893,N_20196);
or U28606 (N_28606,N_24238,N_22959);
or U28607 (N_28607,N_24570,N_21156);
xor U28608 (N_28608,N_20941,N_23678);
xnor U28609 (N_28609,N_23772,N_23770);
nor U28610 (N_28610,N_23195,N_24415);
nand U28611 (N_28611,N_21279,N_24794);
or U28612 (N_28612,N_23426,N_22301);
nand U28613 (N_28613,N_22542,N_20448);
or U28614 (N_28614,N_24757,N_23076);
or U28615 (N_28615,N_20130,N_20996);
nand U28616 (N_28616,N_24293,N_22704);
nor U28617 (N_28617,N_20535,N_22281);
or U28618 (N_28618,N_22048,N_22853);
or U28619 (N_28619,N_24686,N_21398);
nor U28620 (N_28620,N_23502,N_23704);
xor U28621 (N_28621,N_24604,N_24932);
nor U28622 (N_28622,N_20043,N_21442);
xor U28623 (N_28623,N_22100,N_23930);
or U28624 (N_28624,N_24704,N_23789);
and U28625 (N_28625,N_21458,N_21396);
nor U28626 (N_28626,N_20962,N_21911);
or U28627 (N_28627,N_21505,N_21999);
nand U28628 (N_28628,N_24431,N_22370);
or U28629 (N_28629,N_23382,N_20809);
nor U28630 (N_28630,N_23660,N_20408);
and U28631 (N_28631,N_24535,N_22703);
nor U28632 (N_28632,N_22606,N_22600);
nor U28633 (N_28633,N_20261,N_23560);
or U28634 (N_28634,N_23333,N_21071);
or U28635 (N_28635,N_24738,N_24588);
nand U28636 (N_28636,N_21278,N_21146);
nand U28637 (N_28637,N_21625,N_24547);
nand U28638 (N_28638,N_22828,N_22799);
and U28639 (N_28639,N_23763,N_22850);
and U28640 (N_28640,N_20806,N_22912);
nand U28641 (N_28641,N_23124,N_22035);
nand U28642 (N_28642,N_23654,N_23715);
and U28643 (N_28643,N_21677,N_22122);
nand U28644 (N_28644,N_21352,N_23996);
and U28645 (N_28645,N_22317,N_24435);
and U28646 (N_28646,N_24646,N_24629);
or U28647 (N_28647,N_24527,N_24926);
nor U28648 (N_28648,N_21766,N_21866);
nand U28649 (N_28649,N_20691,N_21731);
xnor U28650 (N_28650,N_24873,N_20302);
nand U28651 (N_28651,N_22383,N_21495);
or U28652 (N_28652,N_23214,N_20782);
nor U28653 (N_28653,N_20210,N_21705);
xnor U28654 (N_28654,N_22891,N_20021);
and U28655 (N_28655,N_24192,N_21457);
nor U28656 (N_28656,N_20252,N_24642);
nand U28657 (N_28657,N_24143,N_21532);
or U28658 (N_28658,N_21099,N_24185);
nand U28659 (N_28659,N_23448,N_24256);
and U28660 (N_28660,N_24552,N_23853);
and U28661 (N_28661,N_20692,N_21203);
or U28662 (N_28662,N_24597,N_22130);
nor U28663 (N_28663,N_22368,N_22884);
nor U28664 (N_28664,N_24862,N_22523);
nor U28665 (N_28665,N_22714,N_22021);
nand U28666 (N_28666,N_21417,N_24647);
nand U28667 (N_28667,N_20636,N_22665);
nor U28668 (N_28668,N_24634,N_24279);
or U28669 (N_28669,N_22446,N_21351);
nand U28670 (N_28670,N_21514,N_24287);
nand U28671 (N_28671,N_24692,N_24564);
or U28672 (N_28672,N_22381,N_22137);
and U28673 (N_28673,N_21494,N_21707);
nor U28674 (N_28674,N_20431,N_24850);
nor U28675 (N_28675,N_22883,N_20073);
and U28676 (N_28676,N_21407,N_21749);
nor U28677 (N_28677,N_24925,N_23455);
nand U28678 (N_28678,N_22057,N_23044);
and U28679 (N_28679,N_20028,N_24866);
and U28680 (N_28680,N_21060,N_23415);
nor U28681 (N_28681,N_22415,N_22501);
nor U28682 (N_28682,N_21247,N_21394);
nand U28683 (N_28683,N_23325,N_24477);
or U28684 (N_28684,N_24901,N_21778);
and U28685 (N_28685,N_23962,N_24654);
nor U28686 (N_28686,N_20252,N_21309);
nand U28687 (N_28687,N_22060,N_22114);
nand U28688 (N_28688,N_22304,N_22111);
or U28689 (N_28689,N_22347,N_21455);
nand U28690 (N_28690,N_22681,N_20969);
and U28691 (N_28691,N_24034,N_23851);
nand U28692 (N_28692,N_23954,N_21852);
nor U28693 (N_28693,N_20926,N_22710);
or U28694 (N_28694,N_20914,N_20747);
and U28695 (N_28695,N_23255,N_20344);
nor U28696 (N_28696,N_20026,N_21159);
nand U28697 (N_28697,N_22472,N_20563);
and U28698 (N_28698,N_24564,N_20991);
nand U28699 (N_28699,N_24500,N_23786);
and U28700 (N_28700,N_20135,N_21118);
nand U28701 (N_28701,N_20992,N_24590);
or U28702 (N_28702,N_23232,N_24337);
or U28703 (N_28703,N_23177,N_20628);
or U28704 (N_28704,N_21204,N_22960);
and U28705 (N_28705,N_21716,N_20015);
nor U28706 (N_28706,N_20231,N_23150);
nand U28707 (N_28707,N_22507,N_23053);
or U28708 (N_28708,N_24714,N_20938);
and U28709 (N_28709,N_21888,N_23660);
or U28710 (N_28710,N_20919,N_24980);
or U28711 (N_28711,N_23896,N_20578);
nor U28712 (N_28712,N_21504,N_22416);
nor U28713 (N_28713,N_22373,N_24044);
nand U28714 (N_28714,N_22736,N_22329);
nor U28715 (N_28715,N_23573,N_23045);
xor U28716 (N_28716,N_23359,N_21152);
nor U28717 (N_28717,N_20241,N_22573);
nor U28718 (N_28718,N_21290,N_24993);
and U28719 (N_28719,N_21757,N_24065);
nand U28720 (N_28720,N_20028,N_23573);
and U28721 (N_28721,N_24750,N_22812);
or U28722 (N_28722,N_24031,N_24455);
or U28723 (N_28723,N_22469,N_20226);
nand U28724 (N_28724,N_22294,N_22251);
nand U28725 (N_28725,N_24466,N_23220);
or U28726 (N_28726,N_21638,N_24748);
nand U28727 (N_28727,N_21564,N_21680);
nand U28728 (N_28728,N_24625,N_20587);
nand U28729 (N_28729,N_21917,N_23363);
and U28730 (N_28730,N_20648,N_24576);
nor U28731 (N_28731,N_20868,N_24606);
or U28732 (N_28732,N_20345,N_20444);
or U28733 (N_28733,N_23185,N_20935);
and U28734 (N_28734,N_22913,N_22212);
nor U28735 (N_28735,N_21120,N_24056);
nand U28736 (N_28736,N_23685,N_20207);
and U28737 (N_28737,N_20467,N_20519);
nor U28738 (N_28738,N_21448,N_21459);
nand U28739 (N_28739,N_21630,N_24148);
nor U28740 (N_28740,N_22975,N_22809);
or U28741 (N_28741,N_23582,N_23886);
xor U28742 (N_28742,N_22931,N_23328);
or U28743 (N_28743,N_20237,N_21388);
nor U28744 (N_28744,N_20058,N_22836);
nand U28745 (N_28745,N_20473,N_21874);
nor U28746 (N_28746,N_24735,N_20900);
or U28747 (N_28747,N_24940,N_22218);
and U28748 (N_28748,N_20224,N_23713);
or U28749 (N_28749,N_21390,N_22314);
nand U28750 (N_28750,N_22073,N_24444);
nor U28751 (N_28751,N_23351,N_23173);
nand U28752 (N_28752,N_23682,N_22214);
and U28753 (N_28753,N_20003,N_23464);
or U28754 (N_28754,N_23299,N_20773);
nand U28755 (N_28755,N_24124,N_20007);
nor U28756 (N_28756,N_24210,N_21825);
nand U28757 (N_28757,N_22963,N_23573);
or U28758 (N_28758,N_21434,N_20844);
nor U28759 (N_28759,N_24815,N_22765);
nor U28760 (N_28760,N_23091,N_23420);
and U28761 (N_28761,N_23642,N_20313);
or U28762 (N_28762,N_23001,N_20720);
and U28763 (N_28763,N_23179,N_24341);
nand U28764 (N_28764,N_21899,N_23894);
or U28765 (N_28765,N_22130,N_20802);
and U28766 (N_28766,N_24491,N_24259);
or U28767 (N_28767,N_24222,N_21855);
nand U28768 (N_28768,N_23612,N_20924);
nand U28769 (N_28769,N_24490,N_22238);
xnor U28770 (N_28770,N_23096,N_20521);
nor U28771 (N_28771,N_23405,N_24411);
nor U28772 (N_28772,N_20784,N_21973);
xnor U28773 (N_28773,N_22439,N_24803);
or U28774 (N_28774,N_23076,N_24869);
or U28775 (N_28775,N_24408,N_20701);
nor U28776 (N_28776,N_23141,N_20638);
nand U28777 (N_28777,N_23094,N_20647);
nor U28778 (N_28778,N_23375,N_21936);
nand U28779 (N_28779,N_20392,N_21915);
nor U28780 (N_28780,N_23508,N_20932);
nand U28781 (N_28781,N_24231,N_21707);
and U28782 (N_28782,N_21920,N_23528);
or U28783 (N_28783,N_20081,N_21807);
and U28784 (N_28784,N_20404,N_20513);
or U28785 (N_28785,N_23660,N_20369);
or U28786 (N_28786,N_23530,N_22844);
nand U28787 (N_28787,N_23508,N_24924);
and U28788 (N_28788,N_20206,N_21550);
or U28789 (N_28789,N_24921,N_23822);
xor U28790 (N_28790,N_24288,N_21886);
xor U28791 (N_28791,N_24168,N_22000);
nor U28792 (N_28792,N_21081,N_23874);
or U28793 (N_28793,N_24398,N_21700);
and U28794 (N_28794,N_22293,N_22196);
or U28795 (N_28795,N_23368,N_22837);
nor U28796 (N_28796,N_20001,N_23813);
or U28797 (N_28797,N_24069,N_21959);
nand U28798 (N_28798,N_23721,N_23314);
nor U28799 (N_28799,N_22035,N_22550);
xor U28800 (N_28800,N_21684,N_24752);
nand U28801 (N_28801,N_24527,N_21592);
nor U28802 (N_28802,N_20729,N_22798);
or U28803 (N_28803,N_21093,N_21638);
nor U28804 (N_28804,N_20476,N_23466);
or U28805 (N_28805,N_22785,N_24254);
and U28806 (N_28806,N_24232,N_24507);
nand U28807 (N_28807,N_22320,N_23877);
nand U28808 (N_28808,N_20196,N_21052);
or U28809 (N_28809,N_24697,N_23858);
xor U28810 (N_28810,N_20946,N_20255);
and U28811 (N_28811,N_22618,N_24698);
and U28812 (N_28812,N_24289,N_23202);
nor U28813 (N_28813,N_21796,N_22971);
or U28814 (N_28814,N_24415,N_23826);
or U28815 (N_28815,N_22003,N_24905);
and U28816 (N_28816,N_22769,N_22033);
and U28817 (N_28817,N_24955,N_24099);
or U28818 (N_28818,N_21296,N_23318);
nand U28819 (N_28819,N_20055,N_22191);
nor U28820 (N_28820,N_20382,N_20902);
or U28821 (N_28821,N_24637,N_23958);
and U28822 (N_28822,N_22187,N_23381);
and U28823 (N_28823,N_23106,N_20227);
or U28824 (N_28824,N_24314,N_21189);
nor U28825 (N_28825,N_23015,N_23996);
xnor U28826 (N_28826,N_22489,N_21761);
nand U28827 (N_28827,N_20376,N_22590);
and U28828 (N_28828,N_20922,N_24323);
nor U28829 (N_28829,N_24225,N_23278);
or U28830 (N_28830,N_21256,N_22921);
or U28831 (N_28831,N_22352,N_24392);
and U28832 (N_28832,N_20188,N_21814);
xor U28833 (N_28833,N_23672,N_20711);
xnor U28834 (N_28834,N_23485,N_24015);
and U28835 (N_28835,N_23635,N_21146);
or U28836 (N_28836,N_20905,N_21196);
nor U28837 (N_28837,N_24307,N_23126);
nor U28838 (N_28838,N_20625,N_20145);
nor U28839 (N_28839,N_22895,N_21266);
xor U28840 (N_28840,N_20735,N_24904);
nor U28841 (N_28841,N_21083,N_22191);
or U28842 (N_28842,N_22041,N_24524);
and U28843 (N_28843,N_23306,N_21366);
nand U28844 (N_28844,N_24846,N_20135);
nand U28845 (N_28845,N_22660,N_22772);
or U28846 (N_28846,N_20036,N_20512);
or U28847 (N_28847,N_23995,N_23867);
and U28848 (N_28848,N_21725,N_22922);
nand U28849 (N_28849,N_23738,N_21537);
or U28850 (N_28850,N_23275,N_20214);
nor U28851 (N_28851,N_21443,N_24048);
and U28852 (N_28852,N_24557,N_22167);
and U28853 (N_28853,N_21097,N_22413);
or U28854 (N_28854,N_24842,N_23489);
or U28855 (N_28855,N_23250,N_21562);
or U28856 (N_28856,N_20089,N_22717);
and U28857 (N_28857,N_22371,N_23765);
nand U28858 (N_28858,N_22721,N_22110);
xor U28859 (N_28859,N_21544,N_22902);
and U28860 (N_28860,N_24698,N_21534);
and U28861 (N_28861,N_22463,N_20821);
nand U28862 (N_28862,N_20583,N_22816);
nand U28863 (N_28863,N_20727,N_21597);
nand U28864 (N_28864,N_20561,N_24649);
nand U28865 (N_28865,N_23036,N_22513);
and U28866 (N_28866,N_20304,N_21662);
and U28867 (N_28867,N_23388,N_24690);
xnor U28868 (N_28868,N_22972,N_21401);
or U28869 (N_28869,N_21855,N_23234);
and U28870 (N_28870,N_24770,N_20094);
nand U28871 (N_28871,N_21998,N_23096);
nor U28872 (N_28872,N_22911,N_22038);
nand U28873 (N_28873,N_24711,N_24466);
and U28874 (N_28874,N_21241,N_21448);
nand U28875 (N_28875,N_23477,N_20323);
and U28876 (N_28876,N_23070,N_21735);
nand U28877 (N_28877,N_24528,N_20500);
or U28878 (N_28878,N_24243,N_24764);
nand U28879 (N_28879,N_22590,N_21184);
nand U28880 (N_28880,N_20051,N_20217);
nand U28881 (N_28881,N_24190,N_24050);
or U28882 (N_28882,N_23537,N_24790);
and U28883 (N_28883,N_23428,N_22586);
nand U28884 (N_28884,N_22517,N_22716);
or U28885 (N_28885,N_22495,N_24287);
nand U28886 (N_28886,N_20178,N_22445);
nand U28887 (N_28887,N_21557,N_24162);
xor U28888 (N_28888,N_22758,N_22047);
or U28889 (N_28889,N_22631,N_20119);
nor U28890 (N_28890,N_23865,N_22856);
or U28891 (N_28891,N_20251,N_22891);
nor U28892 (N_28892,N_23549,N_23506);
or U28893 (N_28893,N_21119,N_23239);
nor U28894 (N_28894,N_23166,N_20657);
or U28895 (N_28895,N_22051,N_20614);
and U28896 (N_28896,N_23691,N_24223);
nand U28897 (N_28897,N_22824,N_24609);
nor U28898 (N_28898,N_22857,N_20790);
and U28899 (N_28899,N_22024,N_23957);
nor U28900 (N_28900,N_22414,N_22615);
xnor U28901 (N_28901,N_24948,N_21174);
or U28902 (N_28902,N_20925,N_22807);
nor U28903 (N_28903,N_22762,N_22278);
or U28904 (N_28904,N_24280,N_24115);
nand U28905 (N_28905,N_24786,N_20268);
and U28906 (N_28906,N_23887,N_21317);
nor U28907 (N_28907,N_21406,N_24494);
nor U28908 (N_28908,N_24991,N_23926);
nand U28909 (N_28909,N_20566,N_20654);
nor U28910 (N_28910,N_23928,N_24871);
nor U28911 (N_28911,N_22914,N_22954);
xor U28912 (N_28912,N_23231,N_23847);
nor U28913 (N_28913,N_23398,N_21417);
or U28914 (N_28914,N_23123,N_23236);
xnor U28915 (N_28915,N_23257,N_21614);
and U28916 (N_28916,N_24874,N_24162);
nand U28917 (N_28917,N_24986,N_20844);
nor U28918 (N_28918,N_24088,N_21367);
or U28919 (N_28919,N_21296,N_23091);
nor U28920 (N_28920,N_24767,N_24612);
and U28921 (N_28921,N_24982,N_21446);
nor U28922 (N_28922,N_23598,N_21867);
nand U28923 (N_28923,N_22083,N_24882);
or U28924 (N_28924,N_24275,N_21069);
nor U28925 (N_28925,N_22801,N_24709);
xnor U28926 (N_28926,N_21340,N_20168);
and U28927 (N_28927,N_23382,N_24110);
nand U28928 (N_28928,N_22375,N_21408);
and U28929 (N_28929,N_20950,N_23154);
and U28930 (N_28930,N_22742,N_24317);
or U28931 (N_28931,N_22792,N_20880);
or U28932 (N_28932,N_24628,N_20296);
or U28933 (N_28933,N_22362,N_24253);
or U28934 (N_28934,N_22886,N_22458);
nand U28935 (N_28935,N_22210,N_24986);
nor U28936 (N_28936,N_23870,N_20346);
and U28937 (N_28937,N_23507,N_21921);
nand U28938 (N_28938,N_20042,N_20751);
and U28939 (N_28939,N_23845,N_21266);
or U28940 (N_28940,N_23088,N_21879);
nor U28941 (N_28941,N_22124,N_22335);
nor U28942 (N_28942,N_22019,N_20206);
and U28943 (N_28943,N_21416,N_23156);
or U28944 (N_28944,N_20601,N_22894);
nor U28945 (N_28945,N_21513,N_21929);
or U28946 (N_28946,N_24476,N_24104);
or U28947 (N_28947,N_24915,N_22495);
and U28948 (N_28948,N_24875,N_21266);
and U28949 (N_28949,N_20884,N_23913);
nor U28950 (N_28950,N_24732,N_20200);
nor U28951 (N_28951,N_23368,N_20613);
and U28952 (N_28952,N_23438,N_21322);
and U28953 (N_28953,N_23262,N_20571);
nor U28954 (N_28954,N_24159,N_22865);
or U28955 (N_28955,N_24906,N_24683);
and U28956 (N_28956,N_24846,N_23441);
or U28957 (N_28957,N_22342,N_24024);
nand U28958 (N_28958,N_20940,N_20089);
nor U28959 (N_28959,N_20638,N_20143);
and U28960 (N_28960,N_20537,N_22075);
xnor U28961 (N_28961,N_21933,N_22563);
xnor U28962 (N_28962,N_21053,N_20885);
nor U28963 (N_28963,N_20315,N_23928);
or U28964 (N_28964,N_24711,N_23803);
nand U28965 (N_28965,N_24686,N_23385);
and U28966 (N_28966,N_23195,N_22971);
or U28967 (N_28967,N_21767,N_24623);
and U28968 (N_28968,N_21876,N_20289);
nand U28969 (N_28969,N_24369,N_20095);
nor U28970 (N_28970,N_22027,N_23872);
or U28971 (N_28971,N_24003,N_23914);
nand U28972 (N_28972,N_20334,N_22478);
or U28973 (N_28973,N_21728,N_22410);
or U28974 (N_28974,N_23291,N_22689);
nor U28975 (N_28975,N_22513,N_22618);
xor U28976 (N_28976,N_24981,N_20188);
or U28977 (N_28977,N_23835,N_22311);
nor U28978 (N_28978,N_22581,N_23248);
nor U28979 (N_28979,N_23101,N_24496);
nand U28980 (N_28980,N_22717,N_21257);
nand U28981 (N_28981,N_23341,N_20951);
or U28982 (N_28982,N_21046,N_21452);
xor U28983 (N_28983,N_24621,N_20374);
and U28984 (N_28984,N_24434,N_23399);
nand U28985 (N_28985,N_20862,N_22410);
xor U28986 (N_28986,N_24376,N_21445);
and U28987 (N_28987,N_22116,N_22668);
nor U28988 (N_28988,N_23948,N_23454);
nand U28989 (N_28989,N_21390,N_24297);
and U28990 (N_28990,N_22880,N_24559);
nand U28991 (N_28991,N_22350,N_21273);
and U28992 (N_28992,N_24364,N_20170);
nand U28993 (N_28993,N_22053,N_22095);
and U28994 (N_28994,N_21328,N_22142);
and U28995 (N_28995,N_24827,N_22108);
nor U28996 (N_28996,N_22027,N_20540);
nand U28997 (N_28997,N_23549,N_23762);
nor U28998 (N_28998,N_22266,N_24320);
xnor U28999 (N_28999,N_24626,N_24237);
and U29000 (N_29000,N_24201,N_22954);
and U29001 (N_29001,N_20340,N_24789);
xnor U29002 (N_29002,N_21386,N_20505);
or U29003 (N_29003,N_24021,N_20860);
nand U29004 (N_29004,N_24976,N_22397);
and U29005 (N_29005,N_20299,N_20282);
nand U29006 (N_29006,N_20928,N_24708);
nand U29007 (N_29007,N_23917,N_23435);
nor U29008 (N_29008,N_22439,N_22244);
and U29009 (N_29009,N_22091,N_22802);
or U29010 (N_29010,N_24979,N_22999);
and U29011 (N_29011,N_22575,N_22120);
and U29012 (N_29012,N_22338,N_20179);
and U29013 (N_29013,N_20205,N_22833);
and U29014 (N_29014,N_24369,N_24563);
nand U29015 (N_29015,N_20300,N_21901);
nor U29016 (N_29016,N_21490,N_23321);
nor U29017 (N_29017,N_20846,N_23340);
nor U29018 (N_29018,N_23656,N_21088);
nand U29019 (N_29019,N_21227,N_21945);
or U29020 (N_29020,N_21975,N_24874);
nor U29021 (N_29021,N_20837,N_24524);
nor U29022 (N_29022,N_23525,N_24191);
nand U29023 (N_29023,N_20742,N_24849);
nand U29024 (N_29024,N_22431,N_24729);
nand U29025 (N_29025,N_20747,N_23091);
and U29026 (N_29026,N_24521,N_24858);
and U29027 (N_29027,N_22197,N_22540);
or U29028 (N_29028,N_24535,N_20284);
xnor U29029 (N_29029,N_22812,N_22596);
or U29030 (N_29030,N_24774,N_21488);
or U29031 (N_29031,N_24520,N_23127);
and U29032 (N_29032,N_21233,N_24364);
and U29033 (N_29033,N_21644,N_22208);
and U29034 (N_29034,N_20169,N_22004);
and U29035 (N_29035,N_24387,N_22927);
nor U29036 (N_29036,N_22728,N_22079);
nor U29037 (N_29037,N_21020,N_24408);
nand U29038 (N_29038,N_24263,N_22856);
nor U29039 (N_29039,N_24474,N_24904);
nand U29040 (N_29040,N_23993,N_22102);
nand U29041 (N_29041,N_23117,N_22720);
nand U29042 (N_29042,N_20337,N_22252);
or U29043 (N_29043,N_24750,N_24292);
and U29044 (N_29044,N_20646,N_22506);
and U29045 (N_29045,N_24977,N_24805);
nor U29046 (N_29046,N_24900,N_23902);
nor U29047 (N_29047,N_22328,N_24159);
nor U29048 (N_29048,N_24267,N_21977);
and U29049 (N_29049,N_23134,N_20565);
or U29050 (N_29050,N_22588,N_23275);
or U29051 (N_29051,N_24458,N_22336);
and U29052 (N_29052,N_24624,N_21639);
and U29053 (N_29053,N_20394,N_24899);
or U29054 (N_29054,N_24785,N_20513);
or U29055 (N_29055,N_23049,N_24399);
nor U29056 (N_29056,N_21202,N_24849);
xnor U29057 (N_29057,N_21824,N_23814);
nor U29058 (N_29058,N_23638,N_21000);
nand U29059 (N_29059,N_24031,N_21392);
xnor U29060 (N_29060,N_24864,N_22498);
nor U29061 (N_29061,N_24860,N_20914);
nand U29062 (N_29062,N_20709,N_23329);
nand U29063 (N_29063,N_23566,N_21972);
and U29064 (N_29064,N_22019,N_24347);
nor U29065 (N_29065,N_22510,N_23213);
or U29066 (N_29066,N_24073,N_23152);
nand U29067 (N_29067,N_21766,N_24210);
nor U29068 (N_29068,N_22034,N_21769);
or U29069 (N_29069,N_20117,N_21193);
or U29070 (N_29070,N_21401,N_20810);
or U29071 (N_29071,N_23223,N_21904);
and U29072 (N_29072,N_21057,N_21319);
xor U29073 (N_29073,N_23633,N_24462);
nor U29074 (N_29074,N_24485,N_23253);
and U29075 (N_29075,N_23694,N_23927);
nand U29076 (N_29076,N_22694,N_21558);
and U29077 (N_29077,N_22739,N_23095);
xor U29078 (N_29078,N_23291,N_24063);
xor U29079 (N_29079,N_20779,N_23359);
nand U29080 (N_29080,N_22702,N_24174);
or U29081 (N_29081,N_20906,N_21319);
and U29082 (N_29082,N_20032,N_21765);
nand U29083 (N_29083,N_24405,N_23375);
or U29084 (N_29084,N_21618,N_24935);
nand U29085 (N_29085,N_24281,N_22084);
nand U29086 (N_29086,N_22970,N_23269);
or U29087 (N_29087,N_20909,N_20691);
nor U29088 (N_29088,N_22446,N_24625);
nand U29089 (N_29089,N_24358,N_20986);
nand U29090 (N_29090,N_21120,N_24096);
and U29091 (N_29091,N_22419,N_22079);
xor U29092 (N_29092,N_24990,N_20004);
nor U29093 (N_29093,N_23674,N_22192);
nor U29094 (N_29094,N_20978,N_21483);
xnor U29095 (N_29095,N_20798,N_23164);
nand U29096 (N_29096,N_21092,N_22541);
and U29097 (N_29097,N_22203,N_20893);
and U29098 (N_29098,N_21160,N_24134);
or U29099 (N_29099,N_23540,N_21025);
nor U29100 (N_29100,N_22834,N_20673);
or U29101 (N_29101,N_21900,N_21868);
nor U29102 (N_29102,N_20327,N_24416);
xor U29103 (N_29103,N_22916,N_20413);
xnor U29104 (N_29104,N_22111,N_23371);
nor U29105 (N_29105,N_20460,N_24351);
nand U29106 (N_29106,N_20816,N_23589);
and U29107 (N_29107,N_23168,N_24941);
or U29108 (N_29108,N_23761,N_21425);
or U29109 (N_29109,N_24282,N_24423);
and U29110 (N_29110,N_24652,N_22009);
xor U29111 (N_29111,N_21515,N_24644);
and U29112 (N_29112,N_22465,N_21241);
nor U29113 (N_29113,N_21820,N_21232);
nor U29114 (N_29114,N_22007,N_24188);
nor U29115 (N_29115,N_23616,N_23982);
or U29116 (N_29116,N_21018,N_20598);
nand U29117 (N_29117,N_22130,N_22260);
nor U29118 (N_29118,N_23941,N_24818);
or U29119 (N_29119,N_24451,N_22319);
xor U29120 (N_29120,N_21375,N_20106);
nor U29121 (N_29121,N_21142,N_20376);
nand U29122 (N_29122,N_24448,N_22310);
nand U29123 (N_29123,N_22509,N_23035);
and U29124 (N_29124,N_22769,N_22361);
nand U29125 (N_29125,N_23452,N_21641);
nor U29126 (N_29126,N_21644,N_20797);
xnor U29127 (N_29127,N_23375,N_20635);
or U29128 (N_29128,N_20962,N_20778);
and U29129 (N_29129,N_23665,N_23894);
nor U29130 (N_29130,N_24712,N_24136);
or U29131 (N_29131,N_24170,N_23303);
xnor U29132 (N_29132,N_22108,N_23980);
nor U29133 (N_29133,N_23778,N_23418);
or U29134 (N_29134,N_20212,N_24897);
nand U29135 (N_29135,N_24815,N_23279);
nand U29136 (N_29136,N_23521,N_20022);
or U29137 (N_29137,N_24612,N_24927);
and U29138 (N_29138,N_24712,N_24067);
xor U29139 (N_29139,N_22370,N_24108);
nand U29140 (N_29140,N_22965,N_24822);
or U29141 (N_29141,N_24689,N_21049);
or U29142 (N_29142,N_21697,N_23759);
and U29143 (N_29143,N_22356,N_24970);
and U29144 (N_29144,N_23458,N_21085);
and U29145 (N_29145,N_22814,N_23637);
or U29146 (N_29146,N_24659,N_24827);
or U29147 (N_29147,N_23251,N_21703);
nand U29148 (N_29148,N_24222,N_21510);
and U29149 (N_29149,N_24832,N_23347);
nand U29150 (N_29150,N_20630,N_24442);
nand U29151 (N_29151,N_21015,N_21069);
xnor U29152 (N_29152,N_22617,N_23289);
xor U29153 (N_29153,N_23367,N_22203);
and U29154 (N_29154,N_23351,N_21073);
nor U29155 (N_29155,N_22990,N_20908);
and U29156 (N_29156,N_24346,N_24300);
nor U29157 (N_29157,N_22926,N_22380);
nand U29158 (N_29158,N_22581,N_22081);
xnor U29159 (N_29159,N_24156,N_24936);
and U29160 (N_29160,N_24990,N_22503);
xnor U29161 (N_29161,N_24329,N_20394);
and U29162 (N_29162,N_24889,N_21216);
or U29163 (N_29163,N_21134,N_23793);
nor U29164 (N_29164,N_20374,N_20019);
nor U29165 (N_29165,N_24053,N_22840);
nand U29166 (N_29166,N_22217,N_22032);
nand U29167 (N_29167,N_24446,N_22220);
or U29168 (N_29168,N_23150,N_20371);
or U29169 (N_29169,N_24094,N_23229);
nor U29170 (N_29170,N_20553,N_23232);
and U29171 (N_29171,N_20064,N_23351);
nand U29172 (N_29172,N_22225,N_24938);
xor U29173 (N_29173,N_24336,N_21832);
or U29174 (N_29174,N_24804,N_23585);
nor U29175 (N_29175,N_22197,N_20553);
and U29176 (N_29176,N_23474,N_23256);
xnor U29177 (N_29177,N_22737,N_24601);
or U29178 (N_29178,N_23966,N_23170);
xor U29179 (N_29179,N_23928,N_20933);
nand U29180 (N_29180,N_20083,N_23488);
nand U29181 (N_29181,N_21021,N_23855);
nand U29182 (N_29182,N_23670,N_23906);
xor U29183 (N_29183,N_22108,N_23881);
and U29184 (N_29184,N_21670,N_21227);
and U29185 (N_29185,N_22001,N_20148);
or U29186 (N_29186,N_23267,N_24444);
xnor U29187 (N_29187,N_23301,N_21035);
and U29188 (N_29188,N_24774,N_20252);
nor U29189 (N_29189,N_21640,N_22567);
nor U29190 (N_29190,N_22634,N_24442);
xor U29191 (N_29191,N_22474,N_23111);
nor U29192 (N_29192,N_20018,N_23506);
and U29193 (N_29193,N_23406,N_20990);
nor U29194 (N_29194,N_24025,N_21077);
nand U29195 (N_29195,N_22535,N_20599);
or U29196 (N_29196,N_23042,N_23438);
nand U29197 (N_29197,N_21921,N_23134);
nor U29198 (N_29198,N_24416,N_23770);
nor U29199 (N_29199,N_22177,N_20779);
nor U29200 (N_29200,N_20281,N_22796);
xor U29201 (N_29201,N_24249,N_21969);
nand U29202 (N_29202,N_23912,N_24267);
xnor U29203 (N_29203,N_24797,N_21738);
nor U29204 (N_29204,N_20243,N_23091);
or U29205 (N_29205,N_21630,N_23694);
or U29206 (N_29206,N_20284,N_20157);
and U29207 (N_29207,N_23910,N_20300);
nand U29208 (N_29208,N_24850,N_23989);
or U29209 (N_29209,N_20152,N_23714);
or U29210 (N_29210,N_22132,N_20763);
nor U29211 (N_29211,N_24762,N_20092);
nor U29212 (N_29212,N_22842,N_21366);
or U29213 (N_29213,N_23719,N_22437);
and U29214 (N_29214,N_23909,N_24998);
nand U29215 (N_29215,N_21847,N_24027);
or U29216 (N_29216,N_21767,N_24009);
and U29217 (N_29217,N_21696,N_24768);
xnor U29218 (N_29218,N_23113,N_22867);
nor U29219 (N_29219,N_23993,N_24852);
nor U29220 (N_29220,N_23945,N_20760);
or U29221 (N_29221,N_24008,N_20382);
nor U29222 (N_29222,N_22022,N_20869);
nor U29223 (N_29223,N_23924,N_22143);
nor U29224 (N_29224,N_22423,N_24531);
and U29225 (N_29225,N_22017,N_21356);
nor U29226 (N_29226,N_24190,N_24377);
nor U29227 (N_29227,N_24466,N_20523);
nand U29228 (N_29228,N_24766,N_22992);
nor U29229 (N_29229,N_20721,N_21842);
nor U29230 (N_29230,N_22661,N_21493);
and U29231 (N_29231,N_22835,N_24601);
nand U29232 (N_29232,N_21975,N_20161);
or U29233 (N_29233,N_22375,N_21273);
nand U29234 (N_29234,N_24136,N_24586);
xor U29235 (N_29235,N_22678,N_23343);
xor U29236 (N_29236,N_24122,N_22121);
nand U29237 (N_29237,N_24204,N_21128);
nor U29238 (N_29238,N_24411,N_23694);
nor U29239 (N_29239,N_21544,N_21949);
and U29240 (N_29240,N_24276,N_20869);
nand U29241 (N_29241,N_20296,N_20969);
nor U29242 (N_29242,N_22816,N_23837);
xnor U29243 (N_29243,N_20700,N_23876);
nand U29244 (N_29244,N_23523,N_21860);
nor U29245 (N_29245,N_21575,N_21260);
and U29246 (N_29246,N_23902,N_22403);
and U29247 (N_29247,N_20194,N_22282);
or U29248 (N_29248,N_20333,N_21221);
nand U29249 (N_29249,N_22821,N_24520);
nand U29250 (N_29250,N_24098,N_23766);
or U29251 (N_29251,N_22257,N_22721);
nand U29252 (N_29252,N_24222,N_24860);
nand U29253 (N_29253,N_20776,N_24347);
xor U29254 (N_29254,N_20485,N_21686);
and U29255 (N_29255,N_24343,N_21798);
nor U29256 (N_29256,N_21776,N_21768);
nor U29257 (N_29257,N_23646,N_24486);
nor U29258 (N_29258,N_24216,N_23797);
or U29259 (N_29259,N_20973,N_22473);
xor U29260 (N_29260,N_23302,N_23197);
or U29261 (N_29261,N_21262,N_22049);
and U29262 (N_29262,N_24632,N_22659);
and U29263 (N_29263,N_21169,N_24304);
nand U29264 (N_29264,N_22260,N_20434);
nand U29265 (N_29265,N_22989,N_21173);
nand U29266 (N_29266,N_22752,N_23710);
nand U29267 (N_29267,N_20452,N_22168);
or U29268 (N_29268,N_23309,N_23749);
or U29269 (N_29269,N_24100,N_20396);
nand U29270 (N_29270,N_23202,N_20057);
and U29271 (N_29271,N_20448,N_22068);
nor U29272 (N_29272,N_20507,N_24588);
nand U29273 (N_29273,N_24619,N_23077);
nand U29274 (N_29274,N_23082,N_22318);
nor U29275 (N_29275,N_20880,N_20930);
nor U29276 (N_29276,N_21627,N_20884);
and U29277 (N_29277,N_21570,N_24878);
xnor U29278 (N_29278,N_20217,N_21017);
or U29279 (N_29279,N_22449,N_23788);
xor U29280 (N_29280,N_23109,N_22009);
xnor U29281 (N_29281,N_20621,N_24914);
xnor U29282 (N_29282,N_20878,N_20354);
or U29283 (N_29283,N_24355,N_22756);
nand U29284 (N_29284,N_23014,N_24067);
and U29285 (N_29285,N_20363,N_20386);
or U29286 (N_29286,N_20076,N_21603);
or U29287 (N_29287,N_20951,N_22503);
xor U29288 (N_29288,N_20183,N_24972);
xnor U29289 (N_29289,N_20101,N_20603);
nand U29290 (N_29290,N_24414,N_20732);
and U29291 (N_29291,N_23551,N_24604);
and U29292 (N_29292,N_22640,N_23434);
or U29293 (N_29293,N_21965,N_20496);
or U29294 (N_29294,N_23916,N_21440);
or U29295 (N_29295,N_21207,N_22218);
or U29296 (N_29296,N_22955,N_21232);
or U29297 (N_29297,N_22186,N_20687);
or U29298 (N_29298,N_20066,N_20802);
nand U29299 (N_29299,N_23573,N_21561);
or U29300 (N_29300,N_20631,N_24902);
or U29301 (N_29301,N_22038,N_22643);
or U29302 (N_29302,N_21738,N_23129);
or U29303 (N_29303,N_22824,N_23770);
or U29304 (N_29304,N_23599,N_21864);
or U29305 (N_29305,N_20078,N_21664);
nor U29306 (N_29306,N_22211,N_22186);
and U29307 (N_29307,N_21400,N_23394);
or U29308 (N_29308,N_23821,N_20312);
nor U29309 (N_29309,N_20000,N_21532);
xor U29310 (N_29310,N_22678,N_24215);
or U29311 (N_29311,N_24653,N_22874);
xor U29312 (N_29312,N_20790,N_20068);
nand U29313 (N_29313,N_20910,N_20958);
xnor U29314 (N_29314,N_24599,N_20175);
and U29315 (N_29315,N_23344,N_21879);
nor U29316 (N_29316,N_24375,N_22069);
nand U29317 (N_29317,N_21618,N_21556);
or U29318 (N_29318,N_22404,N_22006);
nor U29319 (N_29319,N_23317,N_22050);
xnor U29320 (N_29320,N_24985,N_21231);
nand U29321 (N_29321,N_22649,N_23212);
or U29322 (N_29322,N_20545,N_20095);
nor U29323 (N_29323,N_24462,N_21485);
nor U29324 (N_29324,N_23074,N_22468);
nand U29325 (N_29325,N_24870,N_21387);
and U29326 (N_29326,N_24768,N_22820);
or U29327 (N_29327,N_23158,N_23219);
or U29328 (N_29328,N_23254,N_23623);
nand U29329 (N_29329,N_20308,N_23735);
nand U29330 (N_29330,N_22024,N_23698);
nand U29331 (N_29331,N_24452,N_24049);
nand U29332 (N_29332,N_20587,N_23561);
and U29333 (N_29333,N_22904,N_23679);
and U29334 (N_29334,N_22351,N_20462);
nand U29335 (N_29335,N_24907,N_24747);
nand U29336 (N_29336,N_22558,N_21287);
or U29337 (N_29337,N_22464,N_24370);
xnor U29338 (N_29338,N_24114,N_20431);
nand U29339 (N_29339,N_22611,N_23957);
nor U29340 (N_29340,N_23076,N_20967);
or U29341 (N_29341,N_21105,N_21494);
and U29342 (N_29342,N_22736,N_24312);
and U29343 (N_29343,N_24474,N_20794);
or U29344 (N_29344,N_23075,N_24074);
or U29345 (N_29345,N_21429,N_23465);
or U29346 (N_29346,N_20322,N_23430);
nor U29347 (N_29347,N_24356,N_20020);
nor U29348 (N_29348,N_23268,N_24005);
nor U29349 (N_29349,N_24333,N_23941);
and U29350 (N_29350,N_23212,N_24290);
or U29351 (N_29351,N_23927,N_24740);
xor U29352 (N_29352,N_20157,N_23305);
nor U29353 (N_29353,N_23615,N_24544);
nand U29354 (N_29354,N_22055,N_22179);
nor U29355 (N_29355,N_20354,N_20999);
or U29356 (N_29356,N_24051,N_24100);
or U29357 (N_29357,N_23639,N_22023);
nor U29358 (N_29358,N_24159,N_23576);
and U29359 (N_29359,N_22832,N_23693);
nor U29360 (N_29360,N_24536,N_24627);
or U29361 (N_29361,N_24888,N_22845);
nor U29362 (N_29362,N_20842,N_21575);
xnor U29363 (N_29363,N_22404,N_20190);
or U29364 (N_29364,N_23738,N_24236);
or U29365 (N_29365,N_22407,N_23324);
and U29366 (N_29366,N_22709,N_21442);
nor U29367 (N_29367,N_21574,N_24396);
nor U29368 (N_29368,N_24623,N_22402);
or U29369 (N_29369,N_24739,N_23942);
or U29370 (N_29370,N_22339,N_22331);
or U29371 (N_29371,N_22955,N_24978);
or U29372 (N_29372,N_21081,N_21027);
or U29373 (N_29373,N_21311,N_23008);
nor U29374 (N_29374,N_24930,N_22927);
nand U29375 (N_29375,N_22256,N_22560);
or U29376 (N_29376,N_22353,N_22009);
and U29377 (N_29377,N_20117,N_24902);
and U29378 (N_29378,N_24777,N_24032);
nor U29379 (N_29379,N_22409,N_21085);
nor U29380 (N_29380,N_24466,N_22455);
nor U29381 (N_29381,N_24911,N_21200);
or U29382 (N_29382,N_21368,N_22741);
or U29383 (N_29383,N_24394,N_23053);
xor U29384 (N_29384,N_23300,N_21635);
nand U29385 (N_29385,N_21089,N_21265);
nor U29386 (N_29386,N_24374,N_21822);
and U29387 (N_29387,N_21321,N_23323);
and U29388 (N_29388,N_21932,N_24562);
and U29389 (N_29389,N_21381,N_22868);
and U29390 (N_29390,N_22121,N_23766);
nor U29391 (N_29391,N_20037,N_22715);
nand U29392 (N_29392,N_21288,N_23767);
or U29393 (N_29393,N_24066,N_22337);
nand U29394 (N_29394,N_20309,N_22473);
and U29395 (N_29395,N_24821,N_22324);
nor U29396 (N_29396,N_24498,N_20806);
xnor U29397 (N_29397,N_21070,N_23288);
nand U29398 (N_29398,N_21153,N_20534);
and U29399 (N_29399,N_23261,N_22797);
nor U29400 (N_29400,N_20713,N_23270);
nand U29401 (N_29401,N_22266,N_21246);
and U29402 (N_29402,N_22964,N_23132);
and U29403 (N_29403,N_20020,N_21204);
nor U29404 (N_29404,N_22417,N_24982);
xor U29405 (N_29405,N_24595,N_21016);
xor U29406 (N_29406,N_23770,N_20235);
and U29407 (N_29407,N_21326,N_24155);
nor U29408 (N_29408,N_23251,N_23453);
or U29409 (N_29409,N_23715,N_21082);
nor U29410 (N_29410,N_21391,N_22049);
nand U29411 (N_29411,N_21539,N_24845);
or U29412 (N_29412,N_22958,N_22064);
nand U29413 (N_29413,N_22457,N_23394);
or U29414 (N_29414,N_23422,N_20955);
and U29415 (N_29415,N_20038,N_21779);
nor U29416 (N_29416,N_24693,N_21953);
or U29417 (N_29417,N_21112,N_20112);
nor U29418 (N_29418,N_21669,N_23326);
nand U29419 (N_29419,N_20769,N_21703);
nor U29420 (N_29420,N_23528,N_21880);
or U29421 (N_29421,N_23780,N_24576);
and U29422 (N_29422,N_22127,N_24862);
or U29423 (N_29423,N_21718,N_23636);
and U29424 (N_29424,N_24899,N_20827);
or U29425 (N_29425,N_24299,N_22231);
xor U29426 (N_29426,N_23626,N_22852);
or U29427 (N_29427,N_21408,N_23997);
or U29428 (N_29428,N_24807,N_23040);
nor U29429 (N_29429,N_22942,N_24061);
or U29430 (N_29430,N_22351,N_20328);
or U29431 (N_29431,N_22408,N_23437);
or U29432 (N_29432,N_21859,N_22269);
or U29433 (N_29433,N_20891,N_21446);
nand U29434 (N_29434,N_21074,N_21609);
or U29435 (N_29435,N_21610,N_20649);
and U29436 (N_29436,N_21141,N_22716);
nor U29437 (N_29437,N_22597,N_21925);
nor U29438 (N_29438,N_24924,N_22301);
or U29439 (N_29439,N_23561,N_21710);
nor U29440 (N_29440,N_21185,N_20342);
nor U29441 (N_29441,N_21740,N_21585);
nor U29442 (N_29442,N_24043,N_20719);
nand U29443 (N_29443,N_22925,N_21073);
and U29444 (N_29444,N_20852,N_24019);
nand U29445 (N_29445,N_22656,N_22670);
or U29446 (N_29446,N_22212,N_24540);
xnor U29447 (N_29447,N_24787,N_22574);
nor U29448 (N_29448,N_23708,N_20923);
nand U29449 (N_29449,N_23028,N_23534);
and U29450 (N_29450,N_24327,N_22506);
nand U29451 (N_29451,N_21231,N_23260);
or U29452 (N_29452,N_22086,N_20967);
or U29453 (N_29453,N_22372,N_20539);
nor U29454 (N_29454,N_23624,N_23572);
and U29455 (N_29455,N_24059,N_21903);
and U29456 (N_29456,N_21028,N_24940);
and U29457 (N_29457,N_24782,N_20970);
or U29458 (N_29458,N_23831,N_23292);
nor U29459 (N_29459,N_24920,N_23137);
nor U29460 (N_29460,N_23749,N_24940);
or U29461 (N_29461,N_24791,N_24269);
or U29462 (N_29462,N_23829,N_23422);
xnor U29463 (N_29463,N_22423,N_24460);
xor U29464 (N_29464,N_21799,N_24541);
nor U29465 (N_29465,N_22576,N_20378);
nand U29466 (N_29466,N_22871,N_23321);
nor U29467 (N_29467,N_23313,N_23834);
nor U29468 (N_29468,N_22987,N_24362);
nor U29469 (N_29469,N_23514,N_21487);
nand U29470 (N_29470,N_22119,N_23395);
nor U29471 (N_29471,N_20412,N_20339);
nor U29472 (N_29472,N_22531,N_21186);
nor U29473 (N_29473,N_24153,N_20541);
or U29474 (N_29474,N_22305,N_23332);
nor U29475 (N_29475,N_21659,N_22462);
and U29476 (N_29476,N_20165,N_22591);
nor U29477 (N_29477,N_20595,N_21702);
nor U29478 (N_29478,N_22236,N_21943);
and U29479 (N_29479,N_23643,N_20702);
nand U29480 (N_29480,N_21299,N_20688);
and U29481 (N_29481,N_23412,N_20318);
or U29482 (N_29482,N_23087,N_20792);
or U29483 (N_29483,N_23142,N_22097);
nor U29484 (N_29484,N_20745,N_21704);
and U29485 (N_29485,N_21713,N_24223);
nor U29486 (N_29486,N_20434,N_24169);
and U29487 (N_29487,N_21690,N_22547);
or U29488 (N_29488,N_21765,N_23925);
nor U29489 (N_29489,N_23436,N_20276);
and U29490 (N_29490,N_20816,N_21722);
xnor U29491 (N_29491,N_22472,N_22085);
nand U29492 (N_29492,N_22646,N_21107);
and U29493 (N_29493,N_22362,N_21773);
or U29494 (N_29494,N_23750,N_23911);
nor U29495 (N_29495,N_24207,N_20737);
and U29496 (N_29496,N_20084,N_22387);
and U29497 (N_29497,N_22677,N_21804);
xnor U29498 (N_29498,N_24518,N_24858);
and U29499 (N_29499,N_24781,N_22817);
nor U29500 (N_29500,N_23429,N_23939);
and U29501 (N_29501,N_21293,N_24029);
and U29502 (N_29502,N_22480,N_20088);
and U29503 (N_29503,N_20533,N_20786);
nor U29504 (N_29504,N_23116,N_20102);
nor U29505 (N_29505,N_21496,N_24215);
xnor U29506 (N_29506,N_24150,N_24221);
nor U29507 (N_29507,N_24233,N_22987);
xnor U29508 (N_29508,N_23009,N_24079);
or U29509 (N_29509,N_23967,N_22549);
xor U29510 (N_29510,N_24649,N_21890);
nor U29511 (N_29511,N_20453,N_21863);
nor U29512 (N_29512,N_22864,N_23759);
and U29513 (N_29513,N_20843,N_23437);
nor U29514 (N_29514,N_23131,N_20605);
and U29515 (N_29515,N_24328,N_22265);
and U29516 (N_29516,N_22049,N_20396);
and U29517 (N_29517,N_20346,N_23408);
nor U29518 (N_29518,N_23471,N_22215);
xnor U29519 (N_29519,N_23145,N_20400);
nor U29520 (N_29520,N_22655,N_23033);
nor U29521 (N_29521,N_20709,N_21510);
or U29522 (N_29522,N_23183,N_22759);
or U29523 (N_29523,N_22136,N_22816);
nor U29524 (N_29524,N_21128,N_22879);
and U29525 (N_29525,N_22659,N_24910);
nor U29526 (N_29526,N_24794,N_21801);
and U29527 (N_29527,N_20021,N_23159);
nand U29528 (N_29528,N_21500,N_21159);
nand U29529 (N_29529,N_22681,N_21673);
and U29530 (N_29530,N_23584,N_20686);
and U29531 (N_29531,N_21858,N_23941);
nor U29532 (N_29532,N_24057,N_22740);
nand U29533 (N_29533,N_23360,N_21865);
nor U29534 (N_29534,N_22550,N_22433);
nand U29535 (N_29535,N_23739,N_20026);
and U29536 (N_29536,N_20646,N_23774);
nor U29537 (N_29537,N_22592,N_22176);
or U29538 (N_29538,N_21551,N_20032);
nor U29539 (N_29539,N_24112,N_23738);
and U29540 (N_29540,N_20226,N_22113);
or U29541 (N_29541,N_23633,N_22096);
or U29542 (N_29542,N_21501,N_24150);
and U29543 (N_29543,N_24425,N_21967);
nand U29544 (N_29544,N_23564,N_22579);
xor U29545 (N_29545,N_24441,N_24002);
nor U29546 (N_29546,N_20625,N_23948);
nor U29547 (N_29547,N_20104,N_22947);
and U29548 (N_29548,N_24240,N_21824);
nor U29549 (N_29549,N_21820,N_23381);
xor U29550 (N_29550,N_20754,N_24865);
and U29551 (N_29551,N_21641,N_21143);
or U29552 (N_29552,N_23467,N_22351);
nor U29553 (N_29553,N_21544,N_23616);
nor U29554 (N_29554,N_21714,N_20420);
nand U29555 (N_29555,N_20451,N_20040);
nor U29556 (N_29556,N_24602,N_21314);
or U29557 (N_29557,N_21127,N_24511);
nand U29558 (N_29558,N_22377,N_20523);
and U29559 (N_29559,N_21987,N_22898);
nand U29560 (N_29560,N_24176,N_20683);
and U29561 (N_29561,N_22378,N_20339);
nor U29562 (N_29562,N_23999,N_20462);
nor U29563 (N_29563,N_20424,N_21574);
and U29564 (N_29564,N_21388,N_21173);
nor U29565 (N_29565,N_24153,N_23700);
and U29566 (N_29566,N_22667,N_20635);
nand U29567 (N_29567,N_20552,N_20657);
or U29568 (N_29568,N_24412,N_22606);
nor U29569 (N_29569,N_21326,N_23964);
nand U29570 (N_29570,N_24501,N_20206);
nand U29571 (N_29571,N_24126,N_23938);
and U29572 (N_29572,N_24270,N_24107);
and U29573 (N_29573,N_22194,N_20791);
nand U29574 (N_29574,N_23595,N_23260);
nor U29575 (N_29575,N_23681,N_22812);
and U29576 (N_29576,N_22179,N_23043);
nand U29577 (N_29577,N_24564,N_21313);
or U29578 (N_29578,N_23358,N_24517);
or U29579 (N_29579,N_24867,N_20036);
nand U29580 (N_29580,N_22194,N_22318);
nand U29581 (N_29581,N_24715,N_24210);
and U29582 (N_29582,N_23415,N_24090);
and U29583 (N_29583,N_21183,N_20366);
nand U29584 (N_29584,N_24818,N_22318);
and U29585 (N_29585,N_22729,N_24292);
and U29586 (N_29586,N_24716,N_21051);
and U29587 (N_29587,N_21099,N_21845);
or U29588 (N_29588,N_21925,N_24556);
nor U29589 (N_29589,N_21767,N_23249);
and U29590 (N_29590,N_20764,N_23573);
or U29591 (N_29591,N_24954,N_22355);
nor U29592 (N_29592,N_22046,N_20596);
and U29593 (N_29593,N_24999,N_21320);
nand U29594 (N_29594,N_22958,N_21168);
nand U29595 (N_29595,N_20494,N_22268);
or U29596 (N_29596,N_20233,N_22943);
nand U29597 (N_29597,N_24430,N_22862);
nor U29598 (N_29598,N_21654,N_23429);
nand U29599 (N_29599,N_23768,N_22183);
and U29600 (N_29600,N_21880,N_24244);
nand U29601 (N_29601,N_24060,N_24822);
xor U29602 (N_29602,N_23158,N_23929);
or U29603 (N_29603,N_24397,N_22556);
and U29604 (N_29604,N_21586,N_24179);
nor U29605 (N_29605,N_23835,N_21646);
nor U29606 (N_29606,N_23791,N_22797);
and U29607 (N_29607,N_23646,N_24281);
nor U29608 (N_29608,N_22505,N_22395);
or U29609 (N_29609,N_20383,N_20521);
and U29610 (N_29610,N_23768,N_22480);
or U29611 (N_29611,N_20629,N_23506);
or U29612 (N_29612,N_23328,N_20307);
nand U29613 (N_29613,N_24089,N_22806);
nor U29614 (N_29614,N_21728,N_23468);
xnor U29615 (N_29615,N_20608,N_24094);
nor U29616 (N_29616,N_22334,N_24691);
nand U29617 (N_29617,N_22656,N_20884);
and U29618 (N_29618,N_23297,N_21575);
and U29619 (N_29619,N_22876,N_23098);
nand U29620 (N_29620,N_21593,N_20919);
nand U29621 (N_29621,N_24121,N_24615);
nor U29622 (N_29622,N_20691,N_20265);
nor U29623 (N_29623,N_20617,N_23920);
nand U29624 (N_29624,N_20934,N_22985);
or U29625 (N_29625,N_23221,N_24873);
xor U29626 (N_29626,N_23901,N_23857);
nor U29627 (N_29627,N_21204,N_23688);
nor U29628 (N_29628,N_21812,N_23973);
and U29629 (N_29629,N_24667,N_23418);
or U29630 (N_29630,N_20791,N_20653);
or U29631 (N_29631,N_22181,N_22407);
nor U29632 (N_29632,N_22546,N_24540);
xnor U29633 (N_29633,N_22484,N_22497);
nand U29634 (N_29634,N_22337,N_22876);
and U29635 (N_29635,N_22525,N_20981);
or U29636 (N_29636,N_20777,N_22310);
nand U29637 (N_29637,N_24072,N_24604);
and U29638 (N_29638,N_20941,N_21683);
nor U29639 (N_29639,N_22152,N_20428);
xor U29640 (N_29640,N_20843,N_23959);
or U29641 (N_29641,N_22969,N_21125);
or U29642 (N_29642,N_21358,N_22329);
nor U29643 (N_29643,N_24690,N_23674);
nand U29644 (N_29644,N_22441,N_24053);
nand U29645 (N_29645,N_23536,N_20305);
nor U29646 (N_29646,N_20572,N_22227);
or U29647 (N_29647,N_24488,N_23923);
xor U29648 (N_29648,N_21737,N_23764);
or U29649 (N_29649,N_20393,N_20007);
or U29650 (N_29650,N_23806,N_23131);
nand U29651 (N_29651,N_24400,N_20863);
or U29652 (N_29652,N_23583,N_21341);
and U29653 (N_29653,N_22206,N_22268);
and U29654 (N_29654,N_23901,N_23802);
or U29655 (N_29655,N_23319,N_22065);
nand U29656 (N_29656,N_24199,N_20646);
and U29657 (N_29657,N_24218,N_22429);
nand U29658 (N_29658,N_20733,N_23295);
nand U29659 (N_29659,N_21806,N_20832);
and U29660 (N_29660,N_23013,N_22599);
or U29661 (N_29661,N_21394,N_21020);
and U29662 (N_29662,N_24248,N_20730);
nor U29663 (N_29663,N_21503,N_23923);
and U29664 (N_29664,N_23283,N_24901);
and U29665 (N_29665,N_20323,N_23645);
nand U29666 (N_29666,N_21844,N_21197);
nand U29667 (N_29667,N_24407,N_23744);
nand U29668 (N_29668,N_21917,N_24396);
xnor U29669 (N_29669,N_21634,N_21211);
and U29670 (N_29670,N_23409,N_22008);
xnor U29671 (N_29671,N_23186,N_20653);
nand U29672 (N_29672,N_22123,N_20034);
and U29673 (N_29673,N_20272,N_24613);
and U29674 (N_29674,N_24101,N_22021);
and U29675 (N_29675,N_23572,N_20076);
and U29676 (N_29676,N_20216,N_21551);
or U29677 (N_29677,N_22351,N_22449);
xnor U29678 (N_29678,N_20917,N_24008);
or U29679 (N_29679,N_23120,N_21403);
or U29680 (N_29680,N_20505,N_23407);
xnor U29681 (N_29681,N_22554,N_23318);
nor U29682 (N_29682,N_24089,N_21372);
xor U29683 (N_29683,N_24784,N_24301);
and U29684 (N_29684,N_21274,N_21994);
and U29685 (N_29685,N_20171,N_23274);
or U29686 (N_29686,N_22217,N_24111);
nor U29687 (N_29687,N_22776,N_23350);
nand U29688 (N_29688,N_24592,N_21627);
nand U29689 (N_29689,N_24789,N_21083);
or U29690 (N_29690,N_24948,N_21618);
nand U29691 (N_29691,N_22323,N_23883);
nor U29692 (N_29692,N_21607,N_20336);
nor U29693 (N_29693,N_23398,N_22800);
nand U29694 (N_29694,N_23265,N_22434);
xnor U29695 (N_29695,N_22601,N_21640);
nand U29696 (N_29696,N_21681,N_24892);
nand U29697 (N_29697,N_24808,N_23222);
nor U29698 (N_29698,N_23028,N_22145);
nand U29699 (N_29699,N_20657,N_24235);
xnor U29700 (N_29700,N_20046,N_21305);
and U29701 (N_29701,N_24645,N_22529);
xor U29702 (N_29702,N_22335,N_21518);
and U29703 (N_29703,N_21208,N_24018);
nand U29704 (N_29704,N_24940,N_23947);
or U29705 (N_29705,N_22938,N_22492);
and U29706 (N_29706,N_23493,N_22833);
nand U29707 (N_29707,N_20367,N_23772);
nand U29708 (N_29708,N_21303,N_22833);
nor U29709 (N_29709,N_23711,N_21252);
or U29710 (N_29710,N_24854,N_21727);
nor U29711 (N_29711,N_23056,N_23736);
nor U29712 (N_29712,N_24243,N_23069);
nand U29713 (N_29713,N_21333,N_23801);
or U29714 (N_29714,N_24577,N_20128);
and U29715 (N_29715,N_21978,N_22634);
or U29716 (N_29716,N_21900,N_20053);
nand U29717 (N_29717,N_22358,N_23120);
nor U29718 (N_29718,N_20884,N_21007);
nor U29719 (N_29719,N_23936,N_20417);
and U29720 (N_29720,N_20126,N_24418);
xnor U29721 (N_29721,N_22611,N_20691);
xor U29722 (N_29722,N_24388,N_21170);
and U29723 (N_29723,N_24688,N_21211);
nand U29724 (N_29724,N_24510,N_22049);
xor U29725 (N_29725,N_22171,N_24125);
nor U29726 (N_29726,N_23736,N_21002);
nor U29727 (N_29727,N_20980,N_20710);
nor U29728 (N_29728,N_24487,N_20207);
xnor U29729 (N_29729,N_24392,N_22815);
or U29730 (N_29730,N_22506,N_21444);
nor U29731 (N_29731,N_23507,N_23296);
nor U29732 (N_29732,N_21017,N_23661);
nand U29733 (N_29733,N_20776,N_21451);
or U29734 (N_29734,N_22840,N_22588);
nor U29735 (N_29735,N_20672,N_23623);
and U29736 (N_29736,N_22451,N_24500);
nand U29737 (N_29737,N_22483,N_20941);
nand U29738 (N_29738,N_23543,N_22813);
nor U29739 (N_29739,N_22237,N_22288);
or U29740 (N_29740,N_21082,N_24505);
nor U29741 (N_29741,N_24156,N_24586);
and U29742 (N_29742,N_20817,N_22874);
nor U29743 (N_29743,N_24118,N_21816);
and U29744 (N_29744,N_23137,N_22656);
or U29745 (N_29745,N_20268,N_23950);
nand U29746 (N_29746,N_23641,N_21486);
and U29747 (N_29747,N_21880,N_21877);
nand U29748 (N_29748,N_20472,N_21695);
or U29749 (N_29749,N_23616,N_23253);
nand U29750 (N_29750,N_22555,N_22824);
nor U29751 (N_29751,N_24222,N_22794);
or U29752 (N_29752,N_21759,N_20400);
nor U29753 (N_29753,N_23497,N_20981);
nand U29754 (N_29754,N_21597,N_23259);
and U29755 (N_29755,N_20943,N_22173);
and U29756 (N_29756,N_23574,N_23575);
nor U29757 (N_29757,N_22037,N_21164);
and U29758 (N_29758,N_24867,N_22906);
or U29759 (N_29759,N_24661,N_21551);
or U29760 (N_29760,N_23253,N_23690);
nor U29761 (N_29761,N_22086,N_22281);
and U29762 (N_29762,N_23546,N_20712);
or U29763 (N_29763,N_23683,N_22504);
or U29764 (N_29764,N_20748,N_21179);
nor U29765 (N_29765,N_23581,N_20856);
nand U29766 (N_29766,N_24275,N_24844);
nor U29767 (N_29767,N_24473,N_23504);
or U29768 (N_29768,N_21566,N_24519);
or U29769 (N_29769,N_21704,N_24197);
and U29770 (N_29770,N_23305,N_20730);
xor U29771 (N_29771,N_22519,N_24483);
nand U29772 (N_29772,N_23566,N_21850);
xnor U29773 (N_29773,N_20501,N_23878);
nand U29774 (N_29774,N_23927,N_23061);
nor U29775 (N_29775,N_20205,N_22616);
and U29776 (N_29776,N_23005,N_21727);
or U29777 (N_29777,N_22213,N_22214);
and U29778 (N_29778,N_24018,N_24679);
or U29779 (N_29779,N_21821,N_21350);
nand U29780 (N_29780,N_23164,N_21207);
nand U29781 (N_29781,N_20151,N_23359);
nand U29782 (N_29782,N_24714,N_23896);
nand U29783 (N_29783,N_24472,N_21443);
and U29784 (N_29784,N_24143,N_20472);
nor U29785 (N_29785,N_22267,N_22552);
and U29786 (N_29786,N_21007,N_20722);
or U29787 (N_29787,N_20331,N_23872);
or U29788 (N_29788,N_24185,N_23622);
nand U29789 (N_29789,N_20638,N_24706);
and U29790 (N_29790,N_22873,N_21166);
or U29791 (N_29791,N_23648,N_22224);
and U29792 (N_29792,N_20547,N_20080);
and U29793 (N_29793,N_24063,N_22779);
nand U29794 (N_29794,N_20174,N_21789);
nand U29795 (N_29795,N_22959,N_23339);
or U29796 (N_29796,N_24688,N_22805);
or U29797 (N_29797,N_23659,N_21474);
or U29798 (N_29798,N_24768,N_23721);
nand U29799 (N_29799,N_23407,N_22987);
or U29800 (N_29800,N_20931,N_21646);
or U29801 (N_29801,N_22331,N_20517);
nor U29802 (N_29802,N_20337,N_21434);
xnor U29803 (N_29803,N_21503,N_21992);
nor U29804 (N_29804,N_22918,N_23997);
nand U29805 (N_29805,N_22514,N_24262);
nor U29806 (N_29806,N_20867,N_22885);
nand U29807 (N_29807,N_24914,N_21407);
xnor U29808 (N_29808,N_20870,N_22764);
nor U29809 (N_29809,N_24413,N_21382);
nand U29810 (N_29810,N_20085,N_21336);
nand U29811 (N_29811,N_24538,N_21217);
nor U29812 (N_29812,N_23937,N_22391);
and U29813 (N_29813,N_24276,N_24045);
nand U29814 (N_29814,N_20206,N_23009);
nand U29815 (N_29815,N_21314,N_20516);
and U29816 (N_29816,N_23873,N_23472);
and U29817 (N_29817,N_22236,N_23443);
and U29818 (N_29818,N_21409,N_24346);
and U29819 (N_29819,N_21185,N_20705);
and U29820 (N_29820,N_23477,N_21345);
nor U29821 (N_29821,N_22276,N_23147);
nor U29822 (N_29822,N_21444,N_22923);
nor U29823 (N_29823,N_24893,N_24604);
xor U29824 (N_29824,N_23234,N_24538);
and U29825 (N_29825,N_21632,N_24352);
nand U29826 (N_29826,N_20987,N_24582);
xor U29827 (N_29827,N_24203,N_22056);
nand U29828 (N_29828,N_23023,N_24939);
xor U29829 (N_29829,N_23640,N_23967);
nor U29830 (N_29830,N_24716,N_20764);
nand U29831 (N_29831,N_24060,N_22208);
nor U29832 (N_29832,N_24248,N_21384);
nand U29833 (N_29833,N_23121,N_23215);
nor U29834 (N_29834,N_21851,N_23944);
or U29835 (N_29835,N_21923,N_23361);
nor U29836 (N_29836,N_22148,N_23727);
nor U29837 (N_29837,N_22586,N_22218);
or U29838 (N_29838,N_22377,N_24439);
or U29839 (N_29839,N_20327,N_24299);
xnor U29840 (N_29840,N_20204,N_20721);
nor U29841 (N_29841,N_20467,N_24166);
nor U29842 (N_29842,N_20534,N_21636);
and U29843 (N_29843,N_22920,N_24103);
or U29844 (N_29844,N_20355,N_21255);
and U29845 (N_29845,N_21063,N_22720);
nand U29846 (N_29846,N_22848,N_21718);
nand U29847 (N_29847,N_23027,N_22704);
nor U29848 (N_29848,N_24342,N_22142);
nand U29849 (N_29849,N_20611,N_24205);
or U29850 (N_29850,N_20261,N_23546);
or U29851 (N_29851,N_20890,N_20528);
xor U29852 (N_29852,N_23738,N_21224);
xnor U29853 (N_29853,N_22124,N_20935);
or U29854 (N_29854,N_21726,N_20099);
nand U29855 (N_29855,N_23879,N_20503);
or U29856 (N_29856,N_21356,N_22958);
and U29857 (N_29857,N_24804,N_21887);
or U29858 (N_29858,N_23938,N_24296);
xor U29859 (N_29859,N_20121,N_20962);
nor U29860 (N_29860,N_24320,N_24933);
nor U29861 (N_29861,N_23140,N_20526);
and U29862 (N_29862,N_20963,N_24445);
nor U29863 (N_29863,N_20701,N_20160);
nor U29864 (N_29864,N_23168,N_21990);
xor U29865 (N_29865,N_20141,N_21625);
nand U29866 (N_29866,N_21823,N_24504);
and U29867 (N_29867,N_24799,N_22289);
and U29868 (N_29868,N_24954,N_24137);
and U29869 (N_29869,N_20728,N_23483);
nand U29870 (N_29870,N_21415,N_24085);
nor U29871 (N_29871,N_22536,N_22709);
or U29872 (N_29872,N_24274,N_23742);
or U29873 (N_29873,N_21915,N_20145);
or U29874 (N_29874,N_22353,N_20354);
nor U29875 (N_29875,N_23872,N_23388);
and U29876 (N_29876,N_23846,N_20926);
nand U29877 (N_29877,N_22994,N_21955);
xor U29878 (N_29878,N_24965,N_20199);
and U29879 (N_29879,N_22931,N_24272);
nor U29880 (N_29880,N_24479,N_20574);
nor U29881 (N_29881,N_23281,N_24657);
and U29882 (N_29882,N_21590,N_24284);
or U29883 (N_29883,N_22575,N_23577);
or U29884 (N_29884,N_24714,N_22539);
or U29885 (N_29885,N_22010,N_22140);
and U29886 (N_29886,N_21197,N_20078);
and U29887 (N_29887,N_20876,N_24393);
or U29888 (N_29888,N_21516,N_24079);
or U29889 (N_29889,N_20658,N_22250);
nor U29890 (N_29890,N_23553,N_21825);
nand U29891 (N_29891,N_22350,N_20649);
nor U29892 (N_29892,N_21278,N_22123);
xnor U29893 (N_29893,N_20548,N_22766);
nand U29894 (N_29894,N_24328,N_23601);
nand U29895 (N_29895,N_22199,N_23861);
nand U29896 (N_29896,N_24593,N_23425);
nand U29897 (N_29897,N_23734,N_23694);
and U29898 (N_29898,N_24033,N_21114);
and U29899 (N_29899,N_21632,N_20279);
nand U29900 (N_29900,N_24600,N_24115);
or U29901 (N_29901,N_22688,N_21584);
nand U29902 (N_29902,N_24234,N_21724);
and U29903 (N_29903,N_22474,N_24954);
nor U29904 (N_29904,N_24994,N_23532);
xor U29905 (N_29905,N_23991,N_22736);
nand U29906 (N_29906,N_23486,N_20562);
nor U29907 (N_29907,N_23424,N_20263);
xnor U29908 (N_29908,N_20732,N_22584);
nor U29909 (N_29909,N_24600,N_23348);
nor U29910 (N_29910,N_20858,N_21633);
and U29911 (N_29911,N_23589,N_21020);
nand U29912 (N_29912,N_24597,N_20575);
nand U29913 (N_29913,N_23778,N_24179);
nor U29914 (N_29914,N_21595,N_20304);
xor U29915 (N_29915,N_22849,N_21892);
and U29916 (N_29916,N_21687,N_23445);
and U29917 (N_29917,N_23183,N_21176);
nor U29918 (N_29918,N_23741,N_21536);
and U29919 (N_29919,N_23756,N_23263);
nand U29920 (N_29920,N_20553,N_20064);
nor U29921 (N_29921,N_24632,N_22365);
and U29922 (N_29922,N_20133,N_22714);
or U29923 (N_29923,N_21712,N_21421);
and U29924 (N_29924,N_20555,N_23631);
nand U29925 (N_29925,N_24232,N_21328);
or U29926 (N_29926,N_21966,N_20349);
nand U29927 (N_29927,N_20401,N_22895);
and U29928 (N_29928,N_22791,N_20465);
or U29929 (N_29929,N_20764,N_24572);
xnor U29930 (N_29930,N_24512,N_20272);
nand U29931 (N_29931,N_21738,N_23285);
nor U29932 (N_29932,N_22580,N_23277);
nor U29933 (N_29933,N_22479,N_20873);
or U29934 (N_29934,N_24759,N_23132);
nor U29935 (N_29935,N_22499,N_20893);
or U29936 (N_29936,N_24200,N_21587);
xor U29937 (N_29937,N_21205,N_24499);
and U29938 (N_29938,N_20479,N_20182);
and U29939 (N_29939,N_24258,N_23035);
or U29940 (N_29940,N_24741,N_21231);
or U29941 (N_29941,N_20948,N_21265);
nor U29942 (N_29942,N_22730,N_20541);
nand U29943 (N_29943,N_22632,N_22704);
nor U29944 (N_29944,N_24103,N_21975);
nor U29945 (N_29945,N_24097,N_22192);
nand U29946 (N_29946,N_20434,N_20686);
and U29947 (N_29947,N_20830,N_24012);
nand U29948 (N_29948,N_24029,N_22959);
nor U29949 (N_29949,N_20514,N_24842);
nor U29950 (N_29950,N_23240,N_24668);
or U29951 (N_29951,N_24550,N_20417);
and U29952 (N_29952,N_23663,N_22152);
nand U29953 (N_29953,N_20553,N_24414);
and U29954 (N_29954,N_24801,N_22196);
and U29955 (N_29955,N_21202,N_21998);
nor U29956 (N_29956,N_21363,N_21886);
nor U29957 (N_29957,N_21683,N_20306);
or U29958 (N_29958,N_22958,N_20940);
xnor U29959 (N_29959,N_24213,N_23967);
nor U29960 (N_29960,N_21508,N_21053);
or U29961 (N_29961,N_20783,N_24025);
nor U29962 (N_29962,N_22170,N_22313);
or U29963 (N_29963,N_23807,N_22356);
nand U29964 (N_29964,N_23502,N_23563);
and U29965 (N_29965,N_21529,N_21689);
nor U29966 (N_29966,N_23902,N_24953);
nor U29967 (N_29967,N_22578,N_24179);
or U29968 (N_29968,N_24529,N_21477);
nand U29969 (N_29969,N_20380,N_20032);
or U29970 (N_29970,N_23930,N_23207);
or U29971 (N_29971,N_24543,N_24932);
or U29972 (N_29972,N_20048,N_20385);
nor U29973 (N_29973,N_20913,N_21535);
nand U29974 (N_29974,N_23444,N_24800);
or U29975 (N_29975,N_21322,N_21944);
xor U29976 (N_29976,N_20659,N_24233);
nand U29977 (N_29977,N_21669,N_23037);
and U29978 (N_29978,N_21305,N_23360);
and U29979 (N_29979,N_21593,N_24270);
nor U29980 (N_29980,N_24396,N_24806);
nand U29981 (N_29981,N_21899,N_21539);
or U29982 (N_29982,N_24187,N_24430);
xor U29983 (N_29983,N_24318,N_20864);
nor U29984 (N_29984,N_23321,N_23707);
and U29985 (N_29985,N_20825,N_24842);
xnor U29986 (N_29986,N_20685,N_24387);
xnor U29987 (N_29987,N_24499,N_23429);
nand U29988 (N_29988,N_21673,N_23724);
and U29989 (N_29989,N_24245,N_20831);
nor U29990 (N_29990,N_20890,N_24266);
nor U29991 (N_29991,N_20689,N_20533);
nand U29992 (N_29992,N_20763,N_23367);
or U29993 (N_29993,N_23480,N_20576);
nand U29994 (N_29994,N_23941,N_20133);
nor U29995 (N_29995,N_21675,N_20984);
nor U29996 (N_29996,N_22478,N_22017);
xnor U29997 (N_29997,N_21278,N_24573);
or U29998 (N_29998,N_21337,N_24227);
nor U29999 (N_29999,N_20193,N_22458);
nand U30000 (N_30000,N_28668,N_27614);
or U30001 (N_30001,N_26312,N_26325);
or U30002 (N_30002,N_26216,N_28399);
nor U30003 (N_30003,N_27991,N_29695);
or U30004 (N_30004,N_25157,N_25235);
xor U30005 (N_30005,N_26439,N_28437);
or U30006 (N_30006,N_29912,N_27325);
and U30007 (N_30007,N_29968,N_27288);
or U30008 (N_30008,N_27535,N_27053);
xor U30009 (N_30009,N_29407,N_29153);
and U30010 (N_30010,N_27407,N_25467);
nor U30011 (N_30011,N_27012,N_27501);
or U30012 (N_30012,N_28949,N_26597);
or U30013 (N_30013,N_27322,N_27323);
nor U30014 (N_30014,N_26875,N_29477);
or U30015 (N_30015,N_28475,N_26829);
nand U30016 (N_30016,N_25876,N_28185);
or U30017 (N_30017,N_25315,N_29907);
or U30018 (N_30018,N_27234,N_29592);
xnor U30019 (N_30019,N_27912,N_28541);
or U30020 (N_30020,N_26672,N_26777);
and U30021 (N_30021,N_27030,N_27090);
nand U30022 (N_30022,N_26964,N_27410);
nand U30023 (N_30023,N_29213,N_28832);
xor U30024 (N_30024,N_28096,N_29406);
nand U30025 (N_30025,N_25763,N_26801);
and U30026 (N_30026,N_27602,N_27633);
or U30027 (N_30027,N_25228,N_25997);
and U30028 (N_30028,N_28895,N_27526);
xor U30029 (N_30029,N_25522,N_28643);
or U30030 (N_30030,N_29783,N_29613);
nor U30031 (N_30031,N_28382,N_28056);
and U30032 (N_30032,N_28615,N_27400);
nor U30033 (N_30033,N_29645,N_27770);
nor U30034 (N_30034,N_27838,N_25286);
or U30035 (N_30035,N_27779,N_28024);
nor U30036 (N_30036,N_28893,N_29403);
nand U30037 (N_30037,N_29004,N_27000);
or U30038 (N_30038,N_27295,N_27514);
nand U30039 (N_30039,N_27853,N_29979);
and U30040 (N_30040,N_25206,N_25111);
nor U30041 (N_30041,N_27125,N_25463);
or U30042 (N_30042,N_28568,N_25555);
or U30043 (N_30043,N_25008,N_29545);
nor U30044 (N_30044,N_27013,N_28301);
nand U30045 (N_30045,N_28520,N_28502);
nand U30046 (N_30046,N_28523,N_27371);
nor U30047 (N_30047,N_28504,N_27472);
nor U30048 (N_30048,N_27861,N_28344);
nand U30049 (N_30049,N_29687,N_29191);
and U30050 (N_30050,N_26102,N_25551);
and U30051 (N_30051,N_27046,N_29696);
and U30052 (N_30052,N_25666,N_29996);
nor U30053 (N_30053,N_29821,N_25149);
or U30054 (N_30054,N_29866,N_27625);
nor U30055 (N_30055,N_26244,N_28148);
or U30056 (N_30056,N_25546,N_28232);
xnor U30057 (N_30057,N_27651,N_29629);
and U30058 (N_30058,N_27554,N_27675);
xnor U30059 (N_30059,N_29003,N_25353);
and U30060 (N_30060,N_27233,N_25490);
or U30061 (N_30061,N_26438,N_28571);
nor U30062 (N_30062,N_29914,N_26568);
nor U30063 (N_30063,N_27668,N_27930);
nand U30064 (N_30064,N_25853,N_29117);
and U30065 (N_30065,N_29539,N_27771);
nand U30066 (N_30066,N_29529,N_26121);
or U30067 (N_30067,N_25545,N_27256);
or U30068 (N_30068,N_26302,N_28273);
nand U30069 (N_30069,N_26646,N_26081);
and U30070 (N_30070,N_29697,N_27852);
and U30071 (N_30071,N_28872,N_28368);
or U30072 (N_30072,N_29279,N_27845);
and U30073 (N_30073,N_26224,N_26936);
and U30074 (N_30074,N_26207,N_25694);
xnor U30075 (N_30075,N_29130,N_29802);
nor U30076 (N_30076,N_26600,N_28076);
xor U30077 (N_30077,N_27654,N_29465);
nor U30078 (N_30078,N_26894,N_28270);
nand U30079 (N_30079,N_29324,N_25476);
and U30080 (N_30080,N_25651,N_27619);
or U30081 (N_30081,N_27333,N_25242);
and U30082 (N_30082,N_25814,N_26677);
nand U30083 (N_30083,N_28563,N_29535);
nand U30084 (N_30084,N_27616,N_26401);
nand U30085 (N_30085,N_25057,N_29329);
or U30086 (N_30086,N_26729,N_25123);
and U30087 (N_30087,N_26410,N_27034);
nor U30088 (N_30088,N_25083,N_26778);
and U30089 (N_30089,N_28440,N_29047);
or U30090 (N_30090,N_27995,N_25882);
nor U30091 (N_30091,N_28445,N_25054);
nand U30092 (N_30092,N_28623,N_25274);
nand U30093 (N_30093,N_26124,N_29152);
nand U30094 (N_30094,N_27883,N_25731);
and U30095 (N_30095,N_25851,N_27927);
nand U30096 (N_30096,N_25475,N_28835);
nor U30097 (N_30097,N_25493,N_27521);
nor U30098 (N_30098,N_26859,N_28091);
nand U30099 (N_30099,N_25167,N_25162);
nor U30100 (N_30100,N_29573,N_26067);
nand U30101 (N_30101,N_25255,N_28870);
nand U30102 (N_30102,N_29876,N_28197);
and U30103 (N_30103,N_28194,N_25841);
nand U30104 (N_30104,N_28791,N_26132);
or U30105 (N_30105,N_27385,N_26549);
nor U30106 (N_30106,N_27279,N_27511);
nand U30107 (N_30107,N_27058,N_27156);
and U30108 (N_30108,N_26363,N_28983);
nand U30109 (N_30109,N_25730,N_29328);
and U30110 (N_30110,N_26079,N_25676);
xnor U30111 (N_30111,N_28287,N_29228);
nand U30112 (N_30112,N_26743,N_27940);
or U30113 (N_30113,N_27271,N_25403);
and U30114 (N_30114,N_25072,N_28579);
and U30115 (N_30115,N_25124,N_25889);
nor U30116 (N_30116,N_27448,N_28325);
nand U30117 (N_30117,N_26021,N_28708);
and U30118 (N_30118,N_29026,N_27674);
nand U30119 (N_30119,N_29286,N_27122);
nand U30120 (N_30120,N_25288,N_28010);
and U30121 (N_30121,N_29584,N_29693);
and U30122 (N_30122,N_25019,N_29437);
xor U30123 (N_30123,N_29146,N_28365);
and U30124 (N_30124,N_26052,N_29079);
nor U30125 (N_30125,N_27782,N_29708);
nand U30126 (N_30126,N_28849,N_25899);
nand U30127 (N_30127,N_25745,N_25334);
nor U30128 (N_30128,N_25070,N_27294);
and U30129 (N_30129,N_29169,N_28514);
and U30130 (N_30130,N_27490,N_27921);
xor U30131 (N_30131,N_28604,N_29461);
nand U30132 (N_30132,N_29847,N_27959);
nand U30133 (N_30133,N_26267,N_27911);
and U30134 (N_30134,N_28317,N_27207);
xnor U30135 (N_30135,N_26058,N_25570);
xnor U30136 (N_30136,N_27438,N_29810);
nand U30137 (N_30137,N_28754,N_26807);
or U30138 (N_30138,N_28155,N_28200);
xor U30139 (N_30139,N_29943,N_28316);
xnor U30140 (N_30140,N_26745,N_26335);
xor U30141 (N_30141,N_25923,N_26557);
and U30142 (N_30142,N_28596,N_29897);
nor U30143 (N_30143,N_27548,N_27937);
and U30144 (N_30144,N_28114,N_26817);
and U30145 (N_30145,N_29910,N_28924);
or U30146 (N_30146,N_25603,N_27834);
or U30147 (N_30147,N_27923,N_25971);
xnor U30148 (N_30148,N_26365,N_29400);
nand U30149 (N_30149,N_29640,N_28733);
or U30150 (N_30150,N_26956,N_28116);
nand U30151 (N_30151,N_29187,N_28865);
or U30152 (N_30152,N_28456,N_26865);
nor U30153 (N_30153,N_28191,N_27855);
and U30154 (N_30154,N_29482,N_29395);
xnor U30155 (N_30155,N_26562,N_25238);
nor U30156 (N_30156,N_25652,N_27813);
or U30157 (N_30157,N_28858,N_28080);
xnor U30158 (N_30158,N_26442,N_28144);
and U30159 (N_30159,N_26272,N_26576);
nand U30160 (N_30160,N_29142,N_27831);
nand U30161 (N_30161,N_27981,N_26403);
and U30162 (N_30162,N_25193,N_27347);
nor U30163 (N_30163,N_28515,N_27127);
or U30164 (N_30164,N_29501,N_27359);
and U30165 (N_30165,N_27310,N_25819);
xnor U30166 (N_30166,N_28166,N_29938);
or U30167 (N_30167,N_27306,N_27904);
nand U30168 (N_30168,N_29772,N_28052);
and U30169 (N_30169,N_28500,N_29918);
nand U30170 (N_30170,N_26627,N_29372);
nor U30171 (N_30171,N_25892,N_29956);
nand U30172 (N_30172,N_25576,N_28640);
nand U30173 (N_30173,N_25950,N_29068);
or U30174 (N_30174,N_25789,N_28731);
nand U30175 (N_30175,N_29426,N_28485);
nand U30176 (N_30176,N_26504,N_25252);
xnor U30177 (N_30177,N_25964,N_26912);
nand U30178 (N_30178,N_27494,N_27055);
nor U30179 (N_30179,N_26113,N_29063);
and U30180 (N_30180,N_26937,N_25588);
nor U30181 (N_30181,N_28262,N_25374);
or U30182 (N_30182,N_28120,N_27048);
and U30183 (N_30183,N_29899,N_25223);
nand U30184 (N_30184,N_26708,N_29973);
and U30185 (N_30185,N_28291,N_28705);
or U30186 (N_30186,N_28066,N_25456);
xnor U30187 (N_30187,N_29417,N_28956);
and U30188 (N_30188,N_26433,N_25535);
or U30189 (N_30189,N_27611,N_29811);
nand U30190 (N_30190,N_28054,N_29302);
or U30191 (N_30191,N_25795,N_27399);
nand U30192 (N_30192,N_29638,N_27082);
nand U30193 (N_30193,N_26001,N_29944);
or U30194 (N_30194,N_28690,N_29633);
nor U30195 (N_30195,N_25412,N_28797);
and U30196 (N_30196,N_28356,N_26157);
xnor U30197 (N_30197,N_25702,N_27748);
nor U30198 (N_30198,N_29649,N_26714);
or U30199 (N_30199,N_28825,N_29744);
nand U30200 (N_30200,N_26934,N_28109);
nor U30201 (N_30201,N_25630,N_26941);
and U30202 (N_30202,N_27255,N_26942);
nor U30203 (N_30203,N_28543,N_25257);
nand U30204 (N_30204,N_28049,N_29340);
and U30205 (N_30205,N_28821,N_28026);
nor U30206 (N_30206,N_27394,N_29591);
nand U30207 (N_30207,N_29597,N_27678);
or U30208 (N_30208,N_27257,N_27142);
nor U30209 (N_30209,N_28810,N_28288);
nand U30210 (N_30210,N_28946,N_28412);
and U30211 (N_30211,N_26542,N_28868);
or U30212 (N_30212,N_27309,N_25655);
nand U30213 (N_30213,N_27725,N_26608);
nand U30214 (N_30214,N_27237,N_29048);
and U30215 (N_30215,N_25345,N_26965);
nor U30216 (N_30216,N_26811,N_27280);
and U30217 (N_30217,N_27499,N_27057);
and U30218 (N_30218,N_27168,N_27839);
nor U30219 (N_30219,N_27003,N_25328);
and U30220 (N_30220,N_28261,N_29136);
or U30221 (N_30221,N_26226,N_26767);
nand U30222 (N_30222,N_25437,N_28777);
or U30223 (N_30223,N_25442,N_28885);
nand U30224 (N_30224,N_29605,N_25880);
nand U30225 (N_30225,N_27327,N_26828);
and U30226 (N_30226,N_29768,N_26285);
and U30227 (N_30227,N_25485,N_28905);
xor U30228 (N_30228,N_25218,N_28195);
nand U30229 (N_30229,N_25126,N_26586);
and U30230 (N_30230,N_28628,N_28510);
xor U30231 (N_30231,N_26200,N_26196);
and U30232 (N_30232,N_26279,N_25216);
nand U30233 (N_30233,N_27235,N_25727);
or U30234 (N_30234,N_29019,N_26169);
nor U30235 (N_30235,N_26088,N_26111);
and U30236 (N_30236,N_26928,N_27020);
xnor U30237 (N_30237,N_29243,N_27687);
and U30238 (N_30238,N_28004,N_26493);
nor U30239 (N_30239,N_26883,N_26949);
or U30240 (N_30240,N_29483,N_26703);
or U30241 (N_30241,N_27968,N_26042);
and U30242 (N_30242,N_27693,N_25616);
and U30243 (N_30243,N_25956,N_28931);
nand U30244 (N_30244,N_26037,N_28855);
and U30245 (N_30245,N_28400,N_25130);
nand U30246 (N_30246,N_27998,N_27364);
or U30247 (N_30247,N_28940,N_26227);
and U30248 (N_30248,N_27740,N_27485);
nand U30249 (N_30249,N_26802,N_28888);
or U30250 (N_30250,N_26149,N_28136);
or U30251 (N_30251,N_26559,N_29497);
nor U30252 (N_30252,N_27598,N_27580);
nand U30253 (N_30253,N_29347,N_27567);
nor U30254 (N_30254,N_28994,N_25679);
nor U30255 (N_30255,N_25253,N_26793);
and U30256 (N_30256,N_25716,N_25271);
nand U30257 (N_30257,N_25842,N_26835);
and U30258 (N_30258,N_29856,N_27713);
nand U30259 (N_30259,N_25532,N_25049);
and U30260 (N_30260,N_27973,N_28724);
nand U30261 (N_30261,N_29904,N_26593);
or U30262 (N_30262,N_27111,N_29265);
nand U30263 (N_30263,N_27964,N_26399);
and U30264 (N_30264,N_28521,N_28404);
or U30265 (N_30265,N_26585,N_29870);
or U30266 (N_30266,N_28844,N_28338);
and U30267 (N_30267,N_27197,N_27115);
nor U30268 (N_30268,N_28496,N_29602);
nor U30269 (N_30269,N_27471,N_28373);
and U30270 (N_30270,N_29257,N_25575);
and U30271 (N_30271,N_25848,N_26718);
and U30272 (N_30272,N_28511,N_28345);
and U30273 (N_30273,N_25232,N_25265);
or U30274 (N_30274,N_27608,N_26023);
nand U30275 (N_30275,N_29746,N_26167);
xnor U30276 (N_30276,N_28419,N_29860);
nand U30277 (N_30277,N_25903,N_29852);
and U30278 (N_30278,N_25395,N_26753);
nor U30279 (N_30279,N_25718,N_28003);
xor U30280 (N_30280,N_26298,N_26156);
nand U30281 (N_30281,N_29014,N_26044);
and U30282 (N_30282,N_25712,N_26693);
nor U30283 (N_30283,N_25658,N_28002);
xnor U30284 (N_30284,N_26142,N_27300);
nor U30285 (N_30285,N_26237,N_27947);
nand U30286 (N_30286,N_28546,N_29727);
nand U30287 (N_30287,N_28472,N_27604);
nand U30288 (N_30288,N_27434,N_27768);
nand U30289 (N_30289,N_29289,N_27769);
and U30290 (N_30290,N_28410,N_26151);
or U30291 (N_30291,N_29678,N_25700);
and U30292 (N_30292,N_26755,N_27832);
or U30293 (N_30293,N_29832,N_27318);
nor U30294 (N_30294,N_26465,N_25947);
and U30295 (N_30295,N_25267,N_29601);
nor U30296 (N_30296,N_25055,N_25349);
and U30297 (N_30297,N_29900,N_29745);
or U30298 (N_30298,N_27252,N_29000);
nor U30299 (N_30299,N_28451,N_28058);
xor U30300 (N_30300,N_27277,N_28603);
nor U30301 (N_30301,N_25972,N_28675);
or U30302 (N_30302,N_26223,N_27098);
nand U30303 (N_30303,N_25317,N_27314);
or U30304 (N_30304,N_25689,N_26725);
nand U30305 (N_30305,N_25553,N_29058);
and U30306 (N_30306,N_29015,N_29258);
nand U30307 (N_30307,N_25583,N_28303);
xor U30308 (N_30308,N_28517,N_26214);
nand U30309 (N_30309,N_25767,N_26491);
nand U30310 (N_30310,N_28182,N_25517);
nand U30311 (N_30311,N_29794,N_25392);
nand U30312 (N_30312,N_25708,N_25806);
and U30313 (N_30313,N_25414,N_28110);
and U30314 (N_30314,N_29728,N_29814);
and U30315 (N_30315,N_29225,N_27649);
and U30316 (N_30316,N_27741,N_27458);
xnor U30317 (N_30317,N_27763,N_26183);
and U30318 (N_30318,N_28219,N_29023);
xor U30319 (N_30319,N_26419,N_29951);
or U30320 (N_30320,N_26686,N_29223);
nor U30321 (N_30321,N_26575,N_29724);
and U30322 (N_30322,N_28359,N_29418);
nand U30323 (N_30323,N_25420,N_29127);
xnor U30324 (N_30324,N_26241,N_29032);
xor U30325 (N_30325,N_26641,N_25015);
and U30326 (N_30326,N_29186,N_28830);
nor U30327 (N_30327,N_26843,N_27274);
nand U30328 (N_30328,N_29361,N_28390);
and U30329 (N_30329,N_25901,N_28130);
or U30330 (N_30330,N_25753,N_29261);
xnor U30331 (N_30331,N_26570,N_28898);
and U30332 (N_30332,N_26440,N_28146);
nand U30333 (N_30333,N_28306,N_28713);
or U30334 (N_30334,N_29123,N_26374);
and U30335 (N_30335,N_27119,N_27095);
and U30336 (N_30336,N_28165,N_28577);
or U30337 (N_30337,N_25134,N_27109);
nor U30338 (N_30338,N_28917,N_26523);
nor U30339 (N_30339,N_29472,N_25687);
xor U30340 (N_30340,N_25991,N_27022);
nand U30341 (N_30341,N_29763,N_29537);
nor U30342 (N_30342,N_27896,N_25635);
and U30343 (N_30343,N_26300,N_25941);
and U30344 (N_30344,N_27663,N_28164);
or U30345 (N_30345,N_27077,N_26616);
nand U30346 (N_30346,N_29466,N_29504);
nor U30347 (N_30347,N_25344,N_28661);
nor U30348 (N_30348,N_26842,N_27146);
nor U30349 (N_30349,N_27129,N_27064);
xor U30350 (N_30350,N_27530,N_27374);
nand U30351 (N_30351,N_26343,N_28282);
nor U30352 (N_30352,N_29614,N_25074);
and U30353 (N_30353,N_28309,N_26806);
nor U30354 (N_30354,N_28285,N_28386);
or U30355 (N_30355,N_28424,N_27751);
or U30356 (N_30356,N_28939,N_25381);
and U30357 (N_30357,N_28237,N_25402);
nand U30358 (N_30358,N_25510,N_27391);
and U30359 (N_30359,N_25574,N_27902);
nor U30360 (N_30360,N_26594,N_29960);
or U30361 (N_30361,N_28216,N_29433);
and U30362 (N_30362,N_29098,N_26235);
or U30363 (N_30363,N_27583,N_29074);
and U30364 (N_30364,N_28240,N_26610);
and U30365 (N_30365,N_25783,N_28245);
nand U30366 (N_30366,N_25106,N_29885);
and U30367 (N_30367,N_29339,N_28297);
or U30368 (N_30368,N_29806,N_28021);
xnor U30369 (N_30369,N_28957,N_25406);
or U30370 (N_30370,N_25781,N_29923);
nand U30371 (N_30371,N_26890,N_25549);
nand U30372 (N_30372,N_27334,N_28747);
nand U30373 (N_30373,N_28207,N_27155);
and U30374 (N_30374,N_27215,N_26952);
nand U30375 (N_30375,N_29519,N_28544);
and U30376 (N_30376,N_28986,N_27384);
nor U30377 (N_30377,N_26376,N_28428);
or U30378 (N_30378,N_25656,N_27764);
nand U30379 (N_30379,N_25204,N_26683);
nor U30380 (N_30380,N_29726,N_25186);
or U30381 (N_30381,N_27958,N_28012);
and U30382 (N_30382,N_29062,N_26069);
or U30383 (N_30383,N_28343,N_27942);
nand U30384 (N_30384,N_26754,N_28457);
nand U30385 (N_30385,N_25075,N_29307);
and U30386 (N_30386,N_25294,N_27868);
or U30387 (N_30387,N_27781,N_25031);
nand U30388 (N_30388,N_26792,N_29589);
or U30389 (N_30389,N_27933,N_27076);
and U30390 (N_30390,N_29654,N_25878);
or U30391 (N_30391,N_25040,N_26996);
and U30392 (N_30392,N_26269,N_28658);
nand U30393 (N_30393,N_26961,N_26915);
and U30394 (N_30394,N_25314,N_29970);
nand U30395 (N_30395,N_28224,N_26876);
or U30396 (N_30396,N_26676,N_26263);
or U30397 (N_30397,N_27085,N_26704);
nor U30398 (N_30398,N_26342,N_29318);
or U30399 (N_30399,N_29809,N_29942);
nor U30400 (N_30400,N_28226,N_26369);
or U30401 (N_30401,N_29121,N_25813);
nor U30402 (N_30402,N_26716,N_26389);
or U30403 (N_30403,N_25980,N_27819);
nor U30404 (N_30404,N_27568,N_27954);
nor U30405 (N_30405,N_28607,N_27081);
nand U30406 (N_30406,N_29366,N_26247);
nor U30407 (N_30407,N_25222,N_28423);
xor U30408 (N_30408,N_26870,N_26667);
or U30409 (N_30409,N_27453,N_26230);
and U30410 (N_30410,N_27996,N_27481);
or U30411 (N_30411,N_29369,N_26741);
nand U30412 (N_30412,N_26946,N_27411);
or U30413 (N_30413,N_29341,N_28599);
and U30414 (N_30414,N_27899,N_25135);
or U30415 (N_30415,N_25062,N_27035);
or U30416 (N_30416,N_26840,N_26662);
nand U30417 (N_30417,N_29830,N_29868);
nand U30418 (N_30418,N_29112,N_29932);
nor U30419 (N_30419,N_27908,N_25478);
nor U30420 (N_30420,N_29757,N_29959);
xnor U30421 (N_30421,N_25618,N_25452);
or U30422 (N_30422,N_29997,N_29698);
or U30423 (N_30423,N_26719,N_26731);
and U30424 (N_30424,N_29540,N_26100);
nand U30425 (N_30425,N_26752,N_27075);
nor U30426 (N_30426,N_26906,N_29270);
or U30427 (N_30427,N_26359,N_27662);
xnor U30428 (N_30428,N_29217,N_29093);
xnor U30429 (N_30429,N_28234,N_29829);
nor U30430 (N_30430,N_25936,N_27375);
or U30431 (N_30431,N_27259,N_26879);
or U30432 (N_30432,N_27049,N_26611);
and U30433 (N_30433,N_27339,N_27823);
nand U30434 (N_30434,N_27766,N_25366);
and U30435 (N_30435,N_25845,N_26854);
nor U30436 (N_30436,N_28582,N_28394);
or U30437 (N_30437,N_29303,N_29424);
and U30438 (N_30438,N_29070,N_26947);
nand U30439 (N_30439,N_25775,N_26799);
nor U30440 (N_30440,N_29616,N_25208);
nand U30441 (N_30441,N_26525,N_29374);
nor U30442 (N_30442,N_27355,N_26295);
and U30443 (N_30443,N_25804,N_28474);
xor U30444 (N_30444,N_27158,N_26138);
or U30445 (N_30445,N_26323,N_29262);
nor U30446 (N_30446,N_27017,N_28536);
nor U30447 (N_30447,N_28086,N_27907);
or U30448 (N_30448,N_28890,N_29521);
and U30449 (N_30449,N_26759,N_28103);
nor U30450 (N_30450,N_29201,N_29679);
nand U30451 (N_30451,N_28757,N_28072);
nand U30452 (N_30452,N_28315,N_26234);
and U30453 (N_30453,N_25400,N_28831);
and U30454 (N_30454,N_29511,N_26978);
nor U30455 (N_30455,N_25047,N_27154);
nor U30456 (N_30456,N_25958,N_27950);
nand U30457 (N_30457,N_26950,N_25102);
and U30458 (N_30458,N_28566,N_26563);
nor U30459 (N_30459,N_26476,N_26039);
or U30460 (N_30460,N_25828,N_29881);
nor U30461 (N_30461,N_25489,N_29385);
nand U30462 (N_30462,N_27424,N_29214);
nor U30463 (N_30463,N_27556,N_26004);
nor U30464 (N_30464,N_26853,N_27767);
nor U30465 (N_30465,N_28214,N_27993);
or U30466 (N_30466,N_25837,N_29087);
or U30467 (N_30467,N_29530,N_26733);
and U30468 (N_30468,N_27532,N_27588);
xor U30469 (N_30469,N_29456,N_29008);
nand U30470 (N_30470,N_28749,N_25087);
or U30471 (N_30471,N_25843,N_26728);
and U30472 (N_30472,N_25965,N_28729);
or U30473 (N_30473,N_29758,N_29204);
and U30474 (N_30474,N_25300,N_25884);
nand U30475 (N_30475,N_25823,N_25338);
and U30476 (N_30476,N_29842,N_26578);
nand U30477 (N_30477,N_29219,N_25132);
nand U30478 (N_30478,N_28498,N_25627);
xor U30479 (N_30479,N_26197,N_27478);
xnor U30480 (N_30480,N_29025,N_28296);
xor U30481 (N_30481,N_28829,N_29484);
nor U30482 (N_30482,N_26836,N_29450);
nand U30483 (N_30483,N_26604,N_28698);
nand U30484 (N_30484,N_25534,N_26109);
and U30485 (N_30485,N_29921,N_26094);
nor U30486 (N_30486,N_27698,N_29609);
or U30487 (N_30487,N_28763,N_29298);
nand U30488 (N_30488,N_27317,N_27380);
nor U30489 (N_30489,N_28095,N_28680);
nand U30490 (N_30490,N_27820,N_26707);
and U30491 (N_30491,N_25784,N_25335);
or U30492 (N_30492,N_26909,N_27412);
nand U30493 (N_30493,N_26756,N_25917);
nor U30494 (N_30494,N_26533,N_29875);
nand U30495 (N_30495,N_26082,N_28249);
or U30496 (N_30496,N_25113,N_25082);
and U30497 (N_30497,N_27623,N_25698);
xor U30498 (N_30498,N_28339,N_26329);
nand U30499 (N_30499,N_25017,N_25127);
or U30500 (N_30500,N_29854,N_28070);
and U30501 (N_30501,N_25231,N_26739);
and U30502 (N_30502,N_27920,N_25359);
nor U30503 (N_30503,N_27586,N_27629);
nand U30504 (N_30504,N_26872,N_25439);
or U30505 (N_30505,N_27824,N_26122);
or U30506 (N_30506,N_25161,N_29065);
nor U30507 (N_30507,N_25750,N_26639);
nor U30508 (N_30508,N_25166,N_25121);
xor U30509 (N_30509,N_27716,N_27979);
or U30510 (N_30510,N_29402,N_26489);
and U30511 (N_30511,N_28828,N_25112);
and U30512 (N_30512,N_25954,N_29132);
nand U30513 (N_30513,N_27343,N_26957);
or U30514 (N_30514,N_26921,N_28375);
or U30515 (N_30515,N_26140,N_29163);
or U30516 (N_30516,N_25939,N_28540);
or U30517 (N_30517,N_26488,N_28793);
xor U30518 (N_30518,N_27204,N_25100);
xor U30519 (N_30519,N_28787,N_28413);
nand U30520 (N_30520,N_25868,N_29946);
or U30521 (N_30521,N_27413,N_27963);
nand U30522 (N_30522,N_26047,N_29976);
nor U30523 (N_30523,N_27903,N_26195);
xnor U30524 (N_30524,N_29651,N_25337);
nand U30525 (N_30525,N_28342,N_28837);
and U30526 (N_30526,N_29884,N_25101);
nor U30527 (N_30527,N_25719,N_25085);
and U30528 (N_30528,N_27225,N_26882);
or U30529 (N_30529,N_29677,N_26596);
nor U30530 (N_30530,N_25262,N_26818);
nor U30531 (N_30531,N_25190,N_28903);
or U30532 (N_30532,N_25474,N_29664);
nand U30533 (N_30533,N_25292,N_29423);
nor U30534 (N_30534,N_27231,N_27179);
xnor U30535 (N_30535,N_28927,N_28463);
nand U30536 (N_30536,N_26571,N_25890);
or U30537 (N_30537,N_28402,N_27479);
or U30538 (N_30538,N_29336,N_25913);
xnor U30539 (N_30539,N_25037,N_26176);
nand U30540 (N_30540,N_28213,N_26400);
or U30541 (N_30541,N_29334,N_27346);
nor U30542 (N_30542,N_29919,N_28970);
or U30543 (N_30543,N_27862,N_27516);
nor U30544 (N_30544,N_28719,N_26322);
nand U30545 (N_30545,N_27040,N_26344);
nor U30546 (N_30546,N_27178,N_27916);
nand U30547 (N_30547,N_26250,N_28387);
xnor U30548 (N_30548,N_28930,N_25409);
xor U30549 (N_30549,N_25289,N_29934);
and U30550 (N_30550,N_29115,N_25654);
nand U30551 (N_30551,N_26724,N_27468);
and U30552 (N_30552,N_26927,N_29165);
nor U30553 (N_30553,N_27607,N_25924);
and U30554 (N_30554,N_29156,N_29428);
and U30555 (N_30555,N_25852,N_27701);
or U30556 (N_30556,N_28826,N_28686);
and U30557 (N_30557,N_25805,N_26904);
or U30558 (N_30558,N_29524,N_28906);
nand U30559 (N_30559,N_26880,N_25026);
and U30560 (N_30560,N_25625,N_26848);
xnor U30561 (N_30561,N_27476,N_27910);
or U30562 (N_30562,N_28716,N_29380);
and U30563 (N_30563,N_26415,N_25771);
and U30564 (N_30564,N_28531,N_26896);
nor U30565 (N_30565,N_28794,N_27537);
nand U30566 (N_30566,N_27007,N_27791);
xor U30567 (N_30567,N_27070,N_28633);
or U30568 (N_30568,N_25361,N_26632);
nor U30569 (N_30569,N_25770,N_29056);
nor U30570 (N_30570,N_27004,N_29050);
and U30571 (N_30571,N_28815,N_25948);
nor U30572 (N_30572,N_25239,N_28174);
nand U30573 (N_30573,N_26080,N_28124);
xor U30574 (N_30574,N_27444,N_28611);
or U30575 (N_30575,N_26057,N_25854);
or U30576 (N_30576,N_26572,N_29297);
and U30577 (N_30577,N_28648,N_29012);
and U30578 (N_30578,N_27794,N_27504);
nand U30579 (N_30579,N_28998,N_29906);
nor U30580 (N_30580,N_28178,N_28391);
and U30581 (N_30581,N_26056,N_25711);
nand U30582 (N_30582,N_28501,N_29268);
nor U30583 (N_30583,N_25530,N_25455);
nand U30584 (N_30584,N_25619,N_29761);
nor U30585 (N_30585,N_26431,N_26698);
and U30586 (N_30586,N_26916,N_28119);
xor U30587 (N_30587,N_28099,N_25628);
nand U30588 (N_30588,N_26114,N_29078);
and U30589 (N_30589,N_27285,N_25639);
nand U30590 (N_30590,N_28693,N_25365);
and U30591 (N_30591,N_25674,N_27732);
and U30592 (N_30592,N_29016,N_25659);
and U30593 (N_30593,N_26159,N_27205);
xnor U30594 (N_30594,N_28861,N_29365);
and U30595 (N_30595,N_29040,N_28327);
and U30596 (N_30596,N_25459,N_29149);
nand U30597 (N_30597,N_26038,N_25301);
nor U30598 (N_30598,N_28133,N_28108);
xor U30599 (N_30599,N_29367,N_25701);
xor U30600 (N_30600,N_25620,N_28703);
and U30601 (N_30601,N_27366,N_25333);
and U30602 (N_30602,N_25696,N_28556);
nor U30603 (N_30603,N_25408,N_26402);
and U30604 (N_30604,N_26198,N_27403);
nor U30605 (N_30605,N_27423,N_27665);
or U30606 (N_30606,N_29389,N_27666);
nor U30607 (N_30607,N_29312,N_26582);
or U30608 (N_30608,N_27867,N_26262);
nor U30609 (N_30609,N_27978,N_26529);
or U30610 (N_30610,N_26606,N_28455);
nor U30611 (N_30611,N_25036,N_28886);
nor U30612 (N_30612,N_25953,N_26863);
or U30613 (N_30613,N_26467,N_26860);
or U30614 (N_30614,N_26814,N_27272);
xor U30615 (N_30615,N_26648,N_29685);
nand U30616 (N_30616,N_25329,N_28177);
or U30617 (N_30617,N_25191,N_27367);
nand U30618 (N_30618,N_25385,N_25084);
and U30619 (N_30619,N_27513,N_26341);
or U30620 (N_30620,N_28781,N_28960);
nand U30621 (N_30621,N_28834,N_27157);
and U30622 (N_30622,N_25371,N_29841);
nor U30623 (N_30623,N_28476,N_26602);
xor U30624 (N_30624,N_26626,N_26135);
and U30625 (N_30625,N_28241,N_28293);
xnor U30626 (N_30626,N_29908,N_29432);
nand U30627 (N_30627,N_25500,N_29416);
or U30628 (N_30628,N_27352,N_27672);
nand U30629 (N_30629,N_26319,N_28326);
or U30630 (N_30630,N_25605,N_28175);
or U30631 (N_30631,N_27603,N_28353);
nand U30632 (N_30632,N_25099,N_26290);
and U30633 (N_30633,N_26583,N_26846);
or U30634 (N_30634,N_25139,N_27550);
xnor U30635 (N_30635,N_25164,N_27073);
xor U30636 (N_30636,N_28600,N_28482);
and U30637 (N_30637,N_25558,N_26540);
nand U30638 (N_30638,N_28711,N_29792);
or U30639 (N_30639,N_29027,N_26178);
nand U30640 (N_30640,N_28920,N_27696);
or U30641 (N_30641,N_27449,N_25496);
nor U30642 (N_30642,N_27436,N_28871);
nor U30643 (N_30643,N_26232,N_29566);
nand U30644 (N_30644,N_27462,N_28535);
nand U30645 (N_30645,N_28206,N_27815);
nor U30646 (N_30646,N_29741,N_29948);
nand U30647 (N_30647,N_26958,N_25983);
and U30648 (N_30648,N_28673,N_25372);
or U30649 (N_30649,N_25388,N_26256);
nand U30650 (N_30650,N_29873,N_27349);
nand U30651 (N_30651,N_26398,N_28059);
and U30652 (N_30652,N_25421,N_29435);
nand U30653 (N_30653,N_29975,N_29503);
or U30654 (N_30654,N_26456,N_27891);
nor U30655 (N_30655,N_25259,N_27645);
and U30656 (N_30656,N_27544,N_25785);
or U30657 (N_30657,N_27528,N_25370);
nor U30658 (N_30658,N_26862,N_28723);
nor U30659 (N_30659,N_25263,N_29791);
and U30660 (N_30660,N_29332,N_28363);
and U30661 (N_30661,N_28032,N_28653);
and U30662 (N_30662,N_26316,N_27615);
nand U30663 (N_30663,N_26991,N_26441);
nor U30664 (N_30664,N_26271,N_25816);
nand U30665 (N_30665,N_27246,N_29736);
or U30666 (N_30666,N_29226,N_29082);
nor U30667 (N_30667,N_29531,N_26395);
nand U30668 (N_30668,N_25988,N_27379);
nand U30669 (N_30669,N_29874,N_27356);
nor U30670 (N_30670,N_26574,N_26763);
xor U30671 (N_30671,N_29415,N_27066);
nand U30672 (N_30672,N_27001,N_29590);
nor U30673 (N_30673,N_28943,N_26680);
nor U30674 (N_30674,N_28159,N_26068);
and U30675 (N_30675,N_28271,N_29205);
or U30676 (N_30676,N_27278,N_28251);
and U30677 (N_30677,N_29722,N_27503);
and U30678 (N_30678,N_29222,N_28803);
and U30679 (N_30679,N_25905,N_25811);
nor U30680 (N_30680,N_26469,N_29060);
nor U30681 (N_30681,N_29734,N_29427);
or U30682 (N_30682,N_28899,N_28618);
xor U30683 (N_30683,N_29317,N_29157);
or U30684 (N_30684,N_28360,N_28751);
or U30685 (N_30685,N_25209,N_27552);
or U30686 (N_30686,N_26179,N_25192);
nand U30687 (N_30687,N_26225,N_26902);
and U30688 (N_30688,N_27268,N_25197);
nor U30689 (N_30689,N_26652,N_29670);
or U30690 (N_30690,N_25859,N_25759);
and U30691 (N_30691,N_26391,N_27447);
or U30692 (N_30692,N_28161,N_28801);
or U30693 (N_30693,N_26348,N_25960);
or U30694 (N_30694,N_25147,N_25907);
nor U30695 (N_30695,N_29913,N_25386);
or U30696 (N_30696,N_29446,N_26353);
nand U30697 (N_30697,N_26722,N_26740);
and U30698 (N_30698,N_26362,N_29804);
nand U30699 (N_30699,N_26202,N_25528);
xnor U30700 (N_30700,N_28732,N_29346);
xnor U30701 (N_30701,N_26637,N_25612);
nor U30702 (N_30702,N_26163,N_26742);
and U30703 (N_30703,N_25815,N_29510);
and U30704 (N_30704,N_28843,N_28193);
and U30705 (N_30705,N_27737,N_25119);
and U30706 (N_30706,N_27785,N_28093);
nor U30707 (N_30707,N_29024,N_25638);
xor U30708 (N_30708,N_25065,N_29049);
xor U30709 (N_30709,N_28471,N_26678);
nand U30710 (N_30710,N_26158,N_29833);
or U30711 (N_30711,N_25449,N_25969);
nand U30712 (N_30712,N_28258,N_25691);
xor U30713 (N_30713,N_25029,N_28684);
and U30714 (N_30714,N_27258,N_27599);
and U30715 (N_30715,N_26473,N_26510);
nor U30716 (N_30716,N_28089,N_28079);
nor U30717 (N_30717,N_29141,N_29978);
and U30718 (N_30718,N_25970,N_29994);
nand U30719 (N_30719,N_29778,N_27213);
or U30720 (N_30720,N_28696,N_28019);
and U30721 (N_30721,N_27120,N_25703);
nor U30722 (N_30722,N_25405,N_28688);
xnor U30723 (N_30723,N_26522,N_27897);
nand U30724 (N_30724,N_25462,N_29246);
and U30725 (N_30725,N_27752,N_29200);
and U30726 (N_30726,N_26816,N_28220);
xor U30727 (N_30727,N_29248,N_26819);
nor U30728 (N_30728,N_29805,N_29309);
or U30729 (N_30729,N_28235,N_29536);
and U30730 (N_30730,N_28743,N_26072);
and U30731 (N_30731,N_29108,N_25743);
nor U30732 (N_30732,N_26289,N_26615);
nand U30733 (N_30733,N_29233,N_25202);
nor U30734 (N_30734,N_26931,N_28230);
xor U30735 (N_30735,N_27547,N_25246);
nand U30736 (N_30736,N_26773,N_28627);
or U30737 (N_30737,N_27775,N_25993);
nor U30738 (N_30738,N_28383,N_25198);
and U30739 (N_30739,N_28346,N_25834);
or U30740 (N_30740,N_25776,N_27390);
nand U30741 (N_30741,N_26910,N_27455);
or U30742 (N_30742,N_26543,N_27784);
xnor U30743 (N_30743,N_29371,N_26372);
nor U30744 (N_30744,N_25397,N_28538);
or U30745 (N_30745,N_29962,N_28160);
and U30746 (N_30746,N_27241,N_29011);
nor U30747 (N_30747,N_28666,N_29940);
and U30748 (N_30748,N_25593,N_25120);
and U30749 (N_30749,N_25554,N_29120);
or U30750 (N_30750,N_28409,N_27953);
nor U30751 (N_30751,N_28184,N_26086);
or U30752 (N_30752,N_26494,N_29825);
nor U30753 (N_30753,N_25316,N_26674);
xor U30754 (N_30754,N_29378,N_26328);
xnor U30755 (N_30755,N_28172,N_29164);
nor U30756 (N_30756,N_29853,N_26715);
and U30757 (N_30757,N_27185,N_29071);
nand U30758 (N_30758,N_26307,N_26841);
and U30759 (N_30759,N_26794,N_28247);
nand U30760 (N_30760,N_25308,N_29144);
or U30761 (N_30761,N_29753,N_27110);
nand U30762 (N_30762,N_27104,N_28497);
xnor U30763 (N_30763,N_28551,N_26008);
and U30764 (N_30764,N_25472,N_28798);
and U30765 (N_30765,N_29512,N_29550);
nand U30766 (N_30766,N_26127,N_29716);
or U30767 (N_30767,N_28547,N_27727);
or U30768 (N_30768,N_26825,N_27491);
and U30769 (N_30769,N_25527,N_28860);
nand U30770 (N_30770,N_28047,N_28961);
nor U30771 (N_30771,N_25145,N_27590);
nand U30772 (N_30772,N_29316,N_27854);
xor U30773 (N_30773,N_25542,N_27089);
nand U30774 (N_30774,N_29211,N_26857);
nand U30775 (N_30775,N_27626,N_28827);
or U30776 (N_30776,N_25347,N_27657);
nor U30777 (N_30777,N_25895,N_27810);
or U30778 (N_30778,N_25798,N_26420);
nor U30779 (N_30779,N_27939,N_25465);
and U30780 (N_30780,N_25597,N_26261);
nand U30781 (N_30781,N_26284,N_29393);
and U30782 (N_30782,N_26356,N_29218);
and U30783 (N_30783,N_25131,N_29296);
or U30784 (N_30784,N_25028,N_25155);
or U30785 (N_30785,N_26333,N_27437);
nand U30786 (N_30786,N_28942,N_28082);
nor U30787 (N_30787,N_27186,N_28955);
and U30788 (N_30788,N_27482,N_29235);
or U30789 (N_30789,N_25063,N_25959);
nand U30790 (N_30790,N_27859,N_26805);
and U30791 (N_30791,N_28818,N_28984);
nor U30792 (N_30792,N_28495,N_28048);
nor U30793 (N_30793,N_27019,N_29905);
nor U30794 (N_30794,N_28588,N_28667);
or U30795 (N_30795,N_26076,N_27315);
or U30796 (N_30796,N_28664,N_27263);
xor U30797 (N_30797,N_28833,N_26516);
nor U30798 (N_30798,N_27783,N_29183);
xnor U30799 (N_30799,N_26097,N_27803);
xor U30800 (N_30800,N_28380,N_27275);
and U30801 (N_30801,N_25448,N_26760);
nand U30802 (N_30802,N_28561,N_26984);
nand U30803 (N_30803,N_29072,N_27652);
and U30804 (N_30804,N_27211,N_28847);
nand U30805 (N_30805,N_26160,N_26887);
and U30806 (N_30806,N_28555,N_26053);
nand U30807 (N_30807,N_29801,N_29872);
nand U30808 (N_30808,N_28977,N_26727);
nor U30809 (N_30809,N_26669,N_26558);
nor U30810 (N_30810,N_27145,N_25794);
or U30811 (N_30811,N_29154,N_27517);
and U30812 (N_30812,N_28617,N_25668);
nand U30813 (N_30813,N_25915,N_26457);
and U30814 (N_30814,N_26141,N_25189);
nand U30815 (N_30815,N_25276,N_25275);
xnor U30816 (N_30816,N_29644,N_28736);
xnor U30817 (N_30817,N_27500,N_27726);
xnor U30818 (N_30818,N_29179,N_29572);
xnor U30819 (N_30819,N_26073,N_29564);
nand U30820 (N_30820,N_28876,N_28037);
nand U30821 (N_30821,N_29630,N_28337);
nand U30822 (N_30822,N_25261,N_27755);
nor U30823 (N_30823,N_27284,N_29507);
or U30824 (N_30824,N_28993,N_25003);
nor U30825 (N_30825,N_25609,N_26917);
or U30826 (N_30826,N_27302,N_27974);
or U30827 (N_30827,N_28490,N_25172);
nand U30828 (N_30828,N_28289,N_26535);
nor U30829 (N_30829,N_27681,N_27282);
or U30830 (N_30830,N_26115,N_26869);
or U30831 (N_30831,N_26547,N_25820);
or U30832 (N_30832,N_28670,N_29505);
and U30833 (N_30833,N_29151,N_25006);
or U30834 (N_30834,N_28468,N_28802);
nor U30835 (N_30835,N_29110,N_27881);
nor U30836 (N_30836,N_29100,N_26809);
nor U30837 (N_30837,N_29965,N_26339);
and U30838 (N_30838,N_25379,N_28900);
xor U30839 (N_30839,N_28115,N_25199);
nand U30840 (N_30840,N_28266,N_29808);
nand U30841 (N_30841,N_27570,N_28145);
or U30842 (N_30842,N_25780,N_27816);
nor U30843 (N_30843,N_25071,N_28506);
nor U30844 (N_30844,N_25007,N_26614);
and U30845 (N_30845,N_25505,N_28411);
or U30846 (N_30846,N_25572,N_27005);
nand U30847 (N_30847,N_28321,N_25396);
or U30848 (N_30848,N_27194,N_26349);
and U30849 (N_30849,N_25821,N_28020);
or U30850 (N_30850,N_25249,N_25247);
nor U30851 (N_30851,N_28722,N_25932);
nor U30852 (N_30852,N_25765,N_28742);
nand U30853 (N_30853,N_29961,N_27773);
or U30854 (N_30854,N_28231,N_27571);
nand U30855 (N_30855,N_25867,N_27305);
nand U30856 (N_30856,N_28770,N_28850);
and U30857 (N_30857,N_25171,N_25035);
and U30858 (N_30858,N_25416,N_25291);
nor U30859 (N_30859,N_27988,N_28460);
nand U30860 (N_30860,N_27538,N_26640);
nor U30861 (N_30861,N_28408,N_25577);
and U30862 (N_30862,N_25863,N_29320);
and U30863 (N_30863,N_27840,N_28188);
nor U30864 (N_30864,N_27797,N_25862);
or U30865 (N_30865,N_29357,N_29569);
nor U30866 (N_30866,N_28884,N_29006);
nand U30867 (N_30867,N_29029,N_26383);
nor U30868 (N_30868,N_27402,N_25080);
or U30869 (N_30869,N_28147,N_27796);
nor U30870 (N_30870,N_27124,N_28660);
nand U30871 (N_30871,N_29053,N_29661);
nand U30872 (N_30872,N_25179,N_26425);
nor U30873 (N_30873,N_25163,N_28741);
nor U30874 (N_30874,N_27103,N_27804);
and U30875 (N_30875,N_25667,N_29044);
nand U30876 (N_30876,N_29349,N_27378);
nor U30877 (N_30877,N_26884,N_28171);
xnor U30878 (N_30878,N_29839,N_27016);
nor U30879 (N_30879,N_25351,N_25977);
and U30880 (N_30880,N_26899,N_27753);
or U30881 (N_30881,N_29735,N_26612);
or U30882 (N_30882,N_27221,N_28128);
and U30883 (N_30883,N_26165,N_29469);
nor U30884 (N_30884,N_27983,N_27062);
nand U30885 (N_30885,N_29061,N_28444);
or U30886 (N_30886,N_25042,N_26002);
nand U30887 (N_30887,N_29915,N_25141);
nand U30888 (N_30888,N_28433,N_26218);
nand U30889 (N_30889,N_26313,N_25399);
nand U30890 (N_30890,N_27428,N_26478);
nor U30891 (N_30891,N_27365,N_26981);
or U30892 (N_30892,N_29673,N_25419);
nand U30893 (N_30893,N_29964,N_27540);
nor U30894 (N_30894,N_29259,N_28557);
nand U30895 (N_30895,N_27351,N_25319);
or U30896 (N_30896,N_25720,N_26595);
nor U30897 (N_30897,N_29348,N_27762);
or U30898 (N_30898,N_25343,N_25030);
and U30899 (N_30899,N_26527,N_25526);
and U30900 (N_30900,N_27269,N_27014);
or U30901 (N_30901,N_25492,N_29294);
or U30902 (N_30902,N_27924,N_27685);
and U30903 (N_30903,N_26308,N_27551);
and U30904 (N_30904,N_25561,N_28462);
and U30905 (N_30905,N_25885,N_28448);
xor U30906 (N_30906,N_26721,N_29720);
nand U30907 (N_30907,N_29711,N_26447);
or U30908 (N_30908,N_25516,N_28313);
or U30909 (N_30909,N_25451,N_29786);
or U30910 (N_30910,N_29398,N_29288);
nand U30911 (N_30911,N_28488,N_28064);
or U30912 (N_30912,N_29751,N_28968);
xnor U30913 (N_30913,N_27160,N_27121);
or U30914 (N_30914,N_25285,N_26550);
or U30915 (N_30915,N_25067,N_28242);
nor U30916 (N_30916,N_29172,N_26025);
nor U30917 (N_30917,N_28549,N_25642);
xnor U30918 (N_30918,N_28882,N_29377);
or U30919 (N_30919,N_25330,N_28721);
nand U30920 (N_30920,N_26242,N_27249);
nor U30921 (N_30921,N_25944,N_29887);
nor U30922 (N_30922,N_27999,N_25999);
or U30923 (N_30923,N_25723,N_27372);
and U30924 (N_30924,N_28759,N_27630);
nor U30925 (N_30925,N_26470,N_25116);
nand U30926 (N_30926,N_26274,N_29359);
and U30927 (N_30927,N_26684,N_29476);
or U30928 (N_30928,N_26345,N_26681);
and U30929 (N_30929,N_29282,N_27262);
and U30930 (N_30930,N_26897,N_28357);
nand U30931 (N_30931,N_29800,N_27184);
nand U30932 (N_30932,N_25016,N_26015);
or U30933 (N_30933,N_27695,N_25107);
or U30934 (N_30934,N_27522,N_27454);
xnor U30935 (N_30935,N_26789,N_27812);
and U30936 (N_30936,N_26734,N_27667);
nand U30937 (N_30937,N_28735,N_27805);
xnor U30938 (N_30938,N_27865,N_25018);
nor U30939 (N_30939,N_25692,N_28951);
or U30940 (N_30940,N_25504,N_26408);
nor U30941 (N_30941,N_27286,N_26087);
nand U30942 (N_30942,N_29855,N_28051);
and U30943 (N_30943,N_26009,N_29344);
nand U30944 (N_30944,N_27175,N_29747);
or U30945 (N_30945,N_29134,N_28028);
nor U30946 (N_30946,N_28078,N_28067);
and U30947 (N_30947,N_26233,N_26309);
and U30948 (N_30948,N_28507,N_26452);
nand U30949 (N_30949,N_25951,N_29857);
nor U30950 (N_30950,N_27414,N_25607);
nand U30951 (N_30951,N_28842,N_29448);
and U30952 (N_30952,N_27152,N_26628);
or U30953 (N_30953,N_28745,N_29345);
xor U30954 (N_30954,N_25341,N_29776);
nand U30955 (N_30955,N_28487,N_27774);
nand U30956 (N_30956,N_27957,N_26744);
or U30957 (N_30957,N_25541,N_25010);
nor U30958 (N_30958,N_29538,N_25644);
xnor U30959 (N_30959,N_26781,N_25987);
nor U30960 (N_30960,N_25717,N_27395);
and U30961 (N_30961,N_29052,N_27613);
nor U30962 (N_30962,N_27134,N_28576);
nand U30963 (N_30963,N_26590,N_27508);
nor U30964 (N_30964,N_29467,N_29878);
nor U30965 (N_30965,N_27170,N_29250);
nor U30966 (N_30966,N_27948,N_26321);
nand U30967 (N_30967,N_26948,N_25431);
nor U30968 (N_30968,N_25760,N_29462);
or U30969 (N_30969,N_28432,N_26273);
and U30970 (N_30970,N_28934,N_29188);
and U30971 (N_30971,N_27648,N_28494);
nand U30972 (N_30972,N_28838,N_28778);
nand U30973 (N_30973,N_29972,N_26866);
nor U30974 (N_30974,N_25488,N_29969);
nand U30975 (N_30975,N_28848,N_28651);
xor U30976 (N_30976,N_28725,N_29859);
or U30977 (N_30977,N_29957,N_28677);
nand U30978 (N_30978,N_27292,N_26324);
nand U30979 (N_30979,N_27620,N_26661);
nor U30980 (N_30980,N_27086,N_29184);
nor U30981 (N_30981,N_26625,N_26155);
nor U30982 (N_30982,N_25248,N_29546);
or U30983 (N_30983,N_26245,N_26320);
nand U30984 (N_30984,N_25604,N_26136);
nand U30985 (N_30985,N_25078,N_27634);
nand U30986 (N_30986,N_25355,N_26914);
and U30987 (N_30987,N_28933,N_28662);
nand U30988 (N_30988,N_25536,N_27582);
nand U30989 (N_30989,N_29022,N_26850);
or U30990 (N_30990,N_29516,N_27063);
nor U30991 (N_30991,N_29816,N_27900);
nand U30992 (N_30992,N_27577,N_27919);
or U30993 (N_30993,N_29680,N_27884);
and U30994 (N_30994,N_29382,N_27208);
nand U30995 (N_30995,N_26022,N_26591);
nor U30996 (N_30996,N_27373,N_25470);
or U30997 (N_30997,N_25581,N_26000);
or U30998 (N_30998,N_26913,N_28489);
nor U30999 (N_30999,N_28385,N_25699);
or U31000 (N_31000,N_25509,N_29498);
or U31001 (N_31001,N_25376,N_28430);
or U31002 (N_31002,N_25595,N_28626);
or U31003 (N_31003,N_25230,N_29480);
or U31004 (N_31004,N_28045,N_28349);
nor U31005 (N_31005,N_25737,N_28347);
nand U31006 (N_31006,N_26430,N_28233);
or U31007 (N_31007,N_29287,N_27818);
and U31008 (N_31008,N_27977,N_29770);
or U31009 (N_31009,N_26458,N_29681);
nand U31010 (N_31010,N_26468,N_25799);
nand U31011 (N_31011,N_27664,N_29933);
nor U31012 (N_31012,N_28405,N_26621);
and U31013 (N_31013,N_29500,N_27894);
and U31014 (N_31014,N_25038,N_28916);
and U31015 (N_31015,N_26503,N_28415);
nor U31016 (N_31016,N_26511,N_25758);
nand U31017 (N_31017,N_25013,N_27460);
or U31018 (N_31018,N_27870,N_29790);
nor U31019 (N_31019,N_26762,N_27833);
or U31020 (N_31020,N_26788,N_26092);
or U31021 (N_31021,N_29684,N_26246);
nand U31022 (N_31022,N_27069,N_27703);
nor U31023 (N_31023,N_27934,N_29850);
and U31024 (N_31024,N_26717,N_28953);
nand U31025 (N_31025,N_26922,N_27710);
nor U31026 (N_31026,N_25825,N_25693);
and U31027 (N_31027,N_29105,N_25060);
xnor U31028 (N_31028,N_27594,N_28982);
nor U31029 (N_31029,N_29264,N_25425);
nor U31030 (N_31030,N_29879,N_27296);
or U31031 (N_31031,N_25053,N_28524);
and U31032 (N_31032,N_29653,N_27381);
and U31033 (N_31033,N_26048,N_28480);
and U31034 (N_31034,N_26886,N_27966);
nand U31035 (N_31035,N_25325,N_26517);
nand U31036 (N_31036,N_29665,N_29656);
nor U31037 (N_31037,N_27426,N_25336);
and U31038 (N_31038,N_25413,N_28964);
or U31039 (N_31039,N_28714,N_28792);
or U31040 (N_31040,N_27451,N_29989);
nand U31041 (N_31041,N_25778,N_28631);
nor U31042 (N_31042,N_28227,N_26579);
nor U31043 (N_31043,N_26103,N_25331);
xor U31044 (N_31044,N_25774,N_26990);
and U31045 (N_31045,N_28006,N_28111);
or U31046 (N_31046,N_26459,N_29595);
nor U31047 (N_31047,N_26638,N_29239);
or U31048 (N_31048,N_29709,N_26536);
or U31049 (N_31049,N_26664,N_26803);
nor U31050 (N_31050,N_26584,N_29612);
nand U31051 (N_31051,N_25384,N_27290);
or U31052 (N_31052,N_29894,N_29543);
or U31053 (N_31053,N_26515,N_29604);
and U31054 (N_31054,N_27393,N_25091);
or U31055 (N_31055,N_27487,N_28376);
nand U31056 (N_31056,N_25921,N_26485);
and U31057 (N_31057,N_26926,N_29635);
xnor U31058 (N_31058,N_27328,N_25320);
or U31059 (N_31059,N_25318,N_29624);
nor U31060 (N_31060,N_27360,N_25299);
or U31061 (N_31061,N_29561,N_28813);
or U31062 (N_31062,N_27340,N_26336);
nor U31063 (N_31063,N_29748,N_28180);
nand U31064 (N_31064,N_27181,N_27293);
nand U31065 (N_31065,N_25482,N_29310);
xnor U31066 (N_31066,N_28131,N_28149);
nor U31067 (N_31067,N_27892,N_26331);
and U31068 (N_31068,N_27313,N_27962);
or U31069 (N_31069,N_27441,N_27336);
nand U31070 (N_31070,N_28367,N_29215);
or U31071 (N_31071,N_27898,N_29486);
nor U31072 (N_31072,N_27440,N_26545);
and U31073 (N_31073,N_26955,N_28533);
or U31074 (N_31074,N_27642,N_27534);
nor U31075 (N_31075,N_26643,N_28978);
or U31076 (N_31076,N_25751,N_29647);
nand U31077 (N_31077,N_28649,N_29077);
or U31078 (N_31078,N_27826,N_27253);
and U31079 (N_31079,N_26286,N_25738);
nand U31080 (N_31080,N_25590,N_29379);
and U31081 (N_31081,N_29603,N_29682);
nor U31082 (N_31082,N_28522,N_28755);
nand U31083 (N_31083,N_29434,N_29780);
nand U31084 (N_31084,N_27926,N_27986);
or U31085 (N_31085,N_29499,N_29224);
nand U31086 (N_31086,N_27470,N_29717);
nor U31087 (N_31087,N_29124,N_25998);
nor U31088 (N_31088,N_29568,N_28921);
xor U31089 (N_31089,N_25772,N_26979);
xor U31090 (N_31090,N_26822,N_29755);
nand U31091 (N_31091,N_26769,N_29606);
nor U31092 (N_31092,N_29442,N_28129);
nand U31093 (N_31093,N_29364,N_26170);
nor U31094 (N_31094,N_25487,N_26785);
xnor U31095 (N_31095,N_25241,N_26706);
xnor U31096 (N_31096,N_29085,N_28769);
and U31097 (N_31097,N_28573,N_25766);
nor U31098 (N_31098,N_26384,N_29209);
nand U31099 (N_31099,N_29391,N_28910);
and U31100 (N_31100,N_29162,N_25556);
nor U31101 (N_31101,N_26479,N_26812);
nor U31102 (N_31102,N_26712,N_27618);
or U31103 (N_31103,N_27099,N_26123);
and U31104 (N_31104,N_29982,N_25380);
xnor U31105 (N_31105,N_26546,N_27332);
nor U31106 (N_31106,N_28127,N_26764);
nor U31107 (N_31107,N_28384,N_26532);
or U31108 (N_31108,N_25450,N_29116);
nand U31109 (N_31109,N_27021,N_29249);
and U31110 (N_31110,N_26477,N_26074);
nor U31111 (N_31111,N_27743,N_26191);
xnor U31112 (N_31112,N_29256,N_29576);
or U31113 (N_31113,N_27051,N_28341);
or U31114 (N_31114,N_29737,N_27361);
and U31115 (N_31115,N_28377,N_26966);
or U31116 (N_31116,N_27592,N_29396);
and U31117 (N_31117,N_25657,N_28612);
nand U31118 (N_31118,N_25610,N_26969);
nor U31119 (N_31119,N_25744,N_25321);
nor U31120 (N_31120,N_28190,N_29386);
xnor U31121 (N_31121,N_27578,N_26653);
xor U31122 (N_31122,N_27038,N_27031);
nor U31123 (N_31123,N_27750,N_29266);
and U31124 (N_31124,N_27843,N_27188);
and U31125 (N_31125,N_27404,N_25095);
or U31126 (N_31126,N_29362,N_25982);
or U31127 (N_31127,N_28017,N_28062);
or U31128 (N_31128,N_26301,N_25309);
xnor U31129 (N_31129,N_29429,N_28892);
or U31130 (N_31130,N_28614,N_29712);
or U31131 (N_31131,N_28074,N_28101);
nand U31132 (N_31132,N_26757,N_26538);
nand U31133 (N_31133,N_29643,N_26623);
nand U31134 (N_31134,N_26702,N_27739);
nand U31135 (N_31135,N_25830,N_29490);
or U31136 (N_31136,N_28971,N_28272);
and U31137 (N_31137,N_26294,N_29752);
or U31138 (N_31138,N_29840,N_26387);
and U31139 (N_31139,N_25981,N_29995);
nand U31140 (N_31140,N_27746,N_28336);
nand U31141 (N_31141,N_28508,N_29594);
nand U31142 (N_31142,N_27096,N_26856);
or U31143 (N_31143,N_27705,N_26282);
nand U31144 (N_31144,N_26849,N_26060);
nand U31145 (N_31145,N_25280,N_25477);
nand U31146 (N_31146,N_27331,N_25979);
or U31147 (N_31147,N_26119,N_29413);
or U31148 (N_31148,N_28138,N_27164);
nand U31149 (N_31149,N_29271,N_27010);
and U31150 (N_31150,N_26976,N_25440);
nor U31151 (N_31151,N_27028,N_28255);
nor U31152 (N_31152,N_29578,N_27078);
or U31153 (N_31153,N_27254,N_27712);
or U31154 (N_31154,N_29725,N_29582);
and U31155 (N_31155,N_28427,N_26932);
and U31156 (N_31156,N_26796,N_27913);
nand U31157 (N_31157,N_25508,N_29749);
and U31158 (N_31158,N_29812,N_27496);
nand U31159 (N_31159,N_25802,N_25032);
nand U31160 (N_31160,N_27987,N_25942);
and U31161 (N_31161,N_29936,N_25908);
xor U31162 (N_31162,N_29542,N_26203);
and U31163 (N_31163,N_25273,N_28913);
or U31164 (N_31164,N_29575,N_29508);
and U31165 (N_31165,N_28550,N_28492);
and U31166 (N_31166,N_26162,N_26746);
nand U31167 (N_31167,N_29861,N_29579);
and U31168 (N_31168,N_29909,N_25857);
and U31169 (N_31169,N_26064,N_26502);
nand U31170 (N_31170,N_27304,N_27817);
nor U31171 (N_31171,N_27825,N_28071);
and U31172 (N_31172,N_29689,N_29892);
nor U31173 (N_31173,N_29733,N_25094);
or U31174 (N_31174,N_29671,N_28084);
or U31175 (N_31175,N_29037,N_26929);
and U31176 (N_31176,N_25326,N_28369);
or U31177 (N_31177,N_25791,N_29180);
nand U31178 (N_31178,N_29076,N_25436);
and U31179 (N_31179,N_29560,N_28765);
and U31180 (N_31180,N_29420,N_26297);
nand U31181 (N_31181,N_25829,N_26514);
and U31182 (N_31182,N_28157,N_29445);
and U31183 (N_31183,N_26605,N_29820);
nor U31184 (N_31184,N_25838,N_27714);
nor U31185 (N_31185,N_26166,N_25494);
nand U31186 (N_31186,N_27533,N_26534);
nor U31187 (N_31187,N_28806,N_27744);
nor U31188 (N_31188,N_26891,N_25817);
or U31189 (N_31189,N_27143,N_29103);
or U31190 (N_31190,N_29101,N_28396);
or U31191 (N_31191,N_25187,N_27106);
and U31192 (N_31192,N_25688,N_26654);
or U31193 (N_31193,N_28450,N_25284);
or U31194 (N_31194,N_27112,N_29704);
nor U31195 (N_31195,N_28584,N_27024);
and U31196 (N_31196,N_26889,N_29705);
or U31197 (N_31197,N_28458,N_29463);
or U31198 (N_31198,N_29672,N_26888);
xnor U31199 (N_31199,N_25479,N_27593);
nor U31200 (N_31200,N_25858,N_27972);
and U31201 (N_31201,N_26026,N_25484);
xnor U31202 (N_31202,N_26905,N_26898);
xor U31203 (N_31203,N_29338,N_28397);
nand U31204 (N_31204,N_26709,N_29148);
nor U31205 (N_31205,N_28094,N_26551);
and U31206 (N_31206,N_29980,N_26361);
nor U31207 (N_31207,N_29496,N_29867);
nand U31208 (N_31208,N_29732,N_28753);
or U31209 (N_31209,N_28308,N_27389);
or U31210 (N_31210,N_25417,N_29721);
nand U31211 (N_31211,N_27828,N_25422);
xnor U31212 (N_31212,N_27601,N_28121);
nand U31213 (N_31213,N_28484,N_26172);
or U31214 (N_31214,N_29113,N_25464);
and U31215 (N_31215,N_26084,N_27071);
nor U31216 (N_31216,N_29766,N_28358);
and U31217 (N_31217,N_29611,N_28300);
nand U31218 (N_31218,N_26520,N_27026);
and U31219 (N_31219,N_29864,N_28795);
or U31220 (N_31220,N_26251,N_25735);
or U31221 (N_31221,N_27217,N_28477);
nor U31222 (N_31222,N_26445,N_29863);
nand U31223 (N_31223,N_29935,N_27497);
nor U31224 (N_31224,N_27435,N_25645);
nand U31225 (N_31225,N_27416,N_27037);
nor U31226 (N_31226,N_28852,N_25756);
nand U31227 (N_31227,N_28486,N_29891);
nor U31228 (N_31228,N_29993,N_25050);
or U31229 (N_31229,N_27050,N_28859);
nand U31230 (N_31230,N_25883,N_26820);
or U31231 (N_31231,N_28275,N_27515);
and U31232 (N_31232,N_29533,N_29703);
and U31233 (N_31233,N_25220,N_29358);
nand U31234 (N_31234,N_28050,N_25226);
and U31235 (N_31235,N_27301,N_28782);
nor U31236 (N_31236,N_29007,N_26471);
nor U31237 (N_31237,N_27708,N_25143);
nand U31238 (N_31238,N_26330,N_25194);
nor U31239 (N_31239,N_28583,N_26055);
or U31240 (N_31240,N_25457,N_29221);
nand U31241 (N_31241,N_25491,N_26375);
nor U31242 (N_31242,N_25650,N_26455);
xor U31243 (N_31243,N_29122,N_26118);
nand U31244 (N_31244,N_29807,N_29627);
nor U31245 (N_31245,N_29208,N_29323);
nor U31246 (N_31246,N_29241,N_25713);
or U31247 (N_31247,N_26426,N_29293);
nand U31248 (N_31248,N_25836,N_28897);
and U31249 (N_31249,N_26561,N_25678);
nand U31250 (N_31250,N_29666,N_25978);
or U31251 (N_31251,N_26635,N_29321);
nand U31252 (N_31252,N_25608,N_25458);
nor U31253 (N_31253,N_27406,N_28790);
or U31254 (N_31254,N_27745,N_27780);
and U31255 (N_31255,N_28307,N_26252);
xnor U31256 (N_31256,N_29114,N_28077);
xor U31257 (N_31257,N_26506,N_25020);
and U31258 (N_31258,N_27858,N_28846);
nor U31259 (N_31259,N_29097,N_25296);
or U31260 (N_31260,N_28209,N_29193);
nor U31261 (N_31261,N_28862,N_26049);
nor U31262 (N_31262,N_28820,N_28707);
or U31263 (N_31263,N_28689,N_27631);
nand U31264 (N_31264,N_26720,N_28936);
or U31265 (N_31265,N_27196,N_26090);
nand U31266 (N_31266,N_28650,N_25706);
xor U31267 (N_31267,N_27761,N_28203);
or U31268 (N_31268,N_28687,N_26730);
and U31269 (N_31269,N_29570,N_29950);
and U31270 (N_31270,N_29553,N_26688);
and U31271 (N_31271,N_25203,N_26393);
nor U31272 (N_31272,N_29667,N_28314);
nor U31273 (N_31273,N_29263,N_29871);
nand U31274 (N_31274,N_29845,N_27624);
or U31275 (N_31275,N_28625,N_26451);
or U31276 (N_31276,N_26580,N_28438);
nor U31277 (N_31277,N_28558,N_28539);
xor U31278 (N_31278,N_26967,N_27431);
and U31279 (N_31279,N_29404,N_27370);
or U31280 (N_31280,N_26409,N_28739);
nand U31281 (N_31281,N_26791,N_28824);
xor U31282 (N_31282,N_25812,N_27276);
or U31283 (N_31283,N_28057,N_28783);
nand U31284 (N_31284,N_29137,N_27486);
nor U31285 (N_31285,N_26751,N_29953);
xor U31286 (N_31286,N_29600,N_27113);
nand U31287 (N_31287,N_25424,N_25827);
nand U31288 (N_31288,N_26075,N_26429);
or U31289 (N_31289,N_28452,N_29771);
nor U31290 (N_31290,N_26110,N_25839);
or U31291 (N_31291,N_28372,N_27409);
nand U31292 (N_31292,N_28656,N_27488);
nand U31293 (N_31293,N_27605,N_27772);
nor U31294 (N_31294,N_27738,N_26474);
or U31295 (N_31295,N_27699,N_25594);
or U31296 (N_31296,N_27362,N_29625);
nand U31297 (N_31297,N_27612,N_25034);
or U31298 (N_31298,N_28530,N_29754);
nand U31299 (N_31299,N_29185,N_27330);
or U31300 (N_31300,N_27956,N_26318);
or U31301 (N_31301,N_29189,N_25562);
nor U31302 (N_31302,N_25069,N_26939);
nand U31303 (N_31303,N_26388,N_28873);
nand U31304 (N_31304,N_27338,N_25871);
and U31305 (N_31305,N_25764,N_28652);
xor U31306 (N_31306,N_29285,N_28389);
nand U31307 (N_31307,N_25739,N_28659);
nor U31308 (N_31308,N_26146,N_26659);
nand U31309 (N_31309,N_25138,N_26834);
or U31310 (N_31310,N_26666,N_25303);
nor U31311 (N_31311,N_26268,N_27869);
nor U31312 (N_31312,N_29194,N_27790);
xor U31313 (N_31313,N_27067,N_28553);
nand U31314 (N_31314,N_28985,N_27159);
nor U31315 (N_31315,N_28205,N_26187);
nor U31316 (N_31316,N_27850,N_27961);
and U31317 (N_31317,N_27531,N_25622);
xnor U31318 (N_31318,N_29774,N_27132);
xnor U31319 (N_31319,N_26258,N_26106);
nand U31320 (N_31320,N_29203,N_27093);
and U31321 (N_31321,N_27507,N_27718);
nor U31322 (N_31322,N_26463,N_25962);
nand U31323 (N_31323,N_26254,N_26182);
nor U31324 (N_31324,N_27461,N_27875);
and U31325 (N_31325,N_25896,N_26554);
nand U31326 (N_31326,N_25710,N_25502);
xnor U31327 (N_31327,N_26275,N_26209);
nor U31328 (N_31328,N_25891,N_29119);
nor U31329 (N_31329,N_29013,N_27786);
nand U31330 (N_31330,N_26620,N_28181);
xor U31331 (N_31331,N_28602,N_25415);
or U31332 (N_31332,N_28025,N_26901);
and U31333 (N_31333,N_28446,N_27166);
and U31334 (N_31334,N_27555,N_29779);
or U31335 (N_31335,N_28196,N_28597);
nor U31336 (N_31336,N_25251,N_27967);
and U31337 (N_31337,N_29176,N_29506);
nand U31338 (N_31338,N_26357,N_26619);
nand U31339 (N_31339,N_26953,N_26249);
or U31340 (N_31340,N_28370,N_27243);
or U31341 (N_31341,N_29232,N_27573);
and U31342 (N_31342,N_27214,N_25514);
and U31343 (N_31343,N_25864,N_26016);
nand U31344 (N_31344,N_28269,N_27938);
xor U31345 (N_31345,N_29888,N_27697);
and U31346 (N_31346,N_28013,N_29941);
nor U31347 (N_31347,N_26054,N_27009);
and U31348 (N_31348,N_28654,N_26521);
or U31349 (N_31349,N_29051,N_25501);
nor U31350 (N_31350,N_26642,N_26629);
nand U31351 (N_31351,N_26972,N_29252);
nand U31352 (N_31352,N_29893,N_29731);
nand U31353 (N_31353,N_26624,N_26696);
nand U31354 (N_31354,N_29088,N_26492);
nor U31355 (N_31355,N_27584,N_28807);
or U31356 (N_31356,N_27265,N_25524);
or U31357 (N_31357,N_25548,N_29534);
or U31358 (N_31358,N_25443,N_29902);
and U31359 (N_31359,N_28775,N_25073);
or U31360 (N_31360,N_29694,N_25680);
and U31361 (N_31361,N_29352,N_27008);
and U31362 (N_31362,N_26093,N_25796);
and U31363 (N_31363,N_26567,N_28908);
nand U31364 (N_31364,N_29327,N_26768);
nor U31365 (N_31365,N_26690,N_25290);
nand U31366 (N_31366,N_25613,N_29822);
or U31367 (N_31367,N_25009,N_26432);
nand U31368 (N_31368,N_27512,N_25503);
nor U31369 (N_31369,N_26587,N_25822);
and U31370 (N_31370,N_27151,N_25564);
nand U31371 (N_31371,N_29333,N_28959);
and U31372 (N_31372,N_27092,N_28104);
nand U31373 (N_31373,N_25306,N_25573);
or U31374 (N_31374,N_25389,N_26134);
and U31375 (N_31375,N_25850,N_28768);
nand U31376 (N_31376,N_27408,N_29046);
nor U31377 (N_31377,N_25840,N_27094);
nor U31378 (N_31378,N_28392,N_26444);
nor U31379 (N_31379,N_27498,N_28107);
nand U31380 (N_31380,N_27694,N_27871);
nand U31381 (N_31381,N_27100,N_25180);
or U31382 (N_31382,N_25846,N_25039);
xnor U31383 (N_31383,N_29527,N_26726);
and U31384 (N_31384,N_29216,N_25624);
or U31385 (N_31385,N_27219,N_25122);
nand U31386 (N_31386,N_26327,N_27116);
and U31387 (N_31387,N_27628,N_29657);
or U31388 (N_31388,N_25833,N_28459);
and U31389 (N_31389,N_25686,N_27133);
nand U31390 (N_31390,N_28158,N_27456);
nand U31391 (N_31391,N_26221,N_25041);
and U31392 (N_31392,N_26975,N_29487);
and U31393 (N_31393,N_28329,N_27432);
nor U31394 (N_31394,N_29311,N_28799);
and U31395 (N_31395,N_25398,N_26980);
nand U31396 (N_31396,N_29230,N_27324);
nor U31397 (N_31397,N_28958,N_25810);
and U31398 (N_31398,N_27140,N_26649);
nand U31399 (N_31399,N_28694,N_25152);
nand U31400 (N_31400,N_25714,N_25807);
nor U31401 (N_31401,N_25000,N_29436);
nor U31402 (N_31402,N_25563,N_29619);
or U31403 (N_31403,N_26782,N_29565);
nand U31404 (N_31404,N_29236,N_28150);
nor U31405 (N_31405,N_25755,N_27457);
nand U31406 (N_31406,N_29438,N_27206);
nand U31407 (N_31407,N_27357,N_26556);
nand U31408 (N_31408,N_27080,N_25363);
or U31409 (N_31409,N_28470,N_27354);
nand U31410 (N_31410,N_29471,N_28229);
and U31411 (N_31411,N_25088,N_27692);
or U31412 (N_31412,N_25109,N_28100);
and U31413 (N_31413,N_26033,N_27250);
nor U31414 (N_31414,N_28965,N_26544);
or U31415 (N_31415,N_28839,N_26462);
nor U31416 (N_31416,N_26776,N_28422);
and U31417 (N_31417,N_28636,N_25495);
and U31418 (N_31418,N_29388,N_26332);
nand U31419 (N_31419,N_27420,N_27477);
xor U31420 (N_31420,N_28598,N_29740);
or U31421 (N_31421,N_28699,N_28183);
nand U31422 (N_31422,N_25150,N_28090);
nor U31423 (N_31423,N_25779,N_27730);
xor U31424 (N_31424,N_25480,N_27220);
and U31425 (N_31425,N_26497,N_25234);
nand U31426 (N_31426,N_26024,N_26091);
nor U31427 (N_31427,N_25205,N_25307);
nand U31428 (N_31428,N_25105,N_29067);
xnor U31429 (N_31429,N_28562,N_26660);
or U31430 (N_31430,N_28000,N_27886);
and U31431 (N_31431,N_27524,N_25803);
or U31432 (N_31432,N_25592,N_29715);
and U31433 (N_31433,N_27707,N_29756);
and U31434 (N_31434,N_29552,N_28981);
or U31435 (N_31435,N_28033,N_26364);
and U31436 (N_31436,N_27415,N_28669);
or U31437 (N_31437,N_29599,N_28092);
or U31438 (N_31438,N_26392,N_29373);
nor U31439 (N_31439,N_29514,N_29796);
or U31440 (N_31440,N_27656,N_29441);
or U31441 (N_31441,N_26827,N_26396);
nand U31442 (N_31442,N_28772,N_25904);
or U31443 (N_31443,N_28663,N_29617);
or U31444 (N_31444,N_28420,N_25404);
nand U31445 (N_31445,N_28854,N_26253);
and U31446 (N_31446,N_25332,N_26089);
and U31447 (N_31447,N_26012,N_26130);
or U31448 (N_31448,N_29196,N_26204);
nand U31449 (N_31449,N_26507,N_28395);
nand U31450 (N_31450,N_29170,N_28362);
nand U31451 (N_31451,N_26607,N_29313);
or U31452 (N_31452,N_28236,N_28973);
nor U31453 (N_31453,N_28311,N_28040);
nor U31454 (N_31454,N_25647,N_29045);
nor U31455 (N_31455,N_28593,N_26786);
nor U31456 (N_31456,N_25683,N_25762);
nand U31457 (N_31457,N_28027,N_28929);
or U31458 (N_31458,N_27297,N_27922);
nand U31459 (N_31459,N_25636,N_25543);
nor U31460 (N_31460,N_25160,N_27893);
and U31461 (N_31461,N_27097,N_29992);
nor U31462 (N_31462,N_25411,N_25058);
nor U31463 (N_31463,N_29557,N_27173);
or U31464 (N_31464,N_25705,N_28102);
nand U31465 (N_31465,N_26636,N_28023);
xor U31466 (N_31466,N_29835,N_28435);
and U31467 (N_31467,N_29464,N_26622);
and U31468 (N_31468,N_28278,N_28135);
xnor U31469 (N_31469,N_28974,N_27032);
and U31470 (N_31470,N_27270,N_28823);
and U31471 (N_31471,N_26847,N_28851);
xor U31472 (N_31472,N_25466,N_25382);
nor U31473 (N_31473,N_25909,N_26790);
or U31474 (N_31474,N_27183,N_26487);
xor U31475 (N_31475,N_26029,N_27052);
nor U31476 (N_31476,N_29474,N_29319);
nand U31477 (N_31477,N_28525,N_25297);
and U31478 (N_31478,N_27591,N_27427);
xor U31479 (N_31479,N_29782,N_27238);
or U31480 (N_31480,N_28378,N_28911);
or U31481 (N_31481,N_28454,N_29743);
nand U31482 (N_31482,N_25324,N_28638);
nand U31483 (N_31483,N_29966,N_25529);
nor U31484 (N_31484,N_25217,N_26117);
and U31485 (N_31485,N_28966,N_27569);
nor U31486 (N_31486,N_26306,N_28286);
nor U31487 (N_31487,N_26735,N_29952);
or U31488 (N_31488,N_25471,N_26541);
or U31489 (N_31489,N_26895,N_27525);
xnor U31490 (N_31490,N_28948,N_27467);
xnor U31491 (N_31491,N_28260,N_27802);
nand U31492 (N_31492,N_26808,N_26999);
nor U31493 (N_31493,N_28976,N_26077);
xnor U31494 (N_31494,N_26701,N_28817);
or U31495 (N_31495,N_29273,N_27632);
nor U31496 (N_31496,N_25089,N_26175);
or U31497 (N_31497,N_27885,N_26264);
nand U31498 (N_31498,N_26685,N_28453);
nand U31499 (N_31499,N_29447,N_26338);
or U31500 (N_31500,N_27542,N_26171);
nand U31501 (N_31501,N_26101,N_28169);
nand U31502 (N_31502,N_27316,N_29107);
and U31503 (N_31503,N_27658,N_27388);
or U31504 (N_31504,N_25391,N_28016);
nand U31505 (N_31505,N_28503,N_25224);
or U31506 (N_31506,N_29255,N_28954);
xor U31507 (N_31507,N_26911,N_26804);
nor U31508 (N_31508,N_28963,N_26923);
xor U31509 (N_31509,N_27419,N_25430);
nor U31510 (N_31510,N_25407,N_25847);
nand U31511 (N_31511,N_28464,N_28264);
and U31512 (N_31512,N_28567,N_28073);
xnor U31513 (N_31513,N_28008,N_29384);
or U31514 (N_31514,N_28869,N_28442);
nand U31515 (N_31515,N_26199,N_26277);
nor U31516 (N_31516,N_25268,N_29202);
xnor U31517 (N_31517,N_26063,N_29240);
nor U31518 (N_31518,N_27949,N_28554);
nand U31519 (N_31519,N_25096,N_25826);
or U31520 (N_31520,N_26647,N_28665);
and U31521 (N_31521,N_29945,N_29147);
and U31522 (N_31522,N_29818,N_28466);
or U31523 (N_31523,N_29977,N_28952);
nor U31524 (N_31524,N_27025,N_27326);
nand U31525 (N_31525,N_25295,N_29596);
nor U31526 (N_31526,N_28516,N_27245);
and U31527 (N_31527,N_29198,N_29274);
or U31528 (N_31528,N_25741,N_26315);
nor U31529 (N_31529,N_27039,N_28044);
and U31530 (N_31530,N_29571,N_25897);
nor U31531 (N_31531,N_29095,N_29554);
or U31532 (N_31532,N_29719,N_29260);
nor U31533 (N_31533,N_29729,N_28589);
and U31534 (N_31534,N_25283,N_26548);
nor U31535 (N_31535,N_29567,N_28075);
nand U31536 (N_31536,N_26577,N_25342);
nor U31537 (N_31537,N_27882,N_26509);
or U31538 (N_31538,N_26311,N_26954);
or U31539 (N_31539,N_28919,N_29690);
nor U31540 (N_31540,N_28605,N_26411);
and U31541 (N_31541,N_28655,N_29306);
xnor U31542 (N_31542,N_28894,N_28879);
nand U31543 (N_31543,N_28734,N_27227);
nor U31544 (N_31544,N_27546,N_29607);
or U31545 (N_31545,N_28630,N_29826);
xor U31546 (N_31546,N_26749,N_26040);
xnor U31547 (N_31547,N_26460,N_29547);
nor U31548 (N_31548,N_28866,N_29843);
nor U31549 (N_31549,N_27126,N_25215);
nand U31550 (N_31550,N_27348,N_26650);
or U31551 (N_31551,N_25369,N_27941);
or U31552 (N_31552,N_25350,N_27148);
and U31553 (N_31553,N_26830,N_28800);
nand U31554 (N_31554,N_28068,N_29280);
xnor U31555 (N_31555,N_28932,N_27398);
nand U31556 (N_31556,N_26765,N_27230);
nor U31557 (N_31557,N_28915,N_29031);
nand U31558 (N_31558,N_25873,N_25086);
and U31559 (N_31559,N_27799,N_26613);
nor U31560 (N_31560,N_29701,N_27529);
or U31561 (N_31561,N_27131,N_26700);
and U31562 (N_31562,N_29517,N_25383);
or U31563 (N_31563,N_28853,N_25729);
or U31564 (N_31564,N_26552,N_25429);
or U31565 (N_31565,N_26908,N_25990);
nand U31566 (N_31566,N_28199,N_26236);
nor U31567 (N_31567,N_25005,N_29858);
and U31568 (N_31568,N_26366,N_25022);
or U31569 (N_31569,N_29742,N_26475);
and U31570 (N_31570,N_28305,N_28937);
nor U31571 (N_31571,N_25233,N_26581);
xnor U31572 (N_31572,N_26892,N_26011);
or U31573 (N_31573,N_29767,N_26815);
or U31574 (N_31574,N_25742,N_26919);
nor U31575 (N_31575,N_28211,N_25125);
or U31576 (N_31576,N_27837,N_25748);
nand U31577 (N_31577,N_27944,N_29523);
nand U31578 (N_31578,N_28139,N_25052);
xor U31579 (N_31579,N_28030,N_29440);
or U31580 (N_31580,N_25938,N_25340);
and U31581 (N_31581,N_29269,N_27749);
or U31582 (N_31582,N_27191,N_28280);
or U31583 (N_31583,N_29588,N_28142);
and U31584 (N_31584,N_29777,N_27224);
nand U31585 (N_31585,N_26148,N_29356);
nand U31586 (N_31586,N_29895,N_27637);
xor U31587 (N_31587,N_27994,N_28697);
and U31588 (N_31588,N_26152,N_25695);
and U31589 (N_31589,N_27888,N_27229);
or U31590 (N_31590,N_26449,N_26347);
nor U31591 (N_31591,N_28679,N_26668);
and U31592 (N_31592,N_27163,N_25533);
nor U31593 (N_31593,N_29691,N_26838);
and U31594 (N_31594,N_25146,N_25824);
nand U31595 (N_31595,N_28967,N_26161);
nor U31596 (N_31596,N_29284,N_26844);
or U31597 (N_31597,N_25521,N_27308);
and U31598 (N_31598,N_29128,N_27576);
and U31599 (N_31599,N_29676,N_27033);
or U31600 (N_31600,N_27600,N_26185);
nand U31601 (N_31601,N_28559,N_27439);
nor U31602 (N_31602,N_27609,N_28519);
xor U31603 (N_31603,N_29267,N_25219);
xnor U31604 (N_31604,N_26861,N_28610);
or U31605 (N_31605,N_26711,N_28776);
and U31606 (N_31606,N_28907,N_26983);
and U31607 (N_31607,N_28709,N_26005);
or U31608 (N_31608,N_29135,N_28750);
or U31609 (N_31609,N_27139,N_26194);
and U31610 (N_31610,N_26299,N_26960);
or U31611 (N_31611,N_27541,N_28587);
and U31612 (N_31612,N_28499,N_26153);
and U31613 (N_31613,N_29718,N_26239);
nand U31614 (N_31614,N_28999,N_25260);
nor U31615 (N_31615,N_27102,N_26826);
nor U31616 (N_31616,N_29674,N_29237);
or U31617 (N_31617,N_27641,N_27579);
nor U31618 (N_31618,N_25092,N_29159);
and U31619 (N_31619,N_27984,N_27493);
and U31620 (N_31620,N_26126,N_29954);
and U31621 (N_31621,N_26083,N_28881);
nor U31622 (N_31622,N_26116,N_26423);
nand U31623 (N_31623,N_25090,N_27844);
nor U31624 (N_31624,N_27267,N_27397);
nand U31625 (N_31625,N_25214,N_29692);
nand U31626 (N_31626,N_28608,N_28575);
or U31627 (N_31627,N_26617,N_25670);
or U31628 (N_31628,N_28018,N_26061);
nand U31629 (N_31629,N_28950,N_27566);
nor U31630 (N_31630,N_28143,N_27982);
nor U31631 (N_31631,N_25401,N_25200);
nor U31632 (N_31632,N_27473,N_25245);
and U31633 (N_31633,N_26404,N_25797);
nand U31634 (N_31634,N_26973,N_26933);
or U31635 (N_31635,N_27505,N_25793);
nor U31636 (N_31636,N_25175,N_29632);
nand U31637 (N_31637,N_25227,N_29525);
and U31638 (N_31638,N_27335,N_26710);
xnor U31639 (N_31639,N_27283,N_27589);
or U31640 (N_31640,N_26974,N_28323);
nor U31641 (N_31641,N_25159,N_27952);
or U31642 (N_31642,N_28418,N_25051);
nor U31643 (N_31643,N_28570,N_25352);
or U31644 (N_31644,N_28548,N_26190);
nand U31645 (N_31645,N_28204,N_26464);
nand U31646 (N_31646,N_27800,N_25922);
or U31647 (N_31647,N_25447,N_25244);
and U31648 (N_31648,N_28085,N_28340);
and U31649 (N_31649,N_28748,N_26495);
nor U31650 (N_31650,N_29443,N_25287);
or U31651 (N_31651,N_29799,N_29489);
xor U31652 (N_31652,N_28756,N_26379);
nor U31653 (N_31653,N_29343,N_28578);
and U31654 (N_31654,N_27466,N_26486);
or U31655 (N_31655,N_29655,N_29314);
or U31656 (N_31656,N_25254,N_25277);
or U31657 (N_31657,N_25104,N_29370);
nand U31658 (N_31658,N_26505,N_29034);
or U31659 (N_31659,N_25264,N_29411);
and U31660 (N_31660,N_29001,N_25142);
nand U31661 (N_31661,N_29659,N_28283);
and U31662 (N_31662,N_28333,N_29623);
and U31663 (N_31663,N_28239,N_28619);
or U31664 (N_31664,N_25869,N_29787);
and U31665 (N_31665,N_28467,N_27341);
nand U31666 (N_31666,N_27640,N_25077);
and U31667 (N_31667,N_29862,N_27483);
nor U31668 (N_31668,N_27787,N_25669);
nand U31669 (N_31669,N_26360,N_26050);
nor U31670 (N_31670,N_29558,N_27539);
nand U31671 (N_31671,N_26174,N_29009);
nand U31672 (N_31672,N_28728,N_27386);
xnor U31673 (N_31673,N_29958,N_26997);
nor U31674 (N_31674,N_26775,N_25027);
xnor U31675 (N_31675,N_26065,N_27647);
nand U31676 (N_31676,N_29544,N_29010);
or U31677 (N_31677,N_25681,N_28875);
and U31678 (N_31678,N_28639,N_29889);
or U31679 (N_31679,N_27138,N_25649);
xnor U31680 (N_31680,N_29662,N_25946);
nand U31681 (N_31681,N_25298,N_25454);
and U31682 (N_31682,N_25648,N_25860);
nor U31683 (N_31683,N_28764,N_29405);
xor U31684 (N_31684,N_29577,N_28479);
and U31685 (N_31685,N_29998,N_26655);
and U31686 (N_31686,N_27856,N_28529);
nand U31687 (N_31687,N_28153,N_25552);
nand U31688 (N_31688,N_27836,N_25598);
or U31689 (N_31689,N_27353,N_25140);
nor U31690 (N_31690,N_28591,N_29788);
and U31691 (N_31691,N_25599,N_28298);
nand U31692 (N_31692,N_28223,N_27932);
or U31693 (N_31693,N_29637,N_26938);
or U31694 (N_31694,N_29253,N_26192);
nand U31695 (N_31695,N_25984,N_26434);
and U31696 (N_31696,N_25968,N_25910);
or U31697 (N_31697,N_27216,N_25940);
or U31698 (N_31698,N_25809,N_25002);
nand U31699 (N_31699,N_29133,N_28154);
nor U31700 (N_31700,N_26147,N_29823);
nor U31701 (N_31701,N_28867,N_28912);
or U31702 (N_31702,N_27639,N_27369);
xor U31703 (N_31703,N_27261,N_29057);
xor U31704 (N_31704,N_28253,N_27422);
nand U31705 (N_31705,N_26228,N_28355);
nand U31706 (N_31706,N_27495,N_25435);
and U31707 (N_31707,N_27835,N_25093);
or U31708 (N_31708,N_29178,N_28996);
xnor U31709 (N_31709,N_28113,N_28312);
or U31710 (N_31710,N_25011,N_29668);
xor U31711 (N_31711,N_26378,N_27887);
nor U31712 (N_31712,N_29928,N_28758);
and U31713 (N_31713,N_28592,N_26903);
and U31714 (N_31714,N_27107,N_25894);
nand U31715 (N_31715,N_26436,N_25682);
nand U31716 (N_31716,N_27795,N_25004);
or U31717 (N_31717,N_27811,N_25646);
and U31718 (N_31718,N_28403,N_28760);
nand U31719 (N_31719,N_29295,N_27895);
nor U31720 (N_31720,N_29618,N_26528);
nand U31721 (N_31721,N_28335,N_25156);
xor U31722 (N_31722,N_27065,N_28276);
and U31723 (N_31723,N_29457,N_26508);
nor U31724 (N_31724,N_25076,N_27877);
nor U31725 (N_31725,N_27171,N_26994);
xnor U31726 (N_31726,N_25064,N_25236);
nor U31727 (N_31727,N_28173,N_28046);
or U31728 (N_31728,N_28740,N_28210);
nand U31729 (N_31729,N_26673,N_27128);
nand U31730 (N_31730,N_26276,N_25626);
nand U31731 (N_31731,N_26618,N_27918);
and U31732 (N_31732,N_25633,N_29615);
xnor U31733 (N_31733,N_28642,N_29583);
and U31734 (N_31734,N_28902,N_27849);
nand U31735 (N_31735,N_25151,N_29688);
or U31736 (N_31736,N_28887,N_27480);
and U31737 (N_31737,N_29886,N_26340);
and U31738 (N_31738,N_27465,N_25974);
and U31739 (N_31739,N_25888,N_26481);
or U31740 (N_31740,N_29541,N_28331);
or U31741 (N_31741,N_26631,N_27162);
or U31742 (N_31742,N_28840,N_28374);
nor U31743 (N_31743,N_27149,N_26208);
nor U31744 (N_31744,N_26386,N_26413);
or U31745 (N_31745,N_25752,N_29815);
and U31746 (N_31746,N_26212,N_27872);
nor U31747 (N_31747,N_25887,N_27248);
xnor U31748 (N_31748,N_28877,N_29453);
nor U31749 (N_31749,N_27765,N_29563);
or U31750 (N_31750,N_29683,N_26125);
and U31751 (N_31751,N_25240,N_29299);
nor U31752 (N_31752,N_27475,N_25358);
and U31753 (N_31753,N_25165,N_25663);
nand U31754 (N_31754,N_25428,N_29981);
or U31755 (N_31755,N_29785,N_25133);
nor U31756 (N_31756,N_25872,N_27617);
and U31757 (N_31757,N_28691,N_28622);
nand U31758 (N_31758,N_28841,N_27610);
or U31759 (N_31759,N_27873,N_25571);
xor U31760 (N_31760,N_26104,N_26713);
nor U31761 (N_31761,N_29555,N_25136);
nand U31762 (N_31762,N_29419,N_27299);
nand U31763 (N_31763,N_26030,N_29559);
or U31764 (N_31764,N_27889,N_27702);
or U31765 (N_31765,N_26303,N_25697);
nand U31766 (N_31766,N_28167,N_27223);
nor U31767 (N_31767,N_27709,N_28328);
nand U31768 (N_31768,N_28935,N_28518);
and U31769 (N_31769,N_28318,N_29479);
nor U31770 (N_31770,N_27056,N_27715);
xnor U31771 (N_31771,N_29234,N_29454);
and U31772 (N_31772,N_26337,N_26691);
nand U31773 (N_31773,N_26346,N_25747);
or U31774 (N_31774,N_25726,N_29104);
or U31775 (N_31775,N_25623,N_28814);
nand U31776 (N_31776,N_25801,N_25898);
xor U31777 (N_31777,N_29663,N_25048);
or U31778 (N_31778,N_29585,N_29916);
nor U31779 (N_31779,N_26694,N_29844);
or U31780 (N_31780,N_27857,N_29473);
nor U31781 (N_31781,N_27671,N_25660);
nor U31782 (N_31782,N_27464,N_29925);
nor U31783 (N_31783,N_29174,N_26314);
and U31784 (N_31784,N_27226,N_28601);
and U31785 (N_31785,N_28702,N_27350);
and U31786 (N_31786,N_27798,N_28580);
xnor U31787 (N_31787,N_28279,N_29363);
nor U31788 (N_31788,N_27264,N_26201);
nand U31789 (N_31789,N_28473,N_26658);
nand U31790 (N_31790,N_27344,N_29430);
nor U31791 (N_31791,N_27636,N_28036);
or U31792 (N_31792,N_26839,N_29231);
and U31793 (N_31793,N_26373,N_29089);
or U31794 (N_31794,N_25539,N_28238);
nor U31795 (N_31795,N_25356,N_26987);
or U31796 (N_31796,N_25906,N_25377);
nor U31797 (N_31797,N_29593,N_27793);
nand U31798 (N_31798,N_28635,N_28063);
and U31799 (N_31799,N_27147,N_28379);
nor U31800 (N_31800,N_28766,N_27239);
and U31801 (N_31801,N_29181,N_25673);
nand U31802 (N_31802,N_27281,N_25768);
nand U31803 (N_31803,N_25662,N_26885);
nor U31804 (N_31804,N_25498,N_29355);
nor U31805 (N_31805,N_28941,N_28212);
nor U31806 (N_31806,N_29781,N_26443);
nand U31807 (N_31807,N_26737,N_29292);
and U31808 (N_31808,N_28590,N_25098);
and U31809 (N_31809,N_25537,N_29707);
nor U31810 (N_31810,N_28644,N_27117);
or U31811 (N_31811,N_29002,N_27980);
or U31812 (N_31812,N_26352,N_26059);
nand U31813 (N_31813,N_25664,N_26243);
nand U31814 (N_31814,N_29099,N_29658);
nor U31815 (N_31815,N_28221,N_28822);
nor U31816 (N_31816,N_26453,N_28909);
nand U31817 (N_31817,N_25881,N_29227);
or U31818 (N_31818,N_25916,N_25211);
nor U31819 (N_31819,N_27733,N_27190);
or U31820 (N_31820,N_27199,N_27955);
and U31821 (N_31821,N_25346,N_25266);
nor U31822 (N_31822,N_29192,N_27489);
nand U31823 (N_31823,N_26985,N_27747);
or U31824 (N_31824,N_25390,N_27677);
xor U31825 (N_31825,N_25926,N_28186);
xnor U31826 (N_31826,N_25632,N_27621);
or U31827 (N_31827,N_27108,N_27925);
nor U31828 (N_31828,N_26007,N_29963);
or U31829 (N_31829,N_27976,N_27969);
or U31830 (N_31830,N_25196,N_28809);
xnor U31831 (N_31831,N_29381,N_25690);
or U31832 (N_31832,N_27342,N_27518);
nand U31833 (N_31833,N_27425,N_26382);
nor U31834 (N_31834,N_28031,N_26031);
nor U31835 (N_31835,N_28891,N_25269);
nor U31836 (N_31836,N_26020,N_28545);
nand U31837 (N_31837,N_28176,N_26428);
or U31838 (N_31838,N_27841,N_28674);
nor U31839 (N_31839,N_26222,N_26483);
nor U31840 (N_31840,N_26210,N_25749);
nor U31841 (N_31841,N_29549,N_26873);
or U31842 (N_31842,N_26128,N_25302);
nor U31843 (N_31843,N_26663,N_25818);
nor U31844 (N_31844,N_25584,N_29242);
nand U31845 (N_31845,N_25728,N_25538);
nand U31846 (N_31846,N_27068,N_25849);
nand U31847 (N_31847,N_28727,N_27169);
and U31848 (N_31848,N_25800,N_26144);
nor U31849 (N_31849,N_29069,N_25996);
nand U31850 (N_31850,N_28700,N_26560);
xnor U31851 (N_31851,N_25629,N_29574);
nor U31852 (N_31852,N_29562,N_28447);
or U31853 (N_31853,N_28938,N_25185);
or U31854 (N_31854,N_28009,N_25661);
nor U31855 (N_31855,N_27890,N_29251);
nor U31856 (N_31856,N_25387,N_27242);
nor U31857 (N_31857,N_28534,N_27192);
or U31858 (N_31858,N_25861,N_25181);
and U31859 (N_31859,N_28320,N_25640);
and U31860 (N_31860,N_27690,N_29738);
nor U31861 (N_31861,N_28215,N_29851);
xnor U31862 (N_31862,N_26539,N_28393);
and U31863 (N_31863,N_29412,N_25225);
nor U31864 (N_31864,N_28156,N_26530);
or U31865 (N_31865,N_28629,N_25757);
xor U31866 (N_31866,N_25671,N_27445);
nand U31867 (N_31867,N_29155,N_26670);
or U31868 (N_31868,N_29901,N_26858);
xor U31869 (N_31869,N_28990,N_29033);
and U31870 (N_31870,N_25129,N_26852);
and U31871 (N_31871,N_28683,N_27808);
and U31872 (N_31872,N_25927,N_28647);
and U31873 (N_31873,N_27105,N_25168);
or U31874 (N_31874,N_28469,N_29846);
or U31875 (N_31875,N_25732,N_27627);
xnor U31876 (N_31876,N_28720,N_28277);
and U31877 (N_31877,N_26260,N_27289);
or U31878 (N_31878,N_29353,N_28786);
or U31879 (N_31879,N_26071,N_27917);
and U31880 (N_31880,N_27655,N_29877);
nor U31881 (N_31881,N_29129,N_25925);
nand U31882 (N_31882,N_29125,N_29987);
or U31883 (N_31883,N_26062,N_26526);
nand U31884 (N_31884,N_26963,N_29551);
nor U31885 (N_31885,N_27563,N_27492);
nand U31886 (N_31886,N_28319,N_27247);
nor U31887 (N_31887,N_26422,N_25986);
or U31888 (N_31888,N_28441,N_29414);
or U31889 (N_31889,N_26351,N_25153);
and U31890 (N_31890,N_25108,N_28988);
or U31891 (N_31891,N_25870,N_25270);
or U31892 (N_31892,N_29580,N_28532);
nand U31893 (N_31893,N_28804,N_28407);
xor U31894 (N_31894,N_29451,N_26188);
nor U31895 (N_31895,N_28443,N_25721);
nand U31896 (N_31896,N_28505,N_26427);
nor U31897 (N_31897,N_26296,N_27150);
nand U31898 (N_31898,N_28304,N_26747);
and U31899 (N_31899,N_29455,N_26358);
nor U31900 (N_31900,N_29283,N_25213);
or U31901 (N_31901,N_28426,N_28126);
or U31902 (N_31902,N_28011,N_25103);
xnor U31903 (N_31903,N_25322,N_29035);
xor U31904 (N_31904,N_28836,N_27575);
nand U31905 (N_31905,N_29493,N_28746);
or U31906 (N_31906,N_29054,N_25746);
nor U31907 (N_31907,N_28595,N_25578);
nor U31908 (N_31908,N_29042,N_25313);
nand U31909 (N_31909,N_28744,N_25014);
nand U31910 (N_31910,N_25056,N_26992);
nor U31911 (N_31911,N_26095,N_29903);
and U31912 (N_31912,N_28125,N_27915);
or U31913 (N_31913,N_28681,N_26105);
nand U31914 (N_31914,N_28388,N_28310);
nor U31915 (N_31915,N_29177,N_25128);
nor U31916 (N_31916,N_28222,N_27443);
nor U31917 (N_31917,N_27203,N_25912);
or U31918 (N_31918,N_29795,N_26292);
or U31919 (N_31919,N_29494,N_29028);
nor U31920 (N_31920,N_29342,N_26120);
xnor U31921 (N_31921,N_29495,N_25761);
or U31922 (N_31922,N_28065,N_27606);
nor U31923 (N_31923,N_27936,N_29509);
or U31924 (N_31924,N_25790,N_26035);
nand U31925 (N_31925,N_25221,N_25606);
nor U31926 (N_31926,N_29937,N_26851);
and U31927 (N_31927,N_28366,N_28324);
or U31928 (N_31928,N_27777,N_28606);
or U31929 (N_31929,N_25615,N_27474);
xor U31930 (N_31930,N_29789,N_25373);
nor U31931 (N_31931,N_25468,N_26013);
nand U31932 (N_31932,N_25441,N_27931);
xor U31933 (N_31933,N_25033,N_26217);
xnor U31934 (N_31934,N_28105,N_26173);
nor U31935 (N_31935,N_29126,N_25453);
nand U31936 (N_31936,N_25602,N_26066);
or U31937 (N_31937,N_28594,N_29773);
or U31938 (N_31938,N_27989,N_27345);
nor U31939 (N_31939,N_28416,N_28997);
or U31940 (N_31940,N_28087,N_28246);
and U31941 (N_31941,N_28944,N_29277);
or U31942 (N_31942,N_26813,N_25506);
and U31943 (N_31943,N_25243,N_25393);
nor U31944 (N_31944,N_27545,N_26998);
and U31945 (N_31945,N_27851,N_29140);
or U31946 (N_31946,N_25210,N_27044);
nand U31947 (N_31947,N_29166,N_29797);
or U31948 (N_31948,N_27878,N_25945);
and U31949 (N_31949,N_26145,N_25438);
nor U31950 (N_31950,N_26215,N_29291);
nand U31951 (N_31951,N_29322,N_28995);
or U31952 (N_31952,N_26028,N_27011);
nor U31953 (N_31953,N_25704,N_29819);
nand U31954 (N_31954,N_25097,N_26019);
and U31955 (N_31955,N_28819,N_29648);
or U31956 (N_31956,N_26143,N_27387);
or U31957 (N_31957,N_26944,N_27997);
nand U31958 (N_31958,N_27814,N_26108);
and U31959 (N_31959,N_26385,N_28928);
or U31960 (N_31960,N_27006,N_25856);
nor U31961 (N_31961,N_28901,N_28586);
nor U31962 (N_31962,N_29880,N_28737);
nor U31963 (N_31963,N_26986,N_29245);
nor U31964 (N_31964,N_28163,N_25591);
xor U31965 (N_31965,N_26450,N_28299);
xor U31966 (N_31966,N_28918,N_25707);
nor U31967 (N_31967,N_29759,N_25773);
or U31968 (N_31968,N_28381,N_27321);
nor U31969 (N_31969,N_29955,N_26394);
and U31970 (N_31970,N_25966,N_28883);
or U31971 (N_31971,N_29335,N_28528);
nor U31972 (N_31972,N_28015,N_25394);
nor U31973 (N_31973,N_28671,N_27088);
or U31974 (N_31974,N_28512,N_27822);
nor U31975 (N_31975,N_29290,N_28904);
nor U31976 (N_31976,N_27661,N_26989);
nand U31977 (N_31977,N_29055,N_28704);
nand U31978 (N_31978,N_25557,N_26354);
and U31979 (N_31979,N_28001,N_29275);
and U31980 (N_31980,N_29139,N_27054);
xor U31981 (N_31981,N_26679,N_28292);
and U31982 (N_31982,N_27788,N_25144);
nor U31983 (N_31983,N_27960,N_28863);
nor U31984 (N_31984,N_27401,N_29784);
nor U31985 (N_31985,N_28785,N_25278);
and U31986 (N_31986,N_25059,N_29175);
or U31987 (N_31987,N_25866,N_27210);
and U31988 (N_31988,N_28187,N_29587);
and U31989 (N_31989,N_26390,N_27643);
and U31990 (N_31990,N_25176,N_26656);
xnor U31991 (N_31991,N_28620,N_28141);
nor U31992 (N_31992,N_29059,N_29798);
or U31993 (N_31993,N_28097,N_25734);
and U31994 (N_31994,N_25855,N_29017);
nor U31995 (N_31995,N_26651,N_29669);
and U31996 (N_31996,N_28225,N_25410);
xor U31997 (N_31997,N_26371,N_29528);
nor U31998 (N_31998,N_29425,N_26657);
nand U31999 (N_31999,N_25001,N_29848);
nor U32000 (N_32000,N_25024,N_27527);
xor U32001 (N_32001,N_26832,N_28980);
nor U32002 (N_32002,N_28117,N_25617);
or U32003 (N_32003,N_26437,N_26995);
nand U32004 (N_32004,N_26424,N_27734);
nor U32005 (N_32005,N_25643,N_29458);
or U32006 (N_32006,N_27928,N_26598);
and U32007 (N_32007,N_27244,N_27042);
xnor U32008 (N_32008,N_28334,N_25201);
nand U32009 (N_32009,N_26665,N_26930);
nand U32010 (N_32010,N_26139,N_28268);
nor U32011 (N_32011,N_27319,N_25634);
nand U32012 (N_32012,N_25684,N_27023);
nor U32013 (N_32013,N_25550,N_25481);
nor U32014 (N_32014,N_29301,N_28701);
and U32015 (N_32015,N_26599,N_26482);
and U32016 (N_32016,N_25831,N_29813);
and U32017 (N_32017,N_26472,N_27754);
nand U32018 (N_32018,N_27669,N_27506);
and U32019 (N_32019,N_28140,N_27757);
xnor U32020 (N_32020,N_28738,N_25832);
and U32021 (N_32021,N_27060,N_26907);
or U32022 (N_32022,N_26377,N_25919);
or U32023 (N_32023,N_26405,N_28788);
or U32024 (N_32024,N_29459,N_29376);
nor U32025 (N_32025,N_26133,N_29150);
xnor U32026 (N_32026,N_29824,N_25182);
and U32027 (N_32027,N_27830,N_26962);
and U32028 (N_32028,N_29985,N_25461);
nand U32029 (N_32029,N_25169,N_27167);
xnor U32030 (N_32030,N_29949,N_27691);
nand U32031 (N_32031,N_28265,N_26180);
and U32032 (N_32032,N_28281,N_27848);
xor U32033 (N_32033,N_28645,N_25989);
and U32034 (N_32034,N_27251,N_28811);
or U32035 (N_32035,N_25782,N_25877);
or U32036 (N_32036,N_29639,N_25025);
nor U32037 (N_32037,N_25310,N_28569);
nor U32038 (N_32038,N_28088,N_28256);
xnor U32039 (N_32039,N_25754,N_28483);
nand U32040 (N_32040,N_29325,N_25596);
or U32041 (N_32041,N_25188,N_27760);
or U32042 (N_32042,N_27312,N_26893);
nor U32043 (N_32043,N_29475,N_29331);
nor U32044 (N_32044,N_26326,N_27029);
and U32045 (N_32045,N_26480,N_26945);
and U32046 (N_32046,N_25158,N_25614);
nand U32047 (N_32047,N_29449,N_26184);
xor U32048 (N_32048,N_28889,N_27165);
xnor U32049 (N_32049,N_28808,N_29634);
nand U32050 (N_32050,N_25724,N_28718);
or U32051 (N_32051,N_29675,N_25788);
nor U32052 (N_32052,N_29195,N_27809);
or U32053 (N_32053,N_29066,N_25184);
or U32054 (N_32054,N_25117,N_27946);
and U32055 (N_32055,N_28947,N_27717);
or U32056 (N_32056,N_29988,N_29409);
xor U32057 (N_32057,N_28081,N_27679);
xor U32058 (N_32058,N_29392,N_28632);
and U32059 (N_32059,N_25568,N_25045);
nand U32060 (N_32060,N_27874,N_25512);
or U32061 (N_32061,N_28042,N_26565);
xnor U32062 (N_32062,N_26466,N_29939);
nand U32063 (N_32063,N_27585,N_25677);
and U32064 (N_32064,N_26498,N_26266);
and U32065 (N_32065,N_29064,N_26555);
nor U32066 (N_32066,N_25423,N_26924);
and U32067 (N_32067,N_28914,N_25835);
nor U32068 (N_32068,N_29803,N_29628);
xnor U32069 (N_32069,N_26943,N_28417);
and U32070 (N_32070,N_28789,N_28796);
nand U32071 (N_32071,N_29439,N_29817);
nor U32072 (N_32072,N_29764,N_25580);
nor U32073 (N_32073,N_29775,N_25769);
and U32074 (N_32074,N_29276,N_27091);
or U32075 (N_32075,N_29145,N_25893);
nand U32076 (N_32076,N_28439,N_26864);
xnor U32077 (N_32077,N_26993,N_26831);
nor U32078 (N_32078,N_26490,N_28685);
or U32079 (N_32079,N_25250,N_27562);
and U32080 (N_32080,N_26407,N_28762);
or U32081 (N_32081,N_28922,N_29173);
or U32082 (N_32082,N_26784,N_25367);
nor U32083 (N_32083,N_25931,N_27273);
and U32084 (N_32084,N_27200,N_27686);
nor U32085 (N_32085,N_28263,N_27182);
nand U32086 (N_32086,N_26051,N_27198);
nand U32087 (N_32087,N_26461,N_27061);
nor U32088 (N_32088,N_25653,N_29631);
and U32089 (N_32089,N_28007,N_28217);
and U32090 (N_32090,N_27821,N_25582);
nand U32091 (N_32091,N_26645,N_29131);
nand U32092 (N_32092,N_25137,N_27706);
and U32093 (N_32093,N_28259,N_27523);
and U32094 (N_32094,N_27084,N_28290);
nor U32095 (N_32095,N_25354,N_28695);
nand U32096 (N_32096,N_25279,N_26736);
nand U32097 (N_32097,N_26406,N_26833);
and U32098 (N_32098,N_29005,N_28923);
or U32099 (N_32099,N_27638,N_29308);
nand U32100 (N_32100,N_27789,N_25585);
nand U32101 (N_32101,N_25046,N_29106);
and U32102 (N_32102,N_27311,N_26868);
nor U32103 (N_32103,N_28228,N_25362);
nor U32104 (N_32104,N_27405,N_25559);
or U32105 (N_32105,N_28710,N_25808);
xnor U32106 (N_32106,N_27417,N_29326);
nand U32107 (N_32107,N_28401,N_25665);
xnor U32108 (N_32108,N_28542,N_27581);
nor U32109 (N_32109,N_25115,N_28151);
nand U32110 (N_32110,N_29769,N_26220);
or U32111 (N_32111,N_25433,N_26569);
nor U32112 (N_32112,N_27560,N_26112);
nand U32113 (N_32113,N_28537,N_26078);
nand U32114 (N_32114,N_28098,N_28041);
and U32115 (N_32115,N_28043,N_29452);
or U32116 (N_32116,N_25879,N_27650);
xnor U32117 (N_32117,N_29220,N_27682);
nor U32118 (N_32118,N_27298,N_27700);
nor U32119 (N_32119,N_27729,N_25178);
xnor U32120 (N_32120,N_27358,N_26287);
or U32121 (N_32121,N_25844,N_29931);
nor U32122 (N_32122,N_26265,N_27520);
nand U32123 (N_32123,N_28682,N_27240);
and U32124 (N_32124,N_27736,N_27776);
nor U32125 (N_32125,N_28371,N_28676);
nor U32126 (N_32126,N_28248,N_28609);
and U32127 (N_32127,N_26512,N_28987);
and U32128 (N_32128,N_29197,N_27459);
nand U32129 (N_32129,N_28038,N_26412);
and U32130 (N_32130,N_27450,N_28243);
and U32131 (N_32131,N_28461,N_25933);
nor U32132 (N_32132,N_26699,N_27728);
xnor U32133 (N_32133,N_25305,N_27153);
and U32134 (N_32134,N_29686,N_29586);
and U32135 (N_32135,N_25589,N_26900);
xnor U32136 (N_32136,N_28034,N_25525);
and U32137 (N_32137,N_25044,N_26920);
nor U32138 (N_32138,N_29837,N_28581);
nand U32139 (N_32139,N_27914,N_28035);
and U32140 (N_32140,N_25961,N_29478);
or U32141 (N_32141,N_25357,N_29460);
nor U32142 (N_32142,N_27724,N_29109);
xnor U32143 (N_32143,N_26705,N_27860);
and U32144 (N_32144,N_28812,N_27945);
nor U32145 (N_32145,N_29350,N_28552);
and U32146 (N_32146,N_29492,N_29073);
nand U32147 (N_32147,N_27363,N_28106);
and U32148 (N_32148,N_25920,N_28481);
nor U32149 (N_32149,N_25364,N_29102);
nor U32150 (N_32150,N_29281,N_29030);
nor U32151 (N_32151,N_29650,N_26592);
nor U32152 (N_32152,N_29927,N_25943);
or U32153 (N_32153,N_29421,N_27622);
and U32154 (N_32154,N_25118,N_29330);
nor U32155 (N_32155,N_28152,N_27383);
nor U32156 (N_32156,N_29039,N_27337);
nor U32157 (N_32157,N_27720,N_25709);
nand U32158 (N_32158,N_26918,N_26758);
or U32159 (N_32159,N_29212,N_29018);
or U32160 (N_32160,N_25348,N_25520);
and U32161 (N_32161,N_26566,N_27377);
nand U32162 (N_32162,N_26416,N_29207);
nand U32163 (N_32163,N_28322,N_29581);
xnor U32164 (N_32164,N_25507,N_29869);
and U32165 (N_32165,N_29300,N_29999);
nand U32166 (N_32166,N_26010,N_27722);
nor U32167 (N_32167,N_29091,N_28991);
and U32168 (N_32168,N_29305,N_29094);
nand U32169 (N_32169,N_28509,N_26982);
nor U32170 (N_32170,N_26738,N_26046);
nand U32171 (N_32171,N_25304,N_28055);
or U32172 (N_32172,N_29702,N_26531);
or U32173 (N_32173,N_29699,N_26355);
xnor U32174 (N_32174,N_28678,N_27876);
xnor U32175 (N_32175,N_27684,N_25777);
xnor U32176 (N_32176,N_29485,N_25170);
or U32177 (N_32177,N_27320,N_28493);
and U32178 (N_32178,N_29491,N_27087);
nand U32179 (N_32179,N_25081,N_27597);
or U32180 (N_32180,N_25994,N_28672);
or U32181 (N_32181,N_26971,N_29399);
or U32182 (N_32182,N_28896,N_29883);
nand U32183 (N_32183,N_27045,N_28351);
nor U32184 (N_32184,N_27564,N_28005);
and U32185 (N_32185,N_26524,N_28039);
nand U32186 (N_32186,N_25195,N_26940);
nand U32187 (N_32187,N_26935,N_29641);
nor U32188 (N_32188,N_26787,N_27901);
nor U32189 (N_32189,N_25427,N_29827);
nor U32190 (N_32190,N_26518,N_25511);
and U32191 (N_32191,N_25911,N_26334);
and U32192 (N_32192,N_27502,N_25177);
and U32193 (N_32193,N_26766,N_27232);
nor U32194 (N_32194,N_27595,N_27721);
nand U32195 (N_32195,N_28646,N_27742);
nand U32196 (N_32196,N_26310,N_28726);
and U32197 (N_32197,N_28634,N_26417);
and U32198 (N_32198,N_27756,N_29383);
nand U32199 (N_32199,N_28354,N_27759);
and U32200 (N_32200,N_26098,N_25740);
or U32201 (N_32201,N_26036,N_26219);
nor U32202 (N_32202,N_28574,N_29084);
nor U32203 (N_32203,N_27382,N_27864);
nand U32204 (N_32204,N_28880,N_25579);
or U32205 (N_32205,N_27303,N_25937);
or U32206 (N_32206,N_28491,N_25256);
xor U32207 (N_32207,N_26270,N_25722);
or U32208 (N_32208,N_28421,N_28657);
and U32209 (N_32209,N_28478,N_28208);
xnor U32210 (N_32210,N_29714,N_28972);
nand U32211 (N_32211,N_28330,N_29244);
or U32212 (N_32212,N_28244,N_27723);
nand U32213 (N_32213,N_25637,N_25360);
nor U32214 (N_32214,N_26397,N_27260);
nand U32215 (N_32215,N_29038,N_29831);
nand U32216 (N_32216,N_29080,N_25631);
and U32217 (N_32217,N_26131,N_25569);
and U32218 (N_32218,N_29739,N_28616);
xor U32219 (N_32219,N_29652,N_29081);
nand U32220 (N_32220,N_27847,N_28925);
or U32221 (N_32221,N_29532,N_27510);
or U32222 (N_32222,N_27118,N_25079);
nand U32223 (N_32223,N_29520,N_29431);
or U32224 (N_32224,N_27863,N_29351);
nand U32225 (N_32225,N_27801,N_29920);
nor U32226 (N_32226,N_27565,N_26107);
or U32227 (N_32227,N_27083,N_25565);
and U32228 (N_32228,N_28715,N_27446);
or U32229 (N_32229,N_27549,N_27827);
and U32230 (N_32230,N_25995,N_26211);
or U32231 (N_32231,N_25874,N_28250);
nand U32232 (N_32232,N_25375,N_25445);
xor U32233 (N_32233,N_28857,N_26988);
nand U32234 (N_32234,N_26032,N_25560);
nor U32235 (N_32235,N_28332,N_28022);
and U32236 (N_32236,N_26281,N_28284);
nor U32237 (N_32237,N_29043,N_25237);
or U32238 (N_32238,N_27236,N_29713);
nor U32239 (N_32239,N_27266,N_26043);
nand U32240 (N_32240,N_27176,N_26770);
xor U32241 (N_32241,N_28069,N_27368);
or U32242 (N_32242,N_27719,N_25154);
or U32243 (N_32243,N_29210,N_26380);
or U32244 (N_32244,N_27218,N_27484);
xnor U32245 (N_32245,N_27135,N_27543);
nor U32246 (N_32246,N_28192,N_29229);
or U32247 (N_32247,N_27842,N_26800);
and U32248 (N_32248,N_29660,N_25418);
and U32249 (N_32249,N_26006,N_29206);
xnor U32250 (N_32250,N_27660,N_25281);
and U32251 (N_32251,N_28449,N_26096);
nand U32252 (N_32252,N_25523,N_26099);
and U32253 (N_32253,N_26537,N_26027);
or U32254 (N_32254,N_28132,N_28979);
nand U32255 (N_32255,N_27587,N_26288);
nor U32256 (N_32256,N_29075,N_25068);
xnor U32257 (N_32257,N_28348,N_29917);
nor U32258 (N_32258,N_27557,N_29849);
or U32259 (N_32259,N_25973,N_26689);
nand U32260 (N_32260,N_26750,N_29422);
or U32261 (N_32261,N_27187,N_26448);
nand U32262 (N_32262,N_27433,N_25378);
xnor U32263 (N_32263,N_27201,N_29337);
and U32264 (N_32264,N_27670,N_28992);
or U32265 (N_32265,N_28429,N_29991);
or U32266 (N_32266,N_25611,N_26774);
xor U32267 (N_32267,N_25229,N_27561);
nand U32268 (N_32268,N_25957,N_27846);
nand U32269 (N_32269,N_26771,N_29254);
nand U32270 (N_32270,N_27463,N_26240);
nor U32271 (N_32271,N_26797,N_26205);
nand U32272 (N_32272,N_26293,N_29984);
and U32273 (N_32273,N_27970,N_27036);
or U32274 (N_32274,N_27144,N_26589);
xnor U32275 (N_32275,N_28122,N_25952);
or U32276 (N_32276,N_29930,N_28465);
or U32277 (N_32277,N_29760,N_27079);
xnor U32278 (N_32278,N_27421,N_28170);
nand U32279 (N_32279,N_26821,N_29621);
nand U32280 (N_32280,N_25148,N_26255);
nand U32281 (N_32281,N_26783,N_29182);
and U32282 (N_32282,N_28878,N_27442);
nor U32283 (N_32283,N_28352,N_27929);
nand U32284 (N_32284,N_26977,N_27287);
or U32285 (N_32285,N_26129,N_26018);
and U32286 (N_32286,N_28717,N_27195);
or U32287 (N_32287,N_27047,N_28989);
and U32288 (N_32288,N_26168,N_27879);
or U32289 (N_32289,N_29636,N_28361);
nand U32290 (N_32290,N_27704,N_29929);
or U32291 (N_32291,N_26181,N_27688);
or U32292 (N_32292,N_26501,N_26278);
nand U32293 (N_32293,N_25928,N_26748);
or U32294 (N_32294,N_29522,N_27951);
nor U32295 (N_32295,N_27174,N_29444);
nand U32296 (N_32296,N_28856,N_29168);
nor U32297 (N_32297,N_25929,N_25272);
or U32298 (N_32298,N_27906,N_29304);
nor U32299 (N_32299,N_25963,N_27043);
and U32300 (N_32300,N_29390,N_26968);
nor U32301 (N_32301,N_26761,N_27376);
and U32302 (N_32302,N_28945,N_27644);
nor U32303 (N_32303,N_28123,N_27676);
or U32304 (N_32304,N_28406,N_28784);
nand U32305 (N_32305,N_26881,N_25426);
or U32306 (N_32306,N_28767,N_29598);
and U32307 (N_32307,N_25918,N_29983);
nand U32308 (N_32308,N_29278,N_25282);
and U32309 (N_32309,N_25715,N_25992);
nor U32310 (N_32310,N_26154,N_26248);
nor U32311 (N_32311,N_25460,N_27180);
nor U32312 (N_32312,N_26970,N_26435);
or U32313 (N_32313,N_26630,N_26014);
or U32314 (N_32314,N_27189,N_26513);
nand U32315 (N_32315,N_29922,N_29971);
nor U32316 (N_32316,N_27123,N_27990);
or U32317 (N_32317,N_27209,N_29401);
or U32318 (N_32318,N_25587,N_29608);
nand U32319 (N_32319,N_27659,N_28779);
nand U32320 (N_32320,N_29247,N_25955);
nor U32321 (N_32321,N_28431,N_25792);
xor U32322 (N_32322,N_25021,N_29986);
and U32323 (N_32323,N_25902,N_28364);
nand U32324 (N_32324,N_25173,N_28112);
nand U32325 (N_32325,N_25621,N_26305);
nor U32326 (N_32326,N_26177,N_25499);
or U32327 (N_32327,N_26925,N_25497);
xor U32328 (N_32328,N_29834,N_26231);
and U32329 (N_32329,N_28137,N_29513);
or U32330 (N_32330,N_29036,N_26041);
or U32331 (N_32331,N_28425,N_29762);
nand U32332 (N_32332,N_26959,N_28712);
and U32333 (N_32333,N_25515,N_25531);
nand U32334 (N_32334,N_27172,N_28201);
and U32335 (N_32335,N_25066,N_29622);
nand U32336 (N_32336,N_29354,N_28526);
nor U32337 (N_32337,N_25886,N_29911);
nor U32338 (N_32338,N_26732,N_28294);
or U32339 (N_32339,N_28257,N_27572);
or U32340 (N_32340,N_29481,N_26164);
or U32341 (N_32341,N_25368,N_27018);
xnor U32342 (N_32342,N_26603,N_26291);
nand U32343 (N_32343,N_26186,N_28218);
nand U32344 (N_32344,N_29171,N_28692);
nand U32345 (N_32345,N_26871,N_28564);
or U32346 (N_32346,N_29394,N_27689);
nor U32347 (N_32347,N_28254,N_25787);
xor U32348 (N_32348,N_25935,N_28168);
or U32349 (N_32349,N_25685,N_27041);
nand U32350 (N_32350,N_25434,N_27731);
and U32351 (N_32351,N_26723,N_28969);
or U32352 (N_32352,N_25985,N_28350);
nand U32353 (N_32353,N_29828,N_25865);
or U32354 (N_32354,N_26280,N_27673);
nor U32355 (N_32355,N_26350,N_28975);
nor U32356 (N_32356,N_27536,N_26045);
or U32357 (N_32357,N_26810,N_26368);
and U32358 (N_32358,N_27735,N_28613);
or U32359 (N_32359,N_27519,N_25327);
or U32360 (N_32360,N_25967,N_27680);
nand U32361 (N_32361,N_25519,N_25725);
xor U32362 (N_32362,N_27212,N_28773);
xnor U32363 (N_32363,N_28805,N_25567);
and U32364 (N_32364,N_29898,N_29620);
nand U32365 (N_32365,N_25061,N_29143);
xor U32366 (N_32366,N_25311,N_29548);
nor U32367 (N_32367,N_29974,N_25875);
nor U32368 (N_32368,N_26878,N_25012);
and U32369 (N_32369,N_26633,N_29610);
xor U32370 (N_32370,N_26609,N_29710);
xnor U32371 (N_32371,N_29161,N_27559);
nand U32372 (N_32372,N_26259,N_29410);
xnor U32373 (N_32373,N_26695,N_26601);
nor U32374 (N_32374,N_25043,N_25258);
and U32375 (N_32375,N_27307,N_27965);
nor U32376 (N_32376,N_26150,N_29750);
or U32377 (N_32377,N_29111,N_29838);
nor U32378 (N_32378,N_25183,N_25023);
nor U32379 (N_32379,N_29730,N_25444);
and U32380 (N_32380,N_29020,N_26229);
nand U32381 (N_32381,N_29315,N_29626);
nand U32382 (N_32382,N_29138,N_27452);
nand U32383 (N_32383,N_29793,N_26070);
nor U32384 (N_32384,N_25786,N_29160);
xnor U32385 (N_32385,N_28398,N_28585);
nor U32386 (N_32386,N_27778,N_26500);
or U32387 (N_32387,N_28527,N_27866);
nand U32388 (N_32388,N_25110,N_27228);
nor U32389 (N_32389,N_29360,N_26573);
nor U32390 (N_32390,N_26553,N_28641);
xor U32391 (N_32391,N_26798,N_28295);
nand U32392 (N_32392,N_26564,N_29515);
nor U32393 (N_32393,N_28513,N_26675);
and U32394 (N_32394,N_27758,N_29083);
and U32395 (N_32395,N_27074,N_27202);
xor U32396 (N_32396,N_28053,N_29947);
nand U32397 (N_32397,N_29556,N_28572);
and U32398 (N_32398,N_27635,N_29096);
nor U32399 (N_32399,N_25544,N_29646);
or U32400 (N_32400,N_26772,N_27161);
nand U32401 (N_32401,N_26367,N_26381);
nand U32402 (N_32402,N_29368,N_28029);
or U32403 (N_32403,N_26823,N_26085);
nor U32404 (N_32404,N_26951,N_28761);
nor U32405 (N_32405,N_28179,N_28274);
xnor U32406 (N_32406,N_29967,N_29765);
or U32407 (N_32407,N_28060,N_28752);
nor U32408 (N_32408,N_27553,N_29041);
nand U32409 (N_32409,N_25293,N_25733);
or U32410 (N_32410,N_26845,N_26682);
or U32411 (N_32411,N_25930,N_29706);
or U32412 (N_32412,N_25339,N_29238);
or U32413 (N_32413,N_25469,N_25174);
or U32414 (N_32414,N_25914,N_27002);
nor U32415 (N_32415,N_25207,N_28162);
nor U32416 (N_32416,N_28202,N_25641);
nand U32417 (N_32417,N_26692,N_26824);
nor U32418 (N_32418,N_29700,N_25600);
or U32419 (N_32419,N_28962,N_27114);
nor U32420 (N_32420,N_25432,N_25518);
or U32421 (N_32421,N_27806,N_27469);
and U32422 (N_32422,N_27880,N_26370);
xnor U32423 (N_32423,N_28780,N_26484);
or U32424 (N_32424,N_25540,N_29468);
or U32425 (N_32425,N_28061,N_26795);
or U32426 (N_32426,N_26304,N_25114);
xnor U32427 (N_32427,N_29836,N_25976);
xnor U32428 (N_32428,N_27291,N_27935);
or U32429 (N_32429,N_27971,N_27392);
xor U32430 (N_32430,N_26213,N_25586);
nand U32431 (N_32431,N_26867,N_28816);
or U32432 (N_32432,N_29526,N_25483);
and U32433 (N_32433,N_26317,N_25312);
nand U32434 (N_32434,N_25675,N_29086);
nand U32435 (N_32435,N_27711,N_27177);
xor U32436 (N_32436,N_26421,N_29924);
nand U32437 (N_32437,N_29167,N_25566);
or U32438 (N_32438,N_27905,N_27909);
or U32439 (N_32439,N_26634,N_27975);
nand U32440 (N_32440,N_28560,N_27992);
or U32441 (N_32441,N_27829,N_26519);
and U32442 (N_32442,N_28637,N_29642);
nand U32443 (N_32443,N_26257,N_27072);
and U32444 (N_32444,N_27101,N_26446);
nor U32445 (N_32445,N_26496,N_28436);
nand U32446 (N_32446,N_25949,N_27683);
nand U32447 (N_32447,N_29158,N_27027);
xnor U32448 (N_32448,N_29896,N_26189);
nand U32449 (N_32449,N_29990,N_26837);
nand U32450 (N_32450,N_26193,N_27653);
nand U32451 (N_32451,N_27059,N_27418);
nand U32452 (N_32452,N_25934,N_27943);
nand U32453 (N_32453,N_25975,N_27596);
nand U32454 (N_32454,N_26671,N_27222);
and U32455 (N_32455,N_28434,N_27985);
nand U32456 (N_32456,N_27509,N_26877);
and U32457 (N_32457,N_28198,N_29199);
and U32458 (N_32458,N_27193,N_26418);
xnor U32459 (N_32459,N_28706,N_26697);
or U32460 (N_32460,N_26779,N_29723);
nor U32461 (N_32461,N_29882,N_26454);
or U32462 (N_32462,N_27646,N_29190);
nor U32463 (N_32463,N_28014,N_29387);
nor U32464 (N_32464,N_29890,N_25323);
nand U32465 (N_32465,N_26644,N_25513);
nor U32466 (N_32466,N_27792,N_26414);
nor U32467 (N_32467,N_29375,N_26874);
or U32468 (N_32468,N_25736,N_27130);
nor U32469 (N_32469,N_26499,N_25446);
nor U32470 (N_32470,N_28267,N_28118);
xnor U32471 (N_32471,N_25212,N_28252);
xor U32472 (N_32472,N_29926,N_28624);
or U32473 (N_32473,N_28414,N_28621);
or U32474 (N_32474,N_26588,N_26137);
and U32475 (N_32475,N_28926,N_27396);
or U32476 (N_32476,N_27430,N_27137);
and U32477 (N_32477,N_26238,N_29865);
or U32478 (N_32478,N_29272,N_27141);
nand U32479 (N_32479,N_28771,N_27429);
nor U32480 (N_32480,N_28134,N_26687);
or U32481 (N_32481,N_25672,N_29408);
and U32482 (N_32482,N_26283,N_25473);
or U32483 (N_32483,N_29092,N_27558);
and U32484 (N_32484,N_28874,N_25900);
and U32485 (N_32485,N_28864,N_26003);
nor U32486 (N_32486,N_26034,N_25601);
nor U32487 (N_32487,N_29518,N_28302);
nor U32488 (N_32488,N_29397,N_28083);
or U32489 (N_32489,N_28774,N_27329);
xor U32490 (N_32490,N_29090,N_27136);
or U32491 (N_32491,N_29021,N_26780);
and U32492 (N_32492,N_27807,N_29502);
or U32493 (N_32493,N_25486,N_26017);
nor U32494 (N_32494,N_28730,N_29488);
and U32495 (N_32495,N_29118,N_26206);
nor U32496 (N_32496,N_26855,N_28189);
nor U32497 (N_32497,N_27574,N_29470);
nand U32498 (N_32498,N_27015,N_25547);
or U32499 (N_32499,N_28845,N_28565);
nand U32500 (N_32500,N_25112,N_27978);
nand U32501 (N_32501,N_27932,N_26753);
and U32502 (N_32502,N_27850,N_26471);
xnor U32503 (N_32503,N_28543,N_26037);
and U32504 (N_32504,N_28840,N_29037);
or U32505 (N_32505,N_27547,N_27115);
or U32506 (N_32506,N_28617,N_26111);
or U32507 (N_32507,N_28782,N_29592);
or U32508 (N_32508,N_27095,N_27433);
or U32509 (N_32509,N_25587,N_28832);
or U32510 (N_32510,N_28151,N_27154);
nand U32511 (N_32511,N_29701,N_29473);
nor U32512 (N_32512,N_27101,N_26748);
and U32513 (N_32513,N_26714,N_29778);
nand U32514 (N_32514,N_25392,N_26986);
nor U32515 (N_32515,N_26499,N_27725);
nor U32516 (N_32516,N_27408,N_26007);
nand U32517 (N_32517,N_27811,N_26750);
nor U32518 (N_32518,N_28341,N_28192);
nand U32519 (N_32519,N_25892,N_25849);
nand U32520 (N_32520,N_29235,N_26715);
nand U32521 (N_32521,N_25230,N_26579);
xnor U32522 (N_32522,N_29525,N_26986);
or U32523 (N_32523,N_28133,N_27770);
or U32524 (N_32524,N_27064,N_25297);
and U32525 (N_32525,N_25544,N_25555);
nand U32526 (N_32526,N_26129,N_25283);
xor U32527 (N_32527,N_25314,N_28739);
nand U32528 (N_32528,N_27871,N_27651);
xor U32529 (N_32529,N_26514,N_25235);
and U32530 (N_32530,N_27692,N_28802);
nand U32531 (N_32531,N_25046,N_28034);
nor U32532 (N_32532,N_27657,N_27521);
nor U32533 (N_32533,N_27775,N_28621);
nor U32534 (N_32534,N_26505,N_28909);
nand U32535 (N_32535,N_28753,N_25961);
and U32536 (N_32536,N_29112,N_28428);
and U32537 (N_32537,N_27735,N_26081);
nor U32538 (N_32538,N_28310,N_29594);
and U32539 (N_32539,N_26626,N_25341);
or U32540 (N_32540,N_27672,N_27659);
and U32541 (N_32541,N_29501,N_27449);
or U32542 (N_32542,N_29799,N_27766);
xnor U32543 (N_32543,N_28990,N_28571);
nor U32544 (N_32544,N_29614,N_27261);
and U32545 (N_32545,N_28130,N_28778);
or U32546 (N_32546,N_29166,N_27675);
nand U32547 (N_32547,N_25044,N_27095);
and U32548 (N_32548,N_25547,N_25360);
and U32549 (N_32549,N_29018,N_27075);
and U32550 (N_32550,N_26175,N_29371);
nand U32551 (N_32551,N_27034,N_26827);
xor U32552 (N_32552,N_29510,N_29375);
nor U32553 (N_32553,N_29250,N_29762);
nor U32554 (N_32554,N_26828,N_28142);
xnor U32555 (N_32555,N_25549,N_25942);
and U32556 (N_32556,N_29566,N_28595);
nor U32557 (N_32557,N_26270,N_28344);
nor U32558 (N_32558,N_26758,N_28854);
nor U32559 (N_32559,N_26016,N_27748);
xnor U32560 (N_32560,N_29335,N_25648);
xor U32561 (N_32561,N_28869,N_25316);
or U32562 (N_32562,N_29263,N_27109);
and U32563 (N_32563,N_25034,N_25173);
or U32564 (N_32564,N_27971,N_28225);
or U32565 (N_32565,N_28128,N_28367);
or U32566 (N_32566,N_26449,N_28333);
and U32567 (N_32567,N_27537,N_29033);
or U32568 (N_32568,N_25475,N_25635);
xnor U32569 (N_32569,N_28424,N_25216);
xnor U32570 (N_32570,N_25403,N_28553);
and U32571 (N_32571,N_29089,N_29583);
nor U32572 (N_32572,N_29785,N_26854);
and U32573 (N_32573,N_26474,N_26244);
nor U32574 (N_32574,N_26890,N_28795);
and U32575 (N_32575,N_27080,N_25607);
and U32576 (N_32576,N_25872,N_27525);
nand U32577 (N_32577,N_29108,N_26630);
and U32578 (N_32578,N_25726,N_27730);
or U32579 (N_32579,N_28883,N_27568);
nor U32580 (N_32580,N_27726,N_25839);
nand U32581 (N_32581,N_29413,N_29529);
xor U32582 (N_32582,N_28719,N_29855);
nor U32583 (N_32583,N_25306,N_26075);
and U32584 (N_32584,N_27754,N_29372);
and U32585 (N_32585,N_29478,N_28908);
or U32586 (N_32586,N_29720,N_26898);
and U32587 (N_32587,N_27520,N_26093);
or U32588 (N_32588,N_29944,N_26006);
and U32589 (N_32589,N_29968,N_25936);
or U32590 (N_32590,N_27194,N_26648);
nor U32591 (N_32591,N_27607,N_25629);
nand U32592 (N_32592,N_28664,N_25253);
nand U32593 (N_32593,N_25477,N_26000);
nor U32594 (N_32594,N_26080,N_29465);
or U32595 (N_32595,N_29071,N_25178);
or U32596 (N_32596,N_27124,N_27015);
and U32597 (N_32597,N_26467,N_28603);
or U32598 (N_32598,N_28037,N_27004);
xor U32599 (N_32599,N_26810,N_28651);
xnor U32600 (N_32600,N_26123,N_25325);
nand U32601 (N_32601,N_29830,N_25647);
or U32602 (N_32602,N_29264,N_25355);
xnor U32603 (N_32603,N_25052,N_29303);
xor U32604 (N_32604,N_28929,N_29699);
nor U32605 (N_32605,N_28506,N_28096);
nor U32606 (N_32606,N_29448,N_26374);
and U32607 (N_32607,N_26959,N_29202);
xnor U32608 (N_32608,N_26333,N_26213);
or U32609 (N_32609,N_28255,N_27926);
or U32610 (N_32610,N_29057,N_27569);
nor U32611 (N_32611,N_29050,N_25423);
nor U32612 (N_32612,N_26818,N_28810);
or U32613 (N_32613,N_28030,N_28736);
or U32614 (N_32614,N_29218,N_29735);
xnor U32615 (N_32615,N_27882,N_27947);
nor U32616 (N_32616,N_29996,N_25064);
nand U32617 (N_32617,N_25681,N_26675);
and U32618 (N_32618,N_29640,N_29834);
or U32619 (N_32619,N_28006,N_26851);
nand U32620 (N_32620,N_28727,N_26729);
and U32621 (N_32621,N_28689,N_27113);
or U32622 (N_32622,N_28603,N_27577);
and U32623 (N_32623,N_27497,N_28780);
or U32624 (N_32624,N_29265,N_28513);
nand U32625 (N_32625,N_28490,N_26755);
or U32626 (N_32626,N_29269,N_29148);
or U32627 (N_32627,N_27602,N_25514);
and U32628 (N_32628,N_29715,N_27626);
and U32629 (N_32629,N_26369,N_27372);
and U32630 (N_32630,N_27123,N_27388);
and U32631 (N_32631,N_27568,N_25543);
or U32632 (N_32632,N_27338,N_28446);
and U32633 (N_32633,N_28581,N_25324);
nand U32634 (N_32634,N_29098,N_28849);
and U32635 (N_32635,N_29826,N_26358);
and U32636 (N_32636,N_25176,N_25033);
or U32637 (N_32637,N_29288,N_27637);
nand U32638 (N_32638,N_25181,N_29317);
and U32639 (N_32639,N_28093,N_25550);
or U32640 (N_32640,N_25741,N_26883);
or U32641 (N_32641,N_26356,N_27021);
nand U32642 (N_32642,N_27928,N_27848);
or U32643 (N_32643,N_26995,N_29463);
nand U32644 (N_32644,N_29976,N_27513);
nand U32645 (N_32645,N_27661,N_25709);
nor U32646 (N_32646,N_25876,N_29833);
nor U32647 (N_32647,N_25781,N_25691);
xnor U32648 (N_32648,N_26783,N_27318);
and U32649 (N_32649,N_29611,N_28298);
nor U32650 (N_32650,N_26446,N_25231);
and U32651 (N_32651,N_25264,N_25407);
or U32652 (N_32652,N_28733,N_28977);
xor U32653 (N_32653,N_27546,N_25018);
nor U32654 (N_32654,N_28408,N_28730);
and U32655 (N_32655,N_26028,N_26474);
and U32656 (N_32656,N_29965,N_26558);
or U32657 (N_32657,N_27773,N_26515);
nand U32658 (N_32658,N_28880,N_29014);
nand U32659 (N_32659,N_25565,N_25984);
nor U32660 (N_32660,N_28267,N_26868);
nor U32661 (N_32661,N_25477,N_29859);
and U32662 (N_32662,N_29358,N_28577);
and U32663 (N_32663,N_28761,N_26857);
xnor U32664 (N_32664,N_26703,N_26100);
nor U32665 (N_32665,N_27586,N_29038);
and U32666 (N_32666,N_28547,N_27119);
and U32667 (N_32667,N_26841,N_29897);
or U32668 (N_32668,N_28059,N_25919);
nand U32669 (N_32669,N_28337,N_25539);
nor U32670 (N_32670,N_29894,N_26818);
nor U32671 (N_32671,N_26085,N_27924);
and U32672 (N_32672,N_28097,N_29616);
or U32673 (N_32673,N_27798,N_29173);
or U32674 (N_32674,N_28504,N_29250);
nand U32675 (N_32675,N_29715,N_27494);
or U32676 (N_32676,N_26725,N_29931);
nand U32677 (N_32677,N_28793,N_28427);
xnor U32678 (N_32678,N_26217,N_25247);
nor U32679 (N_32679,N_25226,N_29861);
or U32680 (N_32680,N_27574,N_26856);
and U32681 (N_32681,N_25932,N_26030);
or U32682 (N_32682,N_27853,N_25636);
nand U32683 (N_32683,N_28442,N_26006);
and U32684 (N_32684,N_29455,N_28040);
nand U32685 (N_32685,N_26066,N_29268);
nor U32686 (N_32686,N_27792,N_28894);
and U32687 (N_32687,N_28960,N_29341);
and U32688 (N_32688,N_25484,N_27436);
and U32689 (N_32689,N_27324,N_25427);
nand U32690 (N_32690,N_25662,N_28350);
xnor U32691 (N_32691,N_26994,N_25781);
nor U32692 (N_32692,N_25692,N_29815);
nand U32693 (N_32693,N_29560,N_25134);
nor U32694 (N_32694,N_25716,N_25429);
nor U32695 (N_32695,N_25184,N_26824);
nand U32696 (N_32696,N_26472,N_29723);
xnor U32697 (N_32697,N_27795,N_28042);
nor U32698 (N_32698,N_27798,N_26080);
nor U32699 (N_32699,N_28945,N_28655);
nand U32700 (N_32700,N_27558,N_25643);
xor U32701 (N_32701,N_29095,N_29677);
nand U32702 (N_32702,N_27370,N_28059);
nand U32703 (N_32703,N_25957,N_25792);
nor U32704 (N_32704,N_29903,N_29139);
nor U32705 (N_32705,N_27188,N_25640);
nand U32706 (N_32706,N_26379,N_25553);
and U32707 (N_32707,N_26772,N_25918);
or U32708 (N_32708,N_26663,N_26599);
or U32709 (N_32709,N_29084,N_27094);
or U32710 (N_32710,N_26984,N_28020);
or U32711 (N_32711,N_26639,N_26038);
and U32712 (N_32712,N_26915,N_27641);
nor U32713 (N_32713,N_26478,N_27628);
nor U32714 (N_32714,N_28708,N_28401);
nand U32715 (N_32715,N_28527,N_26579);
nand U32716 (N_32716,N_27287,N_25871);
nand U32717 (N_32717,N_28430,N_25667);
and U32718 (N_32718,N_26516,N_26235);
and U32719 (N_32719,N_25697,N_27406);
nand U32720 (N_32720,N_29205,N_25330);
or U32721 (N_32721,N_25172,N_26824);
nor U32722 (N_32722,N_25975,N_27438);
nor U32723 (N_32723,N_26591,N_25276);
nand U32724 (N_32724,N_29014,N_25015);
and U32725 (N_32725,N_25351,N_28937);
nor U32726 (N_32726,N_27165,N_26118);
xnor U32727 (N_32727,N_27135,N_25562);
or U32728 (N_32728,N_27154,N_28681);
xnor U32729 (N_32729,N_29644,N_29195);
or U32730 (N_32730,N_29232,N_27111);
nand U32731 (N_32731,N_27146,N_27924);
and U32732 (N_32732,N_29646,N_26766);
nor U32733 (N_32733,N_29467,N_29709);
nor U32734 (N_32734,N_26938,N_26911);
nor U32735 (N_32735,N_27784,N_25619);
or U32736 (N_32736,N_27568,N_28952);
nand U32737 (N_32737,N_25881,N_28578);
nor U32738 (N_32738,N_27768,N_27823);
nand U32739 (N_32739,N_26699,N_25915);
and U32740 (N_32740,N_26414,N_27913);
or U32741 (N_32741,N_29404,N_28307);
nand U32742 (N_32742,N_25172,N_25698);
nor U32743 (N_32743,N_29374,N_25226);
or U32744 (N_32744,N_28428,N_28558);
or U32745 (N_32745,N_29076,N_25403);
nand U32746 (N_32746,N_25199,N_29546);
or U32747 (N_32747,N_27410,N_25207);
nand U32748 (N_32748,N_26946,N_29099);
and U32749 (N_32749,N_25773,N_25410);
or U32750 (N_32750,N_26247,N_28007);
and U32751 (N_32751,N_29501,N_27323);
nor U32752 (N_32752,N_28243,N_27965);
nand U32753 (N_32753,N_26488,N_28319);
nand U32754 (N_32754,N_26668,N_26432);
or U32755 (N_32755,N_29794,N_28761);
and U32756 (N_32756,N_27066,N_29185);
or U32757 (N_32757,N_27697,N_29677);
nor U32758 (N_32758,N_27010,N_28932);
xor U32759 (N_32759,N_27306,N_29636);
nor U32760 (N_32760,N_28867,N_27498);
and U32761 (N_32761,N_27921,N_26820);
or U32762 (N_32762,N_28444,N_25733);
nor U32763 (N_32763,N_28047,N_26292);
nor U32764 (N_32764,N_27468,N_26855);
or U32765 (N_32765,N_26861,N_29712);
nand U32766 (N_32766,N_27241,N_28414);
or U32767 (N_32767,N_28654,N_27124);
and U32768 (N_32768,N_28806,N_27020);
or U32769 (N_32769,N_28508,N_26015);
nand U32770 (N_32770,N_28020,N_26380);
or U32771 (N_32771,N_26181,N_29077);
and U32772 (N_32772,N_25808,N_27717);
nor U32773 (N_32773,N_28095,N_29914);
nand U32774 (N_32774,N_27458,N_26301);
nand U32775 (N_32775,N_25704,N_28068);
nand U32776 (N_32776,N_25188,N_28274);
nor U32777 (N_32777,N_28476,N_28913);
and U32778 (N_32778,N_28354,N_25437);
nor U32779 (N_32779,N_26574,N_28769);
and U32780 (N_32780,N_26126,N_28482);
nand U32781 (N_32781,N_25561,N_26490);
xnor U32782 (N_32782,N_27764,N_26144);
nor U32783 (N_32783,N_27105,N_26031);
nand U32784 (N_32784,N_29576,N_25678);
and U32785 (N_32785,N_25505,N_29252);
and U32786 (N_32786,N_25685,N_28260);
and U32787 (N_32787,N_28435,N_28196);
nor U32788 (N_32788,N_25937,N_26944);
nor U32789 (N_32789,N_27921,N_25553);
nor U32790 (N_32790,N_25994,N_26752);
nand U32791 (N_32791,N_29071,N_29683);
nor U32792 (N_32792,N_28107,N_29553);
nand U32793 (N_32793,N_28118,N_27571);
and U32794 (N_32794,N_25204,N_26594);
nand U32795 (N_32795,N_27468,N_29727);
xnor U32796 (N_32796,N_25929,N_27204);
or U32797 (N_32797,N_27861,N_26853);
or U32798 (N_32798,N_27595,N_26033);
nor U32799 (N_32799,N_25284,N_26737);
nor U32800 (N_32800,N_29427,N_29346);
xnor U32801 (N_32801,N_26544,N_25880);
nor U32802 (N_32802,N_28736,N_29443);
nand U32803 (N_32803,N_26773,N_28081);
nand U32804 (N_32804,N_29694,N_27456);
nand U32805 (N_32805,N_27551,N_29031);
nand U32806 (N_32806,N_27705,N_25269);
nand U32807 (N_32807,N_27176,N_28444);
nand U32808 (N_32808,N_27957,N_29889);
and U32809 (N_32809,N_28778,N_26371);
nand U32810 (N_32810,N_25808,N_27342);
and U32811 (N_32811,N_27314,N_26579);
and U32812 (N_32812,N_27439,N_26339);
nand U32813 (N_32813,N_25988,N_29008);
or U32814 (N_32814,N_29093,N_27915);
and U32815 (N_32815,N_27301,N_29446);
and U32816 (N_32816,N_25589,N_28535);
nand U32817 (N_32817,N_26870,N_28279);
and U32818 (N_32818,N_26980,N_27424);
nor U32819 (N_32819,N_28404,N_28394);
nor U32820 (N_32820,N_29783,N_27710);
or U32821 (N_32821,N_27034,N_28247);
or U32822 (N_32822,N_25970,N_29731);
nand U32823 (N_32823,N_28141,N_26664);
nand U32824 (N_32824,N_29474,N_26368);
or U32825 (N_32825,N_25887,N_27286);
nand U32826 (N_32826,N_27977,N_28781);
nor U32827 (N_32827,N_26211,N_26662);
or U32828 (N_32828,N_25772,N_28671);
or U32829 (N_32829,N_26142,N_28349);
nor U32830 (N_32830,N_26901,N_26919);
nand U32831 (N_32831,N_25744,N_28740);
or U32832 (N_32832,N_28173,N_29584);
and U32833 (N_32833,N_26444,N_27646);
nor U32834 (N_32834,N_27883,N_29575);
or U32835 (N_32835,N_25375,N_28363);
or U32836 (N_32836,N_26929,N_26191);
and U32837 (N_32837,N_27090,N_25679);
and U32838 (N_32838,N_26330,N_25409);
nand U32839 (N_32839,N_29765,N_26885);
nand U32840 (N_32840,N_27439,N_28720);
nor U32841 (N_32841,N_27156,N_27119);
nand U32842 (N_32842,N_28798,N_27387);
or U32843 (N_32843,N_26768,N_28969);
and U32844 (N_32844,N_27697,N_25020);
nor U32845 (N_32845,N_29880,N_29106);
and U32846 (N_32846,N_27476,N_29255);
nand U32847 (N_32847,N_29567,N_25589);
nor U32848 (N_32848,N_28749,N_26355);
nand U32849 (N_32849,N_27294,N_29656);
or U32850 (N_32850,N_28489,N_28824);
nor U32851 (N_32851,N_29907,N_29563);
nor U32852 (N_32852,N_26209,N_27343);
nand U32853 (N_32853,N_29575,N_27135);
or U32854 (N_32854,N_27168,N_26571);
nand U32855 (N_32855,N_25011,N_29951);
nand U32856 (N_32856,N_29550,N_29179);
xor U32857 (N_32857,N_28479,N_25001);
and U32858 (N_32858,N_25819,N_29988);
nor U32859 (N_32859,N_28289,N_29223);
nand U32860 (N_32860,N_25308,N_27107);
nor U32861 (N_32861,N_28422,N_25833);
xor U32862 (N_32862,N_27212,N_29635);
nand U32863 (N_32863,N_28912,N_25191);
xnor U32864 (N_32864,N_29073,N_27400);
nor U32865 (N_32865,N_29879,N_28233);
and U32866 (N_32866,N_27784,N_27148);
nor U32867 (N_32867,N_27206,N_28082);
xor U32868 (N_32868,N_29530,N_27393);
or U32869 (N_32869,N_26752,N_27283);
and U32870 (N_32870,N_25548,N_26931);
and U32871 (N_32871,N_25505,N_26399);
nor U32872 (N_32872,N_25429,N_29442);
nor U32873 (N_32873,N_28246,N_29901);
nor U32874 (N_32874,N_29923,N_26804);
or U32875 (N_32875,N_27499,N_29699);
or U32876 (N_32876,N_27912,N_27197);
nand U32877 (N_32877,N_28326,N_28756);
nand U32878 (N_32878,N_25831,N_26220);
and U32879 (N_32879,N_28607,N_25172);
and U32880 (N_32880,N_26417,N_29420);
nand U32881 (N_32881,N_26451,N_29215);
nor U32882 (N_32882,N_28941,N_29453);
and U32883 (N_32883,N_27565,N_26604);
or U32884 (N_32884,N_27700,N_27648);
nand U32885 (N_32885,N_27831,N_28179);
or U32886 (N_32886,N_26769,N_27126);
xor U32887 (N_32887,N_28937,N_28991);
or U32888 (N_32888,N_25730,N_29079);
nor U32889 (N_32889,N_28565,N_25963);
nand U32890 (N_32890,N_25919,N_25368);
or U32891 (N_32891,N_25469,N_29960);
xnor U32892 (N_32892,N_27520,N_26950);
and U32893 (N_32893,N_28582,N_27814);
and U32894 (N_32894,N_27882,N_26594);
nor U32895 (N_32895,N_27273,N_25690);
and U32896 (N_32896,N_26028,N_28693);
xnor U32897 (N_32897,N_27443,N_29868);
or U32898 (N_32898,N_25638,N_28303);
or U32899 (N_32899,N_28458,N_28530);
and U32900 (N_32900,N_27105,N_29746);
and U32901 (N_32901,N_25956,N_26986);
nand U32902 (N_32902,N_25698,N_27058);
nand U32903 (N_32903,N_29395,N_26242);
or U32904 (N_32904,N_25823,N_27194);
nor U32905 (N_32905,N_25970,N_28923);
xnor U32906 (N_32906,N_29020,N_29791);
nand U32907 (N_32907,N_28518,N_27668);
or U32908 (N_32908,N_25825,N_26731);
or U32909 (N_32909,N_29080,N_26720);
or U32910 (N_32910,N_27933,N_25738);
and U32911 (N_32911,N_25388,N_27989);
and U32912 (N_32912,N_28565,N_26448);
xnor U32913 (N_32913,N_29391,N_25917);
nand U32914 (N_32914,N_27686,N_28634);
and U32915 (N_32915,N_28173,N_26286);
or U32916 (N_32916,N_26035,N_28285);
xnor U32917 (N_32917,N_29240,N_28238);
and U32918 (N_32918,N_28308,N_27536);
and U32919 (N_32919,N_29016,N_28253);
nand U32920 (N_32920,N_28019,N_27568);
and U32921 (N_32921,N_25269,N_29017);
and U32922 (N_32922,N_25899,N_27192);
nand U32923 (N_32923,N_27340,N_29110);
nor U32924 (N_32924,N_25667,N_26590);
and U32925 (N_32925,N_25127,N_25188);
nand U32926 (N_32926,N_26663,N_26662);
nand U32927 (N_32927,N_27695,N_27949);
or U32928 (N_32928,N_28988,N_29509);
or U32929 (N_32929,N_29984,N_29608);
nor U32930 (N_32930,N_26463,N_29683);
or U32931 (N_32931,N_26973,N_26013);
and U32932 (N_32932,N_25773,N_25624);
or U32933 (N_32933,N_26178,N_27654);
xnor U32934 (N_32934,N_27180,N_28122);
nand U32935 (N_32935,N_27884,N_29058);
and U32936 (N_32936,N_27353,N_25003);
xnor U32937 (N_32937,N_29411,N_25310);
xor U32938 (N_32938,N_29111,N_28190);
nor U32939 (N_32939,N_25268,N_25916);
or U32940 (N_32940,N_25589,N_25007);
xnor U32941 (N_32941,N_28902,N_25382);
nor U32942 (N_32942,N_28718,N_26663);
nor U32943 (N_32943,N_26404,N_28031);
and U32944 (N_32944,N_27816,N_27783);
and U32945 (N_32945,N_29009,N_26987);
and U32946 (N_32946,N_28209,N_26713);
and U32947 (N_32947,N_25549,N_27457);
xnor U32948 (N_32948,N_26986,N_29353);
and U32949 (N_32949,N_27796,N_25881);
nand U32950 (N_32950,N_26733,N_25879);
xor U32951 (N_32951,N_27673,N_26780);
nor U32952 (N_32952,N_29965,N_27185);
nand U32953 (N_32953,N_29055,N_26698);
nand U32954 (N_32954,N_25390,N_27957);
nand U32955 (N_32955,N_25638,N_27518);
and U32956 (N_32956,N_27913,N_25608);
nand U32957 (N_32957,N_26307,N_27340);
nor U32958 (N_32958,N_29148,N_25521);
nor U32959 (N_32959,N_29570,N_27045);
xnor U32960 (N_32960,N_26418,N_25343);
nand U32961 (N_32961,N_25037,N_29346);
and U32962 (N_32962,N_25252,N_28701);
xor U32963 (N_32963,N_27725,N_27216);
and U32964 (N_32964,N_25931,N_26108);
xnor U32965 (N_32965,N_27429,N_29409);
xnor U32966 (N_32966,N_25354,N_29516);
nor U32967 (N_32967,N_27418,N_29104);
nor U32968 (N_32968,N_27579,N_27306);
nand U32969 (N_32969,N_27043,N_29490);
nand U32970 (N_32970,N_27058,N_28635);
and U32971 (N_32971,N_26934,N_28895);
or U32972 (N_32972,N_28745,N_28599);
nor U32973 (N_32973,N_28679,N_28308);
and U32974 (N_32974,N_25762,N_26570);
nand U32975 (N_32975,N_27739,N_26019);
and U32976 (N_32976,N_29219,N_26707);
nand U32977 (N_32977,N_27368,N_29965);
and U32978 (N_32978,N_26447,N_25902);
nor U32979 (N_32979,N_28560,N_25108);
nand U32980 (N_32980,N_25072,N_29967);
or U32981 (N_32981,N_27102,N_25306);
or U32982 (N_32982,N_29066,N_28409);
and U32983 (N_32983,N_25810,N_29376);
and U32984 (N_32984,N_28499,N_28571);
nor U32985 (N_32985,N_28577,N_28029);
nor U32986 (N_32986,N_26337,N_27002);
nor U32987 (N_32987,N_29651,N_25405);
and U32988 (N_32988,N_28485,N_29097);
xor U32989 (N_32989,N_25880,N_27816);
xor U32990 (N_32990,N_26227,N_25956);
and U32991 (N_32991,N_29974,N_28546);
nor U32992 (N_32992,N_29154,N_27441);
nand U32993 (N_32993,N_29290,N_26094);
nand U32994 (N_32994,N_29414,N_27066);
nand U32995 (N_32995,N_25312,N_29262);
and U32996 (N_32996,N_29136,N_28980);
nand U32997 (N_32997,N_29352,N_28758);
xor U32998 (N_32998,N_29743,N_27346);
nand U32999 (N_32999,N_27529,N_28663);
or U33000 (N_33000,N_29010,N_26398);
or U33001 (N_33001,N_27765,N_29354);
or U33002 (N_33002,N_26783,N_26647);
nor U33003 (N_33003,N_29520,N_25871);
nor U33004 (N_33004,N_27797,N_27244);
nand U33005 (N_33005,N_28336,N_27576);
xor U33006 (N_33006,N_29081,N_28376);
and U33007 (N_33007,N_27648,N_28044);
and U33008 (N_33008,N_29386,N_29153);
or U33009 (N_33009,N_29885,N_27273);
nor U33010 (N_33010,N_27934,N_29831);
nor U33011 (N_33011,N_29148,N_25471);
xnor U33012 (N_33012,N_25968,N_25073);
xnor U33013 (N_33013,N_25146,N_28806);
xnor U33014 (N_33014,N_28543,N_26670);
nor U33015 (N_33015,N_27994,N_26361);
and U33016 (N_33016,N_26637,N_26040);
nor U33017 (N_33017,N_29240,N_26521);
nand U33018 (N_33018,N_28668,N_26035);
nor U33019 (N_33019,N_25442,N_27885);
or U33020 (N_33020,N_27710,N_26069);
nor U33021 (N_33021,N_27630,N_28187);
or U33022 (N_33022,N_27112,N_25958);
nor U33023 (N_33023,N_29685,N_29250);
xnor U33024 (N_33024,N_27602,N_26139);
and U33025 (N_33025,N_29424,N_29809);
xnor U33026 (N_33026,N_26285,N_26200);
or U33027 (N_33027,N_28952,N_29308);
or U33028 (N_33028,N_25944,N_27811);
nor U33029 (N_33029,N_28949,N_27017);
and U33030 (N_33030,N_29448,N_27628);
xor U33031 (N_33031,N_29607,N_29304);
nor U33032 (N_33032,N_28697,N_25055);
or U33033 (N_33033,N_27044,N_25724);
nor U33034 (N_33034,N_27318,N_26400);
or U33035 (N_33035,N_28391,N_26268);
nand U33036 (N_33036,N_29273,N_26898);
or U33037 (N_33037,N_26761,N_26210);
nor U33038 (N_33038,N_27361,N_27618);
and U33039 (N_33039,N_26843,N_28473);
xnor U33040 (N_33040,N_26082,N_29129);
nor U33041 (N_33041,N_25305,N_26590);
and U33042 (N_33042,N_28263,N_25951);
and U33043 (N_33043,N_29046,N_26142);
or U33044 (N_33044,N_29675,N_25864);
nor U33045 (N_33045,N_25856,N_27658);
xnor U33046 (N_33046,N_28159,N_29594);
or U33047 (N_33047,N_26675,N_25429);
and U33048 (N_33048,N_26212,N_25820);
or U33049 (N_33049,N_27482,N_29812);
nor U33050 (N_33050,N_28884,N_26264);
or U33051 (N_33051,N_26410,N_27992);
and U33052 (N_33052,N_25363,N_27198);
nand U33053 (N_33053,N_27324,N_29961);
xor U33054 (N_33054,N_25706,N_26336);
and U33055 (N_33055,N_28890,N_25408);
or U33056 (N_33056,N_27294,N_29989);
or U33057 (N_33057,N_29810,N_28871);
or U33058 (N_33058,N_26812,N_29190);
and U33059 (N_33059,N_25655,N_28868);
or U33060 (N_33060,N_28527,N_26515);
or U33061 (N_33061,N_26580,N_28855);
or U33062 (N_33062,N_27127,N_26849);
nor U33063 (N_33063,N_27060,N_25233);
and U33064 (N_33064,N_29157,N_27113);
nor U33065 (N_33065,N_28657,N_27055);
or U33066 (N_33066,N_27025,N_27731);
nand U33067 (N_33067,N_26613,N_28095);
nand U33068 (N_33068,N_27098,N_25982);
or U33069 (N_33069,N_26712,N_29145);
nor U33070 (N_33070,N_27180,N_27602);
xnor U33071 (N_33071,N_28368,N_29133);
or U33072 (N_33072,N_29280,N_26089);
nand U33073 (N_33073,N_26555,N_27525);
and U33074 (N_33074,N_26203,N_28085);
nand U33075 (N_33075,N_26156,N_27791);
nand U33076 (N_33076,N_29998,N_29701);
or U33077 (N_33077,N_26449,N_27083);
xnor U33078 (N_33078,N_27067,N_28712);
nor U33079 (N_33079,N_28992,N_25312);
xor U33080 (N_33080,N_25672,N_26974);
nand U33081 (N_33081,N_28940,N_27289);
nor U33082 (N_33082,N_29587,N_25235);
nand U33083 (N_33083,N_25039,N_25395);
or U33084 (N_33084,N_25833,N_26234);
nor U33085 (N_33085,N_28789,N_27325);
xnor U33086 (N_33086,N_26030,N_26643);
nand U33087 (N_33087,N_25792,N_27799);
and U33088 (N_33088,N_26385,N_29056);
nand U33089 (N_33089,N_29505,N_25177);
nor U33090 (N_33090,N_29778,N_25913);
nor U33091 (N_33091,N_26382,N_26359);
or U33092 (N_33092,N_27523,N_25028);
nand U33093 (N_33093,N_29997,N_29710);
and U33094 (N_33094,N_29494,N_26096);
xnor U33095 (N_33095,N_29019,N_28840);
nor U33096 (N_33096,N_26129,N_25538);
and U33097 (N_33097,N_25037,N_29249);
nor U33098 (N_33098,N_25182,N_28815);
and U33099 (N_33099,N_27061,N_27743);
and U33100 (N_33100,N_27520,N_27296);
and U33101 (N_33101,N_28545,N_29993);
nand U33102 (N_33102,N_27724,N_26337);
and U33103 (N_33103,N_28835,N_29325);
xnor U33104 (N_33104,N_29778,N_26928);
and U33105 (N_33105,N_26686,N_26357);
nand U33106 (N_33106,N_25818,N_26185);
nand U33107 (N_33107,N_29982,N_25146);
or U33108 (N_33108,N_27848,N_25040);
and U33109 (N_33109,N_26954,N_27658);
nand U33110 (N_33110,N_26300,N_29899);
or U33111 (N_33111,N_29040,N_25410);
nand U33112 (N_33112,N_28788,N_28149);
nor U33113 (N_33113,N_26031,N_26863);
nor U33114 (N_33114,N_27942,N_25757);
nand U33115 (N_33115,N_28599,N_26002);
and U33116 (N_33116,N_29626,N_27122);
or U33117 (N_33117,N_26128,N_26699);
or U33118 (N_33118,N_29552,N_25469);
and U33119 (N_33119,N_29501,N_27943);
nor U33120 (N_33120,N_26048,N_29757);
nand U33121 (N_33121,N_29768,N_29679);
nor U33122 (N_33122,N_25998,N_29116);
or U33123 (N_33123,N_29127,N_25907);
xnor U33124 (N_33124,N_29744,N_26349);
nor U33125 (N_33125,N_28653,N_29046);
nor U33126 (N_33126,N_27702,N_25748);
nand U33127 (N_33127,N_26799,N_27014);
nand U33128 (N_33128,N_27579,N_25015);
nand U33129 (N_33129,N_25882,N_25740);
nand U33130 (N_33130,N_27676,N_25055);
and U33131 (N_33131,N_29533,N_26140);
nand U33132 (N_33132,N_27990,N_27579);
nor U33133 (N_33133,N_29287,N_26234);
nand U33134 (N_33134,N_29654,N_27613);
and U33135 (N_33135,N_25597,N_28228);
nand U33136 (N_33136,N_28466,N_27369);
nand U33137 (N_33137,N_29648,N_29179);
nand U33138 (N_33138,N_29940,N_27836);
nor U33139 (N_33139,N_26245,N_27961);
nor U33140 (N_33140,N_28721,N_27805);
nor U33141 (N_33141,N_29604,N_26961);
xor U33142 (N_33142,N_25576,N_27685);
nand U33143 (N_33143,N_26212,N_28140);
nor U33144 (N_33144,N_28614,N_27463);
nand U33145 (N_33145,N_28786,N_28337);
nand U33146 (N_33146,N_29182,N_27773);
nand U33147 (N_33147,N_29792,N_25467);
and U33148 (N_33148,N_25246,N_27428);
and U33149 (N_33149,N_29698,N_29452);
and U33150 (N_33150,N_26269,N_25009);
nand U33151 (N_33151,N_27077,N_25367);
nor U33152 (N_33152,N_28710,N_27190);
nand U33153 (N_33153,N_29042,N_27452);
or U33154 (N_33154,N_25564,N_25829);
xnor U33155 (N_33155,N_26678,N_28137);
nand U33156 (N_33156,N_25896,N_26179);
and U33157 (N_33157,N_29712,N_27251);
nor U33158 (N_33158,N_27645,N_28418);
or U33159 (N_33159,N_28911,N_29168);
or U33160 (N_33160,N_26514,N_27476);
nand U33161 (N_33161,N_27822,N_27151);
and U33162 (N_33162,N_26552,N_25993);
nor U33163 (N_33163,N_28714,N_29934);
or U33164 (N_33164,N_25761,N_29646);
or U33165 (N_33165,N_26376,N_26010);
or U33166 (N_33166,N_26699,N_25597);
nand U33167 (N_33167,N_27409,N_25313);
nor U33168 (N_33168,N_25819,N_25386);
and U33169 (N_33169,N_26638,N_26469);
or U33170 (N_33170,N_28885,N_25978);
and U33171 (N_33171,N_25709,N_28693);
nor U33172 (N_33172,N_27626,N_28422);
or U33173 (N_33173,N_26613,N_26072);
or U33174 (N_33174,N_29115,N_29015);
and U33175 (N_33175,N_25086,N_27253);
xor U33176 (N_33176,N_25172,N_29892);
xor U33177 (N_33177,N_29905,N_25761);
xnor U33178 (N_33178,N_28133,N_28754);
or U33179 (N_33179,N_28797,N_27996);
nor U33180 (N_33180,N_29317,N_26838);
nor U33181 (N_33181,N_26289,N_27357);
and U33182 (N_33182,N_25394,N_26975);
nand U33183 (N_33183,N_27577,N_28984);
xnor U33184 (N_33184,N_26420,N_27100);
and U33185 (N_33185,N_25608,N_28043);
nor U33186 (N_33186,N_26793,N_29252);
or U33187 (N_33187,N_26171,N_26808);
and U33188 (N_33188,N_26908,N_28106);
nor U33189 (N_33189,N_28428,N_28316);
and U33190 (N_33190,N_26418,N_25212);
xor U33191 (N_33191,N_26094,N_28304);
or U33192 (N_33192,N_26841,N_29689);
nand U33193 (N_33193,N_25088,N_27921);
and U33194 (N_33194,N_27856,N_27803);
nor U33195 (N_33195,N_29167,N_28280);
nor U33196 (N_33196,N_27290,N_29371);
or U33197 (N_33197,N_28129,N_28734);
or U33198 (N_33198,N_26767,N_27784);
and U33199 (N_33199,N_25357,N_27642);
and U33200 (N_33200,N_29977,N_29797);
xnor U33201 (N_33201,N_28945,N_26717);
or U33202 (N_33202,N_26798,N_29962);
or U33203 (N_33203,N_26206,N_26262);
or U33204 (N_33204,N_25485,N_25157);
and U33205 (N_33205,N_29878,N_27680);
and U33206 (N_33206,N_25207,N_29796);
nand U33207 (N_33207,N_25534,N_26208);
and U33208 (N_33208,N_26135,N_26065);
nor U33209 (N_33209,N_27663,N_28435);
and U33210 (N_33210,N_29781,N_27737);
and U33211 (N_33211,N_25093,N_29736);
xnor U33212 (N_33212,N_29514,N_25972);
nand U33213 (N_33213,N_26416,N_28353);
nor U33214 (N_33214,N_25981,N_26201);
and U33215 (N_33215,N_29887,N_25133);
nor U33216 (N_33216,N_29261,N_28347);
and U33217 (N_33217,N_29050,N_28641);
or U33218 (N_33218,N_29806,N_25312);
or U33219 (N_33219,N_27061,N_26895);
and U33220 (N_33220,N_28545,N_29697);
nor U33221 (N_33221,N_26952,N_28694);
xor U33222 (N_33222,N_27769,N_27043);
nor U33223 (N_33223,N_27785,N_28355);
or U33224 (N_33224,N_27409,N_28018);
or U33225 (N_33225,N_29321,N_25481);
nand U33226 (N_33226,N_25535,N_28986);
and U33227 (N_33227,N_25899,N_25264);
nand U33228 (N_33228,N_25419,N_28015);
nand U33229 (N_33229,N_27237,N_26414);
xor U33230 (N_33230,N_29285,N_27242);
or U33231 (N_33231,N_26450,N_28884);
xor U33232 (N_33232,N_26955,N_28138);
nand U33233 (N_33233,N_27607,N_25866);
and U33234 (N_33234,N_28118,N_25942);
and U33235 (N_33235,N_26742,N_28238);
nand U33236 (N_33236,N_25841,N_26198);
nand U33237 (N_33237,N_26265,N_28366);
or U33238 (N_33238,N_26499,N_28978);
nor U33239 (N_33239,N_29851,N_28710);
nand U33240 (N_33240,N_25310,N_25538);
or U33241 (N_33241,N_25530,N_28554);
or U33242 (N_33242,N_28604,N_27090);
or U33243 (N_33243,N_27122,N_28706);
or U33244 (N_33244,N_29176,N_26206);
nand U33245 (N_33245,N_28671,N_28448);
nand U33246 (N_33246,N_25828,N_28621);
or U33247 (N_33247,N_28516,N_29904);
nor U33248 (N_33248,N_29348,N_27288);
xnor U33249 (N_33249,N_26699,N_26710);
nand U33250 (N_33250,N_27466,N_25447);
and U33251 (N_33251,N_25976,N_26527);
nand U33252 (N_33252,N_27840,N_26014);
or U33253 (N_33253,N_29122,N_26009);
nor U33254 (N_33254,N_27121,N_25331);
or U33255 (N_33255,N_28350,N_27076);
nor U33256 (N_33256,N_26819,N_25429);
and U33257 (N_33257,N_26927,N_29099);
xor U33258 (N_33258,N_27912,N_29924);
nor U33259 (N_33259,N_28109,N_28943);
nand U33260 (N_33260,N_28165,N_27382);
and U33261 (N_33261,N_29844,N_25602);
and U33262 (N_33262,N_29430,N_28160);
and U33263 (N_33263,N_25623,N_28831);
nand U33264 (N_33264,N_25918,N_29393);
nand U33265 (N_33265,N_26739,N_29780);
xor U33266 (N_33266,N_26195,N_26424);
and U33267 (N_33267,N_25785,N_26695);
and U33268 (N_33268,N_26432,N_27692);
and U33269 (N_33269,N_26525,N_27606);
nor U33270 (N_33270,N_29982,N_26297);
nand U33271 (N_33271,N_25557,N_26403);
nand U33272 (N_33272,N_28018,N_29011);
and U33273 (N_33273,N_26023,N_27423);
nand U33274 (N_33274,N_26202,N_27219);
nor U33275 (N_33275,N_29099,N_27548);
and U33276 (N_33276,N_27992,N_29812);
nand U33277 (N_33277,N_29691,N_25711);
and U33278 (N_33278,N_27367,N_25075);
or U33279 (N_33279,N_29371,N_28557);
nand U33280 (N_33280,N_28687,N_28669);
or U33281 (N_33281,N_28206,N_25528);
nor U33282 (N_33282,N_26398,N_28062);
or U33283 (N_33283,N_28727,N_29763);
or U33284 (N_33284,N_25615,N_29969);
and U33285 (N_33285,N_26573,N_29707);
and U33286 (N_33286,N_25108,N_26121);
nor U33287 (N_33287,N_29761,N_29358);
and U33288 (N_33288,N_27675,N_28182);
or U33289 (N_33289,N_28159,N_28643);
nand U33290 (N_33290,N_26157,N_28777);
nor U33291 (N_33291,N_25164,N_27203);
nand U33292 (N_33292,N_27310,N_28716);
nand U33293 (N_33293,N_25638,N_29035);
or U33294 (N_33294,N_29872,N_25770);
nand U33295 (N_33295,N_27117,N_27610);
and U33296 (N_33296,N_25273,N_27963);
and U33297 (N_33297,N_25319,N_27278);
nand U33298 (N_33298,N_25786,N_29776);
or U33299 (N_33299,N_25163,N_27635);
xor U33300 (N_33300,N_28261,N_25642);
or U33301 (N_33301,N_26030,N_26650);
nand U33302 (N_33302,N_25251,N_28486);
nand U33303 (N_33303,N_27844,N_26568);
or U33304 (N_33304,N_28295,N_29277);
or U33305 (N_33305,N_29885,N_26860);
or U33306 (N_33306,N_26880,N_28376);
or U33307 (N_33307,N_25678,N_27512);
and U33308 (N_33308,N_26896,N_25092);
nand U33309 (N_33309,N_25006,N_27843);
nor U33310 (N_33310,N_27865,N_28222);
and U33311 (N_33311,N_28748,N_28222);
and U33312 (N_33312,N_28872,N_27465);
and U33313 (N_33313,N_29152,N_28155);
or U33314 (N_33314,N_26815,N_29588);
nor U33315 (N_33315,N_26216,N_28237);
nand U33316 (N_33316,N_28389,N_29874);
and U33317 (N_33317,N_27126,N_28811);
nor U33318 (N_33318,N_28130,N_26327);
and U33319 (N_33319,N_28113,N_26015);
nor U33320 (N_33320,N_29699,N_25559);
and U33321 (N_33321,N_28873,N_25906);
or U33322 (N_33322,N_28862,N_26406);
nor U33323 (N_33323,N_25280,N_27687);
nand U33324 (N_33324,N_28771,N_29153);
xor U33325 (N_33325,N_29304,N_28399);
nand U33326 (N_33326,N_27561,N_26211);
nor U33327 (N_33327,N_27406,N_28348);
or U33328 (N_33328,N_25644,N_28978);
and U33329 (N_33329,N_25692,N_26943);
xnor U33330 (N_33330,N_25585,N_26755);
or U33331 (N_33331,N_25934,N_29554);
nor U33332 (N_33332,N_26883,N_29002);
nor U33333 (N_33333,N_28687,N_28807);
nor U33334 (N_33334,N_27720,N_29199);
nor U33335 (N_33335,N_26664,N_26602);
nor U33336 (N_33336,N_26043,N_28840);
nand U33337 (N_33337,N_27916,N_29397);
and U33338 (N_33338,N_27203,N_29226);
nor U33339 (N_33339,N_28266,N_26862);
and U33340 (N_33340,N_27564,N_28032);
nand U33341 (N_33341,N_27360,N_25139);
nor U33342 (N_33342,N_27417,N_27675);
or U33343 (N_33343,N_28239,N_28964);
nand U33344 (N_33344,N_26123,N_29908);
nand U33345 (N_33345,N_27805,N_29708);
and U33346 (N_33346,N_26669,N_27241);
and U33347 (N_33347,N_27150,N_25241);
nand U33348 (N_33348,N_25107,N_29882);
nand U33349 (N_33349,N_25874,N_27609);
xor U33350 (N_33350,N_26656,N_27809);
nand U33351 (N_33351,N_28244,N_25213);
and U33352 (N_33352,N_28795,N_28151);
or U33353 (N_33353,N_26994,N_26849);
and U33354 (N_33354,N_28342,N_27351);
nor U33355 (N_33355,N_29235,N_25147);
nand U33356 (N_33356,N_29015,N_27534);
nor U33357 (N_33357,N_27705,N_29938);
and U33358 (N_33358,N_25120,N_27723);
nor U33359 (N_33359,N_27328,N_26562);
or U33360 (N_33360,N_26590,N_25142);
nor U33361 (N_33361,N_28938,N_29161);
nor U33362 (N_33362,N_25920,N_27699);
and U33363 (N_33363,N_28069,N_29302);
xor U33364 (N_33364,N_27090,N_26789);
or U33365 (N_33365,N_29304,N_25541);
and U33366 (N_33366,N_26314,N_25416);
and U33367 (N_33367,N_27182,N_29690);
nand U33368 (N_33368,N_25740,N_27296);
nand U33369 (N_33369,N_27638,N_27233);
and U33370 (N_33370,N_29757,N_28920);
and U33371 (N_33371,N_28493,N_29698);
nor U33372 (N_33372,N_27201,N_25359);
nand U33373 (N_33373,N_28686,N_27854);
nor U33374 (N_33374,N_27298,N_29763);
or U33375 (N_33375,N_27246,N_28664);
and U33376 (N_33376,N_27512,N_26437);
xnor U33377 (N_33377,N_29939,N_28908);
nand U33378 (N_33378,N_26768,N_27314);
and U33379 (N_33379,N_25938,N_29634);
or U33380 (N_33380,N_26105,N_27249);
nor U33381 (N_33381,N_26240,N_25328);
or U33382 (N_33382,N_27905,N_29118);
nand U33383 (N_33383,N_28094,N_27836);
nand U33384 (N_33384,N_29734,N_28916);
nand U33385 (N_33385,N_27851,N_25549);
and U33386 (N_33386,N_29713,N_27188);
or U33387 (N_33387,N_25808,N_26132);
xnor U33388 (N_33388,N_27248,N_25903);
nor U33389 (N_33389,N_26635,N_27400);
nor U33390 (N_33390,N_25276,N_29446);
nand U33391 (N_33391,N_26704,N_25574);
or U33392 (N_33392,N_29243,N_29933);
nand U33393 (N_33393,N_26543,N_26832);
and U33394 (N_33394,N_28733,N_26437);
xnor U33395 (N_33395,N_28878,N_28870);
nor U33396 (N_33396,N_25318,N_25657);
nand U33397 (N_33397,N_26201,N_27846);
xnor U33398 (N_33398,N_29352,N_28218);
or U33399 (N_33399,N_26825,N_25457);
nor U33400 (N_33400,N_27008,N_27381);
nor U33401 (N_33401,N_28306,N_28168);
or U33402 (N_33402,N_28615,N_26692);
nand U33403 (N_33403,N_25083,N_27358);
or U33404 (N_33404,N_28695,N_26877);
nand U33405 (N_33405,N_25672,N_25336);
nand U33406 (N_33406,N_29082,N_25306);
nand U33407 (N_33407,N_26223,N_25498);
nor U33408 (N_33408,N_27456,N_26918);
or U33409 (N_33409,N_29972,N_28510);
nor U33410 (N_33410,N_29062,N_28068);
nor U33411 (N_33411,N_29780,N_26255);
or U33412 (N_33412,N_29866,N_27375);
nand U33413 (N_33413,N_28419,N_27622);
nand U33414 (N_33414,N_27036,N_26488);
xor U33415 (N_33415,N_27520,N_29745);
nor U33416 (N_33416,N_27640,N_28038);
or U33417 (N_33417,N_25947,N_28761);
nand U33418 (N_33418,N_27341,N_29717);
or U33419 (N_33419,N_25368,N_28429);
nand U33420 (N_33420,N_28920,N_27072);
nand U33421 (N_33421,N_28722,N_26109);
or U33422 (N_33422,N_28985,N_25611);
xor U33423 (N_33423,N_28859,N_28350);
nor U33424 (N_33424,N_27915,N_27054);
nand U33425 (N_33425,N_29614,N_29504);
nand U33426 (N_33426,N_27476,N_27028);
nor U33427 (N_33427,N_29862,N_25229);
and U33428 (N_33428,N_28488,N_25100);
nand U33429 (N_33429,N_26226,N_27372);
nand U33430 (N_33430,N_28659,N_25916);
and U33431 (N_33431,N_29330,N_25222);
and U33432 (N_33432,N_28314,N_28381);
nor U33433 (N_33433,N_26782,N_27872);
nand U33434 (N_33434,N_25173,N_29111);
xor U33435 (N_33435,N_26026,N_27861);
xor U33436 (N_33436,N_28989,N_26837);
nand U33437 (N_33437,N_25117,N_25266);
nor U33438 (N_33438,N_26888,N_29270);
nand U33439 (N_33439,N_28513,N_26364);
nand U33440 (N_33440,N_27058,N_28275);
and U33441 (N_33441,N_26637,N_25358);
and U33442 (N_33442,N_27183,N_26031);
and U33443 (N_33443,N_25967,N_26756);
nor U33444 (N_33444,N_25594,N_27167);
nand U33445 (N_33445,N_27377,N_26757);
nand U33446 (N_33446,N_27017,N_25426);
and U33447 (N_33447,N_26375,N_26655);
nor U33448 (N_33448,N_27843,N_27753);
nand U33449 (N_33449,N_28006,N_26266);
nand U33450 (N_33450,N_27228,N_25209);
or U33451 (N_33451,N_25024,N_29317);
nor U33452 (N_33452,N_26189,N_28614);
or U33453 (N_33453,N_26522,N_26132);
nand U33454 (N_33454,N_29670,N_26589);
nor U33455 (N_33455,N_28835,N_26634);
xor U33456 (N_33456,N_28622,N_25476);
nand U33457 (N_33457,N_27976,N_25823);
and U33458 (N_33458,N_29217,N_27699);
and U33459 (N_33459,N_29211,N_26563);
xnor U33460 (N_33460,N_28311,N_26666);
nand U33461 (N_33461,N_28094,N_29443);
or U33462 (N_33462,N_28904,N_28821);
nor U33463 (N_33463,N_26315,N_27594);
xnor U33464 (N_33464,N_28138,N_26607);
nor U33465 (N_33465,N_29854,N_25656);
or U33466 (N_33466,N_29441,N_27097);
nand U33467 (N_33467,N_25015,N_27021);
or U33468 (N_33468,N_29151,N_29716);
or U33469 (N_33469,N_28822,N_27074);
or U33470 (N_33470,N_25692,N_29611);
and U33471 (N_33471,N_29595,N_27662);
nand U33472 (N_33472,N_25608,N_25540);
nand U33473 (N_33473,N_27976,N_25783);
or U33474 (N_33474,N_28034,N_25492);
nor U33475 (N_33475,N_27157,N_25709);
and U33476 (N_33476,N_29799,N_25919);
or U33477 (N_33477,N_29121,N_25706);
and U33478 (N_33478,N_26842,N_28959);
nor U33479 (N_33479,N_29509,N_26609);
or U33480 (N_33480,N_27645,N_28609);
xor U33481 (N_33481,N_25185,N_29327);
and U33482 (N_33482,N_25285,N_27591);
nand U33483 (N_33483,N_25069,N_29110);
nand U33484 (N_33484,N_27122,N_25955);
or U33485 (N_33485,N_29518,N_27230);
or U33486 (N_33486,N_29507,N_26836);
nand U33487 (N_33487,N_25608,N_29252);
nor U33488 (N_33488,N_27296,N_29169);
nor U33489 (N_33489,N_25255,N_29327);
and U33490 (N_33490,N_26345,N_27919);
nor U33491 (N_33491,N_26534,N_26194);
nand U33492 (N_33492,N_29621,N_29544);
or U33493 (N_33493,N_25522,N_26222);
nor U33494 (N_33494,N_27572,N_29219);
and U33495 (N_33495,N_28896,N_25539);
nor U33496 (N_33496,N_27190,N_29542);
nor U33497 (N_33497,N_29629,N_29448);
xnor U33498 (N_33498,N_26935,N_27212);
nor U33499 (N_33499,N_26545,N_29084);
or U33500 (N_33500,N_27830,N_25704);
or U33501 (N_33501,N_28014,N_28827);
nor U33502 (N_33502,N_28336,N_29936);
nor U33503 (N_33503,N_26813,N_29231);
or U33504 (N_33504,N_25697,N_27320);
xor U33505 (N_33505,N_25406,N_26887);
or U33506 (N_33506,N_26513,N_27885);
nand U33507 (N_33507,N_29224,N_25373);
and U33508 (N_33508,N_27401,N_27384);
nand U33509 (N_33509,N_28316,N_28792);
and U33510 (N_33510,N_28326,N_26703);
xnor U33511 (N_33511,N_28120,N_29636);
nor U33512 (N_33512,N_28636,N_28292);
nand U33513 (N_33513,N_27116,N_28615);
or U33514 (N_33514,N_27230,N_29505);
nor U33515 (N_33515,N_26870,N_28267);
or U33516 (N_33516,N_29579,N_28577);
nor U33517 (N_33517,N_26182,N_29515);
and U33518 (N_33518,N_29754,N_25422);
or U33519 (N_33519,N_25078,N_29073);
nand U33520 (N_33520,N_28587,N_27701);
or U33521 (N_33521,N_28595,N_25718);
and U33522 (N_33522,N_27474,N_29776);
and U33523 (N_33523,N_27113,N_25670);
nor U33524 (N_33524,N_28043,N_25422);
and U33525 (N_33525,N_27861,N_28111);
and U33526 (N_33526,N_28705,N_26923);
or U33527 (N_33527,N_28804,N_27272);
or U33528 (N_33528,N_27742,N_29766);
nand U33529 (N_33529,N_28102,N_25378);
nand U33530 (N_33530,N_27526,N_25942);
xnor U33531 (N_33531,N_25236,N_26986);
nor U33532 (N_33532,N_28599,N_27926);
nor U33533 (N_33533,N_27909,N_27982);
nand U33534 (N_33534,N_29577,N_25701);
or U33535 (N_33535,N_25380,N_28006);
nand U33536 (N_33536,N_28325,N_27619);
and U33537 (N_33537,N_27374,N_26892);
nor U33538 (N_33538,N_29070,N_29404);
xnor U33539 (N_33539,N_26852,N_28746);
and U33540 (N_33540,N_28365,N_29676);
or U33541 (N_33541,N_28873,N_25789);
nand U33542 (N_33542,N_29641,N_25449);
nand U33543 (N_33543,N_26835,N_26231);
and U33544 (N_33544,N_29279,N_27451);
and U33545 (N_33545,N_27597,N_27815);
nor U33546 (N_33546,N_25220,N_27783);
nor U33547 (N_33547,N_28679,N_27942);
or U33548 (N_33548,N_28130,N_29481);
and U33549 (N_33549,N_25520,N_27805);
nand U33550 (N_33550,N_26725,N_29546);
or U33551 (N_33551,N_25081,N_25085);
and U33552 (N_33552,N_27976,N_26052);
nand U33553 (N_33553,N_27612,N_29463);
nor U33554 (N_33554,N_27812,N_27118);
and U33555 (N_33555,N_26620,N_29138);
xor U33556 (N_33556,N_26189,N_26174);
nor U33557 (N_33557,N_28059,N_25181);
nand U33558 (N_33558,N_28764,N_26652);
nand U33559 (N_33559,N_28182,N_26053);
and U33560 (N_33560,N_26975,N_26326);
nand U33561 (N_33561,N_26478,N_28620);
or U33562 (N_33562,N_27330,N_25449);
or U33563 (N_33563,N_29641,N_28096);
and U33564 (N_33564,N_27960,N_25790);
or U33565 (N_33565,N_25018,N_27479);
nor U33566 (N_33566,N_29761,N_29896);
nor U33567 (N_33567,N_28377,N_28347);
nor U33568 (N_33568,N_29683,N_27952);
and U33569 (N_33569,N_27028,N_27500);
nand U33570 (N_33570,N_25980,N_29406);
xnor U33571 (N_33571,N_28034,N_26185);
nor U33572 (N_33572,N_27353,N_28801);
nand U33573 (N_33573,N_29241,N_27531);
xnor U33574 (N_33574,N_28864,N_29774);
and U33575 (N_33575,N_25127,N_25407);
and U33576 (N_33576,N_29616,N_28561);
nand U33577 (N_33577,N_29763,N_28035);
or U33578 (N_33578,N_25673,N_27433);
xnor U33579 (N_33579,N_27872,N_25361);
or U33580 (N_33580,N_28570,N_27508);
nand U33581 (N_33581,N_27777,N_26434);
and U33582 (N_33582,N_26733,N_26912);
nor U33583 (N_33583,N_29001,N_28161);
or U33584 (N_33584,N_29724,N_28725);
nand U33585 (N_33585,N_25371,N_25585);
and U33586 (N_33586,N_29567,N_25060);
and U33587 (N_33587,N_27428,N_28242);
nor U33588 (N_33588,N_26828,N_28800);
xnor U33589 (N_33589,N_25803,N_29432);
nand U33590 (N_33590,N_27483,N_29731);
nor U33591 (N_33591,N_28775,N_26296);
or U33592 (N_33592,N_28997,N_29331);
nor U33593 (N_33593,N_27012,N_28266);
nand U33594 (N_33594,N_25177,N_26630);
nor U33595 (N_33595,N_29665,N_27399);
xnor U33596 (N_33596,N_25750,N_27000);
or U33597 (N_33597,N_29538,N_29324);
or U33598 (N_33598,N_27158,N_25320);
nor U33599 (N_33599,N_27149,N_29504);
xor U33600 (N_33600,N_25219,N_26277);
nand U33601 (N_33601,N_27221,N_27190);
and U33602 (N_33602,N_26527,N_29360);
nand U33603 (N_33603,N_25592,N_27314);
or U33604 (N_33604,N_25834,N_27254);
and U33605 (N_33605,N_25571,N_26293);
nand U33606 (N_33606,N_26664,N_29354);
nor U33607 (N_33607,N_25897,N_27718);
and U33608 (N_33608,N_27786,N_25549);
nand U33609 (N_33609,N_28847,N_28263);
nand U33610 (N_33610,N_27512,N_25586);
and U33611 (N_33611,N_27959,N_25401);
and U33612 (N_33612,N_25004,N_26297);
or U33613 (N_33613,N_25122,N_28129);
and U33614 (N_33614,N_29054,N_26986);
nor U33615 (N_33615,N_28608,N_25601);
or U33616 (N_33616,N_28323,N_27727);
and U33617 (N_33617,N_25136,N_26562);
nand U33618 (N_33618,N_26317,N_26762);
nand U33619 (N_33619,N_29617,N_28455);
nand U33620 (N_33620,N_27953,N_28761);
nand U33621 (N_33621,N_27561,N_27458);
nor U33622 (N_33622,N_26659,N_26149);
nor U33623 (N_33623,N_27681,N_25378);
xor U33624 (N_33624,N_25757,N_26295);
nand U33625 (N_33625,N_26230,N_26870);
nor U33626 (N_33626,N_26898,N_27236);
and U33627 (N_33627,N_26978,N_27069);
or U33628 (N_33628,N_28916,N_27869);
or U33629 (N_33629,N_27345,N_29942);
and U33630 (N_33630,N_28573,N_25830);
nand U33631 (N_33631,N_27346,N_29692);
nor U33632 (N_33632,N_29161,N_27736);
nor U33633 (N_33633,N_26525,N_28631);
and U33634 (N_33634,N_25806,N_27817);
or U33635 (N_33635,N_29446,N_25830);
and U33636 (N_33636,N_26049,N_26166);
nor U33637 (N_33637,N_28295,N_26148);
xnor U33638 (N_33638,N_26555,N_26323);
or U33639 (N_33639,N_26696,N_28151);
or U33640 (N_33640,N_29885,N_27475);
or U33641 (N_33641,N_25029,N_26465);
nand U33642 (N_33642,N_27433,N_28643);
xnor U33643 (N_33643,N_28345,N_27045);
xor U33644 (N_33644,N_26233,N_26327);
nand U33645 (N_33645,N_25125,N_27715);
or U33646 (N_33646,N_25367,N_27887);
nor U33647 (N_33647,N_28627,N_27566);
and U33648 (N_33648,N_28981,N_27901);
and U33649 (N_33649,N_28203,N_25945);
and U33650 (N_33650,N_25323,N_27733);
and U33651 (N_33651,N_26988,N_29738);
xnor U33652 (N_33652,N_26816,N_29735);
and U33653 (N_33653,N_27537,N_27590);
nor U33654 (N_33654,N_29298,N_26621);
xnor U33655 (N_33655,N_27596,N_25929);
and U33656 (N_33656,N_29920,N_28265);
nand U33657 (N_33657,N_28021,N_29587);
or U33658 (N_33658,N_29560,N_29508);
and U33659 (N_33659,N_29788,N_29391);
and U33660 (N_33660,N_28557,N_27093);
xor U33661 (N_33661,N_28465,N_26340);
or U33662 (N_33662,N_29577,N_29543);
nor U33663 (N_33663,N_29806,N_28848);
and U33664 (N_33664,N_26798,N_27383);
nand U33665 (N_33665,N_25080,N_29935);
nand U33666 (N_33666,N_26713,N_29533);
and U33667 (N_33667,N_28610,N_29170);
and U33668 (N_33668,N_29099,N_27430);
or U33669 (N_33669,N_25080,N_26426);
and U33670 (N_33670,N_27517,N_27970);
and U33671 (N_33671,N_29880,N_25966);
nand U33672 (N_33672,N_26199,N_25495);
or U33673 (N_33673,N_25134,N_29990);
or U33674 (N_33674,N_27999,N_28683);
nor U33675 (N_33675,N_28412,N_27442);
and U33676 (N_33676,N_25425,N_27603);
nor U33677 (N_33677,N_27557,N_28664);
and U33678 (N_33678,N_25415,N_29503);
xnor U33679 (N_33679,N_26126,N_29851);
or U33680 (N_33680,N_27810,N_26187);
nor U33681 (N_33681,N_28077,N_29869);
or U33682 (N_33682,N_29860,N_25225);
or U33683 (N_33683,N_26915,N_26801);
or U33684 (N_33684,N_29641,N_25819);
xor U33685 (N_33685,N_28647,N_29029);
or U33686 (N_33686,N_29282,N_25352);
nor U33687 (N_33687,N_29127,N_29632);
xnor U33688 (N_33688,N_25225,N_27252);
and U33689 (N_33689,N_26241,N_29924);
nor U33690 (N_33690,N_27406,N_29849);
nand U33691 (N_33691,N_29481,N_25871);
and U33692 (N_33692,N_25867,N_27033);
or U33693 (N_33693,N_27515,N_27551);
and U33694 (N_33694,N_29088,N_25076);
xnor U33695 (N_33695,N_29554,N_28302);
nand U33696 (N_33696,N_29617,N_25059);
and U33697 (N_33697,N_28792,N_26701);
or U33698 (N_33698,N_28220,N_27190);
nand U33699 (N_33699,N_29789,N_27260);
or U33700 (N_33700,N_25097,N_27251);
nand U33701 (N_33701,N_25741,N_27630);
and U33702 (N_33702,N_26490,N_29338);
and U33703 (N_33703,N_25327,N_28234);
or U33704 (N_33704,N_28916,N_28072);
or U33705 (N_33705,N_26654,N_27913);
or U33706 (N_33706,N_25166,N_27662);
nand U33707 (N_33707,N_29306,N_28221);
or U33708 (N_33708,N_27269,N_26890);
and U33709 (N_33709,N_26100,N_25009);
nor U33710 (N_33710,N_28326,N_29817);
or U33711 (N_33711,N_27701,N_25149);
and U33712 (N_33712,N_26940,N_26906);
nor U33713 (N_33713,N_25121,N_27558);
or U33714 (N_33714,N_29431,N_26134);
nand U33715 (N_33715,N_26395,N_29323);
nor U33716 (N_33716,N_25528,N_29147);
nor U33717 (N_33717,N_26424,N_29734);
nor U33718 (N_33718,N_26142,N_27524);
xnor U33719 (N_33719,N_27420,N_27763);
nor U33720 (N_33720,N_29606,N_26826);
or U33721 (N_33721,N_26112,N_29796);
nor U33722 (N_33722,N_29801,N_29734);
or U33723 (N_33723,N_26408,N_26744);
or U33724 (N_33724,N_29300,N_28371);
and U33725 (N_33725,N_28570,N_27256);
or U33726 (N_33726,N_28752,N_29999);
or U33727 (N_33727,N_27595,N_26394);
nor U33728 (N_33728,N_26926,N_25127);
or U33729 (N_33729,N_27990,N_25069);
and U33730 (N_33730,N_29940,N_28488);
nand U33731 (N_33731,N_26386,N_26416);
nand U33732 (N_33732,N_25933,N_29884);
nor U33733 (N_33733,N_26646,N_29986);
or U33734 (N_33734,N_26125,N_28009);
and U33735 (N_33735,N_28704,N_25449);
nor U33736 (N_33736,N_25908,N_29938);
nor U33737 (N_33737,N_29651,N_26581);
or U33738 (N_33738,N_27441,N_28585);
and U33739 (N_33739,N_25446,N_25111);
or U33740 (N_33740,N_25407,N_26688);
or U33741 (N_33741,N_27504,N_27762);
nor U33742 (N_33742,N_29903,N_28520);
or U33743 (N_33743,N_29826,N_29827);
nand U33744 (N_33744,N_29265,N_28822);
nor U33745 (N_33745,N_27463,N_26352);
and U33746 (N_33746,N_28363,N_29046);
and U33747 (N_33747,N_26000,N_29188);
nand U33748 (N_33748,N_28239,N_26955);
and U33749 (N_33749,N_26264,N_28251);
nand U33750 (N_33750,N_27043,N_25997);
xor U33751 (N_33751,N_27165,N_26420);
nor U33752 (N_33752,N_25156,N_27921);
nor U33753 (N_33753,N_28883,N_29625);
and U33754 (N_33754,N_27312,N_26832);
nor U33755 (N_33755,N_27043,N_29672);
and U33756 (N_33756,N_26714,N_28068);
nand U33757 (N_33757,N_25977,N_25604);
and U33758 (N_33758,N_29215,N_29013);
or U33759 (N_33759,N_28076,N_26910);
or U33760 (N_33760,N_28013,N_28240);
nor U33761 (N_33761,N_28140,N_28483);
xnor U33762 (N_33762,N_26134,N_25051);
or U33763 (N_33763,N_25344,N_26459);
nor U33764 (N_33764,N_25478,N_27753);
nor U33765 (N_33765,N_26930,N_26979);
xnor U33766 (N_33766,N_27879,N_27412);
or U33767 (N_33767,N_26874,N_25169);
xnor U33768 (N_33768,N_27726,N_28952);
nor U33769 (N_33769,N_26982,N_26913);
nor U33770 (N_33770,N_29989,N_29424);
nor U33771 (N_33771,N_29417,N_26054);
nand U33772 (N_33772,N_29393,N_27346);
nor U33773 (N_33773,N_28476,N_27760);
nand U33774 (N_33774,N_28996,N_27348);
and U33775 (N_33775,N_25231,N_29491);
nand U33776 (N_33776,N_27382,N_26854);
and U33777 (N_33777,N_26696,N_27093);
nor U33778 (N_33778,N_26880,N_26743);
nor U33779 (N_33779,N_28718,N_28728);
xor U33780 (N_33780,N_26343,N_29741);
xor U33781 (N_33781,N_25964,N_27233);
or U33782 (N_33782,N_28124,N_28525);
nor U33783 (N_33783,N_27373,N_26876);
or U33784 (N_33784,N_25897,N_27473);
xor U33785 (N_33785,N_29487,N_27115);
nor U33786 (N_33786,N_25798,N_28136);
or U33787 (N_33787,N_27620,N_27680);
nand U33788 (N_33788,N_25772,N_28804);
nand U33789 (N_33789,N_26412,N_28351);
and U33790 (N_33790,N_28820,N_26864);
nand U33791 (N_33791,N_28488,N_29047);
nor U33792 (N_33792,N_26673,N_25818);
nand U33793 (N_33793,N_28117,N_29249);
and U33794 (N_33794,N_27248,N_27205);
or U33795 (N_33795,N_29700,N_29053);
nor U33796 (N_33796,N_28666,N_26709);
and U33797 (N_33797,N_25489,N_26193);
xnor U33798 (N_33798,N_27143,N_26879);
and U33799 (N_33799,N_25357,N_29046);
xor U33800 (N_33800,N_28004,N_27129);
or U33801 (N_33801,N_28383,N_26841);
nor U33802 (N_33802,N_29565,N_25348);
xnor U33803 (N_33803,N_25450,N_28696);
nand U33804 (N_33804,N_29133,N_28520);
or U33805 (N_33805,N_26929,N_26012);
or U33806 (N_33806,N_29472,N_29438);
or U33807 (N_33807,N_29842,N_28727);
or U33808 (N_33808,N_28903,N_25366);
and U33809 (N_33809,N_25198,N_25553);
nand U33810 (N_33810,N_26701,N_28404);
nand U33811 (N_33811,N_28623,N_26704);
nor U33812 (N_33812,N_27739,N_25217);
nand U33813 (N_33813,N_25498,N_29803);
or U33814 (N_33814,N_28133,N_28763);
or U33815 (N_33815,N_27001,N_29634);
or U33816 (N_33816,N_25507,N_28722);
nand U33817 (N_33817,N_29222,N_26938);
or U33818 (N_33818,N_26510,N_25098);
xor U33819 (N_33819,N_26382,N_27010);
and U33820 (N_33820,N_28044,N_28444);
and U33821 (N_33821,N_27664,N_29461);
and U33822 (N_33822,N_25987,N_27734);
and U33823 (N_33823,N_27197,N_29472);
nand U33824 (N_33824,N_29786,N_27050);
nor U33825 (N_33825,N_26798,N_26700);
nand U33826 (N_33826,N_29815,N_29612);
xor U33827 (N_33827,N_28885,N_25523);
nand U33828 (N_33828,N_27714,N_27319);
xor U33829 (N_33829,N_25440,N_25742);
and U33830 (N_33830,N_26977,N_26261);
and U33831 (N_33831,N_26377,N_26492);
nor U33832 (N_33832,N_28033,N_25987);
nor U33833 (N_33833,N_25963,N_28488);
or U33834 (N_33834,N_29662,N_26901);
nor U33835 (N_33835,N_26107,N_28008);
and U33836 (N_33836,N_25797,N_29900);
nor U33837 (N_33837,N_28178,N_25808);
and U33838 (N_33838,N_25675,N_25637);
nor U33839 (N_33839,N_25995,N_26180);
nor U33840 (N_33840,N_26032,N_25320);
xnor U33841 (N_33841,N_28560,N_27649);
nor U33842 (N_33842,N_25045,N_25699);
and U33843 (N_33843,N_28701,N_28073);
nor U33844 (N_33844,N_28773,N_28251);
nand U33845 (N_33845,N_25429,N_28331);
nor U33846 (N_33846,N_28972,N_27174);
and U33847 (N_33847,N_25099,N_27072);
and U33848 (N_33848,N_26717,N_27399);
or U33849 (N_33849,N_28751,N_26893);
nor U33850 (N_33850,N_27010,N_28079);
nand U33851 (N_33851,N_28228,N_29377);
nand U33852 (N_33852,N_25455,N_28352);
nor U33853 (N_33853,N_28759,N_29310);
or U33854 (N_33854,N_29844,N_28583);
or U33855 (N_33855,N_25961,N_25234);
nand U33856 (N_33856,N_27151,N_26652);
nand U33857 (N_33857,N_29550,N_26711);
nor U33858 (N_33858,N_28173,N_25140);
or U33859 (N_33859,N_28038,N_27946);
or U33860 (N_33860,N_28536,N_27762);
nor U33861 (N_33861,N_26955,N_27939);
xnor U33862 (N_33862,N_27829,N_29290);
nand U33863 (N_33863,N_26624,N_29997);
or U33864 (N_33864,N_27772,N_25099);
xnor U33865 (N_33865,N_27623,N_25613);
nor U33866 (N_33866,N_25115,N_26317);
or U33867 (N_33867,N_29736,N_27030);
nand U33868 (N_33868,N_27145,N_26150);
or U33869 (N_33869,N_28838,N_27426);
nand U33870 (N_33870,N_26524,N_25121);
and U33871 (N_33871,N_25150,N_29272);
or U33872 (N_33872,N_28753,N_28696);
xnor U33873 (N_33873,N_28250,N_27440);
nor U33874 (N_33874,N_25624,N_28962);
xor U33875 (N_33875,N_25773,N_27493);
xnor U33876 (N_33876,N_27346,N_28031);
xor U33877 (N_33877,N_28261,N_27428);
nor U33878 (N_33878,N_29561,N_27217);
nor U33879 (N_33879,N_28109,N_25582);
and U33880 (N_33880,N_29125,N_27870);
or U33881 (N_33881,N_29241,N_28689);
nor U33882 (N_33882,N_26859,N_28590);
and U33883 (N_33883,N_29875,N_27216);
nand U33884 (N_33884,N_28959,N_26185);
and U33885 (N_33885,N_27142,N_28311);
or U33886 (N_33886,N_26807,N_25723);
and U33887 (N_33887,N_29921,N_25980);
nor U33888 (N_33888,N_29983,N_29166);
and U33889 (N_33889,N_28582,N_26391);
nor U33890 (N_33890,N_26671,N_27953);
nand U33891 (N_33891,N_26208,N_27891);
and U33892 (N_33892,N_29561,N_29079);
nor U33893 (N_33893,N_29273,N_29426);
xor U33894 (N_33894,N_25023,N_28842);
and U33895 (N_33895,N_25204,N_26868);
or U33896 (N_33896,N_26994,N_28345);
or U33897 (N_33897,N_29504,N_26977);
or U33898 (N_33898,N_25141,N_25786);
nand U33899 (N_33899,N_25057,N_26421);
or U33900 (N_33900,N_28418,N_27188);
nor U33901 (N_33901,N_25130,N_29483);
or U33902 (N_33902,N_29597,N_25868);
or U33903 (N_33903,N_25748,N_29074);
nand U33904 (N_33904,N_26082,N_27524);
or U33905 (N_33905,N_25190,N_26300);
nand U33906 (N_33906,N_25499,N_25555);
and U33907 (N_33907,N_25678,N_28164);
nor U33908 (N_33908,N_28657,N_29001);
or U33909 (N_33909,N_27296,N_27519);
nand U33910 (N_33910,N_27283,N_28520);
and U33911 (N_33911,N_29041,N_29628);
xor U33912 (N_33912,N_26954,N_26322);
and U33913 (N_33913,N_29930,N_25679);
nor U33914 (N_33914,N_26106,N_25682);
nand U33915 (N_33915,N_29681,N_26220);
nand U33916 (N_33916,N_26690,N_25993);
nor U33917 (N_33917,N_29570,N_25584);
or U33918 (N_33918,N_29649,N_27197);
or U33919 (N_33919,N_29266,N_25696);
nand U33920 (N_33920,N_25475,N_25681);
or U33921 (N_33921,N_28941,N_29358);
and U33922 (N_33922,N_27096,N_29885);
or U33923 (N_33923,N_28436,N_25301);
nand U33924 (N_33924,N_28265,N_28662);
or U33925 (N_33925,N_29459,N_26296);
nand U33926 (N_33926,N_28109,N_29544);
and U33927 (N_33927,N_25247,N_26772);
or U33928 (N_33928,N_29246,N_28486);
or U33929 (N_33929,N_28529,N_25319);
nor U33930 (N_33930,N_25007,N_27693);
or U33931 (N_33931,N_28607,N_28696);
nand U33932 (N_33932,N_29034,N_28274);
nand U33933 (N_33933,N_27188,N_26741);
or U33934 (N_33934,N_25443,N_27660);
nand U33935 (N_33935,N_25789,N_29050);
or U33936 (N_33936,N_26592,N_27601);
nand U33937 (N_33937,N_29705,N_25324);
or U33938 (N_33938,N_26043,N_27193);
xnor U33939 (N_33939,N_28761,N_29840);
xor U33940 (N_33940,N_28583,N_25345);
or U33941 (N_33941,N_26110,N_27390);
nand U33942 (N_33942,N_29878,N_29252);
or U33943 (N_33943,N_28759,N_25301);
or U33944 (N_33944,N_25963,N_28509);
or U33945 (N_33945,N_26839,N_28792);
nor U33946 (N_33946,N_26263,N_29970);
or U33947 (N_33947,N_27716,N_25603);
and U33948 (N_33948,N_26351,N_27073);
nand U33949 (N_33949,N_25626,N_29776);
nor U33950 (N_33950,N_28844,N_28050);
nor U33951 (N_33951,N_25785,N_25651);
nand U33952 (N_33952,N_28195,N_29780);
nand U33953 (N_33953,N_26106,N_26287);
and U33954 (N_33954,N_26581,N_27427);
nor U33955 (N_33955,N_26271,N_29477);
nor U33956 (N_33956,N_25479,N_29296);
or U33957 (N_33957,N_29852,N_26031);
nand U33958 (N_33958,N_27247,N_27011);
nand U33959 (N_33959,N_26439,N_25306);
nand U33960 (N_33960,N_25691,N_28860);
and U33961 (N_33961,N_25874,N_29996);
nand U33962 (N_33962,N_26212,N_29129);
and U33963 (N_33963,N_26401,N_25680);
nand U33964 (N_33964,N_29114,N_25531);
or U33965 (N_33965,N_28382,N_28755);
nand U33966 (N_33966,N_29353,N_27011);
nand U33967 (N_33967,N_29216,N_27209);
or U33968 (N_33968,N_28459,N_28764);
or U33969 (N_33969,N_29456,N_28526);
xnor U33970 (N_33970,N_25536,N_28924);
or U33971 (N_33971,N_27821,N_25937);
or U33972 (N_33972,N_26833,N_28517);
or U33973 (N_33973,N_27006,N_27749);
or U33974 (N_33974,N_29046,N_29497);
nand U33975 (N_33975,N_28543,N_28480);
nor U33976 (N_33976,N_27950,N_29184);
nand U33977 (N_33977,N_27518,N_27952);
nand U33978 (N_33978,N_27369,N_25253);
or U33979 (N_33979,N_29873,N_26306);
and U33980 (N_33980,N_29885,N_26095);
xor U33981 (N_33981,N_28594,N_29635);
nand U33982 (N_33982,N_26201,N_29691);
and U33983 (N_33983,N_28626,N_25140);
or U33984 (N_33984,N_25673,N_26865);
nand U33985 (N_33985,N_26359,N_28844);
nor U33986 (N_33986,N_26601,N_27700);
and U33987 (N_33987,N_25135,N_26943);
nand U33988 (N_33988,N_28165,N_26896);
nor U33989 (N_33989,N_26935,N_27333);
xnor U33990 (N_33990,N_28170,N_28369);
or U33991 (N_33991,N_27587,N_25901);
nand U33992 (N_33992,N_27100,N_25740);
or U33993 (N_33993,N_26301,N_26563);
or U33994 (N_33994,N_29169,N_26699);
and U33995 (N_33995,N_29713,N_29334);
or U33996 (N_33996,N_28114,N_26230);
or U33997 (N_33997,N_29476,N_27728);
or U33998 (N_33998,N_25592,N_28821);
nand U33999 (N_33999,N_29397,N_28112);
or U34000 (N_34000,N_29631,N_25525);
or U34001 (N_34001,N_26331,N_26842);
or U34002 (N_34002,N_25017,N_27231);
nand U34003 (N_34003,N_28245,N_28055);
xnor U34004 (N_34004,N_27365,N_25520);
and U34005 (N_34005,N_28183,N_28909);
and U34006 (N_34006,N_28553,N_29635);
or U34007 (N_34007,N_28640,N_28259);
nor U34008 (N_34008,N_26760,N_26929);
or U34009 (N_34009,N_27400,N_26657);
and U34010 (N_34010,N_25052,N_29233);
nand U34011 (N_34011,N_25473,N_27732);
nand U34012 (N_34012,N_27363,N_27715);
nand U34013 (N_34013,N_29222,N_25724);
nand U34014 (N_34014,N_28805,N_27467);
and U34015 (N_34015,N_28539,N_28918);
nand U34016 (N_34016,N_26474,N_28516);
nor U34017 (N_34017,N_26221,N_25270);
nor U34018 (N_34018,N_29028,N_28078);
nand U34019 (N_34019,N_26068,N_25952);
nor U34020 (N_34020,N_27855,N_26082);
or U34021 (N_34021,N_25672,N_25360);
or U34022 (N_34022,N_28000,N_29876);
nand U34023 (N_34023,N_27691,N_27487);
nor U34024 (N_34024,N_29987,N_28323);
or U34025 (N_34025,N_26554,N_25728);
and U34026 (N_34026,N_29428,N_27635);
or U34027 (N_34027,N_28007,N_27803);
and U34028 (N_34028,N_26156,N_25711);
nor U34029 (N_34029,N_26403,N_29193);
nor U34030 (N_34030,N_29759,N_29225);
xnor U34031 (N_34031,N_29817,N_27537);
nand U34032 (N_34032,N_26125,N_29350);
nand U34033 (N_34033,N_29486,N_26663);
nor U34034 (N_34034,N_25004,N_27417);
nand U34035 (N_34035,N_26904,N_28984);
nand U34036 (N_34036,N_25349,N_28105);
nor U34037 (N_34037,N_27952,N_27006);
and U34038 (N_34038,N_29072,N_26836);
or U34039 (N_34039,N_28481,N_26485);
and U34040 (N_34040,N_25221,N_29051);
and U34041 (N_34041,N_27302,N_28843);
nor U34042 (N_34042,N_28054,N_29779);
xor U34043 (N_34043,N_27801,N_25316);
xnor U34044 (N_34044,N_25517,N_26786);
nor U34045 (N_34045,N_29641,N_26280);
nand U34046 (N_34046,N_26045,N_25495);
nand U34047 (N_34047,N_27917,N_27753);
nor U34048 (N_34048,N_26792,N_26759);
nand U34049 (N_34049,N_26624,N_26843);
nor U34050 (N_34050,N_27912,N_27726);
and U34051 (N_34051,N_26968,N_25877);
or U34052 (N_34052,N_26702,N_29871);
or U34053 (N_34053,N_25251,N_29013);
nor U34054 (N_34054,N_28497,N_29067);
nand U34055 (N_34055,N_25630,N_29954);
nor U34056 (N_34056,N_25134,N_29626);
nand U34057 (N_34057,N_26012,N_26960);
or U34058 (N_34058,N_27924,N_26992);
or U34059 (N_34059,N_25535,N_26359);
or U34060 (N_34060,N_29985,N_29112);
and U34061 (N_34061,N_27818,N_29036);
or U34062 (N_34062,N_27610,N_25731);
nor U34063 (N_34063,N_29291,N_28635);
or U34064 (N_34064,N_27288,N_27489);
xnor U34065 (N_34065,N_26079,N_25490);
xor U34066 (N_34066,N_25515,N_29953);
nand U34067 (N_34067,N_28992,N_25489);
xnor U34068 (N_34068,N_25486,N_25144);
and U34069 (N_34069,N_26022,N_25358);
or U34070 (N_34070,N_25416,N_26029);
nand U34071 (N_34071,N_25209,N_27451);
nand U34072 (N_34072,N_26886,N_28684);
and U34073 (N_34073,N_26666,N_27254);
or U34074 (N_34074,N_25025,N_29998);
xnor U34075 (N_34075,N_25759,N_28137);
or U34076 (N_34076,N_25905,N_28849);
nor U34077 (N_34077,N_26639,N_25052);
nor U34078 (N_34078,N_29629,N_27471);
and U34079 (N_34079,N_26619,N_26225);
nand U34080 (N_34080,N_29568,N_28018);
or U34081 (N_34081,N_26436,N_26426);
nand U34082 (N_34082,N_28735,N_25058);
or U34083 (N_34083,N_25893,N_29866);
or U34084 (N_34084,N_28979,N_28317);
and U34085 (N_34085,N_25709,N_25282);
or U34086 (N_34086,N_25621,N_26127);
nor U34087 (N_34087,N_26559,N_26125);
and U34088 (N_34088,N_29102,N_29613);
nor U34089 (N_34089,N_29839,N_28306);
nor U34090 (N_34090,N_28017,N_26077);
nand U34091 (N_34091,N_28258,N_28022);
or U34092 (N_34092,N_25837,N_29230);
nand U34093 (N_34093,N_29408,N_27315);
xor U34094 (N_34094,N_27924,N_28498);
nor U34095 (N_34095,N_26949,N_27921);
nand U34096 (N_34096,N_25327,N_29349);
nand U34097 (N_34097,N_25000,N_29699);
xor U34098 (N_34098,N_26535,N_28018);
and U34099 (N_34099,N_26821,N_28970);
nand U34100 (N_34100,N_26285,N_28604);
nor U34101 (N_34101,N_29985,N_28590);
nand U34102 (N_34102,N_27642,N_27940);
nand U34103 (N_34103,N_26251,N_28210);
or U34104 (N_34104,N_28771,N_27683);
or U34105 (N_34105,N_26465,N_26178);
nand U34106 (N_34106,N_27378,N_29936);
nor U34107 (N_34107,N_25034,N_29850);
and U34108 (N_34108,N_27055,N_26896);
nand U34109 (N_34109,N_26532,N_25333);
xor U34110 (N_34110,N_29260,N_25692);
or U34111 (N_34111,N_25859,N_28816);
nor U34112 (N_34112,N_27800,N_27315);
nand U34113 (N_34113,N_25617,N_28405);
or U34114 (N_34114,N_25520,N_25076);
and U34115 (N_34115,N_27429,N_29061);
xnor U34116 (N_34116,N_25207,N_25444);
xor U34117 (N_34117,N_26738,N_28505);
nand U34118 (N_34118,N_28422,N_26067);
and U34119 (N_34119,N_26352,N_27134);
or U34120 (N_34120,N_29318,N_29388);
nand U34121 (N_34121,N_26148,N_29998);
xor U34122 (N_34122,N_25216,N_29330);
and U34123 (N_34123,N_25982,N_29837);
nand U34124 (N_34124,N_26282,N_28975);
and U34125 (N_34125,N_27408,N_26856);
and U34126 (N_34126,N_26377,N_26184);
nor U34127 (N_34127,N_29055,N_29546);
and U34128 (N_34128,N_27719,N_28193);
nand U34129 (N_34129,N_26178,N_26400);
or U34130 (N_34130,N_29678,N_27062);
or U34131 (N_34131,N_25194,N_28805);
or U34132 (N_34132,N_25603,N_25174);
and U34133 (N_34133,N_28309,N_25224);
nor U34134 (N_34134,N_27483,N_27075);
nor U34135 (N_34135,N_29730,N_26466);
xnor U34136 (N_34136,N_26271,N_27986);
nand U34137 (N_34137,N_25975,N_27523);
nand U34138 (N_34138,N_29064,N_25844);
or U34139 (N_34139,N_25472,N_27040);
xor U34140 (N_34140,N_29507,N_26182);
nand U34141 (N_34141,N_29771,N_29808);
xnor U34142 (N_34142,N_25402,N_27083);
and U34143 (N_34143,N_25479,N_26327);
or U34144 (N_34144,N_27921,N_29021);
and U34145 (N_34145,N_27890,N_29597);
and U34146 (N_34146,N_25107,N_25760);
nand U34147 (N_34147,N_26200,N_26769);
nor U34148 (N_34148,N_29833,N_26519);
nand U34149 (N_34149,N_26687,N_29797);
or U34150 (N_34150,N_29012,N_27986);
nor U34151 (N_34151,N_25257,N_27334);
nor U34152 (N_34152,N_28388,N_28020);
and U34153 (N_34153,N_26274,N_29990);
nor U34154 (N_34154,N_29892,N_25812);
and U34155 (N_34155,N_29793,N_29594);
and U34156 (N_34156,N_25661,N_25478);
and U34157 (N_34157,N_26578,N_29517);
nand U34158 (N_34158,N_25065,N_25589);
and U34159 (N_34159,N_26342,N_27090);
and U34160 (N_34160,N_25333,N_28617);
or U34161 (N_34161,N_28248,N_26999);
nor U34162 (N_34162,N_28392,N_27610);
nand U34163 (N_34163,N_28499,N_29211);
nor U34164 (N_34164,N_25772,N_25269);
xor U34165 (N_34165,N_28312,N_27118);
xor U34166 (N_34166,N_26818,N_26925);
nand U34167 (N_34167,N_28832,N_26578);
and U34168 (N_34168,N_28342,N_29782);
or U34169 (N_34169,N_26540,N_29513);
nand U34170 (N_34170,N_26515,N_26302);
and U34171 (N_34171,N_26485,N_29628);
nand U34172 (N_34172,N_29847,N_29505);
or U34173 (N_34173,N_26396,N_26628);
xnor U34174 (N_34174,N_29667,N_26488);
nand U34175 (N_34175,N_25460,N_26824);
xor U34176 (N_34176,N_27849,N_27673);
nand U34177 (N_34177,N_29252,N_27994);
xnor U34178 (N_34178,N_28756,N_29194);
or U34179 (N_34179,N_25072,N_27380);
or U34180 (N_34180,N_26895,N_26088);
nand U34181 (N_34181,N_26340,N_25962);
nor U34182 (N_34182,N_29823,N_29909);
nor U34183 (N_34183,N_25582,N_29918);
and U34184 (N_34184,N_25863,N_25704);
and U34185 (N_34185,N_29546,N_28583);
nor U34186 (N_34186,N_27507,N_28936);
nor U34187 (N_34187,N_27984,N_29692);
and U34188 (N_34188,N_26955,N_27059);
or U34189 (N_34189,N_29385,N_25492);
and U34190 (N_34190,N_25299,N_28251);
nor U34191 (N_34191,N_28418,N_27906);
and U34192 (N_34192,N_26802,N_27412);
nand U34193 (N_34193,N_27861,N_26850);
and U34194 (N_34194,N_29576,N_28011);
nand U34195 (N_34195,N_28862,N_29763);
or U34196 (N_34196,N_27128,N_26872);
xnor U34197 (N_34197,N_29856,N_25921);
nand U34198 (N_34198,N_26418,N_25472);
and U34199 (N_34199,N_28406,N_28515);
and U34200 (N_34200,N_26452,N_29545);
nand U34201 (N_34201,N_26286,N_27301);
and U34202 (N_34202,N_29098,N_26507);
or U34203 (N_34203,N_29690,N_28003);
or U34204 (N_34204,N_28776,N_27958);
or U34205 (N_34205,N_29392,N_28115);
nor U34206 (N_34206,N_25366,N_28385);
and U34207 (N_34207,N_29474,N_29012);
and U34208 (N_34208,N_29137,N_26847);
nand U34209 (N_34209,N_25124,N_25421);
and U34210 (N_34210,N_26781,N_26128);
and U34211 (N_34211,N_29542,N_29649);
and U34212 (N_34212,N_25767,N_28520);
nor U34213 (N_34213,N_27802,N_29582);
and U34214 (N_34214,N_29614,N_28346);
and U34215 (N_34215,N_26370,N_25818);
and U34216 (N_34216,N_28389,N_26772);
and U34217 (N_34217,N_29711,N_26596);
or U34218 (N_34218,N_29731,N_26884);
or U34219 (N_34219,N_25800,N_27492);
nand U34220 (N_34220,N_29092,N_27358);
and U34221 (N_34221,N_28264,N_28768);
and U34222 (N_34222,N_25492,N_27869);
nor U34223 (N_34223,N_29798,N_25444);
nand U34224 (N_34224,N_27191,N_26928);
or U34225 (N_34225,N_27186,N_26830);
nor U34226 (N_34226,N_27356,N_25460);
and U34227 (N_34227,N_28192,N_25782);
or U34228 (N_34228,N_27382,N_29758);
or U34229 (N_34229,N_25647,N_29508);
nand U34230 (N_34230,N_29008,N_27775);
or U34231 (N_34231,N_26718,N_28472);
or U34232 (N_34232,N_27938,N_27215);
and U34233 (N_34233,N_27062,N_25222);
nand U34234 (N_34234,N_27991,N_26062);
nor U34235 (N_34235,N_26538,N_25166);
nor U34236 (N_34236,N_25846,N_27927);
nand U34237 (N_34237,N_25486,N_26692);
nand U34238 (N_34238,N_27996,N_29372);
nand U34239 (N_34239,N_29479,N_29555);
nand U34240 (N_34240,N_28415,N_27410);
nand U34241 (N_34241,N_27826,N_27388);
nand U34242 (N_34242,N_28847,N_26276);
or U34243 (N_34243,N_27695,N_27103);
nor U34244 (N_34244,N_28792,N_29850);
nor U34245 (N_34245,N_29958,N_25151);
nor U34246 (N_34246,N_28481,N_27683);
xnor U34247 (N_34247,N_27781,N_27881);
nand U34248 (N_34248,N_26853,N_25300);
nor U34249 (N_34249,N_26011,N_29236);
nand U34250 (N_34250,N_29256,N_28490);
nor U34251 (N_34251,N_29192,N_25581);
or U34252 (N_34252,N_25852,N_28602);
and U34253 (N_34253,N_26980,N_26556);
nand U34254 (N_34254,N_27993,N_25258);
or U34255 (N_34255,N_25999,N_25586);
or U34256 (N_34256,N_27950,N_26393);
and U34257 (N_34257,N_26273,N_27048);
and U34258 (N_34258,N_28616,N_25838);
nor U34259 (N_34259,N_27211,N_27631);
nor U34260 (N_34260,N_28813,N_25393);
and U34261 (N_34261,N_29488,N_26060);
nand U34262 (N_34262,N_27905,N_29162);
and U34263 (N_34263,N_28373,N_29815);
nand U34264 (N_34264,N_28403,N_28370);
nor U34265 (N_34265,N_25426,N_25966);
nand U34266 (N_34266,N_29210,N_28195);
xor U34267 (N_34267,N_27313,N_27486);
nand U34268 (N_34268,N_26346,N_26738);
or U34269 (N_34269,N_28963,N_27438);
and U34270 (N_34270,N_25013,N_28432);
or U34271 (N_34271,N_27134,N_27694);
and U34272 (N_34272,N_28488,N_27554);
or U34273 (N_34273,N_25094,N_25993);
nor U34274 (N_34274,N_26370,N_28162);
nor U34275 (N_34275,N_29731,N_26694);
and U34276 (N_34276,N_28642,N_28465);
and U34277 (N_34277,N_27948,N_27373);
nand U34278 (N_34278,N_25698,N_29823);
nor U34279 (N_34279,N_26474,N_28320);
or U34280 (N_34280,N_27651,N_25249);
nand U34281 (N_34281,N_29021,N_27625);
or U34282 (N_34282,N_25265,N_28890);
or U34283 (N_34283,N_26781,N_27090);
xnor U34284 (N_34284,N_26421,N_28068);
nand U34285 (N_34285,N_29101,N_27778);
nand U34286 (N_34286,N_29991,N_25473);
or U34287 (N_34287,N_29916,N_26793);
or U34288 (N_34288,N_25194,N_27200);
or U34289 (N_34289,N_28072,N_26212);
or U34290 (N_34290,N_25566,N_27514);
and U34291 (N_34291,N_27647,N_29913);
nor U34292 (N_34292,N_28792,N_25381);
nand U34293 (N_34293,N_29773,N_25756);
or U34294 (N_34294,N_28005,N_27775);
nand U34295 (N_34295,N_27834,N_26022);
xor U34296 (N_34296,N_26586,N_27714);
or U34297 (N_34297,N_28054,N_28481);
and U34298 (N_34298,N_25277,N_25157);
nor U34299 (N_34299,N_27265,N_25375);
nor U34300 (N_34300,N_25464,N_28383);
or U34301 (N_34301,N_28755,N_29283);
nor U34302 (N_34302,N_26511,N_29378);
nor U34303 (N_34303,N_28126,N_27644);
and U34304 (N_34304,N_27589,N_25806);
xnor U34305 (N_34305,N_28106,N_27306);
nand U34306 (N_34306,N_28726,N_26301);
and U34307 (N_34307,N_27415,N_25161);
nor U34308 (N_34308,N_25061,N_27713);
nand U34309 (N_34309,N_28629,N_27690);
nor U34310 (N_34310,N_28112,N_25642);
and U34311 (N_34311,N_29721,N_25158);
and U34312 (N_34312,N_26369,N_25653);
or U34313 (N_34313,N_26407,N_29924);
or U34314 (N_34314,N_28722,N_27059);
and U34315 (N_34315,N_28576,N_29874);
nor U34316 (N_34316,N_28464,N_27434);
nor U34317 (N_34317,N_25349,N_29794);
nand U34318 (N_34318,N_29746,N_26704);
xor U34319 (N_34319,N_25659,N_28876);
nor U34320 (N_34320,N_28090,N_29885);
nand U34321 (N_34321,N_28393,N_25627);
nand U34322 (N_34322,N_27547,N_26784);
nor U34323 (N_34323,N_29670,N_29382);
or U34324 (N_34324,N_26665,N_26037);
or U34325 (N_34325,N_28182,N_27867);
or U34326 (N_34326,N_29574,N_25599);
or U34327 (N_34327,N_26034,N_29434);
and U34328 (N_34328,N_27911,N_29559);
nand U34329 (N_34329,N_25019,N_26081);
or U34330 (N_34330,N_25398,N_26809);
xnor U34331 (N_34331,N_26458,N_26585);
nand U34332 (N_34332,N_26318,N_27327);
nand U34333 (N_34333,N_29603,N_28867);
nor U34334 (N_34334,N_27712,N_27628);
nor U34335 (N_34335,N_29135,N_26651);
nor U34336 (N_34336,N_25771,N_26048);
or U34337 (N_34337,N_26654,N_28149);
and U34338 (N_34338,N_25672,N_25353);
or U34339 (N_34339,N_25881,N_29232);
or U34340 (N_34340,N_29599,N_26562);
or U34341 (N_34341,N_26249,N_26578);
or U34342 (N_34342,N_27252,N_28398);
or U34343 (N_34343,N_27545,N_28166);
or U34344 (N_34344,N_29222,N_26162);
and U34345 (N_34345,N_27166,N_26277);
or U34346 (N_34346,N_28413,N_26624);
nand U34347 (N_34347,N_27368,N_29355);
xnor U34348 (N_34348,N_26824,N_27194);
nand U34349 (N_34349,N_27979,N_29112);
or U34350 (N_34350,N_29151,N_26351);
and U34351 (N_34351,N_26992,N_25211);
and U34352 (N_34352,N_28209,N_25225);
and U34353 (N_34353,N_29722,N_28488);
nand U34354 (N_34354,N_29046,N_27457);
or U34355 (N_34355,N_25247,N_26284);
or U34356 (N_34356,N_27527,N_26236);
nor U34357 (N_34357,N_26178,N_26096);
and U34358 (N_34358,N_27893,N_27793);
nor U34359 (N_34359,N_27682,N_26752);
or U34360 (N_34360,N_29116,N_25961);
or U34361 (N_34361,N_27692,N_25614);
nor U34362 (N_34362,N_26725,N_29072);
or U34363 (N_34363,N_26939,N_29903);
xnor U34364 (N_34364,N_29796,N_26198);
and U34365 (N_34365,N_26950,N_29981);
nand U34366 (N_34366,N_26836,N_25299);
nor U34367 (N_34367,N_26899,N_25507);
nor U34368 (N_34368,N_28467,N_28090);
or U34369 (N_34369,N_29954,N_29249);
or U34370 (N_34370,N_27977,N_27897);
or U34371 (N_34371,N_28079,N_29799);
nand U34372 (N_34372,N_29863,N_28151);
and U34373 (N_34373,N_29198,N_28393);
nor U34374 (N_34374,N_25618,N_29632);
and U34375 (N_34375,N_26959,N_25319);
nand U34376 (N_34376,N_26206,N_28986);
nor U34377 (N_34377,N_27725,N_26423);
nor U34378 (N_34378,N_29796,N_28601);
and U34379 (N_34379,N_27594,N_29994);
nor U34380 (N_34380,N_27384,N_27884);
xor U34381 (N_34381,N_28480,N_28578);
nand U34382 (N_34382,N_27873,N_26505);
xor U34383 (N_34383,N_29363,N_25967);
xnor U34384 (N_34384,N_25341,N_28560);
nor U34385 (N_34385,N_25572,N_28427);
nor U34386 (N_34386,N_25407,N_25182);
and U34387 (N_34387,N_27569,N_27907);
nor U34388 (N_34388,N_29451,N_27146);
nor U34389 (N_34389,N_27812,N_25385);
nor U34390 (N_34390,N_25364,N_27635);
nand U34391 (N_34391,N_29647,N_29707);
or U34392 (N_34392,N_25869,N_26867);
nor U34393 (N_34393,N_25828,N_25045);
or U34394 (N_34394,N_26905,N_27668);
nor U34395 (N_34395,N_29805,N_28226);
and U34396 (N_34396,N_29665,N_27404);
nand U34397 (N_34397,N_25621,N_28187);
and U34398 (N_34398,N_27046,N_25908);
nor U34399 (N_34399,N_28740,N_29004);
xor U34400 (N_34400,N_26853,N_28842);
or U34401 (N_34401,N_26734,N_28951);
nand U34402 (N_34402,N_29747,N_29418);
and U34403 (N_34403,N_28066,N_25005);
xor U34404 (N_34404,N_25236,N_29237);
nor U34405 (N_34405,N_27095,N_29702);
and U34406 (N_34406,N_29429,N_26920);
or U34407 (N_34407,N_25178,N_28261);
or U34408 (N_34408,N_28348,N_26474);
or U34409 (N_34409,N_27586,N_26628);
and U34410 (N_34410,N_26910,N_29063);
xnor U34411 (N_34411,N_27769,N_26240);
or U34412 (N_34412,N_27554,N_27997);
xor U34413 (N_34413,N_29733,N_25430);
and U34414 (N_34414,N_26993,N_28530);
nor U34415 (N_34415,N_27508,N_26290);
xor U34416 (N_34416,N_29951,N_25904);
and U34417 (N_34417,N_28348,N_29830);
nand U34418 (N_34418,N_26692,N_29604);
or U34419 (N_34419,N_25440,N_29833);
or U34420 (N_34420,N_27326,N_27488);
nor U34421 (N_34421,N_28196,N_26684);
nand U34422 (N_34422,N_25567,N_25466);
nand U34423 (N_34423,N_26552,N_29301);
nor U34424 (N_34424,N_26148,N_25754);
or U34425 (N_34425,N_27038,N_28586);
or U34426 (N_34426,N_29408,N_27203);
nand U34427 (N_34427,N_28266,N_29235);
nor U34428 (N_34428,N_29313,N_29618);
nand U34429 (N_34429,N_28832,N_28157);
nand U34430 (N_34430,N_26262,N_26874);
nor U34431 (N_34431,N_29982,N_28564);
nor U34432 (N_34432,N_25237,N_26133);
nand U34433 (N_34433,N_26567,N_28097);
or U34434 (N_34434,N_26736,N_29869);
nor U34435 (N_34435,N_27806,N_26958);
xor U34436 (N_34436,N_27157,N_29609);
or U34437 (N_34437,N_27642,N_27959);
nand U34438 (N_34438,N_27771,N_26377);
nand U34439 (N_34439,N_28722,N_28068);
nand U34440 (N_34440,N_26674,N_29662);
nor U34441 (N_34441,N_25090,N_26182);
nand U34442 (N_34442,N_26487,N_26330);
nand U34443 (N_34443,N_25449,N_26173);
and U34444 (N_34444,N_25244,N_27409);
or U34445 (N_34445,N_29144,N_28057);
or U34446 (N_34446,N_26553,N_25923);
or U34447 (N_34447,N_28133,N_27263);
nor U34448 (N_34448,N_25603,N_25985);
nand U34449 (N_34449,N_27915,N_26784);
or U34450 (N_34450,N_29915,N_26583);
nand U34451 (N_34451,N_25556,N_27616);
nand U34452 (N_34452,N_25886,N_25497);
nor U34453 (N_34453,N_25177,N_28017);
nand U34454 (N_34454,N_28699,N_28213);
nand U34455 (N_34455,N_26276,N_28940);
or U34456 (N_34456,N_29074,N_27727);
nand U34457 (N_34457,N_25875,N_27430);
and U34458 (N_34458,N_28055,N_27649);
nand U34459 (N_34459,N_25911,N_26833);
and U34460 (N_34460,N_25543,N_25855);
and U34461 (N_34461,N_27915,N_26325);
nor U34462 (N_34462,N_25539,N_29241);
or U34463 (N_34463,N_29335,N_27235);
or U34464 (N_34464,N_27016,N_29659);
and U34465 (N_34465,N_26109,N_29261);
xor U34466 (N_34466,N_26692,N_29632);
xor U34467 (N_34467,N_28114,N_26243);
nor U34468 (N_34468,N_26731,N_26419);
nand U34469 (N_34469,N_29130,N_26892);
or U34470 (N_34470,N_28399,N_25605);
nor U34471 (N_34471,N_28215,N_25790);
nor U34472 (N_34472,N_28395,N_25518);
nand U34473 (N_34473,N_26032,N_27503);
or U34474 (N_34474,N_26942,N_29088);
nand U34475 (N_34475,N_26679,N_29408);
and U34476 (N_34476,N_27123,N_25118);
nor U34477 (N_34477,N_25707,N_26261);
or U34478 (N_34478,N_25993,N_25923);
and U34479 (N_34479,N_25635,N_29960);
or U34480 (N_34480,N_26071,N_25789);
and U34481 (N_34481,N_28022,N_27501);
nor U34482 (N_34482,N_27374,N_25538);
nor U34483 (N_34483,N_28621,N_28181);
xnor U34484 (N_34484,N_25425,N_28763);
nor U34485 (N_34485,N_27948,N_25075);
or U34486 (N_34486,N_25283,N_27050);
xor U34487 (N_34487,N_25241,N_29787);
and U34488 (N_34488,N_29868,N_28967);
or U34489 (N_34489,N_26096,N_27877);
nand U34490 (N_34490,N_26992,N_27899);
xor U34491 (N_34491,N_28099,N_28568);
and U34492 (N_34492,N_27079,N_25517);
xor U34493 (N_34493,N_29721,N_27227);
nand U34494 (N_34494,N_25139,N_25241);
nand U34495 (N_34495,N_29424,N_28852);
and U34496 (N_34496,N_29358,N_26459);
nor U34497 (N_34497,N_28642,N_25506);
nor U34498 (N_34498,N_29864,N_28103);
nor U34499 (N_34499,N_28493,N_27037);
nand U34500 (N_34500,N_28738,N_29699);
nor U34501 (N_34501,N_28280,N_26316);
nor U34502 (N_34502,N_25534,N_25830);
or U34503 (N_34503,N_25105,N_25669);
nand U34504 (N_34504,N_28033,N_27191);
nand U34505 (N_34505,N_26944,N_25936);
nand U34506 (N_34506,N_29219,N_26906);
nand U34507 (N_34507,N_26299,N_27745);
nand U34508 (N_34508,N_27410,N_26428);
or U34509 (N_34509,N_25330,N_29807);
or U34510 (N_34510,N_28145,N_29073);
nor U34511 (N_34511,N_26222,N_25219);
and U34512 (N_34512,N_26859,N_27730);
nor U34513 (N_34513,N_28273,N_28129);
or U34514 (N_34514,N_28774,N_27177);
or U34515 (N_34515,N_28771,N_27183);
and U34516 (N_34516,N_26247,N_27931);
or U34517 (N_34517,N_27891,N_26255);
xnor U34518 (N_34518,N_29292,N_25282);
nand U34519 (N_34519,N_29463,N_27861);
nand U34520 (N_34520,N_29281,N_29990);
or U34521 (N_34521,N_26993,N_29392);
nand U34522 (N_34522,N_28893,N_26971);
or U34523 (N_34523,N_29970,N_26726);
nand U34524 (N_34524,N_27696,N_27085);
nand U34525 (N_34525,N_26672,N_27207);
nor U34526 (N_34526,N_29179,N_26491);
and U34527 (N_34527,N_27250,N_27785);
or U34528 (N_34528,N_26813,N_29439);
or U34529 (N_34529,N_26882,N_29191);
xnor U34530 (N_34530,N_25168,N_29537);
and U34531 (N_34531,N_26350,N_27157);
or U34532 (N_34532,N_29721,N_29450);
xor U34533 (N_34533,N_27666,N_27151);
xor U34534 (N_34534,N_27614,N_28266);
nand U34535 (N_34535,N_27926,N_27700);
nand U34536 (N_34536,N_28576,N_26029);
or U34537 (N_34537,N_28661,N_26702);
or U34538 (N_34538,N_27122,N_29749);
nand U34539 (N_34539,N_25946,N_25969);
and U34540 (N_34540,N_28546,N_29898);
nand U34541 (N_34541,N_28774,N_29357);
or U34542 (N_34542,N_28437,N_27407);
and U34543 (N_34543,N_27381,N_26486);
or U34544 (N_34544,N_28854,N_29580);
xnor U34545 (N_34545,N_26117,N_29341);
nor U34546 (N_34546,N_29291,N_27780);
nor U34547 (N_34547,N_25910,N_25833);
nor U34548 (N_34548,N_27214,N_25917);
or U34549 (N_34549,N_28974,N_29216);
and U34550 (N_34550,N_27395,N_25344);
and U34551 (N_34551,N_29735,N_25260);
and U34552 (N_34552,N_29474,N_26990);
and U34553 (N_34553,N_27589,N_26099);
nand U34554 (N_34554,N_26875,N_29133);
or U34555 (N_34555,N_26700,N_25222);
or U34556 (N_34556,N_28150,N_28072);
and U34557 (N_34557,N_27278,N_27084);
xnor U34558 (N_34558,N_28181,N_28666);
nand U34559 (N_34559,N_28579,N_25511);
and U34560 (N_34560,N_27073,N_25660);
nand U34561 (N_34561,N_29119,N_27897);
nor U34562 (N_34562,N_28608,N_25371);
nor U34563 (N_34563,N_26709,N_28824);
xnor U34564 (N_34564,N_29148,N_25060);
or U34565 (N_34565,N_25845,N_25354);
xor U34566 (N_34566,N_26776,N_25844);
nand U34567 (N_34567,N_28471,N_29067);
nand U34568 (N_34568,N_28986,N_25346);
and U34569 (N_34569,N_28435,N_25815);
xor U34570 (N_34570,N_29999,N_28747);
or U34571 (N_34571,N_25839,N_28558);
and U34572 (N_34572,N_26528,N_27722);
nor U34573 (N_34573,N_25510,N_29684);
or U34574 (N_34574,N_28719,N_28834);
and U34575 (N_34575,N_29094,N_29160);
nand U34576 (N_34576,N_27819,N_25982);
or U34577 (N_34577,N_27636,N_28045);
nor U34578 (N_34578,N_28532,N_25275);
nor U34579 (N_34579,N_29868,N_29257);
and U34580 (N_34580,N_27148,N_28787);
nand U34581 (N_34581,N_26748,N_26003);
or U34582 (N_34582,N_27386,N_27460);
nand U34583 (N_34583,N_25379,N_25313);
nand U34584 (N_34584,N_28206,N_26002);
nand U34585 (N_34585,N_27371,N_29025);
xor U34586 (N_34586,N_28884,N_29707);
nand U34587 (N_34587,N_26941,N_25957);
xor U34588 (N_34588,N_25456,N_29766);
nor U34589 (N_34589,N_29485,N_26017);
and U34590 (N_34590,N_26687,N_29066);
and U34591 (N_34591,N_27645,N_25164);
and U34592 (N_34592,N_29035,N_27465);
nand U34593 (N_34593,N_29690,N_25565);
nor U34594 (N_34594,N_27038,N_27456);
and U34595 (N_34595,N_27801,N_28090);
nor U34596 (N_34596,N_27033,N_27267);
and U34597 (N_34597,N_29406,N_27733);
or U34598 (N_34598,N_29656,N_26777);
or U34599 (N_34599,N_29921,N_29840);
nand U34600 (N_34600,N_25335,N_28258);
nand U34601 (N_34601,N_27499,N_27509);
nand U34602 (N_34602,N_25655,N_26238);
xnor U34603 (N_34603,N_25704,N_27101);
and U34604 (N_34604,N_27353,N_25457);
nand U34605 (N_34605,N_28878,N_29588);
or U34606 (N_34606,N_25138,N_28726);
and U34607 (N_34607,N_29304,N_25083);
nand U34608 (N_34608,N_28434,N_27076);
nand U34609 (N_34609,N_27578,N_27751);
and U34610 (N_34610,N_28298,N_25246);
or U34611 (N_34611,N_29782,N_29981);
nand U34612 (N_34612,N_27022,N_28054);
nor U34613 (N_34613,N_28681,N_25413);
nor U34614 (N_34614,N_25650,N_26714);
and U34615 (N_34615,N_28751,N_27552);
or U34616 (N_34616,N_28181,N_26231);
or U34617 (N_34617,N_26221,N_25912);
or U34618 (N_34618,N_26780,N_26775);
nor U34619 (N_34619,N_28680,N_26843);
nand U34620 (N_34620,N_27789,N_26693);
nor U34621 (N_34621,N_25604,N_28148);
nor U34622 (N_34622,N_25040,N_27974);
and U34623 (N_34623,N_25863,N_27099);
and U34624 (N_34624,N_28186,N_26951);
xnor U34625 (N_34625,N_26563,N_29757);
nor U34626 (N_34626,N_26573,N_25598);
and U34627 (N_34627,N_25273,N_28216);
nor U34628 (N_34628,N_25869,N_25360);
and U34629 (N_34629,N_28680,N_29984);
nor U34630 (N_34630,N_27730,N_25333);
and U34631 (N_34631,N_25849,N_25893);
nand U34632 (N_34632,N_27284,N_26745);
and U34633 (N_34633,N_28120,N_26234);
and U34634 (N_34634,N_27311,N_27467);
or U34635 (N_34635,N_26012,N_27316);
nor U34636 (N_34636,N_25201,N_29379);
or U34637 (N_34637,N_27373,N_25256);
xnor U34638 (N_34638,N_27880,N_26339);
nor U34639 (N_34639,N_25661,N_29083);
nand U34640 (N_34640,N_27093,N_29604);
and U34641 (N_34641,N_27597,N_25850);
nor U34642 (N_34642,N_28077,N_29288);
or U34643 (N_34643,N_27466,N_26694);
or U34644 (N_34644,N_27469,N_28731);
or U34645 (N_34645,N_27740,N_25839);
or U34646 (N_34646,N_29186,N_29448);
xnor U34647 (N_34647,N_27776,N_25836);
nor U34648 (N_34648,N_27878,N_29050);
nor U34649 (N_34649,N_27704,N_29994);
or U34650 (N_34650,N_29268,N_29388);
xor U34651 (N_34651,N_28545,N_29782);
and U34652 (N_34652,N_29907,N_25839);
and U34653 (N_34653,N_25761,N_26803);
nor U34654 (N_34654,N_27271,N_26490);
or U34655 (N_34655,N_25205,N_28599);
and U34656 (N_34656,N_26764,N_28166);
or U34657 (N_34657,N_25212,N_26373);
nor U34658 (N_34658,N_25751,N_29488);
or U34659 (N_34659,N_28576,N_25957);
nand U34660 (N_34660,N_26209,N_27227);
or U34661 (N_34661,N_27801,N_28805);
nand U34662 (N_34662,N_29419,N_27333);
nand U34663 (N_34663,N_27802,N_29342);
nand U34664 (N_34664,N_28013,N_25211);
or U34665 (N_34665,N_25092,N_26883);
nand U34666 (N_34666,N_28280,N_27778);
xnor U34667 (N_34667,N_26051,N_26764);
or U34668 (N_34668,N_26150,N_25075);
or U34669 (N_34669,N_27045,N_29719);
nor U34670 (N_34670,N_29799,N_25512);
nor U34671 (N_34671,N_27307,N_25664);
nand U34672 (N_34672,N_25491,N_28143);
nand U34673 (N_34673,N_29367,N_28885);
xnor U34674 (N_34674,N_27415,N_26634);
nor U34675 (N_34675,N_28173,N_27503);
xor U34676 (N_34676,N_25511,N_26545);
or U34677 (N_34677,N_28224,N_29857);
nand U34678 (N_34678,N_25230,N_28026);
and U34679 (N_34679,N_29244,N_26099);
nand U34680 (N_34680,N_25914,N_28414);
nand U34681 (N_34681,N_28054,N_25454);
or U34682 (N_34682,N_29920,N_26459);
nor U34683 (N_34683,N_29371,N_28255);
nor U34684 (N_34684,N_29216,N_28770);
or U34685 (N_34685,N_26455,N_25932);
or U34686 (N_34686,N_27275,N_29429);
or U34687 (N_34687,N_29255,N_26479);
and U34688 (N_34688,N_29123,N_27158);
and U34689 (N_34689,N_29586,N_26851);
xnor U34690 (N_34690,N_27260,N_26767);
nor U34691 (N_34691,N_28877,N_28988);
nor U34692 (N_34692,N_29419,N_28277);
xnor U34693 (N_34693,N_26615,N_27788);
xor U34694 (N_34694,N_29273,N_25733);
or U34695 (N_34695,N_28142,N_25720);
xor U34696 (N_34696,N_27586,N_26539);
and U34697 (N_34697,N_29508,N_25708);
and U34698 (N_34698,N_25913,N_28986);
or U34699 (N_34699,N_29945,N_26319);
nor U34700 (N_34700,N_28839,N_29417);
xor U34701 (N_34701,N_27685,N_25449);
nor U34702 (N_34702,N_27305,N_26044);
and U34703 (N_34703,N_25561,N_26052);
and U34704 (N_34704,N_29595,N_29500);
nor U34705 (N_34705,N_29362,N_25464);
and U34706 (N_34706,N_28525,N_26000);
nor U34707 (N_34707,N_27561,N_29896);
or U34708 (N_34708,N_27539,N_29152);
or U34709 (N_34709,N_25460,N_27153);
or U34710 (N_34710,N_28380,N_29440);
or U34711 (N_34711,N_29644,N_29301);
nor U34712 (N_34712,N_27261,N_27214);
nor U34713 (N_34713,N_26961,N_28248);
or U34714 (N_34714,N_25330,N_28819);
nand U34715 (N_34715,N_25345,N_25047);
and U34716 (N_34716,N_26848,N_27885);
or U34717 (N_34717,N_27621,N_28001);
xor U34718 (N_34718,N_29842,N_27282);
nor U34719 (N_34719,N_26027,N_28779);
or U34720 (N_34720,N_25872,N_25098);
xor U34721 (N_34721,N_25079,N_26000);
or U34722 (N_34722,N_26671,N_25315);
xor U34723 (N_34723,N_26397,N_25518);
nand U34724 (N_34724,N_27215,N_29416);
nand U34725 (N_34725,N_28849,N_25714);
nand U34726 (N_34726,N_29761,N_26661);
xor U34727 (N_34727,N_29011,N_29715);
or U34728 (N_34728,N_28318,N_27572);
or U34729 (N_34729,N_28163,N_26514);
nor U34730 (N_34730,N_29678,N_27107);
nor U34731 (N_34731,N_26881,N_29790);
and U34732 (N_34732,N_25177,N_26126);
nand U34733 (N_34733,N_28181,N_29345);
and U34734 (N_34734,N_29624,N_25955);
nor U34735 (N_34735,N_25756,N_25183);
and U34736 (N_34736,N_29616,N_25151);
nand U34737 (N_34737,N_27192,N_29971);
nand U34738 (N_34738,N_26839,N_29046);
nand U34739 (N_34739,N_27408,N_27399);
nand U34740 (N_34740,N_25810,N_27052);
nor U34741 (N_34741,N_26563,N_26110);
nand U34742 (N_34742,N_29942,N_26030);
nor U34743 (N_34743,N_29454,N_28273);
and U34744 (N_34744,N_25142,N_27605);
or U34745 (N_34745,N_28520,N_27041);
nor U34746 (N_34746,N_28821,N_26555);
and U34747 (N_34747,N_25424,N_26197);
or U34748 (N_34748,N_29408,N_29196);
nor U34749 (N_34749,N_26838,N_25636);
nor U34750 (N_34750,N_29702,N_27568);
nor U34751 (N_34751,N_26179,N_26007);
or U34752 (N_34752,N_28607,N_29913);
nor U34753 (N_34753,N_28545,N_25725);
nand U34754 (N_34754,N_27550,N_28601);
and U34755 (N_34755,N_29813,N_27014);
xnor U34756 (N_34756,N_29089,N_28476);
and U34757 (N_34757,N_25547,N_26560);
nand U34758 (N_34758,N_28739,N_29942);
or U34759 (N_34759,N_25835,N_26421);
nor U34760 (N_34760,N_29006,N_29954);
nor U34761 (N_34761,N_26759,N_29428);
and U34762 (N_34762,N_26691,N_26031);
nand U34763 (N_34763,N_27035,N_26452);
nor U34764 (N_34764,N_29123,N_28410);
xnor U34765 (N_34765,N_29763,N_26368);
nor U34766 (N_34766,N_29024,N_27222);
nand U34767 (N_34767,N_27804,N_28285);
or U34768 (N_34768,N_26470,N_29390);
nand U34769 (N_34769,N_29803,N_28274);
or U34770 (N_34770,N_26877,N_28210);
nor U34771 (N_34771,N_27404,N_27645);
nor U34772 (N_34772,N_25318,N_26888);
or U34773 (N_34773,N_26399,N_25581);
and U34774 (N_34774,N_29909,N_26311);
nand U34775 (N_34775,N_28395,N_29698);
nor U34776 (N_34776,N_26137,N_25184);
or U34777 (N_34777,N_26471,N_25821);
or U34778 (N_34778,N_26024,N_26327);
and U34779 (N_34779,N_27357,N_25046);
and U34780 (N_34780,N_27719,N_25634);
or U34781 (N_34781,N_28706,N_29317);
nand U34782 (N_34782,N_26518,N_25217);
nand U34783 (N_34783,N_25556,N_26658);
nor U34784 (N_34784,N_28031,N_29716);
nor U34785 (N_34785,N_28348,N_27726);
nor U34786 (N_34786,N_29905,N_28876);
and U34787 (N_34787,N_27586,N_29339);
nor U34788 (N_34788,N_25328,N_25768);
nor U34789 (N_34789,N_28577,N_27913);
nand U34790 (N_34790,N_28729,N_28907);
xnor U34791 (N_34791,N_29071,N_25962);
or U34792 (N_34792,N_27335,N_28639);
or U34793 (N_34793,N_26715,N_26360);
nand U34794 (N_34794,N_29035,N_26205);
xnor U34795 (N_34795,N_27095,N_27346);
and U34796 (N_34796,N_26182,N_26135);
nand U34797 (N_34797,N_26738,N_29035);
or U34798 (N_34798,N_26598,N_25739);
nor U34799 (N_34799,N_28388,N_27041);
or U34800 (N_34800,N_25461,N_28763);
or U34801 (N_34801,N_25045,N_27939);
or U34802 (N_34802,N_29579,N_27547);
and U34803 (N_34803,N_28579,N_27355);
or U34804 (N_34804,N_26234,N_28909);
and U34805 (N_34805,N_26218,N_26757);
nor U34806 (N_34806,N_28331,N_28157);
xor U34807 (N_34807,N_29179,N_26035);
and U34808 (N_34808,N_27918,N_26393);
and U34809 (N_34809,N_29195,N_28166);
nand U34810 (N_34810,N_26690,N_26075);
nand U34811 (N_34811,N_26758,N_25650);
or U34812 (N_34812,N_25470,N_27150);
nor U34813 (N_34813,N_28488,N_27740);
xnor U34814 (N_34814,N_25379,N_28737);
nor U34815 (N_34815,N_29315,N_26255);
and U34816 (N_34816,N_29800,N_25343);
and U34817 (N_34817,N_26188,N_25850);
nor U34818 (N_34818,N_29761,N_28125);
nor U34819 (N_34819,N_29416,N_25176);
nor U34820 (N_34820,N_25220,N_27607);
nand U34821 (N_34821,N_29428,N_26002);
nand U34822 (N_34822,N_25006,N_27024);
nand U34823 (N_34823,N_25493,N_28567);
nand U34824 (N_34824,N_25813,N_29557);
nor U34825 (N_34825,N_29690,N_29237);
xor U34826 (N_34826,N_25123,N_26212);
nand U34827 (N_34827,N_28245,N_27175);
xnor U34828 (N_34828,N_25444,N_26538);
nor U34829 (N_34829,N_27860,N_29856);
or U34830 (N_34830,N_25421,N_26941);
and U34831 (N_34831,N_26905,N_28264);
nand U34832 (N_34832,N_27263,N_28601);
nand U34833 (N_34833,N_25941,N_26563);
nor U34834 (N_34834,N_27316,N_27366);
and U34835 (N_34835,N_28211,N_25263);
nand U34836 (N_34836,N_27226,N_29415);
or U34837 (N_34837,N_26044,N_29957);
nor U34838 (N_34838,N_27881,N_26953);
or U34839 (N_34839,N_26935,N_25039);
or U34840 (N_34840,N_29953,N_29691);
nand U34841 (N_34841,N_27020,N_28955);
or U34842 (N_34842,N_27350,N_28345);
nand U34843 (N_34843,N_25511,N_26316);
and U34844 (N_34844,N_29785,N_29399);
and U34845 (N_34845,N_27374,N_28787);
or U34846 (N_34846,N_28902,N_26906);
nand U34847 (N_34847,N_29489,N_28189);
or U34848 (N_34848,N_27009,N_26152);
nand U34849 (N_34849,N_27318,N_29883);
nand U34850 (N_34850,N_29981,N_25999);
nor U34851 (N_34851,N_27435,N_29070);
nor U34852 (N_34852,N_27177,N_26369);
and U34853 (N_34853,N_25925,N_26785);
xnor U34854 (N_34854,N_29799,N_27481);
nand U34855 (N_34855,N_25753,N_26080);
or U34856 (N_34856,N_28374,N_27460);
nand U34857 (N_34857,N_28633,N_26156);
nor U34858 (N_34858,N_29800,N_26287);
and U34859 (N_34859,N_28654,N_25323);
nor U34860 (N_34860,N_29994,N_29769);
or U34861 (N_34861,N_25817,N_25522);
nor U34862 (N_34862,N_28389,N_27367);
or U34863 (N_34863,N_26046,N_26015);
xnor U34864 (N_34864,N_29171,N_29961);
nand U34865 (N_34865,N_29110,N_28616);
nand U34866 (N_34866,N_28938,N_28196);
nand U34867 (N_34867,N_28868,N_27448);
nand U34868 (N_34868,N_29408,N_27627);
nand U34869 (N_34869,N_27028,N_29072);
nand U34870 (N_34870,N_27607,N_26672);
nand U34871 (N_34871,N_28032,N_25947);
nand U34872 (N_34872,N_27440,N_29842);
and U34873 (N_34873,N_29174,N_29024);
or U34874 (N_34874,N_28493,N_28954);
nand U34875 (N_34875,N_29530,N_27725);
xnor U34876 (N_34876,N_25403,N_26615);
or U34877 (N_34877,N_28792,N_25231);
xnor U34878 (N_34878,N_25067,N_25468);
or U34879 (N_34879,N_28306,N_25791);
nor U34880 (N_34880,N_28717,N_26351);
and U34881 (N_34881,N_26206,N_28050);
or U34882 (N_34882,N_27395,N_27193);
and U34883 (N_34883,N_29644,N_29312);
nor U34884 (N_34884,N_28581,N_26180);
nand U34885 (N_34885,N_29614,N_29051);
nand U34886 (N_34886,N_27289,N_26869);
nand U34887 (N_34887,N_27354,N_28792);
nor U34888 (N_34888,N_27769,N_29423);
nand U34889 (N_34889,N_27832,N_26853);
and U34890 (N_34890,N_29796,N_25995);
or U34891 (N_34891,N_26797,N_27192);
nor U34892 (N_34892,N_25983,N_25659);
and U34893 (N_34893,N_27910,N_28830);
nand U34894 (N_34894,N_25211,N_26693);
nor U34895 (N_34895,N_28823,N_29773);
or U34896 (N_34896,N_26594,N_29967);
and U34897 (N_34897,N_26357,N_29170);
and U34898 (N_34898,N_26776,N_26502);
nand U34899 (N_34899,N_25365,N_27495);
and U34900 (N_34900,N_26396,N_25704);
xor U34901 (N_34901,N_28797,N_26634);
nor U34902 (N_34902,N_25183,N_27382);
nor U34903 (N_34903,N_26033,N_27332);
nand U34904 (N_34904,N_28343,N_29631);
nand U34905 (N_34905,N_28075,N_26160);
and U34906 (N_34906,N_27969,N_27877);
nand U34907 (N_34907,N_29775,N_25183);
nor U34908 (N_34908,N_28275,N_28595);
nand U34909 (N_34909,N_25739,N_29178);
nor U34910 (N_34910,N_26441,N_25282);
xnor U34911 (N_34911,N_25574,N_27284);
or U34912 (N_34912,N_28203,N_25251);
or U34913 (N_34913,N_26093,N_29983);
and U34914 (N_34914,N_25376,N_28660);
nor U34915 (N_34915,N_27451,N_25887);
and U34916 (N_34916,N_27099,N_29020);
nor U34917 (N_34917,N_29099,N_26132);
xnor U34918 (N_34918,N_27881,N_27134);
nor U34919 (N_34919,N_27905,N_26812);
nand U34920 (N_34920,N_28389,N_26400);
and U34921 (N_34921,N_27234,N_27500);
nor U34922 (N_34922,N_29541,N_28256);
nor U34923 (N_34923,N_28654,N_26078);
nand U34924 (N_34924,N_28639,N_28939);
or U34925 (N_34925,N_27802,N_29983);
nor U34926 (N_34926,N_25133,N_29412);
nand U34927 (N_34927,N_28139,N_28419);
and U34928 (N_34928,N_26627,N_27087);
nor U34929 (N_34929,N_29406,N_26331);
nand U34930 (N_34930,N_26056,N_26770);
nor U34931 (N_34931,N_25293,N_27509);
nor U34932 (N_34932,N_28390,N_26796);
nand U34933 (N_34933,N_26765,N_27541);
xnor U34934 (N_34934,N_25942,N_29659);
nor U34935 (N_34935,N_29671,N_29404);
nor U34936 (N_34936,N_29897,N_26453);
and U34937 (N_34937,N_29580,N_27228);
nor U34938 (N_34938,N_27849,N_29655);
and U34939 (N_34939,N_27789,N_29394);
or U34940 (N_34940,N_29966,N_27882);
and U34941 (N_34941,N_29436,N_25040);
and U34942 (N_34942,N_29920,N_26992);
nor U34943 (N_34943,N_26382,N_25577);
nor U34944 (N_34944,N_28479,N_25579);
nand U34945 (N_34945,N_26012,N_28192);
xor U34946 (N_34946,N_25020,N_28922);
xor U34947 (N_34947,N_28269,N_26283);
and U34948 (N_34948,N_26769,N_25181);
and U34949 (N_34949,N_28017,N_28880);
nand U34950 (N_34950,N_28483,N_27952);
xor U34951 (N_34951,N_28668,N_26352);
nor U34952 (N_34952,N_26340,N_25451);
nor U34953 (N_34953,N_27891,N_28650);
nor U34954 (N_34954,N_27588,N_27771);
or U34955 (N_34955,N_28005,N_26487);
nand U34956 (N_34956,N_29764,N_28059);
nand U34957 (N_34957,N_27713,N_25776);
nand U34958 (N_34958,N_28707,N_29142);
xnor U34959 (N_34959,N_28219,N_25694);
xor U34960 (N_34960,N_29307,N_28805);
and U34961 (N_34961,N_26107,N_27782);
xnor U34962 (N_34962,N_27395,N_26424);
or U34963 (N_34963,N_27563,N_26346);
and U34964 (N_34964,N_27681,N_28158);
nand U34965 (N_34965,N_29129,N_27046);
xor U34966 (N_34966,N_25935,N_29987);
or U34967 (N_34967,N_29366,N_28090);
or U34968 (N_34968,N_25334,N_27768);
nand U34969 (N_34969,N_25016,N_25157);
and U34970 (N_34970,N_27966,N_28302);
nor U34971 (N_34971,N_26918,N_27762);
and U34972 (N_34972,N_27068,N_27615);
or U34973 (N_34973,N_28348,N_29095);
and U34974 (N_34974,N_25676,N_27026);
or U34975 (N_34975,N_25529,N_27754);
or U34976 (N_34976,N_25563,N_28875);
nor U34977 (N_34977,N_27376,N_28397);
nor U34978 (N_34978,N_25166,N_29511);
and U34979 (N_34979,N_26103,N_26690);
nor U34980 (N_34980,N_26149,N_25463);
nor U34981 (N_34981,N_25501,N_27379);
or U34982 (N_34982,N_27827,N_27397);
and U34983 (N_34983,N_29522,N_29323);
nand U34984 (N_34984,N_29031,N_28960);
nor U34985 (N_34985,N_28204,N_28531);
nand U34986 (N_34986,N_28745,N_26717);
nand U34987 (N_34987,N_27270,N_28982);
or U34988 (N_34988,N_27536,N_27106);
nand U34989 (N_34989,N_28878,N_26687);
and U34990 (N_34990,N_25862,N_29490);
nor U34991 (N_34991,N_29719,N_27197);
nor U34992 (N_34992,N_29355,N_25612);
and U34993 (N_34993,N_25410,N_28630);
and U34994 (N_34994,N_28413,N_26485);
xor U34995 (N_34995,N_28021,N_26612);
nor U34996 (N_34996,N_27314,N_27287);
nor U34997 (N_34997,N_27410,N_26779);
and U34998 (N_34998,N_28149,N_27404);
or U34999 (N_34999,N_26927,N_26131);
or U35000 (N_35000,N_31136,N_30686);
and U35001 (N_35001,N_30697,N_32533);
and U35002 (N_35002,N_30738,N_32849);
and U35003 (N_35003,N_32943,N_31133);
and U35004 (N_35004,N_33371,N_32615);
nand U35005 (N_35005,N_33545,N_33353);
nor U35006 (N_35006,N_34617,N_31478);
nor U35007 (N_35007,N_33413,N_31703);
nand U35008 (N_35008,N_33027,N_32569);
nor U35009 (N_35009,N_31956,N_33290);
or U35010 (N_35010,N_33737,N_31752);
nand U35011 (N_35011,N_34881,N_31104);
or U35012 (N_35012,N_34250,N_30799);
xnor U35013 (N_35013,N_33018,N_34020);
or U35014 (N_35014,N_30129,N_30871);
nor U35015 (N_35015,N_30107,N_34720);
nand U35016 (N_35016,N_34191,N_33478);
nand U35017 (N_35017,N_32237,N_31692);
and U35018 (N_35018,N_32499,N_31489);
and U35019 (N_35019,N_33632,N_34423);
or U35020 (N_35020,N_31100,N_31357);
nand U35021 (N_35021,N_30419,N_31240);
nand U35022 (N_35022,N_31823,N_30263);
nand U35023 (N_35023,N_34450,N_30148);
nand U35024 (N_35024,N_34736,N_32609);
and U35025 (N_35025,N_32730,N_32116);
or U35026 (N_35026,N_32565,N_33655);
nand U35027 (N_35027,N_33380,N_33664);
and U35028 (N_35028,N_31948,N_32011);
or U35029 (N_35029,N_33301,N_33641);
nor U35030 (N_35030,N_32786,N_34282);
or U35031 (N_35031,N_34811,N_33317);
or U35032 (N_35032,N_30549,N_33976);
nand U35033 (N_35033,N_31922,N_30638);
or U35034 (N_35034,N_30334,N_32694);
xor U35035 (N_35035,N_34383,N_34448);
or U35036 (N_35036,N_30389,N_30545);
nor U35037 (N_35037,N_33697,N_32660);
or U35038 (N_35038,N_34748,N_34793);
nor U35039 (N_35039,N_32277,N_31343);
or U35040 (N_35040,N_31095,N_32206);
nor U35041 (N_35041,N_34552,N_32434);
xor U35042 (N_35042,N_30772,N_31660);
and U35043 (N_35043,N_30702,N_31869);
nor U35044 (N_35044,N_32739,N_32412);
or U35045 (N_35045,N_34828,N_34016);
nand U35046 (N_35046,N_31113,N_33077);
or U35047 (N_35047,N_31535,N_32852);
xnor U35048 (N_35048,N_34396,N_31889);
nor U35049 (N_35049,N_30297,N_33538);
nand U35050 (N_35050,N_34353,N_34724);
nand U35051 (N_35051,N_34006,N_30171);
xor U35052 (N_35052,N_33695,N_34208);
or U35053 (N_35053,N_33856,N_30916);
nand U35054 (N_35054,N_31757,N_32029);
nand U35055 (N_35055,N_30596,N_34005);
or U35056 (N_35056,N_30059,N_33091);
nand U35057 (N_35057,N_33034,N_32126);
and U35058 (N_35058,N_32491,N_33733);
nand U35059 (N_35059,N_34656,N_31025);
nor U35060 (N_35060,N_34659,N_31052);
nor U35061 (N_35061,N_34473,N_34510);
or U35062 (N_35062,N_30377,N_31754);
and U35063 (N_35063,N_31542,N_31718);
and U35064 (N_35064,N_34360,N_31039);
nor U35065 (N_35065,N_32428,N_31521);
or U35066 (N_35066,N_33565,N_33765);
nand U35067 (N_35067,N_32610,N_31992);
xnor U35068 (N_35068,N_33523,N_31065);
and U35069 (N_35069,N_33728,N_31828);
and U35070 (N_35070,N_34327,N_31932);
nand U35071 (N_35071,N_33602,N_33908);
xnor U35072 (N_35072,N_30904,N_31780);
nor U35073 (N_35073,N_33834,N_34575);
nand U35074 (N_35074,N_30711,N_32360);
nor U35075 (N_35075,N_30058,N_31014);
nor U35076 (N_35076,N_32181,N_32706);
or U35077 (N_35077,N_34251,N_32909);
nor U35078 (N_35078,N_31848,N_31022);
nand U35079 (N_35079,N_34574,N_34664);
nor U35080 (N_35080,N_30458,N_34771);
nor U35081 (N_35081,N_31677,N_31775);
nor U35082 (N_35082,N_31782,N_33512);
or U35083 (N_35083,N_32151,N_30622);
or U35084 (N_35084,N_33012,N_33485);
nand U35085 (N_35085,N_34606,N_31387);
and U35086 (N_35086,N_32732,N_32130);
nor U35087 (N_35087,N_31329,N_30812);
nand U35088 (N_35088,N_32966,N_30854);
nor U35089 (N_35089,N_30816,N_33238);
or U35090 (N_35090,N_30558,N_30557);
or U35091 (N_35091,N_34760,N_30552);
and U35092 (N_35092,N_31189,N_31410);
and U35093 (N_35093,N_30019,N_32562);
and U35094 (N_35094,N_31833,N_33584);
and U35095 (N_35095,N_32983,N_31227);
xnor U35096 (N_35096,N_32702,N_33937);
nand U35097 (N_35097,N_34807,N_33610);
nand U35098 (N_35098,N_34857,N_32088);
or U35099 (N_35099,N_30333,N_34121);
or U35100 (N_35100,N_34496,N_34925);
and U35101 (N_35101,N_34728,N_30137);
or U35102 (N_35102,N_30996,N_32655);
and U35103 (N_35103,N_32362,N_30763);
nor U35104 (N_35104,N_30039,N_34799);
nand U35105 (N_35105,N_31352,N_34050);
nor U35106 (N_35106,N_30230,N_34745);
nand U35107 (N_35107,N_30994,N_31510);
nand U35108 (N_35108,N_32717,N_33275);
and U35109 (N_35109,N_31683,N_33045);
or U35110 (N_35110,N_30791,N_34902);
xor U35111 (N_35111,N_30840,N_34900);
or U35112 (N_35112,N_33055,N_32023);
nor U35113 (N_35113,N_31438,N_31205);
nor U35114 (N_35114,N_33237,N_34788);
and U35115 (N_35115,N_34822,N_31667);
and U35116 (N_35116,N_32234,N_33945);
nand U35117 (N_35117,N_32244,N_31617);
nor U35118 (N_35118,N_31508,N_32723);
xor U35119 (N_35119,N_32440,N_30864);
nor U35120 (N_35120,N_34403,N_33986);
nor U35121 (N_35121,N_34183,N_32210);
and U35122 (N_35122,N_30568,N_34668);
and U35123 (N_35123,N_33374,N_31358);
nor U35124 (N_35124,N_32289,N_31336);
nand U35125 (N_35125,N_33760,N_31169);
or U35126 (N_35126,N_32322,N_33252);
nor U35127 (N_35127,N_33137,N_34233);
nand U35128 (N_35128,N_31525,N_34585);
and U35129 (N_35129,N_31470,N_31746);
nor U35130 (N_35130,N_31193,N_30834);
or U35131 (N_35131,N_33016,N_32646);
nand U35132 (N_35132,N_32871,N_31821);
or U35133 (N_35133,N_34619,N_33759);
xor U35134 (N_35134,N_33764,N_33284);
nand U35135 (N_35135,N_34068,N_33344);
and U35136 (N_35136,N_30980,N_32245);
xor U35137 (N_35137,N_32182,N_31209);
and U35138 (N_35138,N_30349,N_31079);
nand U35139 (N_35139,N_34297,N_30586);
nand U35140 (N_35140,N_33339,N_34901);
and U35141 (N_35141,N_30920,N_33516);
nand U35142 (N_35142,N_31023,N_30538);
nor U35143 (N_35143,N_34161,N_33044);
or U35144 (N_35144,N_30353,N_30633);
or U35145 (N_35145,N_32999,N_33241);
or U35146 (N_35146,N_31504,N_30838);
and U35147 (N_35147,N_30135,N_30153);
nor U35148 (N_35148,N_31765,N_34678);
nand U35149 (N_35149,N_31618,N_34313);
and U35150 (N_35150,N_30560,N_33308);
nand U35151 (N_35151,N_32617,N_33517);
and U35152 (N_35152,N_34727,N_30508);
and U35153 (N_35153,N_30704,N_32453);
xor U35154 (N_35154,N_33551,N_31407);
or U35155 (N_35155,N_32806,N_33779);
and U35156 (N_35156,N_30530,N_33209);
xnor U35157 (N_35157,N_34525,N_30806);
nand U35158 (N_35158,N_32349,N_33164);
or U35159 (N_35159,N_30144,N_32875);
and U35160 (N_35160,N_33390,N_33983);
xor U35161 (N_35161,N_33453,N_33117);
xor U35162 (N_35162,N_33305,N_32633);
and U35163 (N_35163,N_34468,N_31480);
or U35164 (N_35164,N_32675,N_34498);
nand U35165 (N_35165,N_33744,N_32663);
nand U35166 (N_35166,N_33178,N_33287);
nor U35167 (N_35167,N_33500,N_30793);
xor U35168 (N_35168,N_31653,N_33393);
xor U35169 (N_35169,N_31993,N_33685);
nand U35170 (N_35170,N_34349,N_33964);
and U35171 (N_35171,N_31006,N_32632);
and U35172 (N_35172,N_32055,N_32900);
or U35173 (N_35173,N_34862,N_32910);
nor U35174 (N_35174,N_30173,N_34260);
or U35175 (N_35175,N_32197,N_30052);
nand U35176 (N_35176,N_30490,N_33680);
nand U35177 (N_35177,N_30522,N_31488);
nor U35178 (N_35178,N_30161,N_31225);
and U35179 (N_35179,N_34735,N_34957);
nor U35180 (N_35180,N_32129,N_34528);
or U35181 (N_35181,N_30520,N_30174);
xor U35182 (N_35182,N_34751,N_32457);
and U35183 (N_35183,N_31007,N_33627);
and U35184 (N_35184,N_34329,N_31054);
nor U35185 (N_35185,N_30021,N_33313);
nor U35186 (N_35186,N_31374,N_33195);
and U35187 (N_35187,N_33977,N_33784);
and U35188 (N_35188,N_30086,N_33987);
nor U35189 (N_35189,N_30118,N_31562);
and U35190 (N_35190,N_33471,N_31089);
or U35191 (N_35191,N_30083,N_30617);
nand U35192 (N_35192,N_30740,N_32462);
nor U35193 (N_35193,N_33100,N_32583);
nand U35194 (N_35194,N_34411,N_32337);
and U35195 (N_35195,N_32493,N_32147);
and U35196 (N_35196,N_30483,N_32591);
xor U35197 (N_35197,N_33168,N_32292);
or U35198 (N_35198,N_30542,N_33758);
nor U35199 (N_35199,N_30984,N_30594);
or U35200 (N_35200,N_33597,N_33292);
and U35201 (N_35201,N_33767,N_34713);
nand U35202 (N_35202,N_34884,N_34032);
nor U35203 (N_35203,N_30911,N_33232);
and U35204 (N_35204,N_33033,N_34734);
xnor U35205 (N_35205,N_31224,N_34850);
and U35206 (N_35206,N_31555,N_34135);
and U35207 (N_35207,N_34680,N_31413);
and U35208 (N_35208,N_34247,N_32049);
nand U35209 (N_35209,N_33156,N_31148);
nor U35210 (N_35210,N_34352,N_30737);
nand U35211 (N_35211,N_32082,N_31397);
and U35212 (N_35212,N_32594,N_33488);
or U35213 (N_35213,N_33789,N_30789);
nand U35214 (N_35214,N_32928,N_33753);
or U35215 (N_35215,N_34809,N_34397);
xor U35216 (N_35216,N_34083,N_32693);
or U35217 (N_35217,N_33367,N_32370);
nand U35218 (N_35218,N_34012,N_32375);
nor U35219 (N_35219,N_32919,N_33325);
and U35220 (N_35220,N_31734,N_33483);
and U35221 (N_35221,N_34805,N_30832);
nor U35222 (N_35222,N_33807,N_33429);
and U35223 (N_35223,N_33583,N_34441);
or U35224 (N_35224,N_33190,N_32083);
or U35225 (N_35225,N_32131,N_33053);
and U35226 (N_35226,N_33933,N_34087);
or U35227 (N_35227,N_34265,N_34685);
nand U35228 (N_35228,N_31174,N_34095);
nor U35229 (N_35229,N_34112,N_33494);
nor U35230 (N_35230,N_30723,N_30074);
nand U35231 (N_35231,N_33809,N_32342);
nor U35232 (N_35232,N_34872,N_30796);
nand U35233 (N_35233,N_34681,N_33193);
nand U35234 (N_35234,N_31708,N_32927);
nor U35235 (N_35235,N_31924,N_30371);
nor U35236 (N_35236,N_33480,N_33710);
xor U35237 (N_35237,N_31377,N_31111);
and U35238 (N_35238,N_33050,N_33078);
and U35239 (N_35239,N_33699,N_33578);
nand U35240 (N_35240,N_31305,N_34107);
nand U35241 (N_35241,N_33431,N_30269);
xor U35242 (N_35242,N_34616,N_30771);
or U35243 (N_35243,N_30951,N_33620);
nand U35244 (N_35244,N_30105,N_30294);
nor U35245 (N_35245,N_33177,N_34373);
and U35246 (N_35246,N_32243,N_33771);
nand U35247 (N_35247,N_33795,N_30820);
and U35248 (N_35248,N_30867,N_31854);
nor U35249 (N_35249,N_33061,N_33800);
or U35250 (N_35250,N_34858,N_31511);
nand U35251 (N_35251,N_30134,N_34562);
nor U35252 (N_35252,N_31679,N_32128);
or U35253 (N_35253,N_33071,N_34437);
and U35254 (N_35254,N_31651,N_32820);
nor U35255 (N_35255,N_31951,N_31709);
or U35256 (N_35256,N_31546,N_33057);
nand U35257 (N_35257,N_30880,N_31458);
nand U35258 (N_35258,N_33535,N_31749);
or U35259 (N_35259,N_33444,N_31468);
nand U35260 (N_35260,N_33553,N_33107);
nand U35261 (N_35261,N_32920,N_34970);
nand U35262 (N_35262,N_33386,N_30660);
or U35263 (N_35263,N_33425,N_31856);
xor U35264 (N_35264,N_31669,N_34055);
or U35265 (N_35265,N_31229,N_32500);
and U35266 (N_35266,N_30691,N_31587);
and U35267 (N_35267,N_30561,N_32514);
nor U35268 (N_35268,N_32902,N_34129);
nand U35269 (N_35269,N_30054,N_34491);
and U35270 (N_35270,N_34823,N_31469);
nand U35271 (N_35271,N_34904,N_34148);
nor U35272 (N_35272,N_33132,N_30513);
or U35273 (N_35273,N_33814,N_32962);
or U35274 (N_35274,N_33827,N_34631);
or U35275 (N_35275,N_31384,N_33046);
xor U35276 (N_35276,N_31719,N_32516);
nor U35277 (N_35277,N_30088,N_33592);
nor U35278 (N_35278,N_30967,N_32922);
xor U35279 (N_35279,N_30858,N_30005);
or U35280 (N_35280,N_31099,N_30067);
or U35281 (N_35281,N_34780,N_31817);
nand U35282 (N_35282,N_33625,N_31796);
and U35283 (N_35283,N_32589,N_34110);
or U35284 (N_35284,N_34926,N_30321);
nor U35285 (N_35285,N_31844,N_30865);
nand U35286 (N_35286,N_31447,N_30825);
nand U35287 (N_35287,N_33957,N_31446);
and U35288 (N_35288,N_30332,N_31862);
nor U35289 (N_35289,N_31715,N_33362);
and U35290 (N_35290,N_32228,N_31826);
xnor U35291 (N_35291,N_33970,N_33713);
and U35292 (N_35292,N_33250,N_30494);
nand U35293 (N_35293,N_31676,N_33322);
nor U35294 (N_35294,N_30273,N_33272);
or U35295 (N_35295,N_33159,N_33418);
nand U35296 (N_35296,N_31080,N_31785);
nor U35297 (N_35297,N_34461,N_33120);
xor U35298 (N_35298,N_31547,N_33762);
and U35299 (N_35299,N_33689,N_30512);
nor U35300 (N_35300,N_32051,N_33954);
nor U35301 (N_35301,N_32165,N_34640);
and U35302 (N_35302,N_34676,N_32313);
or U35303 (N_35303,N_31549,N_34429);
nor U35304 (N_35304,N_32486,N_30077);
or U35305 (N_35305,N_34743,N_32879);
and U35306 (N_35306,N_34865,N_30339);
or U35307 (N_35307,N_30471,N_31768);
or U35308 (N_35308,N_33128,N_33183);
and U35309 (N_35309,N_34667,N_30369);
nand U35310 (N_35310,N_30678,N_31942);
or U35311 (N_35311,N_34477,N_33575);
nor U35312 (N_35312,N_33170,N_33104);
nand U35313 (N_35313,N_30057,N_34372);
xnor U35314 (N_35314,N_32532,N_33278);
nand U35315 (N_35315,N_31985,N_32638);
and U35316 (N_35316,N_32213,N_32778);
and U35317 (N_35317,N_32505,N_31273);
and U35318 (N_35318,N_30501,N_32264);
nor U35319 (N_35319,N_30776,N_34092);
and U35320 (N_35320,N_30945,N_30315);
xor U35321 (N_35321,N_33423,N_34182);
or U35322 (N_35322,N_33020,N_33561);
nand U35323 (N_35323,N_30926,N_33581);
nand U35324 (N_35324,N_34144,N_32001);
or U35325 (N_35325,N_33959,N_33477);
or U35326 (N_35326,N_34249,N_31035);
and U35327 (N_35327,N_32052,N_30028);
xnor U35328 (N_35328,N_32117,N_31289);
or U35329 (N_35329,N_31600,N_30846);
nor U35330 (N_35330,N_32599,N_30308);
nor U35331 (N_35331,N_34382,N_34953);
and U35332 (N_35332,N_34915,N_34530);
nand U35333 (N_35333,N_33978,N_31076);
or U35334 (N_35334,N_30034,N_33988);
xor U35335 (N_35335,N_30595,N_31153);
and U35336 (N_35336,N_34142,N_31175);
or U35337 (N_35337,N_30934,N_30261);
nand U35338 (N_35338,N_30326,N_32815);
nor U35339 (N_35339,N_33616,N_30546);
nand U35340 (N_35340,N_33878,N_30953);
and U35341 (N_35341,N_31901,N_32581);
nand U35342 (N_35342,N_32174,N_33158);
nor U35343 (N_35343,N_31353,N_33124);
nor U35344 (N_35344,N_31921,N_32695);
nand U35345 (N_35345,N_31395,N_34169);
and U35346 (N_35346,N_31839,N_32484);
and U35347 (N_35347,N_30290,N_31783);
and U35348 (N_35348,N_30305,N_33938);
nand U35349 (N_35349,N_32823,N_30965);
and U35350 (N_35350,N_33154,N_32015);
or U35351 (N_35351,N_33191,N_30217);
or U35352 (N_35352,N_32293,N_33644);
nand U35353 (N_35353,N_30227,N_31401);
and U35354 (N_35354,N_33385,N_33862);
xor U35355 (N_35355,N_31276,N_30310);
and U35356 (N_35356,N_30424,N_30758);
and U35357 (N_35357,N_33274,N_33788);
nor U35358 (N_35358,N_34325,N_34797);
xor U35359 (N_35359,N_30409,N_33989);
xnor U35360 (N_35360,N_32747,N_31611);
xnor U35361 (N_35361,N_32540,N_33172);
xnor U35362 (N_35362,N_33114,N_31178);
nand U35363 (N_35363,N_32776,N_31712);
xor U35364 (N_35364,N_33778,N_34029);
or U35365 (N_35365,N_34938,N_30550);
nor U35366 (N_35366,N_33083,N_33886);
and U35367 (N_35367,N_34100,N_34154);
and U35368 (N_35368,N_30533,N_30675);
nor U35369 (N_35369,N_32605,N_31723);
and U35370 (N_35370,N_32004,N_30121);
nand U35371 (N_35371,N_30502,N_31863);
nor U35372 (N_35372,N_30189,N_32894);
nand U35373 (N_35373,N_31701,N_30406);
nor U35374 (N_35374,N_32417,N_33473);
nor U35375 (N_35375,N_30673,N_31608);
nand U35376 (N_35376,N_31722,N_32744);
nor U35377 (N_35377,N_33324,N_31337);
and U35378 (N_35378,N_31379,N_34196);
xnor U35379 (N_35379,N_32096,N_33028);
and U35380 (N_35380,N_33615,N_34258);
nand U35381 (N_35381,N_30304,N_32760);
and U35382 (N_35382,N_32733,N_32050);
nor U35383 (N_35383,N_30497,N_34592);
nor U35384 (N_35384,N_34363,N_31559);
xnor U35385 (N_35385,N_34147,N_30923);
nand U35386 (N_35386,N_32832,N_30654);
nor U35387 (N_35387,N_33559,N_31805);
or U35388 (N_35388,N_32895,N_32203);
nor U35389 (N_35389,N_33646,N_30098);
nor U35390 (N_35390,N_33456,N_33703);
nor U35391 (N_35391,N_32265,N_33542);
xnor U35392 (N_35392,N_31228,N_32604);
nor U35393 (N_35393,N_32712,N_33927);
and U35394 (N_35394,N_33410,N_34008);
xor U35395 (N_35395,N_34431,N_30543);
xor U35396 (N_35396,N_33900,N_31540);
nor U35397 (N_35397,N_30681,N_34535);
and U35398 (N_35398,N_34454,N_32560);
nor U35399 (N_35399,N_34428,N_31639);
xnor U35400 (N_35400,N_34746,N_34465);
nor U35401 (N_35401,N_31577,N_30999);
nor U35402 (N_35402,N_34763,N_30102);
or U35403 (N_35403,N_30979,N_33035);
nand U35404 (N_35404,N_30962,N_30156);
and U35405 (N_35405,N_30765,N_30433);
and U35406 (N_35406,N_32474,N_31081);
and U35407 (N_35407,N_32404,N_34200);
and U35408 (N_35408,N_33963,N_34150);
or U35409 (N_35409,N_34764,N_31917);
xnor U35410 (N_35410,N_30044,N_32864);
nor U35411 (N_35411,N_34912,N_33441);
nand U35412 (N_35412,N_32819,N_30410);
or U35413 (N_35413,N_32893,N_32216);
and U35414 (N_35414,N_31331,N_32763);
and U35415 (N_35415,N_32997,N_31340);
and U35416 (N_35416,N_32268,N_30033);
and U35417 (N_35417,N_30170,N_32012);
or U35418 (N_35418,N_33405,N_32970);
nand U35419 (N_35419,N_32179,N_31448);
or U35420 (N_35420,N_30391,N_32750);
and U35421 (N_35421,N_30703,N_33348);
nand U35422 (N_35422,N_33793,N_34149);
or U35423 (N_35423,N_33691,N_34607);
or U35424 (N_35424,N_31943,N_31945);
nor U35425 (N_35425,N_31092,N_31295);
or U35426 (N_35426,N_33026,N_32353);
or U35427 (N_35427,N_30986,N_32305);
and U35428 (N_35428,N_34157,N_34599);
and U35429 (N_35429,N_33346,N_32769);
or U35430 (N_35430,N_30267,N_31852);
nand U35431 (N_35431,N_34484,N_30219);
xor U35432 (N_35432,N_31657,N_31895);
nand U35433 (N_35433,N_32347,N_33701);
nor U35434 (N_35434,N_32557,N_30239);
or U35435 (N_35435,N_31753,N_33504);
and U35436 (N_35436,N_31242,N_31342);
nor U35437 (N_35437,N_30976,N_34755);
nand U35438 (N_35438,N_31571,N_31492);
and U35439 (N_35439,N_34600,N_30635);
nand U35440 (N_35440,N_30632,N_32673);
xor U35441 (N_35441,N_31965,N_30073);
nand U35442 (N_35442,N_34037,N_34941);
and U35443 (N_35443,N_31997,N_30555);
xnor U35444 (N_35444,N_31686,N_32204);
nor U35445 (N_35445,N_31561,N_30469);
nand U35446 (N_35446,N_33184,N_33985);
or U35447 (N_35447,N_30944,N_30445);
or U35448 (N_35448,N_32945,N_34097);
and U35449 (N_35449,N_32000,N_34186);
nand U35450 (N_35450,N_30786,N_32106);
or U35451 (N_35451,N_32914,N_34578);
nor U35452 (N_35452,N_32528,N_33460);
xnor U35453 (N_35453,N_32848,N_32274);
nand U35454 (N_35454,N_31334,N_33163);
nand U35455 (N_35455,N_34344,N_32048);
nor U35456 (N_35456,N_30695,N_30787);
xnor U35457 (N_35457,N_33136,N_32218);
or U35458 (N_35458,N_33918,N_33852);
nand U35459 (N_35459,N_33975,N_31126);
or U35460 (N_35460,N_33540,N_31599);
nand U35461 (N_35461,N_30182,N_30299);
and U35462 (N_35462,N_31988,N_31866);
nand U35463 (N_35463,N_32429,N_30629);
xor U35464 (N_35464,N_32281,N_32758);
and U35465 (N_35465,N_33980,N_32383);
nor U35466 (N_35466,N_30918,N_33484);
nand U35467 (N_35467,N_31583,N_33133);
nand U35468 (N_35468,N_31678,N_30055);
or U35469 (N_35469,N_33668,N_32772);
and U35470 (N_35470,N_34309,N_34217);
nand U35471 (N_35471,N_32377,N_33534);
or U35472 (N_35472,N_32574,N_31010);
or U35473 (N_35473,N_32098,N_32637);
or U35474 (N_35474,N_32199,N_32721);
or U35475 (N_35475,N_32878,N_30836);
or U35476 (N_35476,N_34399,N_34702);
or U35477 (N_35477,N_30237,N_32481);
nand U35478 (N_35478,N_33589,N_30327);
and U35479 (N_35479,N_34610,N_34346);
or U35480 (N_35480,N_30337,N_34773);
or U35481 (N_35481,N_33462,N_34145);
nor U35482 (N_35482,N_31981,N_33155);
nor U35483 (N_35483,N_30685,N_32161);
nor U35484 (N_35484,N_32025,N_33024);
nand U35485 (N_35485,N_30152,N_34266);
or U35486 (N_35486,N_31751,N_33173);
or U35487 (N_35487,N_31246,N_31731);
nor U35488 (N_35488,N_30676,N_32887);
or U35489 (N_35489,N_30255,N_30784);
and U35490 (N_35490,N_30428,N_33215);
or U35491 (N_35491,N_32507,N_31672);
xor U35492 (N_35492,N_33859,N_30091);
nor U35493 (N_35493,N_31641,N_32231);
nand U35494 (N_35494,N_34230,N_34539);
and U35495 (N_35495,N_33436,N_33370);
nor U35496 (N_35496,N_32754,N_34655);
nor U35497 (N_35497,N_30829,N_32634);
and U35498 (N_35498,N_30220,N_30599);
or U35499 (N_35499,N_30722,N_34890);
or U35500 (N_35500,N_34077,N_33387);
xnor U35501 (N_35501,N_34629,N_33279);
or U35502 (N_35502,N_31026,N_33913);
nor U35503 (N_35503,N_34944,N_31758);
and U35504 (N_35504,N_31048,N_32080);
or U35505 (N_35505,N_33902,N_34490);
and U35506 (N_35506,N_30251,N_34398);
and U35507 (N_35507,N_30707,N_32421);
or U35508 (N_35508,N_30043,N_30680);
nand U35509 (N_35509,N_30993,N_31084);
nand U35510 (N_35510,N_34948,N_34318);
and U35511 (N_35511,N_31991,N_32618);
nand U35512 (N_35512,N_31954,N_31778);
xor U35513 (N_35513,N_33727,N_32258);
and U35514 (N_35514,N_34071,N_32075);
nand U35515 (N_35515,N_34166,N_31038);
xor U35516 (N_35516,N_30314,N_33979);
or U35517 (N_35517,N_33427,N_30794);
and U35518 (N_35518,N_34705,N_31834);
or U35519 (N_35519,N_31543,N_34199);
nand U35520 (N_35520,N_30169,N_32222);
nand U35521 (N_35521,N_34483,N_34102);
nand U35522 (N_35522,N_34534,N_31714);
or U35523 (N_35523,N_30526,N_33355);
nor U35524 (N_35524,N_30625,N_30168);
nand U35525 (N_35525,N_32367,N_34789);
or U35526 (N_35526,N_33521,N_32686);
and U35527 (N_35527,N_34877,N_34722);
nor U35528 (N_35528,N_31612,N_34140);
and U35529 (N_35529,N_30061,N_34660);
nand U35530 (N_35530,N_34170,N_31684);
nand U35531 (N_35531,N_32840,N_34011);
nor U35532 (N_35532,N_34332,N_30093);
nand U35533 (N_35533,N_34187,N_32978);
and U35534 (N_35534,N_33569,N_31145);
nand U35535 (N_35535,N_34207,N_30206);
nand U35536 (N_35536,N_30868,N_34976);
nand U35537 (N_35537,N_34605,N_30379);
nor U35538 (N_35538,N_31320,N_30975);
nor U35539 (N_35539,N_32639,N_33048);
and U35540 (N_35540,N_32985,N_32172);
nand U35541 (N_35541,N_31208,N_33130);
and U35542 (N_35542,N_32861,N_32061);
nand U35543 (N_35543,N_33186,N_33863);
and U35544 (N_35544,N_33768,N_33216);
and U35545 (N_35545,N_32194,N_33388);
nor U35546 (N_35546,N_32716,N_30592);
nor U35547 (N_35547,N_34570,N_32938);
xor U35548 (N_35548,N_33426,N_32250);
xnor U35549 (N_35549,N_31254,N_31323);
nand U35550 (N_35550,N_33667,N_34295);
or U35551 (N_35551,N_31648,N_32413);
nor U35552 (N_35552,N_30567,N_34300);
xor U35553 (N_35553,N_30839,N_31290);
or U35554 (N_35554,N_32115,N_34119);
or U35555 (N_35555,N_34375,N_30238);
or U35556 (N_35556,N_32382,N_31245);
or U35557 (N_35557,N_30385,N_34201);
xnor U35558 (N_35558,N_30810,N_32306);
nor U35559 (N_35559,N_33531,N_32257);
xnor U35560 (N_35560,N_31556,N_34028);
nand U35561 (N_35561,N_31151,N_31283);
and U35562 (N_35562,N_34098,N_33347);
and U35563 (N_35563,N_33630,N_32079);
nand U35564 (N_35564,N_30977,N_33919);
nor U35565 (N_35565,N_34898,N_31416);
or U35566 (N_35566,N_32324,N_30484);
and U35567 (N_35567,N_31630,N_32897);
and U35568 (N_35568,N_34267,N_30280);
or U35569 (N_35569,N_33718,N_32789);
nor U35570 (N_35570,N_32690,N_33469);
nand U35571 (N_35571,N_32536,N_32607);
and U35572 (N_35572,N_32579,N_30198);
or U35573 (N_35573,N_31322,N_31004);
nor U35574 (N_35574,N_31801,N_31662);
nand U35575 (N_35575,N_32309,N_30698);
nand U35576 (N_35576,N_32139,N_34175);
and U35577 (N_35577,N_31999,N_31756);
nand U35578 (N_35578,N_32005,N_34075);
or U35579 (N_35579,N_31001,N_33271);
and U35580 (N_35580,N_32333,N_31925);
or U35581 (N_35581,N_31920,N_31811);
and U35582 (N_35582,N_32973,N_34989);
or U35583 (N_35583,N_32326,N_30713);
or U35584 (N_35584,N_33684,N_33613);
or U35585 (N_35585,N_30899,N_32476);
nor U35586 (N_35586,N_34896,N_33448);
and U35587 (N_35587,N_34480,N_32390);
nand U35588 (N_35588,N_32714,N_31388);
or U35589 (N_35589,N_32006,N_32561);
nor U35590 (N_35590,N_31818,N_32214);
and U35591 (N_35591,N_33580,N_31514);
or U35592 (N_35592,N_32899,N_32658);
nor U35593 (N_35593,N_33675,N_32582);
nand U35594 (N_35594,N_31588,N_30666);
and U35595 (N_35595,N_34416,N_31936);
and U35596 (N_35596,N_30049,N_33047);
xnor U35597 (N_35597,N_30296,N_31944);
and U35598 (N_35598,N_34794,N_34004);
nand U35599 (N_35599,N_32135,N_34806);
nor U35600 (N_35600,N_32078,N_34404);
and U35601 (N_35601,N_30655,N_34046);
nor U35602 (N_35602,N_31505,N_30995);
nor U35603 (N_35603,N_31241,N_33996);
nand U35604 (N_35604,N_31275,N_33277);
nor U35605 (N_35605,N_32159,N_30500);
nand U35606 (N_35606,N_32676,N_33860);
nand U35607 (N_35607,N_33302,N_32398);
nor U35608 (N_35608,N_33826,N_34388);
and U35609 (N_35609,N_31259,N_34240);
or U35610 (N_35610,N_30382,N_34911);
or U35611 (N_35611,N_32534,N_33010);
nor U35612 (N_35612,N_33181,N_33502);
and U35613 (N_35613,N_33637,N_30529);
nor U35614 (N_35614,N_30176,N_31923);
xnor U35615 (N_35615,N_33492,N_34307);
and U35616 (N_35616,N_33929,N_30426);
nand U35617 (N_35617,N_30117,N_33161);
and U35618 (N_35618,N_31634,N_32378);
nand U35619 (N_35619,N_34923,N_34776);
nand U35620 (N_35620,N_32502,N_33185);
and U35621 (N_35621,N_34422,N_32363);
nor U35622 (N_35622,N_30416,N_33823);
or U35623 (N_35623,N_34979,N_30618);
xor U35624 (N_35624,N_33230,N_34879);
nand U35625 (N_35625,N_31442,N_30798);
or U35626 (N_35626,N_33672,N_32290);
and U35627 (N_35627,N_30879,N_33101);
xnor U35628 (N_35628,N_31963,N_31150);
and U35629 (N_35629,N_34627,N_33282);
or U35630 (N_35630,N_31106,N_30364);
nand U35631 (N_35631,N_34961,N_30811);
and U35632 (N_35632,N_34426,N_32031);
nor U35633 (N_35633,N_34276,N_34753);
nor U35634 (N_35634,N_30147,N_32859);
nand U35635 (N_35635,N_33375,N_31530);
or U35636 (N_35636,N_34254,N_30048);
and U35637 (N_35637,N_30733,N_32804);
nor U35638 (N_35638,N_32836,N_34213);
xnor U35639 (N_35639,N_33449,N_32196);
and U35640 (N_35640,N_34821,N_31223);
nor U35641 (N_35641,N_33853,N_30201);
nand U35642 (N_35642,N_30075,N_32913);
xnor U35643 (N_35643,N_33907,N_31346);
xor U35644 (N_35644,N_31198,N_34589);
and U35645 (N_35645,N_31324,N_31476);
nand U35646 (N_35646,N_34457,N_31421);
nor U35647 (N_35647,N_30311,N_33123);
and U35648 (N_35648,N_32724,N_34243);
nor U35649 (N_35649,N_31425,N_33941);
or U35650 (N_35650,N_32803,N_33510);
or U35651 (N_35651,N_33121,N_33457);
nor U35652 (N_35652,N_33223,N_30700);
or U35653 (N_35653,N_31268,N_33350);
or U35654 (N_35654,N_33001,N_30835);
nor U35655 (N_35655,N_33847,N_30537);
and U35656 (N_35656,N_33143,N_31539);
nand U35657 (N_35657,N_34151,N_33349);
or U35658 (N_35658,N_31841,N_33304);
or U35659 (N_35659,N_30051,N_30601);
xnor U35660 (N_35660,N_34192,N_31296);
and U35661 (N_35661,N_32158,N_32972);
or U35662 (N_35662,N_32299,N_30166);
nor U35663 (N_35663,N_32566,N_34965);
nor U35664 (N_35664,N_33715,N_34918);
and U35665 (N_35665,N_34687,N_30395);
and U35666 (N_35666,N_31585,N_33949);
nor U35667 (N_35667,N_30874,N_31047);
and U35668 (N_35668,N_34716,N_31451);
or U35669 (N_35669,N_32045,N_30341);
and U35670 (N_35670,N_33931,N_31217);
and U35671 (N_35671,N_33403,N_33135);
and U35672 (N_35672,N_32119,N_30000);
nor U35673 (N_35673,N_30383,N_34273);
and U35674 (N_35674,N_34533,N_30652);
and U35675 (N_35675,N_33635,N_33934);
and U35676 (N_35676,N_30449,N_34856);
or U35677 (N_35677,N_32100,N_32133);
nor U35678 (N_35678,N_34189,N_31138);
nand U35679 (N_35679,N_32954,N_31443);
xor U35680 (N_35680,N_30656,N_31987);
nand U35681 (N_35681,N_31409,N_30080);
or U35682 (N_35682,N_32287,N_32380);
nor U35683 (N_35683,N_31282,N_33628);
nand U35684 (N_35684,N_34524,N_32057);
and U35685 (N_35685,N_34418,N_34917);
and U35686 (N_35686,N_30506,N_31059);
and U35687 (N_35687,N_32826,N_32340);
nand U35688 (N_35688,N_32373,N_31726);
or U35689 (N_35689,N_30828,N_34093);
nor U35690 (N_35690,N_33472,N_32198);
or U35691 (N_35691,N_30919,N_34798);
nor U35692 (N_35692,N_34215,N_34390);
nand U35693 (N_35693,N_30203,N_32066);
nor U35694 (N_35694,N_31251,N_32010);
xnor U35695 (N_35695,N_34237,N_32488);
or U35696 (N_35696,N_31759,N_33554);
nor U35697 (N_35697,N_30716,N_32530);
and U35698 (N_35698,N_34474,N_31972);
nor U35699 (N_35699,N_33486,N_32650);
xor U35700 (N_35700,N_32707,N_32357);
or U35701 (N_35701,N_31415,N_34277);
nor U35702 (N_35702,N_32512,N_32720);
xor U35703 (N_35703,N_32443,N_30495);
nand U35704 (N_35704,N_34648,N_33811);
nand U35705 (N_35705,N_34553,N_32408);
or U35706 (N_35706,N_30841,N_32794);
or U35707 (N_35707,N_32272,N_33004);
and U35708 (N_35708,N_30076,N_34956);
xor U35709 (N_35709,N_30295,N_33574);
nor U35710 (N_35710,N_32246,N_31455);
xnor U35711 (N_35711,N_30204,N_31000);
nor U35712 (N_35712,N_30590,N_32524);
nor U35713 (N_35713,N_34044,N_32492);
nand U35714 (N_35714,N_34314,N_34928);
and U35715 (N_35715,N_31121,N_31391);
or U35716 (N_35716,N_32445,N_34481);
nor U35717 (N_35717,N_30181,N_34502);
nor U35718 (N_35718,N_32085,N_33947);
and U35719 (N_35719,N_30002,N_34766);
xnor U35720 (N_35720,N_30482,N_31112);
or U35721 (N_35721,N_33956,N_34579);
or U35722 (N_35722,N_30946,N_32529);
and U35723 (N_35723,N_33969,N_31063);
or U35724 (N_35724,N_34104,N_34639);
nand U35725 (N_35725,N_32713,N_30591);
or U35726 (N_35726,N_32882,N_34978);
and U35727 (N_35727,N_33731,N_30262);
nand U35728 (N_35728,N_34518,N_31597);
nor U35729 (N_35729,N_30082,N_30476);
nand U35730 (N_35730,N_32480,N_32449);
or U35731 (N_35731,N_33573,N_31799);
nand U35732 (N_35732,N_30626,N_30804);
nand U35733 (N_35733,N_33738,N_34710);
or U35734 (N_35734,N_32042,N_31615);
and U35735 (N_35735,N_32543,N_31781);
or U35736 (N_35736,N_30725,N_34466);
nor U35737 (N_35737,N_33805,N_31728);
and U35738 (N_35738,N_33160,N_33002);
nand U35739 (N_35739,N_30818,N_30336);
nor U35740 (N_35740,N_30040,N_33029);
and U35741 (N_35741,N_34069,N_32120);
nand U35742 (N_35742,N_32847,N_30213);
xor U35743 (N_35743,N_34488,N_33376);
or U35744 (N_35744,N_30809,N_32898);
and U35745 (N_35745,N_31417,N_33310);
xor U35746 (N_35746,N_31969,N_34876);
nand U35747 (N_35747,N_31727,N_34242);
nor U35748 (N_35748,N_31302,N_30573);
nor U35749 (N_35749,N_33881,N_31563);
nand U35750 (N_35750,N_31670,N_31513);
nand U35751 (N_35751,N_34369,N_33782);
nand U35752 (N_35752,N_31533,N_31332);
or U35753 (N_35753,N_33824,N_31333);
nand U35754 (N_35754,N_32186,N_31351);
nor U35755 (N_35755,N_30245,N_32935);
nand U35756 (N_35756,N_32791,N_30813);
xor U35757 (N_35757,N_34176,N_30563);
nand U35758 (N_35758,N_34358,N_30150);
nor U35759 (N_35759,N_33618,N_32344);
xnor U35760 (N_35760,N_30889,N_32584);
nand U35761 (N_35761,N_31506,N_31812);
or U35762 (N_35762,N_30157,N_33253);
nor U35763 (N_35763,N_30065,N_33787);
nor U35764 (N_35764,N_33649,N_30047);
or U35765 (N_35765,N_32929,N_34825);
xor U35766 (N_35766,N_34198,N_32414);
nand U35767 (N_35767,N_31117,N_34962);
and U35768 (N_35768,N_34538,N_34086);
xor U35769 (N_35769,N_33125,N_30046);
and U35770 (N_35770,N_31946,N_34294);
nor U35771 (N_35771,N_32101,N_33153);
or U35772 (N_35772,N_33673,N_34219);
nand U35773 (N_35773,N_32230,N_33221);
and U35774 (N_35774,N_31986,N_30404);
nor U35775 (N_35775,N_34228,N_33082);
and U35776 (N_35776,N_30154,N_33924);
nand U35777 (N_35777,N_31284,N_33867);
nand U35778 (N_35778,N_32511,N_31705);
xnor U35779 (N_35779,N_31810,N_33700);
xor U35780 (N_35780,N_32571,N_30087);
nor U35781 (N_35781,N_31167,N_30001);
nor U35782 (N_35782,N_30196,N_32924);
and U35783 (N_35783,N_32302,N_30572);
or U35784 (N_35784,N_31091,N_33696);
and U35785 (N_35785,N_34573,N_33952);
xor U35786 (N_35786,N_34930,N_32766);
nor U35787 (N_35787,N_30399,N_33769);
xnor U35788 (N_35788,N_30066,N_30588);
nor U35789 (N_35789,N_31603,N_34698);
and U35790 (N_35790,N_32756,N_33960);
and U35791 (N_35791,N_33897,N_31473);
and U35792 (N_35792,N_32588,N_31168);
xor U35793 (N_35793,N_31363,N_34966);
or U35794 (N_35794,N_31884,N_30457);
nor U35795 (N_35795,N_32046,N_32506);
and U35796 (N_35796,N_32388,N_32867);
nand U35797 (N_35797,N_34801,N_33645);
nand U35798 (N_35798,N_31083,N_33334);
nand U35799 (N_35799,N_32842,N_30842);
nand U35800 (N_35800,N_34737,N_32099);
or U35801 (N_35801,N_33679,N_31002);
and U35802 (N_35802,N_34413,N_33377);
xor U35803 (N_35803,N_33797,N_31434);
or U35804 (N_35804,N_33661,N_32361);
nand U35805 (N_35805,N_30440,N_32993);
and U35806 (N_35806,N_31532,N_31347);
and U35807 (N_35807,N_31584,N_31976);
nor U35808 (N_35808,N_32728,N_33608);
nor U35809 (N_35809,N_32286,N_32635);
nor U35810 (N_35810,N_30961,N_33506);
or U35811 (N_35811,N_33930,N_33901);
nor U35812 (N_35812,N_31097,N_32070);
or U35813 (N_35813,N_33775,N_31187);
xor U35814 (N_35814,N_31675,N_31062);
nand U35815 (N_35815,N_31733,N_30013);
and U35816 (N_35816,N_33869,N_30095);
nand U35817 (N_35817,N_31420,N_34871);
nand U35818 (N_35818,N_34133,N_34726);
xnor U35819 (N_35819,N_31085,N_31429);
nand U35820 (N_35820,N_34163,N_30822);
nand U35821 (N_35821,N_30981,N_31843);
and U35822 (N_35822,N_30142,N_34232);
or U35823 (N_35823,N_32981,N_32890);
or U35824 (N_35824,N_32624,N_33330);
nand U35825 (N_35825,N_31319,N_30963);
or U35826 (N_35826,N_31861,N_33481);
or U35827 (N_35827,N_32091,N_32947);
nand U35828 (N_35828,N_33345,N_33257);
or U35829 (N_35829,N_31393,N_31056);
and U35830 (N_35830,N_34367,N_30857);
nand U35831 (N_35831,N_32670,N_33328);
or U35832 (N_35832,N_34124,N_31335);
nor U35833 (N_35833,N_32546,N_31713);
and U35834 (N_35834,N_33849,N_30232);
nor U35835 (N_35835,N_33522,N_31596);
and U35836 (N_35836,N_30580,N_32273);
or U35837 (N_35837,N_32104,N_30659);
nor U35838 (N_35838,N_33605,N_33855);
or U35839 (N_35839,N_32873,N_34692);
or U35840 (N_35840,N_32395,N_32704);
or U35841 (N_35841,N_32021,N_32982);
or U35842 (N_35842,N_30848,N_33776);
or U35843 (N_35843,N_34482,N_34778);
and U35844 (N_35844,N_34334,N_33236);
nand U35845 (N_35845,N_32308,N_34653);
nor U35846 (N_35846,N_31978,N_31716);
nor U35847 (N_35847,N_33915,N_32701);
nand U35848 (N_35848,N_32232,N_33207);
nand U35849 (N_35849,N_30378,N_34696);
and U35850 (N_35850,N_31291,N_31435);
or U35851 (N_35851,N_34889,N_31426);
and U35852 (N_35852,N_33653,N_34410);
nor U35853 (N_35853,N_31979,N_34456);
nand U35854 (N_35854,N_30780,N_34990);
nand U35855 (N_35855,N_34887,N_32314);
nor U35856 (N_35856,N_34996,N_34749);
nand U35857 (N_35857,N_31735,N_32459);
or U35858 (N_35858,N_30570,N_34328);
nor U35859 (N_35859,N_33498,N_33998);
and U35860 (N_35860,N_33674,N_34184);
nor U35861 (N_35861,N_30008,N_34894);
nand U35862 (N_35862,N_30042,N_30877);
or U35863 (N_35863,N_30746,N_33688);
and U35864 (N_35864,N_30190,N_30089);
or U35865 (N_35865,N_33116,N_34204);
or U35866 (N_35866,N_31292,N_31207);
xor U35867 (N_35867,N_30348,N_30260);
or U35868 (N_35868,N_32657,N_33501);
or U35869 (N_35869,N_30587,N_30465);
and U35870 (N_35870,N_34747,N_30960);
nand U35871 (N_35871,N_30833,N_34052);
xnor U35872 (N_35872,N_32577,N_33636);
and U35873 (N_35873,N_34141,N_33935);
and U35874 (N_35874,N_34227,N_30525);
nor U35875 (N_35875,N_31721,N_31238);
nor U35876 (N_35876,N_34910,N_32812);
nor U35877 (N_35877,N_32912,N_32432);
or U35878 (N_35878,N_32545,N_34361);
and U35879 (N_35879,N_32009,N_32424);
nand U35880 (N_35880,N_30209,N_33817);
nand U35881 (N_35881,N_33720,N_31263);
or U35882 (N_35882,N_30356,N_34634);
and U35883 (N_35883,N_32102,N_34622);
nand U35884 (N_35884,N_34427,N_30275);
nand U35885 (N_35885,N_31858,N_32664);
or U35886 (N_35886,N_33249,N_30241);
or U35887 (N_35887,N_31432,N_31300);
and U35888 (N_35888,N_32643,N_31822);
nor U35889 (N_35889,N_31499,N_33669);
and U35890 (N_35890,N_34800,N_31192);
or U35891 (N_35891,N_34003,N_32188);
nand U35892 (N_35892,N_30907,N_31560);
nor U35893 (N_35893,N_32889,N_32784);
nand U35894 (N_35894,N_32183,N_33203);
nand U35895 (N_35895,N_31096,N_32442);
or U35896 (N_35896,N_31200,N_33265);
xor U35897 (N_35897,N_31485,N_30559);
nor U35898 (N_35898,N_30108,N_33866);
nor U35899 (N_35899,N_34638,N_31654);
nand U35900 (N_35900,N_34109,N_34775);
and U35901 (N_35901,N_34495,N_34721);
nand U35902 (N_35902,N_33092,N_33085);
and U35903 (N_35903,N_30444,N_31307);
nor U35904 (N_35904,N_33724,N_30883);
nand U35905 (N_35905,N_32114,N_34072);
or U35906 (N_35906,N_31814,N_30163);
and U35907 (N_35907,N_33730,N_30146);
or U35908 (N_35908,N_30235,N_31591);
and U35909 (N_35909,N_32813,N_32478);
nor U35910 (N_35910,N_34462,N_30264);
xor U35911 (N_35911,N_32678,N_30556);
or U35912 (N_35912,N_30443,N_31687);
nor U35913 (N_35913,N_31906,N_33352);
and U35914 (N_35914,N_31127,N_30701);
xor U35915 (N_35915,N_34336,N_30528);
nand U35916 (N_35916,N_31339,N_33226);
and U35917 (N_35917,N_32869,N_31855);
xnor U35918 (N_35918,N_30761,N_30493);
and U35919 (N_35919,N_31015,N_34603);
or U35920 (N_35920,N_33711,N_32238);
nand U35921 (N_35921,N_34139,N_32397);
nand U35922 (N_35922,N_30427,N_33412);
and U35923 (N_35923,N_30566,N_30205);
nor U35924 (N_35924,N_31520,N_31602);
nor U35925 (N_35925,N_34253,N_31958);
nand U35926 (N_35926,N_30366,N_32278);
nand U35927 (N_35927,N_30347,N_30606);
and U35928 (N_35928,N_32339,N_30875);
and U35929 (N_35929,N_34414,N_34914);
or U35930 (N_35930,N_30411,N_31232);
nor U35931 (N_35931,N_32345,N_31601);
and U35932 (N_35932,N_32156,N_34035);
nand U35933 (N_35933,N_32014,N_34155);
nor U35934 (N_35934,N_32221,N_33885);
and U35935 (N_35935,N_31311,N_33794);
and U35936 (N_35936,N_33951,N_33917);
or U35937 (N_35937,N_30068,N_33475);
or U35938 (N_35938,N_33298,N_33099);
or U35939 (N_35939,N_30721,N_30608);
nor U35940 (N_35940,N_31964,N_30524);
xor U35941 (N_35941,N_34712,N_32544);
or U35942 (N_35942,N_34897,N_30913);
and U35943 (N_35943,N_34331,N_33086);
xor U35944 (N_35944,N_34673,N_32438);
nand U35945 (N_35945,N_31149,N_30607);
nor U35946 (N_35946,N_30895,N_31044);
or U35947 (N_35947,N_33220,N_30989);
or U35948 (N_35948,N_30195,N_33011);
and U35949 (N_35949,N_33102,N_33235);
and U35950 (N_35950,N_30853,N_34281);
xnor U35951 (N_35951,N_34268,N_32746);
and U35952 (N_35952,N_30748,N_32779);
nand U35953 (N_35953,N_30300,N_33665);
nand U35954 (N_35954,N_34783,N_33461);
xnor U35955 (N_35955,N_34636,N_34051);
and U35956 (N_35956,N_32437,N_30488);
xnor U35957 (N_35957,N_32134,N_30467);
or U35958 (N_35958,N_32923,N_34257);
nor U35959 (N_35959,N_32030,N_34838);
or U35960 (N_35960,N_34043,N_32811);
nor U35961 (N_35961,N_33384,N_33180);
nor U35962 (N_35962,N_31813,N_32060);
or U35963 (N_35963,N_33094,N_34479);
nand U35964 (N_35964,N_34855,N_33742);
nor U35965 (N_35965,N_34506,N_30727);
or U35966 (N_35966,N_32266,N_34401);
or U35967 (N_35967,N_31402,N_34967);
nand U35968 (N_35968,N_30320,N_31221);
nor U35969 (N_35969,N_32725,N_34711);
nand U35970 (N_35970,N_30644,N_32426);
and U35971 (N_35971,N_31459,N_33825);
and U35972 (N_35972,N_32835,N_30653);
nand U35973 (N_35973,N_30736,N_32629);
and U35974 (N_35974,N_34137,N_33119);
xor U35975 (N_35975,N_30279,N_34476);
and U35976 (N_35976,N_34041,N_33074);
and U35977 (N_35977,N_30036,N_30459);
or U35978 (N_35978,N_30256,N_31947);
or U35979 (N_35979,N_30234,N_30004);
nand U35980 (N_35980,N_34255,N_34322);
nand U35981 (N_35981,N_30852,N_33365);
nor U35982 (N_35982,N_33297,N_34177);
nand U35983 (N_35983,N_34303,N_32229);
nor U35984 (N_35984,N_34984,N_30693);
or U35985 (N_35985,N_32215,N_33372);
or U35986 (N_35986,N_31016,N_31456);
nand U35987 (N_35987,N_32964,N_33218);
nor U35988 (N_35988,N_33311,N_31313);
and U35989 (N_35989,N_30200,N_34316);
and U35990 (N_35990,N_33443,N_31580);
nor U35991 (N_35991,N_32953,N_32059);
nor U35992 (N_35992,N_32855,N_30097);
nor U35993 (N_35993,N_31287,N_31776);
xnor U35994 (N_35994,N_33846,N_34299);
or U35995 (N_35995,N_32249,N_31141);
xnor U35996 (N_35996,N_34842,N_30453);
xnor U35997 (N_35997,N_30762,N_32814);
nor U35998 (N_35998,N_30432,N_30708);
nor U35999 (N_35999,N_34279,N_34019);
nand U36000 (N_36000,N_31623,N_30509);
and U36001 (N_36001,N_34278,N_30038);
nand U36002 (N_36002,N_33446,N_31024);
and U36003 (N_36003,N_30985,N_34732);
and U36004 (N_36004,N_33445,N_33198);
nand U36005 (N_36005,N_30511,N_31367);
nor U36006 (N_36006,N_33409,N_31934);
nor U36007 (N_36007,N_31120,N_31541);
nand U36008 (N_36008,N_31271,N_34731);
or U36009 (N_36009,N_34136,N_34444);
xnor U36010 (N_36010,N_32212,N_30987);
and U36011 (N_36011,N_30589,N_31461);
or U36012 (N_36012,N_34290,N_33468);
or U36013 (N_36013,N_32058,N_34792);
nor U36014 (N_36014,N_31439,N_33067);
or U36015 (N_36015,N_31748,N_30805);
nand U36016 (N_36016,N_31960,N_33211);
or U36017 (N_36017,N_31706,N_33084);
or U36018 (N_36018,N_32262,N_33594);
and U36019 (N_36019,N_30620,N_32415);
nand U36020 (N_36020,N_32225,N_30990);
nand U36021 (N_36021,N_33268,N_31338);
and U36022 (N_36022,N_32901,N_33875);
nand U36023 (N_36023,N_34741,N_33314);
nand U36024 (N_36024,N_31137,N_32145);
xor U36025 (N_36025,N_34505,N_31794);
nand U36026 (N_36026,N_34125,N_32513);
and U36027 (N_36027,N_33593,N_32606);
and U36028 (N_36028,N_30819,N_31236);
nand U36029 (N_36029,N_32828,N_32743);
and U36030 (N_36030,N_30158,N_34542);
nand U36031 (N_36031,N_32572,N_34866);
nand U36032 (N_36032,N_32227,N_34359);
and U36033 (N_36033,N_31642,N_31030);
or U36034 (N_36034,N_33926,N_33884);
or U36035 (N_36035,N_32960,N_31625);
and U36036 (N_36036,N_32063,N_31215);
nand U36037 (N_36037,N_30094,N_32880);
nor U36038 (N_36038,N_32948,N_31005);
and U36039 (N_36039,N_31400,N_34298);
nand U36040 (N_36040,N_32338,N_33857);
or U36041 (N_36041,N_30307,N_33165);
or U36042 (N_36042,N_31139,N_33739);
or U36043 (N_36043,N_30663,N_34436);
nand U36044 (N_36044,N_31114,N_34819);
or U36045 (N_36045,N_33281,N_31325);
and U36046 (N_36046,N_33525,N_32217);
nand U36047 (N_36047,N_31797,N_33530);
nor U36048 (N_36048,N_32647,N_30376);
nand U36049 (N_36049,N_30582,N_30192);
nor U36050 (N_36050,N_31406,N_30641);
xnor U36051 (N_36051,N_30114,N_34804);
or U36052 (N_36052,N_30630,N_33802);
nand U36053 (N_36053,N_34916,N_31807);
or U36054 (N_36054,N_33822,N_30527);
nand U36055 (N_36055,N_34132,N_33570);
or U36056 (N_36056,N_31517,N_30534);
xor U36057 (N_36057,N_32729,N_32780);
or U36058 (N_36058,N_30988,N_34127);
nor U36059 (N_36059,N_33032,N_30541);
and U36060 (N_36060,N_31072,N_31725);
and U36061 (N_36061,N_31650,N_31695);
or U36062 (N_36062,N_30470,N_33704);
or U36063 (N_36063,N_32471,N_33751);
or U36064 (N_36064,N_33654,N_31481);
nor U36065 (N_36065,N_30429,N_30516);
and U36066 (N_36066,N_32575,N_34864);
nand U36067 (N_36067,N_33707,N_31191);
xnor U36068 (N_36068,N_32295,N_34590);
or U36069 (N_36069,N_31199,N_32251);
or U36070 (N_36070,N_31019,N_34908);
or U36071 (N_36071,N_34214,N_30688);
nand U36072 (N_36072,N_34475,N_32441);
or U36073 (N_36073,N_31278,N_33493);
and U36074 (N_36074,N_32552,N_32235);
xor U36075 (N_36075,N_31693,N_31490);
nor U36076 (N_36076,N_30863,N_31404);
nand U36077 (N_36077,N_31996,N_34703);
or U36078 (N_36078,N_34206,N_31341);
and U36079 (N_36079,N_31524,N_32715);
or U36080 (N_36080,N_31902,N_32327);
and U36081 (N_36081,N_31519,N_33629);
nand U36082 (N_36082,N_33440,N_32193);
or U36083 (N_36083,N_31515,N_34614);
or U36084 (N_36084,N_31659,N_30735);
or U36085 (N_36085,N_33319,N_34647);
and U36086 (N_36086,N_31257,N_30715);
and U36087 (N_36087,N_33883,N_32271);
nand U36088 (N_36088,N_33489,N_34048);
nand U36089 (N_36089,N_32454,N_33819);
and U36090 (N_36090,N_32461,N_31431);
nand U36091 (N_36091,N_34348,N_32795);
or U36092 (N_36092,N_32959,N_32681);
and U36093 (N_36093,N_31008,N_34943);
or U36094 (N_36094,N_31230,N_32745);
or U36095 (N_36095,N_33321,N_34936);
nand U36096 (N_36096,N_33463,N_34026);
or U36097 (N_36097,N_33798,N_34515);
and U36098 (N_36098,N_31957,N_30463);
or U36099 (N_36099,N_32170,N_31326);
nand U36100 (N_36100,N_32567,N_32689);
xor U36101 (N_36101,N_30597,N_33666);
or U36102 (N_36102,N_34859,N_30751);
or U36103 (N_36103,N_30672,N_30532);
nor U36104 (N_36104,N_31256,N_32603);
nor U36105 (N_36105,N_31682,N_34645);
xor U36106 (N_36106,N_30631,N_34852);
and U36107 (N_36107,N_33896,N_31911);
and U36108 (N_36108,N_30922,N_32430);
nand U36109 (N_36109,N_33096,N_34421);
nand U36110 (N_36110,N_33299,N_30861);
nand U36111 (N_36111,N_33396,N_32142);
nor U36112 (N_36112,N_33708,N_32318);
nand U36113 (N_36113,N_33614,N_34354);
or U36114 (N_36114,N_33017,N_32040);
or U36115 (N_36115,N_32541,N_30071);
and U36116 (N_36116,N_32260,N_34870);
nand U36117 (N_36117,N_34091,N_32854);
nor U36118 (N_36118,N_31838,N_33944);
nand U36119 (N_36119,N_31569,N_34909);
nand U36120 (N_36120,N_30343,N_34387);
nand U36121 (N_36121,N_33434,N_32209);
nor U36122 (N_36122,N_31486,N_31607);
xnor U36123 (N_36123,N_30045,N_31500);
and U36124 (N_36124,N_31012,N_32300);
or U36125 (N_36125,N_33638,N_30180);
and U36126 (N_36126,N_34443,N_30360);
and U36127 (N_36127,N_34623,N_30997);
nor U36128 (N_36128,N_32435,N_33950);
and U36129 (N_36129,N_31130,N_31009);
or U36130 (N_36130,N_32409,N_33509);
nor U36131 (N_36131,N_30041,N_34955);
nand U36132 (N_36132,N_34557,N_33065);
nor U36133 (N_36133,N_32885,N_30257);
or U36134 (N_36134,N_31219,N_33722);
and U36135 (N_36135,N_34343,N_30301);
nor U36136 (N_36136,N_31927,N_32026);
or U36137 (N_36137,N_34719,N_32735);
nand U36138 (N_36138,N_32926,N_34706);
nand U36139 (N_36139,N_33063,N_34867);
nor U36140 (N_36140,N_31427,N_32989);
nor U36141 (N_36141,N_30277,N_32024);
xnor U36142 (N_36142,N_31739,N_31916);
nor U36143 (N_36143,N_33204,N_32137);
nand U36144 (N_36144,N_33414,N_32191);
nand U36145 (N_36145,N_30562,N_34762);
nand U36146 (N_36146,N_31793,N_33566);
nand U36147 (N_36147,N_31344,N_34489);
nor U36148 (N_36148,N_33558,N_34088);
and U36149 (N_36149,N_31154,N_34381);
xor U36150 (N_36150,N_30151,N_31011);
and U36151 (N_36151,N_31995,N_30623);
nand U36152 (N_36152,N_31131,N_31390);
nor U36153 (N_36153,N_31663,N_31700);
nor U36154 (N_36154,N_30092,N_31881);
nand U36155 (N_36155,N_30155,N_32269);
nand U36156 (N_36156,N_34569,N_30514);
nor U36157 (N_36157,N_32379,N_30900);
nand U36158 (N_36158,N_34674,N_34848);
nor U36159 (N_36159,N_31885,N_31140);
nor U36160 (N_36160,N_33073,N_30939);
or U36161 (N_36161,N_34153,N_31158);
or U36162 (N_36162,N_32242,N_33626);
or U36163 (N_36163,N_30197,N_31303);
nand U36164 (N_36164,N_34582,N_33518);
nand U36165 (N_36165,N_30286,N_34231);
and U36166 (N_36166,N_31831,N_30891);
nor U36167 (N_36167,N_34854,N_32931);
nand U36168 (N_36168,N_34487,N_33920);
nand U36169 (N_36169,N_31738,N_32202);
nor U36170 (N_36170,N_34921,N_34364);
nor U36171 (N_36171,N_30084,N_33122);
and U36172 (N_36172,N_33533,N_31116);
nor U36173 (N_36173,N_34761,N_31210);
xor U36174 (N_36174,N_34883,N_31928);
nor U36175 (N_36175,N_32123,N_33837);
or U36176 (N_36176,N_32751,N_31018);
xnor U36177 (N_36177,N_34492,N_33761);
and U36178 (N_36178,N_30162,N_33786);
xor U36179 (N_36179,N_30175,N_33152);
or U36180 (N_36180,N_31040,N_33754);
xnor U36181 (N_36181,N_34286,N_30396);
nor U36182 (N_36182,N_31689,N_32891);
or U36183 (N_36183,N_32944,N_32420);
and U36184 (N_36184,N_34922,N_34874);
and U36185 (N_36185,N_30032,N_33598);
nand U36186 (N_36186,N_30937,N_30943);
nand U36187 (N_36187,N_32709,N_34612);
nor U36188 (N_36188,N_31626,N_30344);
or U36189 (N_36189,N_30090,N_32623);
nor U36190 (N_36190,N_31522,N_31049);
nand U36191 (N_36191,N_33487,N_33906);
nor U36192 (N_36192,N_34601,N_33726);
nand U36193 (N_36193,N_30637,N_31220);
nor U36194 (N_36194,N_31368,N_33705);
nand U36195 (N_36195,N_32371,N_32645);
nor U36196 (N_36196,N_32460,N_34555);
or U36197 (N_36197,N_32598,N_31697);
or U36198 (N_36198,N_32297,N_30439);
and U36199 (N_36199,N_32844,N_31661);
nand U36200 (N_36200,N_32554,N_34478);
nand U36201 (N_36201,N_33612,N_31874);
nand U36202 (N_36202,N_33966,N_31467);
nor U36203 (N_36203,N_34814,N_31536);
nor U36204 (N_36204,N_30139,N_34420);
xnor U36205 (N_36205,N_31566,N_34308);
nand U36206 (N_36206,N_32761,N_33921);
or U36207 (N_36207,N_34241,N_30128);
nor U36208 (N_36208,N_31195,N_34446);
nor U36209 (N_36209,N_30669,N_32526);
or U36210 (N_36210,N_30312,N_30649);
nand U36211 (N_36211,N_30571,N_33217);
or U36212 (N_36212,N_33922,N_30978);
nand U36213 (N_36213,N_32490,N_31164);
nand U36214 (N_36214,N_31196,N_32691);
nand U36215 (N_36215,N_30998,N_33206);
nand U36216 (N_36216,N_34301,N_31203);
nand U36217 (N_36217,N_31696,N_32644);
nand U36218 (N_36218,N_31180,N_31235);
and U36219 (N_36219,N_30611,N_31538);
and U36220 (N_36220,N_30610,N_34827);
or U36221 (N_36221,N_32654,N_31935);
nor U36222 (N_36222,N_33080,N_34076);
nor U36223 (N_36223,N_33318,N_33582);
nor U36224 (N_36224,N_34284,N_33360);
and U36225 (N_36225,N_30224,N_33106);
and U36226 (N_36226,N_33040,N_33850);
nor U36227 (N_36227,N_32334,N_34860);
nor U36228 (N_36228,N_33757,N_32356);
or U36229 (N_36229,N_31565,N_33490);
nand U36230 (N_36230,N_33910,N_30442);
and U36231 (N_36231,N_31620,N_34532);
and U36232 (N_36232,N_31845,N_33126);
nor U36233 (N_36233,N_30991,N_30101);
and U36234 (N_36234,N_32665,N_34263);
nand U36235 (N_36235,N_32877,N_31304);
and U36236 (N_36236,N_30710,N_33777);
or U36237 (N_36237,N_31850,N_32301);
xnor U36238 (N_36238,N_30359,N_30064);
and U36239 (N_36239,N_34869,N_33087);
nand U36240 (N_36240,N_31029,N_34920);
nor U36241 (N_36241,N_32659,N_30350);
or U36242 (N_36242,N_32570,N_30750);
and U36243 (N_36243,N_33562,N_30731);
or U36244 (N_36244,N_32679,N_33420);
nand U36245 (N_36245,N_34531,N_32830);
and U36246 (N_36246,N_30354,N_31548);
nor U36247 (N_36247,N_32580,N_34053);
nand U36248 (N_36248,N_32071,N_31045);
or U36249 (N_36249,N_33072,N_30646);
or U36250 (N_36250,N_30925,N_34665);
and U36251 (N_36251,N_31385,N_33038);
and U36252 (N_36252,N_32496,N_33829);
nand U36253 (N_36253,N_31101,N_32614);
nor U36254 (N_36254,N_31170,N_30420);
and U36255 (N_36255,N_30430,N_31529);
nor U36256 (N_36256,N_33576,N_33514);
or U36257 (N_36257,N_34216,N_31747);
and U36258 (N_36258,N_31270,N_31266);
or U36259 (N_36259,N_30795,N_31003);
or U36260 (N_36260,N_34824,N_31163);
xnor U36261 (N_36261,N_32641,N_31741);
nand U36262 (N_36262,N_33693,N_33858);
and U36263 (N_36263,N_30113,N_30531);
or U36264 (N_36264,N_33465,N_31118);
or U36265 (N_36265,N_34010,N_33961);
and U36266 (N_36266,N_32585,N_34497);
nand U36267 (N_36267,N_30125,N_33134);
xnor U36268 (N_36268,N_32821,N_31102);
or U36269 (N_36269,N_34621,N_34464);
xor U36270 (N_36270,N_30029,N_32578);
and U36271 (N_36271,N_33030,N_33895);
xnor U36272 (N_36272,N_34355,N_34058);
nand U36273 (N_36273,N_34803,N_32037);
xor U36274 (N_36274,N_30670,N_34559);
or U36275 (N_36275,N_31980,N_34463);
or U36276 (N_36276,N_31912,N_31575);
nor U36277 (N_36277,N_34919,N_32391);
or U36278 (N_36278,N_34550,N_33194);
nand U36279 (N_36279,N_30317,N_31144);
nand U36280 (N_36280,N_30774,N_32239);
and U36281 (N_36281,N_33394,N_33406);
and U36282 (N_36282,N_32711,N_32111);
and U36283 (N_36283,N_34818,N_31886);
nand U36284 (N_36284,N_33587,N_32905);
xor U36285 (N_36285,N_34085,N_33234);
or U36286 (N_36286,N_34122,N_30742);
and U36287 (N_36287,N_34657,N_31694);
nor U36288 (N_36288,N_30887,N_33965);
nor U36289 (N_36289,N_34998,N_31698);
and U36290 (N_36290,N_30496,N_31389);
nor U36291 (N_36291,N_31082,N_34485);
nor U36292 (N_36292,N_32013,N_31824);
and U36293 (N_36293,N_31226,N_32710);
and U36294 (N_36294,N_32856,N_32402);
and U36295 (N_36295,N_32918,N_32946);
nand U36296 (N_36296,N_30648,N_34417);
nor U36297 (N_36297,N_30886,N_34062);
nor U36298 (N_36298,N_34964,N_30130);
or U36299 (N_36299,N_30603,N_30897);
nor U36300 (N_36300,N_30912,N_30037);
and U36301 (N_36301,N_33076,N_33595);
and U36302 (N_36302,N_32883,N_32807);
and U36303 (N_36303,N_31464,N_31330);
nand U36304 (N_36304,N_32033,N_34167);
nor U36305 (N_36305,N_31636,N_34256);
nand U36306 (N_36306,N_34682,N_34341);
or U36307 (N_36307,N_34469,N_30247);
nor U36308 (N_36308,N_33923,N_33288);
or U36309 (N_36309,N_33541,N_32374);
or U36310 (N_36310,N_32979,N_34335);
nor U36311 (N_36311,N_32044,N_32175);
and U36312 (N_36312,N_30208,N_34604);
nor U36313 (N_36313,N_32121,N_34195);
nor U36314 (N_36314,N_31252,N_33340);
nor U36315 (N_36315,N_30579,N_34954);
nor U36316 (N_36316,N_34400,N_34907);
nor U36317 (N_36317,N_33557,N_30807);
or U36318 (N_36318,N_34985,N_34750);
nor U36319 (N_36319,N_34571,N_30481);
xnor U36320 (N_36320,N_32613,N_31253);
or U36321 (N_36321,N_32587,N_31952);
or U36322 (N_36322,N_34886,N_34234);
xor U36323 (N_36323,N_31247,N_34459);
nor U36324 (N_36324,N_30642,N_30287);
nand U36325 (N_36325,N_31745,N_32089);
nand U36326 (N_36326,N_32936,N_32073);
or U36327 (N_36327,N_30521,N_32568);
nand U36328 (N_36328,N_32620,N_33329);
and U36329 (N_36329,N_33981,N_34440);
and U36330 (N_36330,N_31760,N_30187);
or U36331 (N_36331,N_34846,N_31243);
nand U36332 (N_36332,N_30942,N_34060);
nand U36333 (N_36333,N_31173,N_31777);
nor U36334 (N_36334,N_32531,N_30266);
nor U36335 (N_36335,N_30274,N_33657);
and U36336 (N_36336,N_34997,N_30830);
and U36337 (N_36337,N_31717,N_34433);
nor U36338 (N_36338,N_34808,N_33240);
nand U36339 (N_36339,N_30667,N_33157);
xnor U36340 (N_36340,N_34014,N_34280);
or U36341 (N_36341,N_34040,N_33633);
or U36342 (N_36342,N_34291,N_34831);
nor U36343 (N_36343,N_32275,N_32233);
nand U36344 (N_36344,N_30908,N_30393);
and U36345 (N_36345,N_31903,N_34940);
xor U36346 (N_36346,N_33984,N_34836);
nand U36347 (N_36347,N_30850,N_34593);
xor U36348 (N_36348,N_33815,N_32336);
and U36349 (N_36349,N_32685,N_31929);
nand U36350 (N_36350,N_33812,N_34030);
nand U36351 (N_36351,N_31244,N_33905);
xnor U36352 (N_36352,N_31649,N_34070);
nand U36353 (N_36353,N_32157,N_31462);
and U36354 (N_36354,N_30598,N_33021);
and U36355 (N_36355,N_34264,N_33247);
nand U36356 (N_36356,N_32934,N_30485);
and U36357 (N_36357,N_33442,N_33749);
nor U36358 (N_36358,N_30790,N_31457);
xnor U36359 (N_36359,N_34646,N_31086);
nor U36360 (N_36360,N_34839,N_32881);
nand U36361 (N_36361,N_32627,N_30766);
and U36362 (N_36362,N_30914,N_34642);
and U36363 (N_36363,N_33228,N_34021);
nor U36364 (N_36364,N_34089,N_31372);
nor U36365 (N_36365,N_33326,N_31680);
and U36366 (N_36366,N_33591,N_30063);
nand U36367 (N_36367,N_34270,N_34628);
nor U36368 (N_36368,N_34321,N_32667);
and U36369 (N_36369,N_33142,N_33188);
nand U36370 (N_36370,N_33993,N_33337);
nor U36371 (N_36371,N_32595,N_33607);
and U36372 (N_36372,N_31908,N_33098);
nand U36373 (N_36373,N_33609,N_30268);
nand U36374 (N_36374,N_34576,N_32316);
nor U36375 (N_36375,N_32358,N_31345);
or U36376 (N_36376,N_31234,N_32548);
xor U36377 (N_36377,N_31206,N_33799);
xnor U36378 (N_36378,N_34377,N_30797);
nor U36379 (N_36379,N_31037,N_30933);
nand U36380 (N_36380,N_33202,N_31982);
xnor U36381 (N_36381,N_32800,N_30183);
nand U36382 (N_36382,N_34275,N_34045);
and U36383 (N_36383,N_30243,N_32053);
or U36384 (N_36384,N_34999,N_30112);
and U36385 (N_36385,N_31299,N_30732);
and U36386 (N_36386,N_31820,N_32406);
nand U36387 (N_36387,N_32939,N_32032);
nor U36388 (N_36388,N_31454,N_32470);
and U36389 (N_36389,N_30932,N_31568);
nand U36390 (N_36390,N_31033,N_32590);
or U36391 (N_36391,N_33066,N_31977);
or U36392 (N_36392,N_30140,N_32783);
or U36393 (N_36393,N_34160,N_34022);
nand U36394 (N_36394,N_34777,N_32857);
nor U36395 (N_36395,N_30408,N_34688);
and U36396 (N_36396,N_32539,N_30111);
or U36397 (N_36397,N_34312,N_30866);
and U36398 (N_36398,N_32818,N_32097);
nand U36399 (N_36399,N_32576,N_33064);
nand U36400 (N_36400,N_31132,N_32752);
nor U36401 (N_36401,N_31440,N_33255);
xnor U36402 (N_36402,N_31297,N_32558);
nand U36403 (N_36403,N_32616,N_30634);
nor U36404 (N_36404,N_32307,N_31872);
nor U36405 (N_36405,N_32742,N_32064);
nand U36406 (N_36406,N_31632,N_30745);
and U36407 (N_36407,N_31239,N_32705);
or U36408 (N_36408,N_34672,N_33351);
and U36409 (N_36409,N_30236,N_33916);
nor U36410 (N_36410,N_30849,N_32888);
xor U36411 (N_36411,N_33430,N_32393);
nor U36412 (N_36412,N_31392,N_33940);
nor U36413 (N_36413,N_33601,N_30318);
xor U36414 (N_36414,N_30009,N_30584);
and U36415 (N_36415,N_34853,N_30365);
nand U36416 (N_36416,N_30136,N_31870);
nor U36417 (N_36417,N_32696,N_33640);
and U36418 (N_36418,N_31071,N_30226);
nand U36419 (N_36419,N_32076,N_30728);
and U36420 (N_36420,N_30966,N_33891);
xor U36421 (N_36421,N_33062,N_30699);
nand U36422 (N_36422,N_34156,N_32427);
nor U36423 (N_36423,N_31399,N_32034);
xor U36424 (N_36424,N_34840,N_31310);
nand U36425 (N_36425,N_33373,N_32792);
xnor U36426 (N_36426,N_32834,N_30662);
or U36427 (N_36427,N_32925,N_33031);
nand U36428 (N_36428,N_34849,N_30225);
nand U36429 (N_36429,N_34047,N_33624);
nor U36430 (N_36430,N_31983,N_33864);
nor U36431 (N_36431,N_32153,N_33936);
and U36432 (N_36432,N_31386,N_30160);
and U36433 (N_36433,N_32965,N_34670);
nor U36434 (N_36434,N_34644,N_30576);
xor U36435 (N_36435,N_32749,N_32494);
nand U36436 (N_36436,N_31637,N_31627);
and U36437 (N_36437,N_30284,N_34304);
or U36438 (N_36438,N_31990,N_33464);
and U36439 (N_36439,N_31444,N_31231);
and U36440 (N_36440,N_34288,N_32817);
or U36441 (N_36441,N_32240,N_32846);
or U36442 (N_36442,N_32833,N_32731);
nand U36443 (N_36443,N_30574,N_32255);
nor U36444 (N_36444,N_30329,N_32140);
nor U36445 (N_36445,N_34892,N_30803);
nand U36446 (N_36446,N_30661,N_33245);
nand U36447 (N_36447,N_32452,N_34123);
or U36448 (N_36448,N_31110,N_34516);
nor U36449 (N_36449,N_32138,N_34694);
or U36450 (N_36450,N_30342,N_31362);
nor U36451 (N_36451,N_31119,N_30876);
and U36452 (N_36452,N_30536,N_32473);
nor U36453 (N_36453,N_30971,N_34551);
nor U36454 (N_36454,N_33068,N_33435);
nand U36455 (N_36455,N_34718,N_33171);
xnor U36456 (N_36456,N_34929,N_31194);
nor U36457 (N_36457,N_34017,N_31550);
or U36458 (N_36458,N_30011,N_31528);
nor U36459 (N_36459,N_30696,N_31453);
nand U36460 (N_36460,N_32542,N_32331);
nand U36461 (N_36461,N_33090,N_30968);
nand U36462 (N_36462,N_31237,N_33818);
and U36463 (N_36463,N_32419,N_31261);
nand U36464 (N_36464,N_31825,N_33022);
nor U36465 (N_36465,N_30856,N_32399);
or U36466 (N_36466,N_33816,N_34527);
or U36467 (N_36467,N_34210,N_32827);
and U36468 (N_36468,N_33511,N_34507);
nor U36469 (N_36469,N_33650,N_31317);
nor U36470 (N_36470,N_30291,N_30193);
or U36471 (N_36471,N_34995,N_34202);
nor U36472 (N_36472,N_30164,N_34339);
or U36473 (N_36473,N_31614,N_34554);
nor U36474 (N_36474,N_30138,N_34649);
xor U36475 (N_36475,N_33932,N_32282);
nor U36476 (N_36476,N_30515,N_30473);
or U36477 (N_36477,N_32592,N_33470);
nor U36478 (N_36478,N_34927,N_32195);
and U36479 (N_36479,N_33454,N_34572);
or U36480 (N_36480,N_34271,N_30031);
or U36481 (N_36481,N_34130,N_34238);
nand U36482 (N_36482,N_34905,N_32625);
or U36483 (N_36483,N_34296,N_34547);
nand U36484 (N_36484,N_31621,N_33140);
nand U36485 (N_36485,N_33003,N_31182);
nor U36486 (N_36486,N_34991,N_32254);
nor U36487 (N_36487,N_30438,N_32977);
nand U36488 (N_36488,N_30952,N_34512);
xnor U36489 (N_36489,N_32043,N_34057);
or U36490 (N_36490,N_31655,N_33283);
nand U36491 (N_36491,N_30892,N_31185);
nand U36492 (N_36492,N_33467,N_34899);
nand U36493 (N_36493,N_30362,N_33604);
or U36494 (N_36494,N_33874,N_30581);
nor U36495 (N_36495,N_34738,N_31265);
and U36496 (N_36496,N_32086,N_33174);
and U36497 (N_36497,N_32372,N_30954);
or U36498 (N_36498,N_34969,N_32863);
xor U36499 (N_36499,N_34931,N_31498);
and U36500 (N_36500,N_34595,N_32477);
or U36501 (N_36501,N_32022,N_32423);
and U36502 (N_36502,N_32661,N_33251);
nor U36503 (N_36503,N_30885,N_34686);
nor U36504 (N_36504,N_32241,N_30401);
nand U36505 (N_36505,N_34983,N_30357);
or U36506 (N_36506,N_33060,N_32839);
nor U36507 (N_36507,N_33295,N_30149);
and U36508 (N_36508,N_31699,N_34895);
nor U36509 (N_36509,N_33527,N_34007);
and U36510 (N_36510,N_32267,N_33320);
nand U36511 (N_36511,N_34952,N_31477);
xor U36512 (N_36512,N_32669,N_30127);
nand U36513 (N_36513,N_34882,N_33547);
nand U36514 (N_36514,N_31366,N_31970);
nor U36515 (N_36515,N_32986,N_32458);
nand U36516 (N_36516,N_34677,N_33690);
and U36517 (N_36517,N_31835,N_31847);
nand U36518 (N_36518,N_33681,N_31020);
or U36519 (N_36519,N_30023,N_30565);
and U36520 (N_36520,N_33537,N_30331);
and U36521 (N_36521,N_31115,N_30959);
nor U36522 (N_36522,N_31665,N_33560);
and U36523 (N_36523,N_33109,N_34293);
nor U36524 (N_36524,N_34054,N_34320);
nor U36525 (N_36525,N_34924,N_34521);
or U36526 (N_36526,N_31865,N_31441);
nor U36527 (N_36527,N_31919,N_34379);
nand U36528 (N_36528,N_32976,N_30018);
nor U36529 (N_36529,N_34500,N_30413);
nor U36530 (N_36530,N_30479,N_34376);
nand U36531 (N_36531,N_31124,N_33743);
or U36532 (N_36532,N_32601,N_31779);
xor U36533 (N_36533,N_33368,N_34545);
nor U36534 (N_36534,N_33643,N_33671);
or U36535 (N_36535,N_32328,N_31430);
nand U36536 (N_36536,N_33942,N_34960);
or U36537 (N_36537,N_30815,N_30950);
nor U36538 (N_36538,N_30747,N_32446);
nor U36539 (N_36539,N_33772,N_30434);
nand U36540 (N_36540,N_31643,N_34078);
and U36541 (N_36541,N_33677,N_33105);
nor U36542 (N_36542,N_34049,N_31269);
xnor U36543 (N_36543,N_31105,N_34499);
nor U36544 (N_36544,N_32708,N_33831);
nor U36545 (N_36545,N_33025,N_33568);
nand U36546 (N_36546,N_34832,N_33982);
nand U36547 (N_36547,N_30425,N_30258);
nand U36548 (N_36548,N_31452,N_32942);
or U36549 (N_36549,N_33898,N_34193);
nor U36550 (N_36550,N_30462,N_34031);
xor U36551 (N_36551,N_31050,N_30674);
or U36552 (N_36552,N_31184,N_33258);
nand U36553 (N_36553,N_31354,N_31950);
and U36554 (N_36554,N_31285,N_31487);
nand U36555 (N_36555,N_30709,N_32211);
nand U36556 (N_36556,N_30910,N_30869);
and U36557 (N_36557,N_33479,N_33848);
nor U36558 (N_36558,N_31460,N_34034);
and U36559 (N_36559,N_34018,N_31966);
and U36560 (N_36560,N_31931,N_30099);
nor U36561 (N_36561,N_31074,N_34508);
nor U36562 (N_36562,N_33723,N_32801);
or U36563 (N_36563,N_30056,N_34633);
and U36564 (N_36564,N_30126,N_33438);
or U36565 (N_36565,N_33118,N_32352);
nand U36566 (N_36566,N_33735,N_32987);
and U36567 (N_36567,N_33433,N_33419);
nor U36568 (N_36568,N_31622,N_33088);
and U36569 (N_36569,N_33059,N_31428);
nor U36570 (N_36570,N_34630,N_30254);
nand U36571 (N_36571,N_32619,N_30781);
or U36572 (N_36572,N_31857,N_30802);
xnor U36573 (N_36573,N_31142,N_32190);
or U36574 (N_36574,N_34064,N_32396);
xor U36575 (N_36575,N_30684,N_32132);
xor U36576 (N_36576,N_32683,N_34099);
nand U36577 (N_36577,N_32248,N_34968);
or U36578 (N_36578,N_32740,N_34566);
nor U36579 (N_36579,N_34561,N_30397);
nand U36580 (N_36580,N_30387,N_33332);
and U36581 (N_36581,N_30671,N_30185);
or U36582 (N_36582,N_32984,N_34285);
nor U36583 (N_36583,N_33526,N_32403);
or U36584 (N_36584,N_31905,N_30358);
nor U36585 (N_36585,N_33270,N_33383);
or U36586 (N_36586,N_34815,N_31316);
and U36587 (N_36587,N_31152,N_33791);
nor U36588 (N_36588,N_30288,N_33652);
nor U36589 (N_36589,N_32261,N_30894);
nand U36590 (N_36590,N_32759,N_34371);
nand U36591 (N_36591,N_34165,N_33343);
nand U36592 (N_36592,N_34209,N_31109);
nor U36593 (N_36593,N_34615,N_31628);
nor U36594 (N_36594,N_33719,N_31306);
or U36595 (N_36595,N_34409,N_32521);
nand U36596 (N_36596,N_32553,N_34324);
and U36597 (N_36597,N_32692,N_34096);
nor U36598 (N_36598,N_34025,N_30384);
and U36599 (N_36599,N_33428,N_34784);
nand U36600 (N_36600,N_33842,N_32485);
nand U36601 (N_36601,N_31129,N_31376);
nor U36602 (N_36602,N_31412,N_32862);
and U36603 (N_36603,N_33307,N_31482);
or U36604 (N_36604,N_30862,N_33948);
xor U36605 (N_36605,N_34470,N_34236);
nand U36606 (N_36606,N_32298,N_34178);
nor U36607 (N_36607,N_33179,N_30927);
or U36608 (N_36608,N_34039,N_30188);
nor U36609 (N_36609,N_32285,N_32122);
or U36610 (N_36610,N_32489,N_34974);
nor U36611 (N_36611,N_30517,N_31403);
and U36612 (N_36612,N_31474,N_31423);
nor U36613 (N_36613,N_32785,N_30199);
nand U36614 (N_36614,N_32143,N_34906);
or U36615 (N_36615,N_33285,N_33246);
and U36616 (N_36616,N_32932,N_31497);
nor U36617 (N_36617,N_33361,N_34385);
nand U36618 (N_36618,N_33528,N_32636);
nor U36619 (N_36619,N_33127,N_31157);
and U36620 (N_36620,N_30133,N_32279);
nand U36621 (N_36621,N_31204,N_31349);
nor U36622 (N_36622,N_33113,N_32992);
nor U36623 (N_36623,N_30726,N_34511);
and U36624 (N_36624,N_31371,N_34913);
nand U36625 (N_36625,N_34791,N_34939);
xnor U36626 (N_36626,N_30022,N_34356);
and U36627 (N_36627,N_32831,N_30605);
nand U36628 (N_36628,N_32755,N_34024);
and U36629 (N_36629,N_33075,N_32466);
nand U36630 (N_36630,N_30390,N_31605);
nand U36631 (N_36631,N_33806,N_32503);
or U36632 (N_36632,N_31041,N_34880);
or U36633 (N_36633,N_30281,N_33323);
nor U36634 (N_36634,N_34588,N_34405);
and U36635 (N_36635,N_31859,N_34517);
and U36636 (N_36636,N_31280,N_32173);
nor U36637 (N_36637,N_33838,N_33336);
and U36638 (N_36638,N_31829,N_33543);
nor U36639 (N_36639,N_34611,N_30788);
nand U36640 (N_36640,N_31876,N_32547);
and U36641 (N_36641,N_30131,N_31900);
and U36642 (N_36642,N_32917,N_31155);
nor U36643 (N_36643,N_31892,N_31877);
nand U36644 (N_36644,N_31463,N_30050);
nand U36645 (N_36645,N_31915,N_30627);
nor U36646 (N_36646,N_33725,N_31904);
and U36647 (N_36647,N_34455,N_33928);
or U36648 (N_36648,N_30468,N_32263);
or U36649 (N_36649,N_33622,N_34185);
nand U36650 (N_36650,N_32400,N_34345);
xor U36651 (N_36651,N_32651,N_32008);
nand U36652 (N_36652,N_32149,N_31774);
nand U36653 (N_36653,N_30248,N_30392);
nor U36654 (N_36654,N_31609,N_32799);
nor U36655 (N_36655,N_31887,N_31328);
or U36656 (N_36656,N_34971,N_30739);
and U36657 (N_36657,N_31314,N_34643);
and U36658 (N_36658,N_33182,N_31356);
xor U36659 (N_36659,N_34179,N_32810);
or U36660 (N_36660,N_31691,N_32793);
xor U36661 (N_36661,N_32773,N_33056);
xor U36662 (N_36662,N_30159,N_30335);
or U36663 (N_36663,N_31471,N_32019);
nand U36664 (N_36664,N_34594,N_30451);
nand U36665 (N_36665,N_32184,N_30179);
nor U36666 (N_36666,N_33698,N_33588);
nor U36667 (N_36667,N_32016,N_30882);
or U36668 (N_36668,N_31652,N_33548);
xor U36669 (N_36669,N_31398,N_31233);
nor U36670 (N_36670,N_33036,N_32027);
xnor U36671 (N_36671,N_33097,N_32829);
or U36672 (N_36672,N_31260,N_34596);
nor U36673 (N_36673,N_33437,N_31318);
nor U36674 (N_36674,N_31365,N_34829);
nor U36675 (N_36675,N_32487,N_33712);
nand U36676 (N_36676,N_33721,N_34816);
nand U36677 (N_36677,N_34641,N_33495);
nand U36678 (N_36678,N_34038,N_32559);
and U36679 (N_36679,N_30769,N_30658);
nand U36680 (N_36680,N_32622,N_34235);
or U36681 (N_36681,N_34541,N_31658);
xor U36682 (N_36682,N_34684,N_32090);
nor U36683 (N_36683,N_34056,N_33411);
or U36684 (N_36684,N_32448,N_34451);
nand U36685 (N_36685,N_34565,N_30730);
nand U36686 (N_36686,N_33845,N_31381);
or U36687 (N_36687,N_32038,N_30760);
and U36688 (N_36688,N_33687,N_31491);
and U36689 (N_36689,N_32407,N_31378);
or U36690 (N_36690,N_30982,N_30917);
and U36691 (N_36691,N_32556,N_32095);
nor U36692 (N_36692,N_32684,N_30491);
and U36693 (N_36693,N_30901,N_33686);
and U36694 (N_36694,N_30246,N_30292);
or U36695 (N_36695,N_31635,N_34942);
and U36696 (N_36696,N_33356,N_33972);
nor U36697 (N_36697,N_33840,N_32774);
nand U36698 (N_36698,N_32180,N_34419);
nor U36699 (N_36699,N_30792,N_34693);
and U36700 (N_36700,N_31989,N_34159);
nand U36701 (N_36701,N_30116,N_34172);
nor U36702 (N_36702,N_32355,N_31216);
xor U36703 (N_36703,N_32688,N_31479);
or U36704 (N_36704,N_31878,N_30024);
nand U36705 (N_36705,N_32087,N_30323);
and U36706 (N_36706,N_31789,N_34269);
and U36707 (N_36707,N_32472,N_30859);
and U36708 (N_36708,N_33694,N_30548);
nor U36709 (N_36709,N_32177,N_33804);
nand U36710 (N_36710,N_34707,N_31581);
nor U36711 (N_36711,N_30352,N_31545);
nor U36712 (N_36712,N_34435,N_31424);
or U36713 (N_36713,N_31213,N_34826);
nand U36714 (N_36714,N_31767,N_34120);
and U36715 (N_36715,N_30464,N_30053);
or U36716 (N_36716,N_34637,N_34790);
nand U36717 (N_36717,N_32394,N_33967);
nor U36718 (N_36718,N_30898,N_34987);
or U36719 (N_36719,N_31791,N_33660);
and U36720 (N_36720,N_32418,N_30194);
and U36721 (N_36721,N_34769,N_30289);
nand U36722 (N_36722,N_34613,N_33389);
nand U36723 (N_36723,N_33532,N_30690);
or U36724 (N_36724,N_32330,N_30983);
nor U36725 (N_36725,N_33009,N_33813);
and U36726 (N_36726,N_34128,N_31466);
nor U36727 (N_36727,N_33717,N_34598);
and U36728 (N_36728,N_34168,N_30480);
or U36729 (N_36729,N_32872,N_32738);
nand U36730 (N_36730,N_34584,N_30720);
nor U36731 (N_36731,N_30613,N_30372);
nand U36732 (N_36732,N_30437,N_30593);
nand U36733 (N_36733,N_34620,N_34386);
nand U36734 (N_36734,N_31974,N_33243);
nand U36735 (N_36735,N_32718,N_33379);
or U36736 (N_36736,N_34844,N_32495);
nor U36737 (N_36737,N_30873,N_32384);
or U36738 (N_36738,N_30948,N_32321);
nand U36739 (N_36739,N_34262,N_34951);
nand U36740 (N_36740,N_33990,N_30025);
nand U36741 (N_36741,N_34272,N_33780);
and U36742 (N_36742,N_32930,N_32668);
nand U36743 (N_36743,N_32317,N_30014);
nor U36744 (N_36744,N_32035,N_32020);
nor U36745 (N_36745,N_33315,N_33971);
nor U36746 (N_36746,N_34723,N_30837);
nor U36747 (N_36747,N_32094,N_30276);
nor U36748 (N_36748,N_33792,N_33577);
nor U36749 (N_36749,N_30718,N_30441);
or U36750 (N_36750,N_34486,N_31893);
nor U36751 (N_36751,N_32463,N_32176);
nand U36752 (N_36752,N_30207,N_33692);
or U36753 (N_36753,N_30421,N_32937);
nor U36754 (N_36754,N_34759,N_31645);
and U36755 (N_36755,N_34933,N_33131);
nor U36756 (N_36756,N_32697,N_34203);
xor U36757 (N_36757,N_32608,N_32348);
nor U36758 (N_36758,N_32519,N_30729);
nor U36759 (N_36759,N_31165,N_32921);
or U36760 (N_36760,N_33439,N_31249);
or U36761 (N_36761,N_33955,N_34558);
or U36762 (N_36762,N_31685,N_34977);
nand U36763 (N_36763,N_34730,N_31078);
nor U36764 (N_36764,N_30231,N_30621);
or U36765 (N_36765,N_32350,N_32084);
nand U36766 (N_36766,N_30539,N_32501);
and U36767 (N_36767,N_34445,N_31711);
and U36768 (N_36768,N_30712,N_32369);
or U36769 (N_36769,N_31899,N_31166);
nand U36770 (N_36770,N_34837,N_32523);
and U36771 (N_36771,N_34841,N_33623);
nand U36772 (N_36772,N_33259,N_33590);
and U36773 (N_36773,N_30447,N_34658);
xnor U36774 (N_36774,N_32602,N_30583);
or U36775 (N_36775,N_30970,N_33458);
nand U36776 (N_36776,N_32455,N_32770);
or U36777 (N_36777,N_33925,N_30523);
xnor U36778 (N_36778,N_31737,N_32110);
nor U36779 (N_36779,N_33145,N_30415);
or U36780 (N_36780,N_34224,N_33890);
xor U36781 (N_36781,N_33144,N_33422);
and U36782 (N_36782,N_33953,N_34963);
or U36783 (N_36783,N_33005,N_33392);
nand U36784 (N_36784,N_32475,N_31883);
nand U36785 (N_36785,N_33861,N_34635);
nor U36786 (N_36786,N_33496,N_34812);
and U36787 (N_36787,N_30184,N_32329);
or U36788 (N_36788,N_31800,N_34758);
nand U36789 (N_36789,N_31913,N_33555);
or U36790 (N_36790,N_30551,N_31594);
nor U36791 (N_36791,N_31604,N_30202);
or U36792 (N_36792,N_31183,N_33269);
or U36793 (N_36793,N_30640,N_32642);
or U36794 (N_36794,N_34548,N_31578);
and U36795 (N_36795,N_34066,N_30783);
or U36796 (N_36796,N_32726,N_31732);
or U36797 (N_36797,N_33835,N_30461);
and U36798 (N_36798,N_32385,N_33014);
or U36799 (N_36799,N_32041,N_31766);
xor U36800 (N_36800,N_33015,N_32364);
or U36801 (N_36801,N_34513,N_32764);
and U36802 (N_36802,N_34467,N_33803);
nor U36803 (N_36803,N_31308,N_32666);
and U36804 (N_36804,N_33567,N_32908);
or U36805 (N_36805,N_31509,N_32376);
nand U36806 (N_36806,N_33882,N_33013);
xnor U36807 (N_36807,N_31671,N_31309);
xor U36808 (N_36808,N_31312,N_34080);
and U36809 (N_36809,N_34326,N_34982);
xnor U36810 (N_36810,N_31837,N_34116);
and U36811 (N_36811,N_32444,N_34162);
xor U36812 (N_36812,N_30120,N_32341);
or U36813 (N_36813,N_30764,N_31108);
nand U36814 (N_36814,N_30454,N_31375);
nand U36815 (N_36815,N_31450,N_34033);
nand U36816 (N_36816,N_30860,N_31803);
nand U36817 (N_36817,N_30388,N_33606);
and U36818 (N_36818,N_33832,N_34342);
or U36819 (N_36819,N_33222,N_30645);
and U36820 (N_36820,N_34108,N_33294);
or U36821 (N_36821,N_33354,N_33801);
nor U36822 (N_36822,N_30079,N_31740);
nor U36823 (N_36823,N_34460,N_30285);
and U36824 (N_36824,N_30928,N_32980);
or U36825 (N_36825,N_32320,N_34932);
nand U36826 (N_36826,N_31122,N_30221);
nor U36827 (N_36827,N_32166,N_31058);
and U36828 (N_36828,N_33276,N_32940);
and U36829 (N_36829,N_34001,N_31350);
and U36830 (N_36830,N_30677,N_32652);
nor U36831 (N_36831,N_32640,N_30824);
or U36832 (N_36832,N_33244,N_34143);
or U36833 (N_36833,N_31202,N_30683);
xor U36834 (N_36834,N_31770,N_31590);
nand U36835 (N_36835,N_34090,N_34717);
or U36836 (N_36836,N_34079,N_31616);
nor U36837 (N_36837,N_32941,N_33291);
and U36838 (N_36838,N_34415,N_30186);
or U36839 (N_36839,N_34113,N_33572);
and U36840 (N_36840,N_32067,N_33286);
nand U36841 (N_36841,N_31788,N_34564);
nand U36842 (N_36842,N_30614,N_30119);
or U36843 (N_36843,N_30844,N_30510);
nand U36844 (N_36844,N_31042,N_31809);
nor U36845 (N_36845,N_33515,N_31557);
nand U36846 (N_36846,N_33497,N_33000);
xnor U36847 (N_36847,N_30324,N_33421);
nor U36848 (N_36848,N_30785,N_31619);
and U36849 (N_36849,N_30062,N_32256);
nor U36850 (N_36850,N_34259,N_30616);
nand U36851 (N_36851,N_30778,N_30969);
nand U36852 (N_36852,N_33663,N_32405);
nor U36853 (N_36853,N_34514,N_30823);
xnor U36854 (N_36854,N_31418,N_32169);
nand U36855 (N_36855,N_31034,N_32081);
nand U36856 (N_36856,N_34833,N_30172);
or U36857 (N_36857,N_33810,N_30749);
and U36858 (N_36858,N_34340,N_34520);
xor U36859 (N_36859,N_33939,N_32698);
xor U36860 (N_36860,N_34406,N_33358);
and U36861 (N_36861,N_32093,N_30346);
or U36862 (N_36862,N_31370,N_34394);
or U36863 (N_36863,N_33201,N_33296);
and U36864 (N_36864,N_33147,N_30072);
nor U36865 (N_36865,N_31640,N_32224);
or U36866 (N_36866,N_33197,N_31483);
nand U36867 (N_36867,N_31598,N_33196);
nand U36868 (N_36868,N_34540,N_31077);
and U36869 (N_36869,N_31348,N_30303);
nor U36870 (N_36870,N_33212,N_34934);
nand U36871 (N_36871,N_33151,N_33146);
nor U36872 (N_36872,N_31849,N_33539);
or U36873 (N_36873,N_30924,N_30941);
and U36874 (N_36874,N_34973,N_33404);
or U36875 (N_36875,N_31558,N_30412);
nand U36876 (N_36876,N_34306,N_30370);
and U36877 (N_36877,N_30325,N_32346);
or U36878 (N_36878,N_32809,N_32439);
nor U36879 (N_36879,N_30351,N_33357);
nand U36880 (N_36880,N_31750,N_32906);
and U36881 (N_36881,N_33676,N_34568);
or U36882 (N_36882,N_31069,N_31792);
nand U36883 (N_36883,N_32630,N_33338);
or U36884 (N_36884,N_34988,N_32841);
nor U36885 (N_36885,N_34094,N_34602);
xnor U36886 (N_36886,N_30486,N_34027);
or U36887 (N_36887,N_31552,N_32068);
nor U36888 (N_36888,N_34226,N_33167);
nor U36889 (N_36889,N_31656,N_34608);
nand U36890 (N_36890,N_32757,N_34868);
and U36891 (N_36891,N_30615,N_33333);
and U36892 (N_36892,N_30298,N_31907);
and U36893 (N_36893,N_33359,N_34666);
or U36894 (N_36894,N_33706,N_32187);
xor U36895 (N_36895,N_33872,N_33095);
nand U36896 (N_36896,N_31061,N_34065);
nor U36897 (N_36897,N_31526,N_31188);
and U36898 (N_36898,N_33208,N_32389);
nand U36899 (N_36899,N_34424,N_31422);
xnor U36900 (N_36900,N_31134,N_30639);
nor U36901 (N_36901,N_31211,N_32284);
and U36902 (N_36902,N_31790,N_34197);
nor U36903 (N_36903,N_33415,N_33903);
and U36904 (N_36904,N_32518,N_32853);
nand U36905 (N_36905,N_30283,N_30741);
and U36906 (N_36906,N_32968,N_32236);
or U36907 (N_36907,N_33115,N_34945);
nor U36908 (N_36908,N_34223,N_31940);
nand U36909 (N_36909,N_31624,N_31162);
nor U36910 (N_36910,N_30403,N_30026);
and U36911 (N_36911,N_33459,N_32612);
nand U36912 (N_36912,N_31832,N_34757);
or U36913 (N_36913,N_33746,N_30972);
nand U36914 (N_36914,N_34395,N_30109);
or U36915 (N_36915,N_34544,N_30455);
nor U36916 (N_36916,N_34652,N_34740);
and U36917 (N_36917,N_32775,N_33503);
nand U36918 (N_36918,N_32205,N_32957);
or U36919 (N_36919,N_31909,N_34671);
nor U36920 (N_36920,N_34252,N_32884);
nor U36921 (N_36921,N_31214,N_32762);
and U36922 (N_36922,N_34472,N_33683);
and U36923 (N_36923,N_30405,N_33868);
and U36924 (N_36924,N_34115,N_33342);
or U36925 (N_36925,N_34669,N_34581);
xnor U36926 (N_36926,N_32515,N_31967);
nor U36927 (N_36927,N_34787,N_30915);
nand U36928 (N_36928,N_33611,N_34946);
or U36929 (N_36929,N_30507,N_31093);
nor U36930 (N_36930,N_34081,N_31894);
nor U36931 (N_36931,N_33093,N_33992);
or U36932 (N_36932,N_32312,N_31411);
nand U36933 (N_36933,N_33111,N_30905);
nor U36934 (N_36934,N_34715,N_32551);
nand U36935 (N_36935,N_32062,N_31103);
nor U36936 (N_36936,N_32797,N_30650);
and U36937 (N_36937,N_32028,N_33447);
and U36938 (N_36938,N_33139,N_34384);
nor U36939 (N_36939,N_32304,N_30612);
and U36940 (N_36940,N_34885,N_31840);
nor U36941 (N_36941,N_34292,N_32103);
and U36942 (N_36942,N_30143,N_32148);
nand U36943 (N_36943,N_33049,N_30734);
nor U36944 (N_36944,N_33995,N_30306);
xnor U36945 (N_36945,N_34774,N_30547);
nand U36946 (N_36946,N_34126,N_34023);
or U36947 (N_36947,N_30228,N_33213);
nor U36948 (N_36948,N_31088,N_33596);
and U36949 (N_36949,N_32573,N_30759);
or U36950 (N_36950,N_32178,N_32105);
or U36951 (N_36951,N_34959,N_33233);
xnor U36952 (N_36952,N_33008,N_33058);
nand U36953 (N_36953,N_32002,N_31864);
or U36954 (N_36954,N_34744,N_33499);
nor U36955 (N_36955,N_31755,N_31445);
or U36956 (N_36956,N_32436,N_30636);
or U36957 (N_36957,N_34691,N_30884);
nor U36958 (N_36958,N_33054,N_34986);
nand U36959 (N_36959,N_30706,N_32450);
nor U36960 (N_36960,N_34082,N_32168);
nor U36961 (N_36961,N_31414,N_34509);
nand U36962 (N_36962,N_33880,N_34903);
and U36963 (N_36963,N_30368,N_31816);
nand U36964 (N_36964,N_34246,N_31806);
xnor U36965 (N_36965,N_32843,N_30081);
and U36966 (N_36966,N_32699,N_34563);
nor U36967 (N_36967,N_34391,N_33781);
nand U36968 (N_36968,N_30452,N_33750);
xnor U36969 (N_36969,N_32907,N_30773);
and U36970 (N_36970,N_34770,N_31891);
nand U36971 (N_36971,N_33745,N_32054);
and U36972 (N_36972,N_30302,N_31090);
nor U36973 (N_36973,N_34131,N_30414);
and U36974 (N_36974,N_34586,N_31851);
nor U36975 (N_36975,N_31595,N_31433);
and U36976 (N_36976,N_31274,N_33019);
and U36977 (N_36977,N_30272,N_31060);
and U36978 (N_36978,N_32469,N_34103);
nor U36979 (N_36979,N_30624,N_33039);
nor U36980 (N_36980,N_33312,N_34042);
xnor U36981 (N_36981,N_33851,N_33830);
nor U36982 (N_36982,N_32296,N_31769);
nand U36983 (N_36983,N_34626,N_34000);
or U36984 (N_36984,N_32850,N_34362);
nor U36985 (N_36985,N_32988,N_30381);
or U36986 (N_36986,N_31021,N_31361);
nand U36987 (N_36987,N_31688,N_33051);
or U36988 (N_36988,N_32003,N_30211);
nand U36989 (N_36989,N_30775,N_34338);
or U36990 (N_36990,N_33254,N_30252);
and U36991 (N_36991,N_33888,N_31258);
nand U36992 (N_36992,N_32118,N_32648);
nor U36993 (N_36993,N_30831,N_34245);
or U36994 (N_36994,N_34059,N_31197);
and U36995 (N_36995,N_30070,N_33225);
nand U36996 (N_36996,N_31554,N_30956);
nor U36997 (N_36997,N_31664,N_32247);
nand U36998 (N_36998,N_34408,N_30477);
or U36999 (N_36999,N_34194,N_33303);
nor U37000 (N_37000,N_31998,N_31897);
and U37001 (N_37001,N_30893,N_31070);
and U37002 (N_37002,N_30503,N_33571);
nor U37003 (N_37003,N_31360,N_31592);
and U37004 (N_37004,N_30016,N_30474);
nand U37005 (N_37005,N_31107,N_32765);
nand U37006 (N_37006,N_31579,N_30060);
and U37007 (N_37007,N_30229,N_33893);
or U37008 (N_37008,N_32386,N_31710);
nor U37009 (N_37009,N_30380,N_33242);
and U37010 (N_37010,N_30585,N_31179);
and U37011 (N_37011,N_34958,N_30212);
xnor U37012 (N_37012,N_33843,N_30881);
and U37013 (N_37013,N_33766,N_32874);
nor U37014 (N_37014,N_30992,N_33647);
and U37015 (N_37015,N_34577,N_33162);
and U37016 (N_37016,N_30407,N_33796);
nand U37017 (N_37017,N_33227,N_33264);
and U37018 (N_37018,N_32963,N_30821);
nand U37019 (N_37019,N_32517,N_31930);
nand U37020 (N_37020,N_34714,N_32522);
and U37021 (N_37021,N_34891,N_30499);
nor U37022 (N_37022,N_34754,N_33363);
or U37023 (N_37023,N_32886,N_30422);
nor U37024 (N_37024,N_32303,N_31772);
or U37025 (N_37025,N_32294,N_31798);
nor U37026 (N_37026,N_32737,N_30896);
nand U37027 (N_37027,N_30743,N_30564);
nand U37028 (N_37028,N_31744,N_33662);
xnor U37029 (N_37029,N_34220,N_31742);
nand U37030 (N_37030,N_31250,N_34834);
xor U37031 (N_37031,N_33037,N_32508);
or U37032 (N_37032,N_30940,N_32335);
or U37033 (N_37033,N_31572,N_32065);
and U37034 (N_37034,N_34449,N_34651);
nand U37035 (N_37035,N_31057,N_34708);
or U37036 (N_37036,N_33865,N_34587);
and U37037 (N_37037,N_32822,N_31475);
and U37038 (N_37038,N_31264,N_31405);
or U37039 (N_37039,N_34519,N_30085);
and U37040 (N_37040,N_30643,N_33714);
nor U37041 (N_37041,N_31408,N_30100);
and U37042 (N_37042,N_33946,N_30619);
xor U37043 (N_37043,N_33994,N_34330);
nand U37044 (N_37044,N_30755,N_30817);
or U37045 (N_37045,N_31518,N_33904);
and U37046 (N_37046,N_34434,N_32549);
or U37047 (N_37047,N_32995,N_30973);
or U37048 (N_37048,N_34993,N_31914);
nand U37049 (N_37049,N_31437,N_30651);
and U37050 (N_37050,N_32626,N_33300);
nand U37051 (N_37051,N_31610,N_34888);
nand U37052 (N_37052,N_32270,N_32537);
and U37053 (N_37053,N_30398,N_32431);
and U37054 (N_37054,N_34683,N_32226);
and U37055 (N_37055,N_33732,N_34229);
and U37056 (N_37056,N_33911,N_34310);
and U37057 (N_37057,N_30705,N_33416);
or U37058 (N_37058,N_34471,N_34380);
nand U37059 (N_37059,N_32824,N_30814);
nand U37060 (N_37060,N_33316,N_32798);
nor U37061 (N_37061,N_34845,N_33716);
and U37062 (N_37062,N_34438,N_30478);
nand U37063 (N_37063,N_31359,N_33670);
xor U37064 (N_37064,N_31449,N_34947);
or U37065 (N_37065,N_30123,N_30851);
and U37066 (N_37066,N_32359,N_34289);
nor U37067 (N_37067,N_30518,N_30394);
xor U37068 (N_37068,N_31633,N_34152);
or U37069 (N_37069,N_32447,N_33187);
xnor U37070 (N_37070,N_30374,N_32283);
nand U37071 (N_37071,N_33391,N_34425);
nor U37072 (N_37072,N_33747,N_32223);
or U37073 (N_37073,N_32451,N_32163);
and U37074 (N_37074,N_33603,N_33399);
nor U37075 (N_37075,N_30375,N_32628);
or U37076 (N_37076,N_31293,N_34662);
xnor U37077 (N_37077,N_30017,N_34009);
nand U37078 (N_37078,N_30668,N_31286);
or U37079 (N_37079,N_32771,N_30355);
nor U37080 (N_37080,N_32498,N_33536);
nor U37081 (N_37081,N_33199,N_34975);
nand U37082 (N_37082,N_30472,N_30714);
nand U37083 (N_37083,N_33877,N_34810);
nor U37084 (N_37084,N_34402,N_33508);
nand U37085 (N_37085,N_32974,N_34211);
or U37086 (N_37086,N_33069,N_31272);
nor U37087 (N_37087,N_32600,N_33451);
nand U37088 (N_37088,N_34319,N_30756);
or U37089 (N_37089,N_32911,N_33599);
and U37090 (N_37090,N_34117,N_30110);
nand U37091 (N_37091,N_34212,N_31704);
and U37092 (N_37092,N_34374,N_32845);
nor U37093 (N_37093,N_31808,N_30682);
nor U37094 (N_37094,N_32124,N_34366);
nor U37095 (N_37095,N_31032,N_31690);
or U37096 (N_37096,N_34501,N_34173);
nor U37097 (N_37097,N_32108,N_31527);
nor U37098 (N_37098,N_32220,N_33520);
and U37099 (N_37099,N_30767,N_33267);
xor U37100 (N_37100,N_34218,N_31629);
nor U37101 (N_37101,N_30938,N_33821);
or U37102 (N_37102,N_34782,N_34861);
and U37103 (N_37103,N_34873,N_31013);
or U37104 (N_37104,N_34847,N_33854);
nand U37105 (N_37105,N_30446,N_30007);
nand U37106 (N_37106,N_32150,N_31364);
or U37107 (N_37107,N_31147,N_30215);
or U37108 (N_37108,N_31315,N_32510);
nand U37109 (N_37109,N_34949,N_30418);
xor U37110 (N_37110,N_30779,N_30687);
and U37111 (N_37111,N_33263,N_32680);
or U37112 (N_37112,N_34950,N_32018);
xor U37113 (N_37113,N_33899,N_30929);
nor U37114 (N_37114,N_33808,N_33400);
xor U37115 (N_37115,N_30222,N_34315);
and U37116 (N_37116,N_31281,N_30909);
or U37117 (N_37117,N_32734,N_34013);
or U37118 (N_37118,N_34180,N_31589);
and U37119 (N_37119,N_31890,N_34357);
or U37120 (N_37120,N_30012,N_30845);
nor U37121 (N_37121,N_30316,N_31327);
nand U37122 (N_37122,N_30578,N_31975);
or U37123 (N_37123,N_33709,N_32077);
or U37124 (N_37124,N_34830,N_34567);
nor U37125 (N_37125,N_33432,N_32219);
nor U37126 (N_37126,N_33169,N_34591);
xnor U37127 (N_37127,N_31564,N_34654);
nand U37128 (N_37128,N_31567,N_32354);
xnor U37129 (N_37129,N_34101,N_31181);
xor U37130 (N_37130,N_34248,N_32796);
and U37131 (N_37131,N_34036,N_34549);
and U37132 (N_37132,N_34972,N_30293);
nand U37133 (N_37133,N_34980,N_34772);
nand U37134 (N_37134,N_34796,N_34392);
nor U37135 (N_37135,N_33007,N_33417);
nand U37136 (N_37136,N_31938,N_31248);
and U37137 (N_37137,N_31537,N_33773);
nor U37138 (N_37138,N_33892,N_30216);
nor U37139 (N_37139,N_33991,N_32056);
xnor U37140 (N_37140,N_33138,N_30460);
or U37141 (N_37141,N_32903,N_34937);
xor U37142 (N_37142,N_31815,N_31593);
or U37143 (N_37143,N_33335,N_31298);
or U37144 (N_37144,N_30122,N_34225);
xnor U37145 (N_37145,N_31773,N_30340);
xnor U37146 (N_37146,N_32748,N_32816);
or U37147 (N_37147,N_34412,N_34981);
or U37148 (N_37148,N_30417,N_31668);
or U37149 (N_37149,N_34261,N_32790);
and U37150 (N_37150,N_34106,N_30313);
and U37151 (N_37151,N_32288,N_32596);
and U37152 (N_37152,N_30492,N_32787);
nand U37153 (N_37153,N_30361,N_34146);
nor U37154 (N_37154,N_30271,N_31631);
nand U37155 (N_37155,N_34835,N_32047);
or U37156 (N_37156,N_34493,N_32649);
nand U37157 (N_37157,N_32996,N_33659);
xnor U37158 (N_37158,N_30694,N_30754);
and U37159 (N_37159,N_30242,N_31860);
and U37160 (N_37160,N_33407,N_31973);
nor U37161 (N_37161,N_31161,N_34164);
nor U37162 (N_37162,N_30903,N_33381);
and U37163 (N_37163,N_34221,N_34015);
and U37164 (N_37164,N_34851,N_33524);
and U37165 (N_37165,N_30270,N_30888);
and U37166 (N_37166,N_32781,N_32700);
nor U37167 (N_37167,N_34174,N_32865);
nor U37168 (N_37168,N_30855,N_30540);
nor U37169 (N_37169,N_32107,N_31123);
nor U37170 (N_37170,N_34067,N_33224);
nand U37171 (N_37171,N_30103,N_33914);
nor U37172 (N_37172,N_34526,N_33770);
nand U37173 (N_37173,N_32276,N_34378);
nor U37174 (N_37174,N_31933,N_33999);
or U37175 (N_37175,N_31959,N_32892);
and U37176 (N_37176,N_32007,N_34768);
and U37177 (N_37177,N_34729,N_30808);
or U37178 (N_37178,N_31743,N_30719);
nand U37179 (N_37179,N_33089,N_34795);
and U37180 (N_37180,N_30386,N_33658);
nand U37181 (N_37181,N_32915,N_33968);
nor U37182 (N_37182,N_32777,N_33651);
and U37183 (N_37183,N_32422,N_33505);
nor U37184 (N_37184,N_33175,N_31046);
nor U37185 (N_37185,N_32425,N_32896);
nor U37186 (N_37186,N_33552,N_31586);
or U37187 (N_37187,N_31277,N_32387);
nor U37188 (N_37188,N_30240,N_32467);
nand U37189 (N_37189,N_31681,N_34618);
and U37190 (N_37190,N_31873,N_33544);
and U37191 (N_37191,N_31496,N_30003);
nand U37192 (N_37192,N_34560,N_34543);
and U37193 (N_37193,N_33702,N_33556);
and U37194 (N_37194,N_32315,N_31143);
nor U37195 (N_37195,N_31707,N_32109);
nor U37196 (N_37196,N_30505,N_31736);
or U37197 (N_37197,N_32860,N_34084);
nand U37198 (N_37198,N_31702,N_33262);
nor U37199 (N_37199,N_33619,N_31871);
or U37200 (N_37200,N_31146,N_32586);
or U37201 (N_37201,N_31073,N_32072);
nor U37202 (N_37202,N_34503,N_32564);
and U37203 (N_37203,N_34992,N_30448);
and U37204 (N_37204,N_34158,N_32611);
nor U37205 (N_37205,N_31971,N_31098);
or U37206 (N_37206,N_33306,N_34752);
nor U37207 (N_37207,N_33740,N_33973);
xor U37208 (N_37208,N_32125,N_30717);
and U37209 (N_37209,N_33529,N_34447);
or U37210 (N_37210,N_32208,N_31160);
nand U37211 (N_37211,N_33398,N_33642);
and U37212 (N_37212,N_31771,N_34583);
nand U37213 (N_37213,N_33402,N_34222);
and U37214 (N_37214,N_33617,N_33476);
and U37215 (N_37215,N_30553,N_34813);
nand U37216 (N_37216,N_34546,N_30253);
xnor U37217 (N_37217,N_33382,N_34609);
or U37218 (N_37218,N_31156,N_34786);
nand U37219 (N_37219,N_31724,N_34452);
nand U37220 (N_37220,N_32916,N_30487);
and U37221 (N_37221,N_30800,N_32152);
or U37222 (N_37222,N_30309,N_32504);
and U37223 (N_37223,N_32866,N_30692);
or U37224 (N_37224,N_33912,N_33752);
and U37225 (N_37225,N_33909,N_33293);
or U37226 (N_37226,N_33736,N_31674);
nor U37227 (N_37227,N_32144,N_30191);
or U37228 (N_37228,N_33023,N_31853);
xnor U37229 (N_37229,N_32525,N_34302);
or U37230 (N_37230,N_32171,N_34767);
or U37231 (N_37231,N_32998,N_34111);
nor U37232 (N_37232,N_30132,N_31730);
or U37233 (N_37233,N_33678,N_32767);
nor U37234 (N_37234,N_31055,N_30030);
nand U37235 (N_37235,N_31212,N_30757);
or U37236 (N_37236,N_33229,N_31802);
nor U37237 (N_37237,N_31128,N_33200);
nand U37238 (N_37238,N_32975,N_33079);
or U37239 (N_37239,N_30218,N_34725);
nand U37240 (N_37240,N_34695,N_32433);
nor U37241 (N_37241,N_32280,N_31279);
or U37242 (N_37242,N_34994,N_30890);
and U37243 (N_37243,N_33455,N_33586);
xnor U37244 (N_37244,N_32955,N_34283);
or U37245 (N_37245,N_32671,N_32870);
or U37246 (N_37246,N_34556,N_33042);
nand U37247 (N_37247,N_32971,N_30602);
nand U37248 (N_37248,N_32687,N_33519);
and U37249 (N_37249,N_33150,N_31795);
and U37250 (N_37250,N_32185,N_31953);
nor U37251 (N_37251,N_30770,N_32538);
and U37252 (N_37252,N_30124,N_30665);
nand U37253 (N_37253,N_32154,N_30214);
xnor U37254 (N_37254,N_34935,N_32410);
or U37255 (N_37255,N_31962,N_30870);
xor U37256 (N_37256,N_33248,N_31787);
or U37257 (N_37257,N_33887,N_32951);
xnor U37258 (N_37258,N_34274,N_32782);
nor U37259 (N_37259,N_32167,N_32207);
xnor U37260 (N_37260,N_33261,N_31075);
nor U37261 (N_37261,N_34701,N_30069);
or U37262 (N_37262,N_31301,N_33549);
xnor U37263 (N_37263,N_33656,N_31574);
xnor U37264 (N_37264,N_30535,N_32164);
nand U37265 (N_37265,N_32092,N_30402);
or U37266 (N_37266,N_34337,N_34432);
or U37267 (N_37267,N_30338,N_33231);
and U37268 (N_37268,N_30498,N_32112);
nand U37269 (N_37269,N_33070,N_32563);
or U37270 (N_37270,N_30931,N_31028);
and U37271 (N_37271,N_32366,N_34661);
nor U37272 (N_37272,N_34699,N_31262);
and U37273 (N_37273,N_33507,N_32456);
or U37274 (N_37274,N_32949,N_34863);
and U37275 (N_37275,N_31879,N_34802);
nor U37276 (N_37276,N_30319,N_32802);
or U37277 (N_37277,N_31159,N_32876);
or U37278 (N_37278,N_33450,N_30363);
nand U37279 (N_37279,N_32677,N_34700);
or U37280 (N_37280,N_33879,N_30947);
nor U37281 (N_37281,N_31804,N_30921);
nor U37282 (N_37282,N_34843,N_31087);
nand U37283 (N_37283,N_32416,N_30436);
nand U37284 (N_37284,N_33166,N_31961);
xnor U37285 (N_37285,N_34537,N_30955);
or U37286 (N_37286,N_34370,N_32991);
and U37287 (N_37287,N_30504,N_32593);
nor U37288 (N_37288,N_31553,N_30328);
nand U37289 (N_37289,N_33870,N_33790);
nand U37290 (N_37290,N_34061,N_30958);
nand U37291 (N_37291,N_32837,N_32520);
nand U37292 (N_37292,N_33748,N_32155);
xor U37293 (N_37293,N_33043,N_34523);
nor U37294 (N_37294,N_30223,N_34333);
xor U37295 (N_37295,N_31994,N_34323);
or U37296 (N_37296,N_33341,N_30936);
nand U37297 (N_37297,N_30957,N_31955);
nor U37298 (N_37298,N_33474,N_30265);
nor U37299 (N_37299,N_30141,N_32653);
nor U37300 (N_37300,N_30949,N_30466);
nor U37301 (N_37301,N_32961,N_34709);
xor U37302 (N_37302,N_34244,N_30878);
nand U37303 (N_37303,N_33424,N_31436);
nor U37304 (N_37304,N_33395,N_32113);
and U37305 (N_37305,N_30569,N_34739);
and U37306 (N_37306,N_34442,N_33836);
nor U37307 (N_37307,N_31288,N_34580);
or U37308 (N_37308,N_31534,N_33546);
or U37309 (N_37309,N_31613,N_34063);
xor U37310 (N_37310,N_33873,N_32200);
nor U37311 (N_37311,N_30600,N_32956);
nor U37312 (N_37312,N_34878,N_33482);
and U37313 (N_37313,N_32368,N_31064);
nor U37314 (N_37314,N_32381,N_33401);
nand U37315 (N_37315,N_30964,N_31355);
or U37316 (N_37316,N_30604,N_34494);
nor U37317 (N_37317,N_32259,N_31067);
xor U37318 (N_37318,N_32483,N_34002);
nand U37319 (N_37319,N_33331,N_32703);
or U37320 (N_37320,N_32392,N_31068);
nand U37321 (N_37321,N_33466,N_31176);
or U37322 (N_37322,N_32192,N_34114);
xor U37323 (N_37323,N_30657,N_31135);
or U37324 (N_37324,N_32482,N_31763);
and U37325 (N_37325,N_31383,N_30777);
nand U37326 (N_37326,N_33219,N_30035);
and U37327 (N_37327,N_31888,N_31186);
or U37328 (N_37328,N_34368,N_31493);
and U37329 (N_37329,N_30826,N_32719);
nor U37330 (N_37330,N_33273,N_30724);
and U37331 (N_37331,N_34689,N_30489);
nand U37332 (N_37332,N_31647,N_30282);
nor U37333 (N_37333,N_33755,N_30450);
or U37334 (N_37334,N_33550,N_30906);
nand U37335 (N_37335,N_30456,N_33378);
nand U37336 (N_37336,N_34820,N_33820);
nor U37337 (N_37337,N_30544,N_31218);
and U37338 (N_37338,N_32631,N_34188);
and U37339 (N_37339,N_31380,N_33280);
or U37340 (N_37340,N_31868,N_31027);
and U37341 (N_37341,N_32039,N_32788);
and U37342 (N_37342,N_32291,N_31606);
and U37343 (N_37343,N_30373,N_33585);
nor U37344 (N_37344,N_33844,N_30935);
nor U37345 (N_37345,N_33327,N_32808);
and U37346 (N_37346,N_31644,N_33148);
and U37347 (N_37347,N_33634,N_31720);
xnor U37348 (N_37348,N_34781,N_33041);
nand U37349 (N_37349,N_31673,N_30435);
nor U37350 (N_37350,N_32904,N_32468);
nor U37351 (N_37351,N_30278,N_32838);
nand U37352 (N_37352,N_30027,N_33871);
nor U37353 (N_37353,N_30106,N_31784);
nor U37354 (N_37354,N_31031,N_33889);
or U37355 (N_37355,N_32858,N_31846);
nand U37356 (N_37356,N_34733,N_32550);
or U37357 (N_37357,N_33309,N_32736);
or U37358 (N_37358,N_33364,N_31880);
nor U37359 (N_37359,N_33112,N_31053);
xor U37360 (N_37360,N_30847,N_30167);
xnor U37361 (N_37361,N_33563,N_32136);
or U37362 (N_37362,N_31382,N_32535);
or U37363 (N_37363,N_32805,N_34430);
and U37364 (N_37364,N_34073,N_32741);
and U37365 (N_37365,N_31255,N_34817);
nand U37366 (N_37366,N_34697,N_34458);
xnor U37367 (N_37367,N_34305,N_33052);
xor U37368 (N_37368,N_31761,N_34597);
xnor U37369 (N_37369,N_31830,N_34504);
nand U37370 (N_37370,N_30843,N_30015);
or U37371 (N_37371,N_30744,N_30689);
xor U37372 (N_37372,N_31017,N_31544);
and U37373 (N_37373,N_34632,N_34365);
or U37374 (N_37374,N_33648,N_32252);
or U37375 (N_37375,N_31827,N_31484);
and U37376 (N_37376,N_34756,N_34190);
and U37377 (N_37377,N_34742,N_34624);
nor U37378 (N_37378,N_31503,N_34389);
nand U37379 (N_37379,N_33239,N_33397);
nor U37380 (N_37380,N_31573,N_33894);
nor U37381 (N_37381,N_34134,N_31646);
or U37382 (N_37382,N_34350,N_31875);
or U37383 (N_37383,N_30475,N_30801);
nand U37384 (N_37384,N_32162,N_30020);
or U37385 (N_37385,N_30753,N_31867);
xor U37386 (N_37386,N_32479,N_33600);
or U37387 (N_37387,N_33774,N_30768);
and U37388 (N_37388,N_33452,N_32727);
or U37389 (N_37389,N_30078,N_30104);
nand U37390 (N_37390,N_31638,N_31819);
or U37391 (N_37391,N_31666,N_31939);
xor U37392 (N_37392,N_31764,N_30974);
xnor U37393 (N_37393,N_34311,N_34690);
or U37394 (N_37394,N_31373,N_33214);
nor U37395 (N_37395,N_34118,N_34529);
nor U37396 (N_37396,N_32722,N_32497);
and U37397 (N_37397,N_31582,N_31201);
nand U37398 (N_37398,N_33579,N_33366);
nand U37399 (N_37399,N_32868,N_32069);
nor U37400 (N_37400,N_33081,N_31321);
nand U37401 (N_37401,N_31369,N_30679);
nand U37402 (N_37402,N_32768,N_31267);
nor U37403 (N_37403,N_33149,N_30575);
or U37404 (N_37404,N_30322,N_31926);
or U37405 (N_37405,N_34704,N_33729);
or U37406 (N_37406,N_34765,N_34893);
nand U37407 (N_37407,N_33974,N_31762);
nand U37408 (N_37408,N_33631,N_33491);
or U37409 (N_37409,N_34625,N_34522);
or U37410 (N_37410,N_33639,N_32656);
nor U37411 (N_37411,N_30367,N_31125);
nor U37412 (N_37412,N_31516,N_31494);
nor U37413 (N_37413,N_33176,N_31576);
or U37414 (N_37414,N_34679,N_31523);
and U37415 (N_37415,N_30145,N_32332);
and U37416 (N_37416,N_31910,N_32146);
nor U37417 (N_37417,N_31501,N_32825);
nand U37418 (N_37418,N_31502,N_33141);
and U37419 (N_37419,N_34074,N_33841);
nand U37420 (N_37420,N_30400,N_30647);
and U37421 (N_37421,N_30178,N_33839);
xor U37422 (N_37422,N_34675,N_34317);
and U37423 (N_37423,N_33958,N_32351);
and U37424 (N_37424,N_30782,N_32311);
or U37425 (N_37425,N_31394,N_31066);
or U37426 (N_37426,N_32323,N_31172);
nand U37427 (N_37427,N_30930,N_33756);
or U37428 (N_37428,N_33189,N_34393);
nor U37429 (N_37429,N_32201,N_33192);
nor U37430 (N_37430,N_30609,N_33682);
nor U37431 (N_37431,N_31968,N_31836);
nand U37432 (N_37432,N_30165,N_34875);
nor U37433 (N_37433,N_33741,N_31918);
or U37434 (N_37434,N_33129,N_32310);
nand U37435 (N_37435,N_32325,N_33289);
xnor U37436 (N_37436,N_30115,N_33513);
and U37437 (N_37437,N_32851,N_31396);
and U37438 (N_37438,N_31941,N_33876);
nor U37439 (N_37439,N_32189,N_31842);
nand U37440 (N_37440,N_30249,N_32464);
and U37441 (N_37441,N_33785,N_30010);
nor U37442 (N_37442,N_34453,N_33266);
nor U37443 (N_37443,N_32753,N_34138);
nor U37444 (N_37444,N_30244,N_30577);
nand U37445 (N_37445,N_34439,N_30250);
or U37446 (N_37446,N_34347,N_34239);
and U37447 (N_37447,N_33962,N_32555);
or U37448 (N_37448,N_33763,N_32672);
and U37449 (N_37449,N_33783,N_33006);
nand U37450 (N_37450,N_32036,N_32967);
or U37451 (N_37451,N_32527,N_31495);
nor U37452 (N_37452,N_32674,N_30233);
xnor U37453 (N_37453,N_30519,N_34181);
xor U37454 (N_37454,N_31036,N_32682);
nor U37455 (N_37455,N_30177,N_31937);
nand U37456 (N_37456,N_33564,N_33210);
and U37457 (N_37457,N_32401,N_30259);
and U37458 (N_37458,N_31094,N_32411);
nand U37459 (N_37459,N_34785,N_31882);
nor U37460 (N_37460,N_30431,N_32662);
and U37461 (N_37461,N_33108,N_32253);
nor U37462 (N_37462,N_32127,N_34171);
nor U37463 (N_37463,N_34351,N_32365);
nor U37464 (N_37464,N_31222,N_31512);
or U37465 (N_37465,N_32621,N_32017);
xor U37466 (N_37466,N_33833,N_33943);
xor U37467 (N_37467,N_33103,N_30628);
nand U37468 (N_37468,N_31507,N_34105);
nand U37469 (N_37469,N_31729,N_32933);
or U37470 (N_37470,N_33110,N_32509);
nand U37471 (N_37471,N_30752,N_33828);
or U37472 (N_37472,N_34287,N_31898);
or U37473 (N_37473,N_32343,N_34536);
nor U37474 (N_37474,N_31171,N_31786);
nand U37475 (N_37475,N_30423,N_30554);
and U37476 (N_37476,N_31294,N_32597);
or U37477 (N_37477,N_30096,N_31465);
xor U37478 (N_37478,N_32952,N_31419);
and U37479 (N_37479,N_31570,N_30345);
xnor U37480 (N_37480,N_32074,N_30006);
nand U37481 (N_37481,N_32160,N_32950);
and U37482 (N_37482,N_33205,N_33369);
and U37483 (N_37483,N_32990,N_31472);
nand U37484 (N_37484,N_33621,N_34407);
nand U37485 (N_37485,N_31551,N_33260);
and U37486 (N_37486,N_30872,N_33997);
nand U37487 (N_37487,N_31531,N_30902);
nor U37488 (N_37488,N_33256,N_30827);
and U37489 (N_37489,N_34650,N_33408);
nand U37490 (N_37490,N_30210,N_34663);
and U37491 (N_37491,N_33734,N_31190);
or U37492 (N_37492,N_34779,N_32141);
nor U37493 (N_37493,N_32969,N_31051);
and U37494 (N_37494,N_32319,N_31949);
or U37495 (N_37495,N_31043,N_32958);
and U37496 (N_37496,N_30330,N_32465);
nor U37497 (N_37497,N_30664,N_32994);
nand U37498 (N_37498,N_31984,N_34205);
and U37499 (N_37499,N_31177,N_31896);
xnor U37500 (N_37500,N_33787,N_31979);
and U37501 (N_37501,N_33993,N_32105);
nor U37502 (N_37502,N_34391,N_31687);
nand U37503 (N_37503,N_34751,N_34664);
or U37504 (N_37504,N_30960,N_31274);
nand U37505 (N_37505,N_32841,N_34206);
xnor U37506 (N_37506,N_31888,N_31615);
nand U37507 (N_37507,N_30460,N_34256);
nor U37508 (N_37508,N_31968,N_34659);
or U37509 (N_37509,N_33884,N_33702);
or U37510 (N_37510,N_31282,N_33192);
xor U37511 (N_37511,N_30668,N_31141);
and U37512 (N_37512,N_34474,N_34756);
nor U37513 (N_37513,N_34869,N_34837);
nor U37514 (N_37514,N_32497,N_30772);
nor U37515 (N_37515,N_31686,N_34498);
xnor U37516 (N_37516,N_33977,N_30543);
or U37517 (N_37517,N_33517,N_30506);
nor U37518 (N_37518,N_33381,N_31363);
and U37519 (N_37519,N_33629,N_30061);
and U37520 (N_37520,N_33552,N_33239);
and U37521 (N_37521,N_34690,N_30832);
or U37522 (N_37522,N_32852,N_33491);
and U37523 (N_37523,N_30615,N_31824);
or U37524 (N_37524,N_34173,N_33477);
nand U37525 (N_37525,N_34930,N_33566);
nand U37526 (N_37526,N_32818,N_34533);
nand U37527 (N_37527,N_30515,N_32060);
nor U37528 (N_37528,N_31636,N_34944);
or U37529 (N_37529,N_31686,N_32009);
nor U37530 (N_37530,N_34539,N_30252);
nand U37531 (N_37531,N_34130,N_32567);
or U37532 (N_37532,N_34344,N_30017);
nand U37533 (N_37533,N_30305,N_33124);
and U37534 (N_37534,N_32227,N_31100);
nor U37535 (N_37535,N_32822,N_34751);
and U37536 (N_37536,N_34564,N_31268);
nand U37537 (N_37537,N_32971,N_32883);
nand U37538 (N_37538,N_33464,N_32791);
nand U37539 (N_37539,N_30393,N_31308);
and U37540 (N_37540,N_32298,N_31641);
nor U37541 (N_37541,N_33236,N_31196);
and U37542 (N_37542,N_30683,N_32766);
xnor U37543 (N_37543,N_32757,N_33203);
nor U37544 (N_37544,N_31754,N_34806);
nand U37545 (N_37545,N_32335,N_32638);
xor U37546 (N_37546,N_31106,N_34643);
or U37547 (N_37547,N_31368,N_33021);
nand U37548 (N_37548,N_34330,N_32739);
nand U37549 (N_37549,N_31891,N_34379);
xor U37550 (N_37550,N_32862,N_33670);
and U37551 (N_37551,N_30052,N_31402);
or U37552 (N_37552,N_32240,N_32981);
or U37553 (N_37553,N_32617,N_33776);
nand U37554 (N_37554,N_34941,N_33195);
nor U37555 (N_37555,N_33956,N_34074);
xor U37556 (N_37556,N_31252,N_34127);
nand U37557 (N_37557,N_34181,N_32800);
nand U37558 (N_37558,N_32315,N_32329);
xor U37559 (N_37559,N_33635,N_33907);
and U37560 (N_37560,N_34256,N_34063);
xor U37561 (N_37561,N_30873,N_33124);
nand U37562 (N_37562,N_33836,N_33663);
and U37563 (N_37563,N_34371,N_32543);
nor U37564 (N_37564,N_34216,N_32779);
nor U37565 (N_37565,N_32719,N_31176);
and U37566 (N_37566,N_34673,N_32133);
and U37567 (N_37567,N_32891,N_31592);
or U37568 (N_37568,N_31315,N_30322);
nor U37569 (N_37569,N_32820,N_31149);
and U37570 (N_37570,N_31576,N_34261);
nand U37571 (N_37571,N_34069,N_32368);
nor U37572 (N_37572,N_33898,N_30205);
or U37573 (N_37573,N_30521,N_32370);
nand U37574 (N_37574,N_31840,N_32804);
nor U37575 (N_37575,N_32120,N_32575);
or U37576 (N_37576,N_32988,N_31148);
xor U37577 (N_37577,N_31389,N_34680);
xnor U37578 (N_37578,N_32280,N_31231);
and U37579 (N_37579,N_33040,N_30717);
or U37580 (N_37580,N_33490,N_34282);
or U37581 (N_37581,N_33222,N_32871);
nand U37582 (N_37582,N_31298,N_34250);
nand U37583 (N_37583,N_31705,N_34762);
or U37584 (N_37584,N_30324,N_34177);
or U37585 (N_37585,N_31954,N_33327);
and U37586 (N_37586,N_31876,N_30809);
nor U37587 (N_37587,N_34189,N_32561);
or U37588 (N_37588,N_32325,N_33907);
xor U37589 (N_37589,N_30798,N_31880);
nand U37590 (N_37590,N_32258,N_30329);
nand U37591 (N_37591,N_34673,N_30686);
and U37592 (N_37592,N_31806,N_34721);
or U37593 (N_37593,N_32397,N_34683);
nor U37594 (N_37594,N_32281,N_32292);
nand U37595 (N_37595,N_34458,N_34522);
xor U37596 (N_37596,N_30578,N_31747);
nor U37597 (N_37597,N_30738,N_34232);
and U37598 (N_37598,N_34401,N_33372);
or U37599 (N_37599,N_33013,N_33238);
nand U37600 (N_37600,N_34434,N_31917);
nand U37601 (N_37601,N_31257,N_34903);
nand U37602 (N_37602,N_33243,N_30992);
nand U37603 (N_37603,N_33038,N_33655);
nand U37604 (N_37604,N_32587,N_34796);
nor U37605 (N_37605,N_31122,N_32650);
nand U37606 (N_37606,N_33822,N_32658);
nor U37607 (N_37607,N_30543,N_30678);
nand U37608 (N_37608,N_34845,N_31919);
nor U37609 (N_37609,N_32355,N_33637);
and U37610 (N_37610,N_33912,N_32011);
nand U37611 (N_37611,N_33806,N_33238);
or U37612 (N_37612,N_30044,N_32781);
and U37613 (N_37613,N_34170,N_32071);
or U37614 (N_37614,N_32720,N_31132);
nor U37615 (N_37615,N_32692,N_34979);
xnor U37616 (N_37616,N_30011,N_31894);
nor U37617 (N_37617,N_34489,N_34409);
or U37618 (N_37618,N_32300,N_34575);
nand U37619 (N_37619,N_30692,N_30139);
or U37620 (N_37620,N_33331,N_33978);
xnor U37621 (N_37621,N_32040,N_33741);
nor U37622 (N_37622,N_30664,N_30969);
and U37623 (N_37623,N_34739,N_34690);
and U37624 (N_37624,N_33115,N_30439);
nand U37625 (N_37625,N_33022,N_32555);
nor U37626 (N_37626,N_34539,N_31671);
xnor U37627 (N_37627,N_31334,N_33468);
nand U37628 (N_37628,N_34687,N_33271);
and U37629 (N_37629,N_32518,N_30965);
nor U37630 (N_37630,N_32060,N_31744);
nand U37631 (N_37631,N_32490,N_32057);
and U37632 (N_37632,N_34773,N_32846);
nor U37633 (N_37633,N_30874,N_31724);
or U37634 (N_37634,N_34973,N_33826);
nand U37635 (N_37635,N_32677,N_32678);
or U37636 (N_37636,N_31831,N_30182);
xor U37637 (N_37637,N_30890,N_30246);
and U37638 (N_37638,N_33229,N_32982);
nand U37639 (N_37639,N_31801,N_34036);
or U37640 (N_37640,N_30171,N_32588);
and U37641 (N_37641,N_32032,N_33364);
nor U37642 (N_37642,N_30442,N_32537);
nand U37643 (N_37643,N_34003,N_31137);
or U37644 (N_37644,N_34953,N_31467);
nand U37645 (N_37645,N_31573,N_30297);
or U37646 (N_37646,N_34101,N_31794);
nand U37647 (N_37647,N_32323,N_30696);
nand U37648 (N_37648,N_33667,N_34395);
and U37649 (N_37649,N_31273,N_32536);
or U37650 (N_37650,N_32706,N_31008);
and U37651 (N_37651,N_30515,N_30416);
or U37652 (N_37652,N_34754,N_34282);
xnor U37653 (N_37653,N_30122,N_32470);
or U37654 (N_37654,N_33397,N_32440);
nor U37655 (N_37655,N_31326,N_33806);
or U37656 (N_37656,N_31772,N_34547);
or U37657 (N_37657,N_34718,N_34842);
xor U37658 (N_37658,N_31363,N_34342);
nand U37659 (N_37659,N_33979,N_32788);
nand U37660 (N_37660,N_34740,N_33074);
or U37661 (N_37661,N_30364,N_34418);
and U37662 (N_37662,N_30157,N_33276);
and U37663 (N_37663,N_32059,N_33276);
and U37664 (N_37664,N_30877,N_34567);
nor U37665 (N_37665,N_30096,N_31725);
xor U37666 (N_37666,N_30147,N_33302);
and U37667 (N_37667,N_31306,N_33378);
xor U37668 (N_37668,N_31267,N_31618);
and U37669 (N_37669,N_31080,N_33458);
and U37670 (N_37670,N_32605,N_31085);
nand U37671 (N_37671,N_31102,N_33478);
and U37672 (N_37672,N_30969,N_31909);
or U37673 (N_37673,N_32883,N_32203);
nor U37674 (N_37674,N_33392,N_33501);
nand U37675 (N_37675,N_33523,N_32033);
nor U37676 (N_37676,N_34588,N_33184);
or U37677 (N_37677,N_32474,N_33188);
nand U37678 (N_37678,N_34488,N_32002);
and U37679 (N_37679,N_32682,N_33640);
and U37680 (N_37680,N_31817,N_30051);
nand U37681 (N_37681,N_33404,N_34150);
nor U37682 (N_37682,N_31652,N_32121);
nand U37683 (N_37683,N_30428,N_30679);
nor U37684 (N_37684,N_31581,N_30612);
or U37685 (N_37685,N_31588,N_30557);
nor U37686 (N_37686,N_33719,N_34234);
and U37687 (N_37687,N_32506,N_30439);
or U37688 (N_37688,N_30485,N_33690);
and U37689 (N_37689,N_33427,N_32091);
or U37690 (N_37690,N_30884,N_32546);
or U37691 (N_37691,N_32592,N_31899);
xnor U37692 (N_37692,N_33967,N_32739);
nand U37693 (N_37693,N_32713,N_32218);
or U37694 (N_37694,N_33003,N_33691);
nor U37695 (N_37695,N_30518,N_34979);
xnor U37696 (N_37696,N_33277,N_32943);
nor U37697 (N_37697,N_30992,N_30367);
and U37698 (N_37698,N_33606,N_33556);
and U37699 (N_37699,N_32636,N_30730);
or U37700 (N_37700,N_30259,N_33589);
xnor U37701 (N_37701,N_32172,N_33499);
and U37702 (N_37702,N_30879,N_32397);
nand U37703 (N_37703,N_31870,N_30869);
and U37704 (N_37704,N_32353,N_31432);
nand U37705 (N_37705,N_30814,N_32221);
nand U37706 (N_37706,N_31940,N_33847);
or U37707 (N_37707,N_32201,N_34856);
nand U37708 (N_37708,N_34510,N_33784);
and U37709 (N_37709,N_30948,N_30014);
xor U37710 (N_37710,N_31606,N_30080);
or U37711 (N_37711,N_30354,N_30268);
or U37712 (N_37712,N_34181,N_31928);
nor U37713 (N_37713,N_31783,N_31642);
nor U37714 (N_37714,N_32269,N_31531);
and U37715 (N_37715,N_30397,N_30090);
nand U37716 (N_37716,N_32772,N_34194);
nor U37717 (N_37717,N_32763,N_30924);
nand U37718 (N_37718,N_30257,N_32783);
and U37719 (N_37719,N_30555,N_34852);
nand U37720 (N_37720,N_33633,N_30155);
xor U37721 (N_37721,N_32476,N_30702);
and U37722 (N_37722,N_33988,N_30011);
and U37723 (N_37723,N_31133,N_31177);
nor U37724 (N_37724,N_33280,N_31693);
or U37725 (N_37725,N_34179,N_30006);
nand U37726 (N_37726,N_32416,N_33298);
nor U37727 (N_37727,N_32331,N_33535);
nor U37728 (N_37728,N_33725,N_30497);
nand U37729 (N_37729,N_34672,N_30050);
nor U37730 (N_37730,N_31188,N_30233);
nor U37731 (N_37731,N_34782,N_32951);
or U37732 (N_37732,N_34399,N_30800);
nand U37733 (N_37733,N_34163,N_33740);
and U37734 (N_37734,N_31138,N_31417);
or U37735 (N_37735,N_34581,N_34752);
or U37736 (N_37736,N_30525,N_32690);
nand U37737 (N_37737,N_32459,N_30124);
and U37738 (N_37738,N_33786,N_32496);
or U37739 (N_37739,N_32055,N_31689);
nor U37740 (N_37740,N_33726,N_32249);
or U37741 (N_37741,N_33321,N_30429);
and U37742 (N_37742,N_32304,N_34946);
nor U37743 (N_37743,N_30357,N_33725);
nor U37744 (N_37744,N_34177,N_34197);
nand U37745 (N_37745,N_34298,N_33651);
or U37746 (N_37746,N_32667,N_33383);
nand U37747 (N_37747,N_34968,N_33569);
and U37748 (N_37748,N_33177,N_32957);
xor U37749 (N_37749,N_32499,N_30404);
and U37750 (N_37750,N_31188,N_33947);
nand U37751 (N_37751,N_33297,N_31004);
xor U37752 (N_37752,N_31877,N_33338);
nor U37753 (N_37753,N_31034,N_30218);
nand U37754 (N_37754,N_30121,N_31313);
nor U37755 (N_37755,N_34389,N_34871);
or U37756 (N_37756,N_33009,N_31408);
or U37757 (N_37757,N_33369,N_32621);
and U37758 (N_37758,N_31906,N_31764);
and U37759 (N_37759,N_32195,N_32501);
and U37760 (N_37760,N_30490,N_32737);
nand U37761 (N_37761,N_34977,N_31014);
nand U37762 (N_37762,N_33256,N_33855);
and U37763 (N_37763,N_33453,N_32089);
nand U37764 (N_37764,N_33668,N_31652);
or U37765 (N_37765,N_30420,N_33677);
and U37766 (N_37766,N_32763,N_31347);
or U37767 (N_37767,N_33362,N_32555);
xnor U37768 (N_37768,N_33547,N_31453);
nor U37769 (N_37769,N_31242,N_34057);
or U37770 (N_37770,N_30635,N_30412);
xor U37771 (N_37771,N_30104,N_32915);
and U37772 (N_37772,N_30815,N_31971);
nand U37773 (N_37773,N_30925,N_31489);
nor U37774 (N_37774,N_34791,N_34913);
and U37775 (N_37775,N_34174,N_30622);
nor U37776 (N_37776,N_31830,N_33936);
and U37777 (N_37777,N_34000,N_31338);
nand U37778 (N_37778,N_33709,N_30769);
nand U37779 (N_37779,N_33951,N_31668);
or U37780 (N_37780,N_30296,N_31633);
or U37781 (N_37781,N_31051,N_31332);
and U37782 (N_37782,N_31916,N_32407);
nor U37783 (N_37783,N_31668,N_34691);
nand U37784 (N_37784,N_32844,N_32930);
xor U37785 (N_37785,N_31929,N_31532);
nor U37786 (N_37786,N_34872,N_34521);
nand U37787 (N_37787,N_31698,N_30233);
or U37788 (N_37788,N_30583,N_30459);
nor U37789 (N_37789,N_30536,N_34275);
nor U37790 (N_37790,N_31760,N_34011);
nand U37791 (N_37791,N_31494,N_33714);
and U37792 (N_37792,N_31418,N_31607);
nor U37793 (N_37793,N_30803,N_31927);
nor U37794 (N_37794,N_33210,N_30454);
nand U37795 (N_37795,N_32035,N_30667);
nor U37796 (N_37796,N_32825,N_30581);
or U37797 (N_37797,N_33683,N_31878);
or U37798 (N_37798,N_32016,N_30289);
nand U37799 (N_37799,N_33853,N_34049);
nand U37800 (N_37800,N_30599,N_34091);
nand U37801 (N_37801,N_32339,N_34942);
xnor U37802 (N_37802,N_33387,N_34993);
nor U37803 (N_37803,N_31236,N_34322);
or U37804 (N_37804,N_30471,N_31961);
nand U37805 (N_37805,N_32580,N_33180);
nor U37806 (N_37806,N_33171,N_32658);
nand U37807 (N_37807,N_31879,N_30609);
or U37808 (N_37808,N_31719,N_32751);
nand U37809 (N_37809,N_30859,N_34927);
or U37810 (N_37810,N_31740,N_34916);
or U37811 (N_37811,N_30017,N_33076);
xnor U37812 (N_37812,N_31151,N_30290);
and U37813 (N_37813,N_33367,N_32954);
and U37814 (N_37814,N_34249,N_30190);
nor U37815 (N_37815,N_31487,N_34200);
xnor U37816 (N_37816,N_31136,N_32996);
xor U37817 (N_37817,N_33034,N_32399);
nor U37818 (N_37818,N_31751,N_30301);
or U37819 (N_37819,N_33104,N_33424);
and U37820 (N_37820,N_34404,N_33471);
nor U37821 (N_37821,N_32462,N_30633);
and U37822 (N_37822,N_33500,N_33885);
or U37823 (N_37823,N_30621,N_30401);
and U37824 (N_37824,N_32630,N_33975);
nor U37825 (N_37825,N_30609,N_32640);
and U37826 (N_37826,N_31220,N_33408);
nand U37827 (N_37827,N_30252,N_34983);
nor U37828 (N_37828,N_34011,N_33084);
and U37829 (N_37829,N_33230,N_32547);
and U37830 (N_37830,N_32725,N_33648);
or U37831 (N_37831,N_31643,N_31216);
nor U37832 (N_37832,N_33683,N_32750);
or U37833 (N_37833,N_32691,N_34120);
nand U37834 (N_37834,N_33206,N_32306);
nand U37835 (N_37835,N_33987,N_30388);
and U37836 (N_37836,N_34453,N_31141);
or U37837 (N_37837,N_34407,N_32506);
nor U37838 (N_37838,N_32264,N_30605);
nand U37839 (N_37839,N_34742,N_32348);
and U37840 (N_37840,N_34281,N_31270);
nor U37841 (N_37841,N_32615,N_33040);
or U37842 (N_37842,N_31527,N_31136);
or U37843 (N_37843,N_32481,N_33989);
or U37844 (N_37844,N_32595,N_32299);
or U37845 (N_37845,N_31075,N_32551);
nor U37846 (N_37846,N_34620,N_32559);
and U37847 (N_37847,N_30359,N_33058);
or U37848 (N_37848,N_30766,N_30124);
or U37849 (N_37849,N_30874,N_34072);
xor U37850 (N_37850,N_30537,N_34903);
or U37851 (N_37851,N_31716,N_33147);
and U37852 (N_37852,N_34902,N_33094);
xor U37853 (N_37853,N_31546,N_31402);
nand U37854 (N_37854,N_33213,N_33133);
or U37855 (N_37855,N_34510,N_33979);
and U37856 (N_37856,N_30599,N_30298);
nand U37857 (N_37857,N_33903,N_31616);
nand U37858 (N_37858,N_31426,N_33395);
nor U37859 (N_37859,N_33186,N_33722);
nand U37860 (N_37860,N_34145,N_31400);
xnor U37861 (N_37861,N_31835,N_32627);
or U37862 (N_37862,N_33869,N_32327);
xor U37863 (N_37863,N_34408,N_32154);
nand U37864 (N_37864,N_31551,N_32801);
nor U37865 (N_37865,N_31018,N_32993);
nor U37866 (N_37866,N_31840,N_34868);
xor U37867 (N_37867,N_30665,N_31363);
or U37868 (N_37868,N_32222,N_34134);
or U37869 (N_37869,N_32337,N_33364);
nand U37870 (N_37870,N_33816,N_33104);
or U37871 (N_37871,N_31065,N_30990);
nand U37872 (N_37872,N_33912,N_33478);
nand U37873 (N_37873,N_32470,N_34950);
or U37874 (N_37874,N_33489,N_31417);
nand U37875 (N_37875,N_33495,N_32597);
or U37876 (N_37876,N_33533,N_30075);
and U37877 (N_37877,N_30516,N_32856);
or U37878 (N_37878,N_30487,N_33336);
or U37879 (N_37879,N_34355,N_34811);
nor U37880 (N_37880,N_32387,N_31819);
nand U37881 (N_37881,N_30158,N_30693);
or U37882 (N_37882,N_33272,N_32391);
and U37883 (N_37883,N_31093,N_32044);
and U37884 (N_37884,N_32880,N_30718);
nor U37885 (N_37885,N_31925,N_33754);
or U37886 (N_37886,N_31741,N_34431);
or U37887 (N_37887,N_32595,N_31816);
nand U37888 (N_37888,N_34830,N_30474);
xor U37889 (N_37889,N_31080,N_31017);
xor U37890 (N_37890,N_31740,N_30006);
or U37891 (N_37891,N_30295,N_34015);
xor U37892 (N_37892,N_34920,N_31749);
nor U37893 (N_37893,N_32562,N_34013);
or U37894 (N_37894,N_31816,N_34627);
or U37895 (N_37895,N_31337,N_31152);
or U37896 (N_37896,N_34479,N_32382);
or U37897 (N_37897,N_31365,N_32614);
and U37898 (N_37898,N_30091,N_33262);
or U37899 (N_37899,N_34465,N_32968);
nand U37900 (N_37900,N_34176,N_32928);
or U37901 (N_37901,N_33754,N_31890);
or U37902 (N_37902,N_34834,N_33757);
or U37903 (N_37903,N_31867,N_34489);
or U37904 (N_37904,N_30294,N_32433);
nor U37905 (N_37905,N_30513,N_32610);
or U37906 (N_37906,N_33379,N_34111);
and U37907 (N_37907,N_30985,N_30257);
and U37908 (N_37908,N_30390,N_34757);
or U37909 (N_37909,N_31621,N_31558);
or U37910 (N_37910,N_31761,N_32608);
or U37911 (N_37911,N_31073,N_32424);
nand U37912 (N_37912,N_30167,N_33342);
and U37913 (N_37913,N_34522,N_30645);
xor U37914 (N_37914,N_33190,N_31284);
or U37915 (N_37915,N_34100,N_30626);
nand U37916 (N_37916,N_30903,N_32350);
xor U37917 (N_37917,N_33563,N_32371);
or U37918 (N_37918,N_30786,N_33690);
and U37919 (N_37919,N_33073,N_32318);
and U37920 (N_37920,N_33616,N_30452);
nor U37921 (N_37921,N_32050,N_30411);
nand U37922 (N_37922,N_30057,N_34675);
nand U37923 (N_37923,N_31880,N_34449);
nor U37924 (N_37924,N_31493,N_32724);
nor U37925 (N_37925,N_30924,N_31840);
nand U37926 (N_37926,N_32477,N_34835);
nor U37927 (N_37927,N_33822,N_34841);
and U37928 (N_37928,N_31168,N_32024);
and U37929 (N_37929,N_32370,N_33152);
xnor U37930 (N_37930,N_30555,N_34316);
nor U37931 (N_37931,N_34505,N_33364);
nand U37932 (N_37932,N_31299,N_32862);
nor U37933 (N_37933,N_34634,N_34502);
nor U37934 (N_37934,N_31554,N_32766);
or U37935 (N_37935,N_30029,N_33559);
nor U37936 (N_37936,N_33670,N_34090);
or U37937 (N_37937,N_30991,N_32576);
nand U37938 (N_37938,N_34272,N_32195);
nor U37939 (N_37939,N_33709,N_30193);
and U37940 (N_37940,N_31730,N_34692);
nand U37941 (N_37941,N_30218,N_33264);
nor U37942 (N_37942,N_31387,N_32591);
nand U37943 (N_37943,N_30771,N_34243);
nand U37944 (N_37944,N_34898,N_34260);
nand U37945 (N_37945,N_33648,N_31807);
or U37946 (N_37946,N_30827,N_31989);
and U37947 (N_37947,N_34871,N_31682);
nand U37948 (N_37948,N_31839,N_31798);
and U37949 (N_37949,N_31181,N_32492);
nand U37950 (N_37950,N_30536,N_33287);
and U37951 (N_37951,N_31290,N_31894);
xor U37952 (N_37952,N_34482,N_32606);
and U37953 (N_37953,N_32466,N_32654);
nand U37954 (N_37954,N_33076,N_30302);
nand U37955 (N_37955,N_32442,N_31104);
xnor U37956 (N_37956,N_33342,N_34765);
and U37957 (N_37957,N_31065,N_32464);
or U37958 (N_37958,N_34476,N_32084);
nor U37959 (N_37959,N_30274,N_32649);
nor U37960 (N_37960,N_30152,N_31040);
nand U37961 (N_37961,N_32222,N_32370);
or U37962 (N_37962,N_32378,N_33829);
nor U37963 (N_37963,N_32879,N_31772);
nand U37964 (N_37964,N_32037,N_34739);
nor U37965 (N_37965,N_33356,N_32972);
or U37966 (N_37966,N_31833,N_34019);
nor U37967 (N_37967,N_34914,N_31605);
nand U37968 (N_37968,N_30750,N_33009);
nor U37969 (N_37969,N_34577,N_34345);
nor U37970 (N_37970,N_31848,N_32793);
nor U37971 (N_37971,N_33904,N_34911);
nand U37972 (N_37972,N_30524,N_32229);
nor U37973 (N_37973,N_34727,N_34625);
or U37974 (N_37974,N_31213,N_32618);
and U37975 (N_37975,N_31956,N_30759);
nand U37976 (N_37976,N_33398,N_30486);
nand U37977 (N_37977,N_30172,N_34871);
nand U37978 (N_37978,N_33033,N_31880);
nand U37979 (N_37979,N_33591,N_31983);
nor U37980 (N_37980,N_30355,N_34781);
and U37981 (N_37981,N_34574,N_31857);
nor U37982 (N_37982,N_30959,N_30000);
or U37983 (N_37983,N_30534,N_30847);
or U37984 (N_37984,N_34472,N_32872);
nand U37985 (N_37985,N_32118,N_34151);
nand U37986 (N_37986,N_34908,N_30228);
and U37987 (N_37987,N_32139,N_33921);
nor U37988 (N_37988,N_31290,N_31641);
and U37989 (N_37989,N_34797,N_32769);
or U37990 (N_37990,N_32514,N_30404);
nand U37991 (N_37991,N_30845,N_34948);
nor U37992 (N_37992,N_32497,N_30426);
and U37993 (N_37993,N_31376,N_34581);
and U37994 (N_37994,N_30519,N_30537);
nor U37995 (N_37995,N_31572,N_31373);
and U37996 (N_37996,N_32320,N_31778);
or U37997 (N_37997,N_32340,N_31082);
and U37998 (N_37998,N_31358,N_30249);
and U37999 (N_37999,N_32638,N_34668);
and U38000 (N_38000,N_34460,N_32082);
nand U38001 (N_38001,N_31461,N_33264);
or U38002 (N_38002,N_31373,N_30744);
nand U38003 (N_38003,N_34645,N_34061);
xnor U38004 (N_38004,N_30975,N_34764);
nand U38005 (N_38005,N_32526,N_30795);
nand U38006 (N_38006,N_31373,N_30840);
and U38007 (N_38007,N_32199,N_32659);
nor U38008 (N_38008,N_31908,N_33926);
xnor U38009 (N_38009,N_34795,N_34538);
nand U38010 (N_38010,N_30408,N_30851);
or U38011 (N_38011,N_32895,N_31789);
or U38012 (N_38012,N_34873,N_33418);
nand U38013 (N_38013,N_30831,N_30842);
nand U38014 (N_38014,N_34842,N_33229);
and U38015 (N_38015,N_30956,N_34538);
or U38016 (N_38016,N_30463,N_31741);
nor U38017 (N_38017,N_34148,N_33873);
nor U38018 (N_38018,N_30800,N_34768);
and U38019 (N_38019,N_30288,N_30368);
nand U38020 (N_38020,N_32007,N_31275);
nor U38021 (N_38021,N_32854,N_31730);
nor U38022 (N_38022,N_30880,N_33388);
nand U38023 (N_38023,N_33649,N_32499);
or U38024 (N_38024,N_32204,N_32191);
and U38025 (N_38025,N_34478,N_30521);
and U38026 (N_38026,N_30692,N_32375);
nor U38027 (N_38027,N_33354,N_30341);
nand U38028 (N_38028,N_33981,N_33568);
nor U38029 (N_38029,N_31735,N_33845);
and U38030 (N_38030,N_32336,N_30178);
nor U38031 (N_38031,N_32307,N_30503);
and U38032 (N_38032,N_33889,N_34326);
and U38033 (N_38033,N_31048,N_34009);
and U38034 (N_38034,N_34300,N_30904);
and U38035 (N_38035,N_31030,N_30307);
or U38036 (N_38036,N_30845,N_32136);
nand U38037 (N_38037,N_30994,N_30978);
nand U38038 (N_38038,N_33966,N_32781);
and U38039 (N_38039,N_33645,N_31152);
nand U38040 (N_38040,N_30001,N_31353);
nand U38041 (N_38041,N_33358,N_31893);
nand U38042 (N_38042,N_31217,N_31281);
nand U38043 (N_38043,N_30863,N_31376);
nor U38044 (N_38044,N_32504,N_30691);
xnor U38045 (N_38045,N_32148,N_34093);
nor U38046 (N_38046,N_31752,N_32324);
nand U38047 (N_38047,N_31760,N_33722);
or U38048 (N_38048,N_32262,N_34258);
nor U38049 (N_38049,N_31792,N_31342);
and U38050 (N_38050,N_32878,N_33289);
and U38051 (N_38051,N_30751,N_31692);
nand U38052 (N_38052,N_34711,N_34304);
nand U38053 (N_38053,N_32378,N_31827);
or U38054 (N_38054,N_30736,N_30905);
and U38055 (N_38055,N_30025,N_34911);
nor U38056 (N_38056,N_32628,N_34837);
and U38057 (N_38057,N_32672,N_33049);
and U38058 (N_38058,N_32300,N_32404);
or U38059 (N_38059,N_30216,N_34437);
nand U38060 (N_38060,N_30402,N_32431);
and U38061 (N_38061,N_31389,N_33353);
nor U38062 (N_38062,N_34727,N_34035);
nand U38063 (N_38063,N_31673,N_34176);
nor U38064 (N_38064,N_32387,N_32053);
xnor U38065 (N_38065,N_33521,N_30301);
or U38066 (N_38066,N_31035,N_33947);
nor U38067 (N_38067,N_32536,N_31363);
nand U38068 (N_38068,N_34640,N_34232);
nand U38069 (N_38069,N_33906,N_32477);
xnor U38070 (N_38070,N_32914,N_34274);
and U38071 (N_38071,N_33576,N_32274);
and U38072 (N_38072,N_34175,N_34855);
and U38073 (N_38073,N_30813,N_33177);
nand U38074 (N_38074,N_33051,N_31649);
nor U38075 (N_38075,N_32986,N_30335);
or U38076 (N_38076,N_32574,N_30666);
and U38077 (N_38077,N_32272,N_34617);
xor U38078 (N_38078,N_32377,N_31272);
xnor U38079 (N_38079,N_30991,N_32328);
or U38080 (N_38080,N_33713,N_34111);
xnor U38081 (N_38081,N_30127,N_34221);
and U38082 (N_38082,N_32045,N_30340);
and U38083 (N_38083,N_30553,N_30408);
nand U38084 (N_38084,N_32834,N_32989);
or U38085 (N_38085,N_31136,N_32368);
or U38086 (N_38086,N_31078,N_33292);
nor U38087 (N_38087,N_33761,N_34773);
nor U38088 (N_38088,N_34533,N_34528);
nand U38089 (N_38089,N_31157,N_32580);
nand U38090 (N_38090,N_32784,N_32720);
and U38091 (N_38091,N_32343,N_32196);
or U38092 (N_38092,N_34177,N_32289);
nor U38093 (N_38093,N_30470,N_33466);
and U38094 (N_38094,N_30611,N_33447);
and U38095 (N_38095,N_32796,N_30804);
nand U38096 (N_38096,N_32384,N_34183);
and U38097 (N_38097,N_32056,N_34166);
nor U38098 (N_38098,N_33613,N_31219);
nand U38099 (N_38099,N_30493,N_32837);
nor U38100 (N_38100,N_30063,N_31266);
xnor U38101 (N_38101,N_30887,N_30818);
and U38102 (N_38102,N_34763,N_33882);
or U38103 (N_38103,N_33747,N_30083);
or U38104 (N_38104,N_30980,N_33814);
xnor U38105 (N_38105,N_34481,N_33541);
and U38106 (N_38106,N_32031,N_34800);
and U38107 (N_38107,N_30163,N_31985);
and U38108 (N_38108,N_31469,N_30883);
or U38109 (N_38109,N_31249,N_34217);
xnor U38110 (N_38110,N_34990,N_31759);
nor U38111 (N_38111,N_30814,N_33613);
nand U38112 (N_38112,N_30837,N_31535);
nor U38113 (N_38113,N_33211,N_31834);
xor U38114 (N_38114,N_33145,N_34959);
nand U38115 (N_38115,N_32545,N_31708);
xor U38116 (N_38116,N_30260,N_34102);
or U38117 (N_38117,N_30053,N_33823);
nor U38118 (N_38118,N_30207,N_31613);
or U38119 (N_38119,N_31377,N_30635);
and U38120 (N_38120,N_32911,N_34407);
and U38121 (N_38121,N_31296,N_34403);
nor U38122 (N_38122,N_31549,N_30497);
and U38123 (N_38123,N_30536,N_34086);
and U38124 (N_38124,N_30208,N_30328);
or U38125 (N_38125,N_33543,N_31603);
and U38126 (N_38126,N_33553,N_32822);
nor U38127 (N_38127,N_31658,N_33390);
or U38128 (N_38128,N_34698,N_32464);
nor U38129 (N_38129,N_34230,N_34287);
or U38130 (N_38130,N_31056,N_34507);
and U38131 (N_38131,N_34583,N_33340);
nand U38132 (N_38132,N_32488,N_34788);
nand U38133 (N_38133,N_33965,N_31128);
or U38134 (N_38134,N_33254,N_31375);
or U38135 (N_38135,N_33821,N_34459);
or U38136 (N_38136,N_32460,N_34780);
or U38137 (N_38137,N_30007,N_31273);
or U38138 (N_38138,N_32824,N_33503);
xor U38139 (N_38139,N_32334,N_31801);
or U38140 (N_38140,N_32628,N_31555);
nand U38141 (N_38141,N_34498,N_33216);
nand U38142 (N_38142,N_34337,N_33547);
nand U38143 (N_38143,N_33338,N_34376);
or U38144 (N_38144,N_32201,N_34192);
nand U38145 (N_38145,N_33817,N_30867);
or U38146 (N_38146,N_32625,N_33538);
nand U38147 (N_38147,N_32498,N_30889);
and U38148 (N_38148,N_32318,N_33209);
and U38149 (N_38149,N_30963,N_34051);
or U38150 (N_38150,N_34589,N_32834);
xor U38151 (N_38151,N_33295,N_33452);
or U38152 (N_38152,N_30290,N_30474);
xnor U38153 (N_38153,N_31320,N_32231);
nor U38154 (N_38154,N_33970,N_30191);
or U38155 (N_38155,N_33624,N_30149);
nand U38156 (N_38156,N_30123,N_34534);
and U38157 (N_38157,N_30613,N_30022);
nand U38158 (N_38158,N_34677,N_34075);
nand U38159 (N_38159,N_34616,N_34964);
or U38160 (N_38160,N_31953,N_34136);
nor U38161 (N_38161,N_34463,N_33761);
nand U38162 (N_38162,N_32959,N_30557);
nor U38163 (N_38163,N_33297,N_30421);
nand U38164 (N_38164,N_30506,N_30123);
or U38165 (N_38165,N_31035,N_34473);
nor U38166 (N_38166,N_33098,N_31510);
and U38167 (N_38167,N_33281,N_31213);
and U38168 (N_38168,N_34891,N_34167);
nand U38169 (N_38169,N_31430,N_30086);
and U38170 (N_38170,N_33055,N_30786);
nand U38171 (N_38171,N_34054,N_34018);
xor U38172 (N_38172,N_30904,N_32601);
nor U38173 (N_38173,N_32855,N_33579);
nand U38174 (N_38174,N_33301,N_33048);
or U38175 (N_38175,N_31634,N_33026);
or U38176 (N_38176,N_32085,N_31526);
nand U38177 (N_38177,N_34241,N_31820);
nor U38178 (N_38178,N_34147,N_34617);
and U38179 (N_38179,N_30362,N_34350);
and U38180 (N_38180,N_31384,N_33048);
and U38181 (N_38181,N_31494,N_33595);
and U38182 (N_38182,N_32703,N_32874);
nand U38183 (N_38183,N_32161,N_33847);
nor U38184 (N_38184,N_34909,N_31312);
or U38185 (N_38185,N_34362,N_33548);
nand U38186 (N_38186,N_33668,N_32532);
and U38187 (N_38187,N_32978,N_33682);
and U38188 (N_38188,N_31736,N_31197);
nand U38189 (N_38189,N_30952,N_32449);
nor U38190 (N_38190,N_32320,N_34168);
nor U38191 (N_38191,N_31609,N_30267);
and U38192 (N_38192,N_33055,N_32394);
nand U38193 (N_38193,N_30657,N_34239);
or U38194 (N_38194,N_30549,N_31396);
or U38195 (N_38195,N_30991,N_30785);
or U38196 (N_38196,N_30972,N_32996);
nor U38197 (N_38197,N_30815,N_34035);
xnor U38198 (N_38198,N_30920,N_32348);
nor U38199 (N_38199,N_31719,N_33707);
nand U38200 (N_38200,N_34396,N_31396);
or U38201 (N_38201,N_33934,N_34586);
xor U38202 (N_38202,N_32548,N_31992);
and U38203 (N_38203,N_31988,N_31283);
nor U38204 (N_38204,N_34561,N_32948);
nor U38205 (N_38205,N_34466,N_33264);
or U38206 (N_38206,N_30124,N_34512);
nor U38207 (N_38207,N_31952,N_31837);
nand U38208 (N_38208,N_31771,N_30289);
nor U38209 (N_38209,N_32735,N_31922);
nor U38210 (N_38210,N_31956,N_31434);
or U38211 (N_38211,N_30393,N_34252);
and U38212 (N_38212,N_31899,N_34801);
nand U38213 (N_38213,N_31119,N_30535);
or U38214 (N_38214,N_30882,N_30712);
nor U38215 (N_38215,N_34751,N_34463);
nor U38216 (N_38216,N_33957,N_31490);
xnor U38217 (N_38217,N_34870,N_30838);
and U38218 (N_38218,N_33288,N_33668);
nand U38219 (N_38219,N_33751,N_30436);
xnor U38220 (N_38220,N_30002,N_30894);
nand U38221 (N_38221,N_33927,N_32423);
xnor U38222 (N_38222,N_34122,N_31548);
or U38223 (N_38223,N_31507,N_33025);
nor U38224 (N_38224,N_32075,N_30746);
or U38225 (N_38225,N_31124,N_30858);
nand U38226 (N_38226,N_34199,N_31290);
or U38227 (N_38227,N_33025,N_31140);
or U38228 (N_38228,N_32849,N_33909);
and U38229 (N_38229,N_32549,N_31344);
nand U38230 (N_38230,N_31715,N_31669);
and U38231 (N_38231,N_33913,N_31880);
or U38232 (N_38232,N_30577,N_32989);
nand U38233 (N_38233,N_31818,N_30763);
nand U38234 (N_38234,N_34263,N_32764);
nand U38235 (N_38235,N_30597,N_31973);
or U38236 (N_38236,N_33254,N_32425);
xor U38237 (N_38237,N_30557,N_31862);
and U38238 (N_38238,N_34428,N_34295);
nor U38239 (N_38239,N_30604,N_33240);
xnor U38240 (N_38240,N_30491,N_33667);
nor U38241 (N_38241,N_34556,N_32725);
nand U38242 (N_38242,N_33291,N_30157);
nand U38243 (N_38243,N_31958,N_34284);
and U38244 (N_38244,N_32021,N_34634);
nor U38245 (N_38245,N_34417,N_31921);
xor U38246 (N_38246,N_32583,N_33433);
nor U38247 (N_38247,N_31589,N_32814);
and U38248 (N_38248,N_34898,N_33871);
nand U38249 (N_38249,N_32717,N_30657);
xor U38250 (N_38250,N_33942,N_30616);
or U38251 (N_38251,N_31268,N_31229);
nor U38252 (N_38252,N_34315,N_34845);
or U38253 (N_38253,N_31446,N_32641);
xor U38254 (N_38254,N_31509,N_32265);
and U38255 (N_38255,N_32322,N_33849);
and U38256 (N_38256,N_34454,N_34611);
and U38257 (N_38257,N_32656,N_33285);
or U38258 (N_38258,N_34408,N_32404);
nand U38259 (N_38259,N_32968,N_34244);
xor U38260 (N_38260,N_31716,N_33186);
xor U38261 (N_38261,N_30265,N_32104);
xnor U38262 (N_38262,N_30327,N_34370);
nor U38263 (N_38263,N_31731,N_34925);
xor U38264 (N_38264,N_32112,N_34787);
or U38265 (N_38265,N_30048,N_30237);
or U38266 (N_38266,N_32149,N_30657);
nand U38267 (N_38267,N_30059,N_33484);
nor U38268 (N_38268,N_33779,N_31904);
xnor U38269 (N_38269,N_32410,N_33427);
nor U38270 (N_38270,N_33917,N_31123);
nor U38271 (N_38271,N_31427,N_33818);
nor U38272 (N_38272,N_32250,N_30850);
and U38273 (N_38273,N_32841,N_31226);
and U38274 (N_38274,N_30242,N_31658);
or U38275 (N_38275,N_32613,N_33997);
or U38276 (N_38276,N_32229,N_31115);
nand U38277 (N_38277,N_34191,N_34125);
and U38278 (N_38278,N_31960,N_34285);
and U38279 (N_38279,N_30480,N_30600);
and U38280 (N_38280,N_34173,N_30504);
or U38281 (N_38281,N_30067,N_32891);
and U38282 (N_38282,N_30161,N_33165);
or U38283 (N_38283,N_30480,N_31538);
nand U38284 (N_38284,N_32147,N_32723);
nand U38285 (N_38285,N_33773,N_32158);
nand U38286 (N_38286,N_32130,N_33814);
nor U38287 (N_38287,N_33220,N_30691);
xor U38288 (N_38288,N_34101,N_34358);
or U38289 (N_38289,N_34649,N_32034);
and U38290 (N_38290,N_30761,N_33395);
nor U38291 (N_38291,N_33514,N_32651);
xnor U38292 (N_38292,N_34121,N_34153);
nor U38293 (N_38293,N_34274,N_30042);
and U38294 (N_38294,N_33186,N_32342);
or U38295 (N_38295,N_34467,N_34765);
nor U38296 (N_38296,N_33016,N_34911);
or U38297 (N_38297,N_31758,N_31949);
xor U38298 (N_38298,N_32085,N_33185);
nor U38299 (N_38299,N_34964,N_30180);
nand U38300 (N_38300,N_31048,N_32235);
nor U38301 (N_38301,N_31313,N_32196);
nand U38302 (N_38302,N_31645,N_33357);
and U38303 (N_38303,N_31847,N_31709);
nor U38304 (N_38304,N_30506,N_30238);
and U38305 (N_38305,N_31196,N_30447);
or U38306 (N_38306,N_33995,N_34267);
nand U38307 (N_38307,N_33810,N_34221);
and U38308 (N_38308,N_30377,N_33578);
nand U38309 (N_38309,N_34426,N_30330);
or U38310 (N_38310,N_31684,N_30447);
nor U38311 (N_38311,N_31286,N_32818);
or U38312 (N_38312,N_31240,N_32466);
nand U38313 (N_38313,N_31041,N_33490);
nand U38314 (N_38314,N_32336,N_31496);
nor U38315 (N_38315,N_32811,N_33560);
nor U38316 (N_38316,N_33849,N_31020);
and U38317 (N_38317,N_30396,N_32766);
and U38318 (N_38318,N_33378,N_30895);
nand U38319 (N_38319,N_31300,N_30683);
nor U38320 (N_38320,N_30372,N_30644);
and U38321 (N_38321,N_34218,N_30825);
or U38322 (N_38322,N_30728,N_30119);
or U38323 (N_38323,N_34383,N_34258);
nor U38324 (N_38324,N_32638,N_31551);
nand U38325 (N_38325,N_31860,N_30997);
nand U38326 (N_38326,N_33622,N_33266);
nand U38327 (N_38327,N_30762,N_33963);
and U38328 (N_38328,N_31420,N_31479);
nor U38329 (N_38329,N_34088,N_32482);
nor U38330 (N_38330,N_33723,N_30347);
xnor U38331 (N_38331,N_32251,N_33570);
or U38332 (N_38332,N_33359,N_33886);
nand U38333 (N_38333,N_34706,N_30167);
xor U38334 (N_38334,N_30019,N_32902);
nand U38335 (N_38335,N_32446,N_34672);
nor U38336 (N_38336,N_31828,N_31366);
or U38337 (N_38337,N_34969,N_33102);
and U38338 (N_38338,N_31867,N_34454);
and U38339 (N_38339,N_31650,N_32150);
nand U38340 (N_38340,N_33537,N_32478);
or U38341 (N_38341,N_30646,N_34933);
nand U38342 (N_38342,N_34942,N_34513);
or U38343 (N_38343,N_31465,N_30411);
or U38344 (N_38344,N_30179,N_32389);
xnor U38345 (N_38345,N_31385,N_33283);
or U38346 (N_38346,N_32287,N_34009);
nor U38347 (N_38347,N_30133,N_32566);
nor U38348 (N_38348,N_31001,N_31281);
or U38349 (N_38349,N_32841,N_30412);
nand U38350 (N_38350,N_34598,N_31122);
nor U38351 (N_38351,N_33796,N_30790);
or U38352 (N_38352,N_34179,N_33479);
nand U38353 (N_38353,N_31085,N_31885);
nand U38354 (N_38354,N_30793,N_33104);
or U38355 (N_38355,N_30370,N_34076);
nor U38356 (N_38356,N_31476,N_30021);
and U38357 (N_38357,N_32171,N_33331);
and U38358 (N_38358,N_34187,N_33790);
nor U38359 (N_38359,N_32421,N_34518);
or U38360 (N_38360,N_33900,N_31611);
and U38361 (N_38361,N_32981,N_33402);
nor U38362 (N_38362,N_30529,N_30122);
xnor U38363 (N_38363,N_34012,N_30879);
or U38364 (N_38364,N_30542,N_30275);
and U38365 (N_38365,N_32181,N_34270);
nor U38366 (N_38366,N_30650,N_33654);
nand U38367 (N_38367,N_34996,N_33533);
nand U38368 (N_38368,N_33726,N_33811);
or U38369 (N_38369,N_33003,N_33037);
and U38370 (N_38370,N_31068,N_33308);
and U38371 (N_38371,N_33883,N_30343);
xor U38372 (N_38372,N_31007,N_32698);
and U38373 (N_38373,N_33055,N_34649);
and U38374 (N_38374,N_34943,N_30201);
and U38375 (N_38375,N_31964,N_31290);
nand U38376 (N_38376,N_33183,N_33344);
xor U38377 (N_38377,N_32223,N_30032);
nor U38378 (N_38378,N_33377,N_30595);
nand U38379 (N_38379,N_30004,N_34254);
nor U38380 (N_38380,N_33514,N_34923);
nor U38381 (N_38381,N_34630,N_31301);
nand U38382 (N_38382,N_32879,N_32632);
or U38383 (N_38383,N_33261,N_34478);
and U38384 (N_38384,N_30765,N_30803);
xnor U38385 (N_38385,N_30130,N_30484);
and U38386 (N_38386,N_31605,N_30175);
or U38387 (N_38387,N_34590,N_31476);
nand U38388 (N_38388,N_33116,N_32384);
nand U38389 (N_38389,N_34390,N_30365);
xor U38390 (N_38390,N_33852,N_33105);
nand U38391 (N_38391,N_34246,N_34847);
nand U38392 (N_38392,N_32814,N_32160);
and U38393 (N_38393,N_33990,N_33079);
or U38394 (N_38394,N_30010,N_30857);
nor U38395 (N_38395,N_33376,N_32572);
and U38396 (N_38396,N_34485,N_31800);
nand U38397 (N_38397,N_32657,N_31960);
nor U38398 (N_38398,N_33725,N_33800);
nor U38399 (N_38399,N_33395,N_33023);
xor U38400 (N_38400,N_34462,N_30503);
nand U38401 (N_38401,N_31781,N_30721);
nand U38402 (N_38402,N_31128,N_31267);
and U38403 (N_38403,N_33760,N_31783);
and U38404 (N_38404,N_30683,N_34390);
nand U38405 (N_38405,N_30132,N_32290);
nand U38406 (N_38406,N_34437,N_30797);
nand U38407 (N_38407,N_30374,N_31293);
and U38408 (N_38408,N_32692,N_30263);
xor U38409 (N_38409,N_34398,N_30136);
or U38410 (N_38410,N_34718,N_32003);
nand U38411 (N_38411,N_32957,N_30002);
nor U38412 (N_38412,N_31128,N_34732);
nor U38413 (N_38413,N_30053,N_31698);
and U38414 (N_38414,N_31783,N_30880);
nand U38415 (N_38415,N_33842,N_31639);
or U38416 (N_38416,N_30903,N_30881);
and U38417 (N_38417,N_34791,N_31675);
nor U38418 (N_38418,N_34624,N_33687);
and U38419 (N_38419,N_30646,N_34771);
and U38420 (N_38420,N_30747,N_31357);
and U38421 (N_38421,N_34017,N_30671);
or U38422 (N_38422,N_34000,N_34080);
nor U38423 (N_38423,N_34297,N_30013);
and U38424 (N_38424,N_33125,N_34044);
nand U38425 (N_38425,N_30372,N_34705);
and U38426 (N_38426,N_34637,N_33769);
or U38427 (N_38427,N_33871,N_33423);
xnor U38428 (N_38428,N_32440,N_32827);
nor U38429 (N_38429,N_30296,N_33197);
or U38430 (N_38430,N_30287,N_31866);
nor U38431 (N_38431,N_34926,N_32145);
nand U38432 (N_38432,N_31429,N_31874);
or U38433 (N_38433,N_33036,N_30761);
xnor U38434 (N_38434,N_30238,N_33463);
and U38435 (N_38435,N_30941,N_33135);
nor U38436 (N_38436,N_33745,N_32889);
and U38437 (N_38437,N_30443,N_32086);
nor U38438 (N_38438,N_30820,N_31005);
nor U38439 (N_38439,N_32045,N_30998);
xor U38440 (N_38440,N_30249,N_33235);
nor U38441 (N_38441,N_30331,N_31602);
nor U38442 (N_38442,N_31012,N_32344);
or U38443 (N_38443,N_30453,N_32416);
nand U38444 (N_38444,N_31555,N_34342);
nand U38445 (N_38445,N_33566,N_34018);
and U38446 (N_38446,N_31623,N_30034);
nand U38447 (N_38447,N_33754,N_30055);
nand U38448 (N_38448,N_34737,N_30523);
and U38449 (N_38449,N_34626,N_32345);
or U38450 (N_38450,N_31040,N_34519);
and U38451 (N_38451,N_32829,N_34324);
nand U38452 (N_38452,N_32431,N_31854);
and U38453 (N_38453,N_31135,N_32848);
and U38454 (N_38454,N_33548,N_32401);
nor U38455 (N_38455,N_34211,N_32529);
nor U38456 (N_38456,N_34096,N_30513);
nand U38457 (N_38457,N_31660,N_32543);
xnor U38458 (N_38458,N_33536,N_31108);
xor U38459 (N_38459,N_31834,N_31606);
xnor U38460 (N_38460,N_30347,N_30047);
nand U38461 (N_38461,N_33715,N_33086);
or U38462 (N_38462,N_31558,N_34389);
nand U38463 (N_38463,N_30879,N_31749);
and U38464 (N_38464,N_30962,N_31144);
nand U38465 (N_38465,N_32749,N_33726);
or U38466 (N_38466,N_31700,N_31250);
nand U38467 (N_38467,N_33533,N_34135);
nand U38468 (N_38468,N_32684,N_31024);
nor U38469 (N_38469,N_31865,N_34539);
nand U38470 (N_38470,N_30918,N_31407);
or U38471 (N_38471,N_33296,N_31142);
or U38472 (N_38472,N_34613,N_31320);
and U38473 (N_38473,N_30641,N_33888);
and U38474 (N_38474,N_33671,N_32246);
and U38475 (N_38475,N_34687,N_31463);
and U38476 (N_38476,N_33928,N_30159);
nand U38477 (N_38477,N_34933,N_31654);
nor U38478 (N_38478,N_32599,N_31021);
or U38479 (N_38479,N_33562,N_33467);
and U38480 (N_38480,N_30922,N_32785);
or U38481 (N_38481,N_31104,N_32285);
and U38482 (N_38482,N_32170,N_31657);
or U38483 (N_38483,N_32250,N_31781);
xnor U38484 (N_38484,N_34990,N_31303);
or U38485 (N_38485,N_30354,N_32540);
nor U38486 (N_38486,N_30293,N_30264);
and U38487 (N_38487,N_30666,N_30357);
or U38488 (N_38488,N_32704,N_33223);
or U38489 (N_38489,N_31821,N_30396);
xnor U38490 (N_38490,N_33544,N_32048);
nand U38491 (N_38491,N_33363,N_30042);
or U38492 (N_38492,N_34165,N_34314);
nand U38493 (N_38493,N_31901,N_31173);
or U38494 (N_38494,N_30580,N_31308);
or U38495 (N_38495,N_31705,N_33246);
and U38496 (N_38496,N_32045,N_32253);
or U38497 (N_38497,N_34267,N_30275);
or U38498 (N_38498,N_32750,N_30121);
nor U38499 (N_38499,N_31810,N_31561);
nor U38500 (N_38500,N_33054,N_31439);
nor U38501 (N_38501,N_34740,N_34778);
nand U38502 (N_38502,N_30007,N_33427);
and U38503 (N_38503,N_30980,N_30796);
nor U38504 (N_38504,N_31768,N_33185);
and U38505 (N_38505,N_31008,N_30651);
and U38506 (N_38506,N_32470,N_31266);
or U38507 (N_38507,N_33797,N_30493);
nand U38508 (N_38508,N_34939,N_31581);
nor U38509 (N_38509,N_31615,N_32976);
nor U38510 (N_38510,N_33608,N_31222);
or U38511 (N_38511,N_33708,N_30121);
nor U38512 (N_38512,N_30826,N_34869);
nor U38513 (N_38513,N_34640,N_30264);
or U38514 (N_38514,N_34690,N_33694);
xor U38515 (N_38515,N_30358,N_31735);
nor U38516 (N_38516,N_31402,N_33229);
and U38517 (N_38517,N_31189,N_30133);
nor U38518 (N_38518,N_30716,N_30242);
nand U38519 (N_38519,N_34089,N_31637);
or U38520 (N_38520,N_32989,N_31772);
nor U38521 (N_38521,N_32399,N_34820);
and U38522 (N_38522,N_32578,N_30277);
and U38523 (N_38523,N_33759,N_32011);
nor U38524 (N_38524,N_32755,N_33014);
nor U38525 (N_38525,N_32221,N_30330);
nand U38526 (N_38526,N_31877,N_32787);
and U38527 (N_38527,N_34683,N_34932);
nand U38528 (N_38528,N_30372,N_32901);
and U38529 (N_38529,N_34789,N_34257);
nand U38530 (N_38530,N_30994,N_33962);
nor U38531 (N_38531,N_34937,N_32270);
nand U38532 (N_38532,N_33648,N_33406);
and U38533 (N_38533,N_30665,N_34866);
or U38534 (N_38534,N_31796,N_34140);
nor U38535 (N_38535,N_32970,N_34903);
and U38536 (N_38536,N_33770,N_33714);
nand U38537 (N_38537,N_30828,N_33203);
or U38538 (N_38538,N_31725,N_30264);
or U38539 (N_38539,N_31479,N_33033);
or U38540 (N_38540,N_33376,N_33293);
nor U38541 (N_38541,N_32745,N_34067);
or U38542 (N_38542,N_34722,N_31057);
nor U38543 (N_38543,N_33914,N_32455);
nor U38544 (N_38544,N_34702,N_34731);
or U38545 (N_38545,N_32754,N_30267);
and U38546 (N_38546,N_31100,N_31506);
nor U38547 (N_38547,N_31642,N_34173);
and U38548 (N_38548,N_30284,N_32201);
and U38549 (N_38549,N_33022,N_32828);
nand U38550 (N_38550,N_31126,N_30146);
xnor U38551 (N_38551,N_33883,N_33255);
and U38552 (N_38552,N_32607,N_33319);
nor U38553 (N_38553,N_30079,N_30231);
nand U38554 (N_38554,N_30577,N_31402);
and U38555 (N_38555,N_32399,N_33298);
nand U38556 (N_38556,N_31714,N_32753);
nand U38557 (N_38557,N_33543,N_32511);
xnor U38558 (N_38558,N_31502,N_34442);
nand U38559 (N_38559,N_34541,N_33350);
xnor U38560 (N_38560,N_30279,N_31814);
nand U38561 (N_38561,N_32317,N_30444);
nand U38562 (N_38562,N_34336,N_33748);
and U38563 (N_38563,N_32684,N_33445);
nand U38564 (N_38564,N_34391,N_33434);
or U38565 (N_38565,N_34455,N_30220);
nor U38566 (N_38566,N_34220,N_32760);
or U38567 (N_38567,N_34881,N_32252);
xor U38568 (N_38568,N_31930,N_31350);
nand U38569 (N_38569,N_30033,N_33816);
nor U38570 (N_38570,N_33092,N_34061);
nor U38571 (N_38571,N_32214,N_30864);
nor U38572 (N_38572,N_30624,N_33905);
or U38573 (N_38573,N_34860,N_33763);
nand U38574 (N_38574,N_32752,N_30981);
or U38575 (N_38575,N_32300,N_31239);
nor U38576 (N_38576,N_33352,N_30878);
nand U38577 (N_38577,N_34341,N_33670);
or U38578 (N_38578,N_30368,N_34268);
xor U38579 (N_38579,N_31355,N_34600);
or U38580 (N_38580,N_34416,N_31209);
xnor U38581 (N_38581,N_30940,N_31295);
nor U38582 (N_38582,N_31683,N_30077);
nor U38583 (N_38583,N_33785,N_32957);
or U38584 (N_38584,N_33761,N_31138);
or U38585 (N_38585,N_30378,N_33014);
and U38586 (N_38586,N_30923,N_34980);
nand U38587 (N_38587,N_33618,N_32750);
nand U38588 (N_38588,N_31952,N_32258);
and U38589 (N_38589,N_30241,N_34516);
or U38590 (N_38590,N_30888,N_31394);
nand U38591 (N_38591,N_34508,N_30011);
nor U38592 (N_38592,N_34723,N_34576);
and U38593 (N_38593,N_31236,N_31281);
xnor U38594 (N_38594,N_33603,N_30775);
nand U38595 (N_38595,N_34981,N_32447);
or U38596 (N_38596,N_31069,N_30001);
nand U38597 (N_38597,N_32305,N_31650);
or U38598 (N_38598,N_31743,N_31005);
nand U38599 (N_38599,N_30446,N_32178);
and U38600 (N_38600,N_31203,N_30437);
and U38601 (N_38601,N_34339,N_34782);
nand U38602 (N_38602,N_31171,N_31602);
nand U38603 (N_38603,N_31912,N_33891);
or U38604 (N_38604,N_31179,N_30833);
nand U38605 (N_38605,N_33133,N_34305);
and U38606 (N_38606,N_34415,N_33782);
nor U38607 (N_38607,N_33994,N_34347);
and U38608 (N_38608,N_30981,N_33381);
nand U38609 (N_38609,N_31604,N_32599);
and U38610 (N_38610,N_34458,N_32773);
nor U38611 (N_38611,N_31816,N_30202);
and U38612 (N_38612,N_34119,N_33986);
nor U38613 (N_38613,N_30068,N_30896);
nor U38614 (N_38614,N_31233,N_33758);
nand U38615 (N_38615,N_32269,N_31899);
and U38616 (N_38616,N_31567,N_31153);
nor U38617 (N_38617,N_32141,N_30390);
and U38618 (N_38618,N_34413,N_31766);
nand U38619 (N_38619,N_33703,N_30273);
or U38620 (N_38620,N_31975,N_34683);
or U38621 (N_38621,N_34174,N_34789);
or U38622 (N_38622,N_31832,N_30491);
nor U38623 (N_38623,N_33163,N_34135);
nand U38624 (N_38624,N_33192,N_34656);
and U38625 (N_38625,N_34362,N_33393);
nand U38626 (N_38626,N_34581,N_34982);
nor U38627 (N_38627,N_30311,N_30461);
nor U38628 (N_38628,N_33693,N_33554);
and U38629 (N_38629,N_33762,N_34704);
and U38630 (N_38630,N_34404,N_32848);
and U38631 (N_38631,N_34233,N_34123);
nand U38632 (N_38632,N_30078,N_31580);
and U38633 (N_38633,N_32345,N_31536);
and U38634 (N_38634,N_30044,N_34531);
and U38635 (N_38635,N_32681,N_30136);
nand U38636 (N_38636,N_33007,N_30694);
nor U38637 (N_38637,N_34365,N_32891);
nand U38638 (N_38638,N_33547,N_30786);
xnor U38639 (N_38639,N_34095,N_34449);
xor U38640 (N_38640,N_34185,N_32399);
or U38641 (N_38641,N_30937,N_33011);
xor U38642 (N_38642,N_31900,N_31360);
nand U38643 (N_38643,N_32092,N_30394);
or U38644 (N_38644,N_34619,N_30818);
and U38645 (N_38645,N_34629,N_33548);
nand U38646 (N_38646,N_34900,N_34613);
nand U38647 (N_38647,N_34805,N_30743);
nor U38648 (N_38648,N_30850,N_33504);
or U38649 (N_38649,N_33338,N_33132);
or U38650 (N_38650,N_32032,N_30687);
or U38651 (N_38651,N_30998,N_31233);
nand U38652 (N_38652,N_30632,N_32334);
xor U38653 (N_38653,N_30534,N_31026);
or U38654 (N_38654,N_33255,N_31790);
and U38655 (N_38655,N_32298,N_31200);
nand U38656 (N_38656,N_33173,N_30682);
and U38657 (N_38657,N_34973,N_31814);
nand U38658 (N_38658,N_33065,N_34130);
nor U38659 (N_38659,N_31850,N_32828);
and U38660 (N_38660,N_33026,N_34343);
and U38661 (N_38661,N_31543,N_30732);
and U38662 (N_38662,N_32358,N_30514);
xnor U38663 (N_38663,N_33183,N_31374);
nor U38664 (N_38664,N_31355,N_34206);
nor U38665 (N_38665,N_33119,N_32492);
and U38666 (N_38666,N_32952,N_33431);
or U38667 (N_38667,N_32113,N_32197);
nor U38668 (N_38668,N_34443,N_31563);
and U38669 (N_38669,N_30419,N_30992);
nand U38670 (N_38670,N_30144,N_31391);
nor U38671 (N_38671,N_30291,N_31777);
or U38672 (N_38672,N_33670,N_30886);
or U38673 (N_38673,N_33013,N_30919);
and U38674 (N_38674,N_32221,N_34652);
or U38675 (N_38675,N_34486,N_30705);
and U38676 (N_38676,N_30325,N_33737);
xnor U38677 (N_38677,N_30684,N_33267);
nand U38678 (N_38678,N_34912,N_32584);
nand U38679 (N_38679,N_32696,N_32592);
nand U38680 (N_38680,N_32364,N_31402);
nor U38681 (N_38681,N_32119,N_34421);
xor U38682 (N_38682,N_30740,N_30188);
nand U38683 (N_38683,N_34522,N_30104);
nor U38684 (N_38684,N_30149,N_31962);
or U38685 (N_38685,N_32290,N_33707);
xor U38686 (N_38686,N_33057,N_33546);
and U38687 (N_38687,N_30423,N_31165);
nor U38688 (N_38688,N_32685,N_32767);
and U38689 (N_38689,N_30052,N_31050);
nor U38690 (N_38690,N_30739,N_32974);
and U38691 (N_38691,N_30566,N_34272);
nand U38692 (N_38692,N_33872,N_31988);
or U38693 (N_38693,N_31090,N_34346);
nor U38694 (N_38694,N_32208,N_33246);
nor U38695 (N_38695,N_34499,N_31489);
nand U38696 (N_38696,N_34207,N_31952);
nand U38697 (N_38697,N_32804,N_33340);
or U38698 (N_38698,N_34709,N_33909);
nand U38699 (N_38699,N_31236,N_31148);
xnor U38700 (N_38700,N_31667,N_30304);
or U38701 (N_38701,N_34588,N_31281);
and U38702 (N_38702,N_34979,N_34412);
xnor U38703 (N_38703,N_30220,N_30755);
nor U38704 (N_38704,N_33017,N_31185);
nor U38705 (N_38705,N_31083,N_31622);
or U38706 (N_38706,N_33025,N_34365);
and U38707 (N_38707,N_32137,N_32269);
and U38708 (N_38708,N_34821,N_34295);
nand U38709 (N_38709,N_30245,N_30960);
and U38710 (N_38710,N_33795,N_34153);
or U38711 (N_38711,N_31534,N_34173);
and U38712 (N_38712,N_30529,N_30511);
nor U38713 (N_38713,N_32713,N_34618);
nor U38714 (N_38714,N_31434,N_32775);
or U38715 (N_38715,N_31543,N_33175);
or U38716 (N_38716,N_34091,N_33900);
nand U38717 (N_38717,N_30745,N_32561);
nand U38718 (N_38718,N_32333,N_31516);
nand U38719 (N_38719,N_33594,N_32549);
or U38720 (N_38720,N_33934,N_33765);
nor U38721 (N_38721,N_30560,N_32868);
and U38722 (N_38722,N_34759,N_34807);
or U38723 (N_38723,N_34626,N_32641);
xor U38724 (N_38724,N_33869,N_34511);
nor U38725 (N_38725,N_33515,N_31399);
nand U38726 (N_38726,N_31572,N_30825);
or U38727 (N_38727,N_34565,N_34972);
and U38728 (N_38728,N_32627,N_32402);
nand U38729 (N_38729,N_33942,N_30591);
nor U38730 (N_38730,N_31494,N_33988);
nand U38731 (N_38731,N_31169,N_34017);
nand U38732 (N_38732,N_34953,N_30743);
xor U38733 (N_38733,N_34711,N_34517);
nor U38734 (N_38734,N_33768,N_34270);
or U38735 (N_38735,N_33830,N_33812);
and U38736 (N_38736,N_33297,N_31706);
or U38737 (N_38737,N_32106,N_31822);
and U38738 (N_38738,N_30954,N_33801);
or U38739 (N_38739,N_31512,N_30450);
xor U38740 (N_38740,N_34870,N_34494);
nand U38741 (N_38741,N_32684,N_30202);
nor U38742 (N_38742,N_32104,N_33079);
nor U38743 (N_38743,N_34832,N_32232);
nor U38744 (N_38744,N_32020,N_32286);
nor U38745 (N_38745,N_32319,N_32540);
xor U38746 (N_38746,N_33548,N_33608);
or U38747 (N_38747,N_31588,N_34428);
and U38748 (N_38748,N_33601,N_32560);
and U38749 (N_38749,N_33517,N_32349);
nor U38750 (N_38750,N_34783,N_34029);
or U38751 (N_38751,N_32367,N_31765);
nor U38752 (N_38752,N_30683,N_33646);
nand U38753 (N_38753,N_31421,N_34807);
nor U38754 (N_38754,N_31499,N_31483);
nor U38755 (N_38755,N_31112,N_33740);
xnor U38756 (N_38756,N_34527,N_33865);
or U38757 (N_38757,N_32496,N_30804);
xnor U38758 (N_38758,N_30188,N_32296);
or U38759 (N_38759,N_30660,N_31011);
nor U38760 (N_38760,N_34938,N_34740);
and U38761 (N_38761,N_30250,N_30447);
and U38762 (N_38762,N_31774,N_31299);
or U38763 (N_38763,N_32076,N_32120);
nand U38764 (N_38764,N_31998,N_30660);
or U38765 (N_38765,N_31662,N_32834);
nand U38766 (N_38766,N_34588,N_33840);
and U38767 (N_38767,N_33104,N_33959);
nor U38768 (N_38768,N_32311,N_34812);
xor U38769 (N_38769,N_32389,N_31600);
or U38770 (N_38770,N_32180,N_30377);
xnor U38771 (N_38771,N_32054,N_30195);
nand U38772 (N_38772,N_34893,N_32542);
nor U38773 (N_38773,N_34310,N_34879);
or U38774 (N_38774,N_34228,N_34220);
and U38775 (N_38775,N_32639,N_31966);
or U38776 (N_38776,N_32572,N_30632);
and U38777 (N_38777,N_31561,N_33092);
or U38778 (N_38778,N_31217,N_34990);
and U38779 (N_38779,N_34764,N_32961);
xor U38780 (N_38780,N_32234,N_33467);
xnor U38781 (N_38781,N_30573,N_33106);
or U38782 (N_38782,N_32904,N_34657);
nor U38783 (N_38783,N_30884,N_30422);
or U38784 (N_38784,N_31092,N_32276);
nor U38785 (N_38785,N_30266,N_31048);
nand U38786 (N_38786,N_33088,N_34881);
and U38787 (N_38787,N_33759,N_34735);
and U38788 (N_38788,N_33645,N_30402);
nand U38789 (N_38789,N_34346,N_31595);
and U38790 (N_38790,N_33783,N_34809);
nor U38791 (N_38791,N_33508,N_33060);
xnor U38792 (N_38792,N_34753,N_32382);
and U38793 (N_38793,N_34921,N_33280);
nor U38794 (N_38794,N_32664,N_31907);
or U38795 (N_38795,N_31001,N_31024);
nor U38796 (N_38796,N_31664,N_31788);
xor U38797 (N_38797,N_31969,N_32994);
xnor U38798 (N_38798,N_33585,N_33337);
nor U38799 (N_38799,N_33675,N_33045);
or U38800 (N_38800,N_33077,N_31528);
and U38801 (N_38801,N_30339,N_34898);
nand U38802 (N_38802,N_30449,N_34767);
nand U38803 (N_38803,N_30425,N_32650);
or U38804 (N_38804,N_31501,N_34720);
nor U38805 (N_38805,N_31579,N_30929);
xor U38806 (N_38806,N_30794,N_30082);
and U38807 (N_38807,N_34693,N_34151);
nor U38808 (N_38808,N_31429,N_30051);
nand U38809 (N_38809,N_31512,N_31240);
or U38810 (N_38810,N_30020,N_33252);
and U38811 (N_38811,N_31762,N_34821);
nand U38812 (N_38812,N_31817,N_34759);
nand U38813 (N_38813,N_30088,N_31582);
nor U38814 (N_38814,N_31738,N_30633);
and U38815 (N_38815,N_33901,N_31682);
nor U38816 (N_38816,N_34365,N_34937);
or U38817 (N_38817,N_32499,N_30270);
or U38818 (N_38818,N_33741,N_33526);
or U38819 (N_38819,N_31226,N_30541);
and U38820 (N_38820,N_32308,N_30856);
nor U38821 (N_38821,N_33782,N_31788);
xor U38822 (N_38822,N_33649,N_32886);
nand U38823 (N_38823,N_31197,N_31898);
and U38824 (N_38824,N_33697,N_30223);
nand U38825 (N_38825,N_32324,N_31360);
and U38826 (N_38826,N_32479,N_32514);
xor U38827 (N_38827,N_31597,N_34352);
and U38828 (N_38828,N_32439,N_30811);
xor U38829 (N_38829,N_33862,N_31539);
or U38830 (N_38830,N_32958,N_30344);
and U38831 (N_38831,N_33036,N_30744);
and U38832 (N_38832,N_30363,N_34680);
nor U38833 (N_38833,N_33255,N_31130);
and U38834 (N_38834,N_34665,N_31609);
or U38835 (N_38835,N_30702,N_32562);
nor U38836 (N_38836,N_31072,N_34992);
or U38837 (N_38837,N_31974,N_32637);
and U38838 (N_38838,N_31763,N_31378);
nand U38839 (N_38839,N_30613,N_33335);
nor U38840 (N_38840,N_30279,N_32699);
xor U38841 (N_38841,N_33572,N_33384);
nor U38842 (N_38842,N_31492,N_33320);
nand U38843 (N_38843,N_34817,N_31653);
nor U38844 (N_38844,N_32991,N_34367);
or U38845 (N_38845,N_31044,N_33691);
nor U38846 (N_38846,N_33464,N_30997);
nand U38847 (N_38847,N_32491,N_30496);
nand U38848 (N_38848,N_32467,N_34153);
nand U38849 (N_38849,N_33652,N_32511);
nand U38850 (N_38850,N_31319,N_33838);
xor U38851 (N_38851,N_30325,N_33026);
and U38852 (N_38852,N_32914,N_30641);
nor U38853 (N_38853,N_31504,N_32177);
nor U38854 (N_38854,N_31843,N_31007);
nor U38855 (N_38855,N_31994,N_31397);
xnor U38856 (N_38856,N_32076,N_34492);
or U38857 (N_38857,N_34928,N_31604);
or U38858 (N_38858,N_32321,N_30092);
nand U38859 (N_38859,N_31072,N_33042);
nand U38860 (N_38860,N_33492,N_34019);
and U38861 (N_38861,N_33964,N_32339);
nand U38862 (N_38862,N_32286,N_33354);
nor U38863 (N_38863,N_31776,N_31513);
nor U38864 (N_38864,N_32318,N_30897);
or U38865 (N_38865,N_33539,N_31889);
nand U38866 (N_38866,N_31993,N_32431);
nor U38867 (N_38867,N_30767,N_34546);
nand U38868 (N_38868,N_31021,N_33908);
or U38869 (N_38869,N_32360,N_31018);
or U38870 (N_38870,N_30303,N_32374);
nor U38871 (N_38871,N_34684,N_31492);
nor U38872 (N_38872,N_34582,N_30715);
nand U38873 (N_38873,N_33417,N_30292);
nand U38874 (N_38874,N_30987,N_32097);
and U38875 (N_38875,N_34956,N_33757);
nand U38876 (N_38876,N_30760,N_30420);
nor U38877 (N_38877,N_32462,N_31046);
or U38878 (N_38878,N_32994,N_31336);
and U38879 (N_38879,N_34992,N_32484);
nand U38880 (N_38880,N_31719,N_30243);
or U38881 (N_38881,N_32662,N_33888);
nor U38882 (N_38882,N_33836,N_33965);
or U38883 (N_38883,N_32793,N_33921);
and U38884 (N_38884,N_34694,N_32100);
or U38885 (N_38885,N_32485,N_30751);
nor U38886 (N_38886,N_32963,N_33011);
and U38887 (N_38887,N_30887,N_34471);
and U38888 (N_38888,N_30118,N_30021);
xor U38889 (N_38889,N_30400,N_33890);
and U38890 (N_38890,N_34741,N_32879);
nor U38891 (N_38891,N_34765,N_31285);
nand U38892 (N_38892,N_32554,N_31050);
nand U38893 (N_38893,N_32252,N_34427);
and U38894 (N_38894,N_32096,N_32878);
and U38895 (N_38895,N_32351,N_30343);
xnor U38896 (N_38896,N_34521,N_33669);
or U38897 (N_38897,N_34868,N_33366);
and U38898 (N_38898,N_31938,N_30253);
nand U38899 (N_38899,N_31277,N_31522);
xor U38900 (N_38900,N_32280,N_34356);
nor U38901 (N_38901,N_32396,N_32722);
or U38902 (N_38902,N_30873,N_31385);
or U38903 (N_38903,N_34863,N_33027);
nor U38904 (N_38904,N_30527,N_30584);
nor U38905 (N_38905,N_33242,N_33058);
nor U38906 (N_38906,N_33021,N_34316);
or U38907 (N_38907,N_34808,N_30669);
xor U38908 (N_38908,N_33184,N_30143);
or U38909 (N_38909,N_34194,N_31090);
and U38910 (N_38910,N_31688,N_30717);
or U38911 (N_38911,N_30731,N_34097);
or U38912 (N_38912,N_33591,N_34391);
nand U38913 (N_38913,N_34652,N_32122);
and U38914 (N_38914,N_34400,N_30686);
nand U38915 (N_38915,N_34288,N_34856);
or U38916 (N_38916,N_31244,N_34314);
nor U38917 (N_38917,N_31877,N_32081);
nor U38918 (N_38918,N_33341,N_32671);
nand U38919 (N_38919,N_30407,N_33722);
nor U38920 (N_38920,N_34189,N_32838);
or U38921 (N_38921,N_30637,N_31991);
and U38922 (N_38922,N_32878,N_31371);
xnor U38923 (N_38923,N_33139,N_33495);
nand U38924 (N_38924,N_30877,N_31086);
nor U38925 (N_38925,N_34450,N_32167);
nand U38926 (N_38926,N_31640,N_31938);
or U38927 (N_38927,N_33323,N_31087);
or U38928 (N_38928,N_31964,N_32228);
or U38929 (N_38929,N_31917,N_30076);
or U38930 (N_38930,N_34767,N_31106);
or U38931 (N_38931,N_32232,N_33378);
nand U38932 (N_38932,N_30444,N_33355);
and U38933 (N_38933,N_33042,N_33432);
nor U38934 (N_38934,N_32015,N_32969);
nand U38935 (N_38935,N_34576,N_33978);
nand U38936 (N_38936,N_34588,N_30914);
or U38937 (N_38937,N_30786,N_31815);
nand U38938 (N_38938,N_33658,N_30984);
nor U38939 (N_38939,N_32399,N_33558);
and U38940 (N_38940,N_34122,N_34493);
and U38941 (N_38941,N_32456,N_33744);
and U38942 (N_38942,N_34097,N_34742);
and U38943 (N_38943,N_34682,N_32709);
and U38944 (N_38944,N_32377,N_33983);
nor U38945 (N_38945,N_34078,N_31378);
nor U38946 (N_38946,N_31921,N_30586);
xnor U38947 (N_38947,N_31919,N_32152);
nor U38948 (N_38948,N_31467,N_32454);
xnor U38949 (N_38949,N_31099,N_31860);
xnor U38950 (N_38950,N_32370,N_32023);
or U38951 (N_38951,N_32582,N_33751);
xnor U38952 (N_38952,N_33075,N_32702);
xnor U38953 (N_38953,N_33411,N_30759);
xnor U38954 (N_38954,N_33799,N_34122);
and U38955 (N_38955,N_32088,N_31606);
nor U38956 (N_38956,N_32381,N_32720);
and U38957 (N_38957,N_30900,N_32556);
nor U38958 (N_38958,N_34916,N_30489);
or U38959 (N_38959,N_30518,N_31434);
and U38960 (N_38960,N_32871,N_33262);
xor U38961 (N_38961,N_33080,N_34493);
or U38962 (N_38962,N_32713,N_32052);
xor U38963 (N_38963,N_34540,N_30044);
nor U38964 (N_38964,N_31165,N_33544);
nand U38965 (N_38965,N_32015,N_34916);
xnor U38966 (N_38966,N_32552,N_31060);
and U38967 (N_38967,N_34340,N_32851);
nor U38968 (N_38968,N_30052,N_31429);
nor U38969 (N_38969,N_32806,N_34842);
nand U38970 (N_38970,N_33116,N_33869);
xor U38971 (N_38971,N_32200,N_32111);
nor U38972 (N_38972,N_34421,N_33019);
and U38973 (N_38973,N_30730,N_34371);
xor U38974 (N_38974,N_34631,N_33503);
nor U38975 (N_38975,N_32847,N_30557);
nand U38976 (N_38976,N_31071,N_32291);
nand U38977 (N_38977,N_30048,N_30374);
or U38978 (N_38978,N_30296,N_30120);
nor U38979 (N_38979,N_30794,N_31659);
nand U38980 (N_38980,N_31709,N_33147);
nor U38981 (N_38981,N_30516,N_31207);
and U38982 (N_38982,N_34939,N_32337);
nand U38983 (N_38983,N_34177,N_34106);
nor U38984 (N_38984,N_33195,N_32241);
xor U38985 (N_38985,N_32590,N_33109);
and U38986 (N_38986,N_34403,N_34235);
nor U38987 (N_38987,N_31099,N_31020);
nand U38988 (N_38988,N_32940,N_34077);
or U38989 (N_38989,N_30112,N_31540);
xnor U38990 (N_38990,N_33231,N_30056);
and U38991 (N_38991,N_32769,N_32635);
nor U38992 (N_38992,N_31532,N_34499);
nand U38993 (N_38993,N_34289,N_34928);
and U38994 (N_38994,N_32290,N_31191);
nor U38995 (N_38995,N_33138,N_30955);
and U38996 (N_38996,N_32214,N_31684);
and U38997 (N_38997,N_32121,N_34873);
nor U38998 (N_38998,N_32816,N_32861);
nand U38999 (N_38999,N_31459,N_31046);
nor U39000 (N_39000,N_30728,N_34688);
and U39001 (N_39001,N_32054,N_30630);
or U39002 (N_39002,N_32410,N_31997);
and U39003 (N_39003,N_32584,N_32638);
or U39004 (N_39004,N_33348,N_32852);
nand U39005 (N_39005,N_30414,N_34110);
xnor U39006 (N_39006,N_34939,N_33910);
nor U39007 (N_39007,N_31544,N_30062);
or U39008 (N_39008,N_34977,N_33292);
nand U39009 (N_39009,N_32002,N_32966);
and U39010 (N_39010,N_30389,N_31192);
xor U39011 (N_39011,N_32457,N_33772);
and U39012 (N_39012,N_31801,N_30976);
and U39013 (N_39013,N_31206,N_31247);
nor U39014 (N_39014,N_31425,N_33715);
and U39015 (N_39015,N_34244,N_32138);
or U39016 (N_39016,N_32732,N_33913);
or U39017 (N_39017,N_30051,N_30204);
nand U39018 (N_39018,N_32806,N_30508);
and U39019 (N_39019,N_31937,N_30889);
or U39020 (N_39020,N_30448,N_31589);
and U39021 (N_39021,N_34835,N_32290);
and U39022 (N_39022,N_33251,N_33195);
nand U39023 (N_39023,N_34425,N_34715);
nor U39024 (N_39024,N_31143,N_31254);
nand U39025 (N_39025,N_33672,N_34370);
nand U39026 (N_39026,N_32904,N_34498);
nor U39027 (N_39027,N_31306,N_34170);
nor U39028 (N_39028,N_31945,N_31040);
or U39029 (N_39029,N_32650,N_32194);
nor U39030 (N_39030,N_31617,N_33574);
xor U39031 (N_39031,N_30677,N_32145);
and U39032 (N_39032,N_34888,N_33443);
nor U39033 (N_39033,N_32474,N_31613);
or U39034 (N_39034,N_33801,N_31893);
or U39035 (N_39035,N_33955,N_32605);
nor U39036 (N_39036,N_33750,N_34211);
nor U39037 (N_39037,N_31866,N_31323);
nor U39038 (N_39038,N_30044,N_30109);
or U39039 (N_39039,N_30176,N_34021);
nand U39040 (N_39040,N_34119,N_31024);
or U39041 (N_39041,N_32053,N_31327);
or U39042 (N_39042,N_34110,N_32439);
nor U39043 (N_39043,N_31498,N_34160);
and U39044 (N_39044,N_33461,N_31863);
xnor U39045 (N_39045,N_32776,N_34702);
nor U39046 (N_39046,N_33340,N_31194);
or U39047 (N_39047,N_30445,N_30566);
xor U39048 (N_39048,N_31960,N_34821);
or U39049 (N_39049,N_31529,N_33856);
nand U39050 (N_39050,N_33973,N_33357);
or U39051 (N_39051,N_34953,N_34590);
nor U39052 (N_39052,N_31266,N_32520);
and U39053 (N_39053,N_34743,N_31788);
or U39054 (N_39054,N_31422,N_33380);
or U39055 (N_39055,N_30618,N_32396);
nand U39056 (N_39056,N_30510,N_31291);
or U39057 (N_39057,N_30438,N_32473);
nand U39058 (N_39058,N_34125,N_34810);
nand U39059 (N_39059,N_33949,N_34433);
or U39060 (N_39060,N_31685,N_34102);
nand U39061 (N_39061,N_30818,N_31086);
or U39062 (N_39062,N_32720,N_33157);
and U39063 (N_39063,N_32248,N_34824);
and U39064 (N_39064,N_34704,N_31886);
nand U39065 (N_39065,N_32802,N_33262);
or U39066 (N_39066,N_32126,N_32486);
nand U39067 (N_39067,N_32526,N_31581);
nor U39068 (N_39068,N_34251,N_32775);
or U39069 (N_39069,N_34110,N_31377);
or U39070 (N_39070,N_33236,N_34116);
or U39071 (N_39071,N_34167,N_34523);
xnor U39072 (N_39072,N_33795,N_32410);
nand U39073 (N_39073,N_31250,N_32677);
or U39074 (N_39074,N_30270,N_31298);
and U39075 (N_39075,N_30762,N_33572);
and U39076 (N_39076,N_32786,N_33772);
or U39077 (N_39077,N_30442,N_33458);
xor U39078 (N_39078,N_34860,N_31288);
and U39079 (N_39079,N_34661,N_34714);
and U39080 (N_39080,N_33580,N_32678);
or U39081 (N_39081,N_32000,N_31029);
or U39082 (N_39082,N_31302,N_32664);
and U39083 (N_39083,N_32975,N_30958);
or U39084 (N_39084,N_34136,N_32946);
nor U39085 (N_39085,N_31470,N_30182);
nand U39086 (N_39086,N_31732,N_34298);
and U39087 (N_39087,N_30192,N_32325);
or U39088 (N_39088,N_34021,N_30035);
or U39089 (N_39089,N_30018,N_30939);
nand U39090 (N_39090,N_31478,N_30216);
nor U39091 (N_39091,N_33278,N_30969);
and U39092 (N_39092,N_31357,N_34032);
and U39093 (N_39093,N_31896,N_30797);
and U39094 (N_39094,N_33682,N_32725);
or U39095 (N_39095,N_30967,N_32669);
or U39096 (N_39096,N_31501,N_31772);
and U39097 (N_39097,N_34179,N_32843);
nand U39098 (N_39098,N_30173,N_33692);
nor U39099 (N_39099,N_34302,N_30582);
nand U39100 (N_39100,N_34607,N_31121);
or U39101 (N_39101,N_30952,N_30144);
and U39102 (N_39102,N_30494,N_31396);
or U39103 (N_39103,N_30812,N_32199);
and U39104 (N_39104,N_30946,N_31417);
nor U39105 (N_39105,N_34166,N_32794);
or U39106 (N_39106,N_31675,N_34487);
xor U39107 (N_39107,N_34573,N_32110);
or U39108 (N_39108,N_33141,N_30868);
or U39109 (N_39109,N_31897,N_34101);
or U39110 (N_39110,N_31256,N_30290);
xnor U39111 (N_39111,N_33332,N_33791);
nor U39112 (N_39112,N_34790,N_32507);
and U39113 (N_39113,N_32950,N_33586);
nor U39114 (N_39114,N_32689,N_32355);
and U39115 (N_39115,N_32542,N_31111);
and U39116 (N_39116,N_34042,N_33527);
or U39117 (N_39117,N_34494,N_31544);
nand U39118 (N_39118,N_31320,N_33405);
and U39119 (N_39119,N_31923,N_30887);
and U39120 (N_39120,N_34598,N_30541);
or U39121 (N_39121,N_32080,N_33154);
and U39122 (N_39122,N_33695,N_31483);
or U39123 (N_39123,N_31480,N_32536);
nand U39124 (N_39124,N_31873,N_33533);
nand U39125 (N_39125,N_31139,N_34797);
nand U39126 (N_39126,N_31869,N_33628);
nor U39127 (N_39127,N_33710,N_31877);
and U39128 (N_39128,N_32713,N_30026);
nand U39129 (N_39129,N_33964,N_30362);
or U39130 (N_39130,N_30199,N_31204);
and U39131 (N_39131,N_30864,N_33289);
or U39132 (N_39132,N_30299,N_32378);
nor U39133 (N_39133,N_32041,N_32508);
nor U39134 (N_39134,N_32547,N_31825);
nand U39135 (N_39135,N_30775,N_32295);
nor U39136 (N_39136,N_33425,N_34803);
and U39137 (N_39137,N_30555,N_30219);
or U39138 (N_39138,N_31268,N_30685);
or U39139 (N_39139,N_30564,N_30029);
xnor U39140 (N_39140,N_32196,N_33344);
nor U39141 (N_39141,N_34123,N_33740);
or U39142 (N_39142,N_32757,N_33301);
nand U39143 (N_39143,N_33632,N_30496);
and U39144 (N_39144,N_31061,N_31961);
or U39145 (N_39145,N_34290,N_32211);
nand U39146 (N_39146,N_30152,N_33529);
and U39147 (N_39147,N_31159,N_31508);
nand U39148 (N_39148,N_31904,N_33218);
nand U39149 (N_39149,N_32966,N_33127);
nor U39150 (N_39150,N_31374,N_33335);
or U39151 (N_39151,N_32015,N_31837);
or U39152 (N_39152,N_30689,N_34902);
nor U39153 (N_39153,N_30709,N_31624);
nor U39154 (N_39154,N_31321,N_31292);
and U39155 (N_39155,N_32373,N_33689);
or U39156 (N_39156,N_34243,N_32776);
nor U39157 (N_39157,N_30390,N_33873);
and U39158 (N_39158,N_32891,N_33009);
and U39159 (N_39159,N_31650,N_34933);
nand U39160 (N_39160,N_32655,N_30008);
nor U39161 (N_39161,N_31736,N_30271);
or U39162 (N_39162,N_30166,N_34597);
nor U39163 (N_39163,N_30583,N_33201);
and U39164 (N_39164,N_33750,N_32059);
nor U39165 (N_39165,N_32500,N_33776);
xnor U39166 (N_39166,N_31911,N_31306);
and U39167 (N_39167,N_31255,N_32662);
and U39168 (N_39168,N_32629,N_34753);
nand U39169 (N_39169,N_32784,N_34046);
and U39170 (N_39170,N_34110,N_34716);
or U39171 (N_39171,N_33003,N_32521);
nor U39172 (N_39172,N_32139,N_33545);
and U39173 (N_39173,N_31150,N_31439);
nand U39174 (N_39174,N_33430,N_31121);
nand U39175 (N_39175,N_33053,N_34381);
and U39176 (N_39176,N_31298,N_30344);
xor U39177 (N_39177,N_33180,N_30726);
nand U39178 (N_39178,N_33540,N_34471);
or U39179 (N_39179,N_32801,N_31484);
or U39180 (N_39180,N_31193,N_30566);
nor U39181 (N_39181,N_30511,N_34203);
or U39182 (N_39182,N_34651,N_34163);
and U39183 (N_39183,N_32854,N_30169);
and U39184 (N_39184,N_32889,N_31382);
xor U39185 (N_39185,N_31950,N_34355);
or U39186 (N_39186,N_33127,N_33475);
nand U39187 (N_39187,N_31374,N_30780);
nand U39188 (N_39188,N_32238,N_30200);
and U39189 (N_39189,N_33291,N_33123);
and U39190 (N_39190,N_30390,N_33224);
nor U39191 (N_39191,N_32742,N_34761);
or U39192 (N_39192,N_33126,N_31358);
and U39193 (N_39193,N_33225,N_32466);
nor U39194 (N_39194,N_33280,N_33661);
and U39195 (N_39195,N_34048,N_31506);
nand U39196 (N_39196,N_31800,N_34588);
and U39197 (N_39197,N_31711,N_30832);
nor U39198 (N_39198,N_30420,N_32908);
or U39199 (N_39199,N_31817,N_31095);
or U39200 (N_39200,N_32003,N_34252);
or U39201 (N_39201,N_32489,N_32534);
or U39202 (N_39202,N_30802,N_31709);
or U39203 (N_39203,N_34669,N_31920);
or U39204 (N_39204,N_34026,N_31086);
and U39205 (N_39205,N_32573,N_31882);
nor U39206 (N_39206,N_30351,N_32672);
and U39207 (N_39207,N_31489,N_30299);
or U39208 (N_39208,N_30351,N_31271);
and U39209 (N_39209,N_32656,N_33095);
and U39210 (N_39210,N_33256,N_31361);
nand U39211 (N_39211,N_33129,N_30683);
xnor U39212 (N_39212,N_31562,N_34453);
nand U39213 (N_39213,N_34702,N_30903);
nor U39214 (N_39214,N_30712,N_34442);
and U39215 (N_39215,N_32920,N_32636);
nor U39216 (N_39216,N_33321,N_33866);
or U39217 (N_39217,N_31690,N_33766);
nand U39218 (N_39218,N_30754,N_31555);
nand U39219 (N_39219,N_34211,N_34868);
xnor U39220 (N_39220,N_33913,N_33556);
nor U39221 (N_39221,N_32333,N_31009);
and U39222 (N_39222,N_34302,N_30131);
or U39223 (N_39223,N_30484,N_31537);
nand U39224 (N_39224,N_32947,N_34859);
nand U39225 (N_39225,N_34112,N_33844);
and U39226 (N_39226,N_30164,N_32273);
or U39227 (N_39227,N_33067,N_34440);
and U39228 (N_39228,N_30127,N_31964);
nor U39229 (N_39229,N_33232,N_31631);
or U39230 (N_39230,N_34474,N_30865);
nor U39231 (N_39231,N_32535,N_33410);
nand U39232 (N_39232,N_30575,N_33777);
or U39233 (N_39233,N_33991,N_31972);
nor U39234 (N_39234,N_34062,N_32902);
nor U39235 (N_39235,N_31672,N_32463);
or U39236 (N_39236,N_32066,N_30829);
nor U39237 (N_39237,N_30868,N_33696);
and U39238 (N_39238,N_32559,N_31332);
and U39239 (N_39239,N_34338,N_34973);
nand U39240 (N_39240,N_34979,N_34559);
nor U39241 (N_39241,N_34488,N_31181);
xnor U39242 (N_39242,N_34322,N_32395);
and U39243 (N_39243,N_30933,N_33193);
nor U39244 (N_39244,N_30144,N_30071);
or U39245 (N_39245,N_32448,N_31589);
nand U39246 (N_39246,N_30505,N_34891);
nor U39247 (N_39247,N_33582,N_34609);
xor U39248 (N_39248,N_34411,N_32212);
nor U39249 (N_39249,N_34359,N_30342);
nor U39250 (N_39250,N_32877,N_33821);
or U39251 (N_39251,N_33495,N_34733);
nand U39252 (N_39252,N_33457,N_32448);
nor U39253 (N_39253,N_32366,N_34767);
xnor U39254 (N_39254,N_34152,N_33396);
and U39255 (N_39255,N_33121,N_32492);
nor U39256 (N_39256,N_34561,N_32187);
nand U39257 (N_39257,N_32535,N_31355);
xnor U39258 (N_39258,N_34198,N_34295);
and U39259 (N_39259,N_31204,N_32377);
nor U39260 (N_39260,N_34443,N_32654);
and U39261 (N_39261,N_33794,N_33303);
nor U39262 (N_39262,N_30041,N_31424);
or U39263 (N_39263,N_31224,N_32388);
nor U39264 (N_39264,N_31817,N_31069);
nand U39265 (N_39265,N_33719,N_34143);
and U39266 (N_39266,N_34786,N_32543);
and U39267 (N_39267,N_34192,N_32009);
nor U39268 (N_39268,N_34216,N_33184);
and U39269 (N_39269,N_33221,N_33744);
nor U39270 (N_39270,N_30585,N_33665);
or U39271 (N_39271,N_32759,N_33547);
and U39272 (N_39272,N_31516,N_32133);
nor U39273 (N_39273,N_33825,N_32838);
or U39274 (N_39274,N_31064,N_32618);
nor U39275 (N_39275,N_31167,N_33329);
nor U39276 (N_39276,N_32925,N_34309);
and U39277 (N_39277,N_32843,N_33780);
nor U39278 (N_39278,N_32478,N_30863);
xnor U39279 (N_39279,N_31633,N_32425);
and U39280 (N_39280,N_31668,N_34841);
or U39281 (N_39281,N_32401,N_30629);
nand U39282 (N_39282,N_31358,N_33017);
and U39283 (N_39283,N_33019,N_31201);
nand U39284 (N_39284,N_33740,N_34987);
and U39285 (N_39285,N_32781,N_32702);
and U39286 (N_39286,N_34304,N_30411);
or U39287 (N_39287,N_33142,N_30771);
nand U39288 (N_39288,N_33619,N_31946);
and U39289 (N_39289,N_32489,N_32708);
nor U39290 (N_39290,N_31545,N_34588);
xnor U39291 (N_39291,N_30426,N_32317);
and U39292 (N_39292,N_33831,N_31638);
xor U39293 (N_39293,N_32763,N_33069);
and U39294 (N_39294,N_31184,N_30812);
and U39295 (N_39295,N_34555,N_33951);
nand U39296 (N_39296,N_33732,N_30015);
nand U39297 (N_39297,N_33568,N_32009);
and U39298 (N_39298,N_33688,N_34807);
xnor U39299 (N_39299,N_34400,N_30913);
and U39300 (N_39300,N_34553,N_31966);
nand U39301 (N_39301,N_34290,N_34591);
nor U39302 (N_39302,N_34628,N_33347);
xnor U39303 (N_39303,N_30550,N_30146);
nand U39304 (N_39304,N_31561,N_30444);
nor U39305 (N_39305,N_32821,N_33636);
and U39306 (N_39306,N_34779,N_33170);
or U39307 (N_39307,N_31176,N_31599);
nand U39308 (N_39308,N_31784,N_34240);
nand U39309 (N_39309,N_32121,N_33589);
nor U39310 (N_39310,N_33143,N_32564);
or U39311 (N_39311,N_34166,N_32053);
or U39312 (N_39312,N_33780,N_30822);
and U39313 (N_39313,N_31659,N_32838);
and U39314 (N_39314,N_31858,N_30877);
xnor U39315 (N_39315,N_31250,N_34752);
or U39316 (N_39316,N_31222,N_33636);
and U39317 (N_39317,N_31236,N_31830);
nor U39318 (N_39318,N_34008,N_34368);
nor U39319 (N_39319,N_33262,N_31073);
or U39320 (N_39320,N_31667,N_31551);
nand U39321 (N_39321,N_32639,N_30209);
nand U39322 (N_39322,N_31869,N_34375);
and U39323 (N_39323,N_31947,N_33857);
or U39324 (N_39324,N_33895,N_33557);
and U39325 (N_39325,N_31125,N_32108);
nor U39326 (N_39326,N_33338,N_34155);
nand U39327 (N_39327,N_33323,N_30288);
nor U39328 (N_39328,N_33345,N_34232);
nand U39329 (N_39329,N_34275,N_30441);
and U39330 (N_39330,N_33764,N_30403);
xnor U39331 (N_39331,N_31380,N_33533);
and U39332 (N_39332,N_34954,N_31241);
xor U39333 (N_39333,N_34579,N_33383);
or U39334 (N_39334,N_30910,N_30022);
nand U39335 (N_39335,N_30524,N_30866);
or U39336 (N_39336,N_30433,N_31149);
nor U39337 (N_39337,N_34300,N_32709);
xor U39338 (N_39338,N_30712,N_31033);
and U39339 (N_39339,N_31480,N_31380);
nand U39340 (N_39340,N_33754,N_33189);
or U39341 (N_39341,N_30262,N_34300);
xnor U39342 (N_39342,N_31856,N_30703);
or U39343 (N_39343,N_34287,N_30722);
nand U39344 (N_39344,N_30273,N_30113);
nor U39345 (N_39345,N_33349,N_31570);
nand U39346 (N_39346,N_32611,N_32229);
or U39347 (N_39347,N_30270,N_33642);
nand U39348 (N_39348,N_31924,N_31300);
xor U39349 (N_39349,N_31526,N_33849);
nand U39350 (N_39350,N_33385,N_33887);
and U39351 (N_39351,N_30705,N_30229);
and U39352 (N_39352,N_30142,N_32879);
and U39353 (N_39353,N_33873,N_30720);
xor U39354 (N_39354,N_32418,N_31744);
nor U39355 (N_39355,N_32076,N_32043);
and U39356 (N_39356,N_31452,N_32451);
or U39357 (N_39357,N_33380,N_33286);
and U39358 (N_39358,N_34990,N_31563);
or U39359 (N_39359,N_30276,N_34852);
nand U39360 (N_39360,N_34174,N_31554);
or U39361 (N_39361,N_34897,N_31949);
or U39362 (N_39362,N_33989,N_34316);
nor U39363 (N_39363,N_31414,N_31945);
and U39364 (N_39364,N_32704,N_30899);
and U39365 (N_39365,N_31905,N_30422);
nand U39366 (N_39366,N_33953,N_31167);
nand U39367 (N_39367,N_32052,N_32100);
and U39368 (N_39368,N_31098,N_33759);
and U39369 (N_39369,N_34006,N_30136);
nor U39370 (N_39370,N_31271,N_34837);
nor U39371 (N_39371,N_34656,N_33248);
and U39372 (N_39372,N_30656,N_33326);
xor U39373 (N_39373,N_30183,N_30267);
and U39374 (N_39374,N_33746,N_33066);
nor U39375 (N_39375,N_30802,N_31871);
nor U39376 (N_39376,N_33574,N_33130);
and U39377 (N_39377,N_30061,N_31862);
nor U39378 (N_39378,N_34666,N_30008);
nand U39379 (N_39379,N_32555,N_31304);
nand U39380 (N_39380,N_34918,N_32652);
and U39381 (N_39381,N_33781,N_30709);
nand U39382 (N_39382,N_34756,N_30205);
or U39383 (N_39383,N_30743,N_31654);
or U39384 (N_39384,N_33126,N_32586);
nor U39385 (N_39385,N_30839,N_30956);
xnor U39386 (N_39386,N_32982,N_32860);
and U39387 (N_39387,N_33644,N_32936);
xnor U39388 (N_39388,N_30999,N_33301);
nor U39389 (N_39389,N_31376,N_33926);
nand U39390 (N_39390,N_34723,N_34122);
nand U39391 (N_39391,N_34361,N_34374);
or U39392 (N_39392,N_32782,N_32893);
nor U39393 (N_39393,N_32620,N_33457);
nor U39394 (N_39394,N_31823,N_32167);
and U39395 (N_39395,N_30127,N_33501);
nor U39396 (N_39396,N_31345,N_31924);
and U39397 (N_39397,N_34446,N_33696);
nor U39398 (N_39398,N_33990,N_33611);
nor U39399 (N_39399,N_30085,N_34122);
and U39400 (N_39400,N_31175,N_34328);
or U39401 (N_39401,N_34805,N_32747);
nand U39402 (N_39402,N_30819,N_34558);
nor U39403 (N_39403,N_30411,N_31397);
xnor U39404 (N_39404,N_31823,N_33073);
nand U39405 (N_39405,N_32645,N_31375);
or U39406 (N_39406,N_34246,N_30042);
or U39407 (N_39407,N_31066,N_30887);
nand U39408 (N_39408,N_31440,N_33730);
nor U39409 (N_39409,N_33608,N_30264);
and U39410 (N_39410,N_31667,N_33270);
and U39411 (N_39411,N_33632,N_34614);
nand U39412 (N_39412,N_33871,N_31308);
nand U39413 (N_39413,N_31818,N_32447);
and U39414 (N_39414,N_33248,N_34984);
nor U39415 (N_39415,N_34180,N_33894);
xnor U39416 (N_39416,N_34245,N_34723);
and U39417 (N_39417,N_32864,N_33178);
and U39418 (N_39418,N_31594,N_30229);
or U39419 (N_39419,N_31790,N_33900);
and U39420 (N_39420,N_31704,N_33306);
and U39421 (N_39421,N_32891,N_31195);
or U39422 (N_39422,N_32155,N_31054);
nor U39423 (N_39423,N_34179,N_31917);
nand U39424 (N_39424,N_33501,N_31253);
and U39425 (N_39425,N_30994,N_30310);
nand U39426 (N_39426,N_30296,N_32905);
xor U39427 (N_39427,N_31556,N_31209);
nand U39428 (N_39428,N_32284,N_31187);
or U39429 (N_39429,N_31133,N_30457);
xor U39430 (N_39430,N_32791,N_31142);
nand U39431 (N_39431,N_31256,N_31315);
nand U39432 (N_39432,N_31606,N_32872);
xnor U39433 (N_39433,N_30600,N_30897);
xor U39434 (N_39434,N_32259,N_33119);
or U39435 (N_39435,N_31483,N_30762);
or U39436 (N_39436,N_30252,N_32478);
nand U39437 (N_39437,N_30700,N_32300);
nor U39438 (N_39438,N_32071,N_31219);
nand U39439 (N_39439,N_30777,N_34691);
nor U39440 (N_39440,N_30657,N_33408);
or U39441 (N_39441,N_30804,N_30295);
nand U39442 (N_39442,N_30712,N_30290);
nand U39443 (N_39443,N_32665,N_32609);
nor U39444 (N_39444,N_32966,N_33086);
and U39445 (N_39445,N_34659,N_34823);
nor U39446 (N_39446,N_34318,N_33643);
nand U39447 (N_39447,N_32114,N_34691);
nor U39448 (N_39448,N_31010,N_31875);
nand U39449 (N_39449,N_32020,N_32422);
nor U39450 (N_39450,N_31740,N_32026);
nand U39451 (N_39451,N_30307,N_34591);
and U39452 (N_39452,N_31879,N_33202);
xnor U39453 (N_39453,N_34016,N_34319);
and U39454 (N_39454,N_34209,N_32368);
nand U39455 (N_39455,N_30374,N_30355);
nand U39456 (N_39456,N_30986,N_33224);
or U39457 (N_39457,N_30109,N_32604);
and U39458 (N_39458,N_34464,N_30556);
and U39459 (N_39459,N_33174,N_30114);
nand U39460 (N_39460,N_30158,N_31084);
and U39461 (N_39461,N_31042,N_32765);
and U39462 (N_39462,N_33138,N_30416);
xnor U39463 (N_39463,N_32609,N_33069);
xnor U39464 (N_39464,N_33573,N_32760);
nand U39465 (N_39465,N_32240,N_32791);
or U39466 (N_39466,N_31176,N_32520);
or U39467 (N_39467,N_30859,N_34419);
nor U39468 (N_39468,N_31277,N_33698);
or U39469 (N_39469,N_30372,N_31794);
and U39470 (N_39470,N_32051,N_33192);
nor U39471 (N_39471,N_31563,N_34405);
nor U39472 (N_39472,N_33230,N_31727);
nor U39473 (N_39473,N_33913,N_31087);
and U39474 (N_39474,N_33558,N_34996);
or U39475 (N_39475,N_30262,N_33559);
and U39476 (N_39476,N_33235,N_30378);
nand U39477 (N_39477,N_32471,N_34356);
nand U39478 (N_39478,N_30870,N_30804);
and U39479 (N_39479,N_31990,N_32269);
or U39480 (N_39480,N_33502,N_33998);
nand U39481 (N_39481,N_31411,N_32768);
or U39482 (N_39482,N_34137,N_31669);
and U39483 (N_39483,N_33704,N_32949);
nand U39484 (N_39484,N_32992,N_30832);
nor U39485 (N_39485,N_33812,N_34083);
or U39486 (N_39486,N_33881,N_33474);
and U39487 (N_39487,N_30958,N_30551);
and U39488 (N_39488,N_32695,N_30407);
and U39489 (N_39489,N_31743,N_33121);
and U39490 (N_39490,N_34287,N_32942);
nand U39491 (N_39491,N_32554,N_30585);
nand U39492 (N_39492,N_32267,N_34577);
and U39493 (N_39493,N_30834,N_31087);
or U39494 (N_39494,N_31289,N_33156);
or U39495 (N_39495,N_30505,N_33651);
nor U39496 (N_39496,N_31984,N_30174);
nor U39497 (N_39497,N_34336,N_30283);
nand U39498 (N_39498,N_34987,N_33300);
nor U39499 (N_39499,N_34832,N_32448);
nor U39500 (N_39500,N_33569,N_32485);
nor U39501 (N_39501,N_33116,N_34865);
nor U39502 (N_39502,N_33400,N_33072);
or U39503 (N_39503,N_34603,N_30199);
nand U39504 (N_39504,N_33887,N_30233);
or U39505 (N_39505,N_30627,N_32652);
or U39506 (N_39506,N_33364,N_32563);
nor U39507 (N_39507,N_32634,N_32518);
or U39508 (N_39508,N_31580,N_34187);
or U39509 (N_39509,N_32100,N_32047);
nor U39510 (N_39510,N_32396,N_32176);
or U39511 (N_39511,N_30133,N_30198);
or U39512 (N_39512,N_30067,N_31244);
nand U39513 (N_39513,N_34551,N_32342);
or U39514 (N_39514,N_33080,N_34479);
nor U39515 (N_39515,N_33633,N_34780);
nor U39516 (N_39516,N_32413,N_30721);
nand U39517 (N_39517,N_30143,N_34456);
or U39518 (N_39518,N_31299,N_32878);
and U39519 (N_39519,N_34321,N_31136);
or U39520 (N_39520,N_34859,N_32386);
nor U39521 (N_39521,N_31053,N_30821);
and U39522 (N_39522,N_31831,N_32638);
and U39523 (N_39523,N_32832,N_33946);
nor U39524 (N_39524,N_30398,N_33175);
xnor U39525 (N_39525,N_34201,N_32127);
and U39526 (N_39526,N_33911,N_30051);
or U39527 (N_39527,N_33668,N_31908);
and U39528 (N_39528,N_33899,N_32976);
nor U39529 (N_39529,N_32542,N_34400);
xor U39530 (N_39530,N_33249,N_32531);
and U39531 (N_39531,N_31039,N_32684);
nor U39532 (N_39532,N_32153,N_32081);
or U39533 (N_39533,N_32034,N_33952);
and U39534 (N_39534,N_34952,N_34441);
nor U39535 (N_39535,N_30691,N_33317);
or U39536 (N_39536,N_33119,N_34720);
nor U39537 (N_39537,N_34940,N_31280);
or U39538 (N_39538,N_33562,N_33144);
and U39539 (N_39539,N_30071,N_33474);
nor U39540 (N_39540,N_34752,N_31007);
nor U39541 (N_39541,N_34627,N_33562);
xnor U39542 (N_39542,N_33046,N_33541);
nand U39543 (N_39543,N_32308,N_34053);
nand U39544 (N_39544,N_34601,N_30399);
nor U39545 (N_39545,N_33164,N_32033);
nand U39546 (N_39546,N_32432,N_32631);
and U39547 (N_39547,N_32456,N_34209);
nand U39548 (N_39548,N_30731,N_34142);
nand U39549 (N_39549,N_32075,N_34602);
and U39550 (N_39550,N_31020,N_34786);
and U39551 (N_39551,N_32051,N_34732);
or U39552 (N_39552,N_33193,N_33574);
nor U39553 (N_39553,N_33902,N_33142);
nand U39554 (N_39554,N_30760,N_32534);
nand U39555 (N_39555,N_32300,N_32124);
and U39556 (N_39556,N_32160,N_33509);
and U39557 (N_39557,N_32720,N_34835);
and U39558 (N_39558,N_32494,N_30222);
nor U39559 (N_39559,N_30311,N_31784);
and U39560 (N_39560,N_34287,N_34153);
or U39561 (N_39561,N_34287,N_30931);
or U39562 (N_39562,N_30647,N_31523);
or U39563 (N_39563,N_32358,N_33083);
nor U39564 (N_39564,N_34683,N_33608);
xnor U39565 (N_39565,N_30653,N_30634);
xnor U39566 (N_39566,N_33828,N_31423);
nand U39567 (N_39567,N_30522,N_33291);
xnor U39568 (N_39568,N_34029,N_31028);
nor U39569 (N_39569,N_34378,N_32598);
or U39570 (N_39570,N_34404,N_33143);
xor U39571 (N_39571,N_32081,N_31077);
nand U39572 (N_39572,N_31032,N_33417);
nand U39573 (N_39573,N_32780,N_34506);
nor U39574 (N_39574,N_33782,N_31511);
nand U39575 (N_39575,N_34503,N_33508);
and U39576 (N_39576,N_32368,N_30745);
nor U39577 (N_39577,N_31804,N_31285);
and U39578 (N_39578,N_34293,N_31654);
or U39579 (N_39579,N_31357,N_32874);
nand U39580 (N_39580,N_32180,N_31912);
nand U39581 (N_39581,N_33133,N_30214);
and U39582 (N_39582,N_32151,N_31548);
and U39583 (N_39583,N_30899,N_33687);
and U39584 (N_39584,N_31609,N_31965);
and U39585 (N_39585,N_30035,N_34646);
nor U39586 (N_39586,N_32390,N_30758);
nand U39587 (N_39587,N_30769,N_33812);
nand U39588 (N_39588,N_30033,N_30696);
or U39589 (N_39589,N_30399,N_33692);
or U39590 (N_39590,N_32043,N_31441);
nor U39591 (N_39591,N_33985,N_32709);
nand U39592 (N_39592,N_34712,N_30930);
nor U39593 (N_39593,N_33283,N_31101);
nor U39594 (N_39594,N_31148,N_31844);
nor U39595 (N_39595,N_32777,N_33465);
nand U39596 (N_39596,N_34404,N_34694);
nor U39597 (N_39597,N_34830,N_30070);
and U39598 (N_39598,N_32959,N_34116);
and U39599 (N_39599,N_30229,N_33026);
nor U39600 (N_39600,N_31055,N_32859);
nor U39601 (N_39601,N_33205,N_31120);
or U39602 (N_39602,N_32370,N_33482);
or U39603 (N_39603,N_33623,N_33091);
nor U39604 (N_39604,N_34261,N_32318);
or U39605 (N_39605,N_32394,N_31427);
and U39606 (N_39606,N_33981,N_30875);
xor U39607 (N_39607,N_33167,N_34532);
or U39608 (N_39608,N_34096,N_32172);
nand U39609 (N_39609,N_32483,N_30030);
nand U39610 (N_39610,N_33044,N_34588);
nand U39611 (N_39611,N_32784,N_33236);
or U39612 (N_39612,N_34305,N_33485);
xnor U39613 (N_39613,N_34136,N_34982);
or U39614 (N_39614,N_30291,N_30511);
or U39615 (N_39615,N_32601,N_31636);
nand U39616 (N_39616,N_31407,N_30240);
xnor U39617 (N_39617,N_31247,N_30978);
nand U39618 (N_39618,N_32979,N_32152);
nor U39619 (N_39619,N_31438,N_31094);
and U39620 (N_39620,N_31255,N_34573);
nor U39621 (N_39621,N_31327,N_34343);
or U39622 (N_39622,N_33794,N_31729);
nand U39623 (N_39623,N_30145,N_30118);
and U39624 (N_39624,N_33754,N_31605);
or U39625 (N_39625,N_31827,N_30230);
or U39626 (N_39626,N_34921,N_32863);
xor U39627 (N_39627,N_32563,N_32318);
xnor U39628 (N_39628,N_34223,N_30017);
nor U39629 (N_39629,N_33358,N_34955);
nor U39630 (N_39630,N_34863,N_33988);
nor U39631 (N_39631,N_33680,N_30042);
xnor U39632 (N_39632,N_33886,N_30133);
nor U39633 (N_39633,N_30916,N_32025);
or U39634 (N_39634,N_30144,N_30081);
nor U39635 (N_39635,N_30910,N_30051);
and U39636 (N_39636,N_32956,N_34476);
nor U39637 (N_39637,N_32574,N_34721);
or U39638 (N_39638,N_33299,N_32919);
nor U39639 (N_39639,N_32370,N_32620);
and U39640 (N_39640,N_30179,N_33621);
nand U39641 (N_39641,N_34653,N_33245);
xnor U39642 (N_39642,N_34904,N_31941);
nand U39643 (N_39643,N_33862,N_30228);
or U39644 (N_39644,N_30011,N_33727);
or U39645 (N_39645,N_31251,N_32792);
nor U39646 (N_39646,N_30420,N_31696);
nand U39647 (N_39647,N_31349,N_32953);
xnor U39648 (N_39648,N_31448,N_32622);
or U39649 (N_39649,N_31626,N_34767);
nand U39650 (N_39650,N_34533,N_33818);
nor U39651 (N_39651,N_33980,N_34002);
or U39652 (N_39652,N_32051,N_33097);
nor U39653 (N_39653,N_31320,N_31294);
nand U39654 (N_39654,N_32876,N_31201);
and U39655 (N_39655,N_31901,N_31965);
or U39656 (N_39656,N_34735,N_32299);
nor U39657 (N_39657,N_33131,N_30393);
nand U39658 (N_39658,N_33124,N_34244);
and U39659 (N_39659,N_31852,N_31561);
nor U39660 (N_39660,N_34380,N_34234);
or U39661 (N_39661,N_32465,N_31040);
or U39662 (N_39662,N_33583,N_30456);
and U39663 (N_39663,N_30444,N_30584);
or U39664 (N_39664,N_33305,N_33594);
nand U39665 (N_39665,N_31108,N_33614);
nand U39666 (N_39666,N_33934,N_34651);
or U39667 (N_39667,N_30222,N_34938);
nor U39668 (N_39668,N_31962,N_31135);
nor U39669 (N_39669,N_31294,N_34937);
and U39670 (N_39670,N_31794,N_34789);
nand U39671 (N_39671,N_32271,N_34849);
nor U39672 (N_39672,N_31219,N_31034);
nand U39673 (N_39673,N_30323,N_34212);
and U39674 (N_39674,N_31677,N_31288);
nor U39675 (N_39675,N_33835,N_34756);
nor U39676 (N_39676,N_32255,N_32776);
and U39677 (N_39677,N_33338,N_33559);
and U39678 (N_39678,N_31119,N_33489);
nand U39679 (N_39679,N_33607,N_33709);
and U39680 (N_39680,N_34686,N_30917);
and U39681 (N_39681,N_33621,N_34429);
or U39682 (N_39682,N_33952,N_30795);
nor U39683 (N_39683,N_33466,N_32891);
and U39684 (N_39684,N_30803,N_30395);
and U39685 (N_39685,N_32787,N_32133);
and U39686 (N_39686,N_33631,N_30371);
nand U39687 (N_39687,N_32931,N_32965);
or U39688 (N_39688,N_31538,N_30417);
nor U39689 (N_39689,N_32590,N_32634);
nand U39690 (N_39690,N_32784,N_34767);
nand U39691 (N_39691,N_34802,N_30768);
or U39692 (N_39692,N_34389,N_34520);
and U39693 (N_39693,N_32349,N_33796);
nand U39694 (N_39694,N_34286,N_32820);
xnor U39695 (N_39695,N_32739,N_30335);
and U39696 (N_39696,N_32176,N_34823);
nor U39697 (N_39697,N_31540,N_34123);
nor U39698 (N_39698,N_32980,N_32257);
and U39699 (N_39699,N_33957,N_33536);
nand U39700 (N_39700,N_33051,N_31065);
nor U39701 (N_39701,N_31555,N_32358);
nand U39702 (N_39702,N_30245,N_32330);
and U39703 (N_39703,N_33057,N_34906);
nor U39704 (N_39704,N_34708,N_34175);
and U39705 (N_39705,N_31354,N_31623);
or U39706 (N_39706,N_32104,N_33021);
nand U39707 (N_39707,N_31534,N_33516);
nand U39708 (N_39708,N_30372,N_31659);
nor U39709 (N_39709,N_33965,N_33363);
nor U39710 (N_39710,N_33273,N_31477);
nand U39711 (N_39711,N_31869,N_30174);
nor U39712 (N_39712,N_30688,N_33369);
xor U39713 (N_39713,N_30887,N_31032);
nor U39714 (N_39714,N_33931,N_30833);
nor U39715 (N_39715,N_30169,N_33506);
nor U39716 (N_39716,N_34384,N_34236);
and U39717 (N_39717,N_31984,N_30760);
nor U39718 (N_39718,N_31401,N_33172);
nand U39719 (N_39719,N_32673,N_31510);
or U39720 (N_39720,N_31079,N_33308);
nand U39721 (N_39721,N_30888,N_31799);
nand U39722 (N_39722,N_30566,N_34190);
nor U39723 (N_39723,N_32291,N_30028);
nor U39724 (N_39724,N_31044,N_30550);
nor U39725 (N_39725,N_32534,N_32195);
or U39726 (N_39726,N_32788,N_34935);
nand U39727 (N_39727,N_30385,N_33361);
nand U39728 (N_39728,N_32369,N_31425);
or U39729 (N_39729,N_32604,N_30229);
nand U39730 (N_39730,N_30795,N_34998);
nor U39731 (N_39731,N_34066,N_34521);
or U39732 (N_39732,N_34718,N_31014);
or U39733 (N_39733,N_30699,N_30169);
nor U39734 (N_39734,N_32125,N_30923);
and U39735 (N_39735,N_30959,N_33249);
or U39736 (N_39736,N_32400,N_33724);
xnor U39737 (N_39737,N_32069,N_31426);
nor U39738 (N_39738,N_32467,N_31485);
xnor U39739 (N_39739,N_30028,N_30834);
nand U39740 (N_39740,N_33799,N_32871);
nor U39741 (N_39741,N_31133,N_31958);
nor U39742 (N_39742,N_33669,N_34505);
nor U39743 (N_39743,N_30792,N_31988);
xor U39744 (N_39744,N_33885,N_32063);
nor U39745 (N_39745,N_34835,N_30435);
nand U39746 (N_39746,N_31317,N_33793);
and U39747 (N_39747,N_30444,N_31712);
or U39748 (N_39748,N_32481,N_31813);
nand U39749 (N_39749,N_30524,N_31259);
or U39750 (N_39750,N_33829,N_30011);
and U39751 (N_39751,N_32159,N_34342);
xor U39752 (N_39752,N_31665,N_31596);
and U39753 (N_39753,N_31631,N_32655);
nand U39754 (N_39754,N_30439,N_34996);
and U39755 (N_39755,N_34583,N_30488);
or U39756 (N_39756,N_34903,N_33567);
or U39757 (N_39757,N_33030,N_31366);
or U39758 (N_39758,N_32463,N_33782);
and U39759 (N_39759,N_34356,N_34961);
and U39760 (N_39760,N_33465,N_30432);
nor U39761 (N_39761,N_31451,N_30077);
nor U39762 (N_39762,N_31588,N_34010);
nand U39763 (N_39763,N_33454,N_34952);
and U39764 (N_39764,N_32117,N_33712);
nand U39765 (N_39765,N_32740,N_33301);
and U39766 (N_39766,N_32650,N_30788);
or U39767 (N_39767,N_30895,N_34487);
or U39768 (N_39768,N_31764,N_33342);
and U39769 (N_39769,N_31321,N_31471);
nand U39770 (N_39770,N_30054,N_34008);
and U39771 (N_39771,N_33198,N_30996);
nand U39772 (N_39772,N_34940,N_32124);
or U39773 (N_39773,N_31336,N_33832);
nand U39774 (N_39774,N_34496,N_31141);
nand U39775 (N_39775,N_33034,N_34223);
nand U39776 (N_39776,N_32353,N_34611);
or U39777 (N_39777,N_32258,N_33203);
and U39778 (N_39778,N_33350,N_32131);
nand U39779 (N_39779,N_30877,N_31754);
and U39780 (N_39780,N_34196,N_33989);
nand U39781 (N_39781,N_32270,N_31919);
nand U39782 (N_39782,N_32930,N_31867);
xnor U39783 (N_39783,N_30090,N_30931);
nor U39784 (N_39784,N_33810,N_32639);
nand U39785 (N_39785,N_34568,N_32993);
nand U39786 (N_39786,N_32416,N_34390);
or U39787 (N_39787,N_31922,N_30606);
and U39788 (N_39788,N_31821,N_32759);
xnor U39789 (N_39789,N_31325,N_31073);
and U39790 (N_39790,N_31665,N_32582);
and U39791 (N_39791,N_30955,N_31443);
or U39792 (N_39792,N_33574,N_32775);
nand U39793 (N_39793,N_30528,N_33997);
or U39794 (N_39794,N_34631,N_33270);
or U39795 (N_39795,N_31907,N_33753);
or U39796 (N_39796,N_34430,N_30458);
nor U39797 (N_39797,N_32382,N_30240);
nand U39798 (N_39798,N_32059,N_33067);
or U39799 (N_39799,N_33806,N_31786);
xor U39800 (N_39800,N_32726,N_31153);
and U39801 (N_39801,N_30847,N_34103);
or U39802 (N_39802,N_32671,N_34151);
nor U39803 (N_39803,N_33247,N_31366);
or U39804 (N_39804,N_31084,N_31494);
nand U39805 (N_39805,N_31706,N_33603);
xor U39806 (N_39806,N_32520,N_32991);
and U39807 (N_39807,N_34450,N_32183);
nor U39808 (N_39808,N_34791,N_30936);
nand U39809 (N_39809,N_33816,N_34955);
nor U39810 (N_39810,N_30236,N_31477);
or U39811 (N_39811,N_31128,N_34819);
nand U39812 (N_39812,N_32366,N_34616);
xnor U39813 (N_39813,N_33163,N_31223);
or U39814 (N_39814,N_31849,N_30025);
nor U39815 (N_39815,N_31710,N_32404);
nor U39816 (N_39816,N_30048,N_33250);
and U39817 (N_39817,N_33341,N_32367);
or U39818 (N_39818,N_31156,N_31388);
nor U39819 (N_39819,N_32537,N_34214);
nor U39820 (N_39820,N_30643,N_30147);
nand U39821 (N_39821,N_33308,N_31816);
nand U39822 (N_39822,N_32617,N_31019);
nor U39823 (N_39823,N_34669,N_30611);
and U39824 (N_39824,N_32409,N_33916);
xnor U39825 (N_39825,N_30299,N_32445);
nor U39826 (N_39826,N_30235,N_31896);
nor U39827 (N_39827,N_32672,N_34945);
nor U39828 (N_39828,N_34610,N_33880);
and U39829 (N_39829,N_31969,N_33527);
and U39830 (N_39830,N_34952,N_32340);
nor U39831 (N_39831,N_31686,N_32277);
nand U39832 (N_39832,N_34161,N_34332);
nand U39833 (N_39833,N_30825,N_32220);
or U39834 (N_39834,N_33005,N_31949);
nand U39835 (N_39835,N_34041,N_34188);
nand U39836 (N_39836,N_34683,N_32436);
and U39837 (N_39837,N_31049,N_32987);
or U39838 (N_39838,N_34545,N_34949);
nor U39839 (N_39839,N_33660,N_30782);
nor U39840 (N_39840,N_34366,N_31876);
nand U39841 (N_39841,N_32729,N_32329);
nand U39842 (N_39842,N_31679,N_33802);
nand U39843 (N_39843,N_33560,N_30247);
nand U39844 (N_39844,N_34257,N_33050);
or U39845 (N_39845,N_33764,N_31192);
nand U39846 (N_39846,N_31462,N_30801);
nor U39847 (N_39847,N_34884,N_30824);
and U39848 (N_39848,N_31040,N_34533);
nor U39849 (N_39849,N_31836,N_34308);
nand U39850 (N_39850,N_30081,N_33245);
xor U39851 (N_39851,N_30110,N_32774);
or U39852 (N_39852,N_30745,N_32048);
and U39853 (N_39853,N_31541,N_33377);
nand U39854 (N_39854,N_31659,N_31934);
and U39855 (N_39855,N_33510,N_34245);
and U39856 (N_39856,N_30578,N_30881);
and U39857 (N_39857,N_33588,N_32865);
nand U39858 (N_39858,N_33443,N_32670);
nand U39859 (N_39859,N_33031,N_30792);
or U39860 (N_39860,N_32348,N_30211);
nor U39861 (N_39861,N_34476,N_30302);
and U39862 (N_39862,N_32817,N_32373);
and U39863 (N_39863,N_33557,N_30963);
nand U39864 (N_39864,N_30790,N_33250);
nor U39865 (N_39865,N_32928,N_34910);
or U39866 (N_39866,N_31307,N_30796);
or U39867 (N_39867,N_31176,N_30747);
and U39868 (N_39868,N_30490,N_33225);
nor U39869 (N_39869,N_32707,N_34521);
nor U39870 (N_39870,N_31638,N_34007);
and U39871 (N_39871,N_33151,N_32203);
or U39872 (N_39872,N_30068,N_33156);
nand U39873 (N_39873,N_32365,N_34270);
and U39874 (N_39874,N_31762,N_34922);
or U39875 (N_39875,N_31061,N_31244);
nand U39876 (N_39876,N_31107,N_34001);
and U39877 (N_39877,N_31280,N_34750);
nand U39878 (N_39878,N_33767,N_33125);
or U39879 (N_39879,N_34380,N_34147);
nand U39880 (N_39880,N_33925,N_30374);
nand U39881 (N_39881,N_33306,N_33859);
nor U39882 (N_39882,N_34153,N_34256);
nand U39883 (N_39883,N_32203,N_33628);
nand U39884 (N_39884,N_30741,N_33521);
and U39885 (N_39885,N_34784,N_34666);
nand U39886 (N_39886,N_30430,N_33244);
nand U39887 (N_39887,N_30895,N_34800);
and U39888 (N_39888,N_33520,N_33894);
or U39889 (N_39889,N_33833,N_30430);
or U39890 (N_39890,N_32512,N_33900);
or U39891 (N_39891,N_33472,N_30529);
nor U39892 (N_39892,N_34558,N_30614);
or U39893 (N_39893,N_30895,N_32306);
or U39894 (N_39894,N_31569,N_32488);
and U39895 (N_39895,N_30827,N_33300);
and U39896 (N_39896,N_34355,N_31343);
xor U39897 (N_39897,N_34159,N_32806);
nor U39898 (N_39898,N_30811,N_31299);
nand U39899 (N_39899,N_34810,N_32133);
or U39900 (N_39900,N_34240,N_34604);
nand U39901 (N_39901,N_30422,N_34399);
nand U39902 (N_39902,N_31534,N_31153);
nor U39903 (N_39903,N_30569,N_30409);
or U39904 (N_39904,N_31730,N_31290);
and U39905 (N_39905,N_34416,N_32165);
and U39906 (N_39906,N_33186,N_30665);
nor U39907 (N_39907,N_31677,N_31629);
xnor U39908 (N_39908,N_33890,N_31637);
xnor U39909 (N_39909,N_31519,N_33605);
xor U39910 (N_39910,N_32922,N_32903);
xor U39911 (N_39911,N_31948,N_30490);
or U39912 (N_39912,N_33468,N_34008);
nor U39913 (N_39913,N_33676,N_34782);
nor U39914 (N_39914,N_32482,N_30843);
or U39915 (N_39915,N_32762,N_33752);
or U39916 (N_39916,N_31957,N_32318);
nand U39917 (N_39917,N_33571,N_30400);
or U39918 (N_39918,N_33485,N_30491);
xor U39919 (N_39919,N_34916,N_31611);
nand U39920 (N_39920,N_31027,N_30158);
and U39921 (N_39921,N_31381,N_30307);
nand U39922 (N_39922,N_32023,N_32394);
nor U39923 (N_39923,N_33248,N_34222);
nor U39924 (N_39924,N_32407,N_34660);
nor U39925 (N_39925,N_31907,N_33122);
nand U39926 (N_39926,N_34917,N_30905);
nand U39927 (N_39927,N_34273,N_31742);
xnor U39928 (N_39928,N_32211,N_32923);
and U39929 (N_39929,N_30286,N_34612);
xnor U39930 (N_39930,N_32769,N_32795);
nand U39931 (N_39931,N_32490,N_31612);
xor U39932 (N_39932,N_30903,N_32214);
and U39933 (N_39933,N_31479,N_31534);
xnor U39934 (N_39934,N_30046,N_33299);
and U39935 (N_39935,N_33854,N_33942);
nor U39936 (N_39936,N_30775,N_33877);
nand U39937 (N_39937,N_30279,N_31946);
and U39938 (N_39938,N_30589,N_34942);
nor U39939 (N_39939,N_32417,N_31837);
or U39940 (N_39940,N_34198,N_32358);
and U39941 (N_39941,N_30101,N_32538);
and U39942 (N_39942,N_33780,N_34686);
or U39943 (N_39943,N_33694,N_32175);
and U39944 (N_39944,N_31583,N_31265);
and U39945 (N_39945,N_30492,N_30588);
nor U39946 (N_39946,N_33530,N_33959);
nor U39947 (N_39947,N_33471,N_33127);
and U39948 (N_39948,N_33022,N_34689);
and U39949 (N_39949,N_33547,N_31784);
nand U39950 (N_39950,N_34637,N_32001);
nor U39951 (N_39951,N_31219,N_34992);
and U39952 (N_39952,N_30548,N_31894);
and U39953 (N_39953,N_34498,N_30601);
nor U39954 (N_39954,N_30056,N_32875);
nor U39955 (N_39955,N_32690,N_32549);
or U39956 (N_39956,N_30866,N_34527);
and U39957 (N_39957,N_33982,N_31866);
and U39958 (N_39958,N_32975,N_30051);
or U39959 (N_39959,N_31338,N_31420);
nor U39960 (N_39960,N_32939,N_32082);
nor U39961 (N_39961,N_31824,N_34315);
or U39962 (N_39962,N_32662,N_32056);
or U39963 (N_39963,N_30325,N_33998);
or U39964 (N_39964,N_34731,N_30610);
nand U39965 (N_39965,N_32642,N_31350);
nor U39966 (N_39966,N_30568,N_31949);
nor U39967 (N_39967,N_33439,N_33621);
nor U39968 (N_39968,N_34206,N_30031);
and U39969 (N_39969,N_30154,N_31806);
xor U39970 (N_39970,N_33480,N_31164);
nand U39971 (N_39971,N_33820,N_30625);
nand U39972 (N_39972,N_32746,N_30825);
and U39973 (N_39973,N_32414,N_33890);
and U39974 (N_39974,N_33938,N_30252);
or U39975 (N_39975,N_34758,N_34406);
nand U39976 (N_39976,N_33617,N_30106);
or U39977 (N_39977,N_31567,N_32037);
and U39978 (N_39978,N_31754,N_30958);
and U39979 (N_39979,N_33067,N_33649);
and U39980 (N_39980,N_30710,N_33636);
nor U39981 (N_39981,N_34925,N_34814);
and U39982 (N_39982,N_32178,N_31121);
nor U39983 (N_39983,N_33843,N_32141);
and U39984 (N_39984,N_32610,N_31677);
nor U39985 (N_39985,N_33495,N_34722);
and U39986 (N_39986,N_33694,N_34763);
nand U39987 (N_39987,N_32662,N_31416);
nor U39988 (N_39988,N_34759,N_33678);
nand U39989 (N_39989,N_32773,N_30674);
nor U39990 (N_39990,N_31532,N_33438);
nor U39991 (N_39991,N_30981,N_31039);
nor U39992 (N_39992,N_33558,N_33197);
and U39993 (N_39993,N_34438,N_32214);
nand U39994 (N_39994,N_31335,N_30866);
nor U39995 (N_39995,N_32325,N_34120);
nand U39996 (N_39996,N_30857,N_33420);
nor U39997 (N_39997,N_33083,N_30255);
and U39998 (N_39998,N_34660,N_33003);
or U39999 (N_39999,N_32381,N_31113);
or U40000 (N_40000,N_38959,N_35216);
xnor U40001 (N_40001,N_36392,N_35989);
and U40002 (N_40002,N_36934,N_39893);
nand U40003 (N_40003,N_36091,N_37894);
and U40004 (N_40004,N_37125,N_39872);
and U40005 (N_40005,N_37214,N_35826);
and U40006 (N_40006,N_39430,N_37994);
nand U40007 (N_40007,N_38575,N_37152);
and U40008 (N_40008,N_35528,N_35659);
or U40009 (N_40009,N_38556,N_36185);
nand U40010 (N_40010,N_35918,N_38422);
xor U40011 (N_40011,N_38479,N_35188);
nor U40012 (N_40012,N_37098,N_36378);
and U40013 (N_40013,N_39566,N_35819);
xor U40014 (N_40014,N_35408,N_35060);
nand U40015 (N_40015,N_39353,N_39839);
or U40016 (N_40016,N_36633,N_35822);
and U40017 (N_40017,N_37202,N_36207);
or U40018 (N_40018,N_36066,N_36485);
nor U40019 (N_40019,N_36894,N_37981);
and U40020 (N_40020,N_38610,N_37374);
and U40021 (N_40021,N_35633,N_39331);
nor U40022 (N_40022,N_35264,N_39482);
nor U40023 (N_40023,N_35519,N_35161);
and U40024 (N_40024,N_39514,N_35507);
xnor U40025 (N_40025,N_35075,N_38340);
and U40026 (N_40026,N_38089,N_38909);
nand U40027 (N_40027,N_38223,N_38676);
and U40028 (N_40028,N_36189,N_39373);
nor U40029 (N_40029,N_38313,N_36042);
or U40030 (N_40030,N_35547,N_38647);
nor U40031 (N_40031,N_36942,N_38664);
or U40032 (N_40032,N_35192,N_39875);
nor U40033 (N_40033,N_35213,N_38199);
and U40034 (N_40034,N_39788,N_37944);
nor U40035 (N_40035,N_36447,N_36158);
or U40036 (N_40036,N_37861,N_39238);
and U40037 (N_40037,N_38049,N_37067);
or U40038 (N_40038,N_37762,N_39794);
and U40039 (N_40039,N_38898,N_35808);
xor U40040 (N_40040,N_38881,N_38013);
or U40041 (N_40041,N_35742,N_35476);
nor U40042 (N_40042,N_37901,N_38850);
or U40043 (N_40043,N_35809,N_38969);
nand U40044 (N_40044,N_37524,N_38533);
nor U40045 (N_40045,N_39192,N_35543);
xnor U40046 (N_40046,N_38626,N_36045);
or U40047 (N_40047,N_38245,N_39120);
nor U40048 (N_40048,N_35942,N_38399);
nor U40049 (N_40049,N_38823,N_38987);
and U40050 (N_40050,N_37361,N_36260);
or U40051 (N_40051,N_39254,N_38453);
or U40052 (N_40052,N_35894,N_39079);
and U40053 (N_40053,N_35966,N_36043);
xor U40054 (N_40054,N_36967,N_39235);
xor U40055 (N_40055,N_35522,N_36885);
or U40056 (N_40056,N_39265,N_38853);
or U40057 (N_40057,N_38451,N_37069);
nor U40058 (N_40058,N_38025,N_36837);
and U40059 (N_40059,N_38239,N_36607);
or U40060 (N_40060,N_38638,N_39227);
xor U40061 (N_40061,N_39979,N_38538);
or U40062 (N_40062,N_35860,N_37784);
or U40063 (N_40063,N_35021,N_35748);
xor U40064 (N_40064,N_38941,N_38778);
nand U40065 (N_40065,N_37815,N_38773);
nor U40066 (N_40066,N_36318,N_35234);
xnor U40067 (N_40067,N_37676,N_35278);
nor U40068 (N_40068,N_37555,N_39691);
nor U40069 (N_40069,N_35365,N_36423);
nor U40070 (N_40070,N_37691,N_36245);
and U40071 (N_40071,N_35106,N_36440);
nor U40072 (N_40072,N_35975,N_36491);
nand U40073 (N_40073,N_38158,N_39093);
and U40074 (N_40074,N_39475,N_37681);
nand U40075 (N_40075,N_37454,N_38426);
nand U40076 (N_40076,N_35579,N_36896);
nand U40077 (N_40077,N_39752,N_38989);
xnor U40078 (N_40078,N_35729,N_38143);
xor U40079 (N_40079,N_37550,N_35637);
nor U40080 (N_40080,N_39707,N_37354);
and U40081 (N_40081,N_39047,N_35386);
or U40082 (N_40082,N_37551,N_39680);
and U40083 (N_40083,N_39874,N_37973);
or U40084 (N_40084,N_37032,N_39551);
nand U40085 (N_40085,N_37363,N_36156);
nor U40086 (N_40086,N_36593,N_39730);
and U40087 (N_40087,N_39908,N_35772);
nor U40088 (N_40088,N_35299,N_39134);
or U40089 (N_40089,N_35369,N_36255);
or U40090 (N_40090,N_39746,N_38719);
nand U40091 (N_40091,N_39507,N_39064);
nand U40092 (N_40092,N_36663,N_35739);
or U40093 (N_40093,N_38619,N_38901);
nor U40094 (N_40094,N_39631,N_39028);
nand U40095 (N_40095,N_38916,N_39191);
or U40096 (N_40096,N_38118,N_36925);
and U40097 (N_40097,N_37628,N_39076);
or U40098 (N_40098,N_36792,N_37824);
or U40099 (N_40099,N_38620,N_36386);
or U40100 (N_40100,N_36284,N_38282);
nand U40101 (N_40101,N_37158,N_36930);
or U40102 (N_40102,N_39630,N_39186);
xor U40103 (N_40103,N_38433,N_37780);
xor U40104 (N_40104,N_36664,N_36102);
and U40105 (N_40105,N_37892,N_39199);
or U40106 (N_40106,N_38146,N_36344);
nor U40107 (N_40107,N_37683,N_38267);
nor U40108 (N_40108,N_39768,N_35289);
nor U40109 (N_40109,N_35353,N_35727);
nor U40110 (N_40110,N_38111,N_37800);
nor U40111 (N_40111,N_36522,N_36141);
nor U40112 (N_40112,N_37739,N_36818);
and U40113 (N_40113,N_37207,N_39083);
or U40114 (N_40114,N_39796,N_37289);
nand U40115 (N_40115,N_39489,N_35864);
nand U40116 (N_40116,N_35428,N_38596);
nand U40117 (N_40117,N_35802,N_36254);
nor U40118 (N_40118,N_38600,N_37134);
xnor U40119 (N_40119,N_38960,N_35426);
nand U40120 (N_40120,N_38885,N_38504);
nand U40121 (N_40121,N_37778,N_37868);
or U40122 (N_40122,N_37234,N_36669);
nor U40123 (N_40123,N_37641,N_36501);
and U40124 (N_40124,N_35477,N_39720);
or U40125 (N_40125,N_39498,N_38684);
xor U40126 (N_40126,N_38306,N_35761);
nand U40127 (N_40127,N_37713,N_36272);
nor U40128 (N_40128,N_36907,N_35687);
nor U40129 (N_40129,N_39553,N_38861);
or U40130 (N_40130,N_39367,N_38314);
or U40131 (N_40131,N_35373,N_38474);
nand U40132 (N_40132,N_36547,N_38084);
nor U40133 (N_40133,N_36875,N_35412);
or U40134 (N_40134,N_38765,N_38424);
and U40135 (N_40135,N_37882,N_36073);
and U40136 (N_40136,N_36553,N_38331);
and U40137 (N_40137,N_37849,N_36647);
nor U40138 (N_40138,N_39665,N_35800);
or U40139 (N_40139,N_39442,N_38952);
nor U40140 (N_40140,N_36090,N_38180);
nand U40141 (N_40141,N_36036,N_39841);
and U40142 (N_40142,N_36780,N_39669);
or U40143 (N_40143,N_36484,N_35544);
or U40144 (N_40144,N_39616,N_36481);
and U40145 (N_40145,N_35974,N_36637);
nand U40146 (N_40146,N_36588,N_39488);
nor U40147 (N_40147,N_36106,N_36478);
and U40148 (N_40148,N_35804,N_37660);
and U40149 (N_40149,N_37938,N_39700);
xnor U40150 (N_40150,N_35319,N_37860);
nand U40151 (N_40151,N_35780,N_37675);
nor U40152 (N_40152,N_36829,N_37731);
nand U40153 (N_40153,N_39656,N_38445);
and U40154 (N_40154,N_35360,N_36417);
or U40155 (N_40155,N_37147,N_38269);
or U40156 (N_40156,N_39595,N_37310);
nand U40157 (N_40157,N_39762,N_35720);
and U40158 (N_40158,N_39795,N_35363);
and U40159 (N_40159,N_35602,N_37314);
nand U40160 (N_40160,N_39298,N_37949);
nand U40161 (N_40161,N_36735,N_35431);
and U40162 (N_40162,N_39922,N_35371);
nand U40163 (N_40163,N_39376,N_38648);
or U40164 (N_40164,N_38829,N_39751);
and U40165 (N_40165,N_35122,N_37372);
or U40166 (N_40166,N_38567,N_39101);
nand U40167 (N_40167,N_36049,N_39244);
nand U40168 (N_40168,N_38087,N_39487);
nor U40169 (N_40169,N_35523,N_37364);
and U40170 (N_40170,N_37790,N_38731);
or U40171 (N_40171,N_39767,N_39122);
nor U40172 (N_40172,N_36855,N_39476);
xor U40173 (N_40173,N_39842,N_39117);
and U40174 (N_40174,N_38024,N_36472);
or U40175 (N_40175,N_35596,N_36367);
and U40176 (N_40176,N_38363,N_36923);
nor U40177 (N_40177,N_35166,N_37852);
nor U40178 (N_40178,N_37276,N_39930);
or U40179 (N_40179,N_38098,N_38594);
nor U40180 (N_40180,N_37832,N_36040);
and U40181 (N_40181,N_38542,N_38982);
nor U40182 (N_40182,N_38114,N_39137);
and U40183 (N_40183,N_39995,N_39241);
and U40184 (N_40184,N_37957,N_35463);
nand U40185 (N_40185,N_35741,N_39970);
nand U40186 (N_40186,N_35823,N_39406);
nor U40187 (N_40187,N_35224,N_39902);
and U40188 (N_40188,N_39856,N_39470);
nand U40189 (N_40189,N_37560,N_39947);
nor U40190 (N_40190,N_37086,N_35597);
xnor U40191 (N_40191,N_37175,N_35328);
nor U40192 (N_40192,N_36466,N_39211);
or U40193 (N_40193,N_36198,N_39981);
or U40194 (N_40194,N_38836,N_37444);
nor U40195 (N_40195,N_38782,N_38329);
nand U40196 (N_40196,N_36031,N_38800);
nor U40197 (N_40197,N_38756,N_37963);
or U40198 (N_40198,N_36881,N_35441);
and U40199 (N_40199,N_39151,N_39890);
xnor U40200 (N_40200,N_39864,N_35517);
nor U40201 (N_40201,N_39321,N_37741);
nor U40202 (N_40202,N_37514,N_37678);
or U40203 (N_40203,N_39396,N_35711);
xnor U40204 (N_40204,N_38807,N_36502);
nor U40205 (N_40205,N_38081,N_37584);
nand U40206 (N_40206,N_39703,N_38133);
nor U40207 (N_40207,N_36789,N_37472);
and U40208 (N_40208,N_37260,N_35536);
and U40209 (N_40209,N_37288,N_37631);
and U40210 (N_40210,N_35812,N_38623);
or U40211 (N_40211,N_35880,N_39813);
or U40212 (N_40212,N_36022,N_39814);
nor U40213 (N_40213,N_37462,N_36650);
or U40214 (N_40214,N_39708,N_35691);
xnor U40215 (N_40215,N_35357,N_36579);
nand U40216 (N_40216,N_37577,N_39496);
or U40217 (N_40217,N_38689,N_39517);
nor U40218 (N_40218,N_35871,N_37103);
nand U40219 (N_40219,N_35157,N_35968);
xnor U40220 (N_40220,N_38316,N_35930);
and U40221 (N_40221,N_39757,N_39364);
nand U40222 (N_40222,N_37100,N_37877);
nor U40223 (N_40223,N_38407,N_35946);
nor U40224 (N_40224,N_38880,N_37383);
or U40225 (N_40225,N_35261,N_36528);
or U40226 (N_40226,N_39484,N_35593);
nor U40227 (N_40227,N_38152,N_37291);
nand U40228 (N_40228,N_37992,N_37888);
xnor U40229 (N_40229,N_37677,N_38931);
nand U40230 (N_40230,N_36015,N_37837);
nand U40231 (N_40231,N_38373,N_36731);
nor U40232 (N_40232,N_38443,N_37431);
xnor U40233 (N_40233,N_39977,N_39124);
nand U40234 (N_40234,N_36852,N_37858);
nor U40235 (N_40235,N_39805,N_39026);
nor U40236 (N_40236,N_36152,N_36749);
and U40237 (N_40237,N_37261,N_35086);
or U40238 (N_40238,N_35795,N_36027);
nor U40239 (N_40239,N_39045,N_36068);
nor U40240 (N_40240,N_36455,N_37149);
nor U40241 (N_40241,N_38312,N_39810);
xnor U40242 (N_40242,N_35097,N_39409);
and U40243 (N_40243,N_39775,N_37110);
nand U40244 (N_40244,N_35151,N_37269);
nand U40245 (N_40245,N_35609,N_35305);
and U40246 (N_40246,N_39258,N_39088);
and U40247 (N_40247,N_37498,N_38862);
nor U40248 (N_40248,N_39637,N_35787);
and U40249 (N_40249,N_35337,N_35270);
nand U40250 (N_40250,N_35184,N_35927);
nor U40251 (N_40251,N_39268,N_39857);
nand U40252 (N_40252,N_35650,N_39415);
nor U40253 (N_40253,N_39502,N_37876);
nand U40254 (N_40254,N_36286,N_35423);
xor U40255 (N_40255,N_38318,N_38220);
or U40256 (N_40256,N_38935,N_38883);
or U40257 (N_40257,N_39649,N_37283);
or U40258 (N_40258,N_39313,N_36693);
or U40259 (N_40259,N_36586,N_36836);
nor U40260 (N_40260,N_38785,N_36083);
nor U40261 (N_40261,N_39668,N_37150);
nor U40262 (N_40262,N_39135,N_38032);
xnor U40263 (N_40263,N_39519,N_36825);
and U40264 (N_40264,N_35961,N_36571);
nand U40265 (N_40265,N_38607,N_37210);
nor U40266 (N_40266,N_37836,N_38192);
or U40267 (N_40267,N_39345,N_37557);
xnor U40268 (N_40268,N_35487,N_36161);
and U40269 (N_40269,N_37266,N_36388);
or U40270 (N_40270,N_36424,N_36011);
nor U40271 (N_40271,N_36985,N_37323);
xnor U40272 (N_40272,N_36880,N_35217);
nor U40273 (N_40273,N_35405,N_35503);
or U40274 (N_40274,N_35649,N_38819);
xnor U40275 (N_40275,N_37121,N_38795);
and U40276 (N_40276,N_37763,N_37899);
and U40277 (N_40277,N_39056,N_37567);
nand U40278 (N_40278,N_35012,N_38435);
nand U40279 (N_40279,N_36046,N_37281);
or U40280 (N_40280,N_36492,N_35280);
or U40281 (N_40281,N_39316,N_36312);
or U40282 (N_40282,N_38082,N_39674);
or U40283 (N_40283,N_35652,N_36026);
or U40284 (N_40284,N_38324,N_36389);
nand U40285 (N_40285,N_35446,N_38967);
nor U40286 (N_40286,N_39548,N_36691);
and U40287 (N_40287,N_35955,N_35838);
or U40288 (N_40288,N_35081,N_37297);
nor U40289 (N_40289,N_37966,N_36514);
or U40290 (N_40290,N_37002,N_37629);
and U40291 (N_40291,N_35469,N_38018);
and U40292 (N_40292,N_39343,N_36763);
and U40293 (N_40293,N_36464,N_38436);
xnor U40294 (N_40294,N_37176,N_35453);
nand U40295 (N_40295,N_37996,N_38546);
and U40296 (N_40296,N_39421,N_37510);
nor U40297 (N_40297,N_39765,N_36256);
nand U40298 (N_40298,N_35770,N_35035);
nand U40299 (N_40299,N_39443,N_38653);
or U40300 (N_40300,N_38992,N_36706);
or U40301 (N_40301,N_35554,N_35932);
and U40302 (N_40302,N_38745,N_37914);
nor U40303 (N_40303,N_39275,N_39295);
nand U40304 (N_40304,N_36771,N_35383);
nand U40305 (N_40305,N_35731,N_35121);
nand U40306 (N_40306,N_35817,N_36450);
nand U40307 (N_40307,N_35764,N_39040);
nor U40308 (N_40308,N_37580,N_39726);
nor U40309 (N_40309,N_36899,N_39162);
nor U40310 (N_40310,N_37169,N_36550);
nor U40311 (N_40311,N_36267,N_37268);
and U40312 (N_40312,N_39895,N_35409);
nand U40313 (N_40313,N_39289,N_36694);
or U40314 (N_40314,N_37247,N_38214);
or U40315 (N_40315,N_38516,N_38768);
nand U40316 (N_40316,N_39090,N_35185);
and U40317 (N_40317,N_38561,N_37491);
or U40318 (N_40318,N_38966,N_37620);
or U40319 (N_40319,N_38757,N_38438);
and U40320 (N_40320,N_37519,N_38256);
or U40321 (N_40321,N_35489,N_36546);
or U40322 (N_40322,N_39174,N_37051);
nor U40323 (N_40323,N_38911,N_36774);
or U40324 (N_40324,N_38636,N_35443);
nor U40325 (N_40325,N_38642,N_35972);
and U40326 (N_40326,N_37875,N_37755);
nand U40327 (N_40327,N_37165,N_39536);
or U40328 (N_40328,N_38332,N_39042);
nor U40329 (N_40329,N_37895,N_36609);
nand U40330 (N_40330,N_39339,N_35600);
or U40331 (N_40331,N_37826,N_36847);
nand U40332 (N_40332,N_38156,N_36523);
or U40333 (N_40333,N_36240,N_37467);
nor U40334 (N_40334,N_36956,N_36662);
or U40335 (N_40335,N_35840,N_36728);
and U40336 (N_40336,N_35485,N_36390);
nand U40337 (N_40337,N_39312,N_37265);
nor U40338 (N_40338,N_39449,N_38603);
nor U40339 (N_40339,N_36380,N_35775);
or U40340 (N_40340,N_36163,N_36281);
nor U40341 (N_40341,N_35726,N_39338);
or U40342 (N_40342,N_36902,N_36758);
nor U40343 (N_40343,N_37404,N_37910);
nor U40344 (N_40344,N_35994,N_38174);
xnor U40345 (N_40345,N_38617,N_37346);
and U40346 (N_40346,N_38384,N_36516);
and U40347 (N_40347,N_37828,N_38606);
or U40348 (N_40348,N_36924,N_38608);
xnor U40349 (N_40349,N_35095,N_38691);
nor U40350 (N_40350,N_38350,N_35744);
nand U40351 (N_40351,N_37878,N_36549);
or U40352 (N_40352,N_35288,N_35865);
nand U40353 (N_40353,N_36136,N_39336);
xor U40354 (N_40354,N_38184,N_37694);
nor U40355 (N_40355,N_39604,N_35866);
and U40356 (N_40356,N_38364,N_36603);
nor U40357 (N_40357,N_39713,N_39655);
nor U40358 (N_40358,N_39891,N_35624);
nand U40359 (N_40359,N_38446,N_37232);
xor U40360 (N_40360,N_39354,N_38204);
or U40361 (N_40361,N_39086,N_36870);
and U40362 (N_40362,N_36048,N_35462);
or U40363 (N_40363,N_39413,N_37639);
and U40364 (N_40364,N_36391,N_39204);
and U40365 (N_40365,N_37535,N_39769);
and U40366 (N_40366,N_38042,N_39802);
and U40367 (N_40367,N_35108,N_36080);
nor U40368 (N_40368,N_39948,N_37038);
xor U40369 (N_40369,N_39632,N_35707);
and U40370 (N_40370,N_36329,N_39946);
or U40371 (N_40371,N_39613,N_35322);
nand U40372 (N_40372,N_38609,N_37022);
xnor U40373 (N_40373,N_38587,N_36649);
xor U40374 (N_40374,N_37658,N_37880);
and U40375 (N_40375,N_37080,N_36052);
xnor U40376 (N_40376,N_35300,N_38831);
nand U40377 (N_40377,N_37495,N_38848);
or U40378 (N_40378,N_37795,N_36996);
nor U40379 (N_40379,N_39007,N_36524);
nor U40380 (N_40380,N_39207,N_35790);
nand U40381 (N_40381,N_37831,N_39742);
and U40382 (N_40382,N_35756,N_37757);
nor U40383 (N_40383,N_35259,N_35807);
or U40384 (N_40384,N_36537,N_39851);
or U40385 (N_40385,N_39821,N_38240);
nand U40386 (N_40386,N_38579,N_39942);
and U40387 (N_40387,N_35601,N_37441);
and U40388 (N_40388,N_36505,N_37968);
or U40389 (N_40389,N_36128,N_38794);
and U40390 (N_40390,N_39759,N_36319);
nor U40391 (N_40391,N_38996,N_35361);
and U40392 (N_40392,N_39296,N_39492);
and U40393 (N_40393,N_36743,N_39992);
nor U40394 (N_40394,N_39435,N_37932);
nand U40395 (N_40395,N_39299,N_37744);
or U40396 (N_40396,N_39785,N_39815);
nor U40397 (N_40397,N_35169,N_37039);
nand U40398 (N_40398,N_38251,N_35730);
or U40399 (N_40399,N_37275,N_37839);
nand U40400 (N_40400,N_37023,N_35372);
and U40401 (N_40401,N_37789,N_38733);
and U40402 (N_40402,N_36828,N_39725);
and U40403 (N_40403,N_39279,N_38914);
xor U40404 (N_40404,N_39927,N_37674);
nor U40405 (N_40405,N_38645,N_35938);
nand U40406 (N_40406,N_35675,N_39046);
nand U40407 (N_40407,N_38578,N_36846);
nand U40408 (N_40408,N_37933,N_38791);
nand U40409 (N_40409,N_36697,N_36978);
nand U40410 (N_40410,N_36293,N_35240);
nand U40411 (N_40411,N_39940,N_35530);
and U40412 (N_40412,N_37027,N_38397);
and U40413 (N_40413,N_39812,N_36224);
or U40414 (N_40414,N_36613,N_35498);
or U40415 (N_40415,N_38508,N_38727);
nand U40416 (N_40416,N_39635,N_36791);
and U40417 (N_40417,N_39285,N_35318);
nor U40418 (N_40418,N_35105,N_39879);
nand U40419 (N_40419,N_38978,N_36277);
nand U40420 (N_40420,N_37043,N_39505);
and U40421 (N_40421,N_35221,N_36113);
xnor U40422 (N_40422,N_39580,N_37410);
or U40423 (N_40423,N_38864,N_38704);
nor U40424 (N_40424,N_35951,N_38503);
nor U40425 (N_40425,N_38075,N_36279);
and U40426 (N_40426,N_35402,N_36585);
nor U40427 (N_40427,N_35954,N_38344);
and U40428 (N_40428,N_39378,N_36212);
or U40429 (N_40429,N_35123,N_35380);
and U40430 (N_40430,N_39306,N_38302);
xnor U40431 (N_40431,N_35414,N_39581);
or U40432 (N_40432,N_36414,N_36310);
nor U40433 (N_40433,N_35511,N_36801);
nor U40434 (N_40434,N_39310,N_36954);
or U40435 (N_40435,N_35212,N_36871);
nor U40436 (N_40436,N_38718,N_35018);
and U40437 (N_40437,N_39860,N_36112);
xor U40438 (N_40438,N_36013,N_39926);
nor U40439 (N_40439,N_39850,N_37753);
or U40440 (N_40440,N_39925,N_35987);
nor U40441 (N_40441,N_37217,N_35171);
or U40442 (N_40442,N_37865,N_37459);
or U40443 (N_40443,N_38492,N_35020);
xnor U40444 (N_40444,N_36038,N_37930);
nor U40445 (N_40445,N_35390,N_37195);
or U40446 (N_40446,N_38536,N_39387);
or U40447 (N_40447,N_37610,N_38437);
or U40448 (N_40448,N_36214,N_38303);
and U40449 (N_40449,N_37248,N_37871);
or U40450 (N_40450,N_38126,N_38414);
and U40451 (N_40451,N_38971,N_38040);
nor U40452 (N_40452,N_39740,N_36453);
xor U40453 (N_40453,N_36382,N_38590);
or U40454 (N_40454,N_35642,N_37326);
nand U40455 (N_40455,N_38216,N_39918);
nor U40456 (N_40456,N_36831,N_39799);
nor U40457 (N_40457,N_39834,N_35091);
nand U40458 (N_40458,N_38798,N_35066);
and U40459 (N_40459,N_35606,N_36427);
or U40460 (N_40460,N_37934,N_39542);
nor U40461 (N_40461,N_37614,N_35814);
and U40462 (N_40462,N_36953,N_38710);
nor U40463 (N_40463,N_36988,N_38213);
nor U40464 (N_40464,N_39365,N_36893);
nor U40465 (N_40465,N_37143,N_37701);
xor U40466 (N_40466,N_39508,N_39480);
and U40467 (N_40467,N_39248,N_38457);
nor U40468 (N_40468,N_37097,N_35490);
nand U40469 (N_40469,N_35896,N_36712);
or U40470 (N_40470,N_37976,N_39080);
and U40471 (N_40471,N_39518,N_35314);
nor U40472 (N_40472,N_39897,N_37652);
or U40473 (N_40473,N_38954,N_39729);
or U40474 (N_40474,N_38108,N_39096);
or U40475 (N_40475,N_36781,N_38920);
nand U40476 (N_40476,N_36658,N_37448);
nor U40477 (N_40477,N_38641,N_35702);
nor U40478 (N_40478,N_35957,N_38577);
and U40479 (N_40479,N_39699,N_39924);
nand U40480 (N_40480,N_39394,N_37338);
nand U40481 (N_40481,N_35307,N_35310);
or U40482 (N_40482,N_39390,N_35883);
nor U40483 (N_40483,N_35613,N_39293);
or U40484 (N_40484,N_36530,N_36296);
and U40485 (N_40485,N_36599,N_39383);
or U40486 (N_40486,N_35111,N_39836);
or U40487 (N_40487,N_35899,N_35782);
xor U40488 (N_40488,N_39964,N_37743);
nand U40489 (N_40489,N_38148,N_36258);
or U40490 (N_40490,N_39642,N_39434);
xor U40491 (N_40491,N_37825,N_38060);
xnor U40492 (N_40492,N_38106,N_37405);
nor U40493 (N_40493,N_36800,N_39223);
and U40494 (N_40494,N_37402,N_38847);
and U40495 (N_40495,N_36396,N_37682);
and U40496 (N_40496,N_35368,N_38835);
nor U40497 (N_40497,N_36835,N_35771);
nand U40498 (N_40498,N_36704,N_36077);
nor U40499 (N_40499,N_39678,N_35068);
nor U40500 (N_40500,N_35258,N_35841);
and U40501 (N_40501,N_38672,N_37782);
or U40502 (N_40502,N_37345,N_38804);
nand U40503 (N_40503,N_37397,N_39522);
nor U40504 (N_40504,N_38112,N_38160);
xnor U40505 (N_40505,N_38513,N_37251);
or U40506 (N_40506,N_35906,N_39803);
nor U40507 (N_40507,N_39362,N_35175);
xor U40508 (N_40508,N_37058,N_35296);
nor U40509 (N_40509,N_38611,N_36532);
nand U40510 (N_40510,N_37943,N_35041);
nor U40511 (N_40511,N_38168,N_39176);
and U40512 (N_40512,N_36889,N_35471);
or U40513 (N_40513,N_38377,N_39737);
xnor U40514 (N_40514,N_38449,N_37615);
or U40515 (N_40515,N_39472,N_35323);
xor U40516 (N_40516,N_37257,N_39697);
and U40517 (N_40517,N_37463,N_38932);
nand U40518 (N_40518,N_38716,N_37398);
nor U40519 (N_40519,N_36909,N_36047);
or U40520 (N_40520,N_38028,N_35783);
nor U40521 (N_40521,N_35576,N_35040);
xnor U40522 (N_40522,N_35180,N_39572);
or U40523 (N_40523,N_38305,N_37357);
xor U40524 (N_40524,N_36122,N_37856);
or U40525 (N_40525,N_36186,N_37096);
nand U40526 (N_40526,N_37919,N_35153);
nand U40527 (N_40527,N_35287,N_38279);
nor U40528 (N_40528,N_38855,N_36145);
xor U40529 (N_40529,N_37982,N_39952);
nand U40530 (N_40530,N_35705,N_37295);
nand U40531 (N_40531,N_36057,N_37474);
or U40532 (N_40532,N_38128,N_39690);
or U40533 (N_40533,N_35312,N_39727);
xor U40534 (N_40534,N_37679,N_36111);
nor U40535 (N_40535,N_38588,N_39956);
nand U40536 (N_40536,N_39104,N_36108);
or U40537 (N_40537,N_39395,N_36220);
nor U40538 (N_40538,N_35885,N_36217);
nand U40539 (N_40539,N_38809,N_39242);
nor U40540 (N_40540,N_36583,N_35847);
nand U40541 (N_40541,N_38663,N_35201);
nor U40542 (N_40542,N_38442,N_35445);
nor U40543 (N_40543,N_39847,N_37633);
nor U40544 (N_40544,N_35129,N_39670);
nand U40545 (N_40545,N_37191,N_37813);
nand U40546 (N_40546,N_38917,N_37341);
and U40547 (N_40547,N_39753,N_35862);
and U40548 (N_40548,N_39032,N_37965);
nor U40549 (N_40549,N_36263,N_37686);
or U40550 (N_40550,N_38390,N_37571);
nor U40551 (N_40551,N_39526,N_39676);
or U40552 (N_40552,N_37370,N_36467);
or U40553 (N_40553,N_38092,N_38006);
and U40554 (N_40554,N_35223,N_35695);
nand U40555 (N_40555,N_38002,N_38758);
nor U40556 (N_40556,N_39358,N_38886);
xnor U40557 (N_40557,N_39315,N_36342);
or U40558 (N_40558,N_37174,N_35575);
nand U40559 (N_40559,N_39951,N_38968);
or U40560 (N_40560,N_37016,N_37168);
or U40561 (N_40561,N_35416,N_36572);
xnor U40562 (N_40562,N_37814,N_39084);
or U40563 (N_40563,N_36420,N_38764);
and U40564 (N_40564,N_35411,N_37779);
xor U40565 (N_40565,N_38651,N_36708);
and U40566 (N_40566,N_37812,N_35252);
nand U40567 (N_40567,N_37887,N_37416);
nor U40568 (N_40568,N_35191,N_38463);
and U40569 (N_40569,N_36208,N_36683);
or U40570 (N_40570,N_37235,N_36479);
nand U40571 (N_40571,N_36023,N_37319);
or U40572 (N_40572,N_37126,N_39171);
xnor U40573 (N_40573,N_38991,N_35450);
or U40574 (N_40574,N_39706,N_35331);
nand U40575 (N_40575,N_38134,N_38685);
nor U40576 (N_40576,N_38391,N_38097);
and U40577 (N_40577,N_35850,N_37500);
xor U40578 (N_40578,N_37767,N_37504);
or U40579 (N_40579,N_38080,N_38145);
or U40580 (N_40580,N_35879,N_39214);
or U40581 (N_40581,N_38193,N_37451);
nor U40582 (N_40582,N_39679,N_35359);
nor U40583 (N_40583,N_37029,N_36716);
xnor U40584 (N_40584,N_38510,N_36237);
and U40585 (N_40585,N_39511,N_38372);
or U40586 (N_40586,N_35062,N_38613);
and U40587 (N_40587,N_36715,N_38633);
or U40588 (N_40588,N_35480,N_36710);
and U40589 (N_40589,N_38181,N_36248);
nand U40590 (N_40590,N_37138,N_39590);
nand U40591 (N_40591,N_37026,N_37017);
nand U40592 (N_40592,N_35214,N_36616);
nor U40593 (N_40593,N_35952,N_36443);
nand U40594 (N_40594,N_35902,N_36269);
nor U40595 (N_40595,N_37854,N_39535);
or U40596 (N_40596,N_38345,N_35639);
nor U40597 (N_40597,N_35566,N_36620);
or U40598 (N_40598,N_39340,N_37485);
xor U40599 (N_40599,N_39239,N_37104);
and U40600 (N_40600,N_37187,N_35492);
nand U40601 (N_40601,N_36654,N_36352);
xor U40602 (N_40602,N_39054,N_38368);
and U40603 (N_40603,N_36575,N_38657);
xnor U40604 (N_40604,N_35688,N_36543);
and U40605 (N_40605,N_37237,N_37351);
and U40606 (N_40606,N_36840,N_36150);
and U40607 (N_40607,N_37718,N_36720);
or U40608 (N_40608,N_38544,N_36734);
xor U40609 (N_40609,N_36184,N_39441);
nand U40610 (N_40610,N_39579,N_36025);
nand U40611 (N_40611,N_39377,N_38673);
xor U40612 (N_40612,N_37585,N_37705);
nor U40613 (N_40613,N_39361,N_37563);
nor U40614 (N_40614,N_37386,N_37349);
nand U40615 (N_40615,N_36465,N_36615);
or U40616 (N_40616,N_39436,N_37642);
nor U40617 (N_40617,N_37458,N_39463);
or U40618 (N_40618,N_36307,N_39460);
nand U40619 (N_40619,N_39292,N_35324);
nor U40620 (N_40620,N_37381,N_35749);
and U40621 (N_40621,N_37964,N_36937);
nand U40622 (N_40622,N_39932,N_39352);
and U40623 (N_40623,N_37624,N_36813);
or U40624 (N_40624,N_38473,N_39622);
xnor U40625 (N_40625,N_36331,N_35366);
nand U40626 (N_40626,N_36673,N_39069);
nor U40627 (N_40627,N_35953,N_36685);
nor U40628 (N_40628,N_35126,N_36273);
nor U40629 (N_40629,N_35257,N_35071);
nand U40630 (N_40630,N_37130,N_37801);
or U40631 (N_40631,N_38360,N_36278);
or U40632 (N_40632,N_37011,N_35512);
nor U40633 (N_40633,N_35612,N_38851);
nor U40634 (N_40634,N_35199,N_35589);
nand U40635 (N_40635,N_37533,N_35125);
and U40636 (N_40636,N_35851,N_35005);
xnor U40637 (N_40637,N_38668,N_38859);
or U40638 (N_40638,N_37603,N_39324);
nor U40639 (N_40639,N_37487,N_36508);
nand U40640 (N_40640,N_36103,N_36919);
nor U40641 (N_40641,N_39305,N_39625);
nand U40642 (N_40642,N_39557,N_35120);
and U40643 (N_40643,N_36943,N_37294);
nand U40644 (N_40644,N_38792,N_36518);
and U40645 (N_40645,N_37576,N_39272);
nand U40646 (N_40646,N_35664,N_38170);
nor U40647 (N_40647,N_36655,N_35344);
nand U40648 (N_40648,N_39658,N_35759);
or U40649 (N_40649,N_38321,N_36004);
nor U40650 (N_40650,N_37700,N_39587);
and U40651 (N_40651,N_38121,N_37630);
or U40652 (N_40652,N_36920,N_39705);
xnor U40653 (N_40653,N_37970,N_38053);
nor U40654 (N_40654,N_37623,N_35648);
nand U40655 (N_40655,N_39861,N_36936);
nor U40656 (N_40656,N_37884,N_37324);
nor U40657 (N_40657,N_38076,N_38852);
and U40658 (N_40658,N_36489,N_37714);
and U40659 (N_40659,N_35784,N_39116);
or U40660 (N_40660,N_39866,N_36994);
nor U40661 (N_40661,N_38631,N_39827);
nand U40662 (N_40662,N_39611,N_38871);
nand U40663 (N_40663,N_38994,N_38929);
or U40664 (N_40664,N_35497,N_35430);
and U40665 (N_40665,N_35218,N_39662);
nand U40666 (N_40666,N_38905,N_37863);
nand U40667 (N_40667,N_37254,N_39848);
nand U40668 (N_40668,N_37131,N_39044);
and U40669 (N_40669,N_39816,N_35417);
nor U40670 (N_40670,N_37516,N_39183);
nand U40671 (N_40671,N_38573,N_39963);
and U40672 (N_40672,N_38560,N_39327);
or U40673 (N_40673,N_36159,N_36573);
and U40674 (N_40674,N_36499,N_37118);
and U40675 (N_40675,N_39002,N_38566);
nand U40676 (N_40676,N_36730,N_37547);
nand U40677 (N_40677,N_38278,N_38274);
xnor U40678 (N_40678,N_39754,N_36702);
nor U40679 (N_40679,N_38964,N_36180);
nor U40680 (N_40680,N_37243,N_38827);
and U40681 (N_40681,N_35070,N_36853);
nand U40682 (N_40682,N_38188,N_38257);
nor U40683 (N_40683,N_38292,N_36927);
or U40684 (N_40684,N_35719,N_36640);
and U40685 (N_40685,N_35341,N_38484);
or U40686 (N_40686,N_39433,N_39202);
or U40687 (N_40687,N_37634,N_36033);
and U40688 (N_40688,N_37922,N_36449);
nor U40689 (N_40689,N_36117,N_38925);
nand U40690 (N_40690,N_36678,N_35605);
nor U40691 (N_40691,N_38333,N_37394);
nor U40692 (N_40692,N_35194,N_36299);
or U40693 (N_40693,N_37851,N_38388);
nor U40694 (N_40694,N_38317,N_38173);
and U40695 (N_40695,N_35141,N_37435);
and U40696 (N_40696,N_35542,N_39119);
or U40697 (N_40697,N_39741,N_35072);
or U40698 (N_40698,N_35569,N_39500);
and U40699 (N_40699,N_35713,N_39545);
nand U40700 (N_40700,N_35124,N_38103);
xnor U40701 (N_40701,N_38334,N_35558);
or U40702 (N_40702,N_38614,N_36174);
or U40703 (N_40703,N_36736,N_39224);
nor U40704 (N_40704,N_38205,N_36291);
nor U40705 (N_40705,N_35834,N_39000);
and U40706 (N_40706,N_38824,N_36604);
nor U40707 (N_40707,N_39177,N_39068);
or U40708 (N_40708,N_37137,N_38409);
nor U40709 (N_40709,N_37482,N_39247);
and U40710 (N_40710,N_37241,N_36775);
or U40711 (N_40711,N_35911,N_35346);
nand U40712 (N_40712,N_38039,N_36699);
and U40713 (N_40713,N_38299,N_37956);
and U40714 (N_40714,N_38742,N_37783);
or U40715 (N_40715,N_38654,N_36241);
nor U40716 (N_40716,N_39123,N_37358);
or U40717 (N_40717,N_39182,N_39477);
and U40718 (N_40718,N_37332,N_37479);
and U40719 (N_40719,N_36236,N_39121);
nor U40720 (N_40720,N_37913,N_39618);
nand U40721 (N_40721,N_36938,N_36000);
and U40722 (N_40722,N_36581,N_35116);
nor U40723 (N_40723,N_35007,N_37937);
nand U40724 (N_40724,N_37244,N_37589);
nor U40725 (N_40725,N_38601,N_38309);
or U40726 (N_40726,N_36535,N_39871);
nor U40727 (N_40727,N_39055,N_39546);
or U40728 (N_40728,N_37649,N_39138);
and U40729 (N_40729,N_39983,N_39889);
or U40730 (N_40730,N_38511,N_38477);
nor U40731 (N_40731,N_36239,N_37662);
nor U40732 (N_40732,N_35545,N_35943);
nand U40733 (N_40733,N_38621,N_36428);
nand U40734 (N_40734,N_39774,N_37331);
nor U40735 (N_40735,N_36468,N_37172);
nand U40736 (N_40736,N_37651,N_37129);
and U40737 (N_40737,N_36017,N_39652);
or U40738 (N_40738,N_37393,N_35467);
or U40739 (N_40739,N_39036,N_37796);
and U40740 (N_40740,N_37553,N_36916);
nand U40741 (N_40741,N_36366,N_38666);
nor U40742 (N_40742,N_39953,N_36434);
and U40743 (N_40743,N_38945,N_36997);
or U40744 (N_40744,N_39464,N_35981);
nand U40745 (N_40745,N_37807,N_37565);
and U40746 (N_40746,N_36301,N_38690);
and U40747 (N_40747,N_38744,N_36842);
and U40748 (N_40748,N_38845,N_35617);
nand U40749 (N_40749,N_38072,N_39887);
nor U40750 (N_40750,N_37090,N_38926);
and U40751 (N_40751,N_35699,N_38688);
or U40752 (N_40752,N_38730,N_35061);
and U40753 (N_40753,N_36711,N_35367);
nand U40754 (N_40754,N_39538,N_38369);
and U40755 (N_40755,N_36404,N_35245);
nor U40756 (N_40756,N_36974,N_35815);
or U40757 (N_40757,N_39684,N_35110);
and U40758 (N_40758,N_36362,N_38490);
xor U40759 (N_40759,N_37766,N_35924);
or U40760 (N_40760,N_35375,N_37781);
nor U40761 (N_40761,N_36178,N_39798);
nor U40762 (N_40762,N_37521,N_35971);
nor U40763 (N_40763,N_37632,N_39140);
and U40764 (N_40764,N_37198,N_39143);
nor U40765 (N_40765,N_38837,N_36221);
or U40766 (N_40766,N_36600,N_36409);
nand U40767 (N_40767,N_39592,N_37666);
and U40768 (N_40768,N_38448,N_39232);
and U40769 (N_40769,N_38660,N_37046);
or U40770 (N_40770,N_37798,N_35248);
nor U40771 (N_40771,N_38022,N_37989);
nand U40772 (N_40772,N_35420,N_35557);
nand U40773 (N_40773,N_36506,N_36926);
xnor U40774 (N_40774,N_37199,N_37328);
nor U40775 (N_40775,N_37293,N_37189);
and U40776 (N_40776,N_39523,N_35019);
nor U40777 (N_40777,N_37057,N_35669);
nor U40778 (N_40778,N_39644,N_39671);
nor U40779 (N_40779,N_39414,N_36370);
or U40780 (N_40780,N_38195,N_36977);
nand U40781 (N_40781,N_39584,N_38963);
nor U40782 (N_40782,N_39284,N_36495);
nor U40783 (N_40783,N_39205,N_39901);
and U40784 (N_40784,N_39954,N_35676);
and U40785 (N_40785,N_38362,N_38464);
and U40786 (N_40786,N_38493,N_38661);
or U40787 (N_40787,N_38380,N_37136);
nand U40788 (N_40788,N_36511,N_36336);
nand U40789 (N_40789,N_38330,N_37665);
nor U40790 (N_40790,N_36486,N_37220);
nor U40791 (N_40791,N_36521,N_36540);
nor U40792 (N_40792,N_38523,N_36959);
and U40793 (N_40793,N_36280,N_35050);
or U40794 (N_40794,N_39516,N_36932);
nand U40795 (N_40795,N_36805,N_39139);
or U40796 (N_40796,N_38419,N_36576);
or U40797 (N_40797,N_38752,N_38571);
nand U40798 (N_40798,N_36149,N_39425);
nor U40799 (N_40799,N_37019,N_36628);
nand U40800 (N_40800,N_39278,N_35684);
nand U40801 (N_40801,N_38908,N_38739);
nand U40802 (N_40802,N_35553,N_39465);
nor U40803 (N_40803,N_35253,N_39155);
and U40804 (N_40804,N_35279,N_38777);
nor U40805 (N_40805,N_39854,N_35556);
and U40806 (N_40806,N_37413,N_36405);
nand U40807 (N_40807,N_37347,N_36632);
or U40808 (N_40808,N_36355,N_35578);
nand U40809 (N_40809,N_35581,N_39643);
nand U40810 (N_40810,N_37719,N_36799);
and U40811 (N_40811,N_36262,N_38270);
and U40812 (N_40812,N_39543,N_39896);
and U40813 (N_40813,N_37240,N_35127);
nand U40814 (N_40814,N_35979,N_35769);
nor U40815 (N_40815,N_39081,N_35717);
nand U40816 (N_40816,N_38531,N_35087);
nand U40817 (N_40817,N_38241,N_35660);
xor U40818 (N_40818,N_39939,N_38725);
nand U40819 (N_40819,N_37929,N_37643);
or U40820 (N_40820,N_39418,N_36298);
or U40821 (N_40821,N_36748,N_35900);
xor U40822 (N_40822,N_36591,N_39333);
nor U40823 (N_40823,N_35941,N_37337);
nor U40824 (N_40824,N_37688,N_38142);
or U40825 (N_40825,N_37752,N_39877);
nand U40826 (N_40826,N_38517,N_36552);
and U40827 (N_40827,N_37311,N_37496);
or U40828 (N_40828,N_35447,N_39931);
and U40829 (N_40829,N_35891,N_38030);
nor U40830 (N_40830,N_36175,N_38238);
nand U40831 (N_40831,N_39389,N_39921);
or U40832 (N_40832,N_39562,N_35805);
nor U40833 (N_40833,N_36442,N_36030);
nand U40834 (N_40834,N_35117,N_39153);
and U40835 (N_40835,N_39945,N_38355);
or U40836 (N_40836,N_39852,N_36788);
nor U40837 (N_40837,N_35888,N_35845);
xnor U40838 (N_40838,N_38957,N_37717);
and U40839 (N_40839,N_38656,N_35148);
or U40840 (N_40840,N_39749,N_39282);
and U40841 (N_40841,N_39873,N_38910);
or U40842 (N_40842,N_38502,N_39840);
and U40843 (N_40843,N_35114,N_38014);
nor U40844 (N_40844,N_39220,N_39392);
or U40845 (N_40845,N_39651,N_35959);
nor U40846 (N_40846,N_38748,N_36661);
nand U40847 (N_40847,N_36527,N_37200);
nor U40848 (N_40848,N_36225,N_39495);
nand U40849 (N_40849,N_39677,N_37490);
nand U40850 (N_40850,N_36821,N_39695);
xor U40851 (N_40851,N_39916,N_38583);
nor U40852 (N_40852,N_35824,N_36921);
and U40853 (N_40853,N_38033,N_35614);
or U40854 (N_40854,N_37924,N_38376);
nor U40855 (N_40855,N_38036,N_39374);
nor U40856 (N_40856,N_35832,N_39168);
nand U40857 (N_40857,N_35301,N_39403);
or U40858 (N_40858,N_39573,N_36844);
or U40859 (N_40859,N_37927,N_36983);
nor U40860 (N_40860,N_36981,N_36940);
nor U40861 (N_40861,N_39627,N_37188);
nand U40862 (N_40862,N_35861,N_35694);
and U40863 (N_40863,N_35798,N_39692);
nor U40864 (N_40864,N_37898,N_39941);
and U40865 (N_40865,N_38790,N_39899);
and U40866 (N_40866,N_38310,N_36053);
nor U40867 (N_40867,N_36877,N_36460);
and U40868 (N_40868,N_38382,N_36171);
xor U40869 (N_40869,N_35059,N_36064);
nand U40870 (N_40870,N_35303,N_37723);
or U40871 (N_40871,N_38751,N_35561);
or U40872 (N_40872,N_39898,N_37094);
nand U40873 (N_40873,N_37245,N_38628);
nor U40874 (N_40874,N_36182,N_36786);
nand U40875 (N_40875,N_35458,N_36611);
nor U40876 (N_40876,N_38291,N_35621);
and U40877 (N_40877,N_36623,N_37494);
nand U40878 (N_40878,N_38705,N_36311);
xnor U40879 (N_40879,N_37179,N_37308);
nand U40880 (N_40880,N_39571,N_37033);
xor U40881 (N_40881,N_36767,N_35483);
or U40882 (N_40882,N_37006,N_35183);
xnor U40883 (N_40883,N_36958,N_39458);
nor U40884 (N_40884,N_36228,N_35663);
and U40885 (N_40885,N_35583,N_35452);
nand U40886 (N_40886,N_39858,N_39800);
nand U40887 (N_40887,N_35565,N_39991);
nor U40888 (N_40888,N_35654,N_35472);
nor U40889 (N_40889,N_36398,N_35495);
nand U40890 (N_40890,N_38046,N_38255);
nand U40891 (N_40891,N_37664,N_37221);
nand U40892 (N_40892,N_37879,N_37548);
nand U40893 (N_40893,N_38301,N_35109);
or U40894 (N_40894,N_39074,N_38630);
nor U40895 (N_40895,N_35355,N_36384);
nor U40896 (N_40896,N_36901,N_36261);
nand U40897 (N_40897,N_39391,N_37449);
xnor U40898 (N_40898,N_35128,N_36432);
and U40899 (N_40899,N_39379,N_36249);
or U40900 (N_40900,N_37893,N_37380);
xnor U40901 (N_40901,N_39503,N_38249);
or U40902 (N_40902,N_37917,N_37285);
nor U40903 (N_40903,N_38029,N_36062);
and U40904 (N_40904,N_35836,N_39721);
xor U40905 (N_40905,N_38468,N_37670);
or U40906 (N_40906,N_37447,N_39998);
nor U40907 (N_40907,N_35976,N_39999);
nor U40908 (N_40908,N_39640,N_36177);
or U40909 (N_40909,N_35339,N_39607);
nor U40910 (N_40910,N_38946,N_37921);
and U40911 (N_40911,N_39577,N_36162);
and U40912 (N_40912,N_37471,N_36190);
or U40913 (N_40913,N_37073,N_39471);
nor U40914 (N_40914,N_36206,N_37028);
or U40915 (N_40915,N_39388,N_39359);
nand U40916 (N_40916,N_35947,N_38284);
nand U40917 (N_40917,N_35555,N_36471);
nand U40918 (N_40918,N_38415,N_38863);
or U40919 (N_40919,N_35404,N_39960);
or U40920 (N_40920,N_39666,N_38065);
nand U40921 (N_40921,N_38953,N_37301);
nand U40922 (N_40922,N_35878,N_39131);
xnor U40923 (N_40923,N_37955,N_37313);
nor U40924 (N_40924,N_36671,N_39933);
xor U40925 (N_40925,N_35439,N_36944);
or U40926 (N_40926,N_36784,N_39804);
nor U40927 (N_40927,N_37419,N_39504);
nor U40928 (N_40928,N_39038,N_38206);
nand U40929 (N_40929,N_37437,N_36753);
and U40930 (N_40930,N_36197,N_35856);
and U40931 (N_40931,N_36032,N_35776);
and U40932 (N_40932,N_38627,N_38815);
or U40933 (N_40933,N_38512,N_36863);
or U40934 (N_40934,N_38629,N_39501);
and U40935 (N_40935,N_36770,N_39843);
and U40936 (N_40936,N_36084,N_37998);
or U40937 (N_40937,N_36696,N_39407);
xnor U40938 (N_40938,N_35595,N_38017);
and U40939 (N_40939,N_39111,N_39967);
xnor U40940 (N_40940,N_37274,N_38211);
nor U40941 (N_40941,N_37999,N_38088);
and U40942 (N_40942,N_36176,N_39229);
nand U40943 (N_40943,N_37797,N_38721);
nand U40944 (N_40944,N_36069,N_39828);
nand U40945 (N_40945,N_39417,N_36050);
and U40946 (N_40946,N_36635,N_37593);
nor U40947 (N_40947,N_38677,N_38878);
nand U40948 (N_40948,N_37505,N_35571);
or U40949 (N_40949,N_38894,N_36690);
or U40950 (N_40950,N_37035,N_36827);
xor U40951 (N_40951,N_38649,N_36657);
xnor U40952 (N_40952,N_36862,N_36790);
or U40953 (N_40953,N_36473,N_35594);
nand U40954 (N_40954,N_39323,N_39831);
or U40955 (N_40955,N_36555,N_39167);
and U40956 (N_40956,N_38772,N_36688);
or U40957 (N_40957,N_35534,N_35088);
and U40958 (N_40958,N_37407,N_36793);
nand U40959 (N_40959,N_36946,N_36496);
and U40960 (N_40960,N_38937,N_38139);
nor U40961 (N_40961,N_39006,N_36723);
xnor U40962 (N_40962,N_37818,N_38095);
nand U40963 (N_40963,N_37707,N_36539);
and U40964 (N_40964,N_38010,N_37263);
nand U40965 (N_40965,N_38167,N_35580);
and U40966 (N_40966,N_37154,N_36701);
nor U40967 (N_40967,N_35048,N_36315);
and U40968 (N_40968,N_37434,N_36991);
nand U40969 (N_40969,N_37787,N_39610);
or U40970 (N_40970,N_39567,N_35083);
xor U40971 (N_40971,N_36135,N_38821);
or U40972 (N_40972,N_35723,N_36285);
and U40973 (N_40973,N_38766,N_38454);
nor U40974 (N_40974,N_39585,N_37117);
and U40975 (N_40975,N_37726,N_39540);
nor U40976 (N_40976,N_39541,N_37663);
nand U40977 (N_40977,N_38884,N_38347);
nor U40978 (N_40978,N_35628,N_35820);
nor U40979 (N_40979,N_35884,N_39957);
nor U40980 (N_40980,N_39369,N_37095);
nand U40981 (N_40981,N_38229,N_35740);
and U40982 (N_40982,N_38965,N_35585);
and U40983 (N_40983,N_37192,N_39185);
nor U40984 (N_40984,N_39624,N_39020);
or U40985 (N_40985,N_36879,N_38670);
nand U40986 (N_40986,N_38498,N_35986);
or U40987 (N_40987,N_37945,N_39688);
nor U40988 (N_40988,N_36265,N_38045);
nor U40989 (N_40989,N_35058,N_35317);
and U40990 (N_40990,N_35309,N_36727);
and U40991 (N_40991,N_35249,N_37874);
or U40992 (N_40992,N_38394,N_39029);
or U40993 (N_40993,N_36074,N_37503);
and U40994 (N_40994,N_38995,N_39048);
or U40995 (N_40995,N_35459,N_38869);
nor U40996 (N_40996,N_39600,N_38337);
or U40997 (N_40997,N_36947,N_39178);
or U40998 (N_40998,N_37190,N_38392);
or U40999 (N_40999,N_37193,N_35196);
and U41000 (N_41000,N_39491,N_35389);
nand U41001 (N_41001,N_37208,N_39267);
and U41002 (N_41002,N_36143,N_36962);
and U41003 (N_41003,N_38485,N_35326);
nand U41004 (N_41004,N_35672,N_39989);
or U41005 (N_41005,N_37306,N_38393);
or U41006 (N_41006,N_38728,N_38051);
and U41007 (N_41007,N_38122,N_38734);
xnor U41008 (N_41008,N_35516,N_39467);
nor U41009 (N_41009,N_38326,N_38085);
or U41010 (N_41010,N_39308,N_36477);
nand U41011 (N_41011,N_37520,N_39445);
nor U41012 (N_41012,N_39129,N_36322);
nand U41013 (N_41013,N_38421,N_36915);
nor U41014 (N_41014,N_36952,N_36761);
or U41015 (N_41015,N_39330,N_39719);
and U41016 (N_41016,N_36126,N_36079);
nor U41017 (N_41017,N_39075,N_36019);
or U41018 (N_41018,N_36638,N_37935);
nand U41019 (N_41019,N_38528,N_36202);
and U41020 (N_41020,N_39335,N_37408);
or U41021 (N_41021,N_39823,N_36497);
nand U41022 (N_41022,N_38325,N_38254);
and U41023 (N_41023,N_36339,N_38135);
nor U41024 (N_41024,N_38408,N_36294);
nand U41025 (N_41025,N_39619,N_36563);
nand U41026 (N_41026,N_38527,N_39773);
and U41027 (N_41027,N_37157,N_39058);
nand U41028 (N_41028,N_38736,N_38563);
nand U41029 (N_41029,N_36383,N_39423);
or U41030 (N_41030,N_37151,N_37116);
or U41031 (N_41031,N_37259,N_35665);
nor U41032 (N_41032,N_37991,N_39118);
or U41033 (N_41033,N_36592,N_35520);
nor U41034 (N_41034,N_38323,N_38342);
or U41035 (N_41035,N_38781,N_35225);
or U41036 (N_41036,N_39304,N_36333);
nand U41037 (N_41037,N_36105,N_35488);
or U41038 (N_41038,N_37912,N_35848);
or U41039 (N_41039,N_35432,N_37915);
xor U41040 (N_41040,N_36933,N_36369);
nor U41041 (N_41041,N_39334,N_35235);
or U41042 (N_41042,N_35159,N_35304);
and U41043 (N_41043,N_38525,N_37286);
nor U41044 (N_41044,N_38161,N_36804);
xnor U41045 (N_41045,N_39984,N_37616);
nand U41046 (N_41046,N_39100,N_39092);
or U41047 (N_41047,N_39682,N_37853);
nor U41048 (N_41048,N_36574,N_36076);
and U41049 (N_41049,N_38250,N_35944);
nand U41050 (N_41050,N_37415,N_35623);
and U41051 (N_41051,N_37277,N_35236);
and U41052 (N_41052,N_39621,N_35031);
nand U41053 (N_41053,N_36705,N_39975);
nor U41054 (N_41054,N_35067,N_39822);
nor U41055 (N_41055,N_38172,N_36283);
nor U41056 (N_41056,N_35616,N_35002);
nor U41057 (N_41057,N_39574,N_39937);
nor U41058 (N_41058,N_36114,N_39510);
and U41059 (N_41059,N_39888,N_38225);
nor U41060 (N_41060,N_37350,N_38359);
xor U41061 (N_41061,N_38972,N_37379);
nand U41062 (N_41062,N_36410,N_39019);
and U41063 (N_41063,N_38452,N_38947);
or U41064 (N_41064,N_39094,N_35973);
nor U41065 (N_41065,N_36153,N_36173);
or U41066 (N_41066,N_36971,N_37489);
xor U41067 (N_41067,N_39231,N_36890);
nor U41068 (N_41068,N_37599,N_37751);
nor U41069 (N_41069,N_35905,N_38644);
and U41070 (N_41070,N_39252,N_35158);
or U41071 (N_41071,N_39602,N_36822);
and U41072 (N_41072,N_37442,N_39763);
nor U41073 (N_41073,N_35827,N_39943);
xor U41074 (N_41074,N_37083,N_35098);
nand U41075 (N_41075,N_37897,N_38023);
and U41076 (N_41076,N_38540,N_36922);
nor U41077 (N_41077,N_38506,N_37845);
xnor U41078 (N_41078,N_39870,N_36989);
nand U41079 (N_41079,N_36129,N_35008);
or U41080 (N_41080,N_38882,N_39071);
xnor U41081 (N_41081,N_37145,N_36812);
nor U41082 (N_41082,N_39807,N_39416);
nand U41083 (N_41083,N_39408,N_38434);
nor U41084 (N_41084,N_38153,N_35907);
nor U41085 (N_41085,N_35229,N_37703);
nand U41086 (N_41086,N_38547,N_39057);
nand U41087 (N_41087,N_36618,N_35256);
nor U41088 (N_41088,N_39761,N_35306);
and U41089 (N_41089,N_39809,N_35000);
nand U41090 (N_41090,N_36542,N_36714);
nor U41091 (N_41091,N_39030,N_39133);
nor U41092 (N_41092,N_38810,N_39290);
nor U41093 (N_41093,N_37012,N_38375);
nor U41094 (N_41094,N_38235,N_38828);
and U41095 (N_41095,N_39286,N_36012);
nor U41096 (N_41096,N_35718,N_38311);
and U41097 (N_41097,N_38906,N_36289);
nor U41098 (N_41098,N_36276,N_39370);
and U41099 (N_41099,N_36503,N_36006);
xnor U41100 (N_41100,N_38470,N_36107);
or U41101 (N_41101,N_36809,N_36970);
nor U41102 (N_41102,N_35433,N_37369);
nor U41103 (N_41103,N_37075,N_39328);
nand U41104 (N_41104,N_39127,N_36226);
nand U41105 (N_41105,N_37788,N_36984);
nand U41106 (N_41106,N_37460,N_38100);
and U41107 (N_41107,N_36349,N_38543);
and U41108 (N_41108,N_37153,N_35242);
nand U41109 (N_41109,N_37445,N_37322);
or U41110 (N_41110,N_37842,N_35644);
or U41111 (N_41111,N_39326,N_39758);
nand U41112 (N_41112,N_36762,N_36651);
or U41113 (N_41113,N_39172,N_37750);
and U41114 (N_41114,N_37765,N_36724);
nand U41115 (N_41115,N_37059,N_36334);
nor U41116 (N_41116,N_39620,N_39366);
or U41117 (N_41117,N_38488,N_37436);
or U41118 (N_41118,N_39696,N_39966);
nor U41119 (N_41119,N_37340,N_38413);
xnor U41120 (N_41120,N_35364,N_38120);
and U41121 (N_41121,N_36659,N_35667);
xnor U41122 (N_41122,N_39216,N_39654);
xor U41123 (N_41123,N_35403,N_39011);
nor U41124 (N_41124,N_39145,N_38811);
nor U41125 (N_41125,N_35570,N_38260);
nand U41126 (N_41126,N_35237,N_38482);
nand U41127 (N_41127,N_37053,N_36500);
and U41128 (N_41128,N_36475,N_39859);
nor U41129 (N_41129,N_38090,N_39556);
or U41130 (N_41130,N_37469,N_37960);
xnor U41131 (N_41131,N_39780,N_39494);
or U41132 (N_41132,N_35577,N_37468);
and U41133 (N_41133,N_35484,N_37684);
xor U41134 (N_41134,N_35267,N_35103);
and U41135 (N_41135,N_37473,N_36679);
and U41136 (N_41136,N_37906,N_39351);
nor U41137 (N_41137,N_36760,N_39694);
xnor U41138 (N_41138,N_39073,N_37532);
and U41139 (N_41139,N_35527,N_38052);
or U41140 (N_41140,N_35662,N_39237);
and U41141 (N_41141,N_36218,N_39043);
nor U41142 (N_41142,N_36732,N_35997);
nor U41143 (N_41143,N_39716,N_36807);
or U41144 (N_41144,N_36435,N_39400);
nand U41145 (N_41145,N_38104,N_37673);
and U41146 (N_41146,N_36230,N_36700);
or U41147 (N_41147,N_35022,N_38456);
or U41148 (N_41148,N_37010,N_35033);
nand U41149 (N_41149,N_35228,N_36359);
nand U41150 (N_41150,N_35338,N_38872);
nand U41151 (N_41151,N_35277,N_39468);
and U41152 (N_41152,N_36148,N_35853);
nor U41153 (N_41153,N_38740,N_39004);
nor U41154 (N_41154,N_35268,N_35419);
or U41155 (N_41155,N_39382,N_36610);
nor U41156 (N_41156,N_37926,N_38592);
and U41157 (N_41157,N_38044,N_37591);
and U41158 (N_41158,N_35290,N_35982);
xor U41159 (N_41159,N_35524,N_37773);
nand U41160 (N_41160,N_35643,N_37508);
nor U41161 (N_41161,N_39009,N_37049);
xor U41162 (N_41162,N_37119,N_38417);
or U41163 (N_41163,N_37786,N_39512);
or U41164 (N_41164,N_37792,N_38812);
nor U41165 (N_41165,N_35708,N_38521);
or U41166 (N_41166,N_37296,N_37911);
or U41167 (N_41167,N_39537,N_39776);
and U41168 (N_41168,N_38597,N_39027);
nand U41169 (N_41169,N_37544,N_39077);
and U41170 (N_41170,N_38921,N_37690);
nor U41171 (N_41171,N_39169,N_39024);
nor U41172 (N_41172,N_35939,N_35767);
nor U41173 (N_41173,N_39917,N_36935);
and U41174 (N_41174,N_39698,N_37771);
xor U41175 (N_41175,N_36381,N_36785);
nand U41176 (N_41176,N_37228,N_38956);
nand U41177 (N_41177,N_38598,N_36680);
and U41178 (N_41178,N_39012,N_37432);
nand U41179 (N_41179,N_37114,N_38057);
and U41180 (N_41180,N_39087,N_36729);
and U41181 (N_41181,N_35978,N_39950);
and U41182 (N_41182,N_38796,N_37425);
nor U41183 (N_41183,N_36347,N_37931);
nand U41184 (N_41184,N_37648,N_35753);
or U41185 (N_41185,N_36725,N_38865);
and U41186 (N_41186,N_37905,N_35292);
nor U41187 (N_41187,N_38450,N_35200);
xor U41188 (N_41188,N_36121,N_35077);
xor U41189 (N_41189,N_39319,N_37578);
nor U41190 (N_41190,N_37061,N_39189);
nand U41191 (N_41191,N_38753,N_39156);
or U41192 (N_41192,N_38074,N_36504);
xor U41193 (N_41193,N_37566,N_38858);
and U41194 (N_41194,N_35308,N_37209);
and U41195 (N_41195,N_39082,N_39910);
or U41196 (N_41196,N_38643,N_35284);
nor U41197 (N_41197,N_36619,N_35173);
or U41198 (N_41198,N_37602,N_39778);
nand U41199 (N_41199,N_37627,N_38553);
or U41200 (N_41200,N_35870,N_36887);
or U41201 (N_41201,N_37492,N_36797);
nand U41202 (N_41202,N_36086,N_35043);
nor U41203 (N_41203,N_37162,N_35564);
or U41204 (N_41204,N_35281,N_36098);
nand U41205 (N_41205,N_35438,N_38574);
or U41206 (N_41206,N_37048,N_38154);
and U41207 (N_41207,N_36982,N_36193);
and U41208 (N_41208,N_38061,N_39249);
nand U41209 (N_41209,N_36764,N_35745);
or U41210 (N_41210,N_38487,N_38034);
and U41211 (N_41211,N_38681,N_36843);
or U41212 (N_41212,N_35434,N_37352);
nand U41213 (N_41213,N_36323,N_39878);
and U41214 (N_41214,N_39781,N_36726);
xnor U41215 (N_41215,N_37111,N_35552);
and U41216 (N_41216,N_35980,N_37820);
or U41217 (N_41217,N_39225,N_39246);
xor U41218 (N_41218,N_37389,N_38217);
nor U41219 (N_41219,N_35653,N_38655);
nor U41220 (N_41220,N_39808,N_37984);
and U41221 (N_41221,N_36987,N_39660);
nand U41222 (N_41222,N_35873,N_39318);
and U41223 (N_41223,N_35189,N_37476);
nand U41224 (N_41224,N_39438,N_36247);
xor U41225 (N_41225,N_39212,N_37900);
nor U41226 (N_41226,N_37708,N_38750);
and U41227 (N_41227,N_37205,N_37791);
nor U41228 (N_41228,N_39314,N_35320);
nand U41229 (N_41229,N_38233,N_39337);
and U41230 (N_41230,N_37418,N_38541);
or U41231 (N_41231,N_38754,N_37528);
nor U41232 (N_41232,N_38938,N_36063);
nand U41233 (N_41233,N_36695,N_36216);
nand U41234 (N_41234,N_39280,N_39201);
or U41235 (N_41235,N_39401,N_39219);
and U41236 (N_41236,N_35716,N_39163);
and U41237 (N_41237,N_39673,N_39735);
or U41238 (N_41238,N_35882,N_38702);
xor U41239 (N_41239,N_38041,N_35743);
nand U41240 (N_41240,N_39283,N_36394);
nand U41241 (N_41241,N_35877,N_36259);
and U41242 (N_41242,N_36598,N_37107);
and U41243 (N_41243,N_37348,N_37716);
nand U41244 (N_41244,N_38162,N_37847);
nor U41245 (N_41245,N_35514,N_37805);
nand U41246 (N_41246,N_38021,N_35962);
nor U41247 (N_41247,N_39107,N_36099);
nand U41248 (N_41248,N_38780,N_35297);
nor U41249 (N_41249,N_35101,N_35329);
and U41250 (N_41250,N_39789,N_37227);
nand U41251 (N_41251,N_36782,N_36884);
nand U41252 (N_41252,N_38073,N_35929);
or U41253 (N_41253,N_38817,N_39320);
nand U41254 (N_41254,N_35397,N_38675);
or U41255 (N_41255,N_38441,N_36028);
nor U41256 (N_41256,N_37902,N_39886);
nor U41257 (N_41257,N_39944,N_37769);
nand U41258 (N_41258,N_36709,N_35921);
and U41259 (N_41259,N_36578,N_37339);
or U41260 (N_41260,N_35294,N_38524);
or U41261 (N_41261,N_39355,N_38059);
and U41262 (N_41262,N_38366,N_35010);
nand U41263 (N_41263,N_37873,N_36002);
xor U41264 (N_41264,N_37139,N_36139);
or U41265 (N_41265,N_37292,N_35890);
and U41266 (N_41266,N_37680,N_37948);
and U41267 (N_41267,N_38056,N_38447);
xnor U41268 (N_41268,N_36094,N_37671);
or U41269 (N_41269,N_37712,N_35811);
or U41270 (N_41270,N_38770,N_39663);
and U41271 (N_41271,N_35794,N_38634);
nand U41272 (N_41272,N_35038,N_36519);
or U41273 (N_41273,N_35069,N_37570);
nand U41274 (N_41274,N_36308,N_37222);
nand U41275 (N_41275,N_37600,N_35629);
and U41276 (N_41276,N_39603,N_36430);
and U41277 (N_41277,N_37271,N_36668);
nand U41278 (N_41278,N_39451,N_36510);
or U41279 (N_41279,N_39181,N_37908);
and U41280 (N_41280,N_37396,N_37645);
nor U41281 (N_41281,N_38298,N_39833);
nand U41282 (N_41282,N_35732,N_35026);
and U41283 (N_41283,N_36856,N_37334);
xnor U41284 (N_41284,N_39490,N_38379);
and U41285 (N_41285,N_38833,N_37034);
nand U41286 (N_41286,N_35250,N_37376);
and U41287 (N_41287,N_35525,N_35521);
or U41288 (N_41288,N_36061,N_38197);
and U41289 (N_41289,N_39817,N_35064);
nor U41290 (N_41290,N_38396,N_35327);
and U41291 (N_41291,N_35003,N_36144);
xor U41292 (N_41292,N_35230,N_36656);
nand U41293 (N_41293,N_39968,N_38077);
or U41294 (N_41294,N_37303,N_38808);
nor U41295 (N_41295,N_37513,N_35752);
nand U41296 (N_41296,N_39360,N_39136);
and U41297 (N_41297,N_35275,N_36350);
xnor U41298 (N_41298,N_36713,N_37692);
nand U41299 (N_41299,N_39935,N_36385);
nor U41300 (N_41300,N_38746,N_35546);
or U41301 (N_41301,N_35150,N_39257);
or U41302 (N_41302,N_39732,N_37066);
and U41303 (N_41303,N_38867,N_36097);
nor U41304 (N_41304,N_37087,N_37047);
or U41305 (N_41305,N_39148,N_36850);
nand U41306 (N_41306,N_37526,N_37020);
and U41307 (N_41307,N_37366,N_39787);
nor U41308 (N_41308,N_37164,N_36857);
or U41309 (N_41309,N_38263,N_36582);
xnor U41310 (N_41310,N_37365,N_39715);
and U41311 (N_41311,N_38799,N_36358);
nor U41312 (N_41312,N_39641,N_38079);
nor U41313 (N_41313,N_39576,N_37776);
nor U41314 (N_41314,N_35170,N_37141);
xnor U41315 (N_41315,N_39256,N_38896);
nand U41316 (N_41316,N_39997,N_35155);
or U41317 (N_41317,N_35115,N_39906);
or U41318 (N_41318,N_35674,N_35204);
and U41319 (N_41319,N_36456,N_38475);
nor U41320 (N_41320,N_35913,N_38501);
nor U41321 (N_41321,N_35145,N_35241);
and U41322 (N_41322,N_35774,N_39255);
or U41323 (N_41323,N_36639,N_39209);
or U41324 (N_41324,N_35276,N_39428);
or U41325 (N_41325,N_38296,N_37637);
nor U41326 (N_41326,N_37605,N_36703);
xor U41327 (N_41327,N_39014,N_37777);
nor U41328 (N_41328,N_38069,N_35271);
or U41329 (N_41329,N_38054,N_35825);
and U41330 (N_41330,N_35671,N_38550);
nor U41331 (N_41331,N_35313,N_36980);
and U41332 (N_41332,N_38715,N_38646);
or U41333 (N_41333,N_35945,N_38186);
nor U41334 (N_41334,N_35142,N_38897);
nand U41335 (N_41335,N_35990,N_39687);
nand U41336 (N_41336,N_35140,N_38465);
nand U41337 (N_41337,N_37054,N_35786);
nor U41338 (N_41338,N_38555,N_35136);
and U41339 (N_41339,N_35017,N_37725);
and U41340 (N_41340,N_38755,N_36913);
and U41341 (N_41341,N_35162,N_36067);
and U41342 (N_41342,N_37799,N_36911);
and U41343 (N_41343,N_35168,N_39865);
or U41344 (N_41344,N_39144,N_35889);
and U41345 (N_41345,N_37159,N_38343);
and U41346 (N_41346,N_36231,N_37406);
nand U41347 (N_41347,N_39869,N_36905);
or U41348 (N_41348,N_38237,N_39971);
nand U41349 (N_41349,N_37300,N_39835);
or U41350 (N_41350,N_35548,N_35685);
and U41351 (N_41351,N_35146,N_37273);
or U41352 (N_41352,N_35384,N_36839);
nand U41353 (N_41353,N_38942,N_35231);
or U41354 (N_41354,N_37811,N_38356);
xnor U41355 (N_41355,N_38287,N_39018);
and U41356 (N_41356,N_37160,N_37025);
xor U41357 (N_41357,N_38680,N_36439);
or U41358 (N_41358,N_38683,N_35949);
or U41359 (N_41359,N_39882,N_37573);
and U41360 (N_41360,N_38349,N_36431);
or U41361 (N_41361,N_35988,N_37647);
nor U41362 (N_41362,N_39001,N_38904);
and U41363 (N_41363,N_38389,N_36802);
or U41364 (N_41364,N_38035,N_35046);
or U41365 (N_41365,N_37253,N_39031);
nand U41366 (N_41366,N_36457,N_36667);
nor U41367 (N_41367,N_37181,N_36646);
and U41368 (N_41368,N_36556,N_37618);
nand U41369 (N_41369,N_35686,N_35567);
or U41370 (N_41370,N_38416,N_38846);
and U41371 (N_41371,N_35076,N_37401);
nand U41372 (N_41372,N_37484,N_35936);
nor U41373 (N_41373,N_36252,N_38440);
and U41374 (N_41374,N_37561,N_38275);
nor U41375 (N_41375,N_36577,N_36564);
or U41376 (N_41376,N_38591,N_35448);
nand U41377 (N_41377,N_37942,N_39880);
xor U41378 (N_41378,N_38253,N_38150);
xnor U41379 (N_41379,N_37428,N_36397);
and U41380 (N_41380,N_35917,N_38762);
nor U41381 (N_41381,N_35396,N_39628);
and U41382 (N_41382,N_37378,N_38532);
nand U41383 (N_41383,N_36219,N_37079);
or U41384 (N_41384,N_36811,N_39867);
or U41385 (N_41385,N_39586,N_37018);
nand U41386 (N_41386,N_36756,N_39397);
or U41387 (N_41387,N_36071,N_35291);
and U41388 (N_41388,N_35709,N_39262);
and U41389 (N_41389,N_37774,N_38602);
nor U41390 (N_41390,N_35285,N_38294);
and U41391 (N_41391,N_37659,N_38787);
nand U41392 (N_41392,N_37608,N_36433);
or U41393 (N_41393,N_36512,N_37722);
nand U41394 (N_41394,N_38304,N_38985);
nor U41395 (N_41395,N_36451,N_39106);
nor U41396 (N_41396,N_37746,N_35100);
or U41397 (N_41397,N_39236,N_36545);
nor U41398 (N_41398,N_39646,N_37186);
nand U41399 (N_41399,N_38993,N_37749);
xor U41400 (N_41400,N_37715,N_35455);
or U41401 (N_41401,N_37740,N_38178);
xnor U41402 (N_41402,N_39050,N_36515);
nor U41403 (N_41403,N_35636,N_37399);
nor U41404 (N_41404,N_39437,N_38699);
xor U41405 (N_41405,N_36779,N_39493);
nor U41406 (N_41406,N_35006,N_35029);
nand U41407 (N_41407,N_37867,N_38300);
xnor U41408 (N_41408,N_36740,N_37822);
and U41409 (N_41409,N_39130,N_39876);
or U41410 (N_41410,N_36297,N_37604);
or U41411 (N_41411,N_37078,N_39447);
and U41412 (N_41412,N_39597,N_39483);
nand U41413 (N_41413,N_36060,N_36868);
or U41414 (N_41414,N_37219,N_36020);
and U41415 (N_41415,N_38635,N_39617);
nor U41416 (N_41416,N_36751,N_35466);
and U41417 (N_41417,N_36309,N_37007);
nor U41418 (N_41418,N_35139,N_37185);
nand U41419 (N_41419,N_37772,N_38038);
nor U41420 (N_41420,N_37212,N_36140);
xnor U41421 (N_41421,N_35620,N_37163);
xor U41422 (N_41422,N_37833,N_37997);
or U41423 (N_41423,N_35799,N_35494);
xnor U41424 (N_41424,N_35703,N_36093);
nand U41425 (N_41425,N_38682,N_35187);
nor U41426 (N_41426,N_36343,N_38711);
or U41427 (N_41427,N_35186,N_39294);
nor U41428 (N_41428,N_38348,N_38101);
nand U41429 (N_41429,N_35478,N_39350);
nand U41430 (N_41430,N_36166,N_38462);
and U41431 (N_41431,N_39499,N_39479);
nand U41432 (N_41432,N_37060,N_36963);
and U41433 (N_41433,N_39184,N_37699);
or U41434 (N_41434,N_38055,N_39777);
or U41435 (N_41435,N_38467,N_37497);
nor U41436 (N_41436,N_35854,N_38665);
or U41437 (N_41437,N_38549,N_39782);
and U41438 (N_41438,N_38212,N_35172);
and U41439 (N_41439,N_37085,N_36151);
and U41440 (N_41440,N_36975,N_35055);
nand U41441 (N_41441,N_37305,N_35937);
nor U41442 (N_41442,N_36488,N_38230);
or U41443 (N_41443,N_36534,N_38406);
or U41444 (N_41444,N_39987,N_36059);
nor U41445 (N_41445,N_36687,N_39733);
or U41446 (N_41446,N_39633,N_39159);
or U41447 (N_41447,N_36138,N_38353);
and U41448 (N_41448,N_39766,N_39016);
or U41449 (N_41449,N_39667,N_36462);
and U41450 (N_41450,N_39955,N_37093);
xor U41451 (N_41451,N_38338,N_35781);
nand U41452 (N_41452,N_37590,N_35024);
and U41453 (N_41453,N_39037,N_39709);
nor U41454 (N_41454,N_38277,N_39114);
or U41455 (N_41455,N_37572,N_39420);
nand U41456 (N_41456,N_38564,N_37063);
or U41457 (N_41457,N_37916,N_38723);
or U41458 (N_41458,N_38551,N_38840);
or U41459 (N_41459,N_38489,N_39322);
and U41460 (N_41460,N_38123,N_36559);
or U41461 (N_41461,N_35272,N_35992);
nand U41462 (N_41462,N_38183,N_39786);
nor U41463 (N_41463,N_38866,N_39784);
and U41464 (N_41464,N_39034,N_36229);
nor U41465 (N_41465,N_38119,N_35735);
and U41466 (N_41466,N_37829,N_36009);
and U41467 (N_41467,N_39938,N_37626);
nand U41468 (N_41468,N_38252,N_39748);
xnor U41469 (N_41469,N_37480,N_35551);
or U41470 (N_41470,N_35406,N_36201);
and U41471 (N_41471,N_35931,N_35646);
nand U41472 (N_41472,N_35107,N_36242);
or U41473 (N_41473,N_39710,N_35984);
and U41474 (N_41474,N_36560,N_37466);
nand U41475 (N_41475,N_38732,N_38832);
nand U41476 (N_41476,N_37239,N_35869);
or U41477 (N_41477,N_36413,N_39385);
xnor U41478 (N_41478,N_37990,N_36165);
nor U41479 (N_41479,N_37625,N_37099);
nand U41480 (N_41480,N_39818,N_38769);
and U41481 (N_41481,N_35518,N_36051);
and U41482 (N_41482,N_35893,N_36565);
nand U41483 (N_41483,N_37734,N_36365);
or U41484 (N_41484,N_37656,N_39142);
and U41485 (N_41485,N_36860,N_38093);
nor U41486 (N_41486,N_38378,N_36796);
and U41487 (N_41487,N_38346,N_35683);
nor U41488 (N_41488,N_36429,N_36408);
nand U41489 (N_41489,N_38289,N_36235);
nor U41490 (N_41490,N_39701,N_39846);
or U41491 (N_41491,N_37077,N_38202);
xor U41492 (N_41492,N_38116,N_35473);
nand U41493 (N_41493,N_37885,N_38554);
or U41494 (N_41494,N_39147,N_37132);
nor U41495 (N_41495,N_39575,N_36001);
xor U41496 (N_41496,N_38322,N_37280);
nor U41497 (N_41497,N_36246,N_38175);
nand U41498 (N_41498,N_37538,N_39771);
and U41499 (N_41499,N_38776,N_38520);
nor U41500 (N_41500,N_36627,N_37554);
nand U41501 (N_41501,N_37636,N_39569);
or U41502 (N_41502,N_35233,N_37329);
or U41503 (N_41503,N_38849,N_36950);
and U41504 (N_41504,N_36425,N_35132);
nand U41505 (N_41505,N_35457,N_37817);
nand U41506 (N_41506,N_39988,N_36865);
nand U41507 (N_41507,N_35422,N_37233);
or U41508 (N_41508,N_37252,N_35321);
and U41509 (N_41509,N_36759,N_36474);
nand U41510 (N_41510,N_36035,N_35830);
nor U41511 (N_41511,N_39638,N_39568);
and U41512 (N_41512,N_39564,N_35211);
or U41513 (N_41513,N_36356,N_35436);
nand U41514 (N_41514,N_36999,N_36227);
or U41515 (N_41515,N_36044,N_36452);
or U41516 (N_41516,N_36324,N_39750);
nand U41517 (N_41517,N_38767,N_38398);
or U41518 (N_41518,N_36232,N_35539);
nand U41519 (N_41519,N_37993,N_35415);
and U41520 (N_41520,N_35354,N_37810);
or U41521 (N_41521,N_38749,N_36803);
xor U41522 (N_41522,N_39554,N_35451);
nor U41523 (N_41523,N_36400,N_37881);
nand U41524 (N_41524,N_36567,N_37216);
nand U41525 (N_41525,N_36003,N_39061);
and U41526 (N_41526,N_38944,N_36966);
and U41527 (N_41527,N_37733,N_37974);
nand U41528 (N_41528,N_37928,N_35014);
and U41529 (N_41529,N_39110,N_36513);
nor U41530 (N_41530,N_39961,N_39993);
and U41531 (N_41531,N_37089,N_38860);
and U41532 (N_41532,N_39598,N_37952);
nand U41533 (N_41533,N_36718,N_36878);
or U41534 (N_41534,N_36642,N_38063);
nand U41535 (N_41535,N_37242,N_38078);
nand U41536 (N_41536,N_39832,N_38522);
nand U41537 (N_41537,N_38918,N_35345);
and U41538 (N_41538,N_37422,N_35839);
or U41539 (N_41539,N_38352,N_38922);
or U41540 (N_41540,N_39170,N_37055);
nand U41541 (N_41541,N_39115,N_38802);
and U41542 (N_41542,N_38015,N_37736);
nand U41543 (N_41543,N_36589,N_35950);
and U41544 (N_41544,N_38735,N_38637);
or U41545 (N_41545,N_37834,N_35065);
nor U41546 (N_41546,N_38786,N_36014);
and U41547 (N_41547,N_37619,N_37475);
and U41548 (N_41548,N_35332,N_36133);
xnor U41549 (N_41549,N_37197,N_35311);
and U41550 (N_41550,N_36167,N_38480);
xor U41551 (N_41551,N_38692,N_37122);
nor U41552 (N_41552,N_35442,N_37421);
and U41553 (N_41553,N_36929,N_39820);
nor U41554 (N_41554,N_38198,N_36376);
nand U41555 (N_41555,N_36867,N_35677);
xor U41556 (N_41556,N_37483,N_36395);
xnor U41557 (N_41557,N_39349,N_37515);
and U41558 (N_41558,N_39533,N_39793);
nor U41559 (N_41559,N_37559,N_38244);
and U41560 (N_41560,N_38341,N_37287);
and U41561 (N_41561,N_39065,N_35149);
nor U41562 (N_41562,N_39824,N_38224);
xor U41563 (N_41563,N_39783,N_35715);
or U41564 (N_41564,N_39052,N_35818);
and U41565 (N_41565,N_35881,N_35590);
nand U41566 (N_41566,N_36815,N_35093);
nand U41567 (N_41567,N_35835,N_35025);
nand U41568 (N_41568,N_37523,N_38471);
xor U41569 (N_41569,N_37517,N_39230);
and U41570 (N_41570,N_39629,N_35474);
or U41571 (N_41571,N_35734,N_37709);
nor U41572 (N_41572,N_39685,N_35910);
and U41573 (N_41573,N_37373,N_36742);
nor U41574 (N_41574,N_35690,N_37439);
and U41575 (N_41575,N_39426,N_37539);
and U41576 (N_41576,N_35421,N_39089);
nor U41577 (N_41577,N_38895,N_35842);
or U41578 (N_41578,N_39985,N_35034);
or U41579 (N_41579,N_38701,N_36864);
nor U41580 (N_41580,N_35112,N_36918);
and U41581 (N_41581,N_35657,N_38136);
nand U41582 (N_41582,N_35810,N_37595);
or U41583 (N_41583,N_38268,N_38696);
nand U41584 (N_41584,N_36507,N_37455);
or U41585 (N_41585,N_35970,N_37977);
xnor U41586 (N_41586,N_35392,N_37859);
nand U41587 (N_41587,N_37721,N_36969);
nor U41588 (N_41588,N_36326,N_35903);
nor U41589 (N_41589,N_36684,N_39973);
and U41590 (N_41590,N_37823,N_37655);
and U41591 (N_41591,N_35746,N_36897);
and U41592 (N_41592,N_37031,N_36257);
or U41593 (N_41593,N_37218,N_35247);
nor U41594 (N_41594,N_36058,N_35165);
and U41595 (N_41595,N_36195,N_35377);
xnor U41596 (N_41596,N_36533,N_38165);
nand U41597 (N_41597,N_38336,N_37488);
nor U41598 (N_41598,N_39233,N_35535);
nand U41599 (N_41599,N_35991,N_37971);
xor U41600 (N_41600,N_35526,N_38000);
and U41601 (N_41601,N_35479,N_35246);
or U41602 (N_41602,N_39311,N_37596);
or U41603 (N_41603,N_35208,N_38924);
xnor U41604 (N_41604,N_35933,N_38131);
nand U41605 (N_41605,N_37290,N_37889);
nand U41606 (N_41606,N_35266,N_38395);
and U41607 (N_41607,N_39190,N_38890);
nor U41608 (N_41608,N_36754,N_38110);
nor U41609 (N_41609,N_35130,N_39797);
or U41610 (N_41610,N_37866,N_37041);
nand U41611 (N_41611,N_35393,N_38618);
xor U41612 (N_41612,N_38293,N_36795);
nand U41613 (N_41613,N_39928,N_35791);
or U41614 (N_41614,N_36056,N_35700);
nand U41615 (N_41615,N_36817,N_39645);
xnor U41616 (N_41616,N_39978,N_36851);
nor U41617 (N_41617,N_36303,N_36101);
nor U41618 (N_41618,N_35358,N_36626);
and U41619 (N_41619,N_35550,N_36054);
or U41620 (N_41620,N_38258,N_35347);
and U41621 (N_41621,N_39270,N_36529);
nor U41622 (N_41622,N_35611,N_37403);
and U41623 (N_41623,N_37211,N_36872);
nand U41624 (N_41624,N_36238,N_36194);
or U41625 (N_41625,N_39332,N_35647);
or U41626 (N_41626,N_35627,N_36783);
nand U41627 (N_41627,N_36016,N_35678);
and U41628 (N_41628,N_37123,N_38423);
nand U41629 (N_41629,N_38297,N_37793);
nor U41630 (N_41630,N_36653,N_35855);
xor U41631 (N_41631,N_35013,N_35563);
xnor U41632 (N_41632,N_39986,N_37979);
or U41633 (N_41633,N_39269,N_35538);
nand U41634 (N_41634,N_36794,N_37704);
nand U41635 (N_41635,N_36480,N_38558);
or U41636 (N_41636,N_35205,N_35995);
nand U41637 (N_41637,N_39297,N_38900);
or U41638 (N_41638,N_37056,N_36941);
nor U41639 (N_41639,N_39570,N_36330);
or U41640 (N_41640,N_35598,N_39549);
or U41641 (N_41641,N_36454,N_38058);
or U41642 (N_41642,N_36810,N_35011);
or U41643 (N_41643,N_38164,N_38113);
nor U41644 (N_41644,N_38402,N_37343);
and U41645 (N_41645,N_39051,N_35803);
or U41646 (N_41646,N_35619,N_38990);
and U41647 (N_41647,N_39605,N_38179);
nand U41648 (N_41648,N_35622,N_37855);
or U41649 (N_41649,N_35758,N_37461);
nand U41650 (N_41650,N_35914,N_39555);
xnor U41651 (N_41651,N_35376,N_37896);
nor U41652 (N_41652,N_39736,N_35919);
nand U41653 (N_41653,N_39405,N_35610);
and U41654 (N_41654,N_36769,N_39013);
nor U41655 (N_41655,N_35156,N_36360);
and U41656 (N_41656,N_36744,N_36689);
nor U41657 (N_41657,N_38226,N_39923);
nand U41658 (N_41658,N_35640,N_37638);
nor U41659 (N_41659,N_37315,N_36908);
nand U41660 (N_41660,N_35209,N_39005);
nand U41661 (N_41661,N_35967,N_39738);
xor U41662 (N_41662,N_35696,N_36338);
nand U41663 (N_41663,N_39175,N_38374);
or U41664 (N_41664,N_35792,N_35876);
or U41665 (N_41665,N_38458,N_36419);
xnor U41666 (N_41666,N_38962,N_39724);
nor U41667 (N_41667,N_39097,N_38667);
and U41668 (N_41668,N_39039,N_38999);
nand U41669 (N_41669,N_39203,N_38486);
and U41670 (N_41670,N_38548,N_39547);
nor U41671 (N_41671,N_37693,N_39974);
nand U41672 (N_41672,N_35607,N_39210);
and U41673 (N_41673,N_35895,N_39920);
nand U41674 (N_41674,N_36766,N_38759);
nor U41675 (N_41675,N_37754,N_35925);
or U41676 (N_41676,N_36854,N_39583);
nor U41677 (N_41677,N_36903,N_39194);
nand U41678 (N_41678,N_37816,N_36436);
nor U41679 (N_41679,N_35104,N_35768);
nor U41680 (N_41680,N_39528,N_38286);
or U41681 (N_41681,N_35334,N_35333);
nand U41682 (N_41682,N_38003,N_35385);
and U41683 (N_41683,N_35651,N_37264);
nor U41684 (N_41684,N_36551,N_39559);
xor U41685 (N_41685,N_35904,N_36948);
xor U41686 (N_41686,N_39558,N_35131);
and U41687 (N_41687,N_37758,N_35750);
and U41688 (N_41688,N_38841,N_38125);
nor U41689 (N_41689,N_38115,N_38697);
nand U41690 (N_41690,N_37062,N_35440);
nand U41691 (N_41691,N_35178,N_38401);
nand U41692 (N_41692,N_38545,N_38708);
nor U41693 (N_41693,N_36674,N_38686);
nor U41694 (N_41694,N_37907,N_39723);
nor U41695 (N_41695,N_37201,N_37804);
and U41696 (N_41696,N_36605,N_36314);
nor U41697 (N_41697,N_39303,N_39023);
and U41698 (N_41698,N_38816,N_39439);
or U41699 (N_41699,N_39539,N_38130);
xor U41700 (N_41700,N_35282,N_37735);
and U41701 (N_41701,N_36100,N_35330);
or U41702 (N_41702,N_38713,N_35958);
nor U41703 (N_41703,N_35203,N_39905);
nor U41704 (N_41704,N_38105,N_39675);
and U41705 (N_41705,N_35857,N_37850);
or U41706 (N_41706,N_37215,N_39534);
nor U41707 (N_41707,N_38066,N_38218);
and U41708 (N_41708,N_37024,N_37224);
or U41709 (N_41709,N_36914,N_38094);
or U41710 (N_41710,N_36787,N_35529);
nor U41711 (N_41711,N_38970,N_35506);
nor U41712 (N_41712,N_35464,N_36340);
or U41713 (N_41713,N_39193,N_36337);
nor U41714 (N_41714,N_36509,N_38185);
nand U41715 (N_41715,N_37556,N_35892);
nand U41716 (N_41716,N_39588,N_36548);
nor U41717 (N_41717,N_36755,N_39509);
and U41718 (N_41718,N_38581,N_39478);
and U41719 (N_41719,N_35843,N_35085);
nor U41720 (N_41720,N_37065,N_36459);
xnor U41721 (N_41721,N_38518,N_37262);
or U41722 (N_41722,N_36874,N_37710);
nor U41723 (N_41723,N_38129,N_36869);
and U41724 (N_41724,N_37249,N_35714);
nor U41725 (N_41725,N_39243,N_35023);
and U41726 (N_41726,N_37142,N_38381);
or U41727 (N_41727,N_39772,N_36707);
or U41728 (N_41728,N_38981,N_39021);
and U41729 (N_41729,N_38622,N_37325);
nand U41730 (N_41730,N_39164,N_36199);
nand U41731 (N_41731,N_36328,N_35656);
nand U41732 (N_41732,N_35828,N_38580);
and U41733 (N_41733,N_35335,N_38261);
xor U41734 (N_41734,N_36055,N_37446);
or U41735 (N_41735,N_36305,N_38514);
and U41736 (N_41736,N_36965,N_37728);
or U41737 (N_41737,N_38469,N_37621);
or U41738 (N_41738,N_35999,N_39008);
and U41739 (N_41739,N_35778,N_38455);
and U41740 (N_41740,N_37005,N_37564);
and U41741 (N_41741,N_36757,N_36722);
and U41742 (N_41742,N_36820,N_38612);
xnor U41743 (N_41743,N_39150,N_35681);
nor U41744 (N_41744,N_37574,N_38658);
or U41745 (N_41745,N_35920,N_36858);
and U41746 (N_41746,N_39531,N_35533);
nand U41747 (N_41747,N_35468,N_39325);
xnor U41748 (N_41748,N_37036,N_39250);
nor U41749 (N_41749,N_39264,N_39599);
and U41750 (N_41750,N_39506,N_36181);
or U41751 (N_41751,N_35461,N_36222);
xnor U41752 (N_41752,N_38280,N_37657);
and U41753 (N_41753,N_35532,N_35721);
and U41754 (N_41754,N_37135,N_37606);
nand U41755 (N_41755,N_36531,N_35454);
and U41756 (N_41756,N_35510,N_38182);
nor U41757 (N_41757,N_39404,N_36643);
nor U41758 (N_41758,N_37546,N_38019);
and U41759 (N_41759,N_37857,N_39743);
nor U41760 (N_41760,N_38444,N_39855);
nor U41761 (N_41761,N_36364,N_38189);
or U41762 (N_41762,N_37613,N_39914);
or U41763 (N_41763,N_38998,N_39273);
or U41764 (N_41764,N_38877,N_36594);
nor U41765 (N_41765,N_38159,N_38839);
nor U41766 (N_41766,N_39664,N_36142);
xor U41767 (N_41767,N_38741,N_36972);
or U41768 (N_41768,N_37522,N_36288);
nor U41769 (N_41769,N_38873,N_39764);
xnor U41770 (N_41770,N_37321,N_39849);
and U41771 (N_41771,N_38724,N_37395);
or U41772 (N_41772,N_39532,N_36746);
xnor U41773 (N_41773,N_38695,N_39197);
nand U41774 (N_41774,N_37870,N_38491);
nand U41775 (N_41775,N_35515,N_35813);
nand U41776 (N_41776,N_38509,N_38671);
nor U41777 (N_41777,N_37335,N_36415);
or U41778 (N_41778,N_38420,N_35074);
and U41779 (N_41779,N_37424,N_39217);
and U41780 (N_41780,N_35670,N_36824);
or U41781 (N_41781,N_39561,N_37609);
and U41782 (N_41782,N_39615,N_37430);
or U41783 (N_41783,N_36993,N_36883);
or U41784 (N_41784,N_38194,N_35773);
or U41785 (N_41785,N_37385,N_35983);
nand U41786 (N_41786,N_37225,N_39919);
xor U41787 (N_41787,N_37177,N_39049);
or U41788 (N_41788,N_39066,N_38273);
and U41789 (N_41789,N_35923,N_37745);
and U41790 (N_41790,N_39883,N_37166);
nand U41791 (N_41791,N_36146,N_37764);
or U41792 (N_41792,N_35382,N_36672);
or U41793 (N_41793,N_36250,N_35039);
or U41794 (N_41794,N_39959,N_38083);
and U41795 (N_41795,N_36964,N_38788);
and U41796 (N_41796,N_36317,N_39578);
and U41797 (N_41797,N_39446,N_37862);
nand U41798 (N_41798,N_39560,N_36348);
xor U41799 (N_41799,N_37411,N_37178);
nor U41800 (N_41800,N_36109,N_37148);
nor U41801 (N_41801,N_35680,N_36034);
and U41802 (N_41802,N_36327,N_38200);
or U41803 (N_41803,N_35113,N_36160);
or U41804 (N_41804,N_38495,N_36849);
nand U41805 (N_41805,N_39868,N_38737);
nand U41806 (N_41806,N_39650,N_35232);
nor U41807 (N_41807,N_35343,N_39913);
xnor U41808 (N_41808,N_38351,N_36917);
nor U41809 (N_41809,N_35398,N_39552);
nand U41810 (N_41810,N_36446,N_36393);
nand U41811 (N_41811,N_35816,N_37702);
and U41812 (N_41812,N_35985,N_37890);
and U41813 (N_41813,N_39459,N_38005);
and U41814 (N_41814,N_35413,N_37255);
nand U41815 (N_41815,N_39411,N_37806);
or U41816 (N_41816,N_35679,N_36490);
and U41817 (N_41817,N_37727,N_35852);
nor U41818 (N_41818,N_36244,N_36778);
nor U41819 (N_41819,N_36357,N_37840);
or U41820 (N_41820,N_38067,N_35922);
or U41821 (N_41821,N_36841,N_37390);
or U41822 (N_41822,N_37761,N_37082);
and U41823 (N_41823,N_38961,N_36157);
nor U41824 (N_41824,N_38400,N_39429);
and U41825 (N_41825,N_37972,N_38838);
or U41826 (N_41826,N_35638,N_36580);
nor U41827 (N_41827,N_39770,N_39634);
nor U41828 (N_41828,N_38569,N_36737);
xnor U41829 (N_41829,N_39830,N_38208);
nor U41830 (N_41830,N_39341,N_39161);
and U41831 (N_41831,N_37001,N_35193);
xor U41832 (N_41832,N_35737,N_39791);
nor U41833 (N_41833,N_39606,N_36403);
or U41834 (N_41834,N_37770,N_37661);
nand U41835 (N_41835,N_35243,N_36634);
and U41836 (N_41836,N_37525,N_37644);
nand U41837 (N_41837,N_35269,N_36203);
or U41838 (N_41838,N_39348,N_37417);
or U41839 (N_41839,N_35255,N_38515);
and U41840 (N_41840,N_36561,N_38605);
or U41841 (N_41841,N_37196,N_35493);
and U41842 (N_41842,N_38813,N_36290);
and U41843 (N_41843,N_35134,N_36721);
and U41844 (N_41844,N_37382,N_35868);
nand U41845 (N_41845,N_39302,N_37084);
or U41846 (N_41846,N_36147,N_37886);
nor U41847 (N_41847,N_39356,N_35094);
or U41848 (N_41848,N_38151,N_36306);
and U41849 (N_41849,N_36986,N_37388);
nand U41850 (N_41850,N_35965,N_36660);
nand U41851 (N_41851,N_37980,N_37527);
nand U41852 (N_41852,N_35410,N_36517);
nand U41853 (N_41853,N_36968,N_39158);
xor U41854 (N_41854,N_39911,N_37133);
nor U41855 (N_41855,N_36302,N_38358);
or U41856 (N_41856,N_36205,N_37003);
nand U41857 (N_41857,N_38854,N_38259);
nand U41858 (N_41858,N_36155,N_35588);
xnor U41859 (N_41859,N_39457,N_38774);
and U41860 (N_41860,N_35572,N_37923);
nand U41861 (N_41861,N_36421,N_39909);
or U41862 (N_41862,N_37450,N_39196);
and U41863 (N_41863,N_37299,N_38933);
xor U41864 (N_41864,N_39095,N_36373);
nand U41865 (N_41865,N_38383,N_35177);
nor U41866 (N_41866,N_35349,N_37377);
nor U41867 (N_41867,N_38820,N_35849);
nand U41868 (N_41868,N_36300,N_35047);
nand U41869 (N_41869,N_37967,N_38048);
xnor U41870 (N_41870,N_38137,N_37426);
nor U41871 (N_41871,N_36200,N_38499);
nor U41872 (N_41872,N_39072,N_37838);
or U41873 (N_41873,N_38913,N_35603);
or U41874 (N_41874,N_39524,N_36416);
xor U41875 (N_41875,N_38234,N_35630);
nor U41876 (N_41876,N_39424,N_39160);
and U41877 (N_41877,N_39372,N_39862);
xnor U41878 (N_41878,N_37414,N_35028);
or U41879 (N_41879,N_36612,N_39892);
nor U41880 (N_41880,N_38157,N_35004);
nor U41881 (N_41881,N_39309,N_37848);
nor U41882 (N_41882,N_38700,N_35181);
nand U41883 (N_41883,N_35078,N_37821);
nand U41884 (N_41884,N_38228,N_35697);
nor U41885 (N_41885,N_37711,N_36095);
and U41886 (N_41886,N_37070,N_37320);
nand U41887 (N_41887,N_37987,N_37575);
or U41888 (N_41888,N_35898,N_35908);
and U41889 (N_41889,N_36596,N_36407);
xor U41890 (N_41890,N_35508,N_36608);
nor U41891 (N_41891,N_37995,N_39462);
nand U41892 (N_41892,N_35698,N_35147);
nand U41893 (N_41893,N_39307,N_35226);
or U41894 (N_41894,N_39450,N_39591);
nand U41895 (N_41895,N_39173,N_36538);
and U41896 (N_41896,N_37583,N_37279);
and U41897 (N_41897,N_36597,N_38505);
and U41898 (N_41898,N_39589,N_39661);
xnor U41899 (N_41899,N_36777,N_36738);
or U41900 (N_41900,N_37841,N_35053);
and U41901 (N_41901,N_36039,N_36445);
nor U41902 (N_41902,N_38210,N_38889);
nor U41903 (N_41903,N_37542,N_35874);
or U41904 (N_41904,N_35722,N_39146);
and U41905 (N_41905,N_39711,N_39550);
or U41906 (N_41906,N_38012,N_37756);
nor U41907 (N_41907,N_38231,N_38091);
nand U41908 (N_41908,N_39689,N_37433);
and U41909 (N_41909,N_38432,N_36134);
nor U41910 (N_41910,N_36636,N_36164);
or U41911 (N_41911,N_38169,N_38526);
xor U41912 (N_41912,N_37507,N_39996);
or U41913 (N_41913,N_37506,N_38037);
xnor U41914 (N_41914,N_39025,N_36065);
and U41915 (N_41915,N_38428,N_38387);
and U41916 (N_41916,N_39681,N_36041);
or U41917 (N_41917,N_35704,N_36892);
nand U41918 (N_41918,N_35135,N_37891);
and U41919 (N_41919,N_38893,N_38047);
nand U41920 (N_41920,N_36554,N_35541);
and U41921 (N_41921,N_36110,N_35244);
nand U41922 (N_41922,N_39215,N_37827);
or U41923 (N_41923,N_35079,N_37470);
or U41924 (N_41924,N_38219,N_39845);
xor U41925 (N_41925,N_38979,N_38939);
or U41926 (N_41926,N_39035,N_38365);
xor U41927 (N_41927,N_35875,N_37367);
nor U41928 (N_41928,N_36345,N_36005);
nor U41929 (N_41929,N_36866,N_36120);
nor U41930 (N_41930,N_35666,N_36469);
and U41931 (N_41931,N_39962,N_39287);
nand U41932 (N_41932,N_35501,N_36904);
or U41933 (N_41933,N_38568,N_39734);
or U41934 (N_41934,N_38062,N_37954);
and U41935 (N_41935,N_38940,N_36243);
nor U41936 (N_41936,N_37653,N_36441);
and U41937 (N_41937,N_35210,N_37869);
and U41938 (N_41938,N_38004,N_38977);
xor U41939 (N_41939,N_36621,N_36123);
xor U41940 (N_41940,N_36275,N_35251);
nor U41941 (N_41941,N_37775,N_39976);
and U41942 (N_41942,N_37064,N_37203);
and U41943 (N_41943,N_38266,N_36541);
or U41944 (N_41944,N_37958,N_37534);
nand U41945 (N_41945,N_38481,N_36131);
and U41946 (N_41946,N_37864,N_39582);
or U41947 (N_41947,N_37697,N_36990);
xnor U41948 (N_41948,N_36826,N_36271);
and U41949 (N_41949,N_35496,N_39198);
and U41950 (N_41950,N_38020,N_37231);
nor U41951 (N_41951,N_38572,N_37427);
or U41952 (N_41952,N_38687,N_38674);
nor U41953 (N_41953,N_38822,N_37115);
nand U41954 (N_41954,N_35645,N_38902);
nor U41955 (N_41955,N_37587,N_36776);
and U41956 (N_41956,N_36458,N_36448);
nand U41957 (N_41957,N_38984,N_35779);
nor U41958 (N_41958,N_38196,N_36569);
and U41959 (N_41959,N_39363,N_35316);
nor U41960 (N_41960,N_39801,N_35996);
and U41961 (N_41961,N_39208,N_35102);
nand U41962 (N_41962,N_37872,N_36268);
nor U41963 (N_41963,N_37846,N_39934);
nor U41964 (N_41964,N_38779,N_38191);
and U41965 (N_41965,N_35482,N_39693);
and U41966 (N_41966,N_38763,N_38806);
nand U41967 (N_41967,N_36402,N_36666);
nand U41968 (N_41968,N_37668,N_37835);
and U41969 (N_41969,N_36211,N_39260);
and U41970 (N_41970,N_37420,N_38669);
nand U41971 (N_41971,N_36648,N_39520);
nand U41972 (N_41972,N_39844,N_35926);
nor U41973 (N_41973,N_37536,N_38327);
and U41974 (N_41974,N_35728,N_39702);
and U41975 (N_41975,N_39228,N_37650);
and U41976 (N_41976,N_39276,N_38026);
nand U41977 (N_41977,N_39067,N_38227);
nand U41978 (N_41978,N_35940,N_37978);
nand U41979 (N_41979,N_37336,N_38639);
nand U41980 (N_41980,N_35164,N_37738);
and U41981 (N_41981,N_39317,N_39929);
nor U41982 (N_41982,N_35785,N_39980);
nand U41983 (N_41983,N_39266,N_35362);
and U41984 (N_41984,N_38706,N_35262);
nand U41985 (N_41985,N_35315,N_39686);
and U41986 (N_41986,N_37592,N_35682);
nor U41987 (N_41987,N_38064,N_35867);
or U41988 (N_41988,N_39063,N_39200);
or U41989 (N_41989,N_38500,N_35394);
xnor U41990 (N_41990,N_37569,N_38215);
nor U41991 (N_41991,N_39017,N_37004);
and U41992 (N_41992,N_36313,N_38552);
and U41993 (N_41993,N_38429,N_39187);
or U41994 (N_41994,N_37477,N_39903);
or U41995 (N_41995,N_37256,N_37696);
or U41996 (N_41996,N_37050,N_37113);
or U41997 (N_41997,N_36645,N_38973);
xnor U41998 (N_41998,N_39915,N_37501);
nand U41999 (N_41999,N_36124,N_39626);
nand U42000 (N_42000,N_37456,N_39544);
xnor U42001 (N_42001,N_37091,N_36973);
nor U42002 (N_42002,N_39593,N_36412);
and U42003 (N_42003,N_35491,N_39683);
or U42004 (N_42004,N_38307,N_35797);
nand U42005 (N_42005,N_37183,N_37918);
and U42006 (N_42006,N_36670,N_38803);
xor U42007 (N_42007,N_35449,N_36891);
and U42008 (N_42008,N_35293,N_37737);
or U42009 (N_42009,N_39718,N_35190);
nand U42010 (N_42010,N_38930,N_36125);
nor U42011 (N_42011,N_37127,N_38478);
xnor U42012 (N_42012,N_37272,N_35573);
and U42013 (N_42013,N_36808,N_35054);
and U42014 (N_42014,N_38557,N_35584);
or U42015 (N_42015,N_38007,N_36368);
nor U42016 (N_42016,N_37184,N_37612);
nand U42017 (N_42017,N_38315,N_36498);
and U42018 (N_42018,N_38678,N_36745);
nand U42019 (N_42019,N_35736,N_39853);
and U42020 (N_42020,N_37226,N_37392);
and U42021 (N_42021,N_39994,N_37562);
and U42022 (N_42022,N_35045,N_39907);
or U42023 (N_42023,N_36652,N_39497);
and U42024 (N_42024,N_36196,N_36719);
and U42025 (N_42025,N_35063,N_37582);
and U42026 (N_42026,N_36422,N_35286);
nor U42027 (N_42027,N_37493,N_38016);
nand U42028 (N_42028,N_39154,N_37204);
and U42029 (N_42029,N_38988,N_37173);
nand U42030 (N_42030,N_35137,N_37409);
or U42031 (N_42031,N_38842,N_36798);
nor U42032 (N_42032,N_38276,N_37760);
and U42033 (N_42033,N_37194,N_35641);
nand U42034 (N_42034,N_36223,N_37362);
nor U42035 (N_42035,N_35037,N_36939);
nor U42036 (N_42036,N_38099,N_37258);
xnor U42037 (N_42037,N_35092,N_36945);
or U42038 (N_42038,N_38616,N_38875);
or U42039 (N_42039,N_36928,N_36750);
nor U42040 (N_42040,N_36374,N_37925);
nor U42041 (N_42041,N_35760,N_37541);
nor U42042 (N_42042,N_35424,N_39103);
nand U42043 (N_42043,N_36264,N_36536);
nand U42044 (N_42044,N_35118,N_39530);
and U42045 (N_42045,N_37953,N_37946);
or U42046 (N_42046,N_38264,N_38222);
nor U42047 (N_42047,N_38874,N_35381);
or U42048 (N_42048,N_37170,N_36566);
and U42049 (N_42049,N_39811,N_38265);
nand U42050 (N_42050,N_37549,N_38934);
and U42051 (N_42051,N_36520,N_37654);
or U42052 (N_42052,N_37423,N_35909);
nor U42053 (N_42053,N_36266,N_38385);
nand U42054 (N_42054,N_36876,N_35733);
or U42055 (N_42055,N_35998,N_36584);
xor U42056 (N_42056,N_39386,N_36085);
or U42057 (N_42057,N_36087,N_35182);
nand U42058 (N_42058,N_38288,N_39672);
and U42059 (N_42059,N_38997,N_36406);
nor U42060 (N_42060,N_35274,N_38784);
nor U42061 (N_42061,N_37512,N_35993);
and U42062 (N_42062,N_35693,N_36213);
nand U42063 (N_42063,N_35056,N_35119);
or U42064 (N_42064,N_38472,N_35227);
or U42065 (N_42065,N_35725,N_39829);
or U42066 (N_42066,N_38403,N_38319);
or U42067 (N_42067,N_38650,N_39453);
xor U42068 (N_42068,N_38027,N_37802);
or U42069 (N_42069,N_36168,N_39240);
or U42070 (N_42070,N_35789,N_35499);
nor U42071 (N_42071,N_35352,N_37412);
nand U42072 (N_42072,N_39128,N_39371);
nor U42073 (N_42073,N_38599,N_39402);
nor U42074 (N_42074,N_37109,N_35829);
nand U42075 (N_42075,N_38818,N_38857);
and U42076 (N_42076,N_37105,N_36209);
nor U42077 (N_42077,N_36371,N_39825);
nand U42078 (N_42078,N_37330,N_37360);
and U42079 (N_42079,N_37695,N_35298);
nand U42080 (N_42080,N_39062,N_35206);
xor U42081 (N_42081,N_35509,N_38559);
and U42082 (N_42082,N_38760,N_35505);
or U42083 (N_42083,N_36482,N_35215);
or U42084 (N_42084,N_38899,N_35030);
xnor U42085 (N_42085,N_36686,N_37486);
nor U42086 (N_42086,N_37579,N_35195);
or U42087 (N_42087,N_38915,N_36325);
nor U42088 (N_42088,N_38102,N_35831);
nor U42089 (N_42089,N_35626,N_37045);
nand U42090 (N_42090,N_37072,N_39126);
and U42091 (N_42091,N_38789,N_37986);
or U42092 (N_42092,N_36912,N_37171);
nor U42093 (N_42093,N_37000,N_39885);
nor U42094 (N_42094,N_38308,N_35348);
xnor U42095 (N_42095,N_37502,N_38096);
nor U42096 (N_42096,N_35934,N_38107);
nand U42097 (N_42097,N_39342,N_37904);
nand U42098 (N_42098,N_37429,N_38717);
nand U42099 (N_42099,N_37008,N_37920);
xnor U42100 (N_42100,N_37768,N_37819);
nand U42101 (N_42101,N_38431,N_37327);
nor U42102 (N_42102,N_38285,N_38171);
and U42103 (N_42103,N_38698,N_39221);
nand U42104 (N_42104,N_37640,N_35592);
nor U42105 (N_42105,N_36251,N_35801);
or U42106 (N_42106,N_38425,N_37883);
xnor U42107 (N_42107,N_39357,N_38155);
or U42108 (N_42108,N_35400,N_39469);
and U42109 (N_42109,N_37359,N_36606);
nor U42110 (N_42110,N_36127,N_39744);
nand U42111 (N_42111,N_35133,N_39053);
xor U42112 (N_42112,N_35239,N_38720);
or U42113 (N_42113,N_37400,N_36187);
or U42114 (N_42114,N_36816,N_36115);
nor U42115 (N_42115,N_39022,N_37809);
or U42116 (N_42116,N_37155,N_38693);
and U42117 (N_42117,N_35766,N_38068);
nand U42118 (N_42118,N_35378,N_35886);
nand U42119 (N_42119,N_35608,N_35167);
or U42120 (N_42120,N_38743,N_35388);
nor U42121 (N_42121,N_38703,N_35788);
and U42122 (N_42122,N_37843,N_39108);
or U42123 (N_42123,N_38361,N_38955);
or U42124 (N_42124,N_37568,N_37318);
nor U42125 (N_42125,N_36833,N_38009);
or U42126 (N_42126,N_36832,N_37391);
nand U42127 (N_42127,N_38726,N_38797);
and U42128 (N_42128,N_35295,N_39245);
or U42129 (N_42129,N_39281,N_38370);
or U42130 (N_42130,N_36320,N_39218);
nor U42131 (N_42131,N_39790,N_36848);
and U42132 (N_42132,N_38507,N_37903);
xor U42133 (N_42133,N_35435,N_35901);
nand U42134 (N_42134,N_35668,N_37124);
nand U42135 (N_42135,N_39091,N_35220);
nor U42136 (N_42136,N_38595,N_36438);
nand U42137 (N_42137,N_38589,N_38975);
nand U42138 (N_42138,N_37146,N_36119);
or U42139 (N_42139,N_35263,N_35283);
or U42140 (N_42140,N_37985,N_37074);
and U42141 (N_42141,N_35863,N_39454);
nor U42142 (N_42142,N_36346,N_38207);
xnor U42143 (N_42143,N_35777,N_35084);
nand U42144 (N_42144,N_39958,N_37601);
nand U42145 (N_42145,N_38565,N_39206);
or U42146 (N_42146,N_35655,N_35222);
nand U42147 (N_42147,N_39990,N_38138);
or U42148 (N_42148,N_38466,N_37156);
nand U42149 (N_42149,N_36130,N_37371);
nor U42150 (N_42150,N_39300,N_36886);
nand U42151 (N_42151,N_39614,N_39456);
nor U42152 (N_42152,N_37223,N_39098);
or U42153 (N_42153,N_37951,N_36570);
or U42154 (N_42154,N_37947,N_36372);
nor U42155 (N_42155,N_36739,N_37112);
or U42156 (N_42156,N_39431,N_39274);
nor U42157 (N_42157,N_39792,N_38140);
and U42158 (N_42158,N_37267,N_36210);
nor U42159 (N_42159,N_38722,N_36008);
xnor U42160 (N_42160,N_39712,N_35837);
or U42161 (N_42161,N_35531,N_38868);
nand U42162 (N_42162,N_38534,N_37950);
nand U42163 (N_42163,N_39594,N_36118);
nor U42164 (N_42164,N_39099,N_39612);
and U42165 (N_42165,N_37042,N_39277);
nor U42166 (N_42166,N_37844,N_36494);
nor U42167 (N_42167,N_36132,N_37732);
nand U42168 (N_42168,N_37581,N_38209);
nor U42169 (N_42169,N_39609,N_38652);
and U42170 (N_42170,N_36010,N_39657);
nand U42171 (N_42171,N_38888,N_36354);
xor U42172 (N_42172,N_37622,N_37685);
or U42173 (N_42173,N_39149,N_37803);
nand U42174 (N_42174,N_38951,N_39639);
and U42175 (N_42175,N_39259,N_38801);
nor U42176 (N_42176,N_39234,N_39623);
nand U42177 (N_42177,N_35793,N_36282);
or U42178 (N_42178,N_35562,N_36191);
or U42179 (N_42179,N_36072,N_35342);
or U42180 (N_42180,N_36681,N_38593);
and U42181 (N_42181,N_39863,N_39179);
xnor U42182 (N_42182,N_35977,N_38709);
nor U42183 (N_42183,N_36957,N_39601);
nor U42184 (N_42184,N_36960,N_37284);
and U42185 (N_42185,N_36765,N_37457);
nand U42186 (N_42186,N_37939,N_36955);
nand U42187 (N_42187,N_36768,N_36316);
and U42188 (N_42188,N_36411,N_39375);
or U42189 (N_42189,N_35500,N_35387);
nand U42190 (N_42190,N_39380,N_38176);
nor U42191 (N_42191,N_38679,N_35356);
xnor U42192 (N_42192,N_36444,N_36910);
nand U42193 (N_42193,N_37088,N_38950);
or U42194 (N_42194,N_36361,N_36665);
nor U42195 (N_42195,N_35912,N_36773);
nand U42196 (N_42196,N_37453,N_37206);
and U42197 (N_42197,N_39779,N_37586);
and U42198 (N_42198,N_37081,N_37594);
nor U42199 (N_42199,N_36595,N_35099);
nor U42200 (N_42200,N_39455,N_39410);
or U42201 (N_42201,N_39837,N_38535);
or U42202 (N_42202,N_37140,N_38662);
or U42203 (N_42203,N_35560,N_36353);
nand U42204 (N_42204,N_36192,N_36845);
or U42205 (N_42205,N_36215,N_39180);
and U42206 (N_42206,N_38632,N_38928);
xor U42207 (N_42207,N_38834,N_37759);
xnor U42208 (N_42208,N_36089,N_38271);
or U42209 (N_42209,N_37180,N_36630);
and U42210 (N_42210,N_36104,N_38856);
and U42211 (N_42211,N_37452,N_35049);
nor U42212 (N_42212,N_35090,N_37021);
and U42213 (N_42213,N_39399,N_37037);
xor U42214 (N_42214,N_39608,N_37962);
nand U42215 (N_42215,N_39165,N_39427);
nor U42216 (N_42216,N_39982,N_35152);
nand U42217 (N_42217,N_38190,N_35009);
nand U42218 (N_42218,N_39900,N_35935);
nand U42219 (N_42219,N_37076,N_39717);
nor U42220 (N_42220,N_38738,N_38459);
nand U42221 (N_42221,N_38335,N_35599);
and U42222 (N_42222,N_35615,N_37747);
and U42223 (N_42223,N_36861,N_38974);
and U42224 (N_42224,N_38127,N_39648);
nand U42225 (N_42225,N_37030,N_36461);
nand U42226 (N_42226,N_36096,N_35859);
nand U42227 (N_42227,N_35016,N_35042);
nor U42228 (N_42228,N_39448,N_38923);
nand U42229 (N_42229,N_38793,N_35964);
nand U42230 (N_42230,N_38879,N_36629);
nor U42231 (N_42231,N_38404,N_39474);
nor U42232 (N_42232,N_36558,N_39078);
xnor U42233 (N_42233,N_39747,N_36698);
nor U42234 (N_42234,N_38418,N_35163);
and U42235 (N_42235,N_38248,N_35887);
or U42236 (N_42236,N_39329,N_35260);
nor U42237 (N_42237,N_37102,N_36873);
and U42238 (N_42238,N_35350,N_38496);
xor U42239 (N_42239,N_35872,N_38272);
nand U42240 (N_42240,N_35928,N_37282);
nor U42241 (N_42241,N_37611,N_35219);
or U42242 (N_42242,N_35591,N_35568);
xor U42243 (N_42243,N_35370,N_38427);
and U42244 (N_42244,N_39010,N_36806);
or U42245 (N_42245,N_37545,N_37672);
nor U42246 (N_42246,N_39381,N_37213);
and U42247 (N_42247,N_38843,N_39936);
and U42248 (N_42248,N_38949,N_39949);
and U42249 (N_42249,N_36487,N_38761);
and U42250 (N_42250,N_36931,N_35160);
and U42251 (N_42251,N_37669,N_37537);
nor U42252 (N_42252,N_35481,N_36335);
or U42253 (N_42253,N_36170,N_39513);
or U42254 (N_42254,N_37724,N_39157);
xnor U42255 (N_42255,N_39141,N_36888);
nor U42256 (N_42256,N_39481,N_35401);
or U42257 (N_42257,N_35395,N_37128);
nand U42258 (N_42258,N_36557,N_38497);
or U42259 (N_42259,N_37464,N_39070);
nor U42260 (N_42260,N_37543,N_35618);
nand U42261 (N_42261,N_35143,N_38887);
and U42262 (N_42262,N_36287,N_37540);
or U42263 (N_42263,N_38814,N_38405);
or U42264 (N_42264,N_36602,N_35625);
or U42265 (N_42265,N_37598,N_37785);
or U42266 (N_42266,N_35340,N_36351);
xor U42267 (N_42267,N_39419,N_35948);
or U42268 (N_42268,N_39102,N_36641);
nor U42269 (N_42269,N_38625,N_35096);
nand U42270 (N_42270,N_35504,N_39461);
xnor U42271 (N_42271,N_36622,N_38826);
nor U42272 (N_42272,N_37961,N_38283);
and U42273 (N_42273,N_35057,N_36631);
nor U42274 (N_42274,N_36081,N_38439);
nand U42275 (N_42275,N_39904,N_36677);
nand U42276 (N_42276,N_35634,N_38771);
nand U42277 (N_42277,N_35207,N_36183);
or U42278 (N_42278,N_36321,N_35427);
or U42279 (N_42279,N_39806,N_39636);
nand U42280 (N_42280,N_38177,N_36375);
nor U42281 (N_42281,N_35833,N_39291);
nand U42282 (N_42282,N_36830,N_37440);
xor U42283 (N_42283,N_39432,N_36204);
or U42284 (N_42284,N_39466,N_37481);
and U42285 (N_42285,N_39253,N_35604);
or U42286 (N_42286,N_35537,N_37144);
nand U42287 (N_42287,N_36387,N_38203);
and U42288 (N_42288,N_36295,N_38367);
or U42289 (N_42289,N_37959,N_38412);
and U42290 (N_42290,N_38246,N_35418);
nand U42291 (N_42291,N_37309,N_37808);
or U42292 (N_42292,N_38187,N_36078);
or U42293 (N_42293,N_37068,N_36092);
or U42294 (N_42294,N_39222,N_39112);
or U42295 (N_42295,N_35425,N_36544);
nand U42296 (N_42296,N_37530,N_37936);
nor U42297 (N_42297,N_35273,N_38201);
nor U42298 (N_42298,N_35238,N_36234);
or U42299 (N_42299,N_35658,N_38927);
nor U42300 (N_42300,N_38086,N_38659);
nor U42301 (N_42301,N_39722,N_37748);
nand U42302 (N_42302,N_35751,N_35763);
or U42303 (N_42303,N_39301,N_35754);
and U42304 (N_42304,N_39969,N_39838);
xor U42305 (N_42305,N_38712,N_38001);
or U42306 (N_42306,N_37229,N_37607);
or U42307 (N_42307,N_39188,N_35689);
nand U42308 (N_42308,N_36363,N_38262);
or U42309 (N_42309,N_37617,N_39565);
nand U42310 (N_42310,N_39346,N_37384);
or U42311 (N_42311,N_35198,N_39728);
or U42312 (N_42312,N_36590,N_36752);
and U42313 (N_42313,N_39563,N_36951);
nor U42314 (N_42314,N_38386,N_38519);
nor U42315 (N_42315,N_36772,N_36274);
or U42316 (N_42316,N_38986,N_37312);
nand U42317 (N_42317,N_38483,N_35502);
xor U42318 (N_42318,N_35036,N_39745);
and U42319 (N_42319,N_38339,N_35765);
nor U42320 (N_42320,N_36976,N_37044);
and U42321 (N_42321,N_36399,N_35582);
and U42322 (N_42322,N_35429,N_36493);
or U42323 (N_42323,N_39393,N_39085);
xnor U42324 (N_42324,N_38892,N_38236);
or U42325 (N_42325,N_37368,N_38232);
nor U42326 (N_42326,N_39440,N_35302);
or U42327 (N_42327,N_38912,N_35027);
or U42328 (N_42328,N_35176,N_39105);
nand U42329 (N_42329,N_38586,N_37465);
and U42330 (N_42330,N_36617,N_39739);
nand U42331 (N_42331,N_37478,N_37706);
nor U42332 (N_42332,N_36682,N_37167);
or U42333 (N_42333,N_37355,N_37101);
or U42334 (N_42334,N_39347,N_35559);
nor U42335 (N_42335,N_37236,N_35001);
nor U42336 (N_42336,N_39422,N_37983);
and U42337 (N_42337,N_38163,N_36906);
and U42338 (N_42338,N_38357,N_35692);
xor U42339 (N_42339,N_36253,N_38031);
and U42340 (N_42340,N_38149,N_36088);
or U42341 (N_42341,N_35336,N_36332);
or U42342 (N_42342,N_36624,N_37941);
and U42343 (N_42343,N_39059,N_36717);
nand U42344 (N_42344,N_37246,N_38144);
or U42345 (N_42345,N_36992,N_35540);
nand U42346 (N_42346,N_36834,N_35089);
and U42347 (N_42347,N_39166,N_35391);
and U42348 (N_42348,N_35706,N_39659);
nor U42349 (N_42349,N_38980,N_39527);
and U42350 (N_42350,N_35399,N_37511);
nor U42351 (N_42351,N_35710,N_37794);
nor U42352 (N_42352,N_35486,N_39647);
or U42353 (N_42353,N_39263,N_37529);
or U42354 (N_42354,N_36082,N_36625);
and U42355 (N_42355,N_37438,N_37278);
xnor U42356 (N_42356,N_36379,N_35052);
or U42357 (N_42357,N_37830,N_35374);
and U42358 (N_42358,N_39826,N_36900);
nand U42359 (N_42359,N_37909,N_36814);
xor U42360 (N_42360,N_37730,N_37182);
nand U42361 (N_42361,N_35513,N_35858);
nand U42362 (N_42362,N_36675,N_36483);
xor U42363 (N_42363,N_37071,N_39398);
or U42364 (N_42364,N_36601,N_37344);
nor U42365 (N_42365,N_37342,N_38430);
and U42366 (N_42366,N_39529,N_37307);
and U42367 (N_42367,N_38582,N_38371);
or U42368 (N_42368,N_36895,N_37558);
nand U42369 (N_42369,N_35844,N_35724);
nor U42370 (N_42370,N_35747,N_36037);
nor U42371 (N_42371,N_37443,N_36075);
nand U42372 (N_42372,N_36614,N_38870);
xor U42373 (N_42373,N_35821,N_36882);
nor U42374 (N_42374,N_39444,N_38141);
and U42375 (N_42375,N_37531,N_39515);
xor U42376 (N_42376,N_38604,N_35460);
or U42377 (N_42377,N_37270,N_37635);
nand U42378 (N_42378,N_35265,N_39251);
nor U42379 (N_42379,N_36137,N_39113);
and U42380 (N_42380,N_39003,N_36179);
and U42381 (N_42381,N_38109,N_39033);
or U42382 (N_42382,N_35197,N_38747);
nand U42383 (N_42383,N_38576,N_35051);
or U42384 (N_42384,N_36838,N_37052);
nor U42385 (N_42385,N_39521,N_38562);
or U42386 (N_42386,N_39288,N_39912);
nand U42387 (N_42387,N_35138,N_37108);
and U42388 (N_42388,N_38166,N_37518);
nor U42389 (N_42389,N_39152,N_36188);
and U42390 (N_42390,N_39452,N_38976);
xor U42391 (N_42391,N_38461,N_37499);
nor U42392 (N_42392,N_35916,N_37387);
and U42393 (N_42393,N_36018,N_37040);
xnor U42394 (N_42394,N_38983,N_36401);
nand U42395 (N_42395,N_36024,N_39271);
xnor U42396 (N_42396,N_39485,N_36526);
or U42397 (N_42397,N_39756,N_37375);
and U42398 (N_42398,N_35044,N_37646);
or U42399 (N_42399,N_35456,N_37729);
nor U42400 (N_42400,N_37940,N_36304);
or U42401 (N_42401,N_37687,N_37298);
nand U42402 (N_42402,N_36154,N_36823);
nor U42403 (N_42403,N_35379,N_36116);
and U42404 (N_42404,N_37230,N_38844);
nor U42405 (N_42405,N_35179,N_35738);
nor U42406 (N_42406,N_39384,N_38805);
or U42407 (N_42407,N_37353,N_35202);
nor U42408 (N_42408,N_37975,N_35762);
nor U42409 (N_42409,N_35631,N_35174);
nand U42410 (N_42410,N_36233,N_39731);
or U42411 (N_42411,N_39060,N_38295);
or U42412 (N_42412,N_37509,N_36692);
nand U42413 (N_42413,N_37317,N_36859);
nor U42414 (N_42414,N_37316,N_39714);
and U42415 (N_42415,N_35015,N_35701);
and U42416 (N_42416,N_38328,N_39368);
or U42417 (N_42417,N_38936,N_36470);
nand U42418 (N_42418,N_38221,N_36979);
nand U42419 (N_42419,N_36007,N_37015);
and U42420 (N_42420,N_35635,N_36169);
xor U42421 (N_42421,N_38640,N_38043);
or U42422 (N_42422,N_38011,N_38876);
or U42423 (N_42423,N_36819,N_37238);
and U42424 (N_42424,N_39972,N_37667);
and U42425 (N_42425,N_35673,N_35712);
nand U42426 (N_42426,N_35587,N_37689);
or U42427 (N_42427,N_38615,N_36418);
nand U42428 (N_42428,N_39109,N_38943);
nor U42429 (N_42429,N_38460,N_38830);
xor U42430 (N_42430,N_35574,N_36949);
nand U42431 (N_42431,N_37597,N_35254);
or U42432 (N_42432,N_35632,N_38825);
and U42433 (N_42433,N_39486,N_36172);
nor U42434 (N_42434,N_38529,N_38494);
and U42435 (N_42435,N_39041,N_35325);
and U42436 (N_42436,N_37742,N_35154);
nor U42437 (N_42437,N_36562,N_39132);
and U42438 (N_42438,N_39755,N_39261);
nor U42439 (N_42439,N_36587,N_38783);
and U42440 (N_42440,N_36898,N_38132);
and U42441 (N_42441,N_35549,N_39760);
or U42442 (N_42442,N_38948,N_36998);
nor U42443 (N_42443,N_36437,N_35407);
nand U42444 (N_42444,N_38919,N_35960);
and U42445 (N_42445,N_38714,N_37250);
nor U42446 (N_42446,N_35956,N_38247);
nor U42447 (N_42447,N_37106,N_35757);
nor U42448 (N_42448,N_35470,N_35963);
or U42449 (N_42449,N_35465,N_35806);
and U42450 (N_42450,N_38907,N_39015);
nand U42451 (N_42451,N_38694,N_38707);
or U42452 (N_42452,N_36070,N_36747);
nor U42453 (N_42453,N_38584,N_35437);
or U42454 (N_42454,N_37356,N_37988);
nor U42455 (N_42455,N_38530,N_39412);
nand U42456 (N_42456,N_39344,N_39884);
or U42457 (N_42457,N_37161,N_36426);
nand U42458 (N_42458,N_38476,N_35073);
nand U42459 (N_42459,N_38729,N_38243);
nor U42460 (N_42460,N_38354,N_35755);
and U42461 (N_42461,N_37333,N_37698);
or U42462 (N_42462,N_36292,N_35444);
nor U42463 (N_42463,N_37304,N_36029);
xnor U42464 (N_42464,N_37552,N_38539);
or U42465 (N_42465,N_38008,N_37302);
nand U42466 (N_42466,N_39473,N_36644);
nor U42467 (N_42467,N_35915,N_35082);
nand U42468 (N_42468,N_37014,N_35796);
nor U42469 (N_42469,N_36995,N_38775);
and U42470 (N_42470,N_38242,N_38070);
nand U42471 (N_42471,N_35080,N_38903);
and U42472 (N_42472,N_37120,N_39213);
nor U42473 (N_42473,N_36463,N_35969);
and U42474 (N_42474,N_36021,N_35144);
nand U42475 (N_42475,N_39819,N_39965);
nand U42476 (N_42476,N_37588,N_36733);
nor U42477 (N_42477,N_38320,N_36961);
and U42478 (N_42478,N_35586,N_36270);
nor U42479 (N_42479,N_38624,N_38411);
nand U42480 (N_42480,N_38147,N_36525);
and U42481 (N_42481,N_39894,N_35032);
or U42482 (N_42482,N_38281,N_36476);
and U42483 (N_42483,N_38958,N_38124);
nand U42484 (N_42484,N_38891,N_38071);
nand U42485 (N_42485,N_38117,N_37009);
nand U42486 (N_42486,N_38290,N_36377);
or U42487 (N_42487,N_36341,N_35475);
or U42488 (N_42488,N_36676,N_35351);
or U42489 (N_42489,N_38570,N_36568);
or U42490 (N_42490,N_37013,N_38537);
and U42491 (N_42491,N_38585,N_36741);
nor U42492 (N_42492,N_35846,N_39653);
xor U42493 (N_42493,N_39525,N_37720);
nor U42494 (N_42494,N_39226,N_39596);
nor U42495 (N_42495,N_35661,N_39704);
nor U42496 (N_42496,N_35897,N_39195);
or U42497 (N_42497,N_37092,N_38410);
or U42498 (N_42498,N_39125,N_38050);
nand U42499 (N_42499,N_37969,N_39881);
and U42500 (N_42500,N_35436,N_38256);
or U42501 (N_42501,N_36660,N_36184);
and U42502 (N_42502,N_35042,N_35206);
nand U42503 (N_42503,N_39484,N_38864);
xnor U42504 (N_42504,N_39455,N_37773);
nand U42505 (N_42505,N_36097,N_35836);
nand U42506 (N_42506,N_38451,N_38349);
nor U42507 (N_42507,N_35450,N_39358);
nand U42508 (N_42508,N_35001,N_37567);
or U42509 (N_42509,N_35267,N_37587);
nor U42510 (N_42510,N_35917,N_35208);
nor U42511 (N_42511,N_37816,N_38492);
nor U42512 (N_42512,N_36488,N_37288);
or U42513 (N_42513,N_35057,N_36345);
and U42514 (N_42514,N_36496,N_39839);
xor U42515 (N_42515,N_35370,N_38727);
or U42516 (N_42516,N_35564,N_39424);
and U42517 (N_42517,N_37840,N_36790);
and U42518 (N_42518,N_37518,N_39460);
and U42519 (N_42519,N_35130,N_38965);
nor U42520 (N_42520,N_39795,N_39807);
or U42521 (N_42521,N_38207,N_39693);
nor U42522 (N_42522,N_36450,N_38069);
or U42523 (N_42523,N_38706,N_38485);
or U42524 (N_42524,N_39561,N_39764);
or U42525 (N_42525,N_36843,N_35810);
or U42526 (N_42526,N_36919,N_38713);
nand U42527 (N_42527,N_35311,N_36176);
and U42528 (N_42528,N_39914,N_36542);
or U42529 (N_42529,N_35976,N_35679);
xnor U42530 (N_42530,N_38187,N_35324);
and U42531 (N_42531,N_35134,N_39639);
nand U42532 (N_42532,N_38521,N_35836);
nor U42533 (N_42533,N_37979,N_36344);
or U42534 (N_42534,N_37520,N_39203);
nand U42535 (N_42535,N_35529,N_36869);
nor U42536 (N_42536,N_37307,N_36047);
nor U42537 (N_42537,N_39561,N_36670);
nor U42538 (N_42538,N_39987,N_38048);
and U42539 (N_42539,N_38698,N_38342);
and U42540 (N_42540,N_39308,N_36279);
nand U42541 (N_42541,N_36190,N_38706);
and U42542 (N_42542,N_37020,N_35201);
or U42543 (N_42543,N_39416,N_36307);
xor U42544 (N_42544,N_39062,N_36306);
nor U42545 (N_42545,N_37495,N_38247);
nor U42546 (N_42546,N_35082,N_37723);
nor U42547 (N_42547,N_37836,N_36150);
and U42548 (N_42548,N_39833,N_36225);
or U42549 (N_42549,N_39655,N_39055);
nand U42550 (N_42550,N_38056,N_37189);
nand U42551 (N_42551,N_37927,N_36517);
nor U42552 (N_42552,N_37649,N_35250);
or U42553 (N_42553,N_39973,N_38729);
and U42554 (N_42554,N_37084,N_38615);
or U42555 (N_42555,N_38112,N_36596);
xnor U42556 (N_42556,N_38536,N_37851);
or U42557 (N_42557,N_36085,N_36339);
and U42558 (N_42558,N_39560,N_39131);
and U42559 (N_42559,N_36389,N_39572);
nand U42560 (N_42560,N_39903,N_36211);
nand U42561 (N_42561,N_37650,N_38146);
or U42562 (N_42562,N_35268,N_35596);
or U42563 (N_42563,N_38132,N_37537);
nor U42564 (N_42564,N_37694,N_39125);
nand U42565 (N_42565,N_36003,N_39656);
or U42566 (N_42566,N_39908,N_37181);
xor U42567 (N_42567,N_38260,N_36869);
and U42568 (N_42568,N_36529,N_36017);
nand U42569 (N_42569,N_39880,N_37358);
nor U42570 (N_42570,N_36178,N_35604);
nand U42571 (N_42571,N_39385,N_39131);
or U42572 (N_42572,N_36421,N_39800);
xor U42573 (N_42573,N_35148,N_39707);
or U42574 (N_42574,N_37403,N_36039);
nor U42575 (N_42575,N_37427,N_38218);
nor U42576 (N_42576,N_35545,N_35464);
nand U42577 (N_42577,N_35118,N_38235);
or U42578 (N_42578,N_38746,N_35009);
nand U42579 (N_42579,N_39133,N_39591);
nand U42580 (N_42580,N_38780,N_37816);
nor U42581 (N_42581,N_38061,N_38156);
nand U42582 (N_42582,N_36833,N_35946);
and U42583 (N_42583,N_36079,N_39551);
nor U42584 (N_42584,N_39199,N_39896);
nor U42585 (N_42585,N_39822,N_35928);
nor U42586 (N_42586,N_36520,N_37445);
xnor U42587 (N_42587,N_36082,N_37924);
nor U42588 (N_42588,N_38462,N_35850);
or U42589 (N_42589,N_35195,N_37893);
and U42590 (N_42590,N_35365,N_38426);
and U42591 (N_42591,N_39174,N_38400);
nand U42592 (N_42592,N_36833,N_38422);
nor U42593 (N_42593,N_38162,N_37518);
or U42594 (N_42594,N_39560,N_37738);
nor U42595 (N_42595,N_38910,N_35463);
nand U42596 (N_42596,N_39456,N_39736);
nor U42597 (N_42597,N_37308,N_35103);
nand U42598 (N_42598,N_36489,N_36905);
or U42599 (N_42599,N_37967,N_39425);
and U42600 (N_42600,N_36326,N_35222);
nand U42601 (N_42601,N_38605,N_37335);
and U42602 (N_42602,N_39393,N_37185);
xnor U42603 (N_42603,N_39279,N_36749);
and U42604 (N_42604,N_37429,N_39078);
or U42605 (N_42605,N_35208,N_38483);
or U42606 (N_42606,N_38780,N_39057);
xnor U42607 (N_42607,N_35988,N_36260);
or U42608 (N_42608,N_35180,N_39702);
nand U42609 (N_42609,N_37118,N_37302);
and U42610 (N_42610,N_36047,N_35935);
or U42611 (N_42611,N_35576,N_35044);
xnor U42612 (N_42612,N_36661,N_36244);
nand U42613 (N_42613,N_36148,N_35740);
or U42614 (N_42614,N_37495,N_37411);
nand U42615 (N_42615,N_39544,N_38706);
or U42616 (N_42616,N_39470,N_36523);
nor U42617 (N_42617,N_38981,N_37802);
and U42618 (N_42618,N_38475,N_37233);
and U42619 (N_42619,N_35283,N_37826);
nor U42620 (N_42620,N_35237,N_35158);
nor U42621 (N_42621,N_38024,N_38811);
nor U42622 (N_42622,N_35880,N_36265);
nor U42623 (N_42623,N_38629,N_39558);
and U42624 (N_42624,N_35274,N_36810);
and U42625 (N_42625,N_36978,N_35798);
or U42626 (N_42626,N_37691,N_39277);
nor U42627 (N_42627,N_38249,N_36359);
nand U42628 (N_42628,N_39214,N_38564);
nand U42629 (N_42629,N_39597,N_35063);
nand U42630 (N_42630,N_36458,N_38171);
nor U42631 (N_42631,N_36737,N_37495);
nand U42632 (N_42632,N_35862,N_38182);
or U42633 (N_42633,N_39404,N_35349);
nand U42634 (N_42634,N_38525,N_37023);
or U42635 (N_42635,N_35306,N_35608);
xor U42636 (N_42636,N_37794,N_36146);
or U42637 (N_42637,N_36903,N_37414);
nand U42638 (N_42638,N_37591,N_38144);
nor U42639 (N_42639,N_35503,N_38836);
or U42640 (N_42640,N_39013,N_38744);
and U42641 (N_42641,N_35719,N_37313);
nor U42642 (N_42642,N_37553,N_39916);
or U42643 (N_42643,N_38380,N_37964);
and U42644 (N_42644,N_38580,N_35507);
xnor U42645 (N_42645,N_37723,N_36067);
nand U42646 (N_42646,N_37330,N_38614);
nor U42647 (N_42647,N_35359,N_37598);
nor U42648 (N_42648,N_39816,N_38378);
and U42649 (N_42649,N_37152,N_39000);
and U42650 (N_42650,N_35514,N_39316);
nor U42651 (N_42651,N_39263,N_39218);
nand U42652 (N_42652,N_38776,N_38076);
nand U42653 (N_42653,N_38431,N_37544);
nor U42654 (N_42654,N_38530,N_37989);
nor U42655 (N_42655,N_37849,N_39700);
nor U42656 (N_42656,N_36456,N_38500);
and U42657 (N_42657,N_37180,N_36661);
and U42658 (N_42658,N_37879,N_37159);
xnor U42659 (N_42659,N_39334,N_38294);
nand U42660 (N_42660,N_35697,N_38041);
nor U42661 (N_42661,N_37922,N_35163);
nor U42662 (N_42662,N_37184,N_39860);
and U42663 (N_42663,N_35919,N_39040);
nand U42664 (N_42664,N_35708,N_35581);
and U42665 (N_42665,N_36616,N_37662);
nor U42666 (N_42666,N_39620,N_35130);
nor U42667 (N_42667,N_39125,N_39331);
nand U42668 (N_42668,N_35339,N_39114);
nor U42669 (N_42669,N_35536,N_36259);
nand U42670 (N_42670,N_38885,N_38212);
nand U42671 (N_42671,N_36933,N_35375);
nor U42672 (N_42672,N_38877,N_38629);
nor U42673 (N_42673,N_38381,N_38730);
nor U42674 (N_42674,N_36087,N_37357);
nor U42675 (N_42675,N_38883,N_39689);
or U42676 (N_42676,N_39271,N_35914);
and U42677 (N_42677,N_35678,N_39593);
nor U42678 (N_42678,N_35496,N_39068);
xor U42679 (N_42679,N_38489,N_36744);
nor U42680 (N_42680,N_37565,N_36608);
and U42681 (N_42681,N_37500,N_38546);
nor U42682 (N_42682,N_35900,N_36206);
nor U42683 (N_42683,N_37851,N_38245);
and U42684 (N_42684,N_37579,N_35113);
nand U42685 (N_42685,N_39201,N_36179);
and U42686 (N_42686,N_38757,N_35222);
nor U42687 (N_42687,N_35129,N_37421);
nor U42688 (N_42688,N_35625,N_39052);
nand U42689 (N_42689,N_37947,N_35265);
nor U42690 (N_42690,N_35182,N_36111);
xor U42691 (N_42691,N_35252,N_35411);
nor U42692 (N_42692,N_37847,N_39190);
nor U42693 (N_42693,N_37895,N_39792);
and U42694 (N_42694,N_38461,N_37265);
nand U42695 (N_42695,N_38021,N_35968);
or U42696 (N_42696,N_38332,N_35790);
nand U42697 (N_42697,N_37781,N_39070);
and U42698 (N_42698,N_35247,N_36206);
or U42699 (N_42699,N_36965,N_35147);
or U42700 (N_42700,N_39177,N_35966);
and U42701 (N_42701,N_35284,N_38665);
or U42702 (N_42702,N_38948,N_37348);
nor U42703 (N_42703,N_38351,N_39303);
or U42704 (N_42704,N_37706,N_39873);
nor U42705 (N_42705,N_38940,N_38617);
or U42706 (N_42706,N_39807,N_36023);
and U42707 (N_42707,N_35492,N_37633);
and U42708 (N_42708,N_39001,N_35757);
and U42709 (N_42709,N_38413,N_35804);
and U42710 (N_42710,N_38762,N_39098);
nor U42711 (N_42711,N_38453,N_35430);
nor U42712 (N_42712,N_39192,N_38910);
or U42713 (N_42713,N_39745,N_35911);
and U42714 (N_42714,N_37247,N_35951);
nor U42715 (N_42715,N_37355,N_37302);
xnor U42716 (N_42716,N_37338,N_36708);
and U42717 (N_42717,N_36746,N_35449);
nor U42718 (N_42718,N_36137,N_39168);
xor U42719 (N_42719,N_38233,N_35228);
or U42720 (N_42720,N_35840,N_39950);
nand U42721 (N_42721,N_39614,N_37143);
and U42722 (N_42722,N_39246,N_38780);
nor U42723 (N_42723,N_39338,N_38998);
and U42724 (N_42724,N_36513,N_35093);
and U42725 (N_42725,N_37493,N_37608);
or U42726 (N_42726,N_37883,N_39269);
nand U42727 (N_42727,N_36586,N_37825);
nand U42728 (N_42728,N_39628,N_36197);
or U42729 (N_42729,N_36298,N_39866);
nand U42730 (N_42730,N_39409,N_38512);
and U42731 (N_42731,N_39170,N_36115);
xor U42732 (N_42732,N_38161,N_39553);
nor U42733 (N_42733,N_38535,N_36047);
nand U42734 (N_42734,N_36430,N_38821);
or U42735 (N_42735,N_39095,N_37821);
or U42736 (N_42736,N_35882,N_38460);
and U42737 (N_42737,N_35234,N_38407);
nand U42738 (N_42738,N_37758,N_36402);
nor U42739 (N_42739,N_36308,N_35839);
and U42740 (N_42740,N_39953,N_36942);
nand U42741 (N_42741,N_35789,N_37852);
xnor U42742 (N_42742,N_36431,N_38850);
and U42743 (N_42743,N_35667,N_38153);
and U42744 (N_42744,N_37568,N_37345);
xor U42745 (N_42745,N_37205,N_35610);
or U42746 (N_42746,N_37998,N_38285);
nand U42747 (N_42747,N_36083,N_37631);
nand U42748 (N_42748,N_38426,N_39547);
nor U42749 (N_42749,N_39191,N_36478);
and U42750 (N_42750,N_35338,N_35256);
nand U42751 (N_42751,N_36268,N_36474);
and U42752 (N_42752,N_39028,N_37492);
or U42753 (N_42753,N_39246,N_39658);
or U42754 (N_42754,N_38741,N_37029);
nand U42755 (N_42755,N_37802,N_39158);
and U42756 (N_42756,N_35271,N_38947);
nor U42757 (N_42757,N_39012,N_38973);
xor U42758 (N_42758,N_36454,N_35083);
and U42759 (N_42759,N_37472,N_38775);
or U42760 (N_42760,N_39792,N_38017);
nor U42761 (N_42761,N_36550,N_36251);
nor U42762 (N_42762,N_36063,N_35978);
nor U42763 (N_42763,N_35446,N_37076);
nor U42764 (N_42764,N_38146,N_36371);
nand U42765 (N_42765,N_37759,N_38798);
nand U42766 (N_42766,N_35979,N_36838);
or U42767 (N_42767,N_39008,N_35249);
and U42768 (N_42768,N_36223,N_39754);
nor U42769 (N_42769,N_39762,N_35983);
and U42770 (N_42770,N_39434,N_38349);
and U42771 (N_42771,N_39747,N_37779);
nand U42772 (N_42772,N_36153,N_35532);
nand U42773 (N_42773,N_39375,N_36806);
or U42774 (N_42774,N_36193,N_36012);
or U42775 (N_42775,N_38201,N_35622);
or U42776 (N_42776,N_37192,N_37743);
nand U42777 (N_42777,N_36934,N_36829);
xnor U42778 (N_42778,N_37034,N_35764);
nor U42779 (N_42779,N_37745,N_35939);
and U42780 (N_42780,N_39919,N_39004);
nand U42781 (N_42781,N_37061,N_35316);
xor U42782 (N_42782,N_39911,N_36674);
or U42783 (N_42783,N_39366,N_36952);
and U42784 (N_42784,N_35124,N_36283);
or U42785 (N_42785,N_35004,N_36728);
nand U42786 (N_42786,N_37884,N_36914);
xnor U42787 (N_42787,N_38254,N_37680);
nand U42788 (N_42788,N_36787,N_39639);
or U42789 (N_42789,N_36605,N_36784);
and U42790 (N_42790,N_36592,N_38664);
or U42791 (N_42791,N_37607,N_37026);
nor U42792 (N_42792,N_38353,N_39317);
nor U42793 (N_42793,N_35672,N_35829);
nand U42794 (N_42794,N_37532,N_39450);
nand U42795 (N_42795,N_35160,N_37488);
or U42796 (N_42796,N_39414,N_38279);
nor U42797 (N_42797,N_39712,N_38901);
nor U42798 (N_42798,N_39309,N_38016);
or U42799 (N_42799,N_36152,N_39188);
and U42800 (N_42800,N_39335,N_36932);
nor U42801 (N_42801,N_39748,N_39837);
nand U42802 (N_42802,N_36740,N_35655);
nor U42803 (N_42803,N_39182,N_39074);
or U42804 (N_42804,N_39978,N_36401);
and U42805 (N_42805,N_38356,N_38606);
nand U42806 (N_42806,N_37107,N_39239);
and U42807 (N_42807,N_36291,N_39487);
and U42808 (N_42808,N_36802,N_38778);
and U42809 (N_42809,N_37685,N_38946);
or U42810 (N_42810,N_39767,N_35828);
nand U42811 (N_42811,N_35612,N_38976);
and U42812 (N_42812,N_37887,N_35454);
or U42813 (N_42813,N_39873,N_36415);
nand U42814 (N_42814,N_35414,N_36055);
xor U42815 (N_42815,N_38908,N_36986);
nor U42816 (N_42816,N_37296,N_38891);
or U42817 (N_42817,N_35457,N_36640);
nor U42818 (N_42818,N_36279,N_35088);
nor U42819 (N_42819,N_37534,N_35526);
or U42820 (N_42820,N_39990,N_37648);
nor U42821 (N_42821,N_36554,N_38488);
xor U42822 (N_42822,N_37540,N_36073);
nor U42823 (N_42823,N_37891,N_35843);
or U42824 (N_42824,N_36312,N_39362);
nand U42825 (N_42825,N_36276,N_39321);
or U42826 (N_42826,N_36148,N_35996);
nor U42827 (N_42827,N_36865,N_35674);
nand U42828 (N_42828,N_35887,N_38453);
and U42829 (N_42829,N_38826,N_35083);
xnor U42830 (N_42830,N_35069,N_36467);
and U42831 (N_42831,N_35803,N_36044);
and U42832 (N_42832,N_39617,N_35850);
or U42833 (N_42833,N_38102,N_39075);
or U42834 (N_42834,N_36989,N_38878);
nand U42835 (N_42835,N_36395,N_37021);
and U42836 (N_42836,N_37493,N_37886);
nand U42837 (N_42837,N_38776,N_36765);
or U42838 (N_42838,N_39110,N_35666);
and U42839 (N_42839,N_35827,N_39446);
or U42840 (N_42840,N_38679,N_38599);
or U42841 (N_42841,N_35050,N_37988);
or U42842 (N_42842,N_36162,N_38932);
nor U42843 (N_42843,N_37186,N_36037);
xor U42844 (N_42844,N_36345,N_36852);
nand U42845 (N_42845,N_37201,N_37743);
or U42846 (N_42846,N_37783,N_39786);
xor U42847 (N_42847,N_38160,N_39960);
or U42848 (N_42848,N_39545,N_39227);
xor U42849 (N_42849,N_35366,N_37623);
nand U42850 (N_42850,N_39370,N_38094);
or U42851 (N_42851,N_35675,N_35757);
and U42852 (N_42852,N_37768,N_36364);
or U42853 (N_42853,N_37521,N_37300);
or U42854 (N_42854,N_35671,N_39372);
nor U42855 (N_42855,N_35853,N_38409);
nor U42856 (N_42856,N_39982,N_39914);
nor U42857 (N_42857,N_37261,N_37686);
and U42858 (N_42858,N_36862,N_38572);
and U42859 (N_42859,N_38472,N_38096);
or U42860 (N_42860,N_36962,N_38904);
nand U42861 (N_42861,N_37727,N_36297);
nor U42862 (N_42862,N_39977,N_37025);
xnor U42863 (N_42863,N_36318,N_37889);
and U42864 (N_42864,N_36387,N_38644);
and U42865 (N_42865,N_35079,N_39686);
or U42866 (N_42866,N_35986,N_35439);
or U42867 (N_42867,N_37627,N_35490);
nand U42868 (N_42868,N_36537,N_38942);
nand U42869 (N_42869,N_37322,N_37504);
nand U42870 (N_42870,N_36979,N_36087);
nand U42871 (N_42871,N_37466,N_35736);
nor U42872 (N_42872,N_39040,N_36239);
nand U42873 (N_42873,N_35482,N_38687);
nor U42874 (N_42874,N_37223,N_36105);
nand U42875 (N_42875,N_35648,N_39337);
nand U42876 (N_42876,N_37248,N_36847);
nor U42877 (N_42877,N_38779,N_38269);
nand U42878 (N_42878,N_38109,N_36873);
xor U42879 (N_42879,N_37652,N_35244);
or U42880 (N_42880,N_35115,N_36372);
and U42881 (N_42881,N_36357,N_36837);
or U42882 (N_42882,N_37806,N_39602);
nor U42883 (N_42883,N_38185,N_39107);
nand U42884 (N_42884,N_39094,N_35823);
or U42885 (N_42885,N_36331,N_35365);
nand U42886 (N_42886,N_39095,N_38787);
nor U42887 (N_42887,N_38271,N_37448);
or U42888 (N_42888,N_38730,N_39044);
and U42889 (N_42889,N_39327,N_37945);
xor U42890 (N_42890,N_38807,N_39358);
xnor U42891 (N_42891,N_35274,N_36231);
or U42892 (N_42892,N_38166,N_38169);
and U42893 (N_42893,N_38303,N_38939);
and U42894 (N_42894,N_39235,N_35064);
and U42895 (N_42895,N_37276,N_35179);
and U42896 (N_42896,N_37350,N_37209);
or U42897 (N_42897,N_38793,N_37724);
nand U42898 (N_42898,N_35988,N_39617);
and U42899 (N_42899,N_38371,N_39207);
nand U42900 (N_42900,N_36812,N_39088);
nand U42901 (N_42901,N_38753,N_37027);
nand U42902 (N_42902,N_38806,N_39666);
and U42903 (N_42903,N_35614,N_38185);
nor U42904 (N_42904,N_38990,N_37865);
nand U42905 (N_42905,N_35099,N_36101);
nor U42906 (N_42906,N_35197,N_37116);
xnor U42907 (N_42907,N_38788,N_36261);
nor U42908 (N_42908,N_39101,N_39899);
or U42909 (N_42909,N_35789,N_36015);
and U42910 (N_42910,N_39808,N_38814);
nand U42911 (N_42911,N_39100,N_36479);
or U42912 (N_42912,N_35204,N_37553);
or U42913 (N_42913,N_35286,N_38397);
nor U42914 (N_42914,N_38372,N_37431);
or U42915 (N_42915,N_35649,N_35902);
or U42916 (N_42916,N_39044,N_35178);
or U42917 (N_42917,N_39326,N_35453);
or U42918 (N_42918,N_39413,N_39050);
nand U42919 (N_42919,N_39106,N_38062);
and U42920 (N_42920,N_36566,N_36533);
xor U42921 (N_42921,N_36023,N_35198);
and U42922 (N_42922,N_35326,N_38985);
and U42923 (N_42923,N_37837,N_39594);
and U42924 (N_42924,N_36764,N_37974);
or U42925 (N_42925,N_36345,N_37827);
and U42926 (N_42926,N_38231,N_36239);
and U42927 (N_42927,N_39397,N_36037);
nor U42928 (N_42928,N_35738,N_35885);
nor U42929 (N_42929,N_37472,N_35872);
or U42930 (N_42930,N_35409,N_35977);
or U42931 (N_42931,N_37139,N_37347);
nand U42932 (N_42932,N_35093,N_38692);
nor U42933 (N_42933,N_36404,N_35202);
nand U42934 (N_42934,N_39547,N_38796);
and U42935 (N_42935,N_35385,N_35158);
nand U42936 (N_42936,N_39672,N_37352);
or U42937 (N_42937,N_36938,N_38607);
xor U42938 (N_42938,N_38031,N_35012);
or U42939 (N_42939,N_35900,N_37471);
nor U42940 (N_42940,N_35264,N_39063);
nand U42941 (N_42941,N_36908,N_35878);
xnor U42942 (N_42942,N_36900,N_39510);
or U42943 (N_42943,N_35685,N_39441);
or U42944 (N_42944,N_35397,N_37995);
or U42945 (N_42945,N_38260,N_38008);
or U42946 (N_42946,N_37464,N_38085);
or U42947 (N_42947,N_38762,N_35753);
xnor U42948 (N_42948,N_35168,N_38362);
nor U42949 (N_42949,N_38855,N_35520);
or U42950 (N_42950,N_37779,N_36718);
xnor U42951 (N_42951,N_37590,N_39461);
nor U42952 (N_42952,N_37802,N_35337);
or U42953 (N_42953,N_35765,N_38641);
nor U42954 (N_42954,N_38916,N_38005);
and U42955 (N_42955,N_35911,N_38006);
nor U42956 (N_42956,N_37948,N_35065);
nor U42957 (N_42957,N_36324,N_36239);
nor U42958 (N_42958,N_37180,N_39245);
and U42959 (N_42959,N_38263,N_36114);
nand U42960 (N_42960,N_38480,N_37888);
nor U42961 (N_42961,N_38404,N_36744);
or U42962 (N_42962,N_36377,N_39082);
or U42963 (N_42963,N_35819,N_38334);
and U42964 (N_42964,N_38898,N_37167);
nor U42965 (N_42965,N_38826,N_35523);
or U42966 (N_42966,N_38255,N_38400);
nor U42967 (N_42967,N_38775,N_36039);
xor U42968 (N_42968,N_37872,N_38017);
nand U42969 (N_42969,N_35433,N_35681);
or U42970 (N_42970,N_39171,N_37723);
xor U42971 (N_42971,N_35064,N_38543);
xnor U42972 (N_42972,N_38976,N_36949);
and U42973 (N_42973,N_35648,N_39032);
or U42974 (N_42974,N_38516,N_35032);
and U42975 (N_42975,N_36807,N_39923);
and U42976 (N_42976,N_39026,N_39761);
nor U42977 (N_42977,N_38934,N_38978);
xor U42978 (N_42978,N_39852,N_39850);
nand U42979 (N_42979,N_37049,N_36875);
nor U42980 (N_42980,N_35458,N_38730);
xnor U42981 (N_42981,N_35840,N_38917);
and U42982 (N_42982,N_35558,N_39862);
nand U42983 (N_42983,N_39015,N_39020);
and U42984 (N_42984,N_35917,N_35511);
or U42985 (N_42985,N_39833,N_36440);
or U42986 (N_42986,N_37836,N_37458);
and U42987 (N_42987,N_37682,N_35630);
xor U42988 (N_42988,N_35217,N_39221);
nor U42989 (N_42989,N_39709,N_39496);
xnor U42990 (N_42990,N_39163,N_38600);
nor U42991 (N_42991,N_37203,N_38403);
nand U42992 (N_42992,N_36114,N_38667);
nor U42993 (N_42993,N_38504,N_37027);
xnor U42994 (N_42994,N_35166,N_39185);
nor U42995 (N_42995,N_39653,N_37826);
and U42996 (N_42996,N_35735,N_38708);
xor U42997 (N_42997,N_37432,N_35666);
or U42998 (N_42998,N_39387,N_39759);
nand U42999 (N_42999,N_38578,N_36234);
or U43000 (N_43000,N_38395,N_39457);
nor U43001 (N_43001,N_38921,N_39828);
or U43002 (N_43002,N_35359,N_36716);
and U43003 (N_43003,N_38107,N_36976);
and U43004 (N_43004,N_36674,N_36352);
or U43005 (N_43005,N_37746,N_39387);
nor U43006 (N_43006,N_39440,N_37848);
nand U43007 (N_43007,N_39477,N_38558);
and U43008 (N_43008,N_36120,N_39115);
and U43009 (N_43009,N_36912,N_36302);
and U43010 (N_43010,N_35362,N_38720);
and U43011 (N_43011,N_38524,N_39581);
nand U43012 (N_43012,N_35449,N_39656);
or U43013 (N_43013,N_38010,N_36484);
and U43014 (N_43014,N_36947,N_38692);
xnor U43015 (N_43015,N_38012,N_36622);
nor U43016 (N_43016,N_38686,N_39877);
xor U43017 (N_43017,N_36628,N_39631);
nor U43018 (N_43018,N_37164,N_36179);
nor U43019 (N_43019,N_37951,N_35517);
nor U43020 (N_43020,N_37964,N_35963);
nor U43021 (N_43021,N_37901,N_39642);
and U43022 (N_43022,N_38816,N_37880);
nor U43023 (N_43023,N_38206,N_36742);
nor U43024 (N_43024,N_35132,N_39557);
and U43025 (N_43025,N_37690,N_35893);
nand U43026 (N_43026,N_38194,N_35713);
or U43027 (N_43027,N_37099,N_35244);
or U43028 (N_43028,N_39340,N_39895);
xnor U43029 (N_43029,N_39419,N_36935);
nand U43030 (N_43030,N_37243,N_35723);
and U43031 (N_43031,N_35807,N_35309);
nor U43032 (N_43032,N_36068,N_39624);
and U43033 (N_43033,N_35766,N_35160);
and U43034 (N_43034,N_35495,N_36115);
or U43035 (N_43035,N_39511,N_37485);
or U43036 (N_43036,N_37814,N_35284);
nor U43037 (N_43037,N_37748,N_35755);
nand U43038 (N_43038,N_37757,N_36137);
nand U43039 (N_43039,N_38456,N_38544);
nand U43040 (N_43040,N_37712,N_38524);
and U43041 (N_43041,N_36616,N_38061);
nand U43042 (N_43042,N_36531,N_37531);
xnor U43043 (N_43043,N_39101,N_35709);
and U43044 (N_43044,N_36751,N_35572);
nand U43045 (N_43045,N_38523,N_39053);
nor U43046 (N_43046,N_35581,N_37621);
or U43047 (N_43047,N_39462,N_35240);
nor U43048 (N_43048,N_38439,N_37535);
nand U43049 (N_43049,N_35856,N_36515);
xor U43050 (N_43050,N_36477,N_37414);
nor U43051 (N_43051,N_35263,N_36879);
and U43052 (N_43052,N_35997,N_36585);
nor U43053 (N_43053,N_35189,N_35128);
and U43054 (N_43054,N_36024,N_36627);
xor U43055 (N_43055,N_36829,N_36448);
or U43056 (N_43056,N_36381,N_37417);
nand U43057 (N_43057,N_38803,N_35466);
nand U43058 (N_43058,N_39726,N_38467);
or U43059 (N_43059,N_37113,N_38435);
nand U43060 (N_43060,N_39717,N_39939);
nor U43061 (N_43061,N_35479,N_36201);
nor U43062 (N_43062,N_38797,N_39214);
nand U43063 (N_43063,N_37089,N_36513);
or U43064 (N_43064,N_39732,N_35862);
nor U43065 (N_43065,N_37013,N_35962);
or U43066 (N_43066,N_35755,N_36086);
and U43067 (N_43067,N_38056,N_39484);
nor U43068 (N_43068,N_36055,N_38871);
nor U43069 (N_43069,N_36652,N_37873);
nor U43070 (N_43070,N_37584,N_36473);
and U43071 (N_43071,N_37020,N_38877);
or U43072 (N_43072,N_37440,N_37290);
nor U43073 (N_43073,N_39282,N_38943);
or U43074 (N_43074,N_36512,N_39045);
or U43075 (N_43075,N_36458,N_36528);
and U43076 (N_43076,N_39770,N_38662);
nor U43077 (N_43077,N_35132,N_35084);
nand U43078 (N_43078,N_37867,N_35754);
nor U43079 (N_43079,N_38625,N_36378);
or U43080 (N_43080,N_38455,N_36695);
or U43081 (N_43081,N_37817,N_38359);
nor U43082 (N_43082,N_37019,N_36500);
nor U43083 (N_43083,N_39242,N_39918);
or U43084 (N_43084,N_35958,N_39106);
nor U43085 (N_43085,N_36467,N_38706);
xor U43086 (N_43086,N_39882,N_39496);
or U43087 (N_43087,N_39240,N_37971);
nor U43088 (N_43088,N_38329,N_36587);
nor U43089 (N_43089,N_36768,N_36591);
nor U43090 (N_43090,N_37679,N_39779);
nor U43091 (N_43091,N_37332,N_35862);
nor U43092 (N_43092,N_35962,N_37721);
nor U43093 (N_43093,N_37689,N_39263);
and U43094 (N_43094,N_35453,N_38277);
nor U43095 (N_43095,N_38396,N_39380);
and U43096 (N_43096,N_39471,N_35696);
or U43097 (N_43097,N_37124,N_36310);
nand U43098 (N_43098,N_39327,N_39333);
nor U43099 (N_43099,N_38109,N_36913);
or U43100 (N_43100,N_36619,N_35379);
and U43101 (N_43101,N_36324,N_38578);
or U43102 (N_43102,N_39964,N_36198);
nand U43103 (N_43103,N_38468,N_35448);
nand U43104 (N_43104,N_36574,N_39347);
nor U43105 (N_43105,N_37735,N_39111);
or U43106 (N_43106,N_36737,N_37550);
or U43107 (N_43107,N_38888,N_36105);
or U43108 (N_43108,N_35152,N_35214);
and U43109 (N_43109,N_35343,N_38413);
nand U43110 (N_43110,N_39907,N_38222);
and U43111 (N_43111,N_38743,N_35690);
nand U43112 (N_43112,N_37123,N_37208);
nand U43113 (N_43113,N_37227,N_39630);
nand U43114 (N_43114,N_39462,N_36230);
or U43115 (N_43115,N_35986,N_38616);
or U43116 (N_43116,N_35166,N_36535);
and U43117 (N_43117,N_39112,N_37703);
or U43118 (N_43118,N_37490,N_38167);
or U43119 (N_43119,N_39843,N_39459);
nand U43120 (N_43120,N_39437,N_37176);
and U43121 (N_43121,N_35250,N_35443);
nand U43122 (N_43122,N_37251,N_38895);
nor U43123 (N_43123,N_39432,N_36420);
nand U43124 (N_43124,N_37402,N_35762);
and U43125 (N_43125,N_39345,N_37959);
nor U43126 (N_43126,N_39167,N_39706);
or U43127 (N_43127,N_39073,N_38409);
and U43128 (N_43128,N_35092,N_36780);
and U43129 (N_43129,N_39899,N_35620);
xor U43130 (N_43130,N_37629,N_35383);
nand U43131 (N_43131,N_35538,N_35235);
nand U43132 (N_43132,N_39334,N_35475);
or U43133 (N_43133,N_39615,N_35908);
nand U43134 (N_43134,N_36001,N_38032);
nor U43135 (N_43135,N_36406,N_39936);
or U43136 (N_43136,N_35261,N_38138);
or U43137 (N_43137,N_35354,N_38430);
or U43138 (N_43138,N_37655,N_36571);
nand U43139 (N_43139,N_38823,N_38313);
nand U43140 (N_43140,N_36248,N_35516);
and U43141 (N_43141,N_37262,N_37101);
and U43142 (N_43142,N_37604,N_38958);
or U43143 (N_43143,N_36711,N_39872);
or U43144 (N_43144,N_36691,N_37174);
and U43145 (N_43145,N_35752,N_39487);
nand U43146 (N_43146,N_35300,N_39882);
nor U43147 (N_43147,N_35384,N_35046);
nor U43148 (N_43148,N_35416,N_39572);
nor U43149 (N_43149,N_36938,N_38999);
or U43150 (N_43150,N_38263,N_37296);
nor U43151 (N_43151,N_37335,N_39148);
nand U43152 (N_43152,N_36337,N_36865);
or U43153 (N_43153,N_38224,N_39417);
nor U43154 (N_43154,N_39377,N_36226);
or U43155 (N_43155,N_37611,N_37838);
nor U43156 (N_43156,N_36553,N_39208);
and U43157 (N_43157,N_37281,N_36684);
nor U43158 (N_43158,N_39347,N_36704);
nor U43159 (N_43159,N_38601,N_36505);
nor U43160 (N_43160,N_39284,N_36206);
nor U43161 (N_43161,N_39185,N_37907);
or U43162 (N_43162,N_38478,N_37335);
nand U43163 (N_43163,N_35796,N_36450);
or U43164 (N_43164,N_36927,N_39944);
nor U43165 (N_43165,N_35718,N_39063);
xnor U43166 (N_43166,N_39951,N_38237);
nor U43167 (N_43167,N_37597,N_37200);
xor U43168 (N_43168,N_36420,N_39965);
or U43169 (N_43169,N_39164,N_35367);
xor U43170 (N_43170,N_37270,N_35809);
nand U43171 (N_43171,N_39579,N_39064);
nand U43172 (N_43172,N_37071,N_38634);
xnor U43173 (N_43173,N_39145,N_39427);
nand U43174 (N_43174,N_38072,N_37456);
nand U43175 (N_43175,N_38508,N_39753);
nor U43176 (N_43176,N_36165,N_35202);
xnor U43177 (N_43177,N_35429,N_39622);
xor U43178 (N_43178,N_38522,N_39951);
or U43179 (N_43179,N_38276,N_35034);
and U43180 (N_43180,N_39147,N_35920);
or U43181 (N_43181,N_37063,N_35104);
nor U43182 (N_43182,N_38247,N_37976);
and U43183 (N_43183,N_39897,N_37168);
or U43184 (N_43184,N_38807,N_39367);
or U43185 (N_43185,N_39181,N_36019);
and U43186 (N_43186,N_37800,N_36065);
nor U43187 (N_43187,N_35789,N_37772);
nand U43188 (N_43188,N_37851,N_35436);
or U43189 (N_43189,N_37313,N_37674);
xnor U43190 (N_43190,N_38564,N_36562);
xor U43191 (N_43191,N_38028,N_36624);
xnor U43192 (N_43192,N_35707,N_38708);
or U43193 (N_43193,N_35991,N_37827);
or U43194 (N_43194,N_35547,N_35235);
and U43195 (N_43195,N_39736,N_38422);
or U43196 (N_43196,N_35506,N_36946);
nand U43197 (N_43197,N_35231,N_36310);
or U43198 (N_43198,N_37330,N_37281);
nor U43199 (N_43199,N_36341,N_37286);
nand U43200 (N_43200,N_37129,N_38882);
nor U43201 (N_43201,N_36735,N_36740);
and U43202 (N_43202,N_35437,N_37410);
nor U43203 (N_43203,N_38736,N_36185);
nor U43204 (N_43204,N_39999,N_39129);
and U43205 (N_43205,N_37698,N_35934);
nand U43206 (N_43206,N_35447,N_39888);
or U43207 (N_43207,N_39282,N_37999);
nand U43208 (N_43208,N_36124,N_35431);
or U43209 (N_43209,N_36505,N_38409);
nor U43210 (N_43210,N_37798,N_39082);
and U43211 (N_43211,N_39666,N_38409);
and U43212 (N_43212,N_37351,N_36835);
and U43213 (N_43213,N_36151,N_36435);
and U43214 (N_43214,N_38264,N_36528);
nand U43215 (N_43215,N_36764,N_38440);
nor U43216 (N_43216,N_35014,N_38265);
and U43217 (N_43217,N_37962,N_37080);
nor U43218 (N_43218,N_36094,N_38349);
and U43219 (N_43219,N_36240,N_37879);
or U43220 (N_43220,N_38983,N_37554);
or U43221 (N_43221,N_38463,N_35344);
xnor U43222 (N_43222,N_38347,N_38524);
and U43223 (N_43223,N_36862,N_35862);
xnor U43224 (N_43224,N_37967,N_36509);
xor U43225 (N_43225,N_39714,N_38258);
nor U43226 (N_43226,N_35749,N_35988);
or U43227 (N_43227,N_38044,N_38880);
and U43228 (N_43228,N_35376,N_38616);
xor U43229 (N_43229,N_35545,N_36774);
nand U43230 (N_43230,N_36291,N_38417);
xnor U43231 (N_43231,N_39349,N_36705);
or U43232 (N_43232,N_37568,N_35845);
nand U43233 (N_43233,N_38347,N_37843);
nand U43234 (N_43234,N_39322,N_36580);
xnor U43235 (N_43235,N_36990,N_35165);
or U43236 (N_43236,N_36798,N_39360);
or U43237 (N_43237,N_37273,N_36996);
nor U43238 (N_43238,N_35881,N_36124);
or U43239 (N_43239,N_37969,N_36957);
nand U43240 (N_43240,N_37841,N_36465);
and U43241 (N_43241,N_38652,N_39973);
nand U43242 (N_43242,N_35103,N_38065);
nand U43243 (N_43243,N_39703,N_38081);
or U43244 (N_43244,N_35394,N_39427);
and U43245 (N_43245,N_37733,N_37327);
nor U43246 (N_43246,N_37913,N_35347);
nand U43247 (N_43247,N_39106,N_37808);
or U43248 (N_43248,N_35142,N_36229);
and U43249 (N_43249,N_35963,N_35724);
nand U43250 (N_43250,N_36623,N_37796);
nor U43251 (N_43251,N_39426,N_35163);
nand U43252 (N_43252,N_35662,N_37306);
or U43253 (N_43253,N_36353,N_39436);
nor U43254 (N_43254,N_35591,N_35381);
and U43255 (N_43255,N_37717,N_38216);
nand U43256 (N_43256,N_39505,N_35702);
nor U43257 (N_43257,N_39765,N_37857);
nor U43258 (N_43258,N_38739,N_36709);
nor U43259 (N_43259,N_37663,N_35423);
and U43260 (N_43260,N_36293,N_36669);
nor U43261 (N_43261,N_35854,N_36491);
and U43262 (N_43262,N_35462,N_38445);
and U43263 (N_43263,N_35580,N_37781);
nand U43264 (N_43264,N_37414,N_35549);
nand U43265 (N_43265,N_35535,N_35240);
nand U43266 (N_43266,N_39946,N_35182);
nand U43267 (N_43267,N_36932,N_35007);
or U43268 (N_43268,N_36174,N_37313);
and U43269 (N_43269,N_39357,N_37292);
or U43270 (N_43270,N_38193,N_36310);
nand U43271 (N_43271,N_38555,N_39266);
and U43272 (N_43272,N_39985,N_35888);
xnor U43273 (N_43273,N_39087,N_37231);
and U43274 (N_43274,N_38846,N_35985);
xnor U43275 (N_43275,N_39303,N_37516);
xor U43276 (N_43276,N_39230,N_38668);
or U43277 (N_43277,N_36302,N_37130);
or U43278 (N_43278,N_39924,N_36456);
nand U43279 (N_43279,N_39036,N_36833);
nor U43280 (N_43280,N_38791,N_35378);
xnor U43281 (N_43281,N_39974,N_39465);
or U43282 (N_43282,N_39964,N_36421);
nand U43283 (N_43283,N_39732,N_36193);
and U43284 (N_43284,N_37438,N_38271);
xnor U43285 (N_43285,N_35124,N_38657);
nor U43286 (N_43286,N_35917,N_38133);
nor U43287 (N_43287,N_36242,N_38196);
and U43288 (N_43288,N_39372,N_35296);
nand U43289 (N_43289,N_38569,N_37987);
or U43290 (N_43290,N_38621,N_39841);
and U43291 (N_43291,N_38930,N_37270);
nor U43292 (N_43292,N_39834,N_37716);
nand U43293 (N_43293,N_38727,N_38837);
xnor U43294 (N_43294,N_35124,N_39971);
nand U43295 (N_43295,N_39334,N_36893);
or U43296 (N_43296,N_38958,N_39187);
nor U43297 (N_43297,N_36867,N_37941);
and U43298 (N_43298,N_36506,N_36167);
and U43299 (N_43299,N_35320,N_35374);
xnor U43300 (N_43300,N_37801,N_39104);
nand U43301 (N_43301,N_39545,N_39954);
and U43302 (N_43302,N_36621,N_38230);
and U43303 (N_43303,N_38141,N_37340);
nand U43304 (N_43304,N_37580,N_39217);
nand U43305 (N_43305,N_39518,N_35763);
and U43306 (N_43306,N_38475,N_37489);
or U43307 (N_43307,N_38811,N_37482);
nor U43308 (N_43308,N_37743,N_36667);
or U43309 (N_43309,N_37387,N_35599);
and U43310 (N_43310,N_36608,N_38190);
or U43311 (N_43311,N_39994,N_38829);
nor U43312 (N_43312,N_37081,N_37813);
nor U43313 (N_43313,N_37975,N_36283);
or U43314 (N_43314,N_38070,N_35731);
or U43315 (N_43315,N_37545,N_36143);
nand U43316 (N_43316,N_35240,N_35766);
nand U43317 (N_43317,N_38776,N_35923);
or U43318 (N_43318,N_35198,N_37309);
nand U43319 (N_43319,N_37635,N_38761);
and U43320 (N_43320,N_38067,N_36334);
nand U43321 (N_43321,N_36181,N_35652);
xnor U43322 (N_43322,N_35800,N_37161);
nand U43323 (N_43323,N_37347,N_37924);
nand U43324 (N_43324,N_38709,N_38047);
and U43325 (N_43325,N_37390,N_35645);
or U43326 (N_43326,N_39922,N_35940);
nor U43327 (N_43327,N_38746,N_37591);
xor U43328 (N_43328,N_39837,N_37624);
nand U43329 (N_43329,N_37526,N_37059);
and U43330 (N_43330,N_39298,N_36714);
xor U43331 (N_43331,N_35498,N_35734);
xnor U43332 (N_43332,N_35183,N_36514);
nor U43333 (N_43333,N_38108,N_39532);
and U43334 (N_43334,N_36660,N_38579);
nand U43335 (N_43335,N_35397,N_37486);
xnor U43336 (N_43336,N_37789,N_39127);
xor U43337 (N_43337,N_37818,N_39281);
and U43338 (N_43338,N_37270,N_38583);
nor U43339 (N_43339,N_36046,N_39837);
or U43340 (N_43340,N_37392,N_36410);
nand U43341 (N_43341,N_35362,N_35334);
nor U43342 (N_43342,N_37701,N_39658);
xnor U43343 (N_43343,N_37486,N_38774);
nand U43344 (N_43344,N_39870,N_35509);
nand U43345 (N_43345,N_38273,N_39468);
nor U43346 (N_43346,N_36087,N_35495);
nand U43347 (N_43347,N_35233,N_38834);
nand U43348 (N_43348,N_37500,N_38506);
or U43349 (N_43349,N_35932,N_38282);
nor U43350 (N_43350,N_36447,N_39641);
nor U43351 (N_43351,N_35402,N_35296);
nand U43352 (N_43352,N_37776,N_38042);
and U43353 (N_43353,N_35101,N_38133);
or U43354 (N_43354,N_36036,N_37875);
and U43355 (N_43355,N_36836,N_39497);
or U43356 (N_43356,N_36460,N_37910);
nor U43357 (N_43357,N_39697,N_35632);
nand U43358 (N_43358,N_38846,N_35793);
and U43359 (N_43359,N_35534,N_35925);
or U43360 (N_43360,N_39384,N_38898);
or U43361 (N_43361,N_39496,N_35410);
nand U43362 (N_43362,N_39585,N_36635);
and U43363 (N_43363,N_37706,N_39803);
xnor U43364 (N_43364,N_36203,N_36156);
or U43365 (N_43365,N_38989,N_35160);
and U43366 (N_43366,N_37853,N_37055);
nand U43367 (N_43367,N_36091,N_36984);
nor U43368 (N_43368,N_37689,N_35734);
nor U43369 (N_43369,N_35569,N_37818);
nand U43370 (N_43370,N_38787,N_35335);
or U43371 (N_43371,N_35685,N_37759);
or U43372 (N_43372,N_39219,N_37061);
and U43373 (N_43373,N_39649,N_38059);
nand U43374 (N_43374,N_39725,N_35247);
or U43375 (N_43375,N_35991,N_36720);
nand U43376 (N_43376,N_39949,N_39387);
nand U43377 (N_43377,N_36917,N_36956);
or U43378 (N_43378,N_39425,N_36939);
or U43379 (N_43379,N_38713,N_39466);
nor U43380 (N_43380,N_36648,N_39003);
nand U43381 (N_43381,N_37753,N_39368);
xor U43382 (N_43382,N_38675,N_37039);
and U43383 (N_43383,N_37192,N_38424);
or U43384 (N_43384,N_38048,N_36208);
nor U43385 (N_43385,N_35830,N_39171);
nand U43386 (N_43386,N_39606,N_37625);
xor U43387 (N_43387,N_37754,N_36045);
and U43388 (N_43388,N_39424,N_39925);
or U43389 (N_43389,N_36763,N_37445);
nor U43390 (N_43390,N_35374,N_35377);
nor U43391 (N_43391,N_39924,N_38682);
nand U43392 (N_43392,N_37167,N_38253);
or U43393 (N_43393,N_38556,N_39311);
or U43394 (N_43394,N_37181,N_36740);
xnor U43395 (N_43395,N_37624,N_35884);
nand U43396 (N_43396,N_37046,N_35649);
or U43397 (N_43397,N_38094,N_38410);
nand U43398 (N_43398,N_36760,N_38246);
nor U43399 (N_43399,N_35768,N_37349);
and U43400 (N_43400,N_38492,N_38752);
nor U43401 (N_43401,N_37563,N_39538);
and U43402 (N_43402,N_39896,N_35233);
nor U43403 (N_43403,N_39647,N_39303);
and U43404 (N_43404,N_36387,N_38915);
or U43405 (N_43405,N_38360,N_37055);
nand U43406 (N_43406,N_37128,N_38076);
nand U43407 (N_43407,N_39727,N_39328);
nor U43408 (N_43408,N_37804,N_36069);
xor U43409 (N_43409,N_38271,N_35400);
or U43410 (N_43410,N_35777,N_38525);
nand U43411 (N_43411,N_37499,N_36465);
xor U43412 (N_43412,N_35138,N_37847);
xor U43413 (N_43413,N_35480,N_35525);
nand U43414 (N_43414,N_39290,N_38084);
nand U43415 (N_43415,N_38560,N_37674);
or U43416 (N_43416,N_38046,N_37678);
xnor U43417 (N_43417,N_35734,N_39189);
or U43418 (N_43418,N_35737,N_39990);
or U43419 (N_43419,N_35369,N_39335);
xnor U43420 (N_43420,N_39738,N_39862);
nor U43421 (N_43421,N_36819,N_37038);
nor U43422 (N_43422,N_36313,N_35725);
nand U43423 (N_43423,N_37090,N_35628);
nor U43424 (N_43424,N_37367,N_38180);
and U43425 (N_43425,N_37771,N_38957);
or U43426 (N_43426,N_35119,N_36034);
and U43427 (N_43427,N_39182,N_37837);
nand U43428 (N_43428,N_38982,N_37945);
and U43429 (N_43429,N_39013,N_37767);
or U43430 (N_43430,N_35148,N_39497);
or U43431 (N_43431,N_37814,N_38620);
nand U43432 (N_43432,N_36497,N_39518);
nand U43433 (N_43433,N_37060,N_37035);
nand U43434 (N_43434,N_37530,N_39053);
and U43435 (N_43435,N_38206,N_36707);
or U43436 (N_43436,N_37312,N_39877);
or U43437 (N_43437,N_37158,N_37119);
xor U43438 (N_43438,N_39669,N_38312);
nor U43439 (N_43439,N_35529,N_39488);
or U43440 (N_43440,N_35127,N_39723);
xnor U43441 (N_43441,N_35774,N_39279);
xor U43442 (N_43442,N_39752,N_38064);
xor U43443 (N_43443,N_39032,N_39330);
nand U43444 (N_43444,N_35539,N_38227);
nand U43445 (N_43445,N_36321,N_35437);
or U43446 (N_43446,N_37021,N_37006);
or U43447 (N_43447,N_37829,N_35502);
nand U43448 (N_43448,N_36238,N_37967);
nand U43449 (N_43449,N_36010,N_39340);
nor U43450 (N_43450,N_38243,N_39766);
or U43451 (N_43451,N_37833,N_38439);
or U43452 (N_43452,N_35729,N_35107);
nand U43453 (N_43453,N_36611,N_38228);
nor U43454 (N_43454,N_39008,N_39780);
nand U43455 (N_43455,N_35294,N_39662);
nand U43456 (N_43456,N_38413,N_38150);
nand U43457 (N_43457,N_39803,N_35910);
nor U43458 (N_43458,N_38093,N_35973);
or U43459 (N_43459,N_39529,N_38636);
xor U43460 (N_43460,N_37746,N_35116);
nor U43461 (N_43461,N_35870,N_39670);
and U43462 (N_43462,N_39789,N_38050);
and U43463 (N_43463,N_35112,N_38474);
nand U43464 (N_43464,N_38570,N_38170);
or U43465 (N_43465,N_39998,N_39841);
nor U43466 (N_43466,N_38627,N_37843);
xnor U43467 (N_43467,N_38114,N_36201);
nor U43468 (N_43468,N_35944,N_35957);
or U43469 (N_43469,N_35977,N_38878);
nor U43470 (N_43470,N_35896,N_37019);
nand U43471 (N_43471,N_38606,N_39290);
nor U43472 (N_43472,N_38378,N_35424);
and U43473 (N_43473,N_39577,N_36121);
xnor U43474 (N_43474,N_39254,N_38630);
and U43475 (N_43475,N_39247,N_38659);
and U43476 (N_43476,N_35691,N_37892);
or U43477 (N_43477,N_38844,N_37453);
nor U43478 (N_43478,N_38556,N_35501);
or U43479 (N_43479,N_37764,N_35709);
nand U43480 (N_43480,N_35406,N_38610);
nor U43481 (N_43481,N_37275,N_37251);
nand U43482 (N_43482,N_36052,N_37547);
xnor U43483 (N_43483,N_39736,N_36750);
or U43484 (N_43484,N_39688,N_39733);
and U43485 (N_43485,N_39713,N_38692);
or U43486 (N_43486,N_37618,N_39324);
and U43487 (N_43487,N_39183,N_36924);
or U43488 (N_43488,N_36189,N_36880);
nand U43489 (N_43489,N_38444,N_35664);
and U43490 (N_43490,N_36725,N_38800);
nor U43491 (N_43491,N_39817,N_39693);
xnor U43492 (N_43492,N_35437,N_37577);
or U43493 (N_43493,N_37618,N_35689);
nand U43494 (N_43494,N_35212,N_39918);
xnor U43495 (N_43495,N_36156,N_39539);
nor U43496 (N_43496,N_37678,N_36258);
and U43497 (N_43497,N_36111,N_38870);
nor U43498 (N_43498,N_36841,N_38244);
nand U43499 (N_43499,N_38195,N_37472);
nand U43500 (N_43500,N_38191,N_37052);
nand U43501 (N_43501,N_39162,N_37311);
xnor U43502 (N_43502,N_35216,N_39544);
xor U43503 (N_43503,N_38872,N_37245);
and U43504 (N_43504,N_37156,N_37516);
or U43505 (N_43505,N_39537,N_35945);
and U43506 (N_43506,N_36523,N_36530);
and U43507 (N_43507,N_38222,N_37482);
nor U43508 (N_43508,N_35079,N_39412);
nor U43509 (N_43509,N_36128,N_35039);
nor U43510 (N_43510,N_36642,N_38387);
nor U43511 (N_43511,N_35884,N_39110);
nand U43512 (N_43512,N_36716,N_36400);
nor U43513 (N_43513,N_39219,N_36856);
xor U43514 (N_43514,N_36069,N_35965);
and U43515 (N_43515,N_39285,N_39168);
nand U43516 (N_43516,N_38954,N_35365);
nor U43517 (N_43517,N_37659,N_39970);
or U43518 (N_43518,N_36538,N_38776);
nor U43519 (N_43519,N_39780,N_35140);
xor U43520 (N_43520,N_36071,N_38774);
or U43521 (N_43521,N_39726,N_38874);
nor U43522 (N_43522,N_39584,N_38784);
and U43523 (N_43523,N_38477,N_36233);
and U43524 (N_43524,N_35644,N_36950);
xor U43525 (N_43525,N_39403,N_39923);
nand U43526 (N_43526,N_35797,N_35677);
or U43527 (N_43527,N_38845,N_36659);
nand U43528 (N_43528,N_36390,N_39713);
nor U43529 (N_43529,N_37971,N_38759);
nand U43530 (N_43530,N_38679,N_37070);
or U43531 (N_43531,N_39784,N_37231);
nor U43532 (N_43532,N_39363,N_39732);
nor U43533 (N_43533,N_39781,N_39243);
and U43534 (N_43534,N_36613,N_36809);
and U43535 (N_43535,N_38088,N_39136);
and U43536 (N_43536,N_39579,N_39797);
and U43537 (N_43537,N_37001,N_35838);
nand U43538 (N_43538,N_38031,N_37030);
nand U43539 (N_43539,N_37469,N_39619);
xor U43540 (N_43540,N_35761,N_36900);
or U43541 (N_43541,N_38966,N_39016);
nor U43542 (N_43542,N_38983,N_37339);
nor U43543 (N_43543,N_38262,N_36019);
and U43544 (N_43544,N_38268,N_35138);
and U43545 (N_43545,N_35979,N_36010);
nand U43546 (N_43546,N_38507,N_39960);
and U43547 (N_43547,N_37494,N_39100);
or U43548 (N_43548,N_39508,N_38500);
nand U43549 (N_43549,N_37309,N_37051);
and U43550 (N_43550,N_38618,N_36118);
and U43551 (N_43551,N_35332,N_35952);
nor U43552 (N_43552,N_37251,N_37588);
and U43553 (N_43553,N_38489,N_35134);
nor U43554 (N_43554,N_36428,N_39376);
xnor U43555 (N_43555,N_36746,N_38117);
xor U43556 (N_43556,N_36089,N_38807);
nand U43557 (N_43557,N_37533,N_35934);
or U43558 (N_43558,N_37677,N_39192);
xor U43559 (N_43559,N_37386,N_37333);
nor U43560 (N_43560,N_38819,N_37644);
or U43561 (N_43561,N_39122,N_35662);
xnor U43562 (N_43562,N_36686,N_38779);
nor U43563 (N_43563,N_38501,N_37995);
and U43564 (N_43564,N_38721,N_37272);
nand U43565 (N_43565,N_35771,N_35643);
or U43566 (N_43566,N_35429,N_38921);
nand U43567 (N_43567,N_36285,N_37283);
or U43568 (N_43568,N_39451,N_35990);
nand U43569 (N_43569,N_39594,N_38116);
or U43570 (N_43570,N_35409,N_39402);
and U43571 (N_43571,N_38173,N_38728);
nor U43572 (N_43572,N_36211,N_35891);
nor U43573 (N_43573,N_39336,N_39123);
or U43574 (N_43574,N_37628,N_39486);
nand U43575 (N_43575,N_35746,N_36023);
nand U43576 (N_43576,N_37593,N_35745);
nor U43577 (N_43577,N_35804,N_36803);
and U43578 (N_43578,N_36148,N_37192);
or U43579 (N_43579,N_37149,N_36560);
and U43580 (N_43580,N_36982,N_38260);
nand U43581 (N_43581,N_36126,N_36551);
nand U43582 (N_43582,N_37339,N_35210);
nand U43583 (N_43583,N_38745,N_35986);
or U43584 (N_43584,N_38423,N_38812);
or U43585 (N_43585,N_39170,N_36377);
xor U43586 (N_43586,N_37386,N_36421);
or U43587 (N_43587,N_39720,N_37535);
and U43588 (N_43588,N_36942,N_36929);
nor U43589 (N_43589,N_36473,N_39838);
and U43590 (N_43590,N_39651,N_38399);
and U43591 (N_43591,N_39039,N_37993);
nand U43592 (N_43592,N_38461,N_38326);
or U43593 (N_43593,N_39547,N_35475);
nor U43594 (N_43594,N_36843,N_37182);
or U43595 (N_43595,N_39018,N_35217);
or U43596 (N_43596,N_35964,N_38499);
nand U43597 (N_43597,N_35067,N_35794);
nand U43598 (N_43598,N_36811,N_39513);
and U43599 (N_43599,N_35803,N_39255);
or U43600 (N_43600,N_39294,N_35378);
nand U43601 (N_43601,N_39252,N_35535);
nor U43602 (N_43602,N_35021,N_35037);
or U43603 (N_43603,N_35176,N_36826);
xnor U43604 (N_43604,N_39462,N_36461);
nor U43605 (N_43605,N_38955,N_36561);
and U43606 (N_43606,N_36895,N_37297);
or U43607 (N_43607,N_36517,N_35339);
or U43608 (N_43608,N_38481,N_39803);
or U43609 (N_43609,N_39149,N_38773);
or U43610 (N_43610,N_38194,N_36886);
and U43611 (N_43611,N_39143,N_36029);
nor U43612 (N_43612,N_35071,N_36859);
and U43613 (N_43613,N_39171,N_39163);
nand U43614 (N_43614,N_38568,N_35668);
nor U43615 (N_43615,N_35119,N_37027);
and U43616 (N_43616,N_39496,N_37274);
or U43617 (N_43617,N_36859,N_37832);
nand U43618 (N_43618,N_38201,N_36991);
or U43619 (N_43619,N_35375,N_35571);
and U43620 (N_43620,N_39785,N_36691);
xnor U43621 (N_43621,N_38506,N_37159);
or U43622 (N_43622,N_39392,N_35565);
xor U43623 (N_43623,N_37605,N_35975);
nor U43624 (N_43624,N_37960,N_35274);
nand U43625 (N_43625,N_35811,N_37408);
or U43626 (N_43626,N_39948,N_38779);
nand U43627 (N_43627,N_37520,N_35910);
and U43628 (N_43628,N_39504,N_36378);
or U43629 (N_43629,N_36562,N_38545);
and U43630 (N_43630,N_39197,N_37912);
and U43631 (N_43631,N_39392,N_38926);
nor U43632 (N_43632,N_36323,N_36928);
nand U43633 (N_43633,N_39025,N_37309);
nor U43634 (N_43634,N_38296,N_37090);
and U43635 (N_43635,N_37027,N_37557);
or U43636 (N_43636,N_36639,N_39713);
xor U43637 (N_43637,N_39562,N_38806);
nand U43638 (N_43638,N_38122,N_35318);
xnor U43639 (N_43639,N_38961,N_37650);
nand U43640 (N_43640,N_35401,N_39734);
xor U43641 (N_43641,N_36267,N_37985);
xnor U43642 (N_43642,N_39302,N_35968);
or U43643 (N_43643,N_39674,N_37627);
nand U43644 (N_43644,N_37353,N_39221);
and U43645 (N_43645,N_36469,N_37918);
or U43646 (N_43646,N_36602,N_37987);
and U43647 (N_43647,N_39131,N_39482);
or U43648 (N_43648,N_36805,N_35643);
xnor U43649 (N_43649,N_38426,N_35515);
nor U43650 (N_43650,N_39523,N_38637);
or U43651 (N_43651,N_39570,N_35358);
and U43652 (N_43652,N_39932,N_38784);
and U43653 (N_43653,N_35765,N_37319);
or U43654 (N_43654,N_35675,N_38618);
or U43655 (N_43655,N_35820,N_37141);
and U43656 (N_43656,N_35088,N_35552);
and U43657 (N_43657,N_36534,N_36695);
nand U43658 (N_43658,N_35712,N_37453);
nand U43659 (N_43659,N_37238,N_36229);
nor U43660 (N_43660,N_37321,N_35604);
nor U43661 (N_43661,N_36465,N_38172);
or U43662 (N_43662,N_35076,N_39630);
or U43663 (N_43663,N_36618,N_38667);
or U43664 (N_43664,N_37434,N_37649);
nor U43665 (N_43665,N_39966,N_38192);
and U43666 (N_43666,N_35012,N_37694);
or U43667 (N_43667,N_39443,N_36133);
xor U43668 (N_43668,N_37161,N_39641);
nand U43669 (N_43669,N_35264,N_37382);
nand U43670 (N_43670,N_36988,N_36313);
nor U43671 (N_43671,N_35016,N_35419);
nor U43672 (N_43672,N_37145,N_36480);
and U43673 (N_43673,N_37296,N_37958);
or U43674 (N_43674,N_36401,N_37725);
and U43675 (N_43675,N_39611,N_35204);
or U43676 (N_43676,N_35395,N_37099);
nand U43677 (N_43677,N_36606,N_36918);
nor U43678 (N_43678,N_37460,N_36189);
xnor U43679 (N_43679,N_39623,N_36542);
nand U43680 (N_43680,N_37674,N_36531);
nor U43681 (N_43681,N_35874,N_37580);
nand U43682 (N_43682,N_37233,N_36794);
and U43683 (N_43683,N_36880,N_36021);
or U43684 (N_43684,N_37343,N_36847);
or U43685 (N_43685,N_35332,N_39897);
nand U43686 (N_43686,N_36794,N_39997);
nor U43687 (N_43687,N_35914,N_35176);
or U43688 (N_43688,N_38946,N_38462);
nor U43689 (N_43689,N_37337,N_36557);
nand U43690 (N_43690,N_39622,N_39699);
nand U43691 (N_43691,N_35721,N_36346);
or U43692 (N_43692,N_36081,N_36059);
nor U43693 (N_43693,N_36167,N_38709);
nand U43694 (N_43694,N_39511,N_38089);
or U43695 (N_43695,N_36235,N_36479);
or U43696 (N_43696,N_37140,N_35226);
and U43697 (N_43697,N_36367,N_37399);
nor U43698 (N_43698,N_37949,N_39427);
nor U43699 (N_43699,N_37276,N_35041);
nor U43700 (N_43700,N_37510,N_35933);
nor U43701 (N_43701,N_39789,N_36167);
and U43702 (N_43702,N_35959,N_37944);
nand U43703 (N_43703,N_38878,N_39547);
and U43704 (N_43704,N_39955,N_37813);
or U43705 (N_43705,N_38874,N_37418);
nand U43706 (N_43706,N_35546,N_35363);
or U43707 (N_43707,N_35603,N_36942);
or U43708 (N_43708,N_37313,N_38960);
or U43709 (N_43709,N_35199,N_35729);
or U43710 (N_43710,N_38006,N_38614);
nand U43711 (N_43711,N_35199,N_36494);
nand U43712 (N_43712,N_37119,N_35575);
or U43713 (N_43713,N_39009,N_38440);
nand U43714 (N_43714,N_35850,N_37739);
and U43715 (N_43715,N_35354,N_37378);
and U43716 (N_43716,N_39951,N_35231);
and U43717 (N_43717,N_36353,N_36614);
nor U43718 (N_43718,N_38449,N_37195);
nand U43719 (N_43719,N_39362,N_38330);
and U43720 (N_43720,N_35211,N_39404);
nor U43721 (N_43721,N_37639,N_36101);
and U43722 (N_43722,N_38628,N_38213);
and U43723 (N_43723,N_36583,N_38593);
and U43724 (N_43724,N_37038,N_36442);
and U43725 (N_43725,N_37516,N_37309);
and U43726 (N_43726,N_36639,N_35766);
or U43727 (N_43727,N_36319,N_35506);
xnor U43728 (N_43728,N_37818,N_39571);
or U43729 (N_43729,N_35604,N_39395);
and U43730 (N_43730,N_38072,N_37750);
nor U43731 (N_43731,N_36633,N_37075);
nor U43732 (N_43732,N_36658,N_37773);
and U43733 (N_43733,N_35929,N_37426);
xnor U43734 (N_43734,N_35841,N_36397);
xor U43735 (N_43735,N_36637,N_39026);
nor U43736 (N_43736,N_39930,N_35868);
and U43737 (N_43737,N_38213,N_36616);
xnor U43738 (N_43738,N_39267,N_37533);
or U43739 (N_43739,N_36049,N_38452);
nand U43740 (N_43740,N_36906,N_36464);
or U43741 (N_43741,N_35171,N_38914);
nor U43742 (N_43742,N_37497,N_38009);
and U43743 (N_43743,N_36187,N_35917);
nand U43744 (N_43744,N_35955,N_35552);
or U43745 (N_43745,N_35839,N_38025);
or U43746 (N_43746,N_38423,N_38411);
nor U43747 (N_43747,N_37763,N_38942);
nand U43748 (N_43748,N_37615,N_35365);
nor U43749 (N_43749,N_36250,N_36543);
or U43750 (N_43750,N_37959,N_37357);
nand U43751 (N_43751,N_35995,N_37844);
nand U43752 (N_43752,N_35467,N_35486);
or U43753 (N_43753,N_39617,N_37541);
nand U43754 (N_43754,N_35962,N_39451);
nand U43755 (N_43755,N_38011,N_35356);
nand U43756 (N_43756,N_36109,N_39667);
and U43757 (N_43757,N_39618,N_35784);
or U43758 (N_43758,N_39695,N_37398);
or U43759 (N_43759,N_39531,N_39826);
nor U43760 (N_43760,N_39642,N_38064);
nand U43761 (N_43761,N_38195,N_35512);
nand U43762 (N_43762,N_37585,N_37641);
nor U43763 (N_43763,N_38659,N_35368);
or U43764 (N_43764,N_37047,N_39269);
nor U43765 (N_43765,N_38011,N_36015);
and U43766 (N_43766,N_36051,N_38204);
xnor U43767 (N_43767,N_38886,N_38317);
or U43768 (N_43768,N_39126,N_38346);
and U43769 (N_43769,N_37249,N_36570);
nor U43770 (N_43770,N_36874,N_38519);
nor U43771 (N_43771,N_35712,N_37478);
or U43772 (N_43772,N_38166,N_39739);
nor U43773 (N_43773,N_35344,N_35473);
nand U43774 (N_43774,N_38109,N_39803);
and U43775 (N_43775,N_36905,N_38611);
nor U43776 (N_43776,N_39231,N_39345);
xnor U43777 (N_43777,N_39931,N_38299);
or U43778 (N_43778,N_35352,N_37581);
xor U43779 (N_43779,N_37847,N_36673);
nor U43780 (N_43780,N_37021,N_35860);
nand U43781 (N_43781,N_36523,N_35437);
nand U43782 (N_43782,N_35388,N_36153);
or U43783 (N_43783,N_38452,N_39204);
or U43784 (N_43784,N_36079,N_39402);
and U43785 (N_43785,N_39822,N_35798);
or U43786 (N_43786,N_38843,N_38488);
or U43787 (N_43787,N_36764,N_37766);
and U43788 (N_43788,N_37795,N_35793);
xor U43789 (N_43789,N_38364,N_38043);
and U43790 (N_43790,N_37317,N_36995);
nor U43791 (N_43791,N_38952,N_36339);
nor U43792 (N_43792,N_37227,N_37892);
and U43793 (N_43793,N_35613,N_38123);
nor U43794 (N_43794,N_37668,N_38467);
and U43795 (N_43795,N_37710,N_39347);
or U43796 (N_43796,N_36776,N_39454);
xnor U43797 (N_43797,N_36621,N_38670);
or U43798 (N_43798,N_38549,N_38151);
nor U43799 (N_43799,N_37936,N_36587);
nand U43800 (N_43800,N_38006,N_35110);
nand U43801 (N_43801,N_37025,N_35086);
nand U43802 (N_43802,N_38954,N_39404);
nor U43803 (N_43803,N_36926,N_38614);
and U43804 (N_43804,N_39585,N_39748);
and U43805 (N_43805,N_38285,N_36152);
or U43806 (N_43806,N_38958,N_35243);
nor U43807 (N_43807,N_36890,N_38667);
nand U43808 (N_43808,N_35075,N_36301);
or U43809 (N_43809,N_35200,N_39734);
and U43810 (N_43810,N_35857,N_35830);
and U43811 (N_43811,N_35919,N_35996);
nor U43812 (N_43812,N_37327,N_38832);
nor U43813 (N_43813,N_38548,N_38024);
and U43814 (N_43814,N_36945,N_36952);
nand U43815 (N_43815,N_35916,N_36654);
or U43816 (N_43816,N_36710,N_38396);
nand U43817 (N_43817,N_36177,N_39710);
nand U43818 (N_43818,N_35576,N_36207);
nand U43819 (N_43819,N_35716,N_37837);
nor U43820 (N_43820,N_37652,N_35337);
and U43821 (N_43821,N_37808,N_35456);
nand U43822 (N_43822,N_35180,N_39927);
nor U43823 (N_43823,N_39164,N_35608);
nor U43824 (N_43824,N_35843,N_39887);
nor U43825 (N_43825,N_37156,N_36820);
xnor U43826 (N_43826,N_37680,N_35865);
nand U43827 (N_43827,N_35470,N_36419);
nand U43828 (N_43828,N_38997,N_39909);
or U43829 (N_43829,N_38880,N_37769);
and U43830 (N_43830,N_38107,N_36676);
nand U43831 (N_43831,N_39766,N_37561);
or U43832 (N_43832,N_35538,N_36330);
nor U43833 (N_43833,N_36764,N_38496);
nor U43834 (N_43834,N_37119,N_39553);
or U43835 (N_43835,N_38317,N_37973);
nand U43836 (N_43836,N_36726,N_36175);
and U43837 (N_43837,N_37743,N_35291);
nand U43838 (N_43838,N_37580,N_35069);
nand U43839 (N_43839,N_39548,N_38679);
nor U43840 (N_43840,N_35455,N_35739);
xor U43841 (N_43841,N_39568,N_37153);
and U43842 (N_43842,N_36993,N_35006);
xor U43843 (N_43843,N_39466,N_39487);
or U43844 (N_43844,N_37851,N_39588);
xnor U43845 (N_43845,N_38953,N_38545);
nand U43846 (N_43846,N_39537,N_35664);
nand U43847 (N_43847,N_36491,N_39801);
or U43848 (N_43848,N_35172,N_35036);
or U43849 (N_43849,N_36244,N_36213);
nor U43850 (N_43850,N_36873,N_36569);
and U43851 (N_43851,N_35163,N_37017);
or U43852 (N_43852,N_39070,N_35847);
nor U43853 (N_43853,N_37016,N_36567);
or U43854 (N_43854,N_37015,N_37042);
or U43855 (N_43855,N_35668,N_36918);
nor U43856 (N_43856,N_36709,N_39598);
nor U43857 (N_43857,N_37401,N_38902);
nor U43858 (N_43858,N_37261,N_38210);
and U43859 (N_43859,N_35569,N_39036);
xnor U43860 (N_43860,N_39870,N_35283);
nand U43861 (N_43861,N_38394,N_39241);
nand U43862 (N_43862,N_38391,N_37692);
nand U43863 (N_43863,N_36258,N_37796);
nand U43864 (N_43864,N_35699,N_36845);
and U43865 (N_43865,N_36742,N_37996);
and U43866 (N_43866,N_36651,N_38495);
nor U43867 (N_43867,N_38452,N_37178);
nor U43868 (N_43868,N_36860,N_39810);
nand U43869 (N_43869,N_36582,N_38375);
xor U43870 (N_43870,N_37484,N_38992);
nand U43871 (N_43871,N_38929,N_36556);
nand U43872 (N_43872,N_35961,N_39004);
nor U43873 (N_43873,N_37443,N_35344);
or U43874 (N_43874,N_36069,N_39192);
nand U43875 (N_43875,N_37017,N_37777);
nand U43876 (N_43876,N_35649,N_38291);
and U43877 (N_43877,N_35259,N_35890);
or U43878 (N_43878,N_39075,N_39406);
xnor U43879 (N_43879,N_38038,N_39720);
nor U43880 (N_43880,N_39197,N_39246);
nand U43881 (N_43881,N_39349,N_36766);
nor U43882 (N_43882,N_39079,N_38970);
nand U43883 (N_43883,N_37703,N_36492);
or U43884 (N_43884,N_38216,N_39256);
and U43885 (N_43885,N_38030,N_39068);
or U43886 (N_43886,N_35251,N_38232);
or U43887 (N_43887,N_36925,N_35394);
and U43888 (N_43888,N_35222,N_35616);
nor U43889 (N_43889,N_35680,N_37433);
nor U43890 (N_43890,N_37325,N_35035);
and U43891 (N_43891,N_35983,N_39530);
nand U43892 (N_43892,N_39025,N_39038);
and U43893 (N_43893,N_38224,N_35891);
or U43894 (N_43894,N_36902,N_37430);
and U43895 (N_43895,N_36388,N_38764);
nand U43896 (N_43896,N_39521,N_37195);
nand U43897 (N_43897,N_35787,N_38904);
nand U43898 (N_43898,N_38304,N_38741);
nor U43899 (N_43899,N_35164,N_39115);
and U43900 (N_43900,N_38290,N_39657);
nor U43901 (N_43901,N_38904,N_35493);
nor U43902 (N_43902,N_39980,N_37689);
nor U43903 (N_43903,N_36110,N_38293);
nand U43904 (N_43904,N_38541,N_39730);
or U43905 (N_43905,N_37651,N_36825);
nand U43906 (N_43906,N_39104,N_38137);
nor U43907 (N_43907,N_39355,N_35040);
nand U43908 (N_43908,N_35709,N_35944);
and U43909 (N_43909,N_39164,N_36356);
nor U43910 (N_43910,N_38620,N_37981);
nor U43911 (N_43911,N_39166,N_39742);
xnor U43912 (N_43912,N_35232,N_36206);
nand U43913 (N_43913,N_35170,N_38064);
nand U43914 (N_43914,N_38552,N_39803);
nor U43915 (N_43915,N_36953,N_39156);
and U43916 (N_43916,N_39375,N_38305);
nand U43917 (N_43917,N_37504,N_36148);
nand U43918 (N_43918,N_37081,N_39375);
xor U43919 (N_43919,N_35138,N_38044);
and U43920 (N_43920,N_39348,N_38327);
nand U43921 (N_43921,N_38200,N_36080);
nor U43922 (N_43922,N_37801,N_35890);
nand U43923 (N_43923,N_36051,N_35544);
nand U43924 (N_43924,N_36349,N_35821);
and U43925 (N_43925,N_35760,N_38700);
xor U43926 (N_43926,N_38390,N_39428);
nand U43927 (N_43927,N_35451,N_37385);
nand U43928 (N_43928,N_39244,N_36926);
xnor U43929 (N_43929,N_39420,N_38108);
nand U43930 (N_43930,N_39687,N_35960);
nor U43931 (N_43931,N_35788,N_36830);
nor U43932 (N_43932,N_37091,N_35228);
xor U43933 (N_43933,N_35864,N_35500);
or U43934 (N_43934,N_38038,N_36066);
nand U43935 (N_43935,N_35403,N_37157);
and U43936 (N_43936,N_36819,N_38670);
and U43937 (N_43937,N_35053,N_38317);
and U43938 (N_43938,N_39281,N_38693);
nor U43939 (N_43939,N_39353,N_37531);
xor U43940 (N_43940,N_38039,N_37382);
nand U43941 (N_43941,N_36370,N_37483);
or U43942 (N_43942,N_39788,N_35375);
nor U43943 (N_43943,N_39627,N_38169);
nor U43944 (N_43944,N_35111,N_38050);
and U43945 (N_43945,N_39472,N_36838);
and U43946 (N_43946,N_36382,N_35946);
and U43947 (N_43947,N_35322,N_38880);
xor U43948 (N_43948,N_38915,N_36135);
or U43949 (N_43949,N_36759,N_37793);
nor U43950 (N_43950,N_38288,N_39003);
nor U43951 (N_43951,N_38089,N_39612);
nor U43952 (N_43952,N_38046,N_37820);
and U43953 (N_43953,N_36100,N_35980);
or U43954 (N_43954,N_37292,N_37595);
and U43955 (N_43955,N_35411,N_37480);
nand U43956 (N_43956,N_38278,N_38459);
nand U43957 (N_43957,N_36247,N_39433);
nand U43958 (N_43958,N_38376,N_38507);
and U43959 (N_43959,N_35532,N_38061);
nor U43960 (N_43960,N_35739,N_38837);
and U43961 (N_43961,N_35899,N_37539);
nand U43962 (N_43962,N_37272,N_39737);
or U43963 (N_43963,N_39663,N_37271);
and U43964 (N_43964,N_35322,N_35660);
and U43965 (N_43965,N_35184,N_38827);
and U43966 (N_43966,N_38043,N_38594);
xor U43967 (N_43967,N_35710,N_37380);
nor U43968 (N_43968,N_35206,N_35222);
nor U43969 (N_43969,N_36426,N_39098);
nand U43970 (N_43970,N_39944,N_35474);
nand U43971 (N_43971,N_37935,N_37501);
nor U43972 (N_43972,N_37452,N_36739);
nand U43973 (N_43973,N_36729,N_39450);
and U43974 (N_43974,N_36445,N_36947);
and U43975 (N_43975,N_38880,N_35395);
nand U43976 (N_43976,N_35822,N_35145);
xnor U43977 (N_43977,N_37711,N_38205);
xnor U43978 (N_43978,N_35979,N_37902);
or U43979 (N_43979,N_36091,N_37686);
nor U43980 (N_43980,N_38411,N_35643);
and U43981 (N_43981,N_38957,N_37504);
xor U43982 (N_43982,N_38092,N_37682);
and U43983 (N_43983,N_37460,N_38481);
nand U43984 (N_43984,N_38520,N_36021);
nor U43985 (N_43985,N_39082,N_39284);
nor U43986 (N_43986,N_38241,N_39408);
xor U43987 (N_43987,N_36119,N_38684);
and U43988 (N_43988,N_37252,N_35716);
and U43989 (N_43989,N_38723,N_35204);
or U43990 (N_43990,N_35299,N_38204);
or U43991 (N_43991,N_39520,N_38734);
and U43992 (N_43992,N_39751,N_35397);
and U43993 (N_43993,N_39015,N_39675);
and U43994 (N_43994,N_36782,N_35596);
nor U43995 (N_43995,N_35714,N_38506);
nor U43996 (N_43996,N_36624,N_36848);
xnor U43997 (N_43997,N_37192,N_35738);
xnor U43998 (N_43998,N_39369,N_36005);
nand U43999 (N_43999,N_39197,N_37094);
xor U44000 (N_44000,N_36319,N_39313);
nand U44001 (N_44001,N_37931,N_38221);
nand U44002 (N_44002,N_38312,N_39896);
nor U44003 (N_44003,N_35408,N_37791);
xor U44004 (N_44004,N_36938,N_35252);
nand U44005 (N_44005,N_37469,N_35192);
and U44006 (N_44006,N_38176,N_39650);
or U44007 (N_44007,N_38283,N_38134);
nand U44008 (N_44008,N_37672,N_35491);
or U44009 (N_44009,N_36205,N_35185);
nand U44010 (N_44010,N_36361,N_35985);
and U44011 (N_44011,N_37806,N_38342);
nor U44012 (N_44012,N_39458,N_37579);
or U44013 (N_44013,N_37532,N_38202);
nand U44014 (N_44014,N_36790,N_38276);
or U44015 (N_44015,N_38163,N_36226);
nor U44016 (N_44016,N_39833,N_39554);
nand U44017 (N_44017,N_38949,N_36512);
and U44018 (N_44018,N_36216,N_37310);
and U44019 (N_44019,N_39988,N_38315);
xnor U44020 (N_44020,N_35515,N_35623);
xor U44021 (N_44021,N_36662,N_38215);
nand U44022 (N_44022,N_38053,N_35906);
or U44023 (N_44023,N_35917,N_38518);
or U44024 (N_44024,N_37129,N_39781);
and U44025 (N_44025,N_39244,N_39230);
xor U44026 (N_44026,N_37655,N_38673);
or U44027 (N_44027,N_38794,N_35501);
and U44028 (N_44028,N_35577,N_39576);
and U44029 (N_44029,N_38079,N_38480);
or U44030 (N_44030,N_36610,N_36659);
or U44031 (N_44031,N_37524,N_38804);
and U44032 (N_44032,N_38565,N_39968);
nor U44033 (N_44033,N_36141,N_37012);
or U44034 (N_44034,N_35761,N_38355);
nand U44035 (N_44035,N_37056,N_36049);
nor U44036 (N_44036,N_35354,N_35808);
nand U44037 (N_44037,N_38245,N_36671);
or U44038 (N_44038,N_35250,N_38799);
nor U44039 (N_44039,N_37394,N_39691);
or U44040 (N_44040,N_36577,N_35436);
nand U44041 (N_44041,N_39783,N_39542);
or U44042 (N_44042,N_35243,N_38237);
nand U44043 (N_44043,N_39826,N_38786);
or U44044 (N_44044,N_36731,N_38618);
nor U44045 (N_44045,N_35840,N_36443);
nand U44046 (N_44046,N_36580,N_37562);
or U44047 (N_44047,N_36457,N_36354);
xnor U44048 (N_44048,N_38336,N_35382);
nor U44049 (N_44049,N_36380,N_38642);
or U44050 (N_44050,N_38727,N_35319);
nand U44051 (N_44051,N_38284,N_38960);
and U44052 (N_44052,N_37691,N_37526);
nor U44053 (N_44053,N_39753,N_37355);
nor U44054 (N_44054,N_35398,N_37501);
and U44055 (N_44055,N_39526,N_38059);
nand U44056 (N_44056,N_35283,N_35279);
nor U44057 (N_44057,N_38978,N_35291);
nand U44058 (N_44058,N_39825,N_39504);
nor U44059 (N_44059,N_36332,N_36936);
nor U44060 (N_44060,N_36416,N_36665);
or U44061 (N_44061,N_36266,N_37292);
nand U44062 (N_44062,N_36754,N_36042);
nand U44063 (N_44063,N_39053,N_35211);
nand U44064 (N_44064,N_36435,N_36711);
nand U44065 (N_44065,N_35152,N_38219);
or U44066 (N_44066,N_38803,N_36769);
nor U44067 (N_44067,N_36620,N_39690);
and U44068 (N_44068,N_39255,N_37070);
and U44069 (N_44069,N_36484,N_39920);
and U44070 (N_44070,N_35096,N_35854);
or U44071 (N_44071,N_37773,N_38196);
nand U44072 (N_44072,N_35156,N_37111);
or U44073 (N_44073,N_35976,N_36186);
nand U44074 (N_44074,N_37058,N_35984);
or U44075 (N_44075,N_37407,N_38757);
nand U44076 (N_44076,N_38430,N_36167);
nand U44077 (N_44077,N_39755,N_37285);
nor U44078 (N_44078,N_38518,N_36634);
nor U44079 (N_44079,N_35248,N_37283);
nor U44080 (N_44080,N_36092,N_38045);
and U44081 (N_44081,N_39416,N_37942);
nand U44082 (N_44082,N_36570,N_37995);
and U44083 (N_44083,N_37305,N_37128);
nor U44084 (N_44084,N_37873,N_36658);
xnor U44085 (N_44085,N_36479,N_38106);
nand U44086 (N_44086,N_38173,N_35809);
and U44087 (N_44087,N_38340,N_36447);
and U44088 (N_44088,N_37991,N_37728);
or U44089 (N_44089,N_39717,N_37893);
nor U44090 (N_44090,N_36155,N_35090);
nand U44091 (N_44091,N_36656,N_39541);
nor U44092 (N_44092,N_38457,N_35568);
and U44093 (N_44093,N_39594,N_35893);
and U44094 (N_44094,N_35900,N_36812);
or U44095 (N_44095,N_35744,N_39683);
or U44096 (N_44096,N_39683,N_38758);
and U44097 (N_44097,N_35105,N_38296);
nor U44098 (N_44098,N_35061,N_38878);
xnor U44099 (N_44099,N_35837,N_39260);
nand U44100 (N_44100,N_35167,N_35586);
nor U44101 (N_44101,N_39661,N_38939);
and U44102 (N_44102,N_38796,N_35828);
and U44103 (N_44103,N_35689,N_38330);
nand U44104 (N_44104,N_39997,N_36852);
xnor U44105 (N_44105,N_35110,N_37772);
nor U44106 (N_44106,N_39000,N_39782);
and U44107 (N_44107,N_39571,N_36387);
nor U44108 (N_44108,N_35294,N_37953);
nor U44109 (N_44109,N_38086,N_39087);
nor U44110 (N_44110,N_38102,N_37503);
nand U44111 (N_44111,N_36766,N_38540);
and U44112 (N_44112,N_35013,N_36078);
or U44113 (N_44113,N_38559,N_38063);
nand U44114 (N_44114,N_36034,N_39493);
nand U44115 (N_44115,N_35206,N_35033);
nand U44116 (N_44116,N_36465,N_35775);
and U44117 (N_44117,N_38241,N_38669);
nand U44118 (N_44118,N_39135,N_38215);
and U44119 (N_44119,N_35371,N_35574);
and U44120 (N_44120,N_35949,N_36512);
xnor U44121 (N_44121,N_36965,N_39900);
and U44122 (N_44122,N_35895,N_38267);
xnor U44123 (N_44123,N_39229,N_37359);
nand U44124 (N_44124,N_39386,N_38192);
or U44125 (N_44125,N_39852,N_39725);
or U44126 (N_44126,N_35309,N_38463);
or U44127 (N_44127,N_38231,N_39542);
or U44128 (N_44128,N_38788,N_37673);
nand U44129 (N_44129,N_37133,N_38100);
and U44130 (N_44130,N_36841,N_36761);
or U44131 (N_44131,N_37058,N_37926);
or U44132 (N_44132,N_38857,N_39966);
or U44133 (N_44133,N_38160,N_37213);
xnor U44134 (N_44134,N_39099,N_39685);
nor U44135 (N_44135,N_38374,N_36145);
or U44136 (N_44136,N_38956,N_35566);
or U44137 (N_44137,N_35224,N_38474);
and U44138 (N_44138,N_36350,N_38278);
nand U44139 (N_44139,N_39887,N_36099);
nand U44140 (N_44140,N_37010,N_38254);
nand U44141 (N_44141,N_37538,N_35875);
or U44142 (N_44142,N_36857,N_35253);
or U44143 (N_44143,N_36891,N_39566);
nand U44144 (N_44144,N_35052,N_36206);
nand U44145 (N_44145,N_36682,N_38990);
nor U44146 (N_44146,N_39095,N_35238);
nor U44147 (N_44147,N_36699,N_38372);
nand U44148 (N_44148,N_39161,N_35808);
and U44149 (N_44149,N_38767,N_39468);
and U44150 (N_44150,N_39329,N_39222);
or U44151 (N_44151,N_35883,N_38271);
nand U44152 (N_44152,N_37623,N_35946);
or U44153 (N_44153,N_39752,N_38761);
nand U44154 (N_44154,N_37063,N_38067);
or U44155 (N_44155,N_36051,N_35088);
nand U44156 (N_44156,N_37619,N_35008);
and U44157 (N_44157,N_35715,N_38873);
nor U44158 (N_44158,N_37813,N_35692);
nor U44159 (N_44159,N_36725,N_38843);
nand U44160 (N_44160,N_36834,N_39343);
nand U44161 (N_44161,N_36306,N_36275);
nor U44162 (N_44162,N_38840,N_39023);
nor U44163 (N_44163,N_36220,N_37470);
or U44164 (N_44164,N_37992,N_36515);
and U44165 (N_44165,N_35216,N_35671);
or U44166 (N_44166,N_36997,N_38234);
nor U44167 (N_44167,N_37948,N_38898);
and U44168 (N_44168,N_39086,N_35346);
nand U44169 (N_44169,N_39691,N_37576);
nand U44170 (N_44170,N_36101,N_36631);
nor U44171 (N_44171,N_38958,N_38437);
or U44172 (N_44172,N_35869,N_38356);
nor U44173 (N_44173,N_36121,N_37138);
and U44174 (N_44174,N_35524,N_35273);
and U44175 (N_44175,N_39354,N_35145);
nor U44176 (N_44176,N_38020,N_35330);
nand U44177 (N_44177,N_37852,N_36279);
nor U44178 (N_44178,N_36816,N_39375);
nand U44179 (N_44179,N_38337,N_36300);
or U44180 (N_44180,N_37415,N_35578);
xor U44181 (N_44181,N_37161,N_38620);
and U44182 (N_44182,N_35862,N_38565);
nand U44183 (N_44183,N_37154,N_36994);
or U44184 (N_44184,N_35227,N_38859);
or U44185 (N_44185,N_35389,N_38736);
nor U44186 (N_44186,N_37193,N_36706);
nor U44187 (N_44187,N_39080,N_35739);
nand U44188 (N_44188,N_39381,N_37618);
nand U44189 (N_44189,N_37749,N_36809);
and U44190 (N_44190,N_36662,N_37147);
nand U44191 (N_44191,N_36283,N_39561);
and U44192 (N_44192,N_39825,N_37325);
and U44193 (N_44193,N_37470,N_39020);
xor U44194 (N_44194,N_36585,N_35179);
and U44195 (N_44195,N_39168,N_39816);
nand U44196 (N_44196,N_38082,N_37413);
nor U44197 (N_44197,N_35187,N_38418);
and U44198 (N_44198,N_35608,N_35868);
nor U44199 (N_44199,N_39871,N_36619);
and U44200 (N_44200,N_35134,N_37874);
or U44201 (N_44201,N_37415,N_36882);
nand U44202 (N_44202,N_39918,N_38423);
nor U44203 (N_44203,N_39740,N_35095);
nor U44204 (N_44204,N_36279,N_39462);
or U44205 (N_44205,N_37349,N_37628);
nor U44206 (N_44206,N_38859,N_37050);
nor U44207 (N_44207,N_36449,N_36736);
and U44208 (N_44208,N_36466,N_38443);
or U44209 (N_44209,N_37237,N_37682);
xor U44210 (N_44210,N_39533,N_39960);
nand U44211 (N_44211,N_39496,N_36585);
xor U44212 (N_44212,N_37203,N_35695);
or U44213 (N_44213,N_38369,N_38178);
or U44214 (N_44214,N_36339,N_36643);
and U44215 (N_44215,N_36927,N_37605);
or U44216 (N_44216,N_35260,N_37663);
nor U44217 (N_44217,N_38809,N_36684);
nor U44218 (N_44218,N_36292,N_37360);
nand U44219 (N_44219,N_39465,N_38166);
nor U44220 (N_44220,N_36408,N_36507);
nor U44221 (N_44221,N_36898,N_36376);
or U44222 (N_44222,N_37924,N_36405);
or U44223 (N_44223,N_35124,N_35955);
nand U44224 (N_44224,N_35328,N_39559);
and U44225 (N_44225,N_36149,N_35965);
xnor U44226 (N_44226,N_39282,N_36825);
nor U44227 (N_44227,N_38196,N_39517);
nand U44228 (N_44228,N_36406,N_39259);
nor U44229 (N_44229,N_39514,N_35086);
nor U44230 (N_44230,N_36783,N_38428);
or U44231 (N_44231,N_36905,N_38045);
and U44232 (N_44232,N_38196,N_39622);
nand U44233 (N_44233,N_38239,N_39931);
nor U44234 (N_44234,N_39886,N_35700);
nor U44235 (N_44235,N_39363,N_35733);
or U44236 (N_44236,N_38437,N_35437);
nand U44237 (N_44237,N_39295,N_36915);
nand U44238 (N_44238,N_38469,N_38934);
nand U44239 (N_44239,N_36379,N_35546);
nand U44240 (N_44240,N_35307,N_36871);
nand U44241 (N_44241,N_35904,N_35462);
or U44242 (N_44242,N_35065,N_37255);
or U44243 (N_44243,N_38933,N_38951);
nor U44244 (N_44244,N_39324,N_37364);
nand U44245 (N_44245,N_35800,N_37440);
and U44246 (N_44246,N_37458,N_36576);
or U44247 (N_44247,N_39648,N_36432);
or U44248 (N_44248,N_37425,N_39273);
xor U44249 (N_44249,N_37822,N_35403);
nor U44250 (N_44250,N_35026,N_35499);
nand U44251 (N_44251,N_39304,N_37465);
nor U44252 (N_44252,N_37203,N_39052);
and U44253 (N_44253,N_38570,N_36473);
and U44254 (N_44254,N_36500,N_35856);
and U44255 (N_44255,N_38025,N_35793);
or U44256 (N_44256,N_36852,N_37251);
nor U44257 (N_44257,N_35232,N_39159);
nor U44258 (N_44258,N_38823,N_39912);
nor U44259 (N_44259,N_38710,N_38847);
nand U44260 (N_44260,N_35089,N_36621);
xnor U44261 (N_44261,N_39388,N_38548);
and U44262 (N_44262,N_37383,N_37602);
nand U44263 (N_44263,N_38626,N_39145);
nor U44264 (N_44264,N_38679,N_37122);
nor U44265 (N_44265,N_38073,N_38012);
and U44266 (N_44266,N_39408,N_36696);
and U44267 (N_44267,N_38341,N_35880);
xor U44268 (N_44268,N_37370,N_37460);
or U44269 (N_44269,N_37087,N_35700);
or U44270 (N_44270,N_39949,N_38013);
or U44271 (N_44271,N_39138,N_39585);
nor U44272 (N_44272,N_37468,N_37196);
nand U44273 (N_44273,N_36992,N_35514);
and U44274 (N_44274,N_35962,N_38089);
or U44275 (N_44275,N_37723,N_38517);
or U44276 (N_44276,N_36596,N_37259);
xor U44277 (N_44277,N_35878,N_37794);
or U44278 (N_44278,N_38103,N_39070);
and U44279 (N_44279,N_36788,N_36781);
or U44280 (N_44280,N_35549,N_35626);
xnor U44281 (N_44281,N_39921,N_36478);
nand U44282 (N_44282,N_39975,N_37028);
or U44283 (N_44283,N_36212,N_38565);
nor U44284 (N_44284,N_39924,N_39744);
nor U44285 (N_44285,N_35424,N_36278);
and U44286 (N_44286,N_35171,N_35979);
nor U44287 (N_44287,N_38154,N_35946);
or U44288 (N_44288,N_37470,N_38075);
xor U44289 (N_44289,N_38702,N_35625);
nor U44290 (N_44290,N_38588,N_39493);
or U44291 (N_44291,N_35655,N_39043);
and U44292 (N_44292,N_38035,N_37215);
and U44293 (N_44293,N_38510,N_36926);
or U44294 (N_44294,N_35990,N_38605);
nand U44295 (N_44295,N_38165,N_38972);
and U44296 (N_44296,N_37081,N_37251);
and U44297 (N_44297,N_36584,N_37539);
and U44298 (N_44298,N_39788,N_38880);
nand U44299 (N_44299,N_35845,N_39508);
and U44300 (N_44300,N_35540,N_35664);
nand U44301 (N_44301,N_35195,N_35571);
nand U44302 (N_44302,N_36207,N_36823);
or U44303 (N_44303,N_38329,N_37422);
or U44304 (N_44304,N_36477,N_36826);
nand U44305 (N_44305,N_39759,N_39584);
nor U44306 (N_44306,N_37959,N_38121);
nand U44307 (N_44307,N_36395,N_36254);
or U44308 (N_44308,N_39019,N_38867);
and U44309 (N_44309,N_39724,N_36195);
nand U44310 (N_44310,N_36047,N_38443);
or U44311 (N_44311,N_38964,N_37793);
nand U44312 (N_44312,N_39826,N_36423);
nor U44313 (N_44313,N_35465,N_38832);
nor U44314 (N_44314,N_36617,N_35247);
nor U44315 (N_44315,N_37719,N_38170);
xnor U44316 (N_44316,N_39723,N_38678);
nand U44317 (N_44317,N_39127,N_36555);
nand U44318 (N_44318,N_36442,N_38266);
and U44319 (N_44319,N_37329,N_35079);
and U44320 (N_44320,N_36637,N_37688);
or U44321 (N_44321,N_39733,N_37957);
xnor U44322 (N_44322,N_37201,N_36109);
and U44323 (N_44323,N_37441,N_36460);
and U44324 (N_44324,N_36704,N_39548);
nor U44325 (N_44325,N_39661,N_38166);
and U44326 (N_44326,N_39015,N_37605);
and U44327 (N_44327,N_39161,N_38939);
nand U44328 (N_44328,N_35784,N_35896);
nor U44329 (N_44329,N_36638,N_38985);
nand U44330 (N_44330,N_35286,N_35265);
and U44331 (N_44331,N_39541,N_37771);
or U44332 (N_44332,N_39923,N_37835);
nand U44333 (N_44333,N_36728,N_39416);
or U44334 (N_44334,N_38005,N_35259);
nor U44335 (N_44335,N_39059,N_39630);
and U44336 (N_44336,N_39446,N_38463);
nand U44337 (N_44337,N_39092,N_37316);
nand U44338 (N_44338,N_36378,N_36944);
or U44339 (N_44339,N_36758,N_37007);
or U44340 (N_44340,N_39661,N_35066);
and U44341 (N_44341,N_35215,N_36768);
and U44342 (N_44342,N_38082,N_35831);
xnor U44343 (N_44343,N_38787,N_37894);
xor U44344 (N_44344,N_35817,N_35284);
xnor U44345 (N_44345,N_39945,N_35935);
nor U44346 (N_44346,N_39870,N_35082);
or U44347 (N_44347,N_36927,N_35897);
nor U44348 (N_44348,N_35292,N_39117);
and U44349 (N_44349,N_39560,N_38752);
and U44350 (N_44350,N_35487,N_37743);
or U44351 (N_44351,N_35087,N_38527);
or U44352 (N_44352,N_37345,N_38811);
and U44353 (N_44353,N_36757,N_35612);
or U44354 (N_44354,N_35758,N_35097);
and U44355 (N_44355,N_36684,N_36047);
xnor U44356 (N_44356,N_38204,N_35107);
nand U44357 (N_44357,N_37121,N_39243);
and U44358 (N_44358,N_38124,N_38652);
nand U44359 (N_44359,N_39173,N_35719);
or U44360 (N_44360,N_36305,N_35917);
xnor U44361 (N_44361,N_37180,N_35510);
or U44362 (N_44362,N_36281,N_37963);
nand U44363 (N_44363,N_36897,N_38000);
and U44364 (N_44364,N_38751,N_35810);
and U44365 (N_44365,N_35946,N_39082);
and U44366 (N_44366,N_39084,N_36886);
or U44367 (N_44367,N_38707,N_39357);
or U44368 (N_44368,N_36551,N_35702);
nand U44369 (N_44369,N_37662,N_36426);
nand U44370 (N_44370,N_36672,N_37182);
and U44371 (N_44371,N_35123,N_37900);
and U44372 (N_44372,N_39789,N_39495);
nand U44373 (N_44373,N_35849,N_38374);
nor U44374 (N_44374,N_37856,N_37705);
and U44375 (N_44375,N_38241,N_35129);
nand U44376 (N_44376,N_39989,N_35729);
and U44377 (N_44377,N_39620,N_39492);
and U44378 (N_44378,N_39732,N_36843);
nor U44379 (N_44379,N_39527,N_36491);
nor U44380 (N_44380,N_37315,N_38567);
and U44381 (N_44381,N_39888,N_38928);
or U44382 (N_44382,N_36703,N_37453);
and U44383 (N_44383,N_38969,N_37338);
xnor U44384 (N_44384,N_39210,N_39260);
or U44385 (N_44385,N_37121,N_35432);
nor U44386 (N_44386,N_39451,N_38340);
and U44387 (N_44387,N_37844,N_35422);
or U44388 (N_44388,N_39677,N_38036);
or U44389 (N_44389,N_36387,N_39527);
or U44390 (N_44390,N_36178,N_35630);
or U44391 (N_44391,N_38907,N_37682);
nor U44392 (N_44392,N_39690,N_39547);
xnor U44393 (N_44393,N_35504,N_39389);
nand U44394 (N_44394,N_37690,N_36344);
or U44395 (N_44395,N_36468,N_35291);
or U44396 (N_44396,N_39039,N_36350);
nand U44397 (N_44397,N_37847,N_37070);
nand U44398 (N_44398,N_35346,N_38806);
and U44399 (N_44399,N_39651,N_35428);
nor U44400 (N_44400,N_37259,N_37173);
or U44401 (N_44401,N_37700,N_35927);
and U44402 (N_44402,N_39754,N_37562);
nand U44403 (N_44403,N_36731,N_35905);
or U44404 (N_44404,N_36579,N_35561);
nor U44405 (N_44405,N_36784,N_38077);
and U44406 (N_44406,N_35035,N_39793);
nand U44407 (N_44407,N_39984,N_39373);
nor U44408 (N_44408,N_39682,N_38802);
and U44409 (N_44409,N_36349,N_38074);
nand U44410 (N_44410,N_38675,N_37474);
nand U44411 (N_44411,N_36700,N_36549);
nor U44412 (N_44412,N_39638,N_37597);
nor U44413 (N_44413,N_35069,N_35033);
or U44414 (N_44414,N_39400,N_36834);
or U44415 (N_44415,N_38894,N_35164);
and U44416 (N_44416,N_38831,N_39722);
or U44417 (N_44417,N_37545,N_35047);
and U44418 (N_44418,N_36609,N_35797);
and U44419 (N_44419,N_37824,N_36820);
nor U44420 (N_44420,N_36558,N_36143);
xnor U44421 (N_44421,N_37968,N_37757);
nor U44422 (N_44422,N_35205,N_39800);
nor U44423 (N_44423,N_36971,N_35928);
or U44424 (N_44424,N_36799,N_37287);
nor U44425 (N_44425,N_39794,N_35043);
and U44426 (N_44426,N_37937,N_36909);
and U44427 (N_44427,N_38590,N_37301);
nor U44428 (N_44428,N_37495,N_39292);
xor U44429 (N_44429,N_35793,N_39423);
nand U44430 (N_44430,N_39984,N_38112);
nand U44431 (N_44431,N_35956,N_39493);
xor U44432 (N_44432,N_37262,N_35041);
nand U44433 (N_44433,N_37597,N_36244);
and U44434 (N_44434,N_35805,N_37392);
nand U44435 (N_44435,N_35140,N_35058);
or U44436 (N_44436,N_37230,N_36697);
nand U44437 (N_44437,N_36203,N_38586);
nand U44438 (N_44438,N_36171,N_39492);
and U44439 (N_44439,N_36464,N_37706);
nand U44440 (N_44440,N_36590,N_37129);
or U44441 (N_44441,N_37825,N_36819);
nor U44442 (N_44442,N_39191,N_37095);
nor U44443 (N_44443,N_39189,N_38340);
nand U44444 (N_44444,N_36386,N_39451);
xor U44445 (N_44445,N_35767,N_35952);
and U44446 (N_44446,N_35692,N_39939);
and U44447 (N_44447,N_36690,N_35652);
nand U44448 (N_44448,N_38469,N_39554);
or U44449 (N_44449,N_37208,N_36412);
or U44450 (N_44450,N_36572,N_36879);
nand U44451 (N_44451,N_36903,N_35785);
xor U44452 (N_44452,N_36002,N_38751);
nor U44453 (N_44453,N_39111,N_38698);
xor U44454 (N_44454,N_37207,N_35742);
or U44455 (N_44455,N_36782,N_35379);
nand U44456 (N_44456,N_35717,N_39269);
nand U44457 (N_44457,N_35053,N_39211);
nor U44458 (N_44458,N_37144,N_35194);
and U44459 (N_44459,N_39834,N_38820);
and U44460 (N_44460,N_35725,N_37678);
nor U44461 (N_44461,N_39274,N_38567);
nor U44462 (N_44462,N_37392,N_36202);
and U44463 (N_44463,N_35298,N_37479);
nor U44464 (N_44464,N_36362,N_39950);
nor U44465 (N_44465,N_37045,N_38655);
or U44466 (N_44466,N_36939,N_35103);
or U44467 (N_44467,N_37438,N_35803);
nor U44468 (N_44468,N_35579,N_36356);
nor U44469 (N_44469,N_36627,N_37800);
nor U44470 (N_44470,N_38972,N_35991);
and U44471 (N_44471,N_39961,N_36706);
or U44472 (N_44472,N_35948,N_38935);
and U44473 (N_44473,N_39058,N_39292);
nor U44474 (N_44474,N_36657,N_37832);
and U44475 (N_44475,N_36949,N_35648);
or U44476 (N_44476,N_39888,N_35548);
nand U44477 (N_44477,N_39210,N_36278);
nor U44478 (N_44478,N_36829,N_38266);
nand U44479 (N_44479,N_39630,N_36774);
and U44480 (N_44480,N_35685,N_39149);
nor U44481 (N_44481,N_36109,N_36324);
nor U44482 (N_44482,N_35549,N_38457);
nor U44483 (N_44483,N_35263,N_36798);
or U44484 (N_44484,N_38597,N_35096);
nor U44485 (N_44485,N_39973,N_37199);
nand U44486 (N_44486,N_36028,N_38106);
or U44487 (N_44487,N_36993,N_38456);
nor U44488 (N_44488,N_39234,N_39408);
xnor U44489 (N_44489,N_37493,N_35097);
nor U44490 (N_44490,N_38705,N_35702);
or U44491 (N_44491,N_38830,N_39052);
nor U44492 (N_44492,N_35985,N_38615);
and U44493 (N_44493,N_37762,N_39710);
nor U44494 (N_44494,N_38430,N_39054);
or U44495 (N_44495,N_36130,N_36010);
and U44496 (N_44496,N_38370,N_37954);
and U44497 (N_44497,N_37365,N_38071);
xnor U44498 (N_44498,N_35862,N_36291);
or U44499 (N_44499,N_35082,N_35825);
nand U44500 (N_44500,N_36713,N_35282);
or U44501 (N_44501,N_35763,N_39517);
nor U44502 (N_44502,N_38826,N_36724);
and U44503 (N_44503,N_37560,N_37501);
or U44504 (N_44504,N_37761,N_37120);
and U44505 (N_44505,N_35450,N_37009);
and U44506 (N_44506,N_38843,N_35441);
and U44507 (N_44507,N_37200,N_39976);
xor U44508 (N_44508,N_36163,N_36906);
nor U44509 (N_44509,N_36372,N_39432);
and U44510 (N_44510,N_35453,N_37967);
nand U44511 (N_44511,N_35711,N_38465);
or U44512 (N_44512,N_36961,N_38482);
nor U44513 (N_44513,N_36835,N_36369);
nor U44514 (N_44514,N_35194,N_37224);
nand U44515 (N_44515,N_38978,N_39734);
and U44516 (N_44516,N_36942,N_39850);
or U44517 (N_44517,N_39562,N_35707);
or U44518 (N_44518,N_39367,N_38741);
xnor U44519 (N_44519,N_39744,N_35686);
xor U44520 (N_44520,N_35562,N_36032);
nor U44521 (N_44521,N_35937,N_39340);
nand U44522 (N_44522,N_37918,N_39731);
nor U44523 (N_44523,N_37344,N_38845);
and U44524 (N_44524,N_38145,N_36908);
nor U44525 (N_44525,N_39452,N_39765);
or U44526 (N_44526,N_35549,N_35187);
and U44527 (N_44527,N_36826,N_35150);
nand U44528 (N_44528,N_39917,N_36855);
or U44529 (N_44529,N_38153,N_39005);
or U44530 (N_44530,N_35009,N_39606);
and U44531 (N_44531,N_39451,N_39640);
nor U44532 (N_44532,N_38491,N_36841);
and U44533 (N_44533,N_36493,N_35627);
and U44534 (N_44534,N_39147,N_35181);
and U44535 (N_44535,N_38307,N_39137);
and U44536 (N_44536,N_39048,N_36110);
or U44537 (N_44537,N_37047,N_35214);
nor U44538 (N_44538,N_39551,N_36760);
or U44539 (N_44539,N_38007,N_35931);
nand U44540 (N_44540,N_35806,N_36791);
and U44541 (N_44541,N_36076,N_38147);
and U44542 (N_44542,N_39367,N_38644);
or U44543 (N_44543,N_35973,N_38884);
nor U44544 (N_44544,N_37052,N_35393);
nand U44545 (N_44545,N_39070,N_36705);
nor U44546 (N_44546,N_36542,N_38959);
xnor U44547 (N_44547,N_38246,N_35933);
or U44548 (N_44548,N_35753,N_39575);
nand U44549 (N_44549,N_36546,N_35963);
nor U44550 (N_44550,N_35466,N_38225);
nand U44551 (N_44551,N_37312,N_37271);
nor U44552 (N_44552,N_38138,N_39018);
nand U44553 (N_44553,N_39089,N_36810);
nor U44554 (N_44554,N_37482,N_38864);
or U44555 (N_44555,N_39871,N_35111);
and U44556 (N_44556,N_36549,N_36028);
xnor U44557 (N_44557,N_36294,N_39344);
nor U44558 (N_44558,N_39674,N_35128);
nand U44559 (N_44559,N_35612,N_36670);
and U44560 (N_44560,N_37100,N_35799);
nor U44561 (N_44561,N_37019,N_37218);
nand U44562 (N_44562,N_37702,N_38215);
and U44563 (N_44563,N_36787,N_36373);
xnor U44564 (N_44564,N_38256,N_39733);
nand U44565 (N_44565,N_37462,N_38909);
and U44566 (N_44566,N_36799,N_37845);
nand U44567 (N_44567,N_39092,N_35056);
nor U44568 (N_44568,N_38919,N_38879);
nor U44569 (N_44569,N_35405,N_38204);
nor U44570 (N_44570,N_39149,N_36508);
xnor U44571 (N_44571,N_37310,N_37133);
and U44572 (N_44572,N_39267,N_35707);
nand U44573 (N_44573,N_35892,N_36524);
and U44574 (N_44574,N_35126,N_35021);
and U44575 (N_44575,N_35787,N_37039);
nor U44576 (N_44576,N_38951,N_36962);
nor U44577 (N_44577,N_38956,N_38191);
nor U44578 (N_44578,N_35477,N_36868);
or U44579 (N_44579,N_35962,N_35229);
and U44580 (N_44580,N_37166,N_35808);
or U44581 (N_44581,N_39860,N_37125);
or U44582 (N_44582,N_36989,N_37378);
nor U44583 (N_44583,N_37362,N_39337);
xnor U44584 (N_44584,N_35166,N_38981);
or U44585 (N_44585,N_37472,N_38044);
xor U44586 (N_44586,N_37394,N_38382);
nand U44587 (N_44587,N_36490,N_35154);
nand U44588 (N_44588,N_37560,N_37943);
or U44589 (N_44589,N_36356,N_35150);
nor U44590 (N_44590,N_38360,N_38432);
nand U44591 (N_44591,N_39493,N_37056);
nor U44592 (N_44592,N_37632,N_36445);
or U44593 (N_44593,N_38438,N_35195);
nand U44594 (N_44594,N_37927,N_37906);
nand U44595 (N_44595,N_38044,N_39710);
nor U44596 (N_44596,N_36358,N_39475);
nand U44597 (N_44597,N_38167,N_38346);
or U44598 (N_44598,N_37641,N_36161);
nor U44599 (N_44599,N_35811,N_37225);
nor U44600 (N_44600,N_36645,N_36825);
or U44601 (N_44601,N_35937,N_35322);
or U44602 (N_44602,N_38823,N_38380);
xnor U44603 (N_44603,N_35289,N_36251);
nand U44604 (N_44604,N_37677,N_39576);
nor U44605 (N_44605,N_38524,N_39107);
or U44606 (N_44606,N_39408,N_37090);
nand U44607 (N_44607,N_37068,N_39400);
nand U44608 (N_44608,N_37624,N_37618);
xnor U44609 (N_44609,N_37774,N_38438);
nand U44610 (N_44610,N_38985,N_39049);
nand U44611 (N_44611,N_35485,N_39762);
and U44612 (N_44612,N_37427,N_38442);
or U44613 (N_44613,N_36271,N_39250);
xnor U44614 (N_44614,N_39074,N_37962);
nor U44615 (N_44615,N_37890,N_39433);
or U44616 (N_44616,N_35406,N_37276);
nor U44617 (N_44617,N_39967,N_38418);
nor U44618 (N_44618,N_39495,N_36690);
nand U44619 (N_44619,N_38004,N_37054);
nand U44620 (N_44620,N_38648,N_35908);
and U44621 (N_44621,N_36905,N_36446);
and U44622 (N_44622,N_35099,N_38338);
nor U44623 (N_44623,N_36148,N_37675);
nand U44624 (N_44624,N_39331,N_35055);
or U44625 (N_44625,N_38658,N_36956);
and U44626 (N_44626,N_37283,N_35937);
and U44627 (N_44627,N_37450,N_38288);
xnor U44628 (N_44628,N_37826,N_35444);
and U44629 (N_44629,N_39312,N_35552);
and U44630 (N_44630,N_37124,N_38115);
nand U44631 (N_44631,N_36645,N_36993);
xor U44632 (N_44632,N_38162,N_37676);
and U44633 (N_44633,N_38106,N_39238);
xnor U44634 (N_44634,N_37435,N_38089);
nand U44635 (N_44635,N_39914,N_37777);
nand U44636 (N_44636,N_38382,N_37061);
nor U44637 (N_44637,N_36980,N_37679);
xnor U44638 (N_44638,N_36680,N_35009);
or U44639 (N_44639,N_39149,N_37690);
and U44640 (N_44640,N_39656,N_36659);
nand U44641 (N_44641,N_36691,N_39798);
and U44642 (N_44642,N_39579,N_39206);
nor U44643 (N_44643,N_35529,N_36934);
and U44644 (N_44644,N_36004,N_37232);
nor U44645 (N_44645,N_35340,N_35787);
nor U44646 (N_44646,N_39765,N_37192);
nor U44647 (N_44647,N_39271,N_38983);
and U44648 (N_44648,N_36832,N_38777);
nor U44649 (N_44649,N_39199,N_39354);
nand U44650 (N_44650,N_37673,N_38860);
and U44651 (N_44651,N_35079,N_38956);
and U44652 (N_44652,N_36600,N_38882);
nor U44653 (N_44653,N_35997,N_38313);
nand U44654 (N_44654,N_37843,N_39338);
and U44655 (N_44655,N_35244,N_35719);
and U44656 (N_44656,N_39321,N_36675);
nand U44657 (N_44657,N_35603,N_39636);
nor U44658 (N_44658,N_36343,N_35870);
nand U44659 (N_44659,N_38950,N_38361);
or U44660 (N_44660,N_38257,N_36834);
and U44661 (N_44661,N_38522,N_39421);
nand U44662 (N_44662,N_35096,N_38664);
nand U44663 (N_44663,N_39119,N_35731);
nand U44664 (N_44664,N_37181,N_38048);
nor U44665 (N_44665,N_37152,N_38097);
nor U44666 (N_44666,N_37444,N_36968);
and U44667 (N_44667,N_35232,N_36931);
xnor U44668 (N_44668,N_38600,N_35308);
or U44669 (N_44669,N_37958,N_37832);
or U44670 (N_44670,N_39713,N_39688);
or U44671 (N_44671,N_39979,N_39202);
nor U44672 (N_44672,N_36459,N_38893);
nand U44673 (N_44673,N_37128,N_35709);
nor U44674 (N_44674,N_38238,N_39076);
nand U44675 (N_44675,N_35208,N_37862);
nor U44676 (N_44676,N_38769,N_35635);
or U44677 (N_44677,N_39410,N_36682);
or U44678 (N_44678,N_37966,N_38384);
nand U44679 (N_44679,N_36317,N_37663);
nor U44680 (N_44680,N_39547,N_37210);
nor U44681 (N_44681,N_39106,N_39389);
nand U44682 (N_44682,N_38113,N_36749);
or U44683 (N_44683,N_39833,N_39486);
nand U44684 (N_44684,N_36418,N_39954);
nand U44685 (N_44685,N_37374,N_35800);
xor U44686 (N_44686,N_36952,N_35759);
nor U44687 (N_44687,N_37718,N_36422);
or U44688 (N_44688,N_38542,N_36949);
or U44689 (N_44689,N_38442,N_36475);
or U44690 (N_44690,N_39881,N_37754);
nor U44691 (N_44691,N_39548,N_36342);
and U44692 (N_44692,N_39437,N_36143);
and U44693 (N_44693,N_36955,N_38675);
nand U44694 (N_44694,N_38329,N_38880);
and U44695 (N_44695,N_37836,N_37488);
and U44696 (N_44696,N_35627,N_38345);
nor U44697 (N_44697,N_39795,N_36989);
nand U44698 (N_44698,N_39253,N_36479);
or U44699 (N_44699,N_38540,N_36746);
and U44700 (N_44700,N_39879,N_37581);
and U44701 (N_44701,N_38991,N_37186);
or U44702 (N_44702,N_36584,N_37307);
nand U44703 (N_44703,N_39673,N_36888);
nand U44704 (N_44704,N_38175,N_37350);
xor U44705 (N_44705,N_38841,N_36830);
nand U44706 (N_44706,N_35406,N_36375);
and U44707 (N_44707,N_37864,N_35207);
nor U44708 (N_44708,N_37747,N_39993);
xor U44709 (N_44709,N_37023,N_37732);
nand U44710 (N_44710,N_39671,N_36137);
nor U44711 (N_44711,N_36869,N_38248);
and U44712 (N_44712,N_36932,N_39148);
or U44713 (N_44713,N_39266,N_39020);
and U44714 (N_44714,N_39440,N_35106);
nand U44715 (N_44715,N_37412,N_35144);
and U44716 (N_44716,N_39522,N_38554);
and U44717 (N_44717,N_36203,N_36147);
nand U44718 (N_44718,N_36037,N_36714);
or U44719 (N_44719,N_39018,N_37019);
nand U44720 (N_44720,N_37981,N_35007);
nor U44721 (N_44721,N_36570,N_39862);
nand U44722 (N_44722,N_35947,N_38239);
xnor U44723 (N_44723,N_38058,N_36170);
and U44724 (N_44724,N_35617,N_35972);
nor U44725 (N_44725,N_39521,N_35025);
and U44726 (N_44726,N_38256,N_38222);
or U44727 (N_44727,N_36639,N_36825);
or U44728 (N_44728,N_35993,N_37691);
nor U44729 (N_44729,N_36231,N_36360);
nor U44730 (N_44730,N_39039,N_36377);
or U44731 (N_44731,N_35549,N_37384);
xor U44732 (N_44732,N_36703,N_36518);
xnor U44733 (N_44733,N_39378,N_35330);
or U44734 (N_44734,N_38405,N_38476);
or U44735 (N_44735,N_39829,N_37208);
and U44736 (N_44736,N_38544,N_37121);
and U44737 (N_44737,N_36185,N_36002);
nand U44738 (N_44738,N_35299,N_39922);
and U44739 (N_44739,N_35101,N_38798);
nand U44740 (N_44740,N_38497,N_36632);
and U44741 (N_44741,N_35187,N_39872);
or U44742 (N_44742,N_37581,N_37496);
nand U44743 (N_44743,N_39217,N_37077);
xor U44744 (N_44744,N_37806,N_39201);
nand U44745 (N_44745,N_37439,N_37354);
or U44746 (N_44746,N_39372,N_39979);
and U44747 (N_44747,N_39817,N_36069);
nand U44748 (N_44748,N_36765,N_39259);
or U44749 (N_44749,N_37936,N_36537);
nor U44750 (N_44750,N_36019,N_36340);
nand U44751 (N_44751,N_38261,N_39033);
nor U44752 (N_44752,N_36873,N_35344);
nor U44753 (N_44753,N_36777,N_35727);
nor U44754 (N_44754,N_36096,N_37065);
nand U44755 (N_44755,N_36205,N_38017);
and U44756 (N_44756,N_35818,N_37386);
and U44757 (N_44757,N_39476,N_35203);
xor U44758 (N_44758,N_38106,N_36911);
or U44759 (N_44759,N_37587,N_36132);
or U44760 (N_44760,N_35196,N_39324);
nand U44761 (N_44761,N_38755,N_37317);
and U44762 (N_44762,N_38183,N_37280);
or U44763 (N_44763,N_37636,N_35991);
nor U44764 (N_44764,N_36136,N_37425);
nand U44765 (N_44765,N_35606,N_39835);
nand U44766 (N_44766,N_36259,N_39145);
or U44767 (N_44767,N_39191,N_36336);
and U44768 (N_44768,N_37536,N_35848);
nor U44769 (N_44769,N_39064,N_38013);
xnor U44770 (N_44770,N_37118,N_38494);
and U44771 (N_44771,N_38105,N_38781);
nand U44772 (N_44772,N_36457,N_39299);
and U44773 (N_44773,N_39663,N_35070);
nand U44774 (N_44774,N_36189,N_37122);
xnor U44775 (N_44775,N_35167,N_37267);
and U44776 (N_44776,N_36207,N_35328);
or U44777 (N_44777,N_37684,N_38619);
nor U44778 (N_44778,N_39817,N_37841);
nor U44779 (N_44779,N_37449,N_35489);
and U44780 (N_44780,N_39284,N_35028);
nand U44781 (N_44781,N_37594,N_38603);
xor U44782 (N_44782,N_38226,N_39579);
xnor U44783 (N_44783,N_37883,N_35635);
nor U44784 (N_44784,N_36298,N_38559);
nor U44785 (N_44785,N_38541,N_36053);
and U44786 (N_44786,N_36858,N_38018);
and U44787 (N_44787,N_36990,N_35684);
xnor U44788 (N_44788,N_38660,N_35294);
xor U44789 (N_44789,N_35103,N_39220);
or U44790 (N_44790,N_35427,N_37118);
or U44791 (N_44791,N_38769,N_37281);
nor U44792 (N_44792,N_35896,N_35994);
and U44793 (N_44793,N_36484,N_39945);
nor U44794 (N_44794,N_38454,N_39889);
or U44795 (N_44795,N_35655,N_38339);
nor U44796 (N_44796,N_35172,N_35691);
xor U44797 (N_44797,N_38050,N_35071);
and U44798 (N_44798,N_35476,N_37291);
nand U44799 (N_44799,N_37114,N_37976);
nand U44800 (N_44800,N_39806,N_37377);
or U44801 (N_44801,N_36978,N_36814);
and U44802 (N_44802,N_38033,N_38908);
nor U44803 (N_44803,N_35862,N_35984);
nor U44804 (N_44804,N_38474,N_39850);
nand U44805 (N_44805,N_39446,N_37788);
or U44806 (N_44806,N_39182,N_38690);
and U44807 (N_44807,N_35128,N_36908);
nand U44808 (N_44808,N_35233,N_39615);
and U44809 (N_44809,N_39122,N_39441);
and U44810 (N_44810,N_36698,N_38503);
nor U44811 (N_44811,N_36438,N_37821);
nand U44812 (N_44812,N_35675,N_35615);
or U44813 (N_44813,N_36727,N_37873);
xor U44814 (N_44814,N_35616,N_39634);
or U44815 (N_44815,N_38858,N_39339);
nand U44816 (N_44816,N_35568,N_39277);
or U44817 (N_44817,N_38647,N_37066);
nand U44818 (N_44818,N_36547,N_38924);
xor U44819 (N_44819,N_37215,N_36321);
and U44820 (N_44820,N_38271,N_38632);
xor U44821 (N_44821,N_38490,N_36999);
or U44822 (N_44822,N_36161,N_38309);
nand U44823 (N_44823,N_38346,N_35744);
nor U44824 (N_44824,N_39799,N_38746);
nand U44825 (N_44825,N_36198,N_39408);
nor U44826 (N_44826,N_37298,N_37617);
or U44827 (N_44827,N_39981,N_35095);
and U44828 (N_44828,N_39595,N_36606);
xor U44829 (N_44829,N_36879,N_37999);
or U44830 (N_44830,N_37526,N_39873);
and U44831 (N_44831,N_39796,N_36453);
and U44832 (N_44832,N_37373,N_39415);
xor U44833 (N_44833,N_35185,N_39988);
nor U44834 (N_44834,N_39312,N_36519);
and U44835 (N_44835,N_37462,N_39008);
nor U44836 (N_44836,N_39608,N_36920);
nand U44837 (N_44837,N_37324,N_39506);
or U44838 (N_44838,N_37534,N_39302);
nand U44839 (N_44839,N_39451,N_39207);
xnor U44840 (N_44840,N_38655,N_38461);
nor U44841 (N_44841,N_38546,N_35656);
xnor U44842 (N_44842,N_39973,N_39652);
nor U44843 (N_44843,N_36157,N_37692);
and U44844 (N_44844,N_35417,N_38654);
and U44845 (N_44845,N_37763,N_39609);
or U44846 (N_44846,N_36902,N_37121);
xor U44847 (N_44847,N_39490,N_35894);
xor U44848 (N_44848,N_37326,N_35207);
xor U44849 (N_44849,N_37087,N_39477);
nor U44850 (N_44850,N_37529,N_36072);
nand U44851 (N_44851,N_35703,N_36409);
or U44852 (N_44852,N_38628,N_38140);
xor U44853 (N_44853,N_37503,N_37445);
or U44854 (N_44854,N_38498,N_36219);
nand U44855 (N_44855,N_36464,N_35481);
nor U44856 (N_44856,N_39830,N_36820);
or U44857 (N_44857,N_39998,N_37640);
xnor U44858 (N_44858,N_38089,N_36776);
nand U44859 (N_44859,N_39921,N_35324);
or U44860 (N_44860,N_38561,N_38803);
nor U44861 (N_44861,N_36161,N_37061);
xnor U44862 (N_44862,N_38043,N_36151);
nor U44863 (N_44863,N_37441,N_37778);
nand U44864 (N_44864,N_39384,N_37962);
or U44865 (N_44865,N_39941,N_38138);
nor U44866 (N_44866,N_37558,N_39943);
or U44867 (N_44867,N_37301,N_37719);
or U44868 (N_44868,N_36432,N_35829);
or U44869 (N_44869,N_39340,N_37470);
and U44870 (N_44870,N_35843,N_36017);
and U44871 (N_44871,N_38318,N_38877);
nand U44872 (N_44872,N_38179,N_38199);
or U44873 (N_44873,N_38448,N_35843);
nor U44874 (N_44874,N_36840,N_38261);
nand U44875 (N_44875,N_39283,N_37345);
and U44876 (N_44876,N_39187,N_35965);
and U44877 (N_44877,N_38506,N_35253);
or U44878 (N_44878,N_39256,N_39929);
nor U44879 (N_44879,N_37173,N_36168);
nand U44880 (N_44880,N_37331,N_35613);
and U44881 (N_44881,N_38758,N_38197);
or U44882 (N_44882,N_35502,N_39977);
and U44883 (N_44883,N_35734,N_35917);
nor U44884 (N_44884,N_35112,N_35301);
or U44885 (N_44885,N_39408,N_38435);
xnor U44886 (N_44886,N_36448,N_35049);
nor U44887 (N_44887,N_37125,N_35079);
or U44888 (N_44888,N_38050,N_36122);
nor U44889 (N_44889,N_39754,N_39153);
nor U44890 (N_44890,N_37305,N_39816);
nor U44891 (N_44891,N_37941,N_39981);
or U44892 (N_44892,N_37927,N_36446);
nor U44893 (N_44893,N_36884,N_37412);
or U44894 (N_44894,N_39601,N_37144);
nor U44895 (N_44895,N_37263,N_37431);
nand U44896 (N_44896,N_35940,N_36903);
and U44897 (N_44897,N_39536,N_35716);
nor U44898 (N_44898,N_37489,N_39494);
and U44899 (N_44899,N_37411,N_39656);
and U44900 (N_44900,N_37750,N_38508);
nand U44901 (N_44901,N_38660,N_36249);
nand U44902 (N_44902,N_37884,N_36620);
or U44903 (N_44903,N_39166,N_36165);
and U44904 (N_44904,N_37886,N_37726);
or U44905 (N_44905,N_36975,N_36295);
and U44906 (N_44906,N_36923,N_35332);
and U44907 (N_44907,N_37087,N_36974);
nor U44908 (N_44908,N_36331,N_38530);
and U44909 (N_44909,N_39263,N_35304);
or U44910 (N_44910,N_35072,N_36227);
nand U44911 (N_44911,N_35681,N_39261);
and U44912 (N_44912,N_37209,N_39022);
or U44913 (N_44913,N_38561,N_37917);
nor U44914 (N_44914,N_38242,N_36262);
and U44915 (N_44915,N_39406,N_38250);
xnor U44916 (N_44916,N_39327,N_37908);
and U44917 (N_44917,N_36020,N_35956);
nor U44918 (N_44918,N_37805,N_38847);
nor U44919 (N_44919,N_35572,N_35663);
nor U44920 (N_44920,N_38665,N_38191);
xnor U44921 (N_44921,N_36638,N_38678);
or U44922 (N_44922,N_39919,N_36981);
nor U44923 (N_44923,N_39786,N_36951);
and U44924 (N_44924,N_39125,N_38588);
nand U44925 (N_44925,N_36795,N_39197);
or U44926 (N_44926,N_35295,N_38661);
nand U44927 (N_44927,N_38184,N_36368);
or U44928 (N_44928,N_37000,N_35178);
or U44929 (N_44929,N_38960,N_35141);
or U44930 (N_44930,N_37437,N_39687);
or U44931 (N_44931,N_38945,N_36751);
and U44932 (N_44932,N_38090,N_39419);
and U44933 (N_44933,N_37586,N_36187);
nand U44934 (N_44934,N_35550,N_39212);
xnor U44935 (N_44935,N_36020,N_38203);
xor U44936 (N_44936,N_35713,N_36831);
or U44937 (N_44937,N_35566,N_39137);
xor U44938 (N_44938,N_37410,N_39206);
nor U44939 (N_44939,N_37951,N_35916);
nand U44940 (N_44940,N_38124,N_35050);
or U44941 (N_44941,N_35476,N_35162);
xor U44942 (N_44942,N_37869,N_36119);
nand U44943 (N_44943,N_37410,N_39601);
xnor U44944 (N_44944,N_36296,N_35554);
nor U44945 (N_44945,N_35761,N_39975);
and U44946 (N_44946,N_38898,N_39356);
xnor U44947 (N_44947,N_38898,N_36416);
and U44948 (N_44948,N_38715,N_39656);
or U44949 (N_44949,N_36126,N_38642);
or U44950 (N_44950,N_37831,N_39802);
and U44951 (N_44951,N_35965,N_35385);
or U44952 (N_44952,N_39721,N_38054);
and U44953 (N_44953,N_38020,N_38884);
nand U44954 (N_44954,N_37764,N_37874);
nand U44955 (N_44955,N_36286,N_39838);
nand U44956 (N_44956,N_36140,N_36972);
or U44957 (N_44957,N_36868,N_35174);
or U44958 (N_44958,N_38353,N_38231);
nor U44959 (N_44959,N_37863,N_39212);
and U44960 (N_44960,N_38711,N_39773);
nand U44961 (N_44961,N_35664,N_39691);
and U44962 (N_44962,N_37659,N_37528);
xor U44963 (N_44963,N_36348,N_36796);
and U44964 (N_44964,N_36267,N_36298);
xor U44965 (N_44965,N_37164,N_38943);
or U44966 (N_44966,N_37341,N_35664);
or U44967 (N_44967,N_38578,N_38932);
nand U44968 (N_44968,N_35923,N_37544);
nor U44969 (N_44969,N_36381,N_38079);
and U44970 (N_44970,N_36533,N_36326);
and U44971 (N_44971,N_39061,N_37195);
nor U44972 (N_44972,N_36227,N_36460);
nand U44973 (N_44973,N_39674,N_39806);
nand U44974 (N_44974,N_38774,N_38988);
nor U44975 (N_44975,N_35122,N_38467);
nand U44976 (N_44976,N_39005,N_35177);
nand U44977 (N_44977,N_37903,N_38313);
and U44978 (N_44978,N_35742,N_37875);
nand U44979 (N_44979,N_37472,N_37376);
nand U44980 (N_44980,N_35005,N_38696);
and U44981 (N_44981,N_38250,N_35886);
nand U44982 (N_44982,N_37602,N_37316);
nand U44983 (N_44983,N_36079,N_35836);
and U44984 (N_44984,N_39956,N_36769);
or U44985 (N_44985,N_39215,N_36504);
nand U44986 (N_44986,N_35716,N_35040);
and U44987 (N_44987,N_35562,N_38002);
nand U44988 (N_44988,N_37887,N_37843);
nand U44989 (N_44989,N_35996,N_35771);
or U44990 (N_44990,N_35240,N_36692);
nand U44991 (N_44991,N_37660,N_38714);
and U44992 (N_44992,N_35732,N_36763);
xnor U44993 (N_44993,N_37339,N_36905);
nor U44994 (N_44994,N_35923,N_38942);
xnor U44995 (N_44995,N_38780,N_35529);
and U44996 (N_44996,N_36976,N_35643);
nand U44997 (N_44997,N_37590,N_39422);
and U44998 (N_44998,N_39244,N_36710);
nor U44999 (N_44999,N_37967,N_35952);
and U45000 (N_45000,N_42668,N_44267);
nand U45001 (N_45001,N_40649,N_44289);
nor U45002 (N_45002,N_42860,N_43216);
xnor U45003 (N_45003,N_42269,N_40928);
nor U45004 (N_45004,N_43133,N_43249);
nand U45005 (N_45005,N_44390,N_42270);
nand U45006 (N_45006,N_44833,N_42471);
xor U45007 (N_45007,N_41610,N_41432);
and U45008 (N_45008,N_40781,N_41112);
xor U45009 (N_45009,N_42709,N_41310);
and U45010 (N_45010,N_41061,N_43821);
xnor U45011 (N_45011,N_40432,N_41915);
nand U45012 (N_45012,N_42904,N_43381);
or U45013 (N_45013,N_42392,N_40336);
nand U45014 (N_45014,N_40199,N_42383);
or U45015 (N_45015,N_41047,N_44481);
or U45016 (N_45016,N_44611,N_44311);
or U45017 (N_45017,N_40114,N_42289);
nor U45018 (N_45018,N_42408,N_44728);
and U45019 (N_45019,N_44220,N_41784);
xnor U45020 (N_45020,N_42262,N_40802);
nand U45021 (N_45021,N_42726,N_41360);
nand U45022 (N_45022,N_44351,N_43591);
nor U45023 (N_45023,N_40506,N_42093);
nand U45024 (N_45024,N_43695,N_44786);
or U45025 (N_45025,N_41617,N_41353);
nand U45026 (N_45026,N_40870,N_41918);
and U45027 (N_45027,N_44010,N_44489);
xor U45028 (N_45028,N_41947,N_42189);
or U45029 (N_45029,N_40899,N_41141);
nand U45030 (N_45030,N_44757,N_41337);
nand U45031 (N_45031,N_44046,N_41491);
nand U45032 (N_45032,N_42130,N_44434);
nand U45033 (N_45033,N_44837,N_42237);
or U45034 (N_45034,N_41672,N_42572);
nand U45035 (N_45035,N_41503,N_41127);
nor U45036 (N_45036,N_41680,N_40049);
or U45037 (N_45037,N_43666,N_42939);
nor U45038 (N_45038,N_43322,N_43972);
nor U45039 (N_45039,N_42509,N_43284);
nor U45040 (N_45040,N_41832,N_43977);
nor U45041 (N_45041,N_41072,N_44115);
xor U45042 (N_45042,N_40479,N_42250);
or U45043 (N_45043,N_40373,N_43464);
or U45044 (N_45044,N_44034,N_43251);
nand U45045 (N_45045,N_44697,N_43014);
or U45046 (N_45046,N_40382,N_42979);
nor U45047 (N_45047,N_40339,N_40012);
or U45048 (N_45048,N_42334,N_42720);
nand U45049 (N_45049,N_42527,N_42162);
and U45050 (N_45050,N_40723,N_43350);
and U45051 (N_45051,N_44737,N_42885);
or U45052 (N_45052,N_42390,N_40371);
nand U45053 (N_45053,N_44810,N_44500);
nand U45054 (N_45054,N_40510,N_41845);
xor U45055 (N_45055,N_41062,N_40182);
and U45056 (N_45056,N_42278,N_43910);
xor U45057 (N_45057,N_42481,N_40175);
and U45058 (N_45058,N_40849,N_44771);
nand U45059 (N_45059,N_43810,N_44042);
nor U45060 (N_45060,N_41975,N_43008);
nor U45061 (N_45061,N_42654,N_43545);
nand U45062 (N_45062,N_40467,N_42877);
nand U45063 (N_45063,N_41297,N_42974);
and U45064 (N_45064,N_40514,N_43414);
nor U45065 (N_45065,N_40078,N_40484);
nand U45066 (N_45066,N_43167,N_42550);
nand U45067 (N_45067,N_44406,N_41614);
or U45068 (N_45068,N_43162,N_44859);
nor U45069 (N_45069,N_40240,N_43633);
nor U45070 (N_45070,N_42741,N_41681);
and U45071 (N_45071,N_43253,N_44172);
and U45072 (N_45072,N_42111,N_41490);
nand U45073 (N_45073,N_43484,N_41073);
nor U45074 (N_45074,N_44234,N_40380);
nor U45075 (N_45075,N_43246,N_43646);
and U45076 (N_45076,N_44646,N_42861);
nand U45077 (N_45077,N_40695,N_40197);
nor U45078 (N_45078,N_42625,N_42920);
or U45079 (N_45079,N_42629,N_40153);
or U45080 (N_45080,N_40693,N_42495);
nand U45081 (N_45081,N_44124,N_43779);
or U45082 (N_45082,N_42838,N_40862);
nand U45083 (N_45083,N_41669,N_41540);
and U45084 (N_45084,N_40905,N_43443);
or U45085 (N_45085,N_40566,N_43039);
nor U45086 (N_45086,N_42683,N_44482);
nor U45087 (N_45087,N_40670,N_40256);
nor U45088 (N_45088,N_40702,N_42395);
xor U45089 (N_45089,N_40356,N_43847);
and U45090 (N_45090,N_42248,N_42680);
nand U45091 (N_45091,N_42283,N_44412);
nand U45092 (N_45092,N_41858,N_43586);
nand U45093 (N_45093,N_41560,N_41694);
or U45094 (N_45094,N_42514,N_44447);
or U45095 (N_45095,N_43544,N_44448);
nand U45096 (N_45096,N_40401,N_40044);
or U45097 (N_45097,N_40863,N_42733);
xor U45098 (N_45098,N_40694,N_42833);
or U45099 (N_45099,N_40374,N_44151);
nand U45100 (N_45100,N_41951,N_40599);
or U45101 (N_45101,N_44385,N_44636);
or U45102 (N_45102,N_40174,N_42863);
xor U45103 (N_45103,N_40605,N_40508);
and U45104 (N_45104,N_43129,N_44730);
nand U45105 (N_45105,N_44329,N_41654);
or U45106 (N_45106,N_41087,N_42094);
nand U45107 (N_45107,N_44118,N_43675);
xnor U45108 (N_45108,N_41382,N_43837);
nor U45109 (N_45109,N_41471,N_42449);
nand U45110 (N_45110,N_42172,N_44497);
nand U45111 (N_45111,N_43200,N_43423);
nand U45112 (N_45112,N_40700,N_41443);
or U45113 (N_45113,N_43513,N_41467);
nand U45114 (N_45114,N_41211,N_43025);
nand U45115 (N_45115,N_42988,N_42272);
nand U45116 (N_45116,N_42561,N_42779);
nand U45117 (N_45117,N_41027,N_42465);
nor U45118 (N_45118,N_43517,N_43092);
and U45119 (N_45119,N_43393,N_44718);
or U45120 (N_45120,N_40053,N_41758);
or U45121 (N_45121,N_41812,N_41293);
nand U45122 (N_45122,N_44335,N_43786);
or U45123 (N_45123,N_43702,N_41457);
nand U45124 (N_45124,N_42052,N_40701);
nor U45125 (N_45125,N_41991,N_41330);
nor U45126 (N_45126,N_41469,N_43324);
or U45127 (N_45127,N_43378,N_40833);
nor U45128 (N_45128,N_41902,N_41049);
nor U45129 (N_45129,N_41253,N_44022);
nand U45130 (N_45130,N_42126,N_41071);
nand U45131 (N_45131,N_44824,N_44751);
or U45132 (N_45132,N_42403,N_40455);
nor U45133 (N_45133,N_40419,N_41252);
or U45134 (N_45134,N_43035,N_41786);
nor U45135 (N_45135,N_41871,N_40593);
or U45136 (N_45136,N_43303,N_41348);
and U45137 (N_45137,N_43237,N_41880);
or U45138 (N_45138,N_41128,N_44624);
or U45139 (N_45139,N_41700,N_40301);
nor U45140 (N_45140,N_40763,N_42590);
and U45141 (N_45141,N_40769,N_40105);
and U45142 (N_45142,N_41114,N_42016);
nand U45143 (N_45143,N_42326,N_42540);
nand U45144 (N_45144,N_42933,N_43439);
nor U45145 (N_45145,N_43145,N_40706);
xor U45146 (N_45146,N_41411,N_43996);
or U45147 (N_45147,N_41006,N_42619);
nand U45148 (N_45148,N_41744,N_44093);
or U45149 (N_45149,N_44997,N_43233);
and U45150 (N_45150,N_41030,N_40116);
or U45151 (N_45151,N_43763,N_40493);
or U45152 (N_45152,N_42841,N_42084);
nand U45153 (N_45153,N_41924,N_43385);
or U45154 (N_45154,N_42277,N_44572);
or U45155 (N_45155,N_41788,N_42185);
xor U45156 (N_45156,N_44382,N_40210);
or U45157 (N_45157,N_41295,N_44747);
nand U45158 (N_45158,N_43291,N_41693);
nor U45159 (N_45159,N_41985,N_44127);
nand U45160 (N_45160,N_40363,N_40201);
nor U45161 (N_45161,N_41584,N_44141);
and U45162 (N_45162,N_40840,N_40585);
nand U45163 (N_45163,N_43552,N_43641);
nor U45164 (N_45164,N_40619,N_40686);
nand U45165 (N_45165,N_44047,N_44138);
and U45166 (N_45166,N_40509,N_44806);
xnor U45167 (N_45167,N_42346,N_42207);
nor U45168 (N_45168,N_44764,N_40555);
nor U45169 (N_45169,N_43240,N_42835);
or U45170 (N_45170,N_40716,N_41731);
nand U45171 (N_45171,N_40690,N_44357);
nor U45172 (N_45172,N_42402,N_41450);
and U45173 (N_45173,N_43730,N_44887);
xor U45174 (N_45174,N_42115,N_40047);
nand U45175 (N_45175,N_40776,N_42282);
nand U45176 (N_45176,N_44606,N_44043);
nand U45177 (N_45177,N_42364,N_44233);
and U45178 (N_45178,N_41148,N_43928);
nor U45179 (N_45179,N_43458,N_41419);
or U45180 (N_45180,N_42071,N_40657);
nor U45181 (N_45181,N_40018,N_42826);
nor U45182 (N_45182,N_43841,N_42870);
xnor U45183 (N_45183,N_41369,N_43022);
nor U45184 (N_45184,N_43040,N_41123);
and U45185 (N_45185,N_43561,N_43640);
or U45186 (N_45186,N_40545,N_44437);
and U45187 (N_45187,N_43018,N_44483);
and U45188 (N_45188,N_41989,N_42483);
nand U45189 (N_45189,N_41271,N_41395);
and U45190 (N_45190,N_41955,N_44014);
nor U45191 (N_45191,N_44760,N_43319);
and U45192 (N_45192,N_42158,N_42213);
and U45193 (N_45193,N_44867,N_40359);
or U45194 (N_45194,N_41359,N_41587);
or U45195 (N_45195,N_44809,N_43485);
nand U45196 (N_45196,N_42096,N_40696);
and U45197 (N_45197,N_41098,N_41785);
nand U45198 (N_45198,N_44802,N_42467);
nand U45199 (N_45199,N_43880,N_40972);
and U45200 (N_45200,N_44858,N_40570);
nand U45201 (N_45201,N_41964,N_44963);
nor U45202 (N_45202,N_42500,N_42719);
or U45203 (N_45203,N_41708,N_44324);
nand U45204 (N_45204,N_43542,N_40331);
or U45205 (N_45205,N_42916,N_44977);
nor U45206 (N_45206,N_43348,N_40635);
nand U45207 (N_45207,N_43583,N_44076);
or U45208 (N_45208,N_40150,N_42448);
or U45209 (N_45209,N_42425,N_40154);
and U45210 (N_45210,N_44666,N_42214);
or U45211 (N_45211,N_44223,N_43150);
nand U45212 (N_45212,N_40066,N_44095);
xnor U45213 (N_45213,N_43699,N_42663);
or U45214 (N_45214,N_40854,N_41231);
nand U45215 (N_45215,N_44574,N_41966);
and U45216 (N_45216,N_42792,N_40028);
or U45217 (N_45217,N_44733,N_43355);
and U45218 (N_45218,N_42301,N_44558);
and U45219 (N_45219,N_43416,N_41505);
and U45220 (N_45220,N_40492,N_42636);
xnor U45221 (N_45221,N_42644,N_42868);
and U45222 (N_45222,N_42643,N_40760);
and U45223 (N_45223,N_41579,N_41203);
and U45224 (N_45224,N_43153,N_40722);
xnor U45225 (N_45225,N_41718,N_41398);
and U45226 (N_45226,N_44994,N_41861);
nand U45227 (N_45227,N_40513,N_44071);
and U45228 (N_45228,N_42110,N_42837);
nor U45229 (N_45229,N_44726,N_41798);
nor U45230 (N_45230,N_41448,N_41605);
nor U45231 (N_45231,N_42678,N_40512);
nor U45232 (N_45232,N_41023,N_43475);
xnor U45233 (N_45233,N_41140,N_41220);
nor U45234 (N_45234,N_44471,N_43002);
or U45235 (N_45235,N_43364,N_42795);
nand U45236 (N_45236,N_43985,N_43108);
and U45237 (N_45237,N_43208,N_42241);
and U45238 (N_45238,N_41981,N_40177);
nor U45239 (N_45239,N_40771,N_43907);
or U45240 (N_45240,N_44173,N_40604);
nand U45241 (N_45241,N_42975,N_40612);
nor U45242 (N_45242,N_44620,N_40887);
and U45243 (N_45243,N_43718,N_42151);
or U45244 (N_45244,N_43879,N_42537);
nor U45245 (N_45245,N_40495,N_44560);
or U45246 (N_45246,N_44193,N_40710);
nor U45247 (N_45247,N_40837,N_44523);
or U45248 (N_45248,N_43941,N_44421);
and U45249 (N_45249,N_43234,N_42704);
nor U45250 (N_45250,N_40647,N_43719);
nor U45251 (N_45251,N_41494,N_43388);
nor U45252 (N_45252,N_44298,N_44563);
or U45253 (N_45253,N_42027,N_44512);
nor U45254 (N_45254,N_40788,N_41037);
or U45255 (N_45255,N_42290,N_43321);
nand U45256 (N_45256,N_41263,N_44546);
xor U45257 (N_45257,N_42763,N_43871);
or U45258 (N_45258,N_43973,N_43156);
and U45259 (N_45259,N_40191,N_40074);
and U45260 (N_45260,N_41038,N_42356);
or U45261 (N_45261,N_42171,N_40357);
and U45262 (N_45262,N_43128,N_40660);
nand U45263 (N_45263,N_41408,N_44433);
nand U45264 (N_45264,N_41439,N_44675);
nor U45265 (N_45265,N_42281,N_43235);
or U45266 (N_45266,N_43688,N_41129);
and U45267 (N_45267,N_40257,N_41586);
nor U45268 (N_45268,N_42794,N_41018);
and U45269 (N_45269,N_43952,N_42845);
and U45270 (N_45270,N_44229,N_44402);
and U45271 (N_45271,N_40521,N_40424);
nand U45272 (N_45272,N_43878,N_42308);
nor U45273 (N_45273,N_41775,N_43791);
nor U45274 (N_45274,N_44580,N_42535);
or U45275 (N_45275,N_43992,N_40317);
nand U45276 (N_45276,N_44307,N_41113);
and U45277 (N_45277,N_41233,N_41637);
nor U45278 (N_45278,N_44603,N_42157);
nor U45279 (N_45279,N_42140,N_40857);
or U45280 (N_45280,N_42932,N_40775);
nor U45281 (N_45281,N_44919,N_44792);
and U45282 (N_45282,N_42989,N_41527);
nor U45283 (N_45283,N_43477,N_44197);
and U45284 (N_45284,N_40157,N_41909);
and U45285 (N_45285,N_40135,N_41533);
and U45286 (N_45286,N_43778,N_43957);
and U45287 (N_45287,N_42995,N_42637);
and U45288 (N_45288,N_42080,N_42492);
nand U45289 (N_45289,N_42341,N_41660);
nor U45290 (N_45290,N_43174,N_41109);
nor U45291 (N_45291,N_40740,N_44505);
nand U45292 (N_45292,N_41982,N_40181);
or U45293 (N_45293,N_44213,N_41815);
and U45294 (N_45294,N_41623,N_42472);
nor U45295 (N_45295,N_42015,N_41967);
and U45296 (N_45296,N_44575,N_43021);
nand U45297 (N_45297,N_44460,N_44426);
or U45298 (N_45298,N_44356,N_40103);
and U45299 (N_45299,N_44189,N_41522);
and U45300 (N_45300,N_40858,N_44021);
or U45301 (N_45301,N_44050,N_43041);
nand U45302 (N_45302,N_42307,N_43132);
nand U45303 (N_45303,N_41422,N_40993);
and U45304 (N_45304,N_40678,N_41250);
nand U45305 (N_45305,N_40451,N_44626);
nand U45306 (N_45306,N_42755,N_44451);
and U45307 (N_45307,N_44701,N_44129);
nand U45308 (N_45308,N_44130,N_43333);
nand U45309 (N_45309,N_41963,N_44036);
nor U45310 (N_45310,N_42155,N_43375);
nor U45311 (N_45311,N_40960,N_43672);
xor U45312 (N_45312,N_40312,N_40264);
and U45313 (N_45313,N_44265,N_42173);
nor U45314 (N_45314,N_43437,N_44400);
and U45315 (N_45315,N_42331,N_41303);
or U45316 (N_45316,N_44849,N_44058);
and U45317 (N_45317,N_40294,N_40020);
and U45318 (N_45318,N_41414,N_43680);
or U45319 (N_45319,N_43192,N_42548);
nor U45320 (N_45320,N_44270,N_44261);
or U45321 (N_45321,N_40941,N_44855);
or U45322 (N_45322,N_41142,N_43593);
or U45323 (N_45323,N_41001,N_41756);
nand U45324 (N_45324,N_41447,N_43310);
or U45325 (N_45325,N_42252,N_42413);
nand U45326 (N_45326,N_43600,N_40202);
xor U45327 (N_45327,N_44584,N_44670);
nand U45328 (N_45328,N_41661,N_40507);
nand U45329 (N_45329,N_41243,N_40543);
or U45330 (N_45330,N_40810,N_43667);
nand U45331 (N_45331,N_42831,N_44540);
nor U45332 (N_45332,N_40785,N_43406);
or U45333 (N_45333,N_40586,N_44738);
nor U45334 (N_45334,N_43078,N_40239);
xor U45335 (N_45335,N_41644,N_44326);
xor U45336 (N_45336,N_43172,N_43171);
or U45337 (N_45337,N_42264,N_40265);
xnor U45338 (N_45338,N_40664,N_42693);
nand U45339 (N_45339,N_40395,N_44878);
nand U45340 (N_45340,N_41782,N_43466);
or U45341 (N_45341,N_43264,N_42562);
nor U45342 (N_45342,N_43797,N_41843);
and U45343 (N_45343,N_42638,N_42287);
xnor U45344 (N_45344,N_40063,N_40859);
or U45345 (N_45345,N_41558,N_41913);
and U45346 (N_45346,N_42303,N_41528);
and U45347 (N_45347,N_42856,N_40458);
or U45348 (N_45348,N_40035,N_42593);
nand U45349 (N_45349,N_42817,N_42765);
or U45350 (N_45350,N_41488,N_40703);
nand U45351 (N_45351,N_43061,N_42339);
or U45352 (N_45352,N_44669,N_40290);
or U45353 (N_45353,N_41688,N_41927);
nor U45354 (N_45354,N_43734,N_44827);
nor U45355 (N_45355,N_40777,N_41556);
and U45356 (N_45356,N_44643,N_42288);
nand U45357 (N_45357,N_41514,N_42824);
and U45358 (N_45358,N_41264,N_42642);
nand U45359 (N_45359,N_43570,N_44705);
or U45360 (N_45360,N_44539,N_41853);
nand U45361 (N_45361,N_44692,N_42051);
or U45362 (N_45362,N_44325,N_40141);
nand U45363 (N_45363,N_41232,N_43795);
xor U45364 (N_45364,N_40921,N_43564);
and U45365 (N_45365,N_44299,N_44055);
xor U45366 (N_45366,N_42474,N_43653);
nand U45367 (N_45367,N_43009,N_41643);
nand U45368 (N_45368,N_40821,N_42225);
nand U45369 (N_45369,N_40937,N_44935);
xnor U45370 (N_45370,N_44815,N_42597);
or U45371 (N_45371,N_43494,N_42091);
and U45372 (N_45372,N_44717,N_44340);
or U45373 (N_45373,N_43279,N_41498);
xnor U45374 (N_45374,N_43186,N_44012);
xnor U45375 (N_45375,N_43247,N_43305);
and U45376 (N_45376,N_43384,N_44135);
nor U45377 (N_45377,N_43343,N_40789);
xor U45378 (N_45378,N_43290,N_40940);
nor U45379 (N_45379,N_41905,N_40292);
xor U45380 (N_45380,N_40542,N_42019);
and U45381 (N_45381,N_43742,N_44968);
nand U45382 (N_45382,N_43571,N_40146);
and U45383 (N_45383,N_41230,N_43121);
nand U45384 (N_45384,N_40297,N_42820);
nand U45385 (N_45385,N_44156,N_40911);
and U45386 (N_45386,N_41965,N_40813);
nor U45387 (N_45387,N_41324,N_44667);
nand U45388 (N_45388,N_42120,N_42442);
nor U45389 (N_45389,N_43913,N_41435);
and U45390 (N_45390,N_44085,N_42312);
nor U45391 (N_45391,N_44134,N_43839);
nand U45392 (N_45392,N_41604,N_44147);
xnor U45393 (N_45393,N_43610,N_42022);
nor U45394 (N_45394,N_43851,N_42790);
xor U45395 (N_45395,N_42460,N_43187);
nand U45396 (N_45396,N_43325,N_40398);
or U45397 (N_45397,N_42466,N_40529);
nand U45398 (N_45398,N_42055,N_40828);
and U45399 (N_45399,N_42918,N_43266);
or U45400 (N_45400,N_41002,N_41375);
or U45401 (N_45401,N_41607,N_42108);
xor U45402 (N_45402,N_44182,N_42623);
and U45403 (N_45403,N_42752,N_44936);
nand U45404 (N_45404,N_40107,N_43520);
or U45405 (N_45405,N_43862,N_40076);
and U45406 (N_45406,N_40127,N_43756);
xor U45407 (N_45407,N_44231,N_43920);
xnor U45408 (N_45408,N_41169,N_40073);
or U45409 (N_45409,N_43374,N_44463);
xnor U45410 (N_45410,N_41885,N_42142);
and U45411 (N_45411,N_44762,N_43226);
or U45412 (N_45412,N_43575,N_42854);
nor U45413 (N_45413,N_41152,N_43062);
nor U45414 (N_45414,N_44474,N_42182);
nor U45415 (N_45415,N_44048,N_40386);
xnor U45416 (N_45416,N_40621,N_44080);
nor U45417 (N_45417,N_40303,N_40947);
nor U45418 (N_45418,N_44376,N_41238);
nor U45419 (N_45419,N_41801,N_44821);
nor U45420 (N_45420,N_43842,N_44553);
and U45421 (N_45421,N_40081,N_44441);
and U45422 (N_45422,N_44891,N_43579);
or U45423 (N_45423,N_42422,N_44982);
or U45424 (N_45424,N_41338,N_41642);
or U45425 (N_45425,N_41468,N_41921);
and U45426 (N_45426,N_44978,N_42266);
or U45427 (N_45427,N_40335,N_44257);
or U45428 (N_45428,N_40511,N_44254);
and U45429 (N_45429,N_41896,N_40932);
nand U45430 (N_45430,N_40861,N_41248);
or U45431 (N_45431,N_44202,N_40739);
and U45432 (N_45432,N_44165,N_44845);
or U45433 (N_45433,N_41547,N_41466);
or U45434 (N_45434,N_44423,N_44455);
and U45435 (N_45435,N_40096,N_42586);
nor U45436 (N_45436,N_40643,N_44723);
nor U45437 (N_45437,N_43399,N_43684);
nand U45438 (N_45438,N_43835,N_40125);
nor U45439 (N_45439,N_44088,N_42991);
nor U45440 (N_45440,N_43984,N_40222);
nand U45441 (N_45441,N_40938,N_40563);
nor U45442 (N_45442,N_43244,N_42005);
or U45443 (N_45443,N_42786,N_40169);
nand U45444 (N_45444,N_42784,N_40929);
nor U45445 (N_45445,N_43448,N_41461);
xor U45446 (N_45446,N_44164,N_42063);
or U45447 (N_45447,N_42292,N_43396);
nor U45448 (N_45448,N_40594,N_40254);
or U45449 (N_45449,N_40629,N_41502);
or U45450 (N_45450,N_43904,N_44627);
nand U45451 (N_45451,N_41600,N_42100);
xor U45452 (N_45452,N_41485,N_44567);
nand U45453 (N_45453,N_44053,N_40882);
xnor U45454 (N_45454,N_41313,N_42706);
nand U45455 (N_45455,N_43714,N_43619);
nand U45456 (N_45456,N_40128,N_43481);
and U45457 (N_45457,N_44794,N_42891);
nor U45458 (N_45458,N_44618,N_43769);
and U45459 (N_45459,N_43711,N_44354);
or U45460 (N_45460,N_43772,N_40520);
or U45461 (N_45461,N_41275,N_43678);
nor U45462 (N_45462,N_42197,N_41524);
nand U45463 (N_45463,N_44541,N_41569);
or U45464 (N_45464,N_40568,N_41059);
xnor U45465 (N_45465,N_40001,N_41279);
xnor U45466 (N_45466,N_42404,N_44029);
nor U45467 (N_45467,N_42816,N_40403);
nand U45468 (N_45468,N_44647,N_41489);
or U45469 (N_45469,N_42046,N_40446);
nand U45470 (N_45470,N_42525,N_42216);
and U45471 (N_45471,N_40874,N_42138);
or U45472 (N_45472,N_42992,N_40799);
or U45473 (N_45473,N_43055,N_43151);
nor U45474 (N_45474,N_41299,N_44075);
and U45475 (N_45475,N_40577,N_43152);
nor U45476 (N_45476,N_44305,N_44739);
xnor U45477 (N_45477,N_43277,N_41652);
nand U45478 (N_45478,N_44370,N_44347);
and U45479 (N_45479,N_43193,N_40343);
nand U45480 (N_45480,N_40286,N_41609);
xnor U45481 (N_45481,N_41629,N_42295);
and U45482 (N_45482,N_43456,N_41907);
and U45483 (N_45483,N_40348,N_43894);
nor U45484 (N_45484,N_42223,N_41311);
or U45485 (N_45485,N_41176,N_42737);
xnor U45486 (N_45486,N_41070,N_44149);
or U45487 (N_45487,N_42567,N_40110);
and U45488 (N_45488,N_43721,N_42416);
or U45489 (N_45489,N_43955,N_42691);
or U45490 (N_45490,N_44787,N_40637);
nand U45491 (N_45491,N_41983,N_42280);
and U45492 (N_45492,N_42017,N_41575);
nand U45493 (N_45493,N_44664,N_43093);
nor U45494 (N_45494,N_41576,N_44974);
xor U45495 (N_45495,N_42595,N_42388);
xor U45496 (N_45496,N_43154,N_43969);
nand U45497 (N_45497,N_43001,N_43124);
or U45498 (N_45498,N_40644,N_42166);
xor U45499 (N_45499,N_40425,N_42066);
nor U45500 (N_45500,N_44744,N_43256);
or U45501 (N_45501,N_42074,N_42233);
nor U45502 (N_45502,N_44017,N_42164);
and U45503 (N_45503,N_40838,N_40052);
nor U45504 (N_45504,N_44511,N_44296);
and U45505 (N_45505,N_40600,N_41665);
xor U45506 (N_45506,N_42268,N_41630);
or U45507 (N_45507,N_41701,N_40360);
nand U45508 (N_45508,N_40868,N_40477);
nand U45509 (N_45509,N_43692,N_41667);
and U45510 (N_45510,N_42545,N_44321);
nand U45511 (N_45511,N_41890,N_42532);
xnor U45512 (N_45512,N_41396,N_41732);
or U45513 (N_45513,N_43671,N_43787);
nand U45514 (N_45514,N_41992,N_44896);
or U45515 (N_45515,N_43352,N_43134);
nor U45516 (N_45516,N_44926,N_41988);
nor U45517 (N_45517,N_44294,N_40136);
and U45518 (N_45518,N_44429,N_41133);
nor U45519 (N_45519,N_44313,N_44623);
and U45520 (N_45520,N_42895,N_44244);
and U45521 (N_45521,N_42081,N_43854);
xor U45522 (N_45522,N_40801,N_42818);
nor U45523 (N_45523,N_42659,N_42753);
nand U45524 (N_45524,N_44625,N_42323);
nand U45525 (N_45525,N_43814,N_43726);
or U45526 (N_45526,N_40640,N_43367);
or U45527 (N_45527,N_40697,N_42611);
nand U45528 (N_45528,N_44372,N_43824);
nor U45529 (N_45529,N_41523,N_40148);
xor U45530 (N_45530,N_42137,N_40783);
nand U45531 (N_45531,N_40087,N_44142);
and U45532 (N_45532,N_43991,N_44418);
nand U45533 (N_45533,N_42570,N_40654);
or U45534 (N_45534,N_41096,N_43070);
nor U45535 (N_45535,N_40000,N_44002);
nor U45536 (N_45536,N_40908,N_40140);
nor U45537 (N_45537,N_44155,N_42477);
nor U45538 (N_45538,N_41055,N_41011);
xnor U45539 (N_45539,N_44648,N_42815);
nand U45540 (N_45540,N_42507,N_44020);
nor U45541 (N_45541,N_43184,N_43047);
nor U45542 (N_45542,N_42515,N_42073);
or U45543 (N_45543,N_43522,N_41255);
xnor U45544 (N_45544,N_43116,N_43459);
and U45545 (N_45545,N_43101,N_42279);
nor U45546 (N_45546,N_41107,N_43455);
and U45547 (N_45547,N_42541,N_43607);
or U45548 (N_45548,N_44690,N_43944);
and U45549 (N_45549,N_43773,N_43044);
and U45550 (N_45550,N_44951,N_44224);
or U45551 (N_45551,N_43661,N_41506);
nor U45552 (N_45552,N_42902,N_40850);
and U45553 (N_45553,N_40408,N_40980);
and U45554 (N_45554,N_43389,N_42925);
nand U45555 (N_45555,N_42260,N_41601);
xor U45556 (N_45556,N_44235,N_41887);
and U45557 (N_45557,N_42552,N_40530);
nand U45558 (N_45558,N_41999,N_43519);
nand U45559 (N_45559,N_43013,N_41767);
nand U45560 (N_45560,N_41979,N_44578);
or U45561 (N_45561,N_40376,N_40497);
nand U45562 (N_45562,N_41094,N_44443);
xor U45563 (N_45563,N_43632,N_41945);
xnor U45564 (N_45564,N_44545,N_44404);
and U45565 (N_45565,N_40438,N_40732);
and U45566 (N_45566,N_44823,N_44131);
or U45567 (N_45567,N_43391,N_44399);
or U45568 (N_45568,N_41508,N_40534);
nor U45569 (N_45569,N_41235,N_41010);
nor U45570 (N_45570,N_44013,N_40869);
and U45571 (N_45571,N_44573,N_44549);
or U45572 (N_45572,N_41893,N_41452);
and U45573 (N_45573,N_42699,N_44608);
and U45574 (N_45574,N_44862,N_41846);
or U45575 (N_45575,N_40894,N_41080);
nand U45576 (N_45576,N_41972,N_44924);
nor U45577 (N_45577,N_42314,N_41376);
and U45578 (N_45578,N_41834,N_41682);
nand U45579 (N_45579,N_41941,N_43614);
nand U45580 (N_45580,N_41571,N_42095);
nor U45581 (N_45581,N_44676,N_43693);
nand U45582 (N_45582,N_44362,N_43126);
and U45583 (N_45583,N_40406,N_40429);
nor U45584 (N_45584,N_44405,N_44295);
nand U45585 (N_45585,N_43498,N_42578);
nor U45586 (N_45586,N_40287,N_40068);
or U45587 (N_45587,N_43752,N_43664);
xnor U45588 (N_45588,N_40190,N_43287);
nor U45589 (N_45589,N_41917,N_40305);
and U45590 (N_45590,N_44706,N_42675);
or U45591 (N_45591,N_40755,N_40528);
nor U45592 (N_45592,N_40699,N_42656);
nand U45593 (N_45593,N_43398,N_43729);
nand U45594 (N_45594,N_41568,N_44278);
nand U45595 (N_45595,N_42085,N_44333);
or U45596 (N_45596,N_42827,N_40200);
and U45597 (N_45597,N_40713,N_41768);
or U45598 (N_45598,N_42717,N_40815);
or U45599 (N_45599,N_41325,N_43030);
nand U45600 (N_45600,N_40823,N_40752);
and U45601 (N_45601,N_43948,N_44498);
or U45602 (N_45602,N_41930,N_43085);
or U45603 (N_45603,N_42732,N_44484);
or U45604 (N_45604,N_41792,N_41106);
nor U45605 (N_45605,N_43840,N_42099);
nor U45606 (N_45606,N_44271,N_43068);
xor U45607 (N_45607,N_42814,N_44263);
nor U45608 (N_45608,N_44929,N_41294);
nor U45609 (N_45609,N_43949,N_40981);
or U45610 (N_45610,N_44368,N_42105);
and U45611 (N_45611,N_43883,N_44139);
or U45612 (N_45612,N_41769,N_41445);
nor U45613 (N_45613,N_40805,N_44411);
nor U45614 (N_45614,N_44284,N_44763);
xor U45615 (N_45615,N_43550,N_42729);
nor U45616 (N_45616,N_44880,N_40309);
and U45617 (N_45617,N_44957,N_42770);
nand U45618 (N_45618,N_42231,N_40435);
or U45619 (N_45619,N_40871,N_41839);
nor U45620 (N_45620,N_40969,N_42132);
or U45621 (N_45621,N_42555,N_41676);
and U45622 (N_45622,N_40436,N_40251);
and U45623 (N_45623,N_42156,N_44535);
nand U45624 (N_45624,N_43463,N_43981);
or U45625 (N_45625,N_43903,N_42480);
nor U45626 (N_45626,N_42470,N_44074);
nand U45627 (N_45627,N_40995,N_43708);
and U45628 (N_45628,N_40986,N_41690);
nor U45629 (N_45629,N_42086,N_40248);
nor U45630 (N_45630,N_43541,N_43299);
and U45631 (N_45631,N_43382,N_42235);
xor U45632 (N_45632,N_44210,N_41368);
nand U45633 (N_45633,N_40152,N_41546);
and U45634 (N_45634,N_41168,N_43302);
nor U45635 (N_45635,N_44559,N_40724);
nand U45636 (N_45636,N_44054,N_41266);
nor U45637 (N_45637,N_43701,N_40101);
nand U45638 (N_45638,N_41065,N_40070);
or U45639 (N_45639,N_41875,N_42571);
or U45640 (N_45640,N_44658,N_40648);
nand U45641 (N_45641,N_43569,N_42168);
nand U45642 (N_45642,N_44642,N_40378);
xor U45643 (N_45643,N_43891,N_40002);
and U45644 (N_45644,N_40212,N_40025);
or U45645 (N_45645,N_42796,N_42259);
and U45646 (N_45646,N_41822,N_44677);
nor U45647 (N_45647,N_42106,N_44943);
and U45648 (N_45648,N_41401,N_44166);
nor U45649 (N_45649,N_44521,N_40966);
nand U45650 (N_45650,N_44331,N_41242);
or U45651 (N_45651,N_44711,N_40720);
and U45652 (N_45652,N_43380,N_41103);
nor U45653 (N_45653,N_44207,N_42076);
nor U45654 (N_45654,N_40469,N_42999);
and U45655 (N_45655,N_44799,N_43760);
nor U45656 (N_45656,N_40537,N_44905);
and U45657 (N_45657,N_43023,N_41816);
nand U45658 (N_45658,N_44248,N_43000);
nand U45659 (N_45659,N_43354,N_41134);
nor U45660 (N_45660,N_44516,N_44602);
xor U45661 (N_45661,N_40263,N_40719);
and U45662 (N_45662,N_43634,N_41900);
nand U45663 (N_45663,N_42859,N_42579);
nor U45664 (N_45664,N_41819,N_42774);
and U45665 (N_45665,N_44981,N_40456);
and U45666 (N_45666,N_43874,N_42393);
and U45667 (N_45667,N_43311,N_44640);
nand U45668 (N_45668,N_40291,N_41791);
and U45669 (N_45669,N_43483,N_44663);
or U45670 (N_45670,N_41393,N_42325);
xnor U45671 (N_45671,N_44564,N_42929);
xnor U45672 (N_45672,N_44300,N_41146);
and U45673 (N_45673,N_42843,N_43782);
or U45674 (N_45674,N_44788,N_40728);
and U45675 (N_45675,N_44221,N_41084);
nor U45676 (N_45676,N_40709,N_41458);
and U45677 (N_45677,N_41511,N_40367);
xor U45678 (N_45678,N_41175,N_43543);
and U45679 (N_45679,N_44934,N_43404);
or U45680 (N_45680,N_42688,N_41281);
or U45681 (N_45681,N_42799,N_44432);
and U45682 (N_45682,N_42961,N_40631);
nor U45683 (N_45683,N_44645,N_40400);
or U45684 (N_45684,N_42306,N_43645);
and U45685 (N_45685,N_43524,N_44520);
nand U45686 (N_45686,N_43215,N_42358);
or U45687 (N_45687,N_44673,N_44758);
nand U45688 (N_45688,N_41225,N_44488);
and U45689 (N_45689,N_44912,N_44820);
and U45690 (N_45690,N_41710,N_40244);
xnor U45691 (N_45691,N_43998,N_40372);
and U45692 (N_45692,N_42102,N_42431);
nor U45693 (N_45693,N_41163,N_40443);
and U45694 (N_45694,N_44713,N_40503);
nor U45695 (N_45695,N_41284,N_44875);
nand U45696 (N_45696,N_42559,N_42658);
or U45697 (N_45697,N_42730,N_44748);
xor U45698 (N_45698,N_42682,N_43657);
nand U45699 (N_45699,N_44148,N_41686);
nand U45700 (N_45700,N_44006,N_40867);
nand U45701 (N_45701,N_40794,N_42191);
and U45702 (N_45702,N_41931,N_40320);
and U45703 (N_45703,N_42445,N_42968);
and U45704 (N_45704,N_41628,N_44312);
nor U45705 (N_45705,N_42905,N_42243);
nand U45706 (N_45706,N_40459,N_43229);
and U45707 (N_45707,N_44491,N_43158);
nand U45708 (N_45708,N_41399,N_44282);
and U45709 (N_45709,N_41343,N_41633);
and U45710 (N_45710,N_44344,N_43532);
and U45711 (N_45711,N_40820,N_41976);
nor U45712 (N_45712,N_43441,N_44019);
nor U45713 (N_45713,N_44065,N_44309);
xor U45714 (N_45714,N_44379,N_44766);
and U45715 (N_45715,N_44811,N_41553);
nor U45716 (N_45716,N_42349,N_41429);
nand U45717 (N_45717,N_41319,N_42230);
or U45718 (N_45718,N_41920,N_40682);
xnor U45719 (N_45719,N_41386,N_43856);
nand U45720 (N_45720,N_44007,N_43506);
or U45721 (N_45721,N_44661,N_41205);
or U45722 (N_45722,N_43736,N_43746);
nor U45723 (N_45723,N_40627,N_41515);
or U45724 (N_45724,N_40434,N_42878);
xnor U45725 (N_45725,N_42857,N_41520);
and U45726 (N_45726,N_42830,N_41997);
or U45727 (N_45727,N_43595,N_42897);
xnor U45728 (N_45728,N_40004,N_41512);
and U45729 (N_45729,N_43197,N_44004);
and U45730 (N_45730,N_43978,N_44562);
xor U45731 (N_45731,N_41479,N_44639);
xor U45732 (N_45732,N_41229,N_40472);
nand U45733 (N_45733,N_41124,N_41463);
nand U45734 (N_45734,N_42526,N_40661);
nand U45735 (N_45735,N_44260,N_42821);
and U45736 (N_45736,N_40083,N_44638);
nand U45737 (N_45737,N_44694,N_43628);
nor U45738 (N_45738,N_41809,N_44930);
nor U45739 (N_45739,N_44084,N_41709);
nand U45740 (N_45740,N_41480,N_40334);
nand U45741 (N_45741,N_43515,N_43618);
or U45742 (N_45742,N_40983,N_40971);
nand U45743 (N_45743,N_41442,N_41529);
xor U45744 (N_45744,N_42807,N_40415);
nor U45745 (N_45745,N_40526,N_44551);
nor U45746 (N_45746,N_43652,N_43165);
or U45747 (N_45747,N_43478,N_41585);
and U45748 (N_45748,N_41028,N_41943);
nor U45749 (N_45749,N_44393,N_40705);
or U45750 (N_45750,N_43057,N_43899);
and U45751 (N_45751,N_43548,N_40138);
nor U45752 (N_45752,N_44285,N_42319);
or U45753 (N_45753,N_44023,N_40319);
xnor U45754 (N_45754,N_44119,N_42568);
and U45755 (N_45755,N_44087,N_41327);
or U45756 (N_45756,N_44137,N_43739);
nor U45757 (N_45757,N_44228,N_40160);
and U45758 (N_45758,N_44770,N_42942);
and U45759 (N_45759,N_43426,N_41811);
and U45760 (N_45760,N_43114,N_42518);
or U45761 (N_45761,N_44908,N_41118);
or U45762 (N_45762,N_44297,N_42473);
nor U45763 (N_45763,N_42438,N_44283);
xnor U45764 (N_45764,N_41878,N_42785);
or U45765 (N_45765,N_42622,N_44112);
nand U45766 (N_45766,N_41484,N_44980);
and U45767 (N_45767,N_44719,N_40622);
nand U45768 (N_45768,N_42825,N_41730);
and U45769 (N_45769,N_43710,N_40129);
and U45770 (N_45770,N_43032,N_42199);
or U45771 (N_45771,N_41639,N_42700);
nor U45772 (N_45772,N_41663,N_40045);
nand U45773 (N_45773,N_42385,N_40316);
nor U45774 (N_45774,N_41855,N_41108);
and U45775 (N_45775,N_40677,N_42511);
or U45776 (N_45776,N_42178,N_42998);
nor U45777 (N_45777,N_42446,N_43784);
and U45778 (N_45778,N_43533,N_42372);
and U45779 (N_45779,N_41085,N_40397);
or U45780 (N_45780,N_43968,N_44522);
xnor U45781 (N_45781,N_43276,N_43936);
nor U45782 (N_45782,N_42338,N_41944);
nor U45783 (N_45783,N_40462,N_40959);
nand U45784 (N_45784,N_44597,N_43642);
nand U45785 (N_45785,N_43866,N_41510);
or U45786 (N_45786,N_42776,N_42544);
xnor U45787 (N_45787,N_42276,N_43046);
or U45788 (N_45788,N_42640,N_42309);
or U45789 (N_45789,N_44587,N_41260);
or U45790 (N_45790,N_42001,N_42378);
and U45791 (N_45791,N_41561,N_41863);
and U45792 (N_45792,N_41574,N_40930);
nand U45793 (N_45793,N_41692,N_41402);
or U45794 (N_45794,N_41300,N_40207);
nor U45795 (N_45795,N_44835,N_44798);
or U45796 (N_45796,N_42727,N_41210);
and U45797 (N_45797,N_44860,N_40898);
and U45798 (N_45798,N_42840,N_44086);
nor U45799 (N_45799,N_43762,N_40624);
and U45800 (N_45800,N_44856,N_41820);
and U45801 (N_45801,N_42997,N_43635);
and U45802 (N_45802,N_40026,N_43650);
and U45803 (N_45803,N_43337,N_41385);
or U45804 (N_45804,N_41487,N_42381);
or U45805 (N_45805,N_44192,N_40556);
xor U45806 (N_45806,N_40853,N_42311);
or U45807 (N_45807,N_40653,N_41715);
nand U45808 (N_45808,N_43056,N_41007);
or U45809 (N_45809,N_42749,N_42092);
or U45810 (N_45810,N_40323,N_41164);
or U45811 (N_45811,N_44851,N_43198);
nor U45812 (N_45812,N_41980,N_42454);
and U45813 (N_45813,N_40906,N_44774);
nand U45814 (N_45814,N_44438,N_40846);
or U45815 (N_45815,N_42236,N_42934);
xnor U45816 (N_45816,N_42205,N_40707);
nor U45817 (N_45817,N_43160,N_44796);
nand U45818 (N_45818,N_44591,N_41722);
nand U45819 (N_45819,N_42224,N_41762);
or U45820 (N_45820,N_40476,N_43625);
nor U45821 (N_45821,N_42940,N_42232);
or U45822 (N_45822,N_43735,N_41160);
or U45823 (N_45823,N_40077,N_44683);
or U45824 (N_45824,N_41670,N_42033);
nand U45825 (N_45825,N_41962,N_43143);
nand U45826 (N_45826,N_41060,N_42666);
nand U45827 (N_45827,N_42078,N_43178);
or U45828 (N_45828,N_41807,N_42342);
and U45829 (N_45829,N_44958,N_40687);
and U45830 (N_45830,N_40936,N_42340);
and U45831 (N_45831,N_44146,N_40970);
nor U45832 (N_45832,N_43723,N_42391);
nor U45833 (N_45833,N_44775,N_41388);
or U45834 (N_45834,N_41968,N_42432);
nand U45835 (N_45835,N_43830,N_44941);
nor U45836 (N_45836,N_40229,N_41925);
or U45837 (N_45837,N_43490,N_42047);
or U45838 (N_45838,N_43432,N_40803);
and U45839 (N_45839,N_43248,N_44672);
and U45840 (N_45840,N_43989,N_42058);
and U45841 (N_45841,N_42398,N_40782);
or U45842 (N_45842,N_41110,N_40877);
nand U45843 (N_45843,N_43395,N_40137);
nor U45844 (N_45844,N_44339,N_41328);
and U45845 (N_45845,N_42847,N_40383);
and U45846 (N_45846,N_41831,N_44736);
nand U45847 (N_45847,N_43539,N_43716);
nor U45848 (N_45848,N_41851,N_40131);
nand U45849 (N_45849,N_41509,N_42575);
nand U45850 (N_45850,N_42271,N_44454);
and U45851 (N_45851,N_40418,N_41191);
nand U45852 (N_45852,N_43252,N_41748);
or U45853 (N_45853,N_40968,N_44707);
nand U45854 (N_45854,N_42007,N_44920);
nand U45855 (N_45855,N_42927,N_44776);
or U45856 (N_45856,N_41157,N_40856);
or U45857 (N_45857,N_40571,N_43155);
or U45858 (N_45858,N_41698,N_44268);
or U45859 (N_45859,N_44813,N_43141);
nand U45860 (N_45860,N_40925,N_41695);
or U45861 (N_45861,N_43104,N_42935);
and U45862 (N_45862,N_43826,N_40962);
nand U45863 (N_45863,N_43888,N_43307);
and U45864 (N_45864,N_41499,N_43341);
or U45865 (N_45865,N_42710,N_42803);
or U45866 (N_45866,N_44030,N_43356);
nand U45867 (N_45867,N_41912,N_42439);
or U45868 (N_45868,N_44894,N_43925);
nand U45869 (N_45869,N_41081,N_42502);
and U45870 (N_45870,N_40819,N_44206);
or U45871 (N_45871,N_43914,N_44469);
nor U45872 (N_45872,N_40636,N_40826);
nand U45873 (N_45873,N_42708,N_43181);
nand U45874 (N_45874,N_40060,N_44211);
or U45875 (N_45875,N_43917,N_40646);
or U45876 (N_45876,N_44436,N_43631);
nand U45877 (N_45877,N_44961,N_42134);
xor U45878 (N_45878,N_40895,N_41869);
or U45879 (N_45879,N_44069,N_40133);
or U45880 (N_45880,N_42554,N_44605);
nand U45881 (N_45881,N_41647,N_42149);
or U45882 (N_45882,N_40067,N_40454);
and U45883 (N_45883,N_40321,N_40113);
or U45884 (N_45884,N_40041,N_43605);
and U45885 (N_45885,N_44652,N_42412);
or U45886 (N_45886,N_43554,N_42560);
xnor U45887 (N_45887,N_41223,N_40975);
nor U45888 (N_45888,N_44056,N_41354);
or U45889 (N_45889,N_42912,N_43214);
xnor U45890 (N_45890,N_44703,N_40273);
xnor U45891 (N_45891,N_44225,N_41476);
nor U45892 (N_45892,N_43037,N_40642);
and U45893 (N_45893,N_40885,N_42103);
or U45894 (N_45894,N_42679,N_42211);
xor U45895 (N_45895,N_41470,N_44708);
or U45896 (N_45896,N_42414,N_43829);
nor U45897 (N_45897,N_42123,N_41317);
nand U45898 (N_45898,N_43869,N_43019);
and U45899 (N_45899,N_40912,N_42716);
or U45900 (N_45900,N_40665,N_44060);
or U45901 (N_45901,N_44066,N_40864);
nor U45902 (N_45902,N_40916,N_44439);
nor U45903 (N_45903,N_42551,N_42075);
nor U45904 (N_45904,N_41464,N_43015);
and U45905 (N_45905,N_42482,N_40601);
or U45906 (N_45906,N_41631,N_43613);
xor U45907 (N_45907,N_40878,N_42538);
or U45908 (N_45908,N_41501,N_40950);
nor U45909 (N_45909,N_44772,N_43956);
nand U45910 (N_45910,N_44525,N_43979);
and U45911 (N_45911,N_41344,N_42849);
and U45912 (N_45912,N_41714,N_44883);
or U45913 (N_45913,N_40243,N_40748);
or U45914 (N_45914,N_43789,N_41759);
xnor U45915 (N_45915,N_42589,N_44710);
nor U45916 (N_45916,N_42914,N_40920);
and U45917 (N_45917,N_40439,N_40787);
nand U45918 (N_45918,N_43887,N_44721);
xnor U45919 (N_45919,N_43749,N_42247);
nor U45920 (N_45920,N_42180,N_42946);
and U45921 (N_45921,N_44699,N_40522);
xor U45922 (N_45922,N_43419,N_43875);
xor U45923 (N_45923,N_40351,N_40195);
xor U45924 (N_45924,N_40156,N_44276);
nor U45925 (N_45925,N_43272,N_43806);
nor U45926 (N_45926,N_43081,N_44430);
or U45927 (N_45927,N_44009,N_41451);
nor U45928 (N_45928,N_41953,N_41653);
nand U45929 (N_45929,N_44049,N_40022);
and U45930 (N_45930,N_44687,N_42365);
and U45931 (N_45931,N_43637,N_42209);
or U45932 (N_45932,N_41882,N_43318);
nand U45933 (N_45933,N_43294,N_44416);
nand U45934 (N_45934,N_42738,N_41366);
nand U45935 (N_45935,N_42031,N_42855);
nor U45936 (N_45936,N_43927,N_40250);
nand U45937 (N_45937,N_44999,N_44604);
nand U45938 (N_45938,N_44768,N_40410);
xnor U45939 (N_45939,N_42488,N_43183);
or U45940 (N_45940,N_42969,N_42302);
and U45941 (N_45941,N_42596,N_44033);
nand U45942 (N_45942,N_40270,N_44709);
and U45943 (N_45943,N_44318,N_41035);
xor U45944 (N_45944,N_43526,N_43537);
nand U45945 (N_45945,N_41226,N_44975);
and U45946 (N_45946,N_40062,N_42322);
xnor U45947 (N_45947,N_43421,N_40345);
and U45948 (N_45948,N_41929,N_42848);
nand U45949 (N_45949,N_43268,N_42335);
or U45950 (N_45950,N_40249,N_42655);
nor U45951 (N_45951,N_43612,N_44504);
nand U45952 (N_45952,N_40496,N_40071);
xor U45953 (N_45953,N_40741,N_42304);
nor U45954 (N_45954,N_42936,N_44907);
or U45955 (N_45955,N_40518,N_40967);
or U45956 (N_45956,N_42355,N_42072);
or U45957 (N_45957,N_42725,N_41174);
nor U45958 (N_45958,N_44063,N_43945);
or U45959 (N_45959,N_42698,N_42097);
nor U45960 (N_45960,N_43834,N_43761);
xor U45961 (N_45961,N_44018,N_41161);
xnor U45962 (N_45962,N_42013,N_40187);
xor U45963 (N_45963,N_43142,N_40440);
nor U45964 (N_45964,N_44756,N_43467);
and U45965 (N_45965,N_40460,N_42461);
or U45966 (N_45966,N_44444,N_42775);
nand U45967 (N_45967,N_44094,N_41859);
nand U45968 (N_45968,N_44659,N_40354);
and U45969 (N_45969,N_41481,N_44200);
and U45970 (N_45970,N_43263,N_44816);
nand U45971 (N_45971,N_42429,N_42791);
nor U45972 (N_45972,N_43373,N_40283);
or U45973 (N_45973,N_40681,N_43793);
nor U45974 (N_45974,N_42573,N_42227);
xor U45975 (N_45975,N_44947,N_44322);
nor U45976 (N_45976,N_40839,N_40639);
nor U45977 (N_45977,N_43902,N_40550);
nor U45978 (N_45978,N_42217,N_42018);
and U45979 (N_45979,N_43727,N_44542);
nand U45980 (N_45980,N_41145,N_40151);
xnor U45981 (N_45981,N_43447,N_40108);
and U45982 (N_45982,N_42587,N_41289);
and U45983 (N_45983,N_41155,N_42919);
nor U45984 (N_45984,N_40931,N_42176);
xnor U45985 (N_45985,N_42242,N_41993);
and U45986 (N_45986,N_44461,N_41877);
and U45987 (N_45987,N_40485,N_44279);
or U45988 (N_45988,N_40897,N_40252);
or U45989 (N_45989,N_41804,N_44839);
or U45990 (N_45990,N_44177,N_44682);
nand U45991 (N_45991,N_42496,N_40030);
and U45992 (N_45992,N_44090,N_42324);
nand U45993 (N_45993,N_40385,N_41914);
nor U45994 (N_45994,N_43292,N_41894);
or U45995 (N_45995,N_41873,N_41777);
or U45996 (N_45996,N_40922,N_43180);
and U45997 (N_45997,N_42455,N_44779);
nor U45998 (N_45998,N_44857,N_43939);
xnor U45999 (N_45999,N_43685,N_41190);
nor U46000 (N_46000,N_44377,N_42297);
and U46001 (N_46001,N_43988,N_44161);
nor U46002 (N_46002,N_44741,N_40050);
nand U46003 (N_46003,N_43558,N_41206);
or U46004 (N_46004,N_40606,N_44616);
nor U46005 (N_46005,N_43780,N_41288);
and U46006 (N_46006,N_44116,N_44940);
or U46007 (N_46007,N_43599,N_40226);
and U46008 (N_46008,N_42332,N_43358);
nand U46009 (N_46009,N_43050,N_43079);
and U46010 (N_46010,N_43689,N_40865);
nor U46011 (N_46011,N_42421,N_41626);
nand U46012 (N_46012,N_44219,N_42906);
nor U46013 (N_46013,N_41340,N_43572);
nor U46014 (N_46014,N_43074,N_44035);
nand U46015 (N_46015,N_43765,N_41689);
nand U46016 (N_46016,N_42955,N_40048);
or U46017 (N_46017,N_41301,N_41883);
or U46018 (N_46018,N_44979,N_44547);
and U46019 (N_46019,N_44419,N_43758);
and U46020 (N_46020,N_41954,N_41713);
and U46021 (N_46021,N_42686,N_43703);
or U46022 (N_46022,N_42039,N_42886);
and U46023 (N_46023,N_41156,N_40758);
or U46024 (N_46024,N_44108,N_44678);
and U46025 (N_46025,N_41029,N_44695);
and U46026 (N_46026,N_44369,N_44617);
nand U46027 (N_46027,N_41897,N_40811);
or U46028 (N_46028,N_42165,N_43658);
nor U46029 (N_46029,N_40994,N_42657);
or U46030 (N_46030,N_41197,N_44140);
nor U46031 (N_46031,N_44952,N_41646);
xor U46032 (N_46032,N_41844,N_42661);
nand U46033 (N_46033,N_43065,N_42842);
or U46034 (N_46034,N_40668,N_40092);
or U46035 (N_46035,N_43651,N_44456);
nor U46036 (N_46036,N_43960,N_42882);
nand U46037 (N_46037,N_43656,N_43377);
and U46038 (N_46038,N_44600,N_42440);
nand U46039 (N_46039,N_44320,N_43720);
or U46040 (N_46040,N_43694,N_40123);
xor U46041 (N_46041,N_41850,N_42627);
nor U46042 (N_46042,N_41838,N_42510);
nand U46043 (N_46043,N_42692,N_44301);
and U46044 (N_46044,N_42947,N_40584);
xor U46045 (N_46045,N_43138,N_42788);
nor U46046 (N_46046,N_41668,N_42852);
nor U46047 (N_46047,N_41910,N_44420);
nor U46048 (N_46048,N_40891,N_41212);
and U46049 (N_46049,N_43534,N_41473);
nor U46050 (N_46050,N_42967,N_43051);
nor U46051 (N_46051,N_43069,N_42504);
nand U46052 (N_46052,N_41074,N_42574);
nand U46053 (N_46053,N_40218,N_44515);
nor U46054 (N_46054,N_44252,N_40054);
nor U46055 (N_46055,N_40216,N_43926);
nor U46056 (N_46056,N_41612,N_42060);
or U46057 (N_46057,N_41194,N_42202);
nor U46058 (N_46058,N_40340,N_44556);
and U46059 (N_46059,N_40704,N_42797);
nor U46060 (N_46060,N_43413,N_43861);
nor U46061 (N_46061,N_41020,N_43489);
or U46062 (N_46062,N_42653,N_41261);
and U46063 (N_46063,N_43832,N_40607);
or U46064 (N_46064,N_41287,N_43094);
nor U46065 (N_46065,N_42907,N_40204);
and U46066 (N_46066,N_41876,N_44577);
nand U46067 (N_46067,N_40392,N_44938);
and U46068 (N_46068,N_42713,N_43864);
xnor U46069 (N_46069,N_41557,N_42980);
nor U46070 (N_46070,N_42739,N_40525);
nor U46071 (N_46071,N_40085,N_44946);
and U46072 (N_46072,N_44812,N_40311);
xnor U46073 (N_46073,N_41111,N_43117);
nand U46074 (N_46074,N_40744,N_42089);
nor U46075 (N_46075,N_40746,N_41440);
nand U46076 (N_46076,N_40535,N_44198);
and U46077 (N_46077,N_42246,N_40965);
or U46078 (N_46078,N_43860,N_44988);
and U46079 (N_46079,N_40269,N_44829);
nand U46080 (N_46080,N_43201,N_40910);
xor U46081 (N_46081,N_41555,N_43469);
or U46082 (N_46082,N_43314,N_42888);
nand U46083 (N_46083,N_40344,N_40300);
nand U46084 (N_46084,N_40848,N_41867);
or U46085 (N_46085,N_40358,N_40159);
or U46086 (N_46086,N_42883,N_41497);
and U46087 (N_46087,N_41040,N_41378);
and U46088 (N_46088,N_44746,N_44394);
nand U46089 (N_46089,N_41390,N_42257);
xor U46090 (N_46090,N_43799,N_43482);
and U46091 (N_46091,N_41806,N_43707);
or U46092 (N_46092,N_44782,N_43620);
nand U46093 (N_46093,N_43424,N_43923);
or U46094 (N_46094,N_44303,N_44727);
or U46095 (N_46095,N_44068,N_44671);
nand U46096 (N_46096,N_43951,N_40003);
and U46097 (N_46097,N_44334,N_42447);
xor U46098 (N_46098,N_43687,N_41104);
nor U46099 (N_46099,N_43091,N_43136);
or U46100 (N_46100,N_40698,N_43911);
xor U46101 (N_46101,N_44844,N_43111);
nor U46102 (N_46102,N_40688,N_43422);
nor U46103 (N_46103,N_40088,N_43638);
nand U46104 (N_46104,N_41841,N_41105);
and U46105 (N_46105,N_41678,N_43473);
nor U46106 (N_46106,N_42333,N_41427);
nand U46107 (N_46107,N_41996,N_41625);
and U46108 (N_46108,N_40304,N_41416);
nand U46109 (N_46109,N_41180,N_41620);
xnor U46110 (N_46110,N_43228,N_40893);
xor U46111 (N_46111,N_43523,N_42783);
nor U46112 (N_46112,N_43270,N_44609);
nor U46113 (N_46113,N_41150,N_44176);
and U46114 (N_46114,N_40370,N_40326);
nand U46115 (N_46115,N_43087,N_43425);
nor U46116 (N_46116,N_42366,N_44417);
nor U46117 (N_46117,N_41251,N_44662);
or U46118 (N_46118,N_43468,N_43867);
nor U46119 (N_46119,N_44917,N_44655);
or U46120 (N_46120,N_43179,N_43220);
or U46121 (N_46121,N_43431,N_41935);
nor U46122 (N_46122,N_43360,N_40608);
nand U46123 (N_46123,N_40055,N_42530);
nand U46124 (N_46124,N_40552,N_41864);
nor U46125 (N_46125,N_40333,N_44383);
nand U46126 (N_46126,N_40444,N_43681);
xor U46127 (N_46127,N_41355,N_43012);
nand U46128 (N_46128,N_43194,N_40818);
nor U46129 (N_46129,N_43428,N_43265);
or U46130 (N_46130,N_44532,N_44595);
nor U46131 (N_46131,N_40130,N_44501);
and U46132 (N_46132,N_44003,N_42633);
or U46133 (N_46133,N_40422,N_40258);
nand U46134 (N_46134,N_42344,N_43045);
nor U46135 (N_46135,N_41640,N_42328);
nor U46136 (N_46136,N_41472,N_43863);
or U46137 (N_46137,N_43344,N_41254);
and U46138 (N_46138,N_40582,N_41974);
nand U46139 (N_46139,N_43805,N_43492);
and U46140 (N_46140,N_44954,N_42188);
nor U46141 (N_46141,N_44126,N_40016);
nand U46142 (N_46142,N_40102,N_43261);
or U46143 (N_46143,N_41151,N_41259);
and U46144 (N_46144,N_41998,N_41536);
and U46145 (N_46145,N_43975,N_44038);
nand U46146 (N_46146,N_44925,N_43401);
nand U46147 (N_46147,N_42972,N_43576);
nand U46148 (N_46148,N_42876,N_44530);
or U46149 (N_46149,N_41872,N_41236);
nor U46150 (N_46150,N_43677,N_44226);
nand U46151 (N_46151,N_43203,N_40557);
and U46152 (N_46152,N_41538,N_44114);
or U46153 (N_46153,N_43297,N_40985);
xor U46154 (N_46154,N_43546,N_42893);
and U46155 (N_46155,N_43502,N_40779);
and U46156 (N_46156,N_40416,N_41507);
or U46157 (N_46157,N_43123,N_42065);
nor U46158 (N_46158,N_43006,N_40289);
nor U46159 (N_46159,N_44495,N_44277);
or U46160 (N_46160,N_41000,N_42044);
or U46161 (N_46161,N_40672,N_43017);
nand U46162 (N_46162,N_42664,N_43115);
nor U46163 (N_46163,N_41290,N_44472);
nand U46164 (N_46164,N_40176,N_42605);
or U46165 (N_46165,N_44715,N_42539);
or U46166 (N_46166,N_41444,N_44619);
nand U46167 (N_46167,N_40957,N_43909);
nor U46168 (N_46168,N_42436,N_42760);
and U46169 (N_46169,N_42801,N_44264);
and U46170 (N_46170,N_43994,N_41919);
or U46171 (N_46171,N_43313,N_43402);
or U46172 (N_46172,N_42828,N_44246);
and U46173 (N_46173,N_43334,N_41449);
and U46174 (N_46174,N_42728,N_40812);
nand U46175 (N_46175,N_40449,N_41149);
or U46176 (N_46176,N_43997,N_40964);
nor U46177 (N_46177,N_42667,N_44187);
nand U46178 (N_46178,N_40745,N_40228);
and U46179 (N_46179,N_41373,N_42819);
or U46180 (N_46180,N_41283,N_42762);
nor U46181 (N_46181,N_43118,N_42360);
nand U46182 (N_46182,N_41805,N_43147);
or U46183 (N_46183,N_44304,N_43191);
nor U46184 (N_46184,N_42169,N_44702);
and U46185 (N_46185,N_44754,N_41828);
nor U46186 (N_46186,N_43654,N_44933);
and U46187 (N_46187,N_44863,N_44143);
nand U46188 (N_46188,N_44801,N_40089);
or U46189 (N_46189,N_41790,N_42813);
nor U46190 (N_46190,N_41116,N_42023);
or U46191 (N_46191,N_40998,N_42614);
or U46192 (N_46192,N_42836,N_43884);
and U46193 (N_46193,N_40809,N_43872);
nand U46194 (N_46194,N_43896,N_42812);
or U46195 (N_46195,N_43415,N_43052);
nor U46196 (N_46196,N_44893,N_41039);
nand U46197 (N_46197,N_42778,N_40230);
or U46198 (N_46198,N_42359,N_41729);
nor U46199 (N_46199,N_41372,N_40610);
or U46200 (N_46200,N_43148,N_41304);
xor U46201 (N_46201,N_40549,N_40100);
nor U46202 (N_46202,N_42874,N_44631);
xnor U46203 (N_46203,N_43105,N_43024);
and U46204 (N_46204,N_41772,N_40847);
and U46205 (N_46205,N_42239,N_40675);
nand U46206 (N_46206,N_42565,N_41952);
nor U46207 (N_46207,N_41066,N_42400);
and U46208 (N_46208,N_41234,N_42434);
nand U46209 (N_46209,N_43103,N_42061);
or U46210 (N_46210,N_42256,N_42546);
nor U46211 (N_46211,N_44641,N_43757);
and U46212 (N_46212,N_42681,N_42141);
or U46213 (N_46213,N_44475,N_41089);
or U46214 (N_46214,N_43175,N_44544);
and U46215 (N_46215,N_43135,N_43173);
nor U46216 (N_46216,N_41265,N_42743);
and U46217 (N_46217,N_44024,N_43185);
and U46218 (N_46218,N_43223,N_41456);
and U46219 (N_46219,N_41738,N_44769);
nand U46220 (N_46220,N_42222,N_44195);
and U46221 (N_46221,N_41358,N_44674);
nor U46222 (N_46222,N_43098,N_40038);
nand U46223 (N_46223,N_40122,N_41455);
and U46224 (N_46224,N_42780,N_42600);
nor U46225 (N_46225,N_42789,N_42345);
nand U46226 (N_46226,N_42736,N_41796);
nand U46227 (N_46227,N_40927,N_41032);
nor U46228 (N_46228,N_40134,N_44186);
xor U46229 (N_46229,N_40954,N_41188);
nor U46230 (N_46230,N_42040,N_43930);
nand U46231 (N_46231,N_41679,N_43690);
and U46232 (N_46232,N_44253,N_41582);
nor U46233 (N_46233,N_40006,N_41187);
nand U46234 (N_46234,N_41403,N_44476);
and U46235 (N_46235,N_42261,N_41837);
nand U46236 (N_46236,N_40282,N_42534);
nand U46237 (N_46237,N_41418,N_42957);
nand U46238 (N_46238,N_43403,N_44082);
xor U46239 (N_46239,N_43584,N_42002);
and U46240 (N_46240,N_43504,N_43499);
nand U46241 (N_46241,N_42337,N_43794);
nor U46242 (N_46242,N_41367,N_43849);
and U46243 (N_46243,N_44395,N_41928);
or U46244 (N_46244,N_40946,N_43843);
nor U46245 (N_46245,N_41588,N_43327);
and U46246 (N_46246,N_44272,N_41789);
xor U46247 (N_46247,N_42542,N_43906);
nor U46248 (N_46248,N_44083,N_42941);
nand U46249 (N_46249,N_44555,N_41048);
nor U46250 (N_46250,N_43844,N_40080);
nor U46251 (N_46251,N_41751,N_40268);
and U46252 (N_46252,N_41774,N_43480);
and U46253 (N_46253,N_43336,N_42417);
nor U46254 (N_46254,N_41799,N_44243);
and U46255 (N_46255,N_42616,N_40796);
and U46256 (N_46256,N_41649,N_44104);
nand U46257 (N_46257,N_43691,N_40494);
or U46258 (N_46258,N_42896,N_41423);
and U46259 (N_46259,N_40353,N_44364);
or U46260 (N_46260,N_40632,N_43947);
nor U46261 (N_46261,N_40445,N_42879);
nand U46262 (N_46262,N_43717,N_43982);
and U46263 (N_46263,N_41829,N_41009);
or U46264 (N_46264,N_43807,N_44828);
nand U46265 (N_46265,N_41932,N_42648);
nand U46266 (N_46266,N_40332,N_43900);
nor U46267 (N_46267,N_41577,N_44895);
nor U46268 (N_46268,N_43454,N_43222);
nor U46269 (N_46269,N_43580,N_43655);
nand U46270 (N_46270,N_44785,N_42435);
or U46271 (N_46271,N_41939,N_43540);
and U46272 (N_46272,N_42286,N_43574);
xnor U46273 (N_46273,N_41836,N_41594);
nand U46274 (N_46274,N_42330,N_40939);
nor U46275 (N_46275,N_41840,N_40573);
nand U46276 (N_46276,N_41384,N_41904);
or U46277 (N_46277,N_42793,N_44637);
nand U46278 (N_46278,N_41095,N_44651);
nand U46279 (N_46279,N_41258,N_43258);
or U46280 (N_46280,N_40613,N_42112);
nor U46281 (N_46281,N_41830,N_41724);
or U46282 (N_46282,N_44800,N_40498);
nor U46283 (N_46283,N_40490,N_43405);
and U46284 (N_46284,N_41198,N_43986);
and U46285 (N_46285,N_43232,N_41541);
nand U46286 (N_46286,N_41746,N_40007);
nor U46287 (N_46287,N_40099,N_43788);
nand U46288 (N_46288,N_44807,N_40132);
or U46289 (N_46289,N_41274,N_41821);
xnor U46290 (N_46290,N_40296,N_41054);
nand U46291 (N_46291,N_44537,N_40217);
nand U46292 (N_46292,N_44950,N_42557);
nand U46293 (N_46293,N_41056,N_41833);
or U46294 (N_46294,N_40961,N_41292);
nand U46295 (N_46295,N_42057,N_42009);
and U46296 (N_46296,N_44414,N_44332);
nor U46297 (N_46297,N_40615,N_41413);
or U46298 (N_46298,N_43946,N_43231);
or U46299 (N_46299,N_44258,N_42038);
nand U46300 (N_46300,N_40027,N_44317);
nor U46301 (N_46301,N_44467,N_43195);
and U46302 (N_46302,N_43754,N_42139);
xor U46303 (N_46303,N_44327,N_44927);
and U46304 (N_46304,N_41405,N_43553);
xor U46305 (N_46305,N_41933,N_40236);
xor U46306 (N_46306,N_42298,N_44215);
nand U46307 (N_46307,N_41771,N_44873);
nor U46308 (N_46308,N_41814,N_44524);
nand U46309 (N_46309,N_44528,N_42399);
nor U46310 (N_46310,N_40042,N_42377);
or U46311 (N_46311,N_41970,N_42255);
nand U46312 (N_46312,N_42900,N_42903);
and U46313 (N_46313,N_44910,N_40468);
or U46314 (N_46314,N_41143,N_43146);
or U46315 (N_46315,N_43921,N_42148);
xnor U46316 (N_46316,N_40958,N_40237);
and U46317 (N_46317,N_43609,N_43937);
nand U46318 (N_46318,N_43970,N_40502);
nand U46319 (N_46319,N_44336,N_44465);
and U46320 (N_46320,N_42384,N_44280);
or U46321 (N_46321,N_40235,N_43827);
nand U46322 (N_46322,N_42406,N_41495);
xnor U46323 (N_46323,N_44570,N_40786);
or U46324 (N_46324,N_43815,N_44976);
nand U46325 (N_46325,N_42090,N_42926);
and U46326 (N_46326,N_41938,N_42021);
xnor U46327 (N_46327,N_40822,N_44238);
and U46328 (N_46328,N_40037,N_40996);
nand U46329 (N_46329,N_42506,N_44287);
or U46330 (N_46330,N_42748,N_44101);
nand U46331 (N_46331,N_42418,N_40375);
nand U46332 (N_46332,N_44044,N_44001);
nand U46333 (N_46333,N_41958,N_42068);
xor U46334 (N_46334,N_42119,N_44392);
nand U46335 (N_46335,N_41537,N_43953);
xor U46336 (N_46336,N_44761,N_40662);
nand U46337 (N_46337,N_44487,N_42109);
xor U46338 (N_46338,N_43958,N_40944);
nand U46339 (N_46339,N_40673,N_41426);
and U46340 (N_46340,N_44698,N_41420);
nor U46341 (N_46341,N_44911,N_41696);
xor U46342 (N_46342,N_42212,N_42458);
nor U46343 (N_46343,N_44306,N_43016);
nor U46344 (N_46344,N_42054,N_42566);
nand U46345 (N_46345,N_41711,N_40768);
and U46346 (N_46346,N_42285,N_43386);
nor U46347 (N_46347,N_44700,N_42170);
nand U46348 (N_46348,N_43503,N_40659);
xor U46349 (N_46349,N_43460,N_41595);
nand U46350 (N_46350,N_40145,N_43139);
and U46351 (N_46351,N_44805,N_41333);
and U46352 (N_46352,N_43273,N_44435);
or U46353 (N_46353,N_43682,N_44900);
nand U46354 (N_46354,N_44565,N_43026);
xor U46355 (N_46355,N_41350,N_44693);
and U46356 (N_46356,N_43410,N_43616);
nand U46357 (N_46357,N_44931,N_44830);
nand U46358 (N_46358,N_42953,N_43549);
nor U46359 (N_46359,N_41736,N_41957);
and U46360 (N_46360,N_44470,N_41922);
nor U46361 (N_46361,N_42764,N_43346);
and U46362 (N_46362,N_43053,N_42603);
nor U46363 (N_46363,N_41500,N_43622);
or U46364 (N_46364,N_42420,N_41136);
nand U46365 (N_46365,N_41496,N_40091);
and U46366 (N_46366,N_41717,N_41911);
nor U46367 (N_46367,N_41886,N_44477);
or U46368 (N_46368,N_42136,N_40674);
or U46369 (N_46369,N_41298,N_44274);
nor U46370 (N_46370,N_40189,N_41125);
nor U46371 (N_46371,N_41216,N_42949);
nand U46372 (N_46372,N_41753,N_40835);
and U46373 (N_46373,N_40574,N_41222);
xor U46374 (N_46374,N_44989,N_41153);
or U46375 (N_46375,N_42190,N_42024);
nand U46376 (N_46376,N_42519,N_43420);
and U46377 (N_46377,N_44196,N_43915);
nor U46378 (N_46378,N_40461,N_41492);
xor U46379 (N_46379,N_43938,N_43859);
nand U46380 (N_46380,N_42996,N_43394);
and U46381 (N_46381,N_40592,N_42756);
and U46382 (N_46382,N_42056,N_43363);
nor U46383 (N_46383,N_40179,N_44000);
nand U46384 (N_46384,N_44716,N_43438);
nor U46385 (N_46385,N_44273,N_42649);
nor U46386 (N_46386,N_43295,N_43577);
nor U46387 (N_46387,N_42451,N_40645);
nand U46388 (N_46388,N_44188,N_44884);
and U46389 (N_46389,N_41602,N_43530);
and U46390 (N_46390,N_43790,N_43209);
nand U46391 (N_46391,N_42012,N_43242);
or U46392 (N_46392,N_40750,N_40149);
or U46393 (N_46393,N_41764,N_41664);
nand U46394 (N_46394,N_40824,N_40098);
and U46395 (N_46395,N_40173,N_40094);
xor U46396 (N_46396,N_44509,N_44025);
nand U46397 (N_46397,N_41889,N_44838);
nor U46398 (N_46398,N_41613,N_43846);
and U46399 (N_46399,N_43964,N_40903);
and U46400 (N_46400,N_44725,N_44607);
nor U46401 (N_46401,N_43033,N_40205);
xor U46402 (N_46402,N_42522,N_40186);
nor U46403 (N_46403,N_44654,N_41407);
nor U46404 (N_46404,N_42721,N_43662);
and U46405 (N_46405,N_40515,N_40618);
and U46406 (N_46406,N_43836,N_44759);
nand U46407 (N_46407,N_40196,N_41361);
nor U46408 (N_46408,N_40737,N_44634);
nand U46409 (N_46409,N_40924,N_40109);
nor U46410 (N_46410,N_40193,N_41795);
or U46411 (N_46411,N_44681,N_42943);
nand U46412 (N_46412,N_40238,N_40892);
nand U46413 (N_46413,N_41042,N_44885);
or U46414 (N_46414,N_44897,N_41397);
nor U46415 (N_46415,N_40915,N_41987);
nor U46416 (N_46416,N_41045,N_41566);
and U46417 (N_46417,N_40817,N_44599);
and U46418 (N_46418,N_44783,N_41725);
or U46419 (N_46419,N_41757,N_40772);
or U46420 (N_46420,N_44464,N_44251);
nand U46421 (N_46421,N_41810,N_40298);
nor U46422 (N_46422,N_42909,N_40581);
or U46423 (N_46423,N_44052,N_40591);
nand U46424 (N_46424,N_43131,N_42731);
xor U46425 (N_46425,N_41115,N_41091);
nand U46426 (N_46426,N_41733,N_40178);
xor U46427 (N_46427,N_42107,N_44292);
or U46428 (N_46428,N_40346,N_42948);
xor U46429 (N_46429,N_44804,N_42101);
nand U46430 (N_46430,N_44122,N_41438);
nand U46431 (N_46431,N_40470,N_40399);
nand U46432 (N_46432,N_41567,N_41314);
nor U46433 (N_46433,N_44163,N_40953);
nand U46434 (N_46434,N_43686,N_44724);
nor U46435 (N_46435,N_41421,N_41726);
nand U46436 (N_46436,N_41531,N_41126);
or U46437 (N_46437,N_41581,N_44490);
and U46438 (N_46438,N_44072,N_43496);
and U46439 (N_46439,N_40500,N_43144);
and U46440 (N_46440,N_40816,N_40059);
nand U46441 (N_46441,N_43457,N_43058);
and U46442 (N_46442,N_42201,N_40540);
nor U46443 (N_46443,N_40039,N_41078);
nand U46444 (N_46444,N_42599,N_40227);
nand U46445 (N_46445,N_40168,N_42336);
and U46446 (N_46446,N_42853,N_42804);
xor U46447 (N_46447,N_41638,N_42944);
and U46448 (N_46448,N_40792,N_44644);
and U46449 (N_46449,N_40171,N_43450);
nor U46450 (N_46450,N_41051,N_44817);
nand U46451 (N_46451,N_43738,N_44032);
nor U46452 (N_46452,N_43592,N_43140);
nor U46453 (N_46453,N_43636,N_42293);
xnor U46454 (N_46454,N_43286,N_42626);
nand U46455 (N_46455,N_42200,N_41716);
and U46456 (N_46456,N_44398,N_42475);
nor U46457 (N_46457,N_41827,N_41879);
or U46458 (N_46458,N_43010,N_43931);
or U46459 (N_46459,N_42834,N_44959);
or U46460 (N_46460,N_43581,N_41459);
or U46461 (N_46461,N_41335,N_43741);
nand U46462 (N_46462,N_44790,N_41208);
nand U46463 (N_46463,N_44041,N_40144);
xor U46464 (N_46464,N_40271,N_44653);
xnor U46465 (N_46465,N_41209,N_42175);
nand U46466 (N_46466,N_43371,N_41474);
xor U46467 (N_46467,N_41309,N_42777);
nor U46468 (N_46468,N_43289,N_43557);
and U46469 (N_46469,N_44105,N_42379);
nand U46470 (N_46470,N_41329,N_41135);
or U46471 (N_46471,N_41778,N_40198);
and U46472 (N_46472,N_41195,N_42628);
nand U46473 (N_46473,N_42240,N_43940);
or U46474 (N_46474,N_42711,N_44568);
nand U46475 (N_46475,N_42985,N_40764);
xor U46476 (N_46476,N_40955,N_42950);
nor U46477 (N_46477,N_40793,N_43750);
and U46478 (N_46478,N_44310,N_44803);
or U46479 (N_46479,N_41703,N_41658);
and U46480 (N_46480,N_44853,N_42958);
or U46481 (N_46481,N_43149,N_43338);
nand U46482 (N_46482,N_43811,N_42343);
xor U46483 (N_46483,N_42671,N_42613);
nand U46484 (N_46484,N_42687,N_44389);
and U46485 (N_46485,N_44781,N_43967);
nor U46486 (N_46486,N_43881,N_43159);
nand U46487 (N_46487,N_43725,N_41707);
and U46488 (N_46488,N_40232,N_40481);
nor U46489 (N_46489,N_43950,N_44040);
nor U46490 (N_46490,N_41761,N_41892);
nand U46491 (N_46491,N_42161,N_40538);
and U46492 (N_46492,N_42742,N_42617);
and U46493 (N_46493,N_43369,N_42986);
nand U46494 (N_46494,N_42588,N_44365);
nor U46495 (N_46495,N_40313,N_43559);
xor U46496 (N_46496,N_44256,N_41122);
nor U46497 (N_46497,N_43430,N_41539);
nand U46498 (N_46498,N_42453,N_42098);
nand U46499 (N_46499,N_42064,N_41167);
and U46500 (N_46500,N_42459,N_44070);
nand U46501 (N_46501,N_44635,N_42811);
and U46502 (N_46502,N_41228,N_40214);
and U46503 (N_46503,N_42294,N_44184);
and U46504 (N_46504,N_41763,N_42299);
or U46505 (N_46505,N_44826,N_42368);
and U46506 (N_46506,N_44548,N_44241);
nand U46507 (N_46507,N_40736,N_42426);
nand U46508 (N_46508,N_40327,N_43353);
nor U46509 (N_46509,N_44057,N_44928);
nand U46510 (N_46510,N_42606,N_41934);
and U46511 (N_46511,N_43962,N_44100);
nand U46512 (N_46512,N_42407,N_43089);
or U46513 (N_46513,N_42651,N_44496);
nor U46514 (N_46514,N_43412,N_42576);
or U46515 (N_46515,N_43207,N_41634);
or U46516 (N_46516,N_42758,N_40974);
xnor U46517 (N_46517,N_41622,N_44169);
xor U46518 (N_46518,N_41404,N_44230);
or U46519 (N_46519,N_41884,N_40162);
and U46520 (N_46520,N_42354,N_42781);
nand U46521 (N_46521,N_40338,N_43418);
nand U46522 (N_46522,N_41868,N_43211);
or U46523 (N_46523,N_43004,N_41173);
and U46524 (N_46524,N_44170,N_43095);
nand U46525 (N_46525,N_43737,N_43368);
nor U46526 (N_46526,N_43935,N_43255);
or U46527 (N_46527,N_41215,N_40233);
xor U46528 (N_46528,N_41662,N_44797);
and U46529 (N_46529,N_42035,N_44361);
xnor U46530 (N_46530,N_42973,N_41022);
nor U46531 (N_46531,N_40560,N_40919);
and U46532 (N_46532,N_40474,N_40390);
nand U46533 (N_46533,N_42351,N_42761);
nand U46534 (N_46534,N_44534,N_43073);
nor U46535 (N_46535,N_44073,N_42193);
xnor U46536 (N_46536,N_41099,N_40765);
and U46537 (N_46537,N_44245,N_41285);
nor U46538 (N_46538,N_40471,N_41046);
nand U46539 (N_46539,N_40413,N_44795);
or U46540 (N_46540,N_41687,N_43897);
or U46541 (N_46541,N_41554,N_43831);
nand U46542 (N_46542,N_40547,N_44098);
or U46543 (N_46543,N_41712,N_42585);
or U46544 (N_46544,N_42702,N_41948);
or U46545 (N_46545,N_41406,N_43785);
nor U46546 (N_46546,N_42759,N_42238);
nor U46547 (N_46547,N_40633,N_41493);
nor U46548 (N_46548,N_44113,N_42143);
or U46549 (N_46549,N_44005,N_41545);
and U46550 (N_46550,N_41079,N_40588);
and U46551 (N_46551,N_44949,N_42043);
xor U46552 (N_46552,N_40756,N_41014);
nand U46553 (N_46553,N_40097,N_42690);
xnor U46554 (N_46554,N_42152,N_40589);
and U46555 (N_46555,N_42327,N_42147);
xnor U46556 (N_46556,N_40888,N_44686);
and U46557 (N_46557,N_43316,N_41860);
or U46558 (N_46558,N_41280,N_41371);
nand U46559 (N_46559,N_44367,N_44214);
and U46560 (N_46560,N_42371,N_44819);
nor U46561 (N_46561,N_42577,N_44078);
nor U46562 (N_46562,N_40486,N_42263);
or U46563 (N_46563,N_44346,N_42174);
or U46564 (N_46564,N_41308,N_41825);
and U46565 (N_46565,N_44985,N_44614);
and U46566 (N_46566,N_40531,N_44117);
xnor U46567 (N_46567,N_41268,N_42000);
nand U46568 (N_46568,N_43857,N_40280);
and U46569 (N_46569,N_41808,N_41193);
xnor U46570 (N_46570,N_41139,N_40829);
and U46571 (N_46571,N_44171,N_41336);
nor U46572 (N_46572,N_40023,N_44685);
xnor U46573 (N_46573,N_44995,N_43397);
and U46574 (N_46574,N_43916,N_44818);
nand U46575 (N_46575,N_41891,N_41415);
nand U46576 (N_46576,N_40457,N_44588);
nor U46577 (N_46577,N_43411,N_40634);
nand U46578 (N_46578,N_43751,N_41671);
and U46579 (N_46579,N_42769,N_40979);
and U46580 (N_46580,N_44517,N_44106);
or U46581 (N_46581,N_42582,N_41535);
nand U46582 (N_46582,N_44079,N_43604);
nand U46583 (N_46583,N_40277,N_40163);
nor U46584 (N_46584,N_44848,N_44918);
and U46585 (N_46585,N_40057,N_42468);
nand U46586 (N_46586,N_41417,N_44315);
xnor U46587 (N_46587,N_41580,N_40558);
and U46588 (N_46588,N_41430,N_43031);
or U46589 (N_46589,N_40192,N_41544);
and U46590 (N_46590,N_44338,N_40598);
nor U46591 (N_46591,N_41518,N_42677);
and U46592 (N_46592,N_42050,N_44403);
and U46593 (N_46593,N_41728,N_41326);
and U46594 (N_46594,N_44039,N_41635);
nor U46595 (N_46595,N_40901,N_43110);
nand U46596 (N_46596,N_44765,N_42517);
nand U46597 (N_46597,N_42531,N_40956);
nand U46598 (N_46598,N_40253,N_40733);
nand U46599 (N_46599,N_44401,N_42714);
and U46600 (N_46600,N_40564,N_43034);
nand U46601 (N_46601,N_41727,N_41246);
nor U46602 (N_46602,N_43627,N_41776);
xor U46603 (N_46603,N_42427,N_41296);
xor U46604 (N_46604,N_40019,N_42660);
nand U46605 (N_46605,N_42177,N_44956);
and U46606 (N_46606,N_41144,N_42800);
nor U46607 (N_46607,N_41530,N_41526);
nand U46608 (N_46608,N_41656,N_42805);
and U46609 (N_46609,N_42029,N_41578);
nor U46610 (N_46610,N_43804,N_40617);
and U46611 (N_46611,N_40387,N_41673);
nor U46612 (N_46612,N_44886,N_41519);
and U46613 (N_46613,N_44972,N_42528);
or U46614 (N_46614,N_44015,N_42591);
or U46615 (N_46615,N_44353,N_43740);
and U46616 (N_46616,N_42215,N_41961);
xor U46617 (N_46617,N_41802,N_41132);
nor U46618 (N_46618,N_40272,N_42670);
nor U46619 (N_46619,N_43598,N_42210);
or U46620 (N_46620,N_40505,N_42329);
or U46621 (N_46621,N_42524,N_41754);
nand U46622 (N_46622,N_42966,N_40266);
xnor U46623 (N_46623,N_40184,N_42533);
nor U46624 (N_46624,N_40726,N_41425);
nand U46625 (N_46625,N_42181,N_40949);
and U46626 (N_46626,N_42696,N_42405);
nor U46627 (N_46627,N_42144,N_43227);
nand U46628 (N_46628,N_43820,N_44291);
nor U46629 (N_46629,N_43663,N_41946);
or U46630 (N_46630,N_43870,N_43993);
or U46631 (N_46631,N_43433,N_42430);
nand U46632 (N_46632,N_41779,N_44097);
nand U46633 (N_46633,N_41154,N_44916);
nand U46634 (N_46634,N_40274,N_40650);
nand U46635 (N_46635,N_42032,N_44586);
or U46636 (N_46636,N_43659,N_42983);
and U46637 (N_46637,N_41590,N_40738);
nand U46638 (N_46638,N_42703,N_41766);
xor U46639 (N_46639,N_40896,N_42234);
nand U46640 (N_46640,N_40942,N_40112);
nand U46641 (N_46641,N_44680,N_41171);
nand U46642 (N_46642,N_44825,N_42921);
or U46643 (N_46643,N_40241,N_41272);
nand U46644 (N_46644,N_44971,N_40734);
or U46645 (N_46645,N_44077,N_43508);
xor U46646 (N_46646,N_44167,N_41813);
nor U46647 (N_46647,N_41699,N_42249);
or U46648 (N_46648,N_41818,N_40751);
nor U46649 (N_46649,N_40188,N_40086);
nand U46650 (N_46650,N_44622,N_41068);
nor U46651 (N_46651,N_41589,N_44612);
nor U46652 (N_46652,N_41563,N_44731);
and U46653 (N_46653,N_44067,N_40034);
or U46654 (N_46654,N_44510,N_41770);
and U46655 (N_46655,N_40945,N_43029);
nor U46656 (N_46656,N_40879,N_40115);
nand U46657 (N_46657,N_41400,N_41119);
and U46658 (N_46658,N_43205,N_40259);
nor U46659 (N_46659,N_41182,N_44062);
and U46660 (N_46660,N_43528,N_40747);
and U46661 (N_46661,N_42505,N_44121);
nor U46662 (N_46662,N_43096,N_41092);
nor U46663 (N_46663,N_40361,N_42352);
nand U46664 (N_46664,N_42411,N_44836);
nand U46665 (N_46665,N_41570,N_41024);
xnor U46666 (N_46666,N_40963,N_40120);
and U46667 (N_46667,N_40421,N_42387);
nand U46668 (N_46668,N_41742,N_44259);
or U46669 (N_46669,N_43816,N_44194);
or U46670 (N_46670,N_43036,N_43274);
or U46671 (N_46671,N_40611,N_40881);
and U46672 (N_46672,N_40761,N_44493);
and U46673 (N_46673,N_43767,N_43190);
nor U46674 (N_46674,N_40590,N_43792);
nor U46675 (N_46675,N_41286,N_40679);
and U46676 (N_46676,N_41849,N_44939);
nor U46677 (N_46677,N_40711,N_41172);
nand U46678 (N_46678,N_44866,N_44008);
nand U46679 (N_46679,N_42598,N_43054);
nand U46680 (N_46680,N_40010,N_40951);
nor U46681 (N_46681,N_40616,N_41424);
nand U46682 (N_46682,N_42315,N_41391);
nor U46683 (N_46683,N_42198,N_40717);
nor U46684 (N_46684,N_41513,N_43602);
nand U46685 (N_46685,N_42208,N_42662);
nand U46686 (N_46686,N_42049,N_44286);
or U46687 (N_46687,N_41619,N_41069);
nand U46688 (N_46688,N_44903,N_43243);
and U46689 (N_46689,N_44590,N_41316);
xor U46690 (N_46690,N_42630,N_43309);
nand U46691 (N_46691,N_44503,N_43990);
xor U46692 (N_46692,N_43566,N_43317);
nor U46693 (N_46693,N_41978,N_44937);
xor U46694 (N_46694,N_40325,N_41241);
or U46695 (N_46695,N_44360,N_40652);
xnor U46696 (N_46696,N_41086,N_40832);
xnor U46697 (N_46697,N_42113,N_40909);
nor U46698 (N_46698,N_42251,N_42766);
nor U46699 (N_46699,N_44199,N_41797);
nand U46700 (N_46700,N_43296,N_44621);
nor U46701 (N_46701,N_41706,N_44909);
and U46702 (N_46702,N_44413,N_41276);
nor U46703 (N_46703,N_41453,N_40208);
or U46704 (N_46704,N_42361,N_42296);
and U46705 (N_46705,N_42569,N_40488);
xnor U46706 (N_46706,N_44027,N_43697);
or U46707 (N_46707,N_43712,N_42069);
nor U46708 (N_46708,N_44593,N_43064);
nor U46709 (N_46709,N_40587,N_42610);
nand U46710 (N_46710,N_42433,N_42196);
nor U46711 (N_46711,N_41650,N_42424);
nand U46712 (N_46712,N_43709,N_40147);
nand U46713 (N_46713,N_40342,N_40017);
nand U46714 (N_46714,N_40575,N_40478);
and U46715 (N_46715,N_42938,N_42580);
or U46716 (N_46716,N_43567,N_44037);
nand U46717 (N_46717,N_42890,N_44123);
nand U46718 (N_46718,N_42450,N_44915);
or U46719 (N_46719,N_41342,N_40404);
nor U46720 (N_46720,N_43873,N_42520);
nand U46721 (N_46721,N_41787,N_42127);
xor U46722 (N_46722,N_44458,N_41641);
and U46723 (N_46723,N_41025,N_44486);
nor U46724 (N_46724,N_43306,N_40742);
nor U46725 (N_46725,N_43020,N_42962);
nor U46726 (N_46726,N_43283,N_44396);
and U46727 (N_46727,N_42646,N_40907);
or U46728 (N_46728,N_42864,N_40203);
or U46729 (N_46729,N_42409,N_41147);
nor U46730 (N_46730,N_43269,N_43676);
nor U46731 (N_46731,N_43390,N_41003);
nor U46732 (N_46732,N_42045,N_42956);
nor U46733 (N_46733,N_44016,N_44386);
and U46734 (N_46734,N_40609,N_40255);
and U46735 (N_46735,N_42898,N_43898);
nand U46736 (N_46736,N_43007,N_44942);
nand U46737 (N_46737,N_44598,N_44888);
nor U46738 (N_46738,N_41977,N_40350);
nand U46739 (N_46739,N_44948,N_40036);
or U46740 (N_46740,N_43698,N_41026);
nor U46741 (N_46741,N_41942,N_40396);
nor U46742 (N_46742,N_41940,N_44872);
or U46743 (N_46743,N_43323,N_43573);
nor U46744 (N_46744,N_40111,N_41186);
and U46745 (N_46745,N_44554,N_41101);
nor U46746 (N_46746,N_40014,N_41685);
nand U46747 (N_46747,N_43083,N_44457);
nand U46748 (N_46748,N_44262,N_43218);
and U46749 (N_46749,N_40482,N_42832);
nor U46750 (N_46750,N_43808,N_44011);
or U46751 (N_46751,N_44585,N_42037);
nor U46752 (N_46752,N_41627,N_44255);
xnor U46753 (N_46753,N_43288,N_41179);
nor U46754 (N_46754,N_40165,N_41162);
xor U46755 (N_46755,N_42521,N_42887);
nor U46756 (N_46756,N_43011,N_42003);
or U46757 (N_46757,N_40307,N_41199);
and U46758 (N_46758,N_40691,N_40875);
xnor U46759 (N_46759,N_43049,N_43706);
nor U46760 (N_46760,N_42754,N_43332);
or U46761 (N_46761,N_42543,N_40825);
or U46762 (N_46762,N_43679,N_43067);
and U46763 (N_46763,N_40669,N_43435);
and U46764 (N_46764,N_41159,N_43768);
nand U46765 (N_46765,N_42612,N_40519);
and U46766 (N_46766,N_43959,N_42913);
xnor U46767 (N_46767,N_44789,N_42508);
xnor U46768 (N_46768,N_42025,N_40231);
nand U46769 (N_46769,N_42452,N_40285);
nor U46770 (N_46770,N_41323,N_42363);
or U46771 (N_46771,N_43127,N_41345);
or U46772 (N_46772,N_42665,N_40536);
nand U46773 (N_46773,N_41377,N_44120);
nand U46774 (N_46774,N_40754,N_40161);
nand U46775 (N_46775,N_41177,N_43817);
nor U46776 (N_46776,N_44594,N_40349);
xnor U46777 (N_46777,N_41082,N_40580);
and U46778 (N_46778,N_42088,N_40379);
nand U46779 (N_46779,N_40009,N_40917);
and U46780 (N_46780,N_44507,N_41201);
and U46781 (N_46781,N_41436,N_40808);
and U46782 (N_46782,N_44842,N_42915);
or U46783 (N_46783,N_44773,N_42889);
nor U46784 (N_46784,N_40431,N_40561);
and U46785 (N_46785,N_40553,N_43809);
and U46786 (N_46786,N_41189,N_43326);
nand U46787 (N_46787,N_44366,N_43491);
nand U46788 (N_46788,N_43075,N_41583);
or U46789 (N_46789,N_43434,N_43974);
or U46790 (N_46790,N_43063,N_41593);
nand U46791 (N_46791,N_40923,N_42415);
or U46792 (N_46792,N_43845,N_41200);
and U46793 (N_46793,N_42443,N_41826);
or U46794 (N_46794,N_44468,N_44045);
nand U46795 (N_46795,N_44431,N_41409);
or U46796 (N_46796,N_42806,N_44185);
nor U46797 (N_46797,N_41888,N_41482);
or U46798 (N_46798,N_41747,N_44190);
or U46799 (N_46799,N_43912,N_44136);
xor U46800 (N_46800,N_42067,N_44583);
or U46801 (N_46801,N_43238,N_41170);
or U46802 (N_46802,N_42564,N_40090);
and U46803 (N_46803,N_41857,N_41739);
nand U46804 (N_46804,N_44831,N_44953);
or U46805 (N_46805,N_41572,N_44791);
xor U46806 (N_46806,N_40807,N_40578);
nor U46807 (N_46807,N_44201,N_40943);
xor U46808 (N_46808,N_40021,N_43342);
nor U46809 (N_46809,N_44026,N_43744);
xnor U46810 (N_46810,N_41437,N_44348);
or U46811 (N_46811,N_42745,N_40211);
and U46812 (N_46812,N_43621,N_44890);
and U46813 (N_46813,N_40973,N_40420);
nor U46814 (N_46814,N_42011,N_43351);
nand U46815 (N_46815,N_40501,N_42609);
and U46816 (N_46816,N_42026,N_41899);
xor U46817 (N_46817,N_44064,N_43212);
and U46818 (N_46818,N_44986,N_41720);
xnor U46819 (N_46819,N_41357,N_43161);
and U46820 (N_46820,N_40119,N_42187);
or U46821 (N_46821,N_44323,N_42053);
nand U46822 (N_46822,N_43262,N_43732);
nand U46823 (N_46823,N_44780,N_42652);
or U46824 (N_46824,N_41704,N_40692);
or U46825 (N_46825,N_43429,N_44691);
nand U46826 (N_46826,N_43254,N_41618);
nor U46827 (N_46827,N_43102,N_41908);
nand U46828 (N_46828,N_40414,N_41959);
nor U46829 (N_46829,N_41117,N_44222);
nand U46830 (N_46830,N_43188,N_41005);
and U46831 (N_46831,N_43157,N_43170);
and U46832 (N_46832,N_44889,N_44870);
xnor U46833 (N_46833,N_40987,N_41202);
nor U46834 (N_46834,N_42469,N_40405);
and U46835 (N_46835,N_43206,N_44092);
nor U46836 (N_46836,N_42594,N_42724);
or U46837 (N_46837,N_40394,N_42491);
or U46838 (N_46838,N_40620,N_44581);
and U46839 (N_46839,N_43965,N_42184);
or U46840 (N_46840,N_41374,N_41347);
xor U46841 (N_46841,N_41608,N_40284);
or U46842 (N_46842,N_42809,N_43531);
and U46843 (N_46843,N_41302,N_44753);
nand U46844 (N_46844,N_42757,N_41349);
or U46845 (N_46845,N_44533,N_41050);
nand U46846 (N_46846,N_40364,N_43217);
xnor U46847 (N_46847,N_43119,N_43665);
xor U46848 (N_46848,N_42163,N_44944);
nand U46849 (N_46849,N_40638,N_44494);
nor U46850 (N_46850,N_43176,N_44519);
xnor U46851 (N_46851,N_40516,N_41131);
or U46852 (N_46852,N_43629,N_41677);
and U46853 (N_46853,N_40031,N_40866);
or U46854 (N_46854,N_44478,N_41031);
nand U46855 (N_46855,N_43521,N_42892);
nor U46856 (N_46856,N_43451,N_40299);
nand U46857 (N_46857,N_40275,N_41950);
xnor U46858 (N_46858,N_40676,N_40008);
nand U46859 (N_46859,N_43819,N_43514);
nand U46860 (N_46860,N_43048,N_43298);
nand U46861 (N_46861,N_42010,N_43853);
nand U46862 (N_46862,N_40532,N_44506);
nor U46863 (N_46863,N_43335,N_42373);
and U46864 (N_46864,N_41898,N_43823);
nor U46865 (N_46865,N_44152,N_43759);
and U46866 (N_46866,N_44374,N_44391);
or U46867 (N_46867,N_43753,N_41551);
nand U46868 (N_46868,N_44689,N_40559);
and U46869 (N_46869,N_40952,N_40596);
nor U46870 (N_46870,N_43556,N_41379);
nand U46871 (N_46871,N_43582,N_42608);
or U46872 (N_46872,N_44091,N_44921);
nand U46873 (N_46873,N_43366,N_40337);
nor U46874 (N_46874,N_44734,N_40412);
and U46875 (N_46875,N_43908,N_42114);
and U46876 (N_46876,N_44881,N_43983);
and U46877 (N_46877,N_43486,N_40065);
or U46878 (N_46878,N_44061,N_41043);
nand U46879 (N_46879,N_42079,N_41960);
or U46880 (N_46880,N_41058,N_44998);
nor U46881 (N_46881,N_40712,N_40121);
or U46882 (N_46882,N_41331,N_44428);
xor U46883 (N_46883,N_44415,N_41019);
xnor U46884 (N_46884,N_42116,N_42556);
or U46885 (N_46885,N_42867,N_44740);
xnor U46886 (N_46886,N_43783,N_42154);
nand U46887 (N_46887,N_44408,N_41937);
nand U46888 (N_46888,N_44459,N_43882);
xnor U46889 (N_46889,N_42810,N_41239);
nor U46890 (N_46890,N_44778,N_44714);
and U46891 (N_46891,N_44349,N_41394);
or U46892 (N_46892,N_42028,N_44704);
and U46893 (N_46893,N_44877,N_41075);
nand U46894 (N_46894,N_41370,N_40767);
and U46895 (N_46895,N_42771,N_42750);
and U46896 (N_46896,N_43417,N_44319);
and U46897 (N_46897,N_40032,N_44355);
nor U46898 (N_46898,N_42931,N_41057);
nor U46899 (N_46899,N_40651,N_44227);
nand U46900 (N_46900,N_42536,N_42456);
and U46901 (N_46901,N_44892,N_42160);
nor U46902 (N_46902,N_42275,N_42621);
xnor U46903 (N_46903,N_42722,N_43347);
nor U46904 (N_46904,N_44250,N_44514);
and U46905 (N_46905,N_42798,N_43066);
and U46906 (N_46906,N_42353,N_44913);
and U46907 (N_46907,N_41219,N_40430);
and U46908 (N_46908,N_42823,N_44923);
xor U46909 (N_46909,N_42179,N_44745);
nand U46910 (N_46910,N_42674,N_43890);
nand U46911 (N_46911,N_41835,N_43239);
nand U46912 (N_46912,N_40572,N_40206);
xnor U46913 (N_46913,N_40489,N_41740);
nand U46914 (N_46914,N_43617,N_42204);
nor U46915 (N_46915,N_43449,N_40797);
nor U46916 (N_46916,N_41773,N_40366);
nor U46917 (N_46917,N_40852,N_40730);
or U46918 (N_46918,N_42984,N_42960);
nor U46919 (N_46919,N_43893,N_43624);
nor U46920 (N_46920,N_40427,N_41262);
or U46921 (N_46921,N_41053,N_42862);
nor U46922 (N_46922,N_41158,N_44610);
nor U46923 (N_46923,N_42899,N_41483);
xor U46924 (N_46924,N_43588,N_42369);
nor U46925 (N_46925,N_41017,N_40095);
and U46926 (N_46926,N_43445,N_43590);
and U46927 (N_46927,N_44569,N_41269);
and U46928 (N_46928,N_40759,N_40551);
and U46929 (N_46929,N_41257,N_44180);
nor U46930 (N_46930,N_44508,N_42735);
nor U46931 (N_46931,N_41387,N_41184);
nor U46932 (N_46932,N_44513,N_40155);
nor U46933 (N_46933,N_42498,N_40727);
or U46934 (N_46934,N_40172,N_44203);
nor U46935 (N_46935,N_40448,N_43713);
nand U46936 (N_46936,N_43649,N_43615);
or U46937 (N_46937,N_44628,N_41750);
nand U46938 (N_46938,N_44755,N_44922);
or U46939 (N_46939,N_42305,N_40918);
or U46940 (N_46940,N_40667,N_42464);
nand U46941 (N_46941,N_42494,N_42937);
or U46942 (N_46942,N_44543,N_41842);
nand U46943 (N_46943,N_44249,N_43589);
or U46944 (N_46944,N_42634,N_41856);
nand U46945 (N_46945,N_43043,N_43365);
and U46946 (N_46946,N_42718,N_40084);
nand U46947 (N_46947,N_40411,N_44846);
nor U46948 (N_46948,N_44290,N_43696);
or U46949 (N_46949,N_41267,N_42601);
nor U46950 (N_46950,N_40541,N_42829);
or U46951 (N_46951,N_43501,N_42747);
and U46952 (N_46952,N_44749,N_41270);
nor U46953 (N_46953,N_43120,N_41645);
or U46954 (N_46954,N_43328,N_41036);
or U46955 (N_46955,N_40978,N_43922);
xor U46956 (N_46956,N_41697,N_41183);
and U46957 (N_46957,N_41332,N_44665);
and U46958 (N_46958,N_44843,N_42410);
nor U46959 (N_46959,N_42087,N_43597);
or U46960 (N_46960,N_40391,N_44247);
and U46961 (N_46961,N_42437,N_42221);
xor U46962 (N_46962,N_43800,N_40770);
nor U46963 (N_46963,N_42908,N_41803);
or U46964 (N_46964,N_44442,N_41067);
nor U46965 (N_46965,N_40224,N_40463);
nor U46966 (N_46966,N_43961,N_43408);
or U46967 (N_46967,N_42375,N_43392);
and U46968 (N_46968,N_42869,N_42367);
nor U46969 (N_46969,N_44028,N_40902);
or U46970 (N_46970,N_43077,N_42523);
or U46971 (N_46971,N_42645,N_44876);
nor U46972 (N_46972,N_44218,N_40417);
or U46973 (N_46973,N_41752,N_43304);
and U46974 (N_46974,N_42042,N_40075);
nor U46975 (N_46975,N_42673,N_43510);
nand U46976 (N_46976,N_40302,N_42457);
and U46977 (N_46977,N_44657,N_40757);
nor U46978 (N_46978,N_42873,N_43349);
and U46979 (N_46979,N_41755,N_41655);
nand U46980 (N_46980,N_44178,N_42441);
nand U46981 (N_46981,N_42684,N_40845);
and U46982 (N_46982,N_40126,N_43918);
nand U46983 (N_46983,N_44462,N_44128);
xnor U46984 (N_46984,N_43858,N_42910);
and U46985 (N_46985,N_43585,N_42881);
nor U46986 (N_46986,N_40220,N_41632);
and U46987 (N_46987,N_44378,N_44932);
nor U46988 (N_46988,N_40409,N_43643);
nand U46989 (N_46989,N_43516,N_42976);
nand U46990 (N_46990,N_44808,N_40293);
or U46991 (N_46991,N_44328,N_44882);
or U46992 (N_46992,N_43027,N_43889);
or U46993 (N_46993,N_42994,N_42618);
and U46994 (N_46994,N_40072,N_42641);
xor U46995 (N_46995,N_40583,N_41760);
nand U46996 (N_46996,N_44969,N_44266);
nor U46997 (N_46997,N_42965,N_41599);
or U46998 (N_46998,N_44854,N_43578);
nor U46999 (N_46999,N_41916,N_44529);
or U47000 (N_47000,N_43512,N_42993);
or U47001 (N_47001,N_42004,N_40900);
nand U47002 (N_47002,N_40790,N_43774);
or U47003 (N_47003,N_44531,N_41765);
or U47004 (N_47004,N_41100,N_42723);
nor U47005 (N_47005,N_42254,N_42034);
xnor U47006 (N_47006,N_44732,N_43387);
xnor U47007 (N_47007,N_41517,N_40860);
and U47008 (N_47008,N_41923,N_44479);
or U47009 (N_47009,N_44341,N_44571);
nand U47010 (N_47010,N_43630,N_40762);
nand U47011 (N_47011,N_40851,N_42423);
and U47012 (N_47012,N_41362,N_42930);
or U47013 (N_47013,N_44538,N_43285);
and U47014 (N_47014,N_42228,N_44502);
nor U47015 (N_47015,N_41434,N_44217);
nor U47016 (N_47016,N_42964,N_40441);
nor U47017 (N_47017,N_40185,N_40780);
or U47018 (N_47018,N_44983,N_44350);
or U47019 (N_47019,N_41866,N_42484);
nand U47020 (N_47020,N_40766,N_42990);
or U47021 (N_47021,N_43966,N_41363);
and U47022 (N_47022,N_44107,N_43850);
xnor U47023 (N_47023,N_40830,N_43731);
nor U47024 (N_47024,N_40315,N_43320);
or U47025 (N_47025,N_40491,N_41565);
or U47026 (N_47026,N_40656,N_40180);
nand U47027 (N_47027,N_43359,N_43611);
xnor U47028 (N_47028,N_41549,N_44157);
or U47029 (N_47029,N_41865,N_40164);
nor U47030 (N_47030,N_43282,N_40288);
and U47031 (N_47031,N_40663,N_42153);
or U47032 (N_47032,N_42401,N_40718);
and U47033 (N_47033,N_44150,N_41573);
nor U47034 (N_47034,N_42014,N_42048);
nand U47035 (N_47035,N_41166,N_40093);
nand U47036 (N_47036,N_42374,N_44793);
or U47037 (N_47037,N_40033,N_42226);
or U47038 (N_47038,N_41973,N_40183);
or U47039 (N_47039,N_40883,N_44208);
or U47040 (N_47040,N_41217,N_43555);
nor U47041 (N_47041,N_44822,N_40245);
nand U47042 (N_47042,N_42978,N_40058);
or U47043 (N_47043,N_44871,N_43199);
xor U47044 (N_47044,N_40384,N_42583);
or U47045 (N_47045,N_43042,N_42245);
and U47046 (N_47046,N_43169,N_40517);
nor U47047 (N_47047,N_41278,N_40024);
nor U47048 (N_47048,N_44168,N_42159);
nand U47049 (N_47049,N_41592,N_40051);
and U47050 (N_47050,N_44236,N_43278);
nand U47051 (N_47051,N_40977,N_41949);
nor U47052 (N_47052,N_40355,N_40043);
and U47053 (N_47053,N_44526,N_40533);
nand U47054 (N_47054,N_40795,N_44239);
nand U47055 (N_47055,N_40992,N_44742);
and U47056 (N_47056,N_42150,N_40104);
or U47057 (N_47057,N_44425,N_40219);
nor U47058 (N_47058,N_44422,N_44668);
nor U47059 (N_47059,N_41852,N_41684);
or U47060 (N_47060,N_44209,N_40880);
nand U47061 (N_47061,N_42712,N_40306);
or U47062 (N_47062,N_41691,N_40841);
nand U47063 (N_47063,N_43766,N_44133);
nand U47064 (N_47064,N_42846,N_44743);
and U47065 (N_47065,N_44089,N_40729);
or U47066 (N_47066,N_44375,N_43224);
and U47067 (N_47067,N_43919,N_44996);
or U47068 (N_47068,N_42875,N_43168);
and U47069 (N_47069,N_43260,N_41848);
nor U47070 (N_47070,N_43202,N_44589);
nand U47071 (N_47071,N_41016,N_41615);
nand U47072 (N_47072,N_41083,N_42317);
and U47073 (N_47073,N_41041,N_44212);
or U47074 (N_47074,N_44450,N_41723);
nand U47075 (N_47075,N_43825,N_40407);
and U47076 (N_47076,N_41137,N_42206);
nor U47077 (N_47077,N_43551,N_43980);
or U47078 (N_47078,N_42917,N_40079);
nor U47079 (N_47079,N_41064,N_44582);
nand U47080 (N_47080,N_44371,N_40595);
xnor U47081 (N_47081,N_41441,N_43563);
or U47082 (N_47082,N_40567,N_42428);
and U47083 (N_47083,N_42751,N_44342);
nor U47084 (N_47084,N_40565,N_40800);
and U47085 (N_47085,N_40480,N_43755);
and U47086 (N_47086,N_41462,N_44359);
nor U47087 (N_47087,N_41383,N_42463);
nand U47088 (N_47088,N_42911,N_40504);
and U47089 (N_47089,N_43603,N_41237);
nor U47090 (N_47090,N_43995,N_41013);
nor U47091 (N_47091,N_40246,N_41273);
nor U47092 (N_47092,N_41460,N_40064);
xnor U47093 (N_47093,N_44103,N_42479);
or U47094 (N_47094,N_43400,N_42553);
nand U47095 (N_47095,N_44162,N_41320);
nand U47096 (N_47096,N_41862,N_43801);
or U47097 (N_47097,N_40011,N_40935);
and U47098 (N_47098,N_41121,N_42265);
or U47099 (N_47099,N_43122,N_43300);
or U47100 (N_47100,N_40680,N_41306);
nand U47101 (N_47101,N_43059,N_42977);
or U47102 (N_47102,N_43639,N_43668);
or U47103 (N_47103,N_43587,N_41307);
xor U47104 (N_47104,N_42244,N_43330);
nand U47105 (N_47105,N_44898,N_42685);
and U47106 (N_47106,N_41097,N_42128);
xor U47107 (N_47107,N_40310,N_40773);
nor U47108 (N_47108,N_42258,N_40118);
or U47109 (N_47109,N_41906,N_42981);
and U47110 (N_47110,N_41093,N_41674);
and U47111 (N_47111,N_41562,N_41120);
xnor U47112 (N_47112,N_43452,N_44183);
or U47113 (N_47113,N_43674,N_42310);
and U47114 (N_47114,N_41521,N_40295);
nand U47115 (N_47115,N_42971,N_42951);
nor U47116 (N_47116,N_43493,N_42650);
nand U47117 (N_47117,N_43440,N_41611);
nor U47118 (N_47118,N_41102,N_43905);
nand U47119 (N_47119,N_41389,N_41312);
nor U47120 (N_47120,N_44902,N_43293);
or U47121 (N_47121,N_41648,N_41478);
nor U47122 (N_47122,N_44518,N_41218);
xnor U47123 (N_47123,N_40262,N_44424);
and U47124 (N_47124,N_43813,N_42183);
and U47125 (N_47125,N_43461,N_43308);
nand U47126 (N_47126,N_43943,N_44492);
nand U47127 (N_47127,N_41543,N_44316);
or U47128 (N_47128,N_44473,N_43796);
nor U47129 (N_47129,N_43777,N_43164);
or U47130 (N_47130,N_41936,N_41901);
or U47131 (N_47131,N_41793,N_41185);
xnor U47132 (N_47132,N_41346,N_40798);
and U47133 (N_47133,N_43565,N_41044);
and U47134 (N_47134,N_42129,N_43647);
and U47135 (N_47135,N_40447,N_44550);
or U47136 (N_47136,N_41986,N_40209);
and U47137 (N_47137,N_43345,N_44237);
nor U47138 (N_47138,N_42604,N_40352);
nor U47139 (N_47139,N_44269,N_41341);
and U47140 (N_47140,N_41130,N_43536);
nor U47141 (N_47141,N_40308,N_40791);
xor U47142 (N_47142,N_42922,N_43963);
or U47143 (N_47143,N_44735,N_40554);
xor U47144 (N_47144,N_42008,N_41380);
nand U47145 (N_47145,N_42767,N_40689);
or U47146 (N_47146,N_44649,N_43733);
xnor U47147 (N_47147,N_41675,N_43745);
nor U47148 (N_47148,N_43257,N_43987);
nand U47149 (N_47149,N_43196,N_44992);
or U47150 (N_47150,N_41702,N_40886);
xnor U47151 (N_47151,N_41076,N_43250);
or U47152 (N_47152,N_40666,N_44750);
nand U47153 (N_47153,N_40362,N_43743);
nand U47154 (N_47154,N_42615,N_42963);
nand U47155 (N_47155,N_41192,N_44409);
and U47156 (N_47156,N_43895,N_44081);
or U47157 (N_47157,N_42030,N_42689);
or U47158 (N_47158,N_44592,N_44158);
nor U47159 (N_47159,N_40990,N_40279);
or U47160 (N_47160,N_43538,N_40267);
xnor U47161 (N_47161,N_44679,N_44850);
nor U47162 (N_47162,N_40388,N_41221);
xnor U47163 (N_47163,N_40453,N_40369);
and U47164 (N_47164,N_40466,N_42584);
or U47165 (N_47165,N_43660,N_44330);
and U47166 (N_47166,N_42773,N_40548);
or U47167 (N_47167,N_40630,N_40139);
or U47168 (N_47168,N_43865,N_40827);
or U47169 (N_47169,N_42987,N_41603);
nor U47170 (N_47170,N_41412,N_44096);
and U47171 (N_47171,N_42135,N_42133);
nand U47172 (N_47172,N_43474,N_40683);
nor U47173 (N_47173,N_42124,N_44879);
nand U47174 (N_47174,N_42122,N_41559);
nand U47175 (N_47175,N_41903,N_42419);
and U47176 (N_47176,N_44630,N_43954);
nor U47177 (N_47177,N_40579,N_43601);
and U47178 (N_47178,N_41063,N_41749);
nand U47179 (N_47179,N_42362,N_40158);
nand U47180 (N_47180,N_44174,N_44914);
and U47181 (N_47181,N_41598,N_42389);
nand U47182 (N_47182,N_43372,N_40194);
nor U47183 (N_47183,N_43770,N_41870);
nor U47184 (N_47184,N_41431,N_40056);
nor U47185 (N_47185,N_41516,N_40685);
and U47186 (N_47186,N_42083,N_44240);
or U47187 (N_47187,N_43090,N_41606);
xor U47188 (N_47188,N_42125,N_44232);
nand U47189 (N_47189,N_44656,N_44154);
nor U47190 (N_47190,N_43453,N_41666);
nand U47191 (N_47191,N_43446,N_43670);
nand U47192 (N_47192,N_43076,N_41477);
nand U47193 (N_47193,N_42041,N_40576);
xor U47194 (N_47194,N_43683,N_43236);
or U47195 (N_47195,N_40247,N_42104);
nor U47196 (N_47196,N_42503,N_41995);
or U47197 (N_47197,N_42945,N_43822);
or U47198 (N_47198,N_42880,N_42394);
nand U47199 (N_47199,N_43560,N_41532);
or U47200 (N_47200,N_44632,N_43724);
nand U47201 (N_47201,N_42672,N_43100);
and U47202 (N_47202,N_43177,N_43213);
nor U47203 (N_47203,N_43130,N_43700);
xnor U47204 (N_47204,N_41636,N_40731);
nor U47205 (N_47205,N_40499,N_42062);
nand U47206 (N_47206,N_44987,N_44966);
nor U47207 (N_47207,N_40976,N_42839);
and U47208 (N_47208,N_41138,N_40778);
or U47209 (N_47209,N_41783,N_43099);
and U47210 (N_47210,N_42772,N_40423);
and U47211 (N_47211,N_43669,N_44499);
nand U47212 (N_47212,N_42380,N_41033);
or U47213 (N_47213,N_41247,N_43097);
or U47214 (N_47214,N_43080,N_42740);
and U47215 (N_47215,N_41034,N_40814);
or U47216 (N_47216,N_40142,N_42516);
nand U47217 (N_47217,N_41550,N_43221);
and U47218 (N_47218,N_42734,N_44102);
and U47219 (N_47219,N_44960,N_40544);
nand U47220 (N_47220,N_41021,N_41224);
xor U47221 (N_47221,N_41564,N_44480);
or U47222 (N_47222,N_44840,N_41318);
or U47223 (N_47223,N_40046,N_43848);
nor U47224 (N_47224,N_40948,N_42787);
nand U47225 (N_47225,N_42851,N_42695);
and U47226 (N_47226,N_44864,N_43505);
nor U47227 (N_47227,N_42694,N_43112);
and U47228 (N_47228,N_43932,N_44144);
nand U47229 (N_47229,N_40082,N_41895);
and U47230 (N_47230,N_42320,N_41012);
nand U47231 (N_47231,N_42620,N_40487);
and U47232 (N_47232,N_42274,N_42982);
nand U47233 (N_47233,N_41227,N_40913);
or U47234 (N_47234,N_44242,N_44615);
nand U47235 (N_47235,N_41381,N_42581);
and U47236 (N_47236,N_43038,N_44712);
nor U47237 (N_47237,N_40365,N_40884);
and U47238 (N_47238,N_40402,N_40393);
nand U47239 (N_47239,N_44777,N_42954);
nor U47240 (N_47240,N_43562,N_43071);
nor U47241 (N_47241,N_43976,N_43855);
nand U47242 (N_47242,N_43623,N_40318);
and U47243 (N_47243,N_42901,N_43608);
or U47244 (N_47244,N_42602,N_43125);
or U47245 (N_47245,N_41015,N_44784);
nand U47246 (N_47246,N_42850,N_44110);
or U47247 (N_47247,N_42865,N_42253);
nand U47248 (N_47248,N_41256,N_40381);
and U47249 (N_47249,N_41823,N_40641);
nor U47250 (N_47250,N_40124,N_40215);
xor U47251 (N_47251,N_41847,N_44557);
nor U47252 (N_47252,N_44901,N_44204);
nor U47253 (N_47253,N_42218,N_42347);
and U47254 (N_47254,N_44485,N_40234);
xor U47255 (N_47255,N_40597,N_40328);
and U47256 (N_47256,N_44991,N_44962);
or U47257 (N_47257,N_42192,N_43644);
or U47258 (N_47258,N_44388,N_40523);
and U47259 (N_47259,N_41052,N_41745);
xnor U47260 (N_47260,N_40428,N_41994);
and U47261 (N_47261,N_42444,N_40804);
xor U47262 (N_47262,N_44527,N_43673);
nor U47263 (N_47263,N_41854,N_43868);
and U47264 (N_47264,N_40106,N_40524);
and U47265 (N_47265,N_43210,N_43465);
nand U47266 (N_47266,N_40329,N_41240);
or U47267 (N_47267,N_44407,N_42117);
or U47268 (N_47268,N_43472,N_41352);
xor U47269 (N_47269,N_43301,N_40061);
nand U47270 (N_47270,N_42186,N_44904);
nand U47271 (N_47271,N_44051,N_40831);
and U47272 (N_47272,N_43471,N_43764);
nor U47273 (N_47273,N_43971,N_41204);
or U47274 (N_47274,N_44445,N_43648);
or U47275 (N_47275,N_42676,N_40389);
or U47276 (N_47276,N_41621,N_44160);
xnor U47277 (N_47277,N_44373,N_42705);
xor U47278 (N_47278,N_43933,N_43547);
nor U47279 (N_47279,N_42497,N_43488);
nor U47280 (N_47280,N_43339,N_42529);
xnor U47281 (N_47281,N_40926,N_43003);
nor U47282 (N_47282,N_41356,N_40834);
or U47283 (N_47283,N_40715,N_42146);
nor U47284 (N_47284,N_44865,N_43340);
nor U47285 (N_47285,N_41525,N_41277);
xor U47286 (N_47286,N_44380,N_43509);
or U47287 (N_47287,N_44576,N_40167);
nand U47288 (N_47288,N_44153,N_40562);
or U47289 (N_47289,N_41874,N_41334);
xnor U47290 (N_47290,N_42462,N_44293);
or U47291 (N_47291,N_43626,N_40341);
or U47292 (N_47292,N_41090,N_40844);
xnor U47293 (N_47293,N_42746,N_40437);
or U47294 (N_47294,N_42501,N_41651);
nor U47295 (N_47295,N_41926,N_40753);
and U47296 (N_47296,N_40452,N_42549);
or U47297 (N_47297,N_43107,N_41454);
nor U47298 (N_47298,N_40602,N_43072);
nand U47299 (N_47299,N_40999,N_41446);
and U47300 (N_47300,N_41800,N_42489);
and U47301 (N_47301,N_43511,N_40873);
nor U47302 (N_47302,N_42707,N_44993);
nor U47303 (N_47303,N_43230,N_43225);
and U47304 (N_47304,N_43427,N_43568);
and U47305 (N_47305,N_41596,N_44629);
nor U47306 (N_47306,N_43776,N_43376);
nor U47307 (N_47307,N_43113,N_42635);
nor U47308 (N_47308,N_40473,N_44446);
nor U47309 (N_47309,N_43771,N_43280);
and U47310 (N_47310,N_43086,N_42357);
nand U47311 (N_47311,N_44869,N_44579);
or U47312 (N_47312,N_40721,N_41794);
nand U47313 (N_47313,N_42386,N_42300);
and U47314 (N_47314,N_41504,N_41990);
or U47315 (N_47315,N_43005,N_40658);
and U47316 (N_47316,N_44302,N_44440);
or U47317 (N_47317,N_40242,N_40890);
or U47318 (N_47318,N_43885,N_42871);
nand U47319 (N_47319,N_44397,N_42808);
nand U47320 (N_47320,N_40725,N_40276);
nor U47321 (N_47321,N_42350,N_43060);
nor U47322 (N_47322,N_43082,N_43722);
nor U47323 (N_47323,N_40914,N_43329);
xor U47324 (N_47324,N_42220,N_42647);
and U47325 (N_47325,N_40934,N_42118);
and U47326 (N_47326,N_42631,N_40784);
nand U47327 (N_47327,N_43084,N_40483);
nor U47328 (N_47328,N_41956,N_40069);
nor U47329 (N_47329,N_43812,N_41291);
nand U47330 (N_47330,N_43259,N_42715);
xnor U47331 (N_47331,N_40933,N_43704);
nand U47332 (N_47332,N_44906,N_44650);
or U47333 (N_47333,N_40671,N_43833);
and U47334 (N_47334,N_40330,N_43495);
nand U47335 (N_47335,N_44684,N_44466);
nor U47336 (N_47336,N_43182,N_41780);
xnor U47337 (N_47337,N_42006,N_41705);
nand U47338 (N_47338,N_40281,N_42321);
nor U47339 (N_47339,N_44031,N_42486);
and U47340 (N_47340,N_44841,N_40843);
nand U47341 (N_47341,N_43594,N_42928);
and U47342 (N_47342,N_40426,N_43370);
or U47343 (N_47343,N_41465,N_42592);
or U47344 (N_47344,N_43436,N_42632);
and U47345 (N_47345,N_41657,N_41249);
and U47346 (N_47346,N_40166,N_43901);
or U47347 (N_47347,N_44275,N_42476);
and U47348 (N_47348,N_44179,N_43331);
nand U47349 (N_47349,N_44874,N_40806);
nor U47350 (N_47350,N_41077,N_42291);
or U47351 (N_47351,N_41181,N_40842);
xor U47352 (N_47352,N_41552,N_43028);
and U47353 (N_47353,N_42607,N_43267);
nor U47354 (N_47354,N_44111,N_41004);
nor U47355 (N_47355,N_44561,N_42924);
nor U47356 (N_47356,N_43999,N_43728);
nand U47357 (N_47357,N_42396,N_44964);
or U47358 (N_47358,N_40714,N_40377);
and U47359 (N_47359,N_43924,N_44814);
and U47360 (N_47360,N_42493,N_42768);
or U47361 (N_47361,N_42959,N_42203);
and U47362 (N_47362,N_40117,N_44181);
or U47363 (N_47363,N_41624,N_42512);
xor U47364 (N_47364,N_42370,N_40040);
xor U47365 (N_47365,N_43838,N_41178);
nor U47366 (N_47366,N_43818,N_41165);
and U47367 (N_47367,N_44159,N_44720);
or U47368 (N_47368,N_40005,N_41339);
nand U47369 (N_47369,N_42844,N_41824);
or U47370 (N_47370,N_44387,N_41683);
or U47371 (N_47371,N_44453,N_44834);
and U47372 (N_47372,N_42229,N_43877);
and U47373 (N_47373,N_40603,N_43487);
or U47374 (N_47374,N_44191,N_44688);
and U47375 (N_47375,N_43271,N_43747);
nor U47376 (N_47376,N_41008,N_42547);
nand U47377 (N_47377,N_40988,N_41737);
and U47378 (N_47378,N_43596,N_40464);
or U47379 (N_47379,N_42872,N_44216);
nand U47380 (N_47380,N_43803,N_41591);
xor U47381 (N_47381,N_43315,N_41244);
or U47382 (N_47382,N_42499,N_44601);
nand U47383 (N_47383,N_44660,N_44990);
or U47384 (N_47384,N_43241,N_44099);
nand U47385 (N_47385,N_42697,N_40774);
nor U47386 (N_47386,N_40997,N_43476);
nor U47387 (N_47387,N_43379,N_42884);
nand U47388 (N_47388,N_43383,N_41245);
and U47389 (N_47389,N_42059,N_43798);
and U47390 (N_47390,N_40223,N_43886);
nor U47391 (N_47391,N_40324,N_40655);
nor U47392 (N_47392,N_44566,N_43470);
nor U47393 (N_47393,N_40614,N_41214);
nor U47394 (N_47394,N_40749,N_43219);
or U47395 (N_47395,N_41088,N_42669);
nand U47396 (N_47396,N_44205,N_43245);
or U47397 (N_47397,N_44868,N_44536);
nor U47398 (N_47398,N_40836,N_44109);
and U47399 (N_47399,N_44358,N_41741);
and U47400 (N_47400,N_40170,N_44852);
xnor U47401 (N_47401,N_44337,N_41364);
xnor U47402 (N_47402,N_42490,N_44767);
nand U47403 (N_47403,N_44899,N_44059);
nand U47404 (N_47404,N_40889,N_43462);
and U47405 (N_47405,N_41881,N_43361);
and U47406 (N_47406,N_44314,N_42273);
xnor U47407 (N_47407,N_41984,N_40623);
nand U47408 (N_47408,N_44381,N_42782);
or U47409 (N_47409,N_40546,N_40991);
nand U47410 (N_47410,N_44125,N_42284);
nor U47411 (N_47411,N_42077,N_42894);
and U47412 (N_47412,N_42167,N_43942);
xnor U47413 (N_47413,N_41971,N_43934);
nor U47414 (N_47414,N_40625,N_40735);
nor U47415 (N_47415,N_40569,N_41315);
or U47416 (N_47416,N_44343,N_44281);
xor U47417 (N_47417,N_40213,N_42866);
nor U47418 (N_47418,N_41616,N_44973);
nor U47419 (N_47419,N_40433,N_43529);
xnor U47420 (N_47420,N_44613,N_44847);
and U47421 (N_47421,N_44449,N_40475);
nor U47422 (N_47422,N_42070,N_43275);
and U47423 (N_47423,N_40260,N_40989);
or U47424 (N_47424,N_44861,N_42036);
nand U47425 (N_47425,N_41542,N_42082);
nand U47426 (N_47426,N_40225,N_42313);
and U47427 (N_47427,N_41486,N_43781);
or U47428 (N_47428,N_43705,N_40322);
nor U47429 (N_47429,N_43500,N_40527);
nor U47430 (N_47430,N_43109,N_44970);
nor U47431 (N_47431,N_43407,N_43929);
or U47432 (N_47432,N_42802,N_43527);
nor U47433 (N_47433,N_44427,N_44984);
and U47434 (N_47434,N_44955,N_42267);
nor U47435 (N_47435,N_43479,N_42348);
and U47436 (N_47436,N_43362,N_41305);
and U47437 (N_47437,N_40221,N_41719);
xnor U47438 (N_47438,N_44729,N_42121);
and U47439 (N_47439,N_41735,N_43163);
nand U47440 (N_47440,N_41282,N_42478);
nor U47441 (N_47441,N_42397,N_43189);
nor U47442 (N_47442,N_43281,N_41410);
nor U47443 (N_47443,N_41433,N_41322);
and U47444 (N_47444,N_41781,N_41597);
nor U47445 (N_47445,N_43137,N_44965);
nand U47446 (N_47446,N_41207,N_42376);
nand U47447 (N_47447,N_42382,N_41365);
nand U47448 (N_47448,N_44345,N_40029);
or U47449 (N_47449,N_42952,N_44175);
xor U47450 (N_47450,N_42513,N_44945);
nand U47451 (N_47451,N_43828,N_43357);
or U47452 (N_47452,N_43166,N_44288);
nand U47453 (N_47453,N_42822,N_44145);
and U47454 (N_47454,N_42487,N_44967);
nand U47455 (N_47455,N_40442,N_41534);
nor U47456 (N_47456,N_40347,N_40143);
xnor U47457 (N_47457,N_40465,N_41659);
or U47458 (N_47458,N_43518,N_41351);
nand U47459 (N_47459,N_44552,N_40314);
nand U47460 (N_47460,N_42020,N_44596);
nand U47461 (N_47461,N_41321,N_42558);
and U47462 (N_47462,N_40278,N_42624);
nand U47463 (N_47463,N_41817,N_42219);
nand U47464 (N_47464,N_44832,N_42195);
nor U47465 (N_47465,N_41969,N_40708);
or U47466 (N_47466,N_43444,N_42858);
and U47467 (N_47467,N_43775,N_42923);
nand U47468 (N_47468,N_44384,N_40743);
and U47469 (N_47469,N_43204,N_40539);
nor U47470 (N_47470,N_43088,N_42194);
nor U47471 (N_47471,N_44696,N_43715);
or U47472 (N_47472,N_42316,N_43876);
nor U47473 (N_47473,N_40984,N_40904);
nand U47474 (N_47474,N_41428,N_43312);
xor U47475 (N_47475,N_42744,N_42485);
xor U47476 (N_47476,N_42701,N_44752);
and U47477 (N_47477,N_43535,N_43442);
or U47478 (N_47478,N_43748,N_41392);
and U47479 (N_47479,N_40626,N_42639);
nand U47480 (N_47480,N_43106,N_43497);
nor U47481 (N_47481,N_41196,N_44132);
nor U47482 (N_47482,N_44452,N_41734);
xnor U47483 (N_47483,N_40876,N_43507);
and U47484 (N_47484,N_43409,N_44410);
and U47485 (N_47485,N_44633,N_40872);
nor U47486 (N_47486,N_44308,N_41548);
nand U47487 (N_47487,N_41743,N_44352);
and U47488 (N_47488,N_40368,N_44363);
or U47489 (N_47489,N_40628,N_43892);
nand U47490 (N_47490,N_44722,N_40855);
xnor U47491 (N_47491,N_42970,N_43606);
xor U47492 (N_47492,N_40684,N_40261);
nor U47493 (N_47493,N_43802,N_42563);
nand U47494 (N_47494,N_42145,N_43525);
xor U47495 (N_47495,N_43852,N_40015);
nor U47496 (N_47496,N_40013,N_42318);
nor U47497 (N_47497,N_40982,N_41213);
nand U47498 (N_47498,N_40450,N_41475);
nand U47499 (N_47499,N_41721,N_42131);
nand U47500 (N_47500,N_43941,N_41446);
or U47501 (N_47501,N_42754,N_44090);
nand U47502 (N_47502,N_44758,N_43588);
or U47503 (N_47503,N_40012,N_43236);
and U47504 (N_47504,N_40272,N_40827);
or U47505 (N_47505,N_40463,N_44595);
and U47506 (N_47506,N_41150,N_41723);
and U47507 (N_47507,N_40740,N_41384);
nor U47508 (N_47508,N_44837,N_42084);
or U47509 (N_47509,N_42532,N_41490);
nand U47510 (N_47510,N_41674,N_42645);
nand U47511 (N_47511,N_43787,N_41747);
or U47512 (N_47512,N_44384,N_43040);
nand U47513 (N_47513,N_44571,N_43269);
nor U47514 (N_47514,N_44172,N_40629);
or U47515 (N_47515,N_43409,N_42120);
or U47516 (N_47516,N_44559,N_43290);
or U47517 (N_47517,N_43951,N_43228);
and U47518 (N_47518,N_42787,N_40410);
and U47519 (N_47519,N_41526,N_41924);
xnor U47520 (N_47520,N_43333,N_43500);
and U47521 (N_47521,N_44424,N_44236);
or U47522 (N_47522,N_44310,N_40656);
or U47523 (N_47523,N_44048,N_40539);
nand U47524 (N_47524,N_44608,N_44395);
or U47525 (N_47525,N_42619,N_44266);
nand U47526 (N_47526,N_43045,N_41159);
nor U47527 (N_47527,N_43025,N_40616);
and U47528 (N_47528,N_41907,N_44921);
nor U47529 (N_47529,N_43515,N_41457);
nor U47530 (N_47530,N_43761,N_44790);
or U47531 (N_47531,N_43090,N_43146);
and U47532 (N_47532,N_44874,N_43896);
nand U47533 (N_47533,N_41728,N_42473);
and U47534 (N_47534,N_42398,N_43024);
and U47535 (N_47535,N_43709,N_43772);
and U47536 (N_47536,N_44144,N_42276);
nand U47537 (N_47537,N_40487,N_41963);
xor U47538 (N_47538,N_41005,N_41078);
or U47539 (N_47539,N_42084,N_40293);
nor U47540 (N_47540,N_40643,N_44296);
or U47541 (N_47541,N_44933,N_43517);
nor U47542 (N_47542,N_42580,N_43090);
and U47543 (N_47543,N_42843,N_44474);
or U47544 (N_47544,N_40430,N_40631);
and U47545 (N_47545,N_44458,N_42166);
or U47546 (N_47546,N_44581,N_44819);
xnor U47547 (N_47547,N_44589,N_44414);
or U47548 (N_47548,N_41210,N_41492);
xnor U47549 (N_47549,N_42137,N_41364);
nand U47550 (N_47550,N_44570,N_42883);
nor U47551 (N_47551,N_42814,N_43413);
nor U47552 (N_47552,N_41725,N_44539);
nand U47553 (N_47553,N_40115,N_43080);
nand U47554 (N_47554,N_41841,N_42342);
and U47555 (N_47555,N_41143,N_44875);
xnor U47556 (N_47556,N_43723,N_44681);
nor U47557 (N_47557,N_44924,N_40692);
or U47558 (N_47558,N_43928,N_40140);
nor U47559 (N_47559,N_43964,N_44690);
and U47560 (N_47560,N_44624,N_40840);
and U47561 (N_47561,N_41301,N_40199);
nor U47562 (N_47562,N_42323,N_40573);
or U47563 (N_47563,N_44017,N_41377);
nor U47564 (N_47564,N_42620,N_41432);
nand U47565 (N_47565,N_42727,N_44724);
and U47566 (N_47566,N_40052,N_41378);
and U47567 (N_47567,N_42600,N_42709);
or U47568 (N_47568,N_43573,N_42522);
nor U47569 (N_47569,N_43856,N_41904);
nand U47570 (N_47570,N_43119,N_43553);
nand U47571 (N_47571,N_40054,N_41303);
xnor U47572 (N_47572,N_40131,N_40010);
or U47573 (N_47573,N_40490,N_44331);
and U47574 (N_47574,N_40753,N_44592);
or U47575 (N_47575,N_43447,N_42947);
xnor U47576 (N_47576,N_43503,N_40283);
nor U47577 (N_47577,N_44646,N_44269);
or U47578 (N_47578,N_44993,N_43912);
xor U47579 (N_47579,N_44541,N_42221);
nor U47580 (N_47580,N_40970,N_44354);
or U47581 (N_47581,N_43979,N_41632);
xor U47582 (N_47582,N_43873,N_41547);
or U47583 (N_47583,N_42258,N_43846);
nor U47584 (N_47584,N_41853,N_40407);
or U47585 (N_47585,N_41019,N_42405);
nor U47586 (N_47586,N_41485,N_44824);
nor U47587 (N_47587,N_41126,N_41138);
or U47588 (N_47588,N_43807,N_40778);
and U47589 (N_47589,N_43818,N_42875);
and U47590 (N_47590,N_44199,N_41469);
nor U47591 (N_47591,N_44349,N_44845);
nand U47592 (N_47592,N_42751,N_43143);
or U47593 (N_47593,N_41241,N_43515);
or U47594 (N_47594,N_40663,N_41350);
and U47595 (N_47595,N_42571,N_41552);
or U47596 (N_47596,N_43203,N_43256);
and U47597 (N_47597,N_40882,N_40303);
or U47598 (N_47598,N_40418,N_43307);
or U47599 (N_47599,N_42872,N_44394);
nand U47600 (N_47600,N_44345,N_41826);
nand U47601 (N_47601,N_43166,N_43616);
nor U47602 (N_47602,N_40701,N_43684);
nor U47603 (N_47603,N_43370,N_40746);
nor U47604 (N_47604,N_44944,N_42877);
nand U47605 (N_47605,N_43862,N_40806);
nor U47606 (N_47606,N_41001,N_44256);
xnor U47607 (N_47607,N_43626,N_41531);
nand U47608 (N_47608,N_40194,N_40197);
nor U47609 (N_47609,N_41392,N_41793);
xor U47610 (N_47610,N_40799,N_40462);
nor U47611 (N_47611,N_41909,N_44637);
nor U47612 (N_47612,N_43791,N_44706);
or U47613 (N_47613,N_40804,N_40867);
and U47614 (N_47614,N_43288,N_41189);
or U47615 (N_47615,N_43102,N_43047);
nand U47616 (N_47616,N_41822,N_43332);
and U47617 (N_47617,N_43994,N_43414);
xor U47618 (N_47618,N_40598,N_43877);
nand U47619 (N_47619,N_42308,N_40683);
and U47620 (N_47620,N_40541,N_43065);
and U47621 (N_47621,N_40769,N_42128);
nor U47622 (N_47622,N_41058,N_44994);
and U47623 (N_47623,N_44518,N_41414);
or U47624 (N_47624,N_42818,N_42162);
and U47625 (N_47625,N_43781,N_40611);
nor U47626 (N_47626,N_41302,N_42055);
and U47627 (N_47627,N_44213,N_44006);
nor U47628 (N_47628,N_44697,N_43071);
nor U47629 (N_47629,N_42379,N_41925);
nor U47630 (N_47630,N_41741,N_41743);
nand U47631 (N_47631,N_40713,N_40185);
nand U47632 (N_47632,N_43106,N_41938);
xnor U47633 (N_47633,N_40921,N_41952);
nor U47634 (N_47634,N_40424,N_44264);
and U47635 (N_47635,N_41828,N_43104);
nor U47636 (N_47636,N_42312,N_43026);
nand U47637 (N_47637,N_41106,N_43241);
and U47638 (N_47638,N_41670,N_40923);
and U47639 (N_47639,N_40258,N_40185);
and U47640 (N_47640,N_43518,N_44242);
or U47641 (N_47641,N_43495,N_43469);
and U47642 (N_47642,N_41016,N_44907);
or U47643 (N_47643,N_40209,N_43355);
nor U47644 (N_47644,N_42266,N_43381);
nand U47645 (N_47645,N_44340,N_43486);
nand U47646 (N_47646,N_42898,N_41990);
nor U47647 (N_47647,N_40755,N_44462);
nor U47648 (N_47648,N_42354,N_40156);
and U47649 (N_47649,N_40779,N_43590);
nor U47650 (N_47650,N_41982,N_44245);
and U47651 (N_47651,N_43501,N_43916);
and U47652 (N_47652,N_41115,N_43040);
nor U47653 (N_47653,N_40966,N_44830);
or U47654 (N_47654,N_44723,N_43289);
nand U47655 (N_47655,N_44661,N_41065);
and U47656 (N_47656,N_41697,N_41456);
and U47657 (N_47657,N_44427,N_40281);
nand U47658 (N_47658,N_41310,N_41453);
nand U47659 (N_47659,N_41031,N_40541);
and U47660 (N_47660,N_42193,N_44070);
or U47661 (N_47661,N_41695,N_42808);
or U47662 (N_47662,N_43896,N_42808);
and U47663 (N_47663,N_44740,N_44273);
nand U47664 (N_47664,N_44514,N_43869);
or U47665 (N_47665,N_41684,N_44037);
xnor U47666 (N_47666,N_43000,N_43365);
and U47667 (N_47667,N_44344,N_41242);
nand U47668 (N_47668,N_43946,N_44070);
or U47669 (N_47669,N_40241,N_42298);
and U47670 (N_47670,N_42932,N_42611);
nand U47671 (N_47671,N_43697,N_42188);
or U47672 (N_47672,N_44527,N_44794);
and U47673 (N_47673,N_44665,N_44586);
and U47674 (N_47674,N_43682,N_42388);
and U47675 (N_47675,N_44585,N_40539);
xor U47676 (N_47676,N_42001,N_42395);
xnor U47677 (N_47677,N_40795,N_44797);
or U47678 (N_47678,N_42141,N_42989);
xnor U47679 (N_47679,N_43890,N_40285);
nand U47680 (N_47680,N_41027,N_44925);
nor U47681 (N_47681,N_40581,N_44215);
nand U47682 (N_47682,N_41322,N_40739);
nand U47683 (N_47683,N_44587,N_41955);
xor U47684 (N_47684,N_44225,N_43026);
and U47685 (N_47685,N_41417,N_43793);
nand U47686 (N_47686,N_40796,N_44685);
and U47687 (N_47687,N_42174,N_42935);
or U47688 (N_47688,N_44027,N_44191);
nand U47689 (N_47689,N_43059,N_42571);
xnor U47690 (N_47690,N_41538,N_40741);
or U47691 (N_47691,N_43869,N_40012);
and U47692 (N_47692,N_44607,N_42046);
nor U47693 (N_47693,N_44773,N_43795);
nor U47694 (N_47694,N_42894,N_44233);
nor U47695 (N_47695,N_41554,N_42425);
xor U47696 (N_47696,N_43351,N_41050);
or U47697 (N_47697,N_43757,N_41202);
nor U47698 (N_47698,N_44248,N_41351);
nand U47699 (N_47699,N_43280,N_43489);
or U47700 (N_47700,N_40639,N_44308);
and U47701 (N_47701,N_41111,N_44400);
nand U47702 (N_47702,N_42863,N_42281);
nor U47703 (N_47703,N_40744,N_44748);
nand U47704 (N_47704,N_42733,N_42619);
or U47705 (N_47705,N_43279,N_42184);
nor U47706 (N_47706,N_40488,N_44992);
and U47707 (N_47707,N_42583,N_41171);
nand U47708 (N_47708,N_42282,N_41529);
and U47709 (N_47709,N_41134,N_41117);
nor U47710 (N_47710,N_44398,N_42082);
or U47711 (N_47711,N_41325,N_42545);
xor U47712 (N_47712,N_41392,N_44465);
or U47713 (N_47713,N_43992,N_44174);
and U47714 (N_47714,N_44871,N_42130);
or U47715 (N_47715,N_44193,N_43797);
xor U47716 (N_47716,N_41446,N_43735);
nand U47717 (N_47717,N_41075,N_40726);
and U47718 (N_47718,N_42949,N_44843);
or U47719 (N_47719,N_40922,N_40456);
xnor U47720 (N_47720,N_42453,N_40314);
nor U47721 (N_47721,N_42115,N_43766);
or U47722 (N_47722,N_42950,N_42572);
or U47723 (N_47723,N_43908,N_40598);
or U47724 (N_47724,N_40274,N_42242);
or U47725 (N_47725,N_43350,N_44592);
or U47726 (N_47726,N_44014,N_44800);
xor U47727 (N_47727,N_41063,N_42042);
and U47728 (N_47728,N_42527,N_41472);
nor U47729 (N_47729,N_43845,N_43228);
nand U47730 (N_47730,N_44519,N_40762);
nor U47731 (N_47731,N_41957,N_41617);
nor U47732 (N_47732,N_43517,N_44000);
and U47733 (N_47733,N_43021,N_40024);
and U47734 (N_47734,N_43939,N_41708);
and U47735 (N_47735,N_43000,N_43806);
nor U47736 (N_47736,N_44230,N_44305);
nor U47737 (N_47737,N_41035,N_40252);
and U47738 (N_47738,N_42063,N_44607);
and U47739 (N_47739,N_40919,N_43770);
and U47740 (N_47740,N_40372,N_42498);
or U47741 (N_47741,N_42964,N_42607);
nand U47742 (N_47742,N_41385,N_41367);
nand U47743 (N_47743,N_41565,N_44431);
nand U47744 (N_47744,N_40355,N_40687);
and U47745 (N_47745,N_44458,N_42661);
xnor U47746 (N_47746,N_42043,N_41817);
nand U47747 (N_47747,N_40887,N_41396);
and U47748 (N_47748,N_43062,N_42177);
xor U47749 (N_47749,N_41989,N_43540);
xnor U47750 (N_47750,N_41276,N_44988);
or U47751 (N_47751,N_43603,N_41927);
or U47752 (N_47752,N_43651,N_40011);
nand U47753 (N_47753,N_43088,N_44151);
nand U47754 (N_47754,N_42669,N_41133);
nor U47755 (N_47755,N_43166,N_42437);
or U47756 (N_47756,N_43110,N_42457);
nand U47757 (N_47757,N_41217,N_42545);
and U47758 (N_47758,N_40394,N_42014);
nand U47759 (N_47759,N_44529,N_44700);
nor U47760 (N_47760,N_44734,N_44536);
nor U47761 (N_47761,N_41018,N_40945);
and U47762 (N_47762,N_42656,N_41283);
and U47763 (N_47763,N_42578,N_41947);
xnor U47764 (N_47764,N_42185,N_42901);
nand U47765 (N_47765,N_41868,N_43977);
nor U47766 (N_47766,N_41102,N_43546);
nor U47767 (N_47767,N_40065,N_41665);
nand U47768 (N_47768,N_42616,N_41292);
nor U47769 (N_47769,N_43788,N_44238);
or U47770 (N_47770,N_40024,N_44699);
nor U47771 (N_47771,N_42876,N_41292);
nor U47772 (N_47772,N_42542,N_40980);
nor U47773 (N_47773,N_44459,N_44823);
nor U47774 (N_47774,N_43966,N_40405);
or U47775 (N_47775,N_44369,N_42863);
nand U47776 (N_47776,N_44459,N_43749);
and U47777 (N_47777,N_40984,N_41897);
nand U47778 (N_47778,N_44863,N_43922);
xnor U47779 (N_47779,N_41497,N_43177);
nand U47780 (N_47780,N_43296,N_42894);
or U47781 (N_47781,N_44089,N_41239);
nor U47782 (N_47782,N_40849,N_40826);
nand U47783 (N_47783,N_40528,N_41177);
or U47784 (N_47784,N_43906,N_40492);
nor U47785 (N_47785,N_43970,N_43767);
or U47786 (N_47786,N_40242,N_42415);
nand U47787 (N_47787,N_41133,N_44440);
or U47788 (N_47788,N_42768,N_42439);
nor U47789 (N_47789,N_44081,N_42163);
and U47790 (N_47790,N_42537,N_43741);
nor U47791 (N_47791,N_43237,N_44752);
nand U47792 (N_47792,N_43999,N_44723);
or U47793 (N_47793,N_42535,N_40831);
nor U47794 (N_47794,N_42332,N_40275);
and U47795 (N_47795,N_41453,N_40545);
nand U47796 (N_47796,N_44134,N_43701);
nand U47797 (N_47797,N_40531,N_40803);
nor U47798 (N_47798,N_43343,N_43273);
nand U47799 (N_47799,N_43026,N_42779);
nor U47800 (N_47800,N_43400,N_42113);
nand U47801 (N_47801,N_43217,N_41599);
and U47802 (N_47802,N_42047,N_42434);
and U47803 (N_47803,N_43924,N_42943);
nand U47804 (N_47804,N_43335,N_40671);
nand U47805 (N_47805,N_40056,N_43501);
nand U47806 (N_47806,N_42706,N_43534);
nor U47807 (N_47807,N_44791,N_42647);
xnor U47808 (N_47808,N_40475,N_44001);
nand U47809 (N_47809,N_41706,N_43880);
or U47810 (N_47810,N_44512,N_40076);
or U47811 (N_47811,N_41934,N_43207);
and U47812 (N_47812,N_40748,N_43687);
nor U47813 (N_47813,N_44443,N_43249);
xor U47814 (N_47814,N_40445,N_40543);
xnor U47815 (N_47815,N_44221,N_43410);
nand U47816 (N_47816,N_42018,N_41552);
nor U47817 (N_47817,N_44138,N_40813);
nand U47818 (N_47818,N_41998,N_42330);
nand U47819 (N_47819,N_40860,N_40135);
or U47820 (N_47820,N_44229,N_41045);
or U47821 (N_47821,N_42047,N_44333);
and U47822 (N_47822,N_41685,N_43061);
and U47823 (N_47823,N_42930,N_44887);
xnor U47824 (N_47824,N_44006,N_43635);
and U47825 (N_47825,N_44317,N_43218);
and U47826 (N_47826,N_41837,N_41691);
nor U47827 (N_47827,N_43784,N_40322);
nand U47828 (N_47828,N_44495,N_42819);
nor U47829 (N_47829,N_43196,N_44379);
or U47830 (N_47830,N_43614,N_41202);
nand U47831 (N_47831,N_42818,N_40550);
nor U47832 (N_47832,N_41561,N_43143);
or U47833 (N_47833,N_43860,N_41655);
nand U47834 (N_47834,N_44753,N_41625);
or U47835 (N_47835,N_44624,N_42696);
nor U47836 (N_47836,N_44117,N_44075);
or U47837 (N_47837,N_42597,N_41744);
nand U47838 (N_47838,N_44651,N_42030);
and U47839 (N_47839,N_42018,N_44483);
or U47840 (N_47840,N_44484,N_40216);
nand U47841 (N_47841,N_43896,N_43228);
or U47842 (N_47842,N_40359,N_44775);
nand U47843 (N_47843,N_41689,N_44410);
and U47844 (N_47844,N_44016,N_42535);
nor U47845 (N_47845,N_42014,N_42458);
or U47846 (N_47846,N_42940,N_43278);
or U47847 (N_47847,N_43390,N_42384);
nand U47848 (N_47848,N_40633,N_43005);
nand U47849 (N_47849,N_40394,N_40566);
nand U47850 (N_47850,N_42118,N_44615);
nand U47851 (N_47851,N_43066,N_42842);
nor U47852 (N_47852,N_43330,N_44665);
and U47853 (N_47853,N_40046,N_43030);
nand U47854 (N_47854,N_44171,N_44605);
nand U47855 (N_47855,N_41132,N_42502);
or U47856 (N_47856,N_42729,N_41938);
nor U47857 (N_47857,N_40035,N_44516);
and U47858 (N_47858,N_41722,N_41083);
or U47859 (N_47859,N_41312,N_42095);
or U47860 (N_47860,N_40821,N_40432);
and U47861 (N_47861,N_40344,N_43861);
nand U47862 (N_47862,N_43558,N_41354);
and U47863 (N_47863,N_42028,N_40519);
nor U47864 (N_47864,N_43976,N_44345);
or U47865 (N_47865,N_41955,N_44986);
or U47866 (N_47866,N_43698,N_44303);
or U47867 (N_47867,N_40450,N_40670);
xor U47868 (N_47868,N_42499,N_44881);
and U47869 (N_47869,N_42299,N_44872);
nand U47870 (N_47870,N_40030,N_40827);
nand U47871 (N_47871,N_42750,N_40131);
nand U47872 (N_47872,N_42134,N_41404);
and U47873 (N_47873,N_43504,N_43120);
nor U47874 (N_47874,N_40726,N_42813);
nand U47875 (N_47875,N_42518,N_43598);
nand U47876 (N_47876,N_42924,N_44807);
and U47877 (N_47877,N_43341,N_41814);
and U47878 (N_47878,N_43312,N_44575);
or U47879 (N_47879,N_41066,N_43606);
nand U47880 (N_47880,N_41943,N_40741);
nor U47881 (N_47881,N_44714,N_43532);
xnor U47882 (N_47882,N_41601,N_41613);
or U47883 (N_47883,N_41032,N_43300);
or U47884 (N_47884,N_43544,N_44504);
nor U47885 (N_47885,N_44602,N_44297);
and U47886 (N_47886,N_42601,N_43723);
or U47887 (N_47887,N_42502,N_42160);
nor U47888 (N_47888,N_44535,N_41972);
nor U47889 (N_47889,N_41556,N_41343);
xnor U47890 (N_47890,N_44139,N_42555);
nor U47891 (N_47891,N_43881,N_40959);
xor U47892 (N_47892,N_41909,N_40164);
or U47893 (N_47893,N_42661,N_41863);
nand U47894 (N_47894,N_41281,N_44751);
nand U47895 (N_47895,N_41411,N_40085);
xor U47896 (N_47896,N_43896,N_44218);
or U47897 (N_47897,N_42065,N_42949);
nand U47898 (N_47898,N_41715,N_44168);
or U47899 (N_47899,N_40026,N_44933);
nand U47900 (N_47900,N_41827,N_43974);
nor U47901 (N_47901,N_41354,N_43848);
nand U47902 (N_47902,N_42883,N_41411);
nor U47903 (N_47903,N_41638,N_40475);
and U47904 (N_47904,N_43338,N_44432);
nand U47905 (N_47905,N_43340,N_44650);
nand U47906 (N_47906,N_44711,N_44372);
or U47907 (N_47907,N_43953,N_41658);
nand U47908 (N_47908,N_42681,N_43356);
or U47909 (N_47909,N_42595,N_43828);
nand U47910 (N_47910,N_44720,N_41738);
nand U47911 (N_47911,N_42249,N_44968);
nor U47912 (N_47912,N_41646,N_43076);
nor U47913 (N_47913,N_43999,N_44995);
and U47914 (N_47914,N_42000,N_40566);
nor U47915 (N_47915,N_43997,N_43517);
and U47916 (N_47916,N_44908,N_40680);
or U47917 (N_47917,N_40870,N_41950);
nor U47918 (N_47918,N_43161,N_42569);
xor U47919 (N_47919,N_41368,N_42738);
or U47920 (N_47920,N_44271,N_40358);
or U47921 (N_47921,N_42547,N_42364);
or U47922 (N_47922,N_42387,N_40156);
xnor U47923 (N_47923,N_44980,N_43181);
and U47924 (N_47924,N_40397,N_44659);
or U47925 (N_47925,N_43193,N_42767);
xor U47926 (N_47926,N_43719,N_43691);
and U47927 (N_47927,N_42996,N_44038);
nor U47928 (N_47928,N_43114,N_42567);
nor U47929 (N_47929,N_44175,N_41053);
and U47930 (N_47930,N_41321,N_42194);
xnor U47931 (N_47931,N_41879,N_44261);
nand U47932 (N_47932,N_44608,N_43381);
or U47933 (N_47933,N_41680,N_40747);
and U47934 (N_47934,N_42618,N_44840);
and U47935 (N_47935,N_42240,N_40388);
or U47936 (N_47936,N_42183,N_40456);
xnor U47937 (N_47937,N_44015,N_41935);
and U47938 (N_47938,N_43876,N_40826);
nand U47939 (N_47939,N_43929,N_41334);
nand U47940 (N_47940,N_44495,N_41283);
nand U47941 (N_47941,N_43237,N_44265);
nor U47942 (N_47942,N_43099,N_43651);
or U47943 (N_47943,N_40638,N_41857);
and U47944 (N_47944,N_44256,N_40395);
or U47945 (N_47945,N_44215,N_40917);
nand U47946 (N_47946,N_44418,N_44542);
nor U47947 (N_47947,N_40590,N_42744);
and U47948 (N_47948,N_41881,N_41796);
and U47949 (N_47949,N_40040,N_44821);
nand U47950 (N_47950,N_40968,N_40009);
and U47951 (N_47951,N_43149,N_43198);
nand U47952 (N_47952,N_40496,N_41685);
nand U47953 (N_47953,N_44430,N_41757);
nor U47954 (N_47954,N_40232,N_44838);
nand U47955 (N_47955,N_43490,N_42158);
nand U47956 (N_47956,N_40806,N_42962);
nand U47957 (N_47957,N_44928,N_42546);
and U47958 (N_47958,N_40361,N_41364);
nor U47959 (N_47959,N_40318,N_40291);
xnor U47960 (N_47960,N_44499,N_42568);
nor U47961 (N_47961,N_44546,N_41962);
nand U47962 (N_47962,N_41935,N_44312);
nand U47963 (N_47963,N_40517,N_41376);
nand U47964 (N_47964,N_41799,N_44249);
xnor U47965 (N_47965,N_42823,N_41594);
xnor U47966 (N_47966,N_42101,N_43182);
and U47967 (N_47967,N_42756,N_44677);
nand U47968 (N_47968,N_41079,N_44234);
nand U47969 (N_47969,N_41639,N_42341);
nor U47970 (N_47970,N_42678,N_43929);
nor U47971 (N_47971,N_43169,N_41775);
or U47972 (N_47972,N_43065,N_43349);
and U47973 (N_47973,N_42066,N_43795);
nand U47974 (N_47974,N_44237,N_42164);
nand U47975 (N_47975,N_43721,N_41899);
and U47976 (N_47976,N_43190,N_40158);
nor U47977 (N_47977,N_42942,N_44761);
or U47978 (N_47978,N_43064,N_42494);
or U47979 (N_47979,N_42139,N_41658);
and U47980 (N_47980,N_42530,N_42232);
and U47981 (N_47981,N_42826,N_42249);
nor U47982 (N_47982,N_40119,N_40169);
and U47983 (N_47983,N_42963,N_40763);
xor U47984 (N_47984,N_43629,N_41320);
or U47985 (N_47985,N_40969,N_44100);
or U47986 (N_47986,N_43648,N_40555);
nor U47987 (N_47987,N_44649,N_42029);
nand U47988 (N_47988,N_42865,N_42580);
and U47989 (N_47989,N_44618,N_41825);
nor U47990 (N_47990,N_42397,N_42184);
or U47991 (N_47991,N_44422,N_43601);
nor U47992 (N_47992,N_40221,N_42025);
nand U47993 (N_47993,N_44260,N_43461);
and U47994 (N_47994,N_42652,N_44361);
nand U47995 (N_47995,N_40683,N_42254);
or U47996 (N_47996,N_42436,N_43226);
and U47997 (N_47997,N_43872,N_42846);
nor U47998 (N_47998,N_43141,N_44938);
nor U47999 (N_47999,N_43936,N_41689);
or U48000 (N_48000,N_43904,N_40751);
nor U48001 (N_48001,N_40679,N_44898);
or U48002 (N_48002,N_42532,N_44607);
nor U48003 (N_48003,N_40785,N_43096);
and U48004 (N_48004,N_42827,N_40075);
xor U48005 (N_48005,N_40424,N_42364);
and U48006 (N_48006,N_42943,N_43197);
nand U48007 (N_48007,N_42546,N_40764);
nand U48008 (N_48008,N_42788,N_42612);
nand U48009 (N_48009,N_43194,N_44614);
xnor U48010 (N_48010,N_41681,N_41964);
xnor U48011 (N_48011,N_44416,N_42071);
nor U48012 (N_48012,N_43755,N_42219);
or U48013 (N_48013,N_43517,N_44073);
nor U48014 (N_48014,N_44434,N_44571);
nand U48015 (N_48015,N_40193,N_40397);
nor U48016 (N_48016,N_40035,N_42916);
and U48017 (N_48017,N_43569,N_40601);
or U48018 (N_48018,N_41516,N_42939);
xnor U48019 (N_48019,N_41972,N_44908);
nor U48020 (N_48020,N_40597,N_41617);
nand U48021 (N_48021,N_44947,N_41497);
nor U48022 (N_48022,N_44128,N_43432);
or U48023 (N_48023,N_44466,N_40622);
or U48024 (N_48024,N_41298,N_42895);
nand U48025 (N_48025,N_41398,N_44497);
and U48026 (N_48026,N_44601,N_40524);
and U48027 (N_48027,N_40611,N_41807);
and U48028 (N_48028,N_42343,N_42365);
and U48029 (N_48029,N_41505,N_41606);
nor U48030 (N_48030,N_44638,N_41833);
or U48031 (N_48031,N_44989,N_43157);
and U48032 (N_48032,N_43040,N_40064);
and U48033 (N_48033,N_43641,N_42323);
xnor U48034 (N_48034,N_41625,N_42203);
and U48035 (N_48035,N_43754,N_41377);
and U48036 (N_48036,N_44644,N_42186);
xor U48037 (N_48037,N_40904,N_42746);
or U48038 (N_48038,N_42010,N_43537);
nand U48039 (N_48039,N_41286,N_42239);
nor U48040 (N_48040,N_44558,N_44922);
nor U48041 (N_48041,N_42033,N_42196);
and U48042 (N_48042,N_40023,N_40303);
or U48043 (N_48043,N_41032,N_41530);
or U48044 (N_48044,N_40355,N_41890);
nand U48045 (N_48045,N_42367,N_43418);
xnor U48046 (N_48046,N_44460,N_43528);
or U48047 (N_48047,N_43431,N_42999);
xnor U48048 (N_48048,N_44863,N_40767);
and U48049 (N_48049,N_44871,N_41699);
nor U48050 (N_48050,N_44804,N_44755);
nor U48051 (N_48051,N_44581,N_40726);
or U48052 (N_48052,N_44789,N_41229);
and U48053 (N_48053,N_41829,N_40149);
nand U48054 (N_48054,N_41546,N_41796);
and U48055 (N_48055,N_44924,N_40247);
or U48056 (N_48056,N_40826,N_43614);
and U48057 (N_48057,N_44971,N_41581);
or U48058 (N_48058,N_41748,N_41996);
nand U48059 (N_48059,N_44151,N_42664);
and U48060 (N_48060,N_42562,N_43788);
nor U48061 (N_48061,N_44860,N_43120);
or U48062 (N_48062,N_42203,N_41363);
and U48063 (N_48063,N_41674,N_40403);
and U48064 (N_48064,N_40489,N_43263);
nand U48065 (N_48065,N_42746,N_43825);
and U48066 (N_48066,N_44580,N_44753);
nor U48067 (N_48067,N_40658,N_43093);
nor U48068 (N_48068,N_43889,N_44054);
and U48069 (N_48069,N_43380,N_42109);
or U48070 (N_48070,N_40309,N_43585);
nor U48071 (N_48071,N_43515,N_42520);
and U48072 (N_48072,N_43782,N_44655);
nor U48073 (N_48073,N_44766,N_44152);
nor U48074 (N_48074,N_41755,N_42570);
or U48075 (N_48075,N_43422,N_43122);
and U48076 (N_48076,N_43440,N_43940);
nand U48077 (N_48077,N_41526,N_40572);
nand U48078 (N_48078,N_44675,N_42516);
nand U48079 (N_48079,N_42610,N_44099);
or U48080 (N_48080,N_44165,N_44032);
or U48081 (N_48081,N_44902,N_40737);
and U48082 (N_48082,N_43447,N_41638);
or U48083 (N_48083,N_44900,N_40394);
and U48084 (N_48084,N_40099,N_44892);
and U48085 (N_48085,N_44593,N_40124);
xnor U48086 (N_48086,N_40161,N_43010);
xor U48087 (N_48087,N_42189,N_43349);
and U48088 (N_48088,N_41210,N_43787);
and U48089 (N_48089,N_42527,N_44756);
or U48090 (N_48090,N_42529,N_41290);
and U48091 (N_48091,N_40367,N_40071);
nor U48092 (N_48092,N_42738,N_42869);
and U48093 (N_48093,N_44292,N_44836);
nor U48094 (N_48094,N_40990,N_42873);
xnor U48095 (N_48095,N_44036,N_40173);
xnor U48096 (N_48096,N_41371,N_43802);
nand U48097 (N_48097,N_43054,N_40418);
nand U48098 (N_48098,N_44633,N_43183);
nand U48099 (N_48099,N_42200,N_43338);
nor U48100 (N_48100,N_41958,N_44314);
nor U48101 (N_48101,N_41856,N_42793);
nand U48102 (N_48102,N_41158,N_41096);
nor U48103 (N_48103,N_42373,N_42062);
nand U48104 (N_48104,N_44849,N_41933);
nand U48105 (N_48105,N_42588,N_40644);
or U48106 (N_48106,N_44831,N_40554);
nand U48107 (N_48107,N_42758,N_44862);
and U48108 (N_48108,N_42855,N_43772);
and U48109 (N_48109,N_42910,N_43452);
xor U48110 (N_48110,N_43344,N_44798);
nand U48111 (N_48111,N_40459,N_41813);
nor U48112 (N_48112,N_44863,N_43708);
or U48113 (N_48113,N_43194,N_42172);
and U48114 (N_48114,N_43983,N_41930);
and U48115 (N_48115,N_41562,N_43060);
and U48116 (N_48116,N_43166,N_42256);
nor U48117 (N_48117,N_40972,N_41379);
nor U48118 (N_48118,N_40085,N_43349);
and U48119 (N_48119,N_41528,N_41516);
nor U48120 (N_48120,N_44961,N_42978);
or U48121 (N_48121,N_42723,N_41988);
and U48122 (N_48122,N_40970,N_40654);
and U48123 (N_48123,N_41556,N_40397);
or U48124 (N_48124,N_44432,N_40516);
and U48125 (N_48125,N_43829,N_40299);
or U48126 (N_48126,N_44550,N_42814);
and U48127 (N_48127,N_44023,N_42550);
xnor U48128 (N_48128,N_42484,N_43619);
nor U48129 (N_48129,N_40537,N_43894);
or U48130 (N_48130,N_40129,N_44606);
nand U48131 (N_48131,N_43834,N_40680);
or U48132 (N_48132,N_43222,N_43049);
or U48133 (N_48133,N_41154,N_44189);
or U48134 (N_48134,N_42585,N_42861);
and U48135 (N_48135,N_42389,N_44439);
or U48136 (N_48136,N_43913,N_42883);
nor U48137 (N_48137,N_44562,N_43435);
nor U48138 (N_48138,N_40755,N_44597);
and U48139 (N_48139,N_40350,N_40164);
nor U48140 (N_48140,N_41028,N_43139);
or U48141 (N_48141,N_41697,N_43300);
and U48142 (N_48142,N_44680,N_42389);
or U48143 (N_48143,N_42050,N_40064);
or U48144 (N_48144,N_40437,N_43218);
or U48145 (N_48145,N_43189,N_42455);
nor U48146 (N_48146,N_42410,N_43733);
nand U48147 (N_48147,N_43960,N_44814);
and U48148 (N_48148,N_42361,N_43525);
or U48149 (N_48149,N_44669,N_40584);
nor U48150 (N_48150,N_44897,N_43779);
nor U48151 (N_48151,N_40391,N_40133);
xor U48152 (N_48152,N_40654,N_43743);
and U48153 (N_48153,N_43652,N_40332);
or U48154 (N_48154,N_41074,N_41188);
xor U48155 (N_48155,N_43452,N_43651);
nand U48156 (N_48156,N_41909,N_42020);
xor U48157 (N_48157,N_42329,N_41130);
nand U48158 (N_48158,N_44360,N_44406);
and U48159 (N_48159,N_41839,N_41560);
and U48160 (N_48160,N_41882,N_40371);
nor U48161 (N_48161,N_41630,N_43104);
and U48162 (N_48162,N_44861,N_44089);
nand U48163 (N_48163,N_40912,N_40066);
xor U48164 (N_48164,N_40752,N_42790);
or U48165 (N_48165,N_40707,N_42717);
and U48166 (N_48166,N_43401,N_42959);
nor U48167 (N_48167,N_44355,N_41715);
and U48168 (N_48168,N_43393,N_40292);
and U48169 (N_48169,N_42372,N_40730);
or U48170 (N_48170,N_41462,N_43652);
nand U48171 (N_48171,N_40019,N_43196);
nand U48172 (N_48172,N_41620,N_43249);
xor U48173 (N_48173,N_40789,N_41075);
and U48174 (N_48174,N_40271,N_42250);
nor U48175 (N_48175,N_42493,N_42836);
and U48176 (N_48176,N_42805,N_41321);
xor U48177 (N_48177,N_41172,N_43007);
or U48178 (N_48178,N_44678,N_43956);
or U48179 (N_48179,N_43269,N_44153);
nor U48180 (N_48180,N_43556,N_44582);
nand U48181 (N_48181,N_40529,N_41486);
xor U48182 (N_48182,N_43123,N_44672);
nor U48183 (N_48183,N_41096,N_40815);
nor U48184 (N_48184,N_44777,N_44178);
xor U48185 (N_48185,N_42173,N_43379);
and U48186 (N_48186,N_43842,N_44916);
or U48187 (N_48187,N_41095,N_40237);
and U48188 (N_48188,N_41485,N_42958);
and U48189 (N_48189,N_44857,N_40298);
and U48190 (N_48190,N_44361,N_42623);
and U48191 (N_48191,N_44340,N_40536);
nor U48192 (N_48192,N_42197,N_41698);
nor U48193 (N_48193,N_40099,N_42612);
nor U48194 (N_48194,N_43514,N_41435);
nand U48195 (N_48195,N_44118,N_40163);
nand U48196 (N_48196,N_40356,N_42489);
and U48197 (N_48197,N_41942,N_42688);
and U48198 (N_48198,N_40659,N_44616);
nor U48199 (N_48199,N_44134,N_42971);
nand U48200 (N_48200,N_44431,N_42897);
nand U48201 (N_48201,N_43551,N_42596);
nor U48202 (N_48202,N_41200,N_44352);
or U48203 (N_48203,N_43813,N_42949);
or U48204 (N_48204,N_44887,N_42979);
and U48205 (N_48205,N_42432,N_40926);
or U48206 (N_48206,N_44961,N_44009);
or U48207 (N_48207,N_43681,N_41278);
and U48208 (N_48208,N_44587,N_42009);
nand U48209 (N_48209,N_41093,N_44924);
and U48210 (N_48210,N_40689,N_42601);
nand U48211 (N_48211,N_40584,N_44394);
or U48212 (N_48212,N_41085,N_42366);
or U48213 (N_48213,N_44162,N_41237);
xnor U48214 (N_48214,N_40087,N_43210);
nand U48215 (N_48215,N_42514,N_44873);
nor U48216 (N_48216,N_42394,N_44679);
nor U48217 (N_48217,N_43650,N_40313);
or U48218 (N_48218,N_43642,N_43436);
nor U48219 (N_48219,N_43829,N_44804);
and U48220 (N_48220,N_43941,N_42008);
nor U48221 (N_48221,N_43484,N_44303);
nor U48222 (N_48222,N_44073,N_42776);
nor U48223 (N_48223,N_41839,N_41902);
or U48224 (N_48224,N_42047,N_40330);
nand U48225 (N_48225,N_43924,N_43952);
nand U48226 (N_48226,N_40202,N_44574);
or U48227 (N_48227,N_44235,N_41118);
nand U48228 (N_48228,N_42249,N_42638);
nand U48229 (N_48229,N_44455,N_43748);
or U48230 (N_48230,N_44257,N_41771);
or U48231 (N_48231,N_44887,N_41445);
nand U48232 (N_48232,N_42383,N_44505);
and U48233 (N_48233,N_43737,N_44564);
and U48234 (N_48234,N_41161,N_43606);
xor U48235 (N_48235,N_40063,N_41289);
xnor U48236 (N_48236,N_40018,N_44792);
nand U48237 (N_48237,N_44860,N_44144);
and U48238 (N_48238,N_41818,N_41608);
nor U48239 (N_48239,N_44359,N_41457);
xnor U48240 (N_48240,N_44968,N_41213);
nor U48241 (N_48241,N_41728,N_44339);
nand U48242 (N_48242,N_42711,N_40223);
nand U48243 (N_48243,N_41065,N_43128);
or U48244 (N_48244,N_41291,N_41719);
and U48245 (N_48245,N_40350,N_42515);
and U48246 (N_48246,N_44782,N_44544);
or U48247 (N_48247,N_40103,N_41560);
and U48248 (N_48248,N_44188,N_41114);
or U48249 (N_48249,N_42581,N_40842);
and U48250 (N_48250,N_42498,N_42137);
nand U48251 (N_48251,N_40181,N_40517);
or U48252 (N_48252,N_41903,N_42905);
nand U48253 (N_48253,N_42032,N_40637);
nor U48254 (N_48254,N_42826,N_41696);
and U48255 (N_48255,N_43828,N_42621);
nand U48256 (N_48256,N_41673,N_40556);
xor U48257 (N_48257,N_41010,N_44612);
nand U48258 (N_48258,N_41053,N_40482);
nor U48259 (N_48259,N_42923,N_41440);
nand U48260 (N_48260,N_44506,N_40663);
nand U48261 (N_48261,N_44771,N_43939);
or U48262 (N_48262,N_44668,N_42466);
or U48263 (N_48263,N_40779,N_43039);
nor U48264 (N_48264,N_40137,N_42633);
and U48265 (N_48265,N_43840,N_44261);
and U48266 (N_48266,N_40606,N_43082);
and U48267 (N_48267,N_43045,N_43238);
or U48268 (N_48268,N_40929,N_44541);
and U48269 (N_48269,N_42360,N_43874);
nand U48270 (N_48270,N_40200,N_41127);
and U48271 (N_48271,N_41839,N_44618);
or U48272 (N_48272,N_40099,N_42836);
nor U48273 (N_48273,N_44437,N_41414);
nand U48274 (N_48274,N_43316,N_41159);
and U48275 (N_48275,N_42811,N_40333);
nor U48276 (N_48276,N_43963,N_43097);
or U48277 (N_48277,N_42355,N_43593);
and U48278 (N_48278,N_44737,N_42031);
nor U48279 (N_48279,N_42982,N_41095);
xnor U48280 (N_48280,N_44032,N_42615);
nor U48281 (N_48281,N_44313,N_42858);
or U48282 (N_48282,N_43581,N_40839);
xnor U48283 (N_48283,N_40068,N_40035);
nor U48284 (N_48284,N_40265,N_42841);
and U48285 (N_48285,N_42169,N_41694);
nor U48286 (N_48286,N_40552,N_44360);
nand U48287 (N_48287,N_43630,N_44377);
or U48288 (N_48288,N_40620,N_40314);
nand U48289 (N_48289,N_44143,N_40497);
nor U48290 (N_48290,N_41329,N_40435);
or U48291 (N_48291,N_43636,N_40029);
or U48292 (N_48292,N_44118,N_41537);
nor U48293 (N_48293,N_44489,N_42521);
nand U48294 (N_48294,N_40628,N_42554);
or U48295 (N_48295,N_43471,N_41493);
nand U48296 (N_48296,N_41064,N_43135);
or U48297 (N_48297,N_42056,N_41776);
or U48298 (N_48298,N_43430,N_44271);
and U48299 (N_48299,N_42157,N_40297);
nand U48300 (N_48300,N_43887,N_42640);
or U48301 (N_48301,N_44174,N_41543);
and U48302 (N_48302,N_43056,N_40798);
and U48303 (N_48303,N_44308,N_41430);
and U48304 (N_48304,N_42816,N_44563);
and U48305 (N_48305,N_43987,N_41855);
nor U48306 (N_48306,N_44389,N_40322);
nor U48307 (N_48307,N_40616,N_43669);
or U48308 (N_48308,N_44806,N_43273);
and U48309 (N_48309,N_42536,N_43114);
and U48310 (N_48310,N_43914,N_41332);
and U48311 (N_48311,N_43117,N_43603);
nor U48312 (N_48312,N_41331,N_40414);
xor U48313 (N_48313,N_42842,N_41124);
and U48314 (N_48314,N_40301,N_42689);
nor U48315 (N_48315,N_42690,N_44818);
or U48316 (N_48316,N_44375,N_40990);
or U48317 (N_48317,N_43559,N_44062);
or U48318 (N_48318,N_40257,N_44599);
nor U48319 (N_48319,N_42388,N_40650);
nand U48320 (N_48320,N_41743,N_40929);
nor U48321 (N_48321,N_40529,N_40921);
nor U48322 (N_48322,N_43399,N_44552);
nor U48323 (N_48323,N_40083,N_44200);
nand U48324 (N_48324,N_43974,N_41548);
nand U48325 (N_48325,N_44540,N_42205);
nand U48326 (N_48326,N_44674,N_41015);
nor U48327 (N_48327,N_43405,N_42579);
xnor U48328 (N_48328,N_41308,N_41289);
nor U48329 (N_48329,N_40368,N_41905);
or U48330 (N_48330,N_42295,N_40953);
or U48331 (N_48331,N_43406,N_43403);
and U48332 (N_48332,N_40762,N_41638);
and U48333 (N_48333,N_43604,N_40765);
and U48334 (N_48334,N_41355,N_42233);
and U48335 (N_48335,N_43720,N_43420);
and U48336 (N_48336,N_41576,N_42248);
and U48337 (N_48337,N_43410,N_41945);
xnor U48338 (N_48338,N_42699,N_42231);
and U48339 (N_48339,N_41292,N_40496);
nand U48340 (N_48340,N_43909,N_42401);
and U48341 (N_48341,N_41083,N_42528);
or U48342 (N_48342,N_40958,N_42451);
nor U48343 (N_48343,N_43576,N_44407);
nor U48344 (N_48344,N_44698,N_44973);
nand U48345 (N_48345,N_44618,N_44040);
nor U48346 (N_48346,N_41977,N_43936);
nor U48347 (N_48347,N_40112,N_41741);
nand U48348 (N_48348,N_41898,N_41618);
nand U48349 (N_48349,N_41552,N_43104);
nor U48350 (N_48350,N_41537,N_44323);
and U48351 (N_48351,N_40049,N_43866);
nand U48352 (N_48352,N_44335,N_40069);
or U48353 (N_48353,N_42049,N_43753);
and U48354 (N_48354,N_40651,N_40881);
xor U48355 (N_48355,N_43134,N_41074);
or U48356 (N_48356,N_41394,N_42519);
and U48357 (N_48357,N_41813,N_41805);
nor U48358 (N_48358,N_40383,N_43718);
and U48359 (N_48359,N_43462,N_40565);
and U48360 (N_48360,N_40250,N_40213);
xnor U48361 (N_48361,N_43507,N_42256);
or U48362 (N_48362,N_40736,N_43142);
nand U48363 (N_48363,N_44502,N_40056);
nand U48364 (N_48364,N_43574,N_44246);
and U48365 (N_48365,N_41278,N_41581);
and U48366 (N_48366,N_43628,N_44802);
or U48367 (N_48367,N_41473,N_43184);
and U48368 (N_48368,N_42307,N_42599);
nor U48369 (N_48369,N_42098,N_41651);
and U48370 (N_48370,N_43725,N_43233);
and U48371 (N_48371,N_41497,N_43145);
or U48372 (N_48372,N_43259,N_43340);
and U48373 (N_48373,N_41274,N_42010);
or U48374 (N_48374,N_42059,N_41272);
or U48375 (N_48375,N_40910,N_40528);
or U48376 (N_48376,N_40936,N_41668);
nor U48377 (N_48377,N_41707,N_42513);
and U48378 (N_48378,N_43162,N_40726);
nor U48379 (N_48379,N_43726,N_40982);
nor U48380 (N_48380,N_41399,N_41515);
nand U48381 (N_48381,N_42186,N_42999);
or U48382 (N_48382,N_44542,N_40872);
or U48383 (N_48383,N_42354,N_40399);
nand U48384 (N_48384,N_42976,N_41961);
or U48385 (N_48385,N_40740,N_43064);
nor U48386 (N_48386,N_43803,N_44507);
nand U48387 (N_48387,N_42252,N_41125);
xnor U48388 (N_48388,N_43596,N_40287);
nor U48389 (N_48389,N_40140,N_42647);
nand U48390 (N_48390,N_41781,N_43821);
nand U48391 (N_48391,N_44693,N_41648);
xnor U48392 (N_48392,N_44016,N_40567);
nand U48393 (N_48393,N_40224,N_44622);
nand U48394 (N_48394,N_40940,N_44893);
nor U48395 (N_48395,N_44491,N_42195);
nor U48396 (N_48396,N_43506,N_40845);
nor U48397 (N_48397,N_40222,N_42500);
nor U48398 (N_48398,N_44371,N_44248);
nand U48399 (N_48399,N_41678,N_41399);
xor U48400 (N_48400,N_43674,N_44951);
and U48401 (N_48401,N_44874,N_44200);
nand U48402 (N_48402,N_42330,N_43772);
nand U48403 (N_48403,N_44792,N_40436);
nor U48404 (N_48404,N_44475,N_43508);
and U48405 (N_48405,N_44308,N_42421);
nand U48406 (N_48406,N_42239,N_40727);
nand U48407 (N_48407,N_41307,N_43250);
nand U48408 (N_48408,N_44990,N_40293);
nand U48409 (N_48409,N_43504,N_43836);
nor U48410 (N_48410,N_43969,N_44544);
nand U48411 (N_48411,N_40943,N_42658);
nor U48412 (N_48412,N_43796,N_44453);
nand U48413 (N_48413,N_40898,N_41828);
and U48414 (N_48414,N_43172,N_40036);
or U48415 (N_48415,N_42431,N_44231);
or U48416 (N_48416,N_43688,N_43627);
or U48417 (N_48417,N_44406,N_42232);
and U48418 (N_48418,N_42050,N_44533);
or U48419 (N_48419,N_40426,N_43621);
nand U48420 (N_48420,N_40371,N_40370);
or U48421 (N_48421,N_43266,N_43757);
nand U48422 (N_48422,N_40434,N_44119);
nor U48423 (N_48423,N_40984,N_44374);
and U48424 (N_48424,N_40000,N_42421);
or U48425 (N_48425,N_41008,N_43924);
and U48426 (N_48426,N_43339,N_42271);
nand U48427 (N_48427,N_43651,N_44641);
nand U48428 (N_48428,N_43016,N_41773);
and U48429 (N_48429,N_41137,N_42017);
nor U48430 (N_48430,N_40997,N_40780);
nand U48431 (N_48431,N_40533,N_41650);
nand U48432 (N_48432,N_41365,N_42533);
or U48433 (N_48433,N_44217,N_44305);
or U48434 (N_48434,N_41831,N_43765);
nand U48435 (N_48435,N_41870,N_41005);
nor U48436 (N_48436,N_41685,N_43209);
nand U48437 (N_48437,N_41081,N_42292);
and U48438 (N_48438,N_41513,N_43019);
xnor U48439 (N_48439,N_44485,N_40450);
nand U48440 (N_48440,N_43147,N_43915);
and U48441 (N_48441,N_43277,N_40815);
nand U48442 (N_48442,N_41470,N_42476);
nor U48443 (N_48443,N_44740,N_43296);
and U48444 (N_48444,N_41862,N_43944);
nand U48445 (N_48445,N_43558,N_40145);
or U48446 (N_48446,N_40587,N_43734);
xnor U48447 (N_48447,N_40013,N_44754);
nand U48448 (N_48448,N_43321,N_41511);
nand U48449 (N_48449,N_40557,N_43235);
and U48450 (N_48450,N_42704,N_41718);
and U48451 (N_48451,N_41736,N_41535);
and U48452 (N_48452,N_41762,N_41547);
nor U48453 (N_48453,N_42382,N_40211);
or U48454 (N_48454,N_40133,N_44775);
nor U48455 (N_48455,N_41551,N_40796);
or U48456 (N_48456,N_41604,N_43810);
or U48457 (N_48457,N_42488,N_42638);
or U48458 (N_48458,N_43470,N_40914);
xnor U48459 (N_48459,N_41830,N_44423);
nand U48460 (N_48460,N_40949,N_42331);
and U48461 (N_48461,N_42010,N_43123);
nand U48462 (N_48462,N_42027,N_40882);
or U48463 (N_48463,N_43159,N_44081);
or U48464 (N_48464,N_40698,N_44210);
and U48465 (N_48465,N_40781,N_43616);
xnor U48466 (N_48466,N_42455,N_43128);
or U48467 (N_48467,N_44852,N_42487);
nand U48468 (N_48468,N_40656,N_41650);
and U48469 (N_48469,N_44345,N_41591);
or U48470 (N_48470,N_41510,N_40119);
nand U48471 (N_48471,N_42414,N_41187);
nand U48472 (N_48472,N_42087,N_43862);
nor U48473 (N_48473,N_41440,N_42422);
or U48474 (N_48474,N_43676,N_44948);
or U48475 (N_48475,N_40499,N_41447);
nand U48476 (N_48476,N_41578,N_41969);
xor U48477 (N_48477,N_41934,N_40413);
and U48478 (N_48478,N_41853,N_44300);
and U48479 (N_48479,N_41331,N_43407);
and U48480 (N_48480,N_41955,N_41213);
nor U48481 (N_48481,N_42342,N_41312);
nor U48482 (N_48482,N_42651,N_40008);
nand U48483 (N_48483,N_44046,N_40652);
nand U48484 (N_48484,N_42662,N_44494);
nor U48485 (N_48485,N_40996,N_43848);
nand U48486 (N_48486,N_44916,N_43105);
xnor U48487 (N_48487,N_42475,N_43699);
nand U48488 (N_48488,N_44865,N_41891);
nand U48489 (N_48489,N_42742,N_42623);
nand U48490 (N_48490,N_41606,N_42473);
and U48491 (N_48491,N_43564,N_44750);
and U48492 (N_48492,N_40283,N_44634);
and U48493 (N_48493,N_40565,N_43004);
or U48494 (N_48494,N_40016,N_43900);
nand U48495 (N_48495,N_43849,N_43926);
nor U48496 (N_48496,N_40488,N_43489);
xor U48497 (N_48497,N_40716,N_42872);
nor U48498 (N_48498,N_43778,N_43797);
and U48499 (N_48499,N_43367,N_43677);
and U48500 (N_48500,N_43993,N_42389);
or U48501 (N_48501,N_42727,N_44732);
nor U48502 (N_48502,N_41170,N_40391);
nor U48503 (N_48503,N_41442,N_42036);
xor U48504 (N_48504,N_43639,N_41865);
nor U48505 (N_48505,N_41454,N_44793);
and U48506 (N_48506,N_42976,N_40512);
or U48507 (N_48507,N_42587,N_44025);
nor U48508 (N_48508,N_40459,N_43486);
nor U48509 (N_48509,N_44091,N_41226);
nand U48510 (N_48510,N_44975,N_42681);
xnor U48511 (N_48511,N_44473,N_41142);
nand U48512 (N_48512,N_41513,N_44973);
or U48513 (N_48513,N_40873,N_40052);
or U48514 (N_48514,N_43060,N_42956);
or U48515 (N_48515,N_40560,N_42310);
or U48516 (N_48516,N_43941,N_43504);
and U48517 (N_48517,N_40062,N_42124);
nor U48518 (N_48518,N_40496,N_41998);
nor U48519 (N_48519,N_42583,N_40915);
or U48520 (N_48520,N_42198,N_41895);
nor U48521 (N_48521,N_44040,N_43958);
nand U48522 (N_48522,N_43997,N_43220);
nand U48523 (N_48523,N_41622,N_42445);
and U48524 (N_48524,N_40089,N_41475);
or U48525 (N_48525,N_41198,N_41296);
nand U48526 (N_48526,N_42819,N_42460);
nor U48527 (N_48527,N_41604,N_43374);
or U48528 (N_48528,N_41654,N_40788);
xnor U48529 (N_48529,N_42466,N_43711);
xor U48530 (N_48530,N_42119,N_40483);
and U48531 (N_48531,N_44193,N_44307);
and U48532 (N_48532,N_41301,N_43354);
nor U48533 (N_48533,N_41526,N_42302);
xnor U48534 (N_48534,N_44474,N_41280);
nand U48535 (N_48535,N_43982,N_44302);
nor U48536 (N_48536,N_44905,N_43031);
nand U48537 (N_48537,N_40250,N_41132);
nand U48538 (N_48538,N_43851,N_44757);
and U48539 (N_48539,N_40849,N_41003);
nor U48540 (N_48540,N_41484,N_40200);
nor U48541 (N_48541,N_40049,N_43798);
nor U48542 (N_48542,N_43344,N_42968);
or U48543 (N_48543,N_42586,N_41573);
nor U48544 (N_48544,N_40172,N_43574);
nand U48545 (N_48545,N_41709,N_40272);
and U48546 (N_48546,N_44242,N_44057);
nor U48547 (N_48547,N_42161,N_40555);
nor U48548 (N_48548,N_41479,N_42743);
nor U48549 (N_48549,N_43894,N_44442);
or U48550 (N_48550,N_42131,N_40767);
xor U48551 (N_48551,N_43138,N_43024);
nor U48552 (N_48552,N_40818,N_41190);
and U48553 (N_48553,N_44795,N_40287);
nand U48554 (N_48554,N_44065,N_43965);
nor U48555 (N_48555,N_44243,N_43918);
and U48556 (N_48556,N_41674,N_40264);
nand U48557 (N_48557,N_42030,N_41659);
nand U48558 (N_48558,N_41404,N_40191);
nor U48559 (N_48559,N_44282,N_43185);
nand U48560 (N_48560,N_43549,N_44251);
nor U48561 (N_48561,N_43791,N_40533);
nor U48562 (N_48562,N_42735,N_42085);
nor U48563 (N_48563,N_42121,N_42620);
or U48564 (N_48564,N_44037,N_43405);
and U48565 (N_48565,N_44808,N_44298);
nor U48566 (N_48566,N_40440,N_42235);
xor U48567 (N_48567,N_44571,N_44257);
or U48568 (N_48568,N_42465,N_41975);
and U48569 (N_48569,N_41940,N_44932);
nand U48570 (N_48570,N_41426,N_44234);
nand U48571 (N_48571,N_40739,N_43291);
nand U48572 (N_48572,N_40981,N_42564);
and U48573 (N_48573,N_41241,N_43283);
nor U48574 (N_48574,N_43943,N_42849);
or U48575 (N_48575,N_43277,N_40892);
nor U48576 (N_48576,N_42691,N_43225);
and U48577 (N_48577,N_44927,N_40424);
and U48578 (N_48578,N_41191,N_41046);
nor U48579 (N_48579,N_43000,N_43645);
or U48580 (N_48580,N_43226,N_44239);
or U48581 (N_48581,N_42812,N_44138);
nand U48582 (N_48582,N_44287,N_44810);
or U48583 (N_48583,N_41648,N_42335);
nor U48584 (N_48584,N_43492,N_44123);
xor U48585 (N_48585,N_42868,N_44498);
or U48586 (N_48586,N_44481,N_44169);
or U48587 (N_48587,N_42716,N_43500);
or U48588 (N_48588,N_42786,N_44328);
nor U48589 (N_48589,N_43328,N_41067);
or U48590 (N_48590,N_42403,N_41995);
nor U48591 (N_48591,N_41243,N_40781);
xor U48592 (N_48592,N_44667,N_43054);
nand U48593 (N_48593,N_41401,N_42619);
nand U48594 (N_48594,N_42098,N_43053);
or U48595 (N_48595,N_43020,N_40236);
or U48596 (N_48596,N_44788,N_44155);
nand U48597 (N_48597,N_43370,N_40954);
nand U48598 (N_48598,N_42732,N_43797);
xnor U48599 (N_48599,N_43822,N_40509);
and U48600 (N_48600,N_40698,N_42275);
nor U48601 (N_48601,N_43979,N_44674);
or U48602 (N_48602,N_43323,N_42457);
nor U48603 (N_48603,N_41253,N_44986);
and U48604 (N_48604,N_43640,N_41394);
and U48605 (N_48605,N_44154,N_40648);
and U48606 (N_48606,N_40299,N_41134);
and U48607 (N_48607,N_40721,N_43416);
nand U48608 (N_48608,N_42191,N_42032);
or U48609 (N_48609,N_43269,N_41678);
or U48610 (N_48610,N_43241,N_41487);
and U48611 (N_48611,N_44108,N_41571);
or U48612 (N_48612,N_40384,N_41069);
nand U48613 (N_48613,N_40930,N_43856);
and U48614 (N_48614,N_41846,N_41742);
and U48615 (N_48615,N_40425,N_44172);
and U48616 (N_48616,N_42031,N_42916);
nand U48617 (N_48617,N_40172,N_44829);
or U48618 (N_48618,N_41785,N_44431);
and U48619 (N_48619,N_44574,N_44605);
or U48620 (N_48620,N_41236,N_41523);
nand U48621 (N_48621,N_42809,N_44800);
and U48622 (N_48622,N_40854,N_41035);
nand U48623 (N_48623,N_43265,N_40122);
and U48624 (N_48624,N_44105,N_42139);
nand U48625 (N_48625,N_41443,N_42055);
or U48626 (N_48626,N_42543,N_41020);
and U48627 (N_48627,N_40401,N_44249);
or U48628 (N_48628,N_44553,N_43424);
nor U48629 (N_48629,N_43070,N_40927);
and U48630 (N_48630,N_41607,N_41944);
or U48631 (N_48631,N_44030,N_42113);
and U48632 (N_48632,N_42174,N_42000);
or U48633 (N_48633,N_43171,N_40143);
xor U48634 (N_48634,N_43025,N_43939);
nand U48635 (N_48635,N_43636,N_42353);
or U48636 (N_48636,N_41823,N_44850);
and U48637 (N_48637,N_42497,N_42864);
nor U48638 (N_48638,N_44144,N_40272);
or U48639 (N_48639,N_43691,N_42179);
nor U48640 (N_48640,N_40285,N_42244);
nand U48641 (N_48641,N_40034,N_44054);
nand U48642 (N_48642,N_40970,N_41392);
xnor U48643 (N_48643,N_44294,N_42484);
nor U48644 (N_48644,N_44877,N_44972);
nor U48645 (N_48645,N_43352,N_44517);
and U48646 (N_48646,N_44186,N_43423);
nor U48647 (N_48647,N_44265,N_42229);
or U48648 (N_48648,N_44261,N_40058);
and U48649 (N_48649,N_40741,N_43899);
and U48650 (N_48650,N_41240,N_42958);
and U48651 (N_48651,N_41867,N_40865);
and U48652 (N_48652,N_41991,N_40821);
and U48653 (N_48653,N_41316,N_44780);
and U48654 (N_48654,N_43782,N_41562);
and U48655 (N_48655,N_40647,N_44322);
nor U48656 (N_48656,N_41865,N_44738);
and U48657 (N_48657,N_43570,N_41107);
or U48658 (N_48658,N_43854,N_40465);
xor U48659 (N_48659,N_41236,N_41326);
xor U48660 (N_48660,N_42136,N_42974);
or U48661 (N_48661,N_43990,N_44891);
nand U48662 (N_48662,N_40740,N_43986);
xor U48663 (N_48663,N_44634,N_41926);
xor U48664 (N_48664,N_42658,N_40966);
or U48665 (N_48665,N_41850,N_42300);
and U48666 (N_48666,N_43456,N_41411);
nand U48667 (N_48667,N_40233,N_40329);
nor U48668 (N_48668,N_43640,N_40180);
and U48669 (N_48669,N_43349,N_40459);
nand U48670 (N_48670,N_42520,N_41896);
nand U48671 (N_48671,N_41029,N_40854);
and U48672 (N_48672,N_44961,N_44540);
xor U48673 (N_48673,N_40130,N_43681);
nor U48674 (N_48674,N_40307,N_43504);
xnor U48675 (N_48675,N_44874,N_44613);
and U48676 (N_48676,N_40663,N_41205);
nand U48677 (N_48677,N_44193,N_44180);
xnor U48678 (N_48678,N_42536,N_42102);
nand U48679 (N_48679,N_40846,N_43355);
nand U48680 (N_48680,N_41226,N_44852);
xor U48681 (N_48681,N_40911,N_43505);
nand U48682 (N_48682,N_44054,N_43920);
xnor U48683 (N_48683,N_44746,N_41766);
nand U48684 (N_48684,N_43152,N_44768);
and U48685 (N_48685,N_40683,N_41361);
nand U48686 (N_48686,N_40430,N_43716);
and U48687 (N_48687,N_41131,N_43241);
nor U48688 (N_48688,N_42364,N_40259);
nor U48689 (N_48689,N_43771,N_40519);
nor U48690 (N_48690,N_44972,N_41726);
nor U48691 (N_48691,N_40164,N_41088);
xor U48692 (N_48692,N_44227,N_40509);
or U48693 (N_48693,N_43879,N_44348);
xor U48694 (N_48694,N_41534,N_40231);
and U48695 (N_48695,N_42082,N_40698);
nand U48696 (N_48696,N_44422,N_42067);
nand U48697 (N_48697,N_40984,N_41442);
or U48698 (N_48698,N_40288,N_44935);
nand U48699 (N_48699,N_43794,N_42965);
and U48700 (N_48700,N_42674,N_43295);
nor U48701 (N_48701,N_44733,N_42970);
nor U48702 (N_48702,N_44424,N_44281);
nand U48703 (N_48703,N_42677,N_41489);
and U48704 (N_48704,N_44426,N_43729);
or U48705 (N_48705,N_41031,N_42979);
nand U48706 (N_48706,N_42103,N_44165);
nand U48707 (N_48707,N_41948,N_44182);
and U48708 (N_48708,N_41252,N_40606);
nand U48709 (N_48709,N_40679,N_44816);
and U48710 (N_48710,N_44451,N_43122);
nor U48711 (N_48711,N_44625,N_41392);
xor U48712 (N_48712,N_43954,N_43884);
xor U48713 (N_48713,N_42346,N_42935);
and U48714 (N_48714,N_44926,N_40005);
nor U48715 (N_48715,N_44028,N_43677);
xor U48716 (N_48716,N_44963,N_42654);
nand U48717 (N_48717,N_41901,N_40901);
nor U48718 (N_48718,N_43400,N_41943);
nand U48719 (N_48719,N_41865,N_43764);
or U48720 (N_48720,N_40671,N_44827);
nand U48721 (N_48721,N_42226,N_43543);
or U48722 (N_48722,N_43287,N_40337);
nand U48723 (N_48723,N_44896,N_40214);
or U48724 (N_48724,N_43719,N_43295);
or U48725 (N_48725,N_42819,N_41754);
nand U48726 (N_48726,N_42522,N_42225);
nor U48727 (N_48727,N_42014,N_44007);
xnor U48728 (N_48728,N_43448,N_40870);
or U48729 (N_48729,N_42485,N_40550);
and U48730 (N_48730,N_40004,N_41772);
xor U48731 (N_48731,N_40979,N_42772);
nand U48732 (N_48732,N_43368,N_42372);
or U48733 (N_48733,N_40417,N_40179);
and U48734 (N_48734,N_43145,N_44778);
nand U48735 (N_48735,N_40540,N_44988);
or U48736 (N_48736,N_44864,N_42421);
or U48737 (N_48737,N_43183,N_44773);
nand U48738 (N_48738,N_42026,N_40513);
and U48739 (N_48739,N_42012,N_43286);
or U48740 (N_48740,N_40911,N_40503);
nand U48741 (N_48741,N_43146,N_42665);
and U48742 (N_48742,N_41077,N_42777);
and U48743 (N_48743,N_40644,N_40960);
or U48744 (N_48744,N_44465,N_41149);
nor U48745 (N_48745,N_44141,N_42857);
nor U48746 (N_48746,N_43184,N_40836);
and U48747 (N_48747,N_43450,N_40730);
or U48748 (N_48748,N_41156,N_42608);
and U48749 (N_48749,N_42708,N_42113);
nand U48750 (N_48750,N_43097,N_41908);
nand U48751 (N_48751,N_43026,N_40712);
nand U48752 (N_48752,N_41699,N_44414);
or U48753 (N_48753,N_43509,N_41896);
or U48754 (N_48754,N_44772,N_44322);
nand U48755 (N_48755,N_43904,N_41983);
or U48756 (N_48756,N_44161,N_43103);
or U48757 (N_48757,N_41690,N_41077);
nor U48758 (N_48758,N_42666,N_40570);
nand U48759 (N_48759,N_41425,N_43735);
nor U48760 (N_48760,N_42022,N_42047);
or U48761 (N_48761,N_42307,N_44504);
and U48762 (N_48762,N_43825,N_42543);
or U48763 (N_48763,N_43928,N_44191);
or U48764 (N_48764,N_43935,N_42613);
and U48765 (N_48765,N_40738,N_40904);
nor U48766 (N_48766,N_43870,N_40149);
and U48767 (N_48767,N_44051,N_44253);
and U48768 (N_48768,N_42118,N_41528);
nand U48769 (N_48769,N_40228,N_43301);
xnor U48770 (N_48770,N_41391,N_41885);
nor U48771 (N_48771,N_41842,N_43966);
or U48772 (N_48772,N_40629,N_40111);
nand U48773 (N_48773,N_40072,N_43880);
nor U48774 (N_48774,N_44203,N_40116);
nor U48775 (N_48775,N_44222,N_43655);
nand U48776 (N_48776,N_43379,N_42094);
nand U48777 (N_48777,N_42541,N_44045);
and U48778 (N_48778,N_44081,N_40988);
and U48779 (N_48779,N_41464,N_41381);
nor U48780 (N_48780,N_40034,N_42879);
and U48781 (N_48781,N_41733,N_44819);
and U48782 (N_48782,N_40285,N_44224);
nand U48783 (N_48783,N_43070,N_41197);
nand U48784 (N_48784,N_44335,N_40861);
xor U48785 (N_48785,N_41599,N_43202);
or U48786 (N_48786,N_41988,N_42372);
nor U48787 (N_48787,N_43933,N_42686);
nor U48788 (N_48788,N_42122,N_41076);
or U48789 (N_48789,N_44791,N_44262);
nand U48790 (N_48790,N_42668,N_44371);
nor U48791 (N_48791,N_44343,N_42716);
xor U48792 (N_48792,N_43731,N_43348);
nor U48793 (N_48793,N_44796,N_40077);
nand U48794 (N_48794,N_43031,N_41606);
or U48795 (N_48795,N_44221,N_42612);
and U48796 (N_48796,N_42160,N_40960);
and U48797 (N_48797,N_43665,N_44678);
xor U48798 (N_48798,N_41686,N_44822);
nand U48799 (N_48799,N_41634,N_42209);
nor U48800 (N_48800,N_44759,N_44860);
nor U48801 (N_48801,N_42342,N_44794);
or U48802 (N_48802,N_42964,N_44290);
nor U48803 (N_48803,N_43926,N_44163);
nor U48804 (N_48804,N_43580,N_42936);
nor U48805 (N_48805,N_42493,N_44742);
or U48806 (N_48806,N_41318,N_42346);
and U48807 (N_48807,N_44072,N_44686);
or U48808 (N_48808,N_44134,N_41147);
nor U48809 (N_48809,N_43952,N_42055);
xor U48810 (N_48810,N_43278,N_43661);
nand U48811 (N_48811,N_41668,N_40949);
or U48812 (N_48812,N_40641,N_40238);
nand U48813 (N_48813,N_42129,N_42375);
and U48814 (N_48814,N_44553,N_40834);
nor U48815 (N_48815,N_41384,N_40381);
and U48816 (N_48816,N_40203,N_42052);
nand U48817 (N_48817,N_43040,N_44355);
nor U48818 (N_48818,N_40329,N_41875);
or U48819 (N_48819,N_41340,N_41082);
nor U48820 (N_48820,N_40158,N_41477);
nand U48821 (N_48821,N_43016,N_41879);
nor U48822 (N_48822,N_44121,N_44654);
or U48823 (N_48823,N_43256,N_42667);
and U48824 (N_48824,N_43709,N_43198);
xnor U48825 (N_48825,N_43252,N_44385);
or U48826 (N_48826,N_40116,N_41653);
nor U48827 (N_48827,N_42100,N_42659);
nand U48828 (N_48828,N_42435,N_40179);
or U48829 (N_48829,N_41471,N_40988);
or U48830 (N_48830,N_42237,N_43432);
nand U48831 (N_48831,N_40255,N_40832);
or U48832 (N_48832,N_40966,N_43022);
nor U48833 (N_48833,N_44088,N_43083);
and U48834 (N_48834,N_44791,N_42611);
xor U48835 (N_48835,N_40514,N_42978);
or U48836 (N_48836,N_44178,N_43389);
nand U48837 (N_48837,N_40753,N_43638);
or U48838 (N_48838,N_42013,N_42548);
nor U48839 (N_48839,N_44009,N_40375);
and U48840 (N_48840,N_43963,N_44758);
nor U48841 (N_48841,N_43818,N_41923);
or U48842 (N_48842,N_41119,N_41957);
nand U48843 (N_48843,N_41427,N_43095);
nor U48844 (N_48844,N_40868,N_44934);
xnor U48845 (N_48845,N_43535,N_43231);
nand U48846 (N_48846,N_41565,N_44032);
and U48847 (N_48847,N_43156,N_40982);
nor U48848 (N_48848,N_40577,N_42688);
or U48849 (N_48849,N_42418,N_41009);
nor U48850 (N_48850,N_40932,N_40734);
or U48851 (N_48851,N_42159,N_42188);
nor U48852 (N_48852,N_40271,N_44228);
or U48853 (N_48853,N_42746,N_41757);
nor U48854 (N_48854,N_40794,N_44649);
nand U48855 (N_48855,N_41185,N_41251);
nor U48856 (N_48856,N_40026,N_41448);
and U48857 (N_48857,N_42515,N_44170);
nand U48858 (N_48858,N_44188,N_42426);
nand U48859 (N_48859,N_40410,N_43821);
nand U48860 (N_48860,N_44130,N_42660);
and U48861 (N_48861,N_40643,N_41627);
and U48862 (N_48862,N_42579,N_41701);
or U48863 (N_48863,N_40054,N_43721);
nand U48864 (N_48864,N_44359,N_43770);
and U48865 (N_48865,N_44157,N_41392);
or U48866 (N_48866,N_43344,N_44167);
nor U48867 (N_48867,N_44467,N_44655);
and U48868 (N_48868,N_40052,N_41821);
nor U48869 (N_48869,N_44452,N_42077);
nand U48870 (N_48870,N_41174,N_40865);
nand U48871 (N_48871,N_41349,N_44781);
nor U48872 (N_48872,N_41129,N_42014);
xnor U48873 (N_48873,N_41666,N_40733);
and U48874 (N_48874,N_43579,N_41085);
nor U48875 (N_48875,N_41437,N_40101);
and U48876 (N_48876,N_43338,N_40082);
xnor U48877 (N_48877,N_40295,N_43379);
xnor U48878 (N_48878,N_44236,N_43745);
or U48879 (N_48879,N_44931,N_40581);
nand U48880 (N_48880,N_42323,N_44409);
nand U48881 (N_48881,N_44751,N_41707);
nand U48882 (N_48882,N_43832,N_41226);
nand U48883 (N_48883,N_41958,N_40453);
nand U48884 (N_48884,N_42386,N_44453);
and U48885 (N_48885,N_40300,N_41362);
nor U48886 (N_48886,N_44691,N_42513);
or U48887 (N_48887,N_40319,N_44505);
or U48888 (N_48888,N_40427,N_43448);
and U48889 (N_48889,N_44391,N_42911);
nor U48890 (N_48890,N_42783,N_41569);
and U48891 (N_48891,N_40536,N_43804);
and U48892 (N_48892,N_40010,N_41985);
xnor U48893 (N_48893,N_42909,N_44124);
or U48894 (N_48894,N_40623,N_44552);
nand U48895 (N_48895,N_44171,N_44830);
nor U48896 (N_48896,N_42953,N_43922);
nor U48897 (N_48897,N_41740,N_42678);
and U48898 (N_48898,N_41077,N_44732);
or U48899 (N_48899,N_41222,N_43279);
nor U48900 (N_48900,N_40834,N_42523);
nor U48901 (N_48901,N_40667,N_44101);
nor U48902 (N_48902,N_43882,N_41243);
and U48903 (N_48903,N_40662,N_42510);
and U48904 (N_48904,N_43787,N_44105);
nor U48905 (N_48905,N_43308,N_43292);
nor U48906 (N_48906,N_42622,N_41566);
nor U48907 (N_48907,N_42146,N_44730);
nor U48908 (N_48908,N_44897,N_44357);
nand U48909 (N_48909,N_43014,N_43198);
and U48910 (N_48910,N_44275,N_43228);
or U48911 (N_48911,N_44966,N_44761);
nor U48912 (N_48912,N_44546,N_43157);
nor U48913 (N_48913,N_42800,N_43002);
or U48914 (N_48914,N_43281,N_44739);
nand U48915 (N_48915,N_41687,N_44453);
nor U48916 (N_48916,N_43473,N_40889);
xnor U48917 (N_48917,N_40211,N_41424);
and U48918 (N_48918,N_43315,N_42527);
xor U48919 (N_48919,N_43589,N_42786);
and U48920 (N_48920,N_44467,N_44079);
nor U48921 (N_48921,N_40510,N_43409);
or U48922 (N_48922,N_42709,N_40306);
nor U48923 (N_48923,N_42203,N_43534);
and U48924 (N_48924,N_44028,N_43139);
xor U48925 (N_48925,N_44073,N_40267);
nor U48926 (N_48926,N_41743,N_42429);
and U48927 (N_48927,N_44349,N_43343);
or U48928 (N_48928,N_41144,N_41442);
nand U48929 (N_48929,N_41248,N_41012);
nor U48930 (N_48930,N_42919,N_42883);
or U48931 (N_48931,N_44263,N_43319);
or U48932 (N_48932,N_41287,N_42415);
or U48933 (N_48933,N_42176,N_41211);
xnor U48934 (N_48934,N_42640,N_41834);
and U48935 (N_48935,N_41398,N_43000);
or U48936 (N_48936,N_41213,N_41502);
or U48937 (N_48937,N_41591,N_40990);
or U48938 (N_48938,N_41718,N_41934);
nand U48939 (N_48939,N_43995,N_41401);
xnor U48940 (N_48940,N_43006,N_44103);
xnor U48941 (N_48941,N_41622,N_40133);
xnor U48942 (N_48942,N_41341,N_40737);
xnor U48943 (N_48943,N_41463,N_41098);
nor U48944 (N_48944,N_44344,N_44758);
nor U48945 (N_48945,N_40554,N_42045);
nor U48946 (N_48946,N_40811,N_42614);
nand U48947 (N_48947,N_43873,N_41233);
nor U48948 (N_48948,N_43954,N_42506);
nand U48949 (N_48949,N_44735,N_42436);
nor U48950 (N_48950,N_43935,N_40096);
and U48951 (N_48951,N_42397,N_44978);
nand U48952 (N_48952,N_40637,N_41738);
and U48953 (N_48953,N_41354,N_43968);
nor U48954 (N_48954,N_43010,N_44925);
nor U48955 (N_48955,N_43746,N_40524);
and U48956 (N_48956,N_42337,N_42471);
or U48957 (N_48957,N_41429,N_43996);
nor U48958 (N_48958,N_41072,N_42345);
and U48959 (N_48959,N_41364,N_44323);
nor U48960 (N_48960,N_41247,N_41786);
nand U48961 (N_48961,N_40234,N_42096);
and U48962 (N_48962,N_44730,N_43494);
or U48963 (N_48963,N_40332,N_44434);
and U48964 (N_48964,N_43388,N_43159);
and U48965 (N_48965,N_44703,N_41369);
or U48966 (N_48966,N_41030,N_43360);
nand U48967 (N_48967,N_41168,N_40826);
and U48968 (N_48968,N_40570,N_44603);
nor U48969 (N_48969,N_43611,N_42361);
and U48970 (N_48970,N_43924,N_42031);
nor U48971 (N_48971,N_40015,N_43205);
or U48972 (N_48972,N_44919,N_40943);
nand U48973 (N_48973,N_43442,N_42111);
nor U48974 (N_48974,N_41258,N_43910);
nor U48975 (N_48975,N_42251,N_41305);
and U48976 (N_48976,N_44012,N_40565);
nor U48977 (N_48977,N_44805,N_42824);
nor U48978 (N_48978,N_41371,N_40334);
and U48979 (N_48979,N_44485,N_40003);
or U48980 (N_48980,N_41713,N_42549);
nand U48981 (N_48981,N_43590,N_40762);
nand U48982 (N_48982,N_43899,N_42987);
nand U48983 (N_48983,N_44501,N_41249);
nor U48984 (N_48984,N_42370,N_43238);
or U48985 (N_48985,N_42058,N_43033);
nand U48986 (N_48986,N_41049,N_41308);
and U48987 (N_48987,N_41076,N_41313);
nand U48988 (N_48988,N_41454,N_43226);
nand U48989 (N_48989,N_41712,N_43729);
and U48990 (N_48990,N_44871,N_40981);
or U48991 (N_48991,N_43159,N_42019);
or U48992 (N_48992,N_42392,N_44746);
and U48993 (N_48993,N_41011,N_43701);
nor U48994 (N_48994,N_42172,N_42826);
nor U48995 (N_48995,N_42760,N_42159);
or U48996 (N_48996,N_42093,N_44503);
or U48997 (N_48997,N_42054,N_42707);
nor U48998 (N_48998,N_43500,N_43160);
xor U48999 (N_48999,N_43002,N_43392);
and U49000 (N_49000,N_44695,N_43084);
nor U49001 (N_49001,N_40065,N_42783);
nand U49002 (N_49002,N_41004,N_42003);
or U49003 (N_49003,N_41800,N_44568);
and U49004 (N_49004,N_44139,N_42951);
or U49005 (N_49005,N_41791,N_41674);
xnor U49006 (N_49006,N_44660,N_43063);
nand U49007 (N_49007,N_44096,N_44816);
nand U49008 (N_49008,N_40016,N_43290);
or U49009 (N_49009,N_43454,N_43863);
or U49010 (N_49010,N_40610,N_44432);
nand U49011 (N_49011,N_42777,N_42515);
or U49012 (N_49012,N_43509,N_41564);
or U49013 (N_49013,N_43508,N_44905);
or U49014 (N_49014,N_40051,N_42148);
and U49015 (N_49015,N_43417,N_42971);
xnor U49016 (N_49016,N_41554,N_41094);
and U49017 (N_49017,N_42832,N_41458);
or U49018 (N_49018,N_42444,N_43286);
xnor U49019 (N_49019,N_44350,N_41110);
nand U49020 (N_49020,N_42047,N_40046);
nor U49021 (N_49021,N_41171,N_43303);
nand U49022 (N_49022,N_43705,N_44536);
or U49023 (N_49023,N_40723,N_40935);
or U49024 (N_49024,N_41162,N_41067);
and U49025 (N_49025,N_40119,N_41990);
nand U49026 (N_49026,N_44204,N_41553);
and U49027 (N_49027,N_43296,N_44328);
nand U49028 (N_49028,N_43230,N_44198);
nand U49029 (N_49029,N_40962,N_43397);
nand U49030 (N_49030,N_44867,N_44101);
or U49031 (N_49031,N_40118,N_41605);
or U49032 (N_49032,N_44336,N_42528);
and U49033 (N_49033,N_43612,N_42421);
or U49034 (N_49034,N_41082,N_41114);
nand U49035 (N_49035,N_42386,N_41376);
xor U49036 (N_49036,N_44620,N_41571);
and U49037 (N_49037,N_40721,N_42004);
nor U49038 (N_49038,N_42686,N_44039);
nand U49039 (N_49039,N_41685,N_42944);
and U49040 (N_49040,N_40277,N_44554);
and U49041 (N_49041,N_44793,N_42430);
nand U49042 (N_49042,N_44598,N_41951);
or U49043 (N_49043,N_42075,N_43641);
nor U49044 (N_49044,N_44108,N_41359);
nand U49045 (N_49045,N_42821,N_42977);
nor U49046 (N_49046,N_44585,N_43708);
and U49047 (N_49047,N_41508,N_44757);
xor U49048 (N_49048,N_44027,N_41454);
nand U49049 (N_49049,N_44415,N_43200);
nor U49050 (N_49050,N_44189,N_44646);
nand U49051 (N_49051,N_43980,N_44896);
nor U49052 (N_49052,N_40900,N_40310);
nor U49053 (N_49053,N_40403,N_41025);
and U49054 (N_49054,N_42383,N_40698);
nor U49055 (N_49055,N_43100,N_44326);
nor U49056 (N_49056,N_44764,N_41690);
and U49057 (N_49057,N_43993,N_40674);
or U49058 (N_49058,N_42747,N_40063);
nor U49059 (N_49059,N_44437,N_43218);
and U49060 (N_49060,N_43598,N_41356);
nor U49061 (N_49061,N_40834,N_44712);
xnor U49062 (N_49062,N_44089,N_43284);
nand U49063 (N_49063,N_40773,N_42376);
and U49064 (N_49064,N_43500,N_44043);
nand U49065 (N_49065,N_40897,N_40396);
nand U49066 (N_49066,N_43640,N_42567);
and U49067 (N_49067,N_43112,N_42834);
and U49068 (N_49068,N_40304,N_44371);
or U49069 (N_49069,N_42449,N_42961);
nor U49070 (N_49070,N_44157,N_43282);
nand U49071 (N_49071,N_40348,N_44868);
and U49072 (N_49072,N_43313,N_44667);
and U49073 (N_49073,N_44486,N_40030);
nor U49074 (N_49074,N_44768,N_44782);
nor U49075 (N_49075,N_40866,N_42124);
nor U49076 (N_49076,N_41392,N_40607);
or U49077 (N_49077,N_42250,N_40905);
or U49078 (N_49078,N_41754,N_41414);
or U49079 (N_49079,N_41494,N_40390);
nor U49080 (N_49080,N_42022,N_44836);
xnor U49081 (N_49081,N_40206,N_42871);
nand U49082 (N_49082,N_43504,N_44203);
and U49083 (N_49083,N_40311,N_41948);
and U49084 (N_49084,N_43309,N_43458);
nand U49085 (N_49085,N_43185,N_42961);
and U49086 (N_49086,N_42310,N_42712);
nor U49087 (N_49087,N_43641,N_42419);
nor U49088 (N_49088,N_43338,N_41919);
nand U49089 (N_49089,N_41446,N_40745);
nor U49090 (N_49090,N_41349,N_41943);
and U49091 (N_49091,N_43121,N_44205);
and U49092 (N_49092,N_43895,N_44666);
and U49093 (N_49093,N_43681,N_44086);
or U49094 (N_49094,N_44845,N_43738);
and U49095 (N_49095,N_44088,N_40412);
nand U49096 (N_49096,N_41334,N_40960);
nor U49097 (N_49097,N_44249,N_42948);
nand U49098 (N_49098,N_41343,N_42137);
nor U49099 (N_49099,N_42903,N_43217);
or U49100 (N_49100,N_44818,N_41668);
nor U49101 (N_49101,N_43628,N_42325);
nor U49102 (N_49102,N_42042,N_43680);
nor U49103 (N_49103,N_42265,N_40719);
or U49104 (N_49104,N_42781,N_44430);
xor U49105 (N_49105,N_40856,N_42684);
nand U49106 (N_49106,N_41205,N_43855);
and U49107 (N_49107,N_41130,N_43219);
and U49108 (N_49108,N_43182,N_42476);
and U49109 (N_49109,N_44035,N_42789);
or U49110 (N_49110,N_40487,N_40038);
and U49111 (N_49111,N_41683,N_40679);
or U49112 (N_49112,N_41838,N_41393);
xnor U49113 (N_49113,N_42053,N_44834);
nand U49114 (N_49114,N_42650,N_44939);
nor U49115 (N_49115,N_42912,N_42346);
and U49116 (N_49116,N_43030,N_40900);
and U49117 (N_49117,N_44700,N_40793);
xnor U49118 (N_49118,N_44262,N_44192);
or U49119 (N_49119,N_41821,N_42404);
xor U49120 (N_49120,N_42480,N_40095);
nor U49121 (N_49121,N_43030,N_43725);
and U49122 (N_49122,N_43106,N_40416);
or U49123 (N_49123,N_41425,N_40723);
nand U49124 (N_49124,N_42002,N_43311);
nor U49125 (N_49125,N_40987,N_41219);
nor U49126 (N_49126,N_41562,N_40497);
nand U49127 (N_49127,N_44685,N_40531);
nand U49128 (N_49128,N_43539,N_40073);
or U49129 (N_49129,N_41605,N_43358);
xnor U49130 (N_49130,N_40888,N_44472);
nand U49131 (N_49131,N_43730,N_43347);
xnor U49132 (N_49132,N_40225,N_41862);
and U49133 (N_49133,N_41080,N_43488);
or U49134 (N_49134,N_40153,N_43554);
or U49135 (N_49135,N_42186,N_44391);
nand U49136 (N_49136,N_44680,N_44195);
nand U49137 (N_49137,N_42472,N_41248);
nand U49138 (N_49138,N_43934,N_42773);
nand U49139 (N_49139,N_43661,N_44309);
nand U49140 (N_49140,N_44824,N_40565);
nor U49141 (N_49141,N_43686,N_40421);
nand U49142 (N_49142,N_44826,N_40716);
nand U49143 (N_49143,N_40124,N_41416);
or U49144 (N_49144,N_42938,N_44705);
xor U49145 (N_49145,N_44560,N_44372);
and U49146 (N_49146,N_43488,N_41411);
nand U49147 (N_49147,N_42370,N_43359);
and U49148 (N_49148,N_40500,N_41001);
nand U49149 (N_49149,N_44719,N_44264);
nor U49150 (N_49150,N_42828,N_44173);
nand U49151 (N_49151,N_42034,N_44382);
nand U49152 (N_49152,N_43709,N_44833);
and U49153 (N_49153,N_42698,N_41802);
nand U49154 (N_49154,N_44110,N_44214);
nor U49155 (N_49155,N_41672,N_44689);
or U49156 (N_49156,N_44433,N_43538);
nor U49157 (N_49157,N_43977,N_41440);
xnor U49158 (N_49158,N_42555,N_43065);
nand U49159 (N_49159,N_41750,N_41492);
nor U49160 (N_49160,N_42358,N_41703);
or U49161 (N_49161,N_40311,N_43420);
and U49162 (N_49162,N_42923,N_40285);
nor U49163 (N_49163,N_40601,N_42656);
nor U49164 (N_49164,N_40118,N_40986);
or U49165 (N_49165,N_43506,N_43123);
or U49166 (N_49166,N_41899,N_44083);
and U49167 (N_49167,N_44254,N_42513);
nand U49168 (N_49168,N_41355,N_43225);
nand U49169 (N_49169,N_40409,N_40838);
nor U49170 (N_49170,N_41981,N_43851);
xnor U49171 (N_49171,N_43285,N_44874);
or U49172 (N_49172,N_42261,N_41682);
and U49173 (N_49173,N_43519,N_40559);
and U49174 (N_49174,N_41252,N_44679);
and U49175 (N_49175,N_41657,N_41010);
or U49176 (N_49176,N_44146,N_44533);
nand U49177 (N_49177,N_40911,N_41242);
or U49178 (N_49178,N_41605,N_42545);
or U49179 (N_49179,N_42458,N_41020);
or U49180 (N_49180,N_43977,N_44771);
nand U49181 (N_49181,N_43605,N_44919);
and U49182 (N_49182,N_43096,N_44208);
nor U49183 (N_49183,N_43143,N_40729);
and U49184 (N_49184,N_43860,N_43241);
nand U49185 (N_49185,N_40619,N_43077);
nor U49186 (N_49186,N_41881,N_43895);
or U49187 (N_49187,N_41377,N_42100);
and U49188 (N_49188,N_42322,N_40771);
and U49189 (N_49189,N_43171,N_44936);
nor U49190 (N_49190,N_42331,N_43845);
xor U49191 (N_49191,N_40142,N_41295);
nand U49192 (N_49192,N_40406,N_43786);
nor U49193 (N_49193,N_43489,N_43347);
nand U49194 (N_49194,N_43873,N_43473);
or U49195 (N_49195,N_40747,N_42722);
nor U49196 (N_49196,N_42900,N_40336);
xnor U49197 (N_49197,N_43269,N_40226);
and U49198 (N_49198,N_44416,N_40159);
nand U49199 (N_49199,N_43634,N_41355);
and U49200 (N_49200,N_40248,N_43368);
or U49201 (N_49201,N_44969,N_43456);
nor U49202 (N_49202,N_41546,N_43294);
and U49203 (N_49203,N_40005,N_41349);
nand U49204 (N_49204,N_41004,N_42267);
nand U49205 (N_49205,N_40545,N_44901);
nand U49206 (N_49206,N_43018,N_42167);
nand U49207 (N_49207,N_44196,N_42004);
or U49208 (N_49208,N_42570,N_42673);
and U49209 (N_49209,N_43874,N_43951);
and U49210 (N_49210,N_42490,N_42375);
nor U49211 (N_49211,N_41579,N_41555);
nor U49212 (N_49212,N_43032,N_42338);
nand U49213 (N_49213,N_42846,N_44060);
nor U49214 (N_49214,N_40351,N_43550);
and U49215 (N_49215,N_41330,N_44101);
and U49216 (N_49216,N_42105,N_44499);
nor U49217 (N_49217,N_40669,N_40862);
and U49218 (N_49218,N_41472,N_44798);
nor U49219 (N_49219,N_44102,N_43168);
nand U49220 (N_49220,N_43764,N_42960);
and U49221 (N_49221,N_43920,N_43309);
and U49222 (N_49222,N_42544,N_43806);
or U49223 (N_49223,N_43079,N_43309);
and U49224 (N_49224,N_41369,N_44661);
or U49225 (N_49225,N_41523,N_40439);
and U49226 (N_49226,N_43121,N_41514);
or U49227 (N_49227,N_44518,N_43924);
nand U49228 (N_49228,N_40703,N_40208);
and U49229 (N_49229,N_42653,N_43998);
xnor U49230 (N_49230,N_40517,N_40394);
nor U49231 (N_49231,N_43444,N_40123);
and U49232 (N_49232,N_40157,N_42633);
and U49233 (N_49233,N_44501,N_43477);
nor U49234 (N_49234,N_41993,N_44039);
and U49235 (N_49235,N_42070,N_43091);
or U49236 (N_49236,N_42665,N_43820);
or U49237 (N_49237,N_41895,N_41880);
nand U49238 (N_49238,N_44501,N_43648);
or U49239 (N_49239,N_44924,N_40380);
nand U49240 (N_49240,N_40268,N_44209);
or U49241 (N_49241,N_43427,N_44886);
and U49242 (N_49242,N_42575,N_43177);
nand U49243 (N_49243,N_43488,N_40684);
nor U49244 (N_49244,N_43355,N_41683);
nor U49245 (N_49245,N_40824,N_44733);
nand U49246 (N_49246,N_42835,N_40956);
nand U49247 (N_49247,N_41540,N_44547);
or U49248 (N_49248,N_43415,N_42256);
xor U49249 (N_49249,N_44758,N_44237);
xor U49250 (N_49250,N_41747,N_44020);
or U49251 (N_49251,N_41101,N_41077);
or U49252 (N_49252,N_40077,N_40427);
xnor U49253 (N_49253,N_41008,N_43549);
and U49254 (N_49254,N_41618,N_44459);
nor U49255 (N_49255,N_44769,N_41762);
xor U49256 (N_49256,N_42478,N_40336);
nand U49257 (N_49257,N_41272,N_41688);
nor U49258 (N_49258,N_40269,N_40133);
nand U49259 (N_49259,N_43517,N_44757);
and U49260 (N_49260,N_42541,N_40230);
or U49261 (N_49261,N_43526,N_42944);
or U49262 (N_49262,N_41752,N_40131);
or U49263 (N_49263,N_42732,N_42127);
nor U49264 (N_49264,N_42161,N_42936);
xor U49265 (N_49265,N_43633,N_42008);
nor U49266 (N_49266,N_41551,N_40170);
nor U49267 (N_49267,N_42041,N_44450);
nand U49268 (N_49268,N_44820,N_40328);
and U49269 (N_49269,N_43074,N_41842);
and U49270 (N_49270,N_44796,N_41780);
or U49271 (N_49271,N_42049,N_41744);
nand U49272 (N_49272,N_43353,N_42763);
nor U49273 (N_49273,N_44436,N_44388);
or U49274 (N_49274,N_44318,N_40994);
or U49275 (N_49275,N_42278,N_44687);
xnor U49276 (N_49276,N_41051,N_41049);
or U49277 (N_49277,N_40894,N_41838);
nor U49278 (N_49278,N_42865,N_41246);
nand U49279 (N_49279,N_42161,N_43751);
and U49280 (N_49280,N_41493,N_44794);
nor U49281 (N_49281,N_42077,N_40078);
xnor U49282 (N_49282,N_42578,N_42831);
nand U49283 (N_49283,N_44800,N_42162);
xor U49284 (N_49284,N_41680,N_42046);
and U49285 (N_49285,N_42732,N_42187);
and U49286 (N_49286,N_44569,N_40503);
nand U49287 (N_49287,N_42013,N_42845);
nand U49288 (N_49288,N_42740,N_44446);
or U49289 (N_49289,N_44206,N_44314);
nor U49290 (N_49290,N_41487,N_40146);
nor U49291 (N_49291,N_42966,N_44673);
and U49292 (N_49292,N_42410,N_42379);
or U49293 (N_49293,N_44225,N_42100);
nor U49294 (N_49294,N_41249,N_41248);
nand U49295 (N_49295,N_42467,N_44340);
and U49296 (N_49296,N_40203,N_42234);
and U49297 (N_49297,N_43767,N_40586);
or U49298 (N_49298,N_44024,N_43268);
nand U49299 (N_49299,N_42300,N_40293);
and U49300 (N_49300,N_43700,N_42263);
nor U49301 (N_49301,N_41744,N_40923);
nand U49302 (N_49302,N_41613,N_43175);
nand U49303 (N_49303,N_43280,N_41431);
nor U49304 (N_49304,N_42574,N_44570);
or U49305 (N_49305,N_40201,N_43580);
and U49306 (N_49306,N_42143,N_44777);
nor U49307 (N_49307,N_43342,N_44092);
nand U49308 (N_49308,N_42069,N_44095);
or U49309 (N_49309,N_44835,N_40513);
and U49310 (N_49310,N_41867,N_43494);
nand U49311 (N_49311,N_41189,N_40864);
nand U49312 (N_49312,N_42816,N_40149);
and U49313 (N_49313,N_40745,N_41225);
and U49314 (N_49314,N_44408,N_42158);
nor U49315 (N_49315,N_42319,N_40982);
xnor U49316 (N_49316,N_42020,N_43996);
nor U49317 (N_49317,N_40428,N_43725);
or U49318 (N_49318,N_43030,N_41666);
nor U49319 (N_49319,N_42636,N_42353);
nor U49320 (N_49320,N_43873,N_44715);
and U49321 (N_49321,N_41104,N_41731);
nand U49322 (N_49322,N_42654,N_44803);
or U49323 (N_49323,N_42303,N_43901);
nand U49324 (N_49324,N_44569,N_44149);
and U49325 (N_49325,N_40323,N_44142);
or U49326 (N_49326,N_43631,N_43260);
nor U49327 (N_49327,N_44152,N_41870);
xor U49328 (N_49328,N_40002,N_42047);
nand U49329 (N_49329,N_44022,N_41180);
or U49330 (N_49330,N_42617,N_40589);
or U49331 (N_49331,N_41173,N_43760);
and U49332 (N_49332,N_43056,N_42813);
and U49333 (N_49333,N_43589,N_40074);
and U49334 (N_49334,N_41909,N_40299);
nand U49335 (N_49335,N_40360,N_43784);
nor U49336 (N_49336,N_43593,N_44718);
nor U49337 (N_49337,N_43455,N_42585);
or U49338 (N_49338,N_43871,N_43481);
nand U49339 (N_49339,N_40510,N_40323);
nor U49340 (N_49340,N_40572,N_44989);
or U49341 (N_49341,N_43256,N_40053);
xor U49342 (N_49342,N_43005,N_43781);
nor U49343 (N_49343,N_44082,N_41130);
nand U49344 (N_49344,N_41696,N_40202);
and U49345 (N_49345,N_41478,N_42183);
nand U49346 (N_49346,N_41353,N_43705);
and U49347 (N_49347,N_40825,N_44131);
or U49348 (N_49348,N_42005,N_42352);
nor U49349 (N_49349,N_44697,N_44809);
and U49350 (N_49350,N_42884,N_43981);
nand U49351 (N_49351,N_43023,N_42441);
and U49352 (N_49352,N_43208,N_43300);
nor U49353 (N_49353,N_44731,N_40734);
nand U49354 (N_49354,N_40387,N_40459);
nor U49355 (N_49355,N_44256,N_41668);
and U49356 (N_49356,N_40483,N_43630);
xnor U49357 (N_49357,N_43380,N_41110);
nand U49358 (N_49358,N_40938,N_44719);
xor U49359 (N_49359,N_43050,N_41888);
nand U49360 (N_49360,N_41146,N_42062);
nor U49361 (N_49361,N_44816,N_41215);
and U49362 (N_49362,N_43299,N_41508);
and U49363 (N_49363,N_41406,N_44283);
or U49364 (N_49364,N_43315,N_40121);
nor U49365 (N_49365,N_40731,N_44229);
and U49366 (N_49366,N_42693,N_43136);
nand U49367 (N_49367,N_41627,N_43972);
nor U49368 (N_49368,N_40644,N_41547);
nor U49369 (N_49369,N_40496,N_44558);
nand U49370 (N_49370,N_44241,N_41935);
and U49371 (N_49371,N_42032,N_41676);
nor U49372 (N_49372,N_40380,N_42782);
nor U49373 (N_49373,N_43641,N_40795);
xnor U49374 (N_49374,N_40849,N_43795);
or U49375 (N_49375,N_44412,N_40098);
or U49376 (N_49376,N_40175,N_41611);
nand U49377 (N_49377,N_42197,N_43574);
nor U49378 (N_49378,N_42918,N_44105);
nand U49379 (N_49379,N_40660,N_41717);
or U49380 (N_49380,N_44574,N_44446);
or U49381 (N_49381,N_40497,N_43056);
and U49382 (N_49382,N_41782,N_40915);
nand U49383 (N_49383,N_41904,N_42527);
nand U49384 (N_49384,N_41218,N_41345);
or U49385 (N_49385,N_43349,N_40763);
nor U49386 (N_49386,N_41091,N_44210);
nor U49387 (N_49387,N_42464,N_40834);
and U49388 (N_49388,N_43211,N_44472);
and U49389 (N_49389,N_44183,N_41322);
and U49390 (N_49390,N_41247,N_40350);
or U49391 (N_49391,N_42438,N_41257);
and U49392 (N_49392,N_42684,N_41475);
and U49393 (N_49393,N_43470,N_40525);
nand U49394 (N_49394,N_41145,N_44901);
xor U49395 (N_49395,N_44452,N_41291);
nor U49396 (N_49396,N_40357,N_44353);
and U49397 (N_49397,N_44354,N_40989);
or U49398 (N_49398,N_44159,N_42913);
nor U49399 (N_49399,N_43376,N_40537);
or U49400 (N_49400,N_42852,N_44031);
nor U49401 (N_49401,N_42205,N_41877);
and U49402 (N_49402,N_44043,N_42052);
and U49403 (N_49403,N_42191,N_43035);
nand U49404 (N_49404,N_42608,N_41189);
and U49405 (N_49405,N_41669,N_42491);
xnor U49406 (N_49406,N_41298,N_40637);
xor U49407 (N_49407,N_44267,N_42062);
or U49408 (N_49408,N_41229,N_40587);
nor U49409 (N_49409,N_44781,N_40991);
and U49410 (N_49410,N_42890,N_43816);
or U49411 (N_49411,N_44552,N_40595);
and U49412 (N_49412,N_43121,N_42397);
or U49413 (N_49413,N_41488,N_43456);
or U49414 (N_49414,N_43626,N_42635);
and U49415 (N_49415,N_43790,N_42540);
nand U49416 (N_49416,N_41811,N_44051);
nand U49417 (N_49417,N_41051,N_44401);
or U49418 (N_49418,N_41489,N_43541);
nor U49419 (N_49419,N_41842,N_40308);
nand U49420 (N_49420,N_41046,N_43917);
or U49421 (N_49421,N_42911,N_44001);
nand U49422 (N_49422,N_40252,N_44348);
nand U49423 (N_49423,N_42792,N_44412);
nand U49424 (N_49424,N_43345,N_44865);
and U49425 (N_49425,N_43562,N_43826);
nor U49426 (N_49426,N_42907,N_43764);
or U49427 (N_49427,N_42593,N_44900);
nand U49428 (N_49428,N_44133,N_40506);
nor U49429 (N_49429,N_42085,N_41775);
and U49430 (N_49430,N_41357,N_41913);
or U49431 (N_49431,N_40567,N_44519);
nor U49432 (N_49432,N_41186,N_44237);
nand U49433 (N_49433,N_41577,N_42461);
nor U49434 (N_49434,N_43914,N_44687);
nand U49435 (N_49435,N_44301,N_43593);
and U49436 (N_49436,N_44970,N_42301);
nand U49437 (N_49437,N_43134,N_44114);
or U49438 (N_49438,N_44789,N_42708);
or U49439 (N_49439,N_43163,N_42136);
xor U49440 (N_49440,N_42159,N_42907);
and U49441 (N_49441,N_44564,N_43514);
nor U49442 (N_49442,N_41908,N_40092);
nor U49443 (N_49443,N_44692,N_40442);
nand U49444 (N_49444,N_41394,N_41564);
nor U49445 (N_49445,N_43627,N_44319);
and U49446 (N_49446,N_40144,N_41606);
and U49447 (N_49447,N_42520,N_40458);
nand U49448 (N_49448,N_44658,N_41107);
nand U49449 (N_49449,N_44781,N_44425);
or U49450 (N_49450,N_43599,N_40003);
and U49451 (N_49451,N_42064,N_41503);
nand U49452 (N_49452,N_44673,N_44816);
nand U49453 (N_49453,N_43136,N_41547);
and U49454 (N_49454,N_42744,N_42081);
nand U49455 (N_49455,N_41540,N_42567);
nor U49456 (N_49456,N_44993,N_41304);
nand U49457 (N_49457,N_43048,N_40938);
and U49458 (N_49458,N_41001,N_43075);
and U49459 (N_49459,N_42770,N_40771);
and U49460 (N_49460,N_43430,N_42691);
and U49461 (N_49461,N_41242,N_42640);
xnor U49462 (N_49462,N_42990,N_41836);
nor U49463 (N_49463,N_40097,N_44241);
nor U49464 (N_49464,N_41281,N_41217);
and U49465 (N_49465,N_44267,N_42355);
and U49466 (N_49466,N_43152,N_40807);
and U49467 (N_49467,N_44278,N_40285);
and U49468 (N_49468,N_44910,N_43894);
nand U49469 (N_49469,N_40190,N_41390);
and U49470 (N_49470,N_43874,N_44606);
nor U49471 (N_49471,N_43744,N_43096);
nor U49472 (N_49472,N_40649,N_41493);
and U49473 (N_49473,N_43520,N_41649);
or U49474 (N_49474,N_40295,N_43158);
and U49475 (N_49475,N_44415,N_44533);
or U49476 (N_49476,N_42518,N_42244);
nand U49477 (N_49477,N_40018,N_43389);
or U49478 (N_49478,N_40643,N_41848);
and U49479 (N_49479,N_41102,N_42214);
and U49480 (N_49480,N_41234,N_43383);
and U49481 (N_49481,N_41242,N_43078);
and U49482 (N_49482,N_41016,N_40622);
xor U49483 (N_49483,N_42500,N_41656);
and U49484 (N_49484,N_43679,N_41565);
nand U49485 (N_49485,N_44360,N_41539);
xnor U49486 (N_49486,N_43585,N_44316);
nor U49487 (N_49487,N_44193,N_42045);
nor U49488 (N_49488,N_42174,N_44305);
nand U49489 (N_49489,N_44688,N_41216);
nor U49490 (N_49490,N_44143,N_44383);
and U49491 (N_49491,N_40866,N_43011);
or U49492 (N_49492,N_44795,N_42219);
nor U49493 (N_49493,N_40235,N_40048);
or U49494 (N_49494,N_40984,N_43900);
or U49495 (N_49495,N_42341,N_43355);
nand U49496 (N_49496,N_42949,N_40404);
nor U49497 (N_49497,N_43750,N_41819);
nand U49498 (N_49498,N_44526,N_42265);
nor U49499 (N_49499,N_43753,N_42888);
xor U49500 (N_49500,N_42644,N_44889);
nor U49501 (N_49501,N_42776,N_44558);
or U49502 (N_49502,N_42435,N_40581);
and U49503 (N_49503,N_41276,N_41436);
or U49504 (N_49504,N_41671,N_43049);
xor U49505 (N_49505,N_41524,N_44034);
nand U49506 (N_49506,N_42664,N_41401);
nand U49507 (N_49507,N_43638,N_40537);
or U49508 (N_49508,N_40844,N_44149);
or U49509 (N_49509,N_42061,N_40252);
nand U49510 (N_49510,N_40564,N_40190);
nand U49511 (N_49511,N_41229,N_43701);
and U49512 (N_49512,N_42412,N_43176);
xnor U49513 (N_49513,N_42072,N_40810);
xor U49514 (N_49514,N_40917,N_44465);
nand U49515 (N_49515,N_41833,N_43000);
and U49516 (N_49516,N_42691,N_40963);
nand U49517 (N_49517,N_40075,N_40440);
or U49518 (N_49518,N_41385,N_40620);
and U49519 (N_49519,N_40327,N_40080);
nand U49520 (N_49520,N_43455,N_43537);
nor U49521 (N_49521,N_42967,N_43000);
xnor U49522 (N_49522,N_44730,N_41065);
nor U49523 (N_49523,N_42350,N_41984);
nand U49524 (N_49524,N_41194,N_40799);
or U49525 (N_49525,N_40583,N_41396);
or U49526 (N_49526,N_42866,N_44616);
nand U49527 (N_49527,N_43241,N_43170);
nand U49528 (N_49528,N_44216,N_40217);
nand U49529 (N_49529,N_41739,N_42370);
or U49530 (N_49530,N_41017,N_40784);
and U49531 (N_49531,N_42238,N_43781);
or U49532 (N_49532,N_40448,N_42064);
xor U49533 (N_49533,N_44882,N_40114);
and U49534 (N_49534,N_40304,N_40718);
or U49535 (N_49535,N_42148,N_42732);
nor U49536 (N_49536,N_41021,N_42345);
nand U49537 (N_49537,N_44438,N_44045);
nor U49538 (N_49538,N_41914,N_44827);
nand U49539 (N_49539,N_43957,N_42849);
xnor U49540 (N_49540,N_41341,N_40010);
and U49541 (N_49541,N_40450,N_41755);
nor U49542 (N_49542,N_40101,N_40485);
nand U49543 (N_49543,N_41596,N_41205);
nand U49544 (N_49544,N_43963,N_43576);
nor U49545 (N_49545,N_40781,N_43467);
or U49546 (N_49546,N_41420,N_40069);
xnor U49547 (N_49547,N_40339,N_43251);
nor U49548 (N_49548,N_42748,N_42676);
and U49549 (N_49549,N_40725,N_40785);
nand U49550 (N_49550,N_42186,N_41525);
or U49551 (N_49551,N_42010,N_44200);
or U49552 (N_49552,N_42269,N_41835);
nand U49553 (N_49553,N_41321,N_44299);
or U49554 (N_49554,N_42040,N_44317);
nor U49555 (N_49555,N_43476,N_41941);
nand U49556 (N_49556,N_42189,N_43574);
nand U49557 (N_49557,N_41541,N_40800);
nand U49558 (N_49558,N_40814,N_40324);
nor U49559 (N_49559,N_41239,N_42407);
or U49560 (N_49560,N_42188,N_40835);
nor U49561 (N_49561,N_42872,N_41235);
or U49562 (N_49562,N_42920,N_44137);
nand U49563 (N_49563,N_41801,N_40724);
and U49564 (N_49564,N_41007,N_43005);
nand U49565 (N_49565,N_44156,N_44127);
and U49566 (N_49566,N_40426,N_42661);
and U49567 (N_49567,N_41528,N_41606);
or U49568 (N_49568,N_43170,N_44704);
nand U49569 (N_49569,N_42793,N_44890);
or U49570 (N_49570,N_40723,N_44159);
nand U49571 (N_49571,N_41870,N_40145);
and U49572 (N_49572,N_40592,N_42209);
or U49573 (N_49573,N_40127,N_42359);
nand U49574 (N_49574,N_43040,N_41801);
and U49575 (N_49575,N_40567,N_43660);
or U49576 (N_49576,N_41233,N_40674);
nor U49577 (N_49577,N_40359,N_40672);
and U49578 (N_49578,N_43373,N_40260);
and U49579 (N_49579,N_41878,N_40685);
xnor U49580 (N_49580,N_40689,N_40417);
nor U49581 (N_49581,N_44814,N_42903);
or U49582 (N_49582,N_40828,N_42906);
and U49583 (N_49583,N_43847,N_44994);
and U49584 (N_49584,N_41995,N_40369);
or U49585 (N_49585,N_42307,N_41754);
or U49586 (N_49586,N_44978,N_41766);
or U49587 (N_49587,N_42138,N_40951);
nor U49588 (N_49588,N_42975,N_44777);
and U49589 (N_49589,N_43057,N_43847);
nand U49590 (N_49590,N_44730,N_40669);
or U49591 (N_49591,N_40974,N_40675);
and U49592 (N_49592,N_41854,N_41124);
or U49593 (N_49593,N_43424,N_40356);
or U49594 (N_49594,N_41911,N_43822);
nor U49595 (N_49595,N_43987,N_43422);
xnor U49596 (N_49596,N_43457,N_40600);
or U49597 (N_49597,N_40244,N_44555);
and U49598 (N_49598,N_40797,N_44995);
nand U49599 (N_49599,N_40024,N_40893);
and U49600 (N_49600,N_42396,N_42607);
nor U49601 (N_49601,N_44519,N_42748);
and U49602 (N_49602,N_44666,N_42312);
nor U49603 (N_49603,N_44555,N_41157);
nor U49604 (N_49604,N_43509,N_43401);
xor U49605 (N_49605,N_42864,N_44866);
nor U49606 (N_49606,N_40871,N_43580);
nor U49607 (N_49607,N_40457,N_41181);
nand U49608 (N_49608,N_44153,N_43220);
and U49609 (N_49609,N_43728,N_41835);
or U49610 (N_49610,N_40626,N_43260);
nand U49611 (N_49611,N_44585,N_44137);
xor U49612 (N_49612,N_41383,N_40546);
nor U49613 (N_49613,N_40668,N_41370);
or U49614 (N_49614,N_40406,N_42738);
nand U49615 (N_49615,N_42774,N_40272);
or U49616 (N_49616,N_43107,N_40050);
nand U49617 (N_49617,N_41049,N_43714);
or U49618 (N_49618,N_42957,N_41629);
nand U49619 (N_49619,N_43279,N_41424);
or U49620 (N_49620,N_40768,N_44938);
nand U49621 (N_49621,N_43890,N_44158);
nor U49622 (N_49622,N_42981,N_42359);
xnor U49623 (N_49623,N_43017,N_43330);
or U49624 (N_49624,N_40281,N_41850);
xnor U49625 (N_49625,N_41880,N_41606);
nand U49626 (N_49626,N_43164,N_40588);
or U49627 (N_49627,N_44162,N_44498);
xor U49628 (N_49628,N_44935,N_42037);
nand U49629 (N_49629,N_43099,N_43328);
nand U49630 (N_49630,N_40111,N_40066);
and U49631 (N_49631,N_44587,N_41604);
and U49632 (N_49632,N_43656,N_41914);
or U49633 (N_49633,N_41899,N_43466);
xor U49634 (N_49634,N_40482,N_42779);
nor U49635 (N_49635,N_41452,N_40253);
or U49636 (N_49636,N_42850,N_40088);
nand U49637 (N_49637,N_40266,N_44635);
or U49638 (N_49638,N_42478,N_43112);
nor U49639 (N_49639,N_43693,N_42431);
nand U49640 (N_49640,N_44939,N_44222);
or U49641 (N_49641,N_43103,N_42507);
and U49642 (N_49642,N_41649,N_42865);
nor U49643 (N_49643,N_43049,N_40181);
and U49644 (N_49644,N_42081,N_40461);
nand U49645 (N_49645,N_40062,N_44185);
or U49646 (N_49646,N_40977,N_41894);
and U49647 (N_49647,N_44903,N_43766);
xor U49648 (N_49648,N_41574,N_40461);
xor U49649 (N_49649,N_42941,N_44049);
or U49650 (N_49650,N_44406,N_43346);
nand U49651 (N_49651,N_40863,N_40716);
nand U49652 (N_49652,N_40667,N_43472);
nor U49653 (N_49653,N_44277,N_42182);
and U49654 (N_49654,N_44665,N_44478);
nand U49655 (N_49655,N_41893,N_40959);
nor U49656 (N_49656,N_41478,N_44234);
nand U49657 (N_49657,N_43906,N_40946);
nor U49658 (N_49658,N_43820,N_42042);
nor U49659 (N_49659,N_40032,N_42457);
nand U49660 (N_49660,N_44337,N_41926);
or U49661 (N_49661,N_42839,N_41420);
and U49662 (N_49662,N_40782,N_40592);
and U49663 (N_49663,N_44176,N_43650);
or U49664 (N_49664,N_41672,N_42296);
xor U49665 (N_49665,N_44902,N_42191);
nand U49666 (N_49666,N_44684,N_43755);
nor U49667 (N_49667,N_43086,N_41030);
nor U49668 (N_49668,N_41161,N_41997);
nand U49669 (N_49669,N_40794,N_43971);
and U49670 (N_49670,N_44309,N_44651);
xnor U49671 (N_49671,N_43849,N_44321);
or U49672 (N_49672,N_42377,N_43115);
nor U49673 (N_49673,N_44310,N_44447);
and U49674 (N_49674,N_40826,N_40605);
nor U49675 (N_49675,N_41576,N_44649);
xnor U49676 (N_49676,N_40481,N_40855);
or U49677 (N_49677,N_43534,N_40281);
xnor U49678 (N_49678,N_41522,N_42557);
xor U49679 (N_49679,N_42865,N_41332);
or U49680 (N_49680,N_42697,N_44199);
or U49681 (N_49681,N_40869,N_43146);
and U49682 (N_49682,N_41951,N_40280);
and U49683 (N_49683,N_41898,N_42751);
and U49684 (N_49684,N_44050,N_44658);
xnor U49685 (N_49685,N_44848,N_41995);
and U49686 (N_49686,N_40951,N_41468);
nor U49687 (N_49687,N_44278,N_44535);
nand U49688 (N_49688,N_41559,N_41580);
nand U49689 (N_49689,N_44244,N_42398);
and U49690 (N_49690,N_43901,N_40329);
nor U49691 (N_49691,N_43126,N_42034);
xnor U49692 (N_49692,N_40305,N_43933);
nor U49693 (N_49693,N_40279,N_41218);
nand U49694 (N_49694,N_40551,N_40283);
xor U49695 (N_49695,N_44056,N_43012);
nor U49696 (N_49696,N_43214,N_42755);
nand U49697 (N_49697,N_41376,N_41831);
nand U49698 (N_49698,N_40296,N_42993);
nor U49699 (N_49699,N_41455,N_41351);
nand U49700 (N_49700,N_41378,N_40500);
nand U49701 (N_49701,N_40658,N_40133);
xnor U49702 (N_49702,N_43882,N_44761);
nor U49703 (N_49703,N_41455,N_42495);
nor U49704 (N_49704,N_43848,N_43808);
nand U49705 (N_49705,N_41598,N_44160);
xor U49706 (N_49706,N_44727,N_44165);
nand U49707 (N_49707,N_44860,N_41293);
nand U49708 (N_49708,N_40646,N_42963);
nor U49709 (N_49709,N_41120,N_40818);
nand U49710 (N_49710,N_43702,N_41166);
xor U49711 (N_49711,N_40492,N_42360);
or U49712 (N_49712,N_41401,N_42352);
and U49713 (N_49713,N_44667,N_41635);
nand U49714 (N_49714,N_40135,N_40847);
or U49715 (N_49715,N_41161,N_42720);
and U49716 (N_49716,N_44675,N_42486);
nand U49717 (N_49717,N_41200,N_41939);
nand U49718 (N_49718,N_43429,N_40272);
or U49719 (N_49719,N_40710,N_43823);
xnor U49720 (N_49720,N_44187,N_43345);
nand U49721 (N_49721,N_42422,N_42566);
nor U49722 (N_49722,N_41618,N_42894);
nand U49723 (N_49723,N_40333,N_40112);
nor U49724 (N_49724,N_43176,N_40268);
and U49725 (N_49725,N_42118,N_43782);
and U49726 (N_49726,N_44941,N_43699);
or U49727 (N_49727,N_44448,N_43970);
nor U49728 (N_49728,N_44933,N_44507);
nor U49729 (N_49729,N_42972,N_43656);
nand U49730 (N_49730,N_42224,N_42078);
or U49731 (N_49731,N_41776,N_40771);
or U49732 (N_49732,N_40764,N_42640);
or U49733 (N_49733,N_44502,N_42833);
or U49734 (N_49734,N_42305,N_40084);
and U49735 (N_49735,N_41269,N_42160);
nand U49736 (N_49736,N_41353,N_44110);
xnor U49737 (N_49737,N_43367,N_44314);
or U49738 (N_49738,N_41107,N_40674);
and U49739 (N_49739,N_44526,N_40191);
xor U49740 (N_49740,N_42880,N_41002);
nand U49741 (N_49741,N_41361,N_42416);
nand U49742 (N_49742,N_41216,N_43438);
nor U49743 (N_49743,N_42354,N_40366);
xor U49744 (N_49744,N_41946,N_40785);
or U49745 (N_49745,N_42808,N_44589);
xnor U49746 (N_49746,N_44470,N_44950);
and U49747 (N_49747,N_44391,N_41525);
nand U49748 (N_49748,N_42032,N_44242);
or U49749 (N_49749,N_43907,N_43842);
or U49750 (N_49750,N_40837,N_44613);
nand U49751 (N_49751,N_41185,N_44913);
nand U49752 (N_49752,N_43722,N_42024);
and U49753 (N_49753,N_40213,N_42787);
xor U49754 (N_49754,N_43621,N_43382);
nand U49755 (N_49755,N_41888,N_42112);
or U49756 (N_49756,N_40335,N_44353);
nor U49757 (N_49757,N_44437,N_40660);
and U49758 (N_49758,N_44652,N_40396);
nor U49759 (N_49759,N_41495,N_42524);
and U49760 (N_49760,N_42668,N_44393);
nand U49761 (N_49761,N_40509,N_41752);
nand U49762 (N_49762,N_44106,N_42832);
and U49763 (N_49763,N_42325,N_40982);
nor U49764 (N_49764,N_40148,N_43699);
and U49765 (N_49765,N_44187,N_41129);
nand U49766 (N_49766,N_40336,N_41124);
nor U49767 (N_49767,N_40861,N_41240);
and U49768 (N_49768,N_40820,N_44035);
nand U49769 (N_49769,N_40189,N_43706);
or U49770 (N_49770,N_41815,N_44538);
and U49771 (N_49771,N_42571,N_42123);
and U49772 (N_49772,N_42300,N_42243);
or U49773 (N_49773,N_42613,N_43752);
or U49774 (N_49774,N_42820,N_42064);
and U49775 (N_49775,N_40698,N_44511);
or U49776 (N_49776,N_44210,N_41661);
nor U49777 (N_49777,N_40243,N_44476);
or U49778 (N_49778,N_44965,N_41161);
xor U49779 (N_49779,N_43054,N_42080);
and U49780 (N_49780,N_44284,N_40629);
nor U49781 (N_49781,N_42447,N_42910);
nor U49782 (N_49782,N_40840,N_42486);
or U49783 (N_49783,N_40052,N_40507);
or U49784 (N_49784,N_44799,N_43676);
or U49785 (N_49785,N_43425,N_44003);
xnor U49786 (N_49786,N_40977,N_44397);
or U49787 (N_49787,N_42192,N_40008);
nand U49788 (N_49788,N_40084,N_40079);
xor U49789 (N_49789,N_44003,N_40843);
nor U49790 (N_49790,N_40094,N_41522);
nor U49791 (N_49791,N_40693,N_43745);
or U49792 (N_49792,N_43841,N_43405);
and U49793 (N_49793,N_43670,N_44919);
and U49794 (N_49794,N_41591,N_40964);
nor U49795 (N_49795,N_41280,N_41891);
nand U49796 (N_49796,N_41752,N_43178);
xor U49797 (N_49797,N_44338,N_43740);
nand U49798 (N_49798,N_40875,N_41517);
nand U49799 (N_49799,N_42350,N_40100);
xor U49800 (N_49800,N_42321,N_40102);
nor U49801 (N_49801,N_43800,N_41387);
nand U49802 (N_49802,N_42210,N_42331);
nor U49803 (N_49803,N_44767,N_44231);
nor U49804 (N_49804,N_41055,N_42599);
nor U49805 (N_49805,N_43921,N_40766);
xor U49806 (N_49806,N_42572,N_44683);
nor U49807 (N_49807,N_44830,N_43266);
nand U49808 (N_49808,N_41110,N_43331);
nand U49809 (N_49809,N_42926,N_44194);
or U49810 (N_49810,N_41954,N_44807);
or U49811 (N_49811,N_40104,N_42344);
nor U49812 (N_49812,N_43680,N_44125);
and U49813 (N_49813,N_44353,N_41097);
or U49814 (N_49814,N_44371,N_41619);
or U49815 (N_49815,N_44518,N_44877);
nand U49816 (N_49816,N_40720,N_40469);
or U49817 (N_49817,N_41505,N_42391);
or U49818 (N_49818,N_44756,N_44080);
xnor U49819 (N_49819,N_44208,N_42124);
or U49820 (N_49820,N_42861,N_43224);
nand U49821 (N_49821,N_44208,N_43025);
and U49822 (N_49822,N_43052,N_40597);
xor U49823 (N_49823,N_40459,N_44064);
nand U49824 (N_49824,N_44951,N_43209);
nand U49825 (N_49825,N_40918,N_42179);
and U49826 (N_49826,N_43742,N_43663);
and U49827 (N_49827,N_44088,N_43961);
or U49828 (N_49828,N_41392,N_41847);
nor U49829 (N_49829,N_42228,N_44403);
nor U49830 (N_49830,N_41392,N_40459);
and U49831 (N_49831,N_42557,N_41788);
or U49832 (N_49832,N_40557,N_40265);
or U49833 (N_49833,N_40927,N_41617);
nand U49834 (N_49834,N_43181,N_40519);
nand U49835 (N_49835,N_43601,N_41442);
or U49836 (N_49836,N_40899,N_41173);
nor U49837 (N_49837,N_44627,N_43132);
nand U49838 (N_49838,N_42215,N_42538);
nand U49839 (N_49839,N_44816,N_43530);
or U49840 (N_49840,N_42197,N_41058);
and U49841 (N_49841,N_44436,N_43563);
or U49842 (N_49842,N_44088,N_44449);
xnor U49843 (N_49843,N_40044,N_44709);
and U49844 (N_49844,N_40616,N_40034);
or U49845 (N_49845,N_41357,N_42859);
or U49846 (N_49846,N_43677,N_42468);
or U49847 (N_49847,N_44917,N_43955);
and U49848 (N_49848,N_43248,N_44865);
nor U49849 (N_49849,N_41170,N_40360);
xor U49850 (N_49850,N_42670,N_43214);
nand U49851 (N_49851,N_42160,N_40476);
nor U49852 (N_49852,N_41054,N_44299);
nor U49853 (N_49853,N_41581,N_43652);
xnor U49854 (N_49854,N_44482,N_43079);
nor U49855 (N_49855,N_44159,N_42848);
xnor U49856 (N_49856,N_44798,N_41447);
xor U49857 (N_49857,N_42659,N_43184);
nor U49858 (N_49858,N_43647,N_40941);
nand U49859 (N_49859,N_43655,N_40668);
nor U49860 (N_49860,N_41210,N_40517);
nand U49861 (N_49861,N_42583,N_42336);
nand U49862 (N_49862,N_40129,N_42283);
or U49863 (N_49863,N_40016,N_42508);
or U49864 (N_49864,N_43239,N_43328);
or U49865 (N_49865,N_43705,N_43800);
or U49866 (N_49866,N_42767,N_43167);
or U49867 (N_49867,N_42028,N_42891);
nor U49868 (N_49868,N_42880,N_42177);
nor U49869 (N_49869,N_44975,N_43127);
nor U49870 (N_49870,N_43529,N_43932);
and U49871 (N_49871,N_41646,N_43163);
or U49872 (N_49872,N_43975,N_41640);
nor U49873 (N_49873,N_43560,N_42298);
nand U49874 (N_49874,N_42263,N_43484);
nor U49875 (N_49875,N_42509,N_44600);
xnor U49876 (N_49876,N_40364,N_43440);
and U49877 (N_49877,N_40020,N_43675);
nor U49878 (N_49878,N_43560,N_44918);
nand U49879 (N_49879,N_43164,N_41987);
xnor U49880 (N_49880,N_40062,N_43710);
or U49881 (N_49881,N_43899,N_44393);
nand U49882 (N_49882,N_42650,N_40122);
nor U49883 (N_49883,N_44268,N_41090);
nand U49884 (N_49884,N_41427,N_44697);
xor U49885 (N_49885,N_44268,N_41235);
nand U49886 (N_49886,N_42279,N_44890);
xnor U49887 (N_49887,N_43647,N_43040);
and U49888 (N_49888,N_43478,N_44320);
and U49889 (N_49889,N_40032,N_42315);
or U49890 (N_49890,N_44811,N_42375);
nand U49891 (N_49891,N_41670,N_43645);
nor U49892 (N_49892,N_41224,N_44550);
nor U49893 (N_49893,N_43979,N_43935);
nor U49894 (N_49894,N_43812,N_42266);
nor U49895 (N_49895,N_40806,N_42387);
or U49896 (N_49896,N_40197,N_40247);
nand U49897 (N_49897,N_44062,N_41922);
or U49898 (N_49898,N_42322,N_41796);
nor U49899 (N_49899,N_43740,N_44527);
nand U49900 (N_49900,N_43110,N_40834);
nand U49901 (N_49901,N_41698,N_40915);
or U49902 (N_49902,N_42014,N_41778);
nand U49903 (N_49903,N_42311,N_42511);
and U49904 (N_49904,N_40013,N_40499);
nand U49905 (N_49905,N_41073,N_42784);
xor U49906 (N_49906,N_40644,N_40430);
and U49907 (N_49907,N_40578,N_42846);
nor U49908 (N_49908,N_42826,N_44585);
nand U49909 (N_49909,N_42475,N_43560);
nand U49910 (N_49910,N_41120,N_41853);
or U49911 (N_49911,N_42248,N_40830);
or U49912 (N_49912,N_43332,N_42648);
xor U49913 (N_49913,N_41857,N_44967);
nand U49914 (N_49914,N_43246,N_44792);
and U49915 (N_49915,N_40279,N_41789);
xor U49916 (N_49916,N_44734,N_43305);
or U49917 (N_49917,N_42709,N_44946);
nor U49918 (N_49918,N_43673,N_40092);
nor U49919 (N_49919,N_44813,N_42960);
nand U49920 (N_49920,N_41181,N_43247);
or U49921 (N_49921,N_42142,N_41931);
and U49922 (N_49922,N_42529,N_41720);
xor U49923 (N_49923,N_44320,N_44455);
nand U49924 (N_49924,N_41901,N_43208);
and U49925 (N_49925,N_41499,N_40390);
and U49926 (N_49926,N_44501,N_44398);
nor U49927 (N_49927,N_44749,N_43484);
nor U49928 (N_49928,N_43863,N_40381);
and U49929 (N_49929,N_40330,N_42699);
nor U49930 (N_49930,N_42137,N_41685);
nand U49931 (N_49931,N_41958,N_43717);
nor U49932 (N_49932,N_42793,N_42729);
nand U49933 (N_49933,N_44558,N_41423);
xor U49934 (N_49934,N_43038,N_44992);
or U49935 (N_49935,N_44214,N_40143);
and U49936 (N_49936,N_43794,N_43148);
and U49937 (N_49937,N_41136,N_44163);
or U49938 (N_49938,N_40618,N_41379);
nor U49939 (N_49939,N_44236,N_44075);
and U49940 (N_49940,N_41841,N_41979);
or U49941 (N_49941,N_40279,N_42982);
nor U49942 (N_49942,N_42152,N_41050);
nor U49943 (N_49943,N_43477,N_43751);
and U49944 (N_49944,N_41669,N_42041);
or U49945 (N_49945,N_44732,N_42376);
nand U49946 (N_49946,N_42369,N_42886);
and U49947 (N_49947,N_41352,N_44504);
nand U49948 (N_49948,N_42402,N_43246);
nor U49949 (N_49949,N_44387,N_42950);
nand U49950 (N_49950,N_41124,N_41595);
xnor U49951 (N_49951,N_40380,N_43885);
and U49952 (N_49952,N_43907,N_44391);
nand U49953 (N_49953,N_40332,N_40584);
nand U49954 (N_49954,N_42660,N_40260);
nand U49955 (N_49955,N_40632,N_40282);
nand U49956 (N_49956,N_43067,N_43326);
and U49957 (N_49957,N_41565,N_43315);
nand U49958 (N_49958,N_42935,N_40961);
nand U49959 (N_49959,N_43135,N_44697);
nand U49960 (N_49960,N_41828,N_41453);
nor U49961 (N_49961,N_43081,N_43706);
nor U49962 (N_49962,N_42115,N_40171);
or U49963 (N_49963,N_40292,N_44373);
or U49964 (N_49964,N_44262,N_44113);
and U49965 (N_49965,N_42236,N_43632);
nand U49966 (N_49966,N_43683,N_44632);
or U49967 (N_49967,N_40802,N_40536);
xnor U49968 (N_49968,N_41569,N_43856);
nor U49969 (N_49969,N_42029,N_42450);
nor U49970 (N_49970,N_44182,N_44207);
nand U49971 (N_49971,N_42537,N_43750);
nand U49972 (N_49972,N_40558,N_43790);
nand U49973 (N_49973,N_41049,N_41346);
nor U49974 (N_49974,N_42633,N_43191);
or U49975 (N_49975,N_44827,N_41827);
or U49976 (N_49976,N_42794,N_44597);
or U49977 (N_49977,N_41817,N_42916);
and U49978 (N_49978,N_42112,N_40471);
or U49979 (N_49979,N_44598,N_40142);
nand U49980 (N_49980,N_42965,N_43247);
and U49981 (N_49981,N_42515,N_40157);
nand U49982 (N_49982,N_40518,N_43356);
or U49983 (N_49983,N_43360,N_44606);
and U49984 (N_49984,N_44387,N_42645);
nor U49985 (N_49985,N_41239,N_42121);
nor U49986 (N_49986,N_40435,N_42060);
nand U49987 (N_49987,N_41183,N_41382);
or U49988 (N_49988,N_43293,N_41702);
or U49989 (N_49989,N_44750,N_44078);
nor U49990 (N_49990,N_44085,N_40509);
and U49991 (N_49991,N_42264,N_41325);
xnor U49992 (N_49992,N_42045,N_40948);
and U49993 (N_49993,N_43861,N_43438);
nor U49994 (N_49994,N_42642,N_43438);
nand U49995 (N_49995,N_42451,N_44106);
nor U49996 (N_49996,N_41157,N_44468);
nand U49997 (N_49997,N_42718,N_44723);
nor U49998 (N_49998,N_41709,N_40161);
nand U49999 (N_49999,N_40171,N_40944);
or UO_0 (O_0,N_47599,N_47549);
nor UO_1 (O_1,N_48649,N_49761);
nor UO_2 (O_2,N_45682,N_45672);
xor UO_3 (O_3,N_46904,N_49784);
or UO_4 (O_4,N_46040,N_49732);
nor UO_5 (O_5,N_48993,N_49988);
nand UO_6 (O_6,N_46277,N_45983);
nand UO_7 (O_7,N_49886,N_47334);
nor UO_8 (O_8,N_47193,N_48684);
xnor UO_9 (O_9,N_46764,N_48417);
and UO_10 (O_10,N_45918,N_47878);
nand UO_11 (O_11,N_46418,N_47881);
nand UO_12 (O_12,N_46821,N_47759);
nand UO_13 (O_13,N_46987,N_46025);
nand UO_14 (O_14,N_49464,N_45778);
xnor UO_15 (O_15,N_47895,N_46725);
and UO_16 (O_16,N_46644,N_49891);
nand UO_17 (O_17,N_46034,N_46107);
nor UO_18 (O_18,N_49984,N_46917);
xor UO_19 (O_19,N_49162,N_45388);
nor UO_20 (O_20,N_48552,N_48999);
nand UO_21 (O_21,N_48835,N_46640);
nand UO_22 (O_22,N_49963,N_49204);
and UO_23 (O_23,N_46466,N_49830);
nor UO_24 (O_24,N_49871,N_45344);
nand UO_25 (O_25,N_48168,N_48010);
nand UO_26 (O_26,N_45158,N_46355);
nand UO_27 (O_27,N_49471,N_47966);
or UO_28 (O_28,N_48498,N_46512);
or UO_29 (O_29,N_45600,N_46125);
nor UO_30 (O_30,N_47134,N_45591);
or UO_31 (O_31,N_47150,N_45973);
nor UO_32 (O_32,N_46656,N_49236);
nor UO_33 (O_33,N_48695,N_48826);
nor UO_34 (O_34,N_49759,N_46063);
or UO_35 (O_35,N_46488,N_45130);
and UO_36 (O_36,N_48917,N_48584);
nand UO_37 (O_37,N_47489,N_45382);
nor UO_38 (O_38,N_46704,N_47924);
or UO_39 (O_39,N_45022,N_48182);
or UO_40 (O_40,N_49645,N_47778);
and UO_41 (O_41,N_46156,N_46915);
or UO_42 (O_42,N_48633,N_48631);
or UO_43 (O_43,N_46619,N_49073);
and UO_44 (O_44,N_47686,N_45222);
nor UO_45 (O_45,N_46335,N_46455);
xnor UO_46 (O_46,N_49509,N_46302);
or UO_47 (O_47,N_49198,N_47927);
xor UO_48 (O_48,N_46187,N_47469);
or UO_49 (O_49,N_48735,N_45792);
nor UO_50 (O_50,N_47710,N_45034);
nand UO_51 (O_51,N_46627,N_46651);
nor UO_52 (O_52,N_45519,N_48200);
xor UO_53 (O_53,N_48817,N_47561);
or UO_54 (O_54,N_46555,N_45385);
or UO_55 (O_55,N_45796,N_48583);
or UO_56 (O_56,N_47567,N_47975);
nor UO_57 (O_57,N_49630,N_47991);
xor UO_58 (O_58,N_48858,N_46816);
or UO_59 (O_59,N_45744,N_48592);
xor UO_60 (O_60,N_47220,N_49681);
or UO_61 (O_61,N_45430,N_49866);
xnor UO_62 (O_62,N_45096,N_45131);
or UO_63 (O_63,N_45989,N_49373);
and UO_64 (O_64,N_46007,N_48230);
nand UO_65 (O_65,N_46090,N_47266);
nor UO_66 (O_66,N_49102,N_49133);
and UO_67 (O_67,N_47781,N_45758);
nand UO_68 (O_68,N_45129,N_49975);
or UO_69 (O_69,N_49539,N_48074);
xnor UO_70 (O_70,N_46254,N_48945);
and UO_71 (O_71,N_46606,N_49206);
or UO_72 (O_72,N_48235,N_45785);
or UO_73 (O_73,N_47641,N_47373);
nor UO_74 (O_74,N_46210,N_46120);
nand UO_75 (O_75,N_48034,N_48895);
or UO_76 (O_76,N_46127,N_48832);
nand UO_77 (O_77,N_46909,N_47337);
nor UO_78 (O_78,N_47733,N_46746);
or UO_79 (O_79,N_49309,N_49483);
and UO_80 (O_80,N_49056,N_49097);
or UO_81 (O_81,N_45482,N_46085);
and UO_82 (O_82,N_45206,N_46133);
xnor UO_83 (O_83,N_49864,N_46828);
or UO_84 (O_84,N_48605,N_48171);
or UO_85 (O_85,N_46486,N_45243);
or UO_86 (O_86,N_45802,N_48717);
xnor UO_87 (O_87,N_45146,N_45378);
xor UO_88 (O_88,N_47069,N_46345);
or UO_89 (O_89,N_46485,N_47465);
nand UO_90 (O_90,N_48428,N_45551);
nand UO_91 (O_91,N_47956,N_47973);
and UO_92 (O_92,N_49424,N_46883);
nor UO_93 (O_93,N_49149,N_45756);
or UO_94 (O_94,N_47533,N_45358);
and UO_95 (O_95,N_47617,N_46944);
or UO_96 (O_96,N_46313,N_46172);
nor UO_97 (O_97,N_48862,N_45760);
or UO_98 (O_98,N_46255,N_49142);
and UO_99 (O_99,N_46557,N_48956);
nand UO_100 (O_100,N_46093,N_47814);
or UO_101 (O_101,N_47718,N_49797);
nor UO_102 (O_102,N_45850,N_46657);
nor UO_103 (O_103,N_45588,N_48547);
or UO_104 (O_104,N_46241,N_46011);
and UO_105 (O_105,N_47873,N_47809);
xnor UO_106 (O_106,N_47464,N_45687);
nor UO_107 (O_107,N_46398,N_48914);
or UO_108 (O_108,N_48921,N_47245);
nand UO_109 (O_109,N_45263,N_45090);
nor UO_110 (O_110,N_46042,N_48276);
or UO_111 (O_111,N_49333,N_49846);
nor UO_112 (O_112,N_46267,N_45091);
or UO_113 (O_113,N_45714,N_47003);
nor UO_114 (O_114,N_48787,N_48983);
xnor UO_115 (O_115,N_46033,N_46899);
nor UO_116 (O_116,N_47648,N_49092);
nand UO_117 (O_117,N_49727,N_46414);
or UO_118 (O_118,N_48431,N_45543);
nor UO_119 (O_119,N_49958,N_47278);
nand UO_120 (O_120,N_45992,N_48282);
nor UO_121 (O_121,N_46896,N_47195);
or UO_122 (O_122,N_48432,N_47336);
and UO_123 (O_123,N_47537,N_46213);
nand UO_124 (O_124,N_48634,N_48868);
nand UO_125 (O_125,N_47925,N_48941);
nor UO_126 (O_126,N_49752,N_45638);
xor UO_127 (O_127,N_49881,N_49240);
or UO_128 (O_128,N_49554,N_46908);
nor UO_129 (O_129,N_48725,N_47139);
nor UO_130 (O_130,N_45563,N_47044);
or UO_131 (O_131,N_46248,N_46989);
or UO_132 (O_132,N_46684,N_46434);
nand UO_133 (O_133,N_48389,N_49691);
nand UO_134 (O_134,N_45401,N_48121);
nand UO_135 (O_135,N_46715,N_46779);
and UO_136 (O_136,N_48287,N_45320);
nand UO_137 (O_137,N_47971,N_47581);
and UO_138 (O_138,N_46312,N_48091);
xor UO_139 (O_139,N_49129,N_47214);
nor UO_140 (O_140,N_46551,N_49716);
nand UO_141 (O_141,N_48032,N_49758);
xnor UO_142 (O_142,N_45287,N_49628);
nor UO_143 (O_143,N_46641,N_47661);
and UO_144 (O_144,N_47328,N_48562);
or UO_145 (O_145,N_45587,N_47673);
nand UO_146 (O_146,N_46538,N_46785);
nor UO_147 (O_147,N_46667,N_47777);
nand UO_148 (O_148,N_45311,N_45858);
and UO_149 (O_149,N_47452,N_49640);
nand UO_150 (O_150,N_46101,N_45979);
nor UO_151 (O_151,N_49100,N_48071);
and UO_152 (O_152,N_46502,N_47346);
nor UO_153 (O_153,N_46415,N_45408);
nand UO_154 (O_154,N_45708,N_48775);
or UO_155 (O_155,N_47575,N_48643);
and UO_156 (O_156,N_47475,N_45295);
or UO_157 (O_157,N_49955,N_49754);
and UO_158 (O_158,N_45377,N_46868);
or UO_159 (O_159,N_47590,N_48095);
and UO_160 (O_160,N_45361,N_45655);
and UO_161 (O_161,N_47815,N_46546);
nand UO_162 (O_162,N_49485,N_49633);
nand UO_163 (O_163,N_49592,N_48240);
nand UO_164 (O_164,N_45380,N_45322);
and UO_165 (O_165,N_48163,N_46996);
nor UO_166 (O_166,N_46013,N_49989);
and UO_167 (O_167,N_49232,N_48384);
nand UO_168 (O_168,N_46349,N_46372);
nor UO_169 (O_169,N_45530,N_49636);
and UO_170 (O_170,N_46479,N_47384);
nand UO_171 (O_171,N_49532,N_47841);
nand UO_172 (O_172,N_47622,N_49831);
and UO_173 (O_173,N_46561,N_49849);
and UO_174 (O_174,N_45610,N_49012);
nand UO_175 (O_175,N_47602,N_45908);
xnor UO_176 (O_176,N_45168,N_47845);
or UO_177 (O_177,N_45851,N_46665);
or UO_178 (O_178,N_48538,N_45447);
nor UO_179 (O_179,N_47058,N_48535);
and UO_180 (O_180,N_46597,N_46648);
or UO_181 (O_181,N_48679,N_47591);
and UO_182 (O_182,N_48724,N_46171);
and UO_183 (O_183,N_49036,N_45968);
nor UO_184 (O_184,N_48000,N_48064);
or UO_185 (O_185,N_49230,N_45808);
xnor UO_186 (O_186,N_47912,N_48756);
and UO_187 (O_187,N_49480,N_48776);
nor UO_188 (O_188,N_46795,N_47621);
nor UO_189 (O_189,N_47577,N_45095);
and UO_190 (O_190,N_46921,N_45565);
nand UO_191 (O_191,N_46450,N_46406);
nor UO_192 (O_192,N_47920,N_49974);
and UO_193 (O_193,N_46198,N_47664);
or UO_194 (O_194,N_47131,N_47172);
and UO_195 (O_195,N_48516,N_48117);
or UO_196 (O_196,N_46006,N_46189);
nor UO_197 (O_197,N_48310,N_48434);
and UO_198 (O_198,N_49644,N_47541);
nand UO_199 (O_199,N_45703,N_45293);
nand UO_200 (O_200,N_46226,N_48124);
or UO_201 (O_201,N_48228,N_45170);
nand UO_202 (O_202,N_49621,N_45470);
and UO_203 (O_203,N_47862,N_48367);
nand UO_204 (O_204,N_47800,N_48707);
xor UO_205 (O_205,N_49283,N_45728);
and UO_206 (O_206,N_47163,N_47649);
nand UO_207 (O_207,N_47199,N_47851);
nand UO_208 (O_208,N_49419,N_46065);
or UO_209 (O_209,N_47442,N_47053);
nor UO_210 (O_210,N_47239,N_45451);
or UO_211 (O_211,N_49577,N_48073);
or UO_212 (O_212,N_46353,N_45546);
or UO_213 (O_213,N_47268,N_45435);
and UO_214 (O_214,N_46519,N_45651);
or UO_215 (O_215,N_45348,N_49346);
nor UO_216 (O_216,N_45313,N_49626);
nor UO_217 (O_217,N_45173,N_45794);
xor UO_218 (O_218,N_47834,N_48588);
or UO_219 (O_219,N_46338,N_47564);
xnor UO_220 (O_220,N_47688,N_47883);
xor UO_221 (O_221,N_46926,N_49513);
or UO_222 (O_222,N_45337,N_46762);
xor UO_223 (O_223,N_49153,N_46977);
xor UO_224 (O_224,N_47740,N_46283);
and UO_225 (O_225,N_48167,N_47273);
xnor UO_226 (O_226,N_49748,N_46811);
nand UO_227 (O_227,N_48852,N_47595);
xor UO_228 (O_228,N_48100,N_48386);
and UO_229 (O_229,N_45357,N_47116);
or UO_230 (O_230,N_46583,N_45192);
xor UO_231 (O_231,N_48648,N_46492);
and UO_232 (O_232,N_45428,N_47780);
xor UO_233 (O_233,N_48352,N_48833);
and UO_234 (O_234,N_46276,N_46686);
nor UO_235 (O_235,N_48493,N_45353);
or UO_236 (O_236,N_47856,N_45548);
nand UO_237 (O_237,N_46882,N_45406);
or UO_238 (O_238,N_45272,N_47510);
nand UO_239 (O_239,N_45120,N_49550);
xnor UO_240 (O_240,N_47865,N_47518);
xor UO_241 (O_241,N_49120,N_47506);
nand UO_242 (O_242,N_48441,N_48258);
nand UO_243 (O_243,N_49410,N_45397);
or UO_244 (O_244,N_49132,N_45869);
nor UO_245 (O_245,N_47093,N_46251);
nand UO_246 (O_246,N_49286,N_45103);
nor UO_247 (O_247,N_48654,N_47863);
nand UO_248 (O_248,N_48264,N_45070);
nor UO_249 (O_249,N_45661,N_45880);
or UO_250 (O_250,N_49937,N_47939);
nor UO_251 (O_251,N_49836,N_45038);
and UO_252 (O_252,N_47747,N_48655);
and UO_253 (O_253,N_46885,N_49816);
and UO_254 (O_254,N_47584,N_49319);
and UO_255 (O_255,N_46881,N_45152);
xnor UO_256 (O_256,N_46878,N_46293);
nand UO_257 (O_257,N_45019,N_47000);
and UO_258 (O_258,N_45885,N_45855);
nor UO_259 (O_259,N_47766,N_48120);
nor UO_260 (O_260,N_48323,N_46887);
or UO_261 (O_261,N_49391,N_47704);
nor UO_262 (O_262,N_48901,N_48334);
and UO_263 (O_263,N_46717,N_49562);
nand UO_264 (O_264,N_49794,N_45485);
nand UO_265 (O_265,N_46253,N_46716);
nand UO_266 (O_266,N_46559,N_45440);
nor UO_267 (O_267,N_45912,N_46257);
and UO_268 (O_268,N_48070,N_48361);
or UO_269 (O_269,N_47548,N_49436);
nand UO_270 (O_270,N_47596,N_48873);
nor UO_271 (O_271,N_47158,N_48140);
nor UO_272 (O_272,N_48995,N_46945);
or UO_273 (O_273,N_49903,N_45659);
nor UO_274 (O_274,N_47663,N_49964);
and UO_275 (O_275,N_47821,N_45788);
nor UO_276 (O_276,N_49750,N_48006);
and UO_277 (O_277,N_49641,N_49468);
or UO_278 (O_278,N_46736,N_49940);
and UO_279 (O_279,N_47221,N_46131);
and UO_280 (O_280,N_49725,N_46015);
or UO_281 (O_281,N_46815,N_47657);
and UO_282 (O_282,N_46081,N_45167);
xnor UO_283 (O_283,N_49247,N_48730);
or UO_284 (O_284,N_49529,N_49452);
or UO_285 (O_285,N_48878,N_48482);
nor UO_286 (O_286,N_47887,N_49388);
nor UO_287 (O_287,N_45270,N_45066);
or UO_288 (O_288,N_49445,N_46083);
nor UO_289 (O_289,N_49163,N_48532);
nand UO_290 (O_290,N_49067,N_49598);
nor UO_291 (O_291,N_49269,N_45474);
nor UO_292 (O_292,N_45073,N_45278);
or UO_293 (O_293,N_48785,N_47007);
or UO_294 (O_294,N_48269,N_49001);
nand UO_295 (O_295,N_48906,N_47313);
xor UO_296 (O_296,N_45372,N_46838);
nand UO_297 (O_297,N_47418,N_46625);
or UO_298 (O_298,N_48700,N_49858);
nand UO_299 (O_299,N_48030,N_48143);
nor UO_300 (O_300,N_49345,N_45685);
nand UO_301 (O_301,N_46316,N_47324);
nor UO_302 (O_302,N_49684,N_45631);
or UO_303 (O_303,N_47751,N_49608);
xnor UO_304 (O_304,N_45843,N_47232);
nor UO_305 (O_305,N_48455,N_48626);
or UO_306 (O_306,N_49216,N_49257);
nor UO_307 (O_307,N_48561,N_45284);
nor UO_308 (O_308,N_49076,N_46347);
and UO_309 (O_309,N_48677,N_47121);
or UO_310 (O_310,N_48273,N_47762);
and UO_311 (O_311,N_47035,N_49173);
or UO_312 (O_312,N_47861,N_45697);
or UO_313 (O_313,N_45327,N_47600);
xnor UO_314 (O_314,N_47919,N_48297);
nor UO_315 (O_315,N_45571,N_47329);
and UO_316 (O_316,N_47258,N_47372);
nand UO_317 (O_317,N_46928,N_46537);
and UO_318 (O_318,N_48861,N_46028);
and UO_319 (O_319,N_46884,N_45352);
xnor UO_320 (O_320,N_47047,N_47285);
nand UO_321 (O_321,N_49826,N_46106);
nor UO_322 (O_322,N_46853,N_46339);
nand UO_323 (O_323,N_48129,N_47793);
xor UO_324 (O_324,N_45314,N_45879);
and UO_325 (O_325,N_48157,N_46258);
and UO_326 (O_326,N_45411,N_48514);
nand UO_327 (O_327,N_48439,N_45305);
nor UO_328 (O_328,N_47619,N_46818);
and UO_329 (O_329,N_46201,N_45394);
nor UO_330 (O_330,N_48736,N_47011);
nor UO_331 (O_331,N_46966,N_47957);
nor UO_332 (O_332,N_45585,N_46721);
and UO_333 (O_333,N_45472,N_46023);
or UO_334 (O_334,N_46491,N_47536);
nor UO_335 (O_335,N_45508,N_49088);
or UO_336 (O_336,N_47060,N_49046);
nand UO_337 (O_337,N_46672,N_49602);
and UO_338 (O_338,N_45139,N_49544);
nand UO_339 (O_339,N_47931,N_47036);
nor UO_340 (O_340,N_49209,N_46786);
nand UO_341 (O_341,N_48748,N_48714);
or UO_342 (O_342,N_47752,N_47148);
nand UO_343 (O_343,N_47909,N_46741);
nor UO_344 (O_344,N_49774,N_46370);
and UO_345 (O_345,N_46906,N_48198);
nor UO_346 (O_346,N_45198,N_47910);
xor UO_347 (O_347,N_48892,N_45230);
nand UO_348 (O_348,N_49276,N_46021);
nor UO_349 (O_349,N_49938,N_48250);
and UO_350 (O_350,N_48824,N_48027);
nor UO_351 (O_351,N_45200,N_49508);
xor UO_352 (O_352,N_47198,N_48078);
or UO_353 (O_353,N_48268,N_49946);
xor UO_354 (O_354,N_46054,N_48982);
and UO_355 (O_355,N_48279,N_48666);
and UO_356 (O_356,N_48485,N_45718);
and UO_357 (O_357,N_45975,N_46582);
and UO_358 (O_358,N_47070,N_45183);
or UO_359 (O_359,N_45569,N_46891);
and UO_360 (O_360,N_45861,N_48739);
nand UO_361 (O_361,N_48313,N_49907);
nor UO_362 (O_362,N_49859,N_49025);
nor UO_363 (O_363,N_45684,N_48587);
nand UO_364 (O_364,N_48507,N_45241);
and UO_365 (O_365,N_49800,N_49540);
or UO_366 (O_366,N_49870,N_48019);
nor UO_367 (O_367,N_49069,N_47553);
and UO_368 (O_368,N_48769,N_46150);
nor UO_369 (O_369,N_49143,N_47106);
nor UO_370 (O_370,N_46529,N_48663);
nand UO_371 (O_371,N_48308,N_48497);
nand UO_372 (O_372,N_48068,N_49459);
or UO_373 (O_373,N_45719,N_47297);
and UO_374 (O_374,N_47120,N_47430);
xor UO_375 (O_375,N_49809,N_46104);
nand UO_376 (O_376,N_48871,N_47043);
nor UO_377 (O_377,N_48363,N_49837);
or UO_378 (O_378,N_49087,N_46751);
nand UO_379 (O_379,N_45823,N_48151);
nor UO_380 (O_380,N_47932,N_45627);
and UO_381 (O_381,N_47226,N_45537);
xor UO_382 (O_382,N_47374,N_46634);
nand UO_383 (O_383,N_49901,N_49446);
and UO_384 (O_384,N_47331,N_46074);
nand UO_385 (O_385,N_46279,N_48162);
nor UO_386 (O_386,N_49358,N_46870);
nor UO_387 (O_387,N_49953,N_48123);
or UO_388 (O_388,N_49293,N_45265);
or UO_389 (O_389,N_48454,N_47321);
or UO_390 (O_390,N_49998,N_45902);
nor UO_391 (O_391,N_47946,N_48238);
or UO_392 (O_392,N_46413,N_47213);
xnor UO_393 (O_393,N_49364,N_49976);
nand UO_394 (O_394,N_49245,N_49611);
nand UO_395 (O_395,N_45803,N_46206);
or UO_396 (O_396,N_47715,N_45498);
and UO_397 (O_397,N_47354,N_48533);
nand UO_398 (O_398,N_47259,N_47967);
nor UO_399 (O_399,N_49743,N_45877);
nor UO_400 (O_400,N_49267,N_48590);
and UO_401 (O_401,N_45653,N_45478);
nor UO_402 (O_402,N_48630,N_48150);
nor UO_403 (O_403,N_45824,N_45196);
or UO_404 (O_404,N_48551,N_47359);
nand UO_405 (O_405,N_47791,N_46427);
and UO_406 (O_406,N_47059,N_46620);
and UO_407 (O_407,N_48373,N_49880);
and UO_408 (O_408,N_45298,N_45942);
nand UO_409 (O_409,N_48261,N_48412);
or UO_410 (O_410,N_49655,N_47155);
and UO_411 (O_411,N_49710,N_45024);
or UO_412 (O_412,N_46673,N_45874);
and UO_413 (O_413,N_49217,N_48734);
nand UO_414 (O_414,N_46389,N_45257);
and UO_415 (O_415,N_47667,N_46941);
nand UO_416 (O_416,N_47170,N_45807);
xnor UO_417 (O_417,N_48368,N_48328);
and UO_418 (O_418,N_45547,N_47065);
nor UO_419 (O_419,N_46790,N_45110);
nor UO_420 (O_420,N_49574,N_48229);
nand UO_421 (O_421,N_47654,N_48615);
or UO_422 (O_422,N_46742,N_48499);
nand UO_423 (O_423,N_45396,N_49768);
or UO_424 (O_424,N_46831,N_47787);
nand UO_425 (O_425,N_46278,N_49737);
or UO_426 (O_426,N_46523,N_45817);
nor UO_427 (O_427,N_46628,N_48608);
nor UO_428 (O_428,N_47795,N_48336);
and UO_429 (O_429,N_48476,N_46348);
or UO_430 (O_430,N_46117,N_49549);
or UO_431 (O_431,N_47246,N_45643);
and UO_432 (O_432,N_46056,N_45893);
and UO_433 (O_433,N_47128,N_45267);
or UO_434 (O_434,N_49028,N_46315);
xnor UO_435 (O_435,N_45087,N_49004);
or UO_436 (O_436,N_47698,N_48622);
and UO_437 (O_437,N_46985,N_46140);
xnor UO_438 (O_438,N_47938,N_47414);
nor UO_439 (O_439,N_48620,N_49488);
nand UO_440 (O_440,N_47251,N_45233);
nand UO_441 (O_441,N_49924,N_46393);
nand UO_442 (O_442,N_47524,N_48281);
nand UO_443 (O_443,N_46378,N_47560);
or UO_444 (O_444,N_45692,N_47243);
and UO_445 (O_445,N_47831,N_45738);
nand UO_446 (O_446,N_49458,N_47869);
nor UO_447 (O_447,N_49160,N_49141);
xnor UO_448 (O_448,N_45012,N_49921);
nor UO_449 (O_449,N_48968,N_46281);
xor UO_450 (O_450,N_45189,N_49020);
nand UO_451 (O_451,N_48502,N_48043);
xnor UO_452 (O_452,N_48192,N_47257);
or UO_453 (O_453,N_45938,N_48761);
or UO_454 (O_454,N_45504,N_49631);
or UO_455 (O_455,N_47828,N_45341);
nor UO_456 (O_456,N_45641,N_46699);
nor UO_457 (O_457,N_48844,N_48733);
or UO_458 (O_458,N_48014,N_49987);
nand UO_459 (O_459,N_47992,N_48395);
nor UO_460 (O_460,N_49791,N_45321);
nand UO_461 (O_461,N_49895,N_45094);
and UO_462 (O_462,N_49499,N_45705);
nor UO_463 (O_463,N_45354,N_47314);
nand UO_464 (O_464,N_47725,N_47377);
nand UO_465 (O_465,N_45391,N_47731);
and UO_466 (O_466,N_47703,N_45882);
or UO_467 (O_467,N_47854,N_45424);
nand UO_468 (O_468,N_48789,N_46032);
nand UO_469 (O_469,N_47225,N_45201);
or UO_470 (O_470,N_47849,N_45619);
xnor UO_471 (O_471,N_49706,N_47995);
nor UO_472 (O_472,N_48042,N_45965);
or UO_473 (O_473,N_45266,N_46144);
or UO_474 (O_474,N_49158,N_46859);
and UO_475 (O_475,N_49000,N_48191);
nor UO_476 (O_476,N_48480,N_49969);
nand UO_477 (O_477,N_49646,N_45667);
nor UO_478 (O_478,N_48948,N_48097);
nand UO_479 (O_479,N_47391,N_49049);
xor UO_480 (O_480,N_48029,N_45870);
or UO_481 (O_481,N_45828,N_47889);
or UO_482 (O_482,N_46431,N_46708);
xor UO_483 (O_483,N_46473,N_45590);
xnor UO_484 (O_484,N_48357,N_49270);
xor UO_485 (O_485,N_45507,N_48614);
nor UO_486 (O_486,N_48465,N_45299);
nor UO_487 (O_487,N_46515,N_46739);
or UO_488 (O_488,N_47678,N_45153);
xor UO_489 (O_489,N_48463,N_45015);
nand UO_490 (O_490,N_46452,N_46695);
and UO_491 (O_491,N_45421,N_46540);
or UO_492 (O_492,N_48344,N_46865);
and UO_493 (O_493,N_48773,N_48617);
or UO_494 (O_494,N_48854,N_47392);
nor UO_495 (O_495,N_46128,N_49287);
nor UO_496 (O_496,N_47467,N_49571);
nand UO_497 (O_497,N_48472,N_45499);
nand UO_498 (O_498,N_48996,N_48672);
nand UO_499 (O_499,N_46577,N_46616);
and UO_500 (O_500,N_48184,N_47272);
nor UO_501 (O_501,N_47371,N_47395);
and UO_502 (O_502,N_45510,N_45890);
and UO_503 (O_503,N_49729,N_48098);
nand UO_504 (O_504,N_47990,N_45488);
or UO_505 (O_505,N_45124,N_49022);
and UO_506 (O_506,N_48863,N_46659);
and UO_507 (O_507,N_45252,N_45209);
nor UO_508 (O_508,N_49029,N_49199);
and UO_509 (O_509,N_46802,N_45042);
xor UO_510 (O_510,N_48604,N_47502);
nand UO_511 (O_511,N_49956,N_47015);
nand UO_512 (O_512,N_47933,N_46099);
or UO_513 (O_513,N_45941,N_47741);
or UO_514 (O_514,N_48205,N_49168);
xnor UO_515 (O_515,N_48049,N_46132);
nand UO_516 (O_516,N_49239,N_48138);
and UO_517 (O_517,N_48656,N_48815);
and UO_518 (O_518,N_46436,N_48959);
nor UO_519 (O_519,N_46998,N_46357);
and UO_520 (O_520,N_45202,N_47802);
nand UO_521 (O_521,N_47839,N_49515);
xnor UO_522 (O_522,N_46876,N_46841);
or UO_523 (O_523,N_49847,N_48460);
and UO_524 (O_524,N_46712,N_49190);
xnor UO_525 (O_525,N_46940,N_47159);
nand UO_526 (O_526,N_45645,N_48834);
and UO_527 (O_527,N_45349,N_49438);
nand UO_528 (O_528,N_45141,N_45346);
nor UO_529 (O_529,N_49083,N_47078);
xor UO_530 (O_530,N_48423,N_49527);
and UO_531 (O_531,N_46075,N_47875);
and UO_532 (O_532,N_48188,N_49226);
nor UO_533 (O_533,N_49294,N_46318);
nor UO_534 (O_534,N_47764,N_49212);
and UO_535 (O_535,N_48637,N_48462);
and UO_536 (O_536,N_48011,N_48757);
or UO_537 (O_537,N_48415,N_45193);
nand UO_538 (O_538,N_45678,N_46176);
and UO_539 (O_539,N_49165,N_47864);
nand UO_540 (O_540,N_47668,N_46103);
and UO_541 (O_541,N_48145,N_46527);
or UO_542 (O_542,N_48348,N_45647);
nand UO_543 (O_543,N_46806,N_46680);
xor UO_544 (O_544,N_45525,N_49543);
xnor UO_545 (O_545,N_46602,N_45274);
and UO_546 (O_546,N_45984,N_49802);
or UO_547 (O_547,N_49823,N_49653);
and UO_548 (O_548,N_46775,N_48008);
and UO_549 (O_549,N_49612,N_45669);
or UO_550 (O_550,N_48706,N_46905);
nand UO_551 (O_551,N_47840,N_48541);
and UO_552 (O_552,N_48353,N_49161);
nor UO_553 (O_553,N_48795,N_47633);
or UO_554 (O_554,N_49815,N_48131);
nand UO_555 (O_555,N_47087,N_47707);
nor UO_556 (O_556,N_46873,N_47072);
and UO_557 (O_557,N_48888,N_45520);
nand UO_558 (O_558,N_47737,N_49009);
nand UO_559 (O_559,N_48937,N_47153);
nor UO_560 (O_560,N_45863,N_48744);
or UO_561 (O_561,N_49814,N_49825);
nand UO_562 (O_562,N_48400,N_47355);
or UO_563 (O_563,N_47202,N_48671);
or UO_564 (O_564,N_48572,N_46256);
nand UO_565 (O_565,N_48259,N_46728);
nor UO_566 (O_566,N_45114,N_49344);
and UO_567 (O_567,N_48146,N_48942);
and UO_568 (O_568,N_45921,N_47811);
and UO_569 (O_569,N_46780,N_46542);
or UO_570 (O_570,N_45261,N_48193);
and UO_571 (O_571,N_45497,N_46073);
or UO_572 (O_572,N_46541,N_49429);
and UO_573 (O_573,N_49131,N_48132);
nand UO_574 (O_574,N_47436,N_45336);
or UO_575 (O_575,N_45514,N_49408);
or UO_576 (O_576,N_48437,N_48216);
and UO_577 (O_577,N_48063,N_46967);
xnor UO_578 (O_578,N_49443,N_49365);
nor UO_579 (O_579,N_47262,N_47398);
or UO_580 (O_580,N_47082,N_45674);
xor UO_581 (O_581,N_48044,N_45920);
nor UO_582 (O_582,N_46237,N_48810);
nand UO_583 (O_583,N_46026,N_49994);
or UO_584 (O_584,N_49674,N_45283);
or UO_585 (O_585,N_47568,N_47941);
xnor UO_586 (O_586,N_47525,N_47857);
xnor UO_587 (O_587,N_48084,N_45092);
and UO_588 (O_588,N_47746,N_49561);
and UO_589 (O_589,N_48404,N_45306);
nand UO_590 (O_590,N_49151,N_45089);
nor UO_591 (O_591,N_49548,N_47196);
and UO_592 (O_592,N_47389,N_46982);
or UO_593 (O_593,N_45213,N_45771);
nor UO_594 (O_594,N_45473,N_47269);
nand UO_595 (O_595,N_47680,N_48303);
nand UO_596 (O_596,N_45325,N_49152);
nand UO_597 (O_597,N_48953,N_48926);
and UO_598 (O_598,N_46757,N_47915);
nand UO_599 (O_599,N_49578,N_47025);
or UO_600 (O_600,N_48305,N_49398);
nor UO_601 (O_601,N_48113,N_49297);
or UO_602 (O_602,N_45464,N_47276);
nand UO_603 (O_603,N_45580,N_49547);
and UO_604 (O_604,N_48177,N_49538);
or UO_605 (O_605,N_48822,N_45745);
and UO_606 (O_606,N_49930,N_47642);
nor UO_607 (O_607,N_47645,N_48515);
and UO_608 (O_608,N_47706,N_45560);
nand UO_609 (O_609,N_48378,N_46292);
xnor UO_610 (O_610,N_48952,N_47527);
or UO_611 (O_611,N_45522,N_45021);
nor UO_612 (O_612,N_45556,N_45007);
nand UO_613 (O_613,N_45997,N_47205);
and UO_614 (O_614,N_46988,N_45664);
nor UO_615 (O_615,N_47461,N_48309);
and UO_616 (O_616,N_47112,N_48265);
and UO_617 (O_617,N_48005,N_47643);
and UO_618 (O_618,N_48130,N_48271);
nor UO_619 (O_619,N_45126,N_46965);
nor UO_620 (O_620,N_48758,N_49780);
nor UO_621 (O_621,N_46914,N_46707);
nor UO_622 (O_622,N_46984,N_48424);
and UO_623 (O_623,N_49126,N_46186);
or UO_624 (O_624,N_49546,N_48807);
and UO_625 (O_625,N_49957,N_47001);
and UO_626 (O_626,N_45549,N_45431);
or UO_627 (O_627,N_47056,N_48045);
and UO_628 (O_628,N_45174,N_46211);
or UO_629 (O_629,N_45106,N_47504);
or UO_630 (O_630,N_46810,N_45969);
nor UO_631 (O_631,N_47566,N_49530);
nor UO_632 (O_632,N_48199,N_45704);
xnor UO_633 (O_633,N_47903,N_49356);
and UO_634 (O_634,N_45462,N_47375);
nand UO_635 (O_635,N_49699,N_46911);
nor UO_636 (O_636,N_49195,N_45698);
xnor UO_637 (O_637,N_49031,N_45531);
and UO_638 (O_638,N_45512,N_46191);
nor UO_639 (O_639,N_49308,N_48488);
or UO_640 (O_640,N_47311,N_45539);
nand UO_641 (O_641,N_45212,N_47485);
nand UO_642 (O_642,N_49418,N_47681);
or UO_643 (O_643,N_47094,N_47891);
and UO_644 (O_644,N_47702,N_45301);
nor UO_645 (O_645,N_46861,N_46823);
or UO_646 (O_646,N_45262,N_47726);
or UO_647 (O_647,N_48522,N_47383);
xor UO_648 (O_648,N_45964,N_49449);
or UO_649 (O_649,N_47241,N_49995);
or UO_650 (O_650,N_45848,N_47135);
nand UO_651 (O_651,N_45163,N_49068);
or UO_652 (O_652,N_48595,N_48779);
or UO_653 (O_653,N_45730,N_48893);
and UO_654 (O_654,N_48705,N_47911);
nor UO_655 (O_655,N_49868,N_46461);
and UO_656 (O_656,N_48274,N_45433);
nand UO_657 (O_657,N_47937,N_46192);
xnor UO_658 (O_658,N_49834,N_45323);
nand UO_659 (O_659,N_45300,N_46297);
or UO_660 (O_660,N_47338,N_48886);
or UO_661 (O_661,N_46774,N_46750);
nand UO_662 (O_662,N_48664,N_49861);
and UO_663 (O_663,N_49500,N_49015);
nand UO_664 (O_664,N_47468,N_45273);
or UO_665 (O_665,N_48754,N_45953);
nor UO_666 (O_666,N_49749,N_48716);
and UO_667 (O_667,N_46401,N_47387);
nor UO_668 (O_668,N_49041,N_49227);
and UO_669 (O_669,N_49330,N_49788);
or UO_670 (O_670,N_48185,N_46010);
and UO_671 (O_671,N_47792,N_49374);
nor UO_672 (O_672,N_46138,N_46285);
and UO_673 (O_673,N_49558,N_47368);
nor UO_674 (O_674,N_47360,N_49769);
nand UO_675 (O_675,N_45109,N_49043);
nand UO_676 (O_676,N_47417,N_45706);
xnor UO_677 (O_677,N_46243,N_45621);
nand UO_678 (O_678,N_47008,N_49667);
nor UO_679 (O_679,N_46465,N_47717);
or UO_680 (O_680,N_45415,N_46096);
xnor UO_681 (O_681,N_47625,N_45832);
nor UO_682 (O_682,N_45303,N_45822);
nand UO_683 (O_683,N_45416,N_48164);
or UO_684 (O_684,N_46346,N_47801);
nor UO_685 (O_685,N_45905,N_45691);
nor UO_686 (O_686,N_45132,N_49016);
and UO_687 (O_687,N_45339,N_45916);
and UO_688 (O_688,N_48372,N_46428);
nor UO_689 (O_689,N_49677,N_45988);
xnor UO_690 (O_690,N_45335,N_45294);
nor UO_691 (O_691,N_47123,N_47038);
and UO_692 (O_692,N_48195,N_49496);
nand UO_693 (O_693,N_47289,N_45605);
nor UO_694 (O_694,N_45679,N_49576);
xor UO_695 (O_695,N_47308,N_45936);
and UO_696 (O_696,N_46677,N_49878);
or UO_697 (O_697,N_47624,N_45057);
or UO_698 (O_698,N_45460,N_46307);
nor UO_699 (O_699,N_48461,N_45254);
or UO_700 (O_700,N_45841,N_49511);
and UO_701 (O_701,N_48172,N_48977);
nand UO_702 (O_702,N_49923,N_47608);
nand UO_703 (O_703,N_48907,N_46995);
nand UO_704 (O_704,N_45444,N_49887);
or UO_705 (O_705,N_48981,N_48857);
nor UO_706 (O_706,N_49839,N_47118);
or UO_707 (O_707,N_47413,N_48035);
nor UO_708 (O_708,N_46306,N_45063);
xor UO_709 (O_709,N_46484,N_46204);
nor UO_710 (O_710,N_48718,N_49248);
and UO_711 (O_711,N_47753,N_48877);
nand UO_712 (O_712,N_49627,N_49114);
nand UO_713 (O_713,N_45515,N_47460);
nand UO_714 (O_714,N_47785,N_47034);
or UO_715 (O_715,N_48170,N_49615);
nand UO_716 (O_716,N_46886,N_46380);
nand UO_717 (O_717,N_46678,N_48850);
or UO_718 (O_718,N_45948,N_45943);
nor UO_719 (O_719,N_49139,N_47409);
or UO_720 (O_720,N_45500,N_46260);
nor UO_721 (O_721,N_49589,N_47209);
xor UO_722 (O_722,N_46614,N_45383);
or UO_723 (O_723,N_48911,N_48846);
nor UO_724 (O_724,N_46869,N_46999);
xnor UO_725 (O_725,N_45423,N_49741);
nand UO_726 (O_726,N_45345,N_48089);
or UO_727 (O_727,N_49192,N_48209);
nand UO_728 (O_728,N_49397,N_46747);
nor UO_729 (O_729,N_49740,N_48780);
and UO_730 (O_730,N_48582,N_48266);
or UO_731 (O_731,N_46638,N_48652);
and UO_732 (O_732,N_46740,N_46425);
nand UO_733 (O_733,N_45800,N_47769);
nor UO_734 (O_734,N_45404,N_45449);
nor UO_735 (O_735,N_46671,N_45100);
xnor UO_736 (O_736,N_48984,N_47904);
and UO_737 (O_737,N_48494,N_49763);
and UO_738 (O_738,N_45471,N_49798);
nand UO_739 (O_739,N_48681,N_49035);
or UO_740 (O_740,N_49263,N_48659);
or UO_741 (O_741,N_48467,N_49188);
or UO_742 (O_742,N_46900,N_45575);
xnor UO_743 (O_743,N_45194,N_47124);
xor UO_744 (O_744,N_48116,N_48430);
xor UO_745 (O_745,N_49282,N_47190);
nor UO_746 (O_746,N_49117,N_47972);
nand UO_747 (O_747,N_46396,N_47721);
nand UO_748 (O_748,N_48359,N_47421);
nor UO_749 (O_749,N_46135,N_47361);
nand UO_750 (O_750,N_49591,N_46877);
or UO_751 (O_751,N_49796,N_46799);
or UO_752 (O_752,N_49570,N_48838);
or UO_753 (O_753,N_46758,N_48225);
and UO_754 (O_754,N_47054,N_49805);
nand UO_755 (O_755,N_45518,N_46698);
or UO_756 (O_756,N_47587,N_45169);
xor UO_757 (O_757,N_49916,N_45955);
or UO_758 (O_758,N_48451,N_49516);
and UO_759 (O_759,N_49221,N_46618);
nor UO_760 (O_760,N_46122,N_45809);
or UO_761 (O_761,N_45443,N_46937);
or UO_762 (O_762,N_48223,N_46834);
or UO_763 (O_763,N_46895,N_45523);
nand UO_764 (O_764,N_45597,N_47400);
and UO_765 (O_765,N_49738,N_45442);
nor UO_766 (O_766,N_47088,N_47411);
or UO_767 (O_767,N_46469,N_47394);
nor UO_768 (O_768,N_48054,N_48568);
and UO_769 (O_769,N_49119,N_47606);
xor UO_770 (O_770,N_46164,N_49360);
xnor UO_771 (O_771,N_48174,N_46621);
or UO_772 (O_772,N_46690,N_49137);
xor UO_773 (O_773,N_47495,N_46710);
and UO_774 (O_774,N_46719,N_46992);
nor UO_775 (O_775,N_47825,N_47748);
nand UO_776 (O_776,N_46888,N_45533);
nor UO_777 (O_777,N_46091,N_48453);
and UO_778 (O_778,N_48843,N_45002);
and UO_779 (O_779,N_45052,N_46119);
nor UO_780 (O_780,N_49795,N_46400);
and UO_781 (O_781,N_48237,N_46196);
or UO_782 (O_782,N_47237,N_46696);
nand UO_783 (O_783,N_47913,N_47534);
xor UO_784 (O_784,N_46954,N_45316);
nor UO_785 (O_785,N_48385,N_49882);
nor UO_786 (O_786,N_46729,N_46654);
xnor UO_787 (O_787,N_47526,N_45180);
nand UO_788 (O_788,N_48289,N_49051);
nor UO_789 (O_789,N_47228,N_45524);
or UO_790 (O_790,N_49697,N_48056);
or UO_791 (O_791,N_46874,N_45720);
and UO_792 (O_792,N_46072,N_48676);
nor UO_793 (O_793,N_46317,N_49605);
nand UO_794 (O_794,N_47168,N_49093);
and UO_795 (O_795,N_46272,N_49492);
nand UO_796 (O_796,N_47445,N_47675);
and UO_797 (O_797,N_45368,N_45282);
nand UO_798 (O_798,N_48570,N_45573);
xnor UO_799 (O_799,N_49841,N_48760);
and UO_800 (O_800,N_48413,N_49252);
or UO_801 (O_801,N_48890,N_49298);
and UO_802 (O_802,N_45888,N_45010);
nor UO_803 (O_803,N_47114,N_49523);
nand UO_804 (O_804,N_45892,N_47694);
and UO_805 (O_805,N_46922,N_46748);
nand UO_806 (O_806,N_48211,N_48203);
nor UO_807 (O_807,N_46018,N_47101);
or UO_808 (O_808,N_46296,N_46807);
or UO_809 (O_809,N_49253,N_47415);
xnor UO_810 (O_810,N_45386,N_45650);
and UO_811 (O_811,N_49692,N_46145);
or UO_812 (O_812,N_49472,N_48082);
nor UO_813 (O_813,N_45072,N_46392);
xnor UO_814 (O_814,N_49448,N_48260);
xor UO_815 (O_815,N_49619,N_49183);
and UO_816 (O_816,N_47040,N_46022);
xnor UO_817 (O_817,N_45995,N_45332);
and UO_818 (O_818,N_48632,N_48702);
nand UO_819 (O_819,N_46071,N_46102);
nand UO_820 (O_820,N_47353,N_45977);
nor UO_821 (O_821,N_48445,N_48459);
and UO_822 (O_822,N_48371,N_47773);
and UO_823 (O_823,N_48102,N_46703);
or UO_824 (O_824,N_46794,N_49860);
nand UO_825 (O_825,N_46734,N_46282);
xnor UO_826 (O_826,N_47157,N_46646);
and UO_827 (O_827,N_47129,N_46507);
or UO_828 (O_828,N_45974,N_45179);
or UO_829 (O_829,N_46482,N_46863);
or UO_830 (O_830,N_45023,N_47576);
xnor UO_831 (O_831,N_46217,N_48784);
nand UO_832 (O_832,N_45351,N_47836);
and UO_833 (O_833,N_47563,N_46426);
or UO_834 (O_834,N_49829,N_48537);
and UO_835 (O_835,N_48396,N_48866);
and UO_836 (O_836,N_49191,N_49785);
nor UO_837 (O_837,N_48165,N_47750);
nor UO_838 (O_838,N_46531,N_47071);
or UO_839 (O_839,N_47345,N_45972);
or UO_840 (O_840,N_49134,N_49292);
and UO_841 (O_841,N_49476,N_47265);
and UO_842 (O_842,N_45970,N_48546);
or UO_843 (O_843,N_46483,N_46294);
nand UO_844 (O_844,N_47727,N_49334);
or UO_845 (O_845,N_46956,N_49623);
nand UO_846 (O_846,N_47730,N_46049);
nand UO_847 (O_847,N_48954,N_46441);
nand UO_848 (O_848,N_49904,N_45668);
and UO_849 (O_849,N_49745,N_48919);
nand UO_850 (O_850,N_47640,N_49599);
nor UO_851 (O_851,N_46359,N_48362);
nand UO_852 (O_852,N_49587,N_49075);
and UO_853 (O_853,N_48732,N_46299);
or UO_854 (O_854,N_47294,N_47914);
or UO_855 (O_855,N_48814,N_49896);
and UO_856 (O_856,N_46639,N_45033);
and UO_857 (O_857,N_46649,N_47719);
xor UO_858 (O_858,N_48128,N_45614);
nor UO_859 (O_859,N_47256,N_45636);
and UO_860 (O_860,N_49325,N_46844);
or UO_861 (O_861,N_46978,N_47483);
nand UO_862 (O_862,N_45616,N_48215);
and UO_863 (O_863,N_49403,N_49551);
and UO_864 (O_864,N_48477,N_48985);
nor UO_865 (O_865,N_48242,N_47098);
or UO_866 (O_866,N_46266,N_48998);
nand UO_867 (O_867,N_47646,N_45118);
or UO_868 (O_868,N_45450,N_48311);
or UO_869 (O_869,N_45403,N_49279);
nand UO_870 (O_870,N_47610,N_48031);
nor UO_871 (O_871,N_49624,N_45789);
xor UO_872 (O_872,N_45777,N_48379);
and UO_873 (O_873,N_47396,N_49219);
or UO_874 (O_874,N_49342,N_47367);
or UO_875 (O_875,N_49926,N_48470);
xnor UO_876 (O_876,N_49686,N_46416);
and UO_877 (O_877,N_48178,N_49058);
or UO_878 (O_878,N_48374,N_46756);
nor UO_879 (O_879,N_47550,N_45176);
or UO_880 (O_880,N_49369,N_45429);
nor UO_881 (O_881,N_48206,N_49469);
nor UO_882 (O_882,N_47080,N_49912);
xnor UO_883 (O_883,N_49648,N_49256);
nand UO_884 (O_884,N_48096,N_45887);
or UO_885 (O_885,N_48628,N_48908);
nor UO_886 (O_886,N_48322,N_49575);
and UO_887 (O_887,N_49179,N_47014);
nor UO_888 (O_888,N_49213,N_48913);
nor UO_889 (O_889,N_45220,N_45245);
nor UO_890 (O_890,N_46364,N_48013);
nand UO_891 (O_891,N_47685,N_48646);
nand UO_892 (O_892,N_48601,N_48275);
or UO_893 (O_893,N_47929,N_47890);
or UO_894 (O_894,N_49728,N_46070);
or UO_895 (O_895,N_48550,N_46005);
nand UO_896 (O_896,N_45776,N_49259);
xnor UO_897 (O_897,N_47950,N_49156);
nand UO_898 (O_898,N_47146,N_49560);
and UO_899 (O_899,N_47739,N_49054);
or UO_900 (O_900,N_46303,N_48489);
and UO_901 (O_901,N_46724,N_48107);
xnor UO_902 (O_902,N_46569,N_47630);
and UO_903 (O_903,N_45359,N_45438);
nand UO_904 (O_904,N_46770,N_46141);
or UO_905 (O_905,N_45469,N_46675);
nor UO_906 (O_906,N_47161,N_48081);
nor UO_907 (O_907,N_49447,N_46358);
xnor UO_908 (O_908,N_46932,N_45465);
xor UO_909 (O_909,N_48899,N_46064);
and UO_910 (O_910,N_49996,N_47829);
or UO_911 (O_911,N_49254,N_49872);
nor UO_912 (O_912,N_46566,N_47974);
nor UO_913 (O_913,N_49962,N_45147);
xnor UO_914 (O_914,N_48290,N_46233);
nand UO_915 (O_915,N_45987,N_49382);
nor UO_916 (O_916,N_49047,N_45924);
nand UO_917 (O_917,N_45203,N_46517);
xor UO_918 (O_918,N_47143,N_46535);
and UO_919 (O_919,N_48351,N_49840);
nor UO_920 (O_920,N_48526,N_45389);
and UO_921 (O_921,N_49353,N_47980);
nor UO_922 (O_922,N_49299,N_46080);
xnor UO_923 (O_923,N_45680,N_47200);
or UO_924 (O_924,N_47637,N_45061);
or UO_925 (O_925,N_45896,N_46694);
or UO_926 (O_926,N_47562,N_49489);
nand UO_927 (O_927,N_45527,N_45098);
nand UO_928 (O_928,N_47026,N_49722);
or UO_929 (O_929,N_47344,N_49108);
xnor UO_930 (O_930,N_47907,N_46446);
or UO_931 (O_931,N_47760,N_46793);
or UO_932 (O_932,N_48518,N_47186);
and UO_933 (O_933,N_45982,N_47644);
nand UO_934 (O_934,N_48175,N_45934);
or UO_935 (O_935,N_45554,N_49712);
nor UO_936 (O_936,N_49122,N_46298);
nor UO_937 (O_937,N_48105,N_46368);
nand UO_938 (O_938,N_49537,N_45991);
and UO_939 (O_939,N_47162,N_45121);
or UO_940 (O_940,N_45071,N_45783);
nand UO_941 (O_941,N_48298,N_49182);
nor UO_942 (O_942,N_46613,N_45279);
nor UO_943 (O_943,N_46417,N_45134);
nand UO_944 (O_944,N_49702,N_49920);
nand UO_945 (O_945,N_47450,N_48418);
xor UO_946 (O_946,N_46162,N_49652);
nor UO_947 (O_947,N_46429,N_45812);
or UO_948 (O_948,N_48422,N_48731);
and UO_949 (O_949,N_49228,N_45615);
or UO_950 (O_950,N_46421,N_45561);
and UO_951 (O_951,N_46617,N_46763);
nand UO_952 (O_952,N_49597,N_47349);
or UO_953 (O_953,N_48285,N_47319);
or UO_954 (O_954,N_46477,N_47898);
or UO_955 (O_955,N_47222,N_49968);
nor UO_956 (O_956,N_48487,N_45049);
nand UO_957 (O_957,N_45739,N_46139);
nand UO_958 (O_958,N_45020,N_46456);
nor UO_959 (O_959,N_45137,N_48508);
and UO_960 (O_960,N_47055,N_46812);
and UO_961 (O_961,N_45402,N_49949);
and UO_962 (O_962,N_45452,N_46784);
and UO_963 (O_963,N_47532,N_45175);
and UO_964 (O_964,N_47555,N_48816);
or UO_965 (O_965,N_46650,N_49793);
or UO_966 (O_966,N_46897,N_49874);
nand UO_967 (O_967,N_46509,N_48239);
nor UO_968 (O_968,N_47514,N_45933);
nor UO_969 (O_969,N_45253,N_46097);
nor UO_970 (O_970,N_45135,N_49932);
and UO_971 (O_971,N_45816,N_48066);
xnor UO_972 (O_972,N_47031,N_48057);
xor UO_973 (O_973,N_46369,N_48636);
nor UO_974 (O_974,N_47876,N_46605);
nor UO_975 (O_975,N_49672,N_46182);
or UO_976 (O_976,N_48925,N_46275);
nand UO_977 (O_977,N_48111,N_49999);
and UO_978 (O_978,N_48966,N_49435);
nor UO_979 (O_979,N_46608,N_48651);
or UO_980 (O_980,N_48625,N_49898);
and UO_981 (O_981,N_45328,N_46468);
xor UO_982 (O_982,N_48544,N_45779);
nor UO_983 (O_983,N_48183,N_48364);
and UO_984 (O_984,N_46094,N_47224);
and UO_985 (O_985,N_49534,N_45790);
nor UO_986 (O_986,N_46367,N_46753);
or UO_987 (O_987,N_45929,N_49072);
nor UO_988 (O_988,N_49867,N_48321);
or UO_989 (O_989,N_47057,N_48746);
nor UO_990 (O_990,N_45754,N_46445);
nand UO_991 (O_991,N_47776,N_45940);
xor UO_992 (O_992,N_47738,N_47545);
or UO_993 (O_993,N_49386,N_46754);
nand UO_994 (O_994,N_49125,N_49456);
or UO_995 (O_995,N_45740,N_49899);
or UO_996 (O_996,N_47019,N_47953);
xnor UO_997 (O_997,N_48141,N_46449);
nor UO_998 (O_998,N_47099,N_46076);
or UO_999 (O_999,N_48947,N_49804);
nor UO_1000 (O_1000,N_47083,N_48503);
nand UO_1001 (O_1001,N_45506,N_47136);
nand UO_1002 (O_1002,N_45364,N_48204);
nor UO_1003 (O_1003,N_49944,N_46668);
or UO_1004 (O_1004,N_45801,N_48840);
xor UO_1005 (O_1005,N_48798,N_49581);
and UO_1006 (O_1006,N_46513,N_49024);
and UO_1007 (O_1007,N_47300,N_49010);
nand UO_1008 (O_1008,N_46397,N_46108);
nand UO_1009 (O_1009,N_48317,N_45044);
nor UO_1010 (O_1010,N_48767,N_45162);
nand UO_1011 (O_1011,N_46825,N_48821);
or UO_1012 (O_1012,N_48075,N_46797);
xnor UO_1013 (O_1013,N_48166,N_49517);
or UO_1014 (O_1014,N_48860,N_49819);
nor UO_1015 (O_1015,N_47884,N_46448);
nand UO_1016 (O_1016,N_46124,N_49064);
or UO_1017 (O_1017,N_45418,N_46161);
and UO_1018 (O_1018,N_47253,N_49144);
nand UO_1019 (O_1019,N_48161,N_46842);
nand UO_1020 (O_1020,N_49321,N_48155);
nor UO_1021 (O_1021,N_45324,N_46250);
or UO_1022 (O_1022,N_45577,N_47579);
and UO_1023 (O_1023,N_48427,N_46951);
nand UO_1024 (O_1024,N_49082,N_46112);
nor UO_1025 (O_1025,N_45657,N_46500);
nand UO_1026 (O_1026,N_45384,N_47437);
nand UO_1027 (O_1027,N_45891,N_47935);
nand UO_1028 (O_1028,N_49065,N_49430);
and UO_1029 (O_1029,N_48023,N_45207);
xor UO_1030 (O_1030,N_46088,N_49314);
nand UO_1031 (O_1031,N_49665,N_48224);
and UO_1032 (O_1032,N_48823,N_49417);
or UO_1033 (O_1033,N_49462,N_47638);
and UO_1034 (O_1034,N_45503,N_48438);
nand UO_1035 (O_1035,N_49306,N_49961);
or UO_1036 (O_1036,N_46304,N_45099);
nor UO_1037 (O_1037,N_45675,N_45711);
nand UO_1038 (O_1038,N_45355,N_48512);
or UO_1039 (O_1039,N_46701,N_45111);
nand UO_1040 (O_1040,N_48345,N_49531);
nand UO_1041 (O_1041,N_49170,N_45333);
nand UO_1042 (O_1042,N_49231,N_49595);
nor UO_1043 (O_1043,N_45628,N_46342);
or UO_1044 (O_1044,N_45446,N_45642);
and UO_1045 (O_1045,N_46849,N_49440);
or UO_1046 (O_1046,N_45317,N_45032);
and UO_1047 (O_1047,N_45999,N_48015);
or UO_1048 (O_1048,N_49673,N_47393);
nand UO_1049 (O_1049,N_48065,N_47104);
nand UO_1050 (O_1050,N_47944,N_46852);
and UO_1051 (O_1051,N_46137,N_48973);
xor UO_1052 (O_1052,N_48125,N_46875);
nand UO_1053 (O_1053,N_45795,N_46371);
xnor UO_1054 (O_1054,N_47166,N_46636);
or UO_1055 (O_1055,N_49086,N_45821);
xor UO_1056 (O_1056,N_45763,N_49307);
or UO_1057 (O_1057,N_46029,N_47979);
or UO_1058 (O_1058,N_49787,N_49166);
nand UO_1059 (O_1059,N_49281,N_45937);
nor UO_1060 (O_1060,N_47156,N_46570);
or UO_1061 (O_1061,N_49713,N_47351);
or UO_1062 (O_1062,N_48606,N_45928);
and UO_1063 (O_1063,N_45208,N_46377);
and UO_1064 (O_1064,N_46839,N_49657);
nor UO_1065 (O_1065,N_45787,N_45743);
and UO_1066 (O_1066,N_49148,N_49146);
nor UO_1067 (O_1067,N_46223,N_45574);
nand UO_1068 (O_1068,N_46344,N_49782);
xnor UO_1069 (O_1069,N_48435,N_49979);
nor UO_1070 (O_1070,N_48567,N_49735);
and UO_1071 (O_1071,N_47716,N_48803);
or UO_1072 (O_1072,N_45077,N_46180);
and UO_1073 (O_1073,N_45055,N_47574);
nand UO_1074 (O_1074,N_47295,N_48004);
xor UO_1075 (O_1075,N_46270,N_45399);
nand UO_1076 (O_1076,N_45735,N_46249);
and UO_1077 (O_1077,N_49018,N_48090);
and UO_1078 (O_1078,N_45054,N_46310);
xnor UO_1079 (O_1079,N_47233,N_45027);
nor UO_1080 (O_1080,N_47711,N_46584);
nand UO_1081 (O_1081,N_46731,N_45853);
nand UO_1082 (O_1082,N_45637,N_45056);
or UO_1083 (O_1083,N_49427,N_46361);
nand UO_1084 (O_1084,N_49184,N_45029);
or UO_1085 (O_1085,N_45699,N_45494);
and UO_1086 (O_1086,N_45990,N_48726);
nand UO_1087 (O_1087,N_48012,N_48388);
nand UO_1088 (O_1088,N_49507,N_48912);
nand UO_1089 (O_1089,N_49753,N_49568);
and UO_1090 (O_1090,N_45074,N_46178);
nand UO_1091 (O_1091,N_46722,N_49304);
and UO_1092 (O_1092,N_49573,N_49522);
or UO_1093 (O_1093,N_45255,N_45646);
and UO_1094 (O_1094,N_47255,N_47219);
or UO_1095 (O_1095,N_47629,N_48156);
nor UO_1096 (O_1096,N_47817,N_49971);
nor UO_1097 (O_1097,N_47317,N_46326);
or UO_1098 (O_1098,N_49017,N_49381);
nand UO_1099 (O_1099,N_45875,N_47985);
and UO_1100 (O_1100,N_47318,N_49324);
xor UO_1101 (O_1101,N_46305,N_47988);
and UO_1102 (O_1102,N_47105,N_48936);
and UO_1103 (O_1103,N_49196,N_45729);
nor UO_1104 (O_1104,N_49167,N_45876);
nand UO_1105 (O_1105,N_49328,N_48771);
xnor UO_1106 (O_1106,N_49105,N_49193);
and UO_1107 (O_1107,N_48720,N_47208);
nand UO_1108 (O_1108,N_47125,N_49862);
or UO_1109 (O_1109,N_49413,N_49366);
xor UO_1110 (O_1110,N_45856,N_47540);
or UO_1111 (O_1111,N_45362,N_45733);
nor UO_1112 (O_1112,N_48882,N_47842);
or UO_1113 (O_1113,N_49739,N_49742);
or UO_1114 (O_1114,N_48797,N_47832);
nand UO_1115 (O_1115,N_47492,N_49552);
nor UO_1116 (O_1116,N_46997,N_47539);
and UO_1117 (O_1117,N_46020,N_48961);
nor UO_1118 (O_1118,N_46167,N_49038);
nand UO_1119 (O_1119,N_49302,N_47432);
nor UO_1120 (O_1120,N_45097,N_48179);
nand UO_1121 (O_1121,N_46320,N_47451);
xor UO_1122 (O_1122,N_46385,N_49609);
or UO_1123 (O_1123,N_45825,N_48520);
and UO_1124 (O_1124,N_48381,N_48638);
nor UO_1125 (O_1125,N_49567,N_46530);
and UO_1126 (O_1126,N_48369,N_48329);
nand UO_1127 (O_1127,N_49407,N_49564);
nand UO_1128 (O_1128,N_47175,N_46787);
nand UO_1129 (O_1129,N_48661,N_49197);
nor UO_1130 (O_1130,N_48420,N_48028);
or UO_1131 (O_1131,N_49433,N_45903);
or UO_1132 (O_1132,N_49487,N_45011);
nand UO_1133 (O_1133,N_49331,N_48398);
xnor UO_1134 (O_1134,N_46723,N_48683);
nand UO_1135 (O_1135,N_49078,N_45453);
nand UO_1136 (O_1136,N_49123,N_45897);
or UO_1137 (O_1137,N_45652,N_47434);
nand UO_1138 (O_1138,N_45083,N_45475);
nor UO_1139 (O_1139,N_46019,N_46129);
or UO_1140 (O_1140,N_47916,N_47847);
and UO_1141 (O_1141,N_49174,N_48403);
nand UO_1142 (O_1142,N_45166,N_45392);
or UO_1143 (O_1143,N_48088,N_47103);
and UO_1144 (O_1144,N_45370,N_49385);
or UO_1145 (O_1145,N_49490,N_45978);
nand UO_1146 (O_1146,N_47188,N_49201);
nand UO_1147 (O_1147,N_48173,N_49734);
and UO_1148 (O_1148,N_47048,N_47470);
or UO_1149 (O_1149,N_48811,N_45798);
or UO_1150 (O_1150,N_47052,N_46024);
nor UO_1151 (O_1151,N_49526,N_46175);
or UO_1152 (O_1152,N_49268,N_46003);
nor UO_1153 (O_1153,N_46612,N_49801);
nor UO_1154 (O_1154,N_47167,N_49110);
or UO_1155 (O_1155,N_49050,N_48093);
and UO_1156 (O_1156,N_45901,N_45966);
nand UO_1157 (O_1157,N_49442,N_47390);
and UO_1158 (O_1158,N_48292,N_48474);
nor UO_1159 (O_1159,N_48492,N_45834);
nand UO_1160 (O_1160,N_45064,N_45594);
and UO_1161 (O_1161,N_49135,N_49285);
or UO_1162 (O_1162,N_47176,N_49647);
or UO_1163 (O_1163,N_49929,N_46245);
nor UO_1164 (O_1164,N_47201,N_48149);
nor UO_1165 (O_1165,N_47819,N_49260);
nor UO_1166 (O_1166,N_47656,N_49877);
nand UO_1167 (O_1167,N_47771,N_49832);
or UO_1168 (O_1168,N_49032,N_46955);
and UO_1169 (O_1169,N_48778,N_48891);
or UO_1170 (O_1170,N_46950,N_48135);
and UO_1171 (O_1171,N_45018,N_47660);
and UO_1172 (O_1172,N_47408,N_46048);
nor UO_1173 (O_1173,N_46169,N_47930);
and UO_1174 (O_1174,N_48870,N_49951);
and UO_1175 (O_1175,N_47511,N_48326);
nor UO_1176 (O_1176,N_47089,N_47812);
nor UO_1177 (O_1177,N_49229,N_49208);
or UO_1178 (O_1178,N_45417,N_48994);
or UO_1179 (O_1179,N_48148,N_45996);
and UO_1180 (O_1180,N_45840,N_46765);
and UO_1181 (O_1181,N_48442,N_46373);
or UO_1182 (O_1182,N_46264,N_46588);
nand UO_1183 (O_1183,N_45107,N_45770);
or UO_1184 (O_1184,N_47012,N_46521);
or UO_1185 (O_1185,N_45085,N_47126);
nor UO_1186 (O_1186,N_47115,N_46840);
nor UO_1187 (O_1187,N_47594,N_48086);
and UO_1188 (O_1188,N_47456,N_49055);
nor UO_1189 (O_1189,N_49865,N_45599);
or UO_1190 (O_1190,N_49404,N_48039);
nand UO_1191 (O_1191,N_49687,N_47519);
nor UO_1192 (O_1192,N_47439,N_49011);
and UO_1193 (O_1193,N_49844,N_49863);
nor UO_1194 (O_1194,N_45593,N_49883);
and UO_1195 (O_1195,N_46038,N_45371);
and UO_1196 (O_1196,N_46166,N_48245);
nand UO_1197 (O_1197,N_46350,N_47261);
and UO_1198 (O_1198,N_48755,N_48801);
nor UO_1199 (O_1199,N_45602,N_45171);
and UO_1200 (O_1200,N_47189,N_48900);
and UO_1201 (O_1201,N_45584,N_48080);
nor UO_1202 (O_1202,N_47874,N_48443);
nor UO_1203 (O_1203,N_45218,N_45489);
nor UO_1204 (O_1204,N_46462,N_49948);
and UO_1205 (O_1205,N_46340,N_48449);
nand UO_1206 (O_1206,N_48067,N_45625);
or UO_1207 (O_1207,N_46943,N_47723);
nor UO_1208 (O_1208,N_47758,N_47358);
nand UO_1209 (O_1209,N_45712,N_48446);
nor UO_1210 (O_1210,N_48115,N_48549);
and UO_1211 (O_1211,N_49662,N_47538);
and UO_1212 (O_1212,N_45477,N_49370);
or UO_1213 (O_1213,N_45490,N_48603);
xnor UO_1214 (O_1214,N_49237,N_45239);
nor UO_1215 (O_1215,N_48880,N_47807);
xor UO_1216 (O_1216,N_47782,N_47433);
nand UO_1217 (O_1217,N_48219,N_45782);
nand UO_1218 (O_1218,N_45839,N_47037);
or UO_1219 (O_1219,N_47666,N_48909);
xor UO_1220 (O_1220,N_49074,N_47498);
or UO_1221 (O_1221,N_49347,N_49113);
or UO_1222 (O_1222,N_49233,N_48394);
nor UO_1223 (O_1223,N_48241,N_47963);
nor UO_1224 (O_1224,N_46981,N_45884);
nor UO_1225 (O_1225,N_49262,N_49792);
nor UO_1226 (O_1226,N_45078,N_47611);
nor UO_1227 (O_1227,N_48715,N_46114);
nor UO_1228 (O_1228,N_48377,N_49705);
nand UO_1229 (O_1229,N_47705,N_47381);
and UO_1230 (O_1230,N_49851,N_46409);
nor UO_1231 (O_1231,N_46534,N_46860);
nand UO_1232 (O_1232,N_47076,N_47264);
nand UO_1233 (O_1233,N_45915,N_47844);
and UO_1234 (O_1234,N_47544,N_49339);
and UO_1235 (O_1235,N_48291,N_47917);
nand UO_1236 (O_1236,N_45781,N_48048);
or UO_1237 (O_1237,N_48296,N_46759);
or UO_1238 (O_1238,N_48682,N_48874);
or UO_1239 (O_1239,N_47612,N_47712);
and UO_1240 (O_1240,N_49335,N_46314);
or UO_1241 (O_1241,N_45224,N_49066);
nand UO_1242 (O_1242,N_45741,N_48267);
nor UO_1243 (O_1243,N_45717,N_45360);
and UO_1244 (O_1244,N_46457,N_49721);
nand UO_1245 (O_1245,N_49894,N_49214);
nand UO_1246 (O_1246,N_49811,N_45811);
nor UO_1247 (O_1247,N_48783,N_49654);
and UO_1248 (O_1248,N_49525,N_49145);
nand UO_1249 (O_1249,N_46391,N_46730);
nor UO_1250 (O_1250,N_49934,N_48669);
nand UO_1251 (O_1251,N_47435,N_46789);
xor UO_1252 (O_1252,N_48693,N_49157);
xnor UO_1253 (O_1253,N_46454,N_47250);
or UO_1254 (O_1254,N_45557,N_47515);
nor UO_1255 (O_1255,N_45164,N_46012);
or UO_1256 (O_1256,N_46126,N_47281);
or UO_1257 (O_1257,N_45102,N_48923);
and UO_1258 (O_1258,N_46604,N_45456);
nand UO_1259 (O_1259,N_46532,N_48794);
xnor UO_1260 (O_1260,N_45145,N_46432);
nand UO_1261 (O_1261,N_47696,N_46594);
nor UO_1262 (O_1262,N_49985,N_46847);
and UO_1263 (O_1263,N_47682,N_46631);
nor UO_1264 (O_1264,N_48915,N_49265);
and UO_1265 (O_1265,N_49109,N_47102);
xnor UO_1266 (O_1266,N_47177,N_49856);
nand UO_1267 (O_1267,N_46437,N_46769);
and UO_1268 (O_1268,N_46323,N_46974);
nor UO_1269 (O_1269,N_45466,N_46289);
nand UO_1270 (O_1270,N_48517,N_49514);
and UO_1271 (O_1271,N_49821,N_46912);
and UO_1272 (O_1272,N_47356,N_47772);
and UO_1273 (O_1273,N_48257,N_48578);
xor UO_1274 (O_1274,N_47097,N_46560);
nand UO_1275 (O_1275,N_45117,N_46949);
or UO_1276 (O_1276,N_45014,N_45422);
or UO_1277 (O_1277,N_48792,N_48770);
nand UO_1278 (O_1278,N_45286,N_47323);
nand UO_1279 (O_1279,N_48690,N_48703);
nor UO_1280 (O_1280,N_49779,N_45051);
nand UO_1281 (O_1281,N_46545,N_47305);
or UO_1282 (O_1282,N_45844,N_49053);
xor UO_1283 (O_1283,N_47333,N_45872);
xnor UO_1284 (O_1284,N_46052,N_48975);
or UO_1285 (O_1285,N_49960,N_48597);
or UO_1286 (O_1286,N_47755,N_47254);
and UO_1287 (O_1287,N_47111,N_48645);
nor UO_1288 (O_1288,N_47493,N_48727);
nand UO_1289 (O_1289,N_45161,N_47027);
and UO_1290 (O_1290,N_49579,N_48104);
or UO_1291 (O_1291,N_48327,N_49348);
or UO_1292 (O_1292,N_49967,N_45757);
nand UO_1293 (O_1293,N_49731,N_49906);
or UO_1294 (O_1294,N_45058,N_47743);
or UO_1295 (O_1295,N_48304,N_46833);
nand UO_1296 (O_1296,N_48790,N_45606);
nor UO_1297 (O_1297,N_46630,N_45838);
and UO_1298 (O_1298,N_45732,N_45945);
xnor UO_1299 (O_1299,N_45967,N_49318);
xnor UO_1300 (O_1300,N_45749,N_45104);
and UO_1301 (O_1301,N_45769,N_48003);
or UO_1302 (O_1302,N_46405,N_49596);
xnor UO_1303 (O_1303,N_46615,N_49402);
and UO_1304 (O_1304,N_45632,N_45746);
or UO_1305 (O_1305,N_49607,N_46263);
nand UO_1306 (O_1306,N_45128,N_49701);
nand UO_1307 (O_1307,N_47218,N_48468);
nor UO_1308 (O_1308,N_47480,N_46309);
and UO_1309 (O_1309,N_45528,N_48610);
nand UO_1310 (O_1310,N_47977,N_45608);
or UO_1311 (O_1311,N_48263,N_45150);
nor UO_1312 (O_1312,N_48406,N_49533);
nand UO_1313 (O_1313,N_45356,N_46412);
nand UO_1314 (O_1314,N_46202,N_48988);
xor UO_1315 (O_1315,N_48644,N_48376);
and UO_1316 (O_1316,N_49897,N_46813);
xor UO_1317 (O_1317,N_46737,N_48576);
or UO_1318 (O_1318,N_48346,N_48101);
nor UO_1319 (O_1319,N_47315,N_45846);
and UO_1320 (O_1320,N_49422,N_48607);
and UO_1321 (O_1321,N_48144,N_47850);
nand UO_1322 (O_1322,N_47270,N_47021);
nor UO_1323 (O_1323,N_48350,N_48092);
or UO_1324 (O_1324,N_48830,N_49289);
xnor UO_1325 (O_1325,N_45455,N_47820);
xor UO_1326 (O_1326,N_46587,N_49019);
nand UO_1327 (O_1327,N_45334,N_48674);
nor UO_1328 (O_1328,N_47074,N_47578);
or UO_1329 (O_1329,N_47423,N_47978);
and UO_1330 (O_1330,N_47184,N_45509);
nand UO_1331 (O_1331,N_45913,N_49693);
and UO_1332 (O_1332,N_45835,N_46060);
or UO_1333 (O_1333,N_49205,N_46354);
nand UO_1334 (O_1334,N_45618,N_48613);
or UO_1335 (O_1335,N_49760,N_49103);
nand UO_1336 (O_1336,N_45240,N_49757);
and UO_1337 (O_1337,N_48496,N_48708);
nor UO_1338 (O_1338,N_47499,N_46420);
and UO_1339 (O_1339,N_48217,N_49154);
nand UO_1340 (O_1340,N_46179,N_49420);
or UO_1341 (O_1341,N_48246,N_49629);
or UO_1342 (O_1342,N_48099,N_45113);
or UO_1343 (O_1343,N_46039,N_47144);
and UO_1344 (O_1344,N_45108,N_46647);
or UO_1345 (O_1345,N_47713,N_46585);
nor UO_1346 (O_1346,N_47284,N_48457);
nor UO_1347 (O_1347,N_46826,N_48231);
or UO_1348 (O_1348,N_47477,N_45028);
nor UO_1349 (O_1349,N_49244,N_48951);
and UO_1350 (O_1350,N_47263,N_49003);
or UO_1351 (O_1351,N_46510,N_45961);
and UO_1352 (O_1352,N_46554,N_45214);
and UO_1353 (O_1353,N_45144,N_48383);
and UO_1354 (O_1354,N_48059,N_46045);
xor UO_1355 (O_1355,N_48278,N_47786);
or UO_1356 (O_1356,N_48938,N_47808);
or UO_1357 (O_1357,N_48190,N_47589);
xor UO_1358 (O_1358,N_49977,N_49696);
and UO_1359 (O_1359,N_48751,N_46498);
and UO_1360 (O_1360,N_47827,N_48272);
nand UO_1361 (O_1361,N_45562,N_48557);
nand UO_1362 (O_1362,N_45784,N_47342);
nor UO_1363 (O_1363,N_47352,N_47822);
or UO_1364 (O_1364,N_49666,N_45909);
nand UO_1365 (O_1365,N_47191,N_49437);
xor UO_1366 (O_1366,N_49211,N_46440);
or UO_1367 (O_1367,N_48629,N_45747);
nor UO_1368 (O_1368,N_45666,N_48548);
nand UO_1369 (O_1369,N_45393,N_46352);
or UO_1370 (O_1370,N_48196,N_48898);
nor UO_1371 (O_1371,N_45395,N_46194);
xor UO_1372 (O_1372,N_47406,N_49663);
nand UO_1373 (O_1373,N_49918,N_49777);
nand UO_1374 (O_1374,N_47479,N_49101);
xor UO_1375 (O_1375,N_47987,N_47952);
and UO_1376 (O_1376,N_45644,N_45958);
and UO_1377 (O_1377,N_49601,N_46290);
nor UO_1378 (O_1378,N_45670,N_47486);
nand UO_1379 (O_1379,N_45040,N_49890);
nor UO_1380 (O_1380,N_46511,N_47846);
and UO_1381 (O_1381,N_48050,N_45190);
nand UO_1382 (O_1382,N_48380,N_45773);
and UO_1383 (O_1383,N_48698,N_46188);
or UO_1384 (O_1384,N_48108,N_49224);
xor UO_1385 (O_1385,N_49246,N_49034);
and UO_1386 (O_1386,N_45250,N_49136);
nand UO_1387 (O_1387,N_45148,N_45234);
nand UO_1388 (O_1388,N_47017,N_45716);
nand UO_1389 (O_1389,N_49194,N_46490);
and UO_1390 (O_1390,N_45269,N_46662);
xor UO_1391 (O_1391,N_46867,N_47790);
xnor UO_1392 (O_1392,N_46771,N_46732);
and UO_1393 (O_1393,N_47062,N_49720);
nand UO_1394 (O_1394,N_47137,N_46287);
nand UO_1395 (O_1395,N_45555,N_46991);
nor UO_1396 (O_1396,N_47620,N_48139);
nand UO_1397 (O_1397,N_46232,N_48774);
or UO_1398 (O_1398,N_45251,N_45375);
xnor UO_1399 (O_1399,N_45907,N_48475);
nor UO_1400 (O_1400,N_49467,N_47466);
and UO_1401 (O_1401,N_48691,N_49091);
and UO_1402 (O_1402,N_49400,N_46927);
and UO_1403 (O_1403,N_49588,N_45654);
xor UO_1404 (O_1404,N_48529,N_49978);
nor UO_1405 (O_1405,N_45157,N_49822);
nand UO_1406 (O_1406,N_48542,N_49723);
nor UO_1407 (O_1407,N_49614,N_48565);
or UO_1408 (O_1408,N_45694,N_45570);
and UO_1409 (O_1409,N_49312,N_47006);
nand UO_1410 (O_1410,N_49747,N_45258);
and UO_1411 (O_1411,N_46209,N_48444);
or UO_1412 (O_1412,N_45951,N_48158);
and UO_1413 (O_1413,N_47296,N_46711);
nand UO_1414 (O_1414,N_49375,N_45818);
nand UO_1415 (O_1415,N_45000,N_45544);
and UO_1416 (O_1416,N_48244,N_45842);
or UO_1417 (O_1417,N_46782,N_46681);
and UO_1418 (O_1418,N_48314,N_49642);
nand UO_1419 (O_1419,N_47806,N_46030);
or UO_1420 (O_1420,N_49708,N_47529);
xor UO_1421 (O_1421,N_49618,N_46611);
and UO_1422 (O_1422,N_49059,N_46240);
and UO_1423 (O_1423,N_49258,N_48931);
nor UO_1424 (O_1424,N_47279,N_49428);
and UO_1425 (O_1425,N_47613,N_46607);
or UO_1426 (O_1426,N_47976,N_47478);
and UO_1427 (O_1427,N_49494,N_48972);
nor UO_1428 (O_1428,N_46533,N_48722);
nand UO_1429 (O_1429,N_45343,N_46803);
nor UO_1430 (O_1430,N_47626,N_46092);
xnor UO_1431 (O_1431,N_45673,N_45831);
nand UO_1432 (O_1432,N_45326,N_45737);
or UO_1433 (O_1433,N_49541,N_45911);
or UO_1434 (O_1434,N_47249,N_48944);
nand UO_1435 (O_1435,N_47079,N_45276);
or UO_1436 (O_1436,N_48555,N_46973);
and UO_1437 (O_1437,N_47609,N_49726);
nand UO_1438 (O_1438,N_48670,N_49461);
xor UO_1439 (O_1439,N_48447,N_49061);
nor UO_1440 (O_1440,N_46508,N_45799);
or UO_1441 (O_1441,N_45568,N_48114);
or UO_1442 (O_1442,N_46691,N_49070);
nand UO_1443 (O_1443,N_46590,N_45535);
nor UO_1444 (O_1444,N_45715,N_47113);
nand UO_1445 (O_1445,N_49966,N_46653);
or UO_1446 (O_1446,N_46942,N_46622);
nor UO_1447 (O_1447,N_45281,N_49730);
and UO_1448 (O_1448,N_45288,N_49390);
nand UO_1449 (O_1449,N_46572,N_45868);
and UO_1450 (O_1450,N_49505,N_49583);
and UO_1451 (O_1451,N_49378,N_47068);
and UO_1452 (O_1452,N_47260,N_48220);
or UO_1453 (O_1453,N_49085,N_46971);
nor UO_1454 (O_1454,N_46953,N_46903);
and UO_1455 (O_1455,N_48270,N_47803);
xor UO_1456 (O_1456,N_46744,N_47364);
and UO_1457 (O_1457,N_47659,N_47085);
nor UO_1458 (O_1458,N_48922,N_46688);
nand UO_1459 (O_1459,N_48650,N_48692);
nor UO_1460 (O_1460,N_45688,N_45285);
and UO_1461 (O_1461,N_46547,N_46645);
nand UO_1462 (O_1462,N_48856,N_45806);
and UO_1463 (O_1463,N_48053,N_45035);
nor UO_1464 (O_1464,N_46552,N_45138);
nand UO_1465 (O_1465,N_48728,N_45814);
xor UO_1466 (O_1466,N_45467,N_47843);
nor UO_1467 (O_1467,N_49603,N_45199);
xnor UO_1468 (O_1468,N_49463,N_48704);
xor UO_1469 (O_1469,N_48040,N_47677);
nand UO_1470 (O_1470,N_49927,N_46205);
and UO_1471 (O_1471,N_48208,N_49556);
nand UO_1472 (O_1472,N_47770,N_49185);
nor UO_1473 (O_1473,N_47605,N_48024);
and UO_1474 (O_1474,N_49992,N_45400);
nor UO_1475 (O_1475,N_49764,N_46404);
nor UO_1476 (O_1476,N_46220,N_49945);
nor UO_1477 (O_1477,N_45302,N_48106);
nor UO_1478 (O_1478,N_45867,N_48602);
nand UO_1479 (O_1479,N_46983,N_47283);
or UO_1480 (O_1480,N_45696,N_46766);
nor UO_1481 (O_1481,N_49042,N_46219);
and UO_1482 (O_1482,N_46858,N_47075);
nand UO_1483 (O_1483,N_46475,N_47302);
or UO_1484 (O_1484,N_45105,N_46489);
or UO_1485 (O_1485,N_46598,N_49223);
nand UO_1486 (O_1486,N_47379,N_46043);
nor UO_1487 (O_1487,N_47607,N_46386);
xnor UO_1488 (O_1488,N_46760,N_46506);
xor UO_1489 (O_1489,N_46444,N_46286);
nand UO_1490 (O_1490,N_48839,N_45541);
and UO_1491 (O_1491,N_47554,N_47757);
nor UO_1492 (O_1492,N_45043,N_47446);
and UO_1493 (O_1493,N_46907,N_45581);
xor UO_1494 (O_1494,N_45205,N_46727);
nand UO_1495 (O_1495,N_46655,N_46165);
and UO_1496 (O_1496,N_46565,N_48176);
and UO_1497 (O_1497,N_48360,N_45484);
or UO_1498 (O_1498,N_49121,N_47962);
nand UO_1499 (O_1499,N_45981,N_49519);
or UO_1500 (O_1500,N_48504,N_47788);
nor UO_1501 (O_1501,N_45481,N_49790);
nand UO_1502 (O_1502,N_47949,N_45101);
nand UO_1503 (O_1503,N_46332,N_47968);
xor UO_1504 (O_1504,N_49563,N_47109);
and UO_1505 (O_1505,N_47127,N_46225);
nand UO_1506 (O_1506,N_45331,N_45219);
and UO_1507 (O_1507,N_48016,N_47385);
nor UO_1508 (O_1508,N_47662,N_46268);
or UO_1509 (O_1509,N_45127,N_45613);
nor UO_1510 (O_1510,N_49278,N_45526);
xnor UO_1511 (O_1511,N_46061,N_48247);
and UO_1512 (O_1512,N_46986,N_45289);
or UO_1513 (O_1513,N_45432,N_48036);
or UO_1514 (O_1514,N_47947,N_47585);
nand UO_1515 (O_1515,N_47674,N_49524);
or UO_1516 (O_1516,N_45004,N_46963);
xnor UO_1517 (O_1517,N_48153,N_48284);
or UO_1518 (O_1518,N_49416,N_45833);
nor UO_1519 (O_1519,N_49671,N_48976);
and UO_1520 (O_1520,N_49919,N_46363);
nor UO_1521 (O_1521,N_47709,N_47634);
xnor UO_1522 (O_1522,N_45271,N_47628);
nor UO_1523 (O_1523,N_46976,N_48827);
nand UO_1524 (O_1524,N_46642,N_46068);
or UO_1525 (O_1525,N_47724,N_46726);
nand UO_1526 (O_1526,N_47899,N_46637);
and UO_1527 (O_1527,N_46854,N_49719);
nor UO_1528 (O_1528,N_49040,N_49271);
or UO_1529 (O_1529,N_47900,N_47796);
xor UO_1530 (O_1530,N_45318,N_48227);
or UO_1531 (O_1531,N_45188,N_48112);
and UO_1532 (O_1532,N_49683,N_49338);
nor UO_1533 (O_1533,N_49751,N_46783);
nor UO_1534 (O_1534,N_45725,N_46920);
and UO_1535 (O_1535,N_47427,N_47299);
or UO_1536 (O_1536,N_46778,N_47689);
or UO_1537 (O_1537,N_49255,N_48885);
nand UO_1538 (O_1538,N_48884,N_49186);
or UO_1539 (O_1539,N_47983,N_49947);
or UO_1540 (O_1540,N_46408,N_48791);
nor UO_1541 (O_1541,N_46197,N_48989);
nand UO_1542 (O_1542,N_48366,N_49981);
and UO_1543 (O_1543,N_46925,N_48122);
and UO_1544 (O_1544,N_47520,N_48665);
and UO_1545 (O_1545,N_49320,N_47236);
and UO_1546 (O_1546,N_49613,N_47754);
and UO_1547 (O_1547,N_45277,N_46913);
nand UO_1548 (O_1548,N_49337,N_45873);
nor UO_1549 (O_1549,N_48347,N_46836);
and UO_1550 (O_1550,N_45649,N_48387);
or UO_1551 (O_1551,N_48534,N_49332);
and UO_1552 (O_1552,N_49799,N_46077);
nor UO_1553 (O_1553,N_49039,N_47853);
and UO_1554 (O_1554,N_49094,N_46543);
xor UO_1555 (O_1555,N_46633,N_49089);
or UO_1556 (O_1556,N_46214,N_48987);
or UO_1557 (O_1557,N_46705,N_46185);
nand UO_1558 (O_1558,N_47923,N_47443);
and UO_1559 (O_1559,N_47095,N_45813);
nand UO_1560 (O_1560,N_45567,N_47407);
and UO_1561 (O_1561,N_47132,N_45702);
and UO_1562 (O_1562,N_48991,N_49733);
nand UO_1563 (O_1563,N_47024,N_45031);
nand UO_1564 (O_1564,N_45249,N_49905);
nand UO_1565 (O_1565,N_49555,N_49582);
and UO_1566 (O_1566,N_49367,N_46549);
nand UO_1567 (O_1567,N_47140,N_49288);
nor UO_1568 (O_1568,N_49421,N_46679);
xor UO_1569 (O_1569,N_46801,N_47298);
and UO_1570 (O_1570,N_48471,N_48405);
and UO_1571 (O_1571,N_48545,N_47211);
and UO_1572 (O_1572,N_49773,N_49885);
or UO_1573 (O_1573,N_46556,N_45603);
and UO_1574 (O_1574,N_46084,N_46105);
or UO_1575 (O_1575,N_49439,N_49033);
or UO_1576 (O_1576,N_46573,N_46460);
or UO_1577 (O_1577,N_49305,N_49771);
nor UO_1578 (O_1578,N_46356,N_45700);
or UO_1579 (O_1579,N_46247,N_47837);
nor UO_1580 (O_1580,N_45558,N_48277);
nor UO_1581 (O_1581,N_49715,N_49486);
nor UO_1582 (O_1582,N_48753,N_45665);
nor UO_1583 (O_1583,N_46497,N_45724);
nor UO_1584 (O_1584,N_47926,N_46745);
and UO_1585 (O_1585,N_46274,N_46337);
nand UO_1586 (O_1586,N_47601,N_46952);
xnor UO_1587 (O_1587,N_48222,N_48339);
or UO_1588 (O_1588,N_49854,N_49127);
nor UO_1589 (O_1589,N_48786,N_47138);
or UO_1590 (O_1590,N_49670,N_48411);
xnor UO_1591 (O_1591,N_47798,N_45487);
or UO_1592 (O_1592,N_47320,N_49704);
nor UO_1593 (O_1593,N_48627,N_48781);
xor UO_1594 (O_1594,N_45686,N_48294);
nand UO_1595 (O_1595,N_46078,N_49986);
nor UO_1596 (O_1596,N_45439,N_48052);
or UO_1597 (O_1597,N_46031,N_48254);
and UO_1598 (O_1598,N_47286,N_46228);
nand UO_1599 (O_1599,N_47227,N_45648);
or UO_1600 (O_1600,N_45883,N_46516);
and UO_1601 (O_1601,N_47906,N_45003);
xnor UO_1602 (O_1602,N_48062,N_47350);
nor UO_1603 (O_1603,N_48077,N_48828);
or UO_1604 (O_1604,N_46524,N_48147);
nand UO_1605 (O_1605,N_46975,N_45701);
nor UO_1606 (O_1606,N_47880,N_48025);
and UO_1607 (O_1607,N_48667,N_46478);
nor UO_1608 (O_1608,N_49980,N_45026);
nand UO_1609 (O_1609,N_45904,N_48397);
and UO_1610 (O_1610,N_45363,N_48623);
xnor UO_1611 (O_1611,N_46008,N_49590);
xor UO_1612 (O_1612,N_45826,N_45766);
nand UO_1613 (O_1613,N_49501,N_48436);
or UO_1614 (O_1614,N_45136,N_45133);
or UO_1615 (O_1615,N_47960,N_48251);
xnor UO_1616 (O_1616,N_46147,N_49414);
and UO_1617 (O_1617,N_46109,N_48286);
or UO_1618 (O_1618,N_47799,N_45412);
and UO_1619 (O_1619,N_47708,N_45859);
and UO_1620 (O_1620,N_49264,N_47982);
nor UO_1621 (O_1621,N_46069,N_48566);
nand UO_1622 (O_1622,N_48699,N_48187);
or UO_1623 (O_1623,N_48928,N_47516);
nand UO_1624 (O_1624,N_49336,N_48478);
xnor UO_1625 (O_1625,N_45041,N_48302);
nor UO_1626 (O_1626,N_45036,N_46693);
and UO_1627 (O_1627,N_46111,N_47197);
or UO_1628 (O_1628,N_46382,N_45376);
and UO_1629 (O_1629,N_45660,N_46901);
or UO_1630 (O_1630,N_45340,N_45764);
nand UO_1631 (O_1631,N_46658,N_48809);
or UO_1632 (O_1632,N_45865,N_49394);
or UO_1633 (O_1633,N_46004,N_48647);
nor UO_1634 (O_1634,N_45836,N_47756);
or UO_1635 (O_1635,N_49409,N_48349);
or UO_1636 (O_1636,N_47603,N_45448);
nand UO_1637 (O_1637,N_47867,N_47639);
nand UO_1638 (O_1638,N_49970,N_45583);
nand UO_1639 (O_1639,N_46471,N_48358);
or UO_1640 (O_1640,N_46499,N_49638);
nor UO_1641 (O_1641,N_46155,N_46244);
nor UO_1642 (O_1642,N_49027,N_49290);
nor UO_1643 (O_1643,N_48152,N_46504);
nand UO_1644 (O_1644,N_48600,N_46624);
nor UO_1645 (O_1645,N_49380,N_47149);
or UO_1646 (O_1646,N_46777,N_46115);
nand UO_1647 (O_1647,N_49423,N_47248);
nor UO_1648 (O_1648,N_47028,N_48932);
or UO_1649 (O_1649,N_45050,N_47523);
nor UO_1650 (O_1650,N_46334,N_45677);
nor UO_1651 (O_1651,N_49620,N_48109);
and UO_1652 (O_1652,N_49806,N_46383);
nand UO_1653 (O_1653,N_49326,N_45663);
nor UO_1654 (O_1654,N_48662,N_49474);
nand UO_1655 (O_1655,N_48579,N_46265);
and UO_1656 (O_1656,N_49301,N_46862);
nand UO_1657 (O_1657,N_49116,N_49393);
nand UO_1658 (O_1658,N_46235,N_49475);
nor UO_1659 (O_1659,N_46193,N_49914);
nand UO_1660 (O_1660,N_49766,N_47774);
and UO_1661 (O_1661,N_49425,N_46451);
and UO_1662 (O_1662,N_46814,N_47453);
and UO_1663 (O_1663,N_49383,N_46366);
or UO_1664 (O_1664,N_46850,N_46496);
nor UO_1665 (O_1665,N_46972,N_45046);
nand UO_1666 (O_1666,N_48712,N_49057);
and UO_1667 (O_1667,N_47735,N_45767);
nor UO_1668 (O_1668,N_45962,N_46476);
and UO_1669 (O_1669,N_47855,N_49694);
nand UO_1670 (O_1670,N_47999,N_47816);
nor UO_1671 (O_1671,N_45236,N_49643);
and UO_1672 (O_1672,N_48399,N_45820);
and UO_1673 (O_1673,N_45309,N_48137);
and UO_1674 (O_1674,N_48426,N_48910);
and UO_1675 (O_1675,N_46058,N_46798);
nor UO_1676 (O_1676,N_48765,N_49765);
and UO_1677 (O_1677,N_49454,N_45191);
xor UO_1678 (O_1678,N_47357,N_47405);
nor UO_1679 (O_1679,N_47897,N_49107);
nand UO_1680 (O_1680,N_45016,N_46116);
nor UO_1681 (O_1681,N_47277,N_46804);
or UO_1682 (O_1682,N_47425,N_48159);
nand UO_1683 (O_1683,N_49625,N_49470);
nor UO_1684 (O_1684,N_45081,N_49465);
or UO_1685 (O_1685,N_45248,N_49635);
nor UO_1686 (O_1686,N_46036,N_48986);
nand UO_1687 (O_1687,N_48934,N_48635);
nand UO_1688 (O_1688,N_46121,N_48723);
nor UO_1689 (O_1689,N_47623,N_45917);
xor UO_1690 (O_1690,N_48594,N_47185);
or UO_1691 (O_1691,N_49357,N_46578);
nand UO_1692 (O_1692,N_45143,N_47501);
nor UO_1693 (O_1693,N_46151,N_49481);
nor UO_1694 (O_1694,N_45622,N_46629);
nand UO_1695 (O_1695,N_46827,N_45954);
nand UO_1696 (O_1696,N_45182,N_48598);
nand UO_1697 (O_1697,N_45534,N_46222);
and UO_1698 (O_1698,N_45181,N_47203);
xnor UO_1699 (O_1699,N_49676,N_46872);
or UO_1700 (O_1700,N_46231,N_48924);
and UO_1701 (O_1701,N_47092,N_49833);
and UO_1702 (O_1702,N_45748,N_49317);
nand UO_1703 (O_1703,N_48020,N_46082);
nor UO_1704 (O_1704,N_49510,N_49111);
nor UO_1705 (O_1705,N_47484,N_47552);
and UO_1706 (O_1706,N_46216,N_47422);
nor UO_1707 (O_1707,N_45935,N_46331);
and UO_1708 (O_1708,N_45187,N_46227);
and UO_1709 (O_1709,N_45993,N_49007);
nand UO_1710 (O_1710,N_45900,N_47521);
or UO_1711 (O_1711,N_48589,N_49503);
or UO_1712 (O_1712,N_45604,N_45232);
nand UO_1713 (O_1713,N_47582,N_47077);
nor UO_1714 (O_1714,N_46273,N_45881);
nand UO_1715 (O_1715,N_48678,N_46300);
or UO_1716 (O_1716,N_49077,N_49095);
xor UO_1717 (O_1717,N_48207,N_48341);
nor UO_1718 (O_1718,N_48657,N_45695);
or UO_1719 (O_1719,N_47986,N_48575);
or UO_1720 (O_1720,N_49724,N_47067);
nor UO_1721 (O_1721,N_47505,N_49200);
nand UO_1722 (O_1722,N_46493,N_48085);
or UO_1723 (O_1723,N_46224,N_45086);
nor UO_1724 (O_1724,N_49313,N_48046);
nor UO_1725 (O_1725,N_47081,N_46059);
xnor UO_1726 (O_1726,N_46095,N_45629);
and UO_1727 (O_1727,N_45315,N_47376);
or UO_1728 (O_1728,N_46791,N_49817);
xnor UO_1729 (O_1729,N_47955,N_45815);
nor UO_1730 (O_1730,N_48960,N_49327);
nand UO_1731 (O_1731,N_49518,N_47122);
or UO_1732 (O_1732,N_47152,N_49013);
xnor UO_1733 (O_1733,N_46181,N_45247);
and UO_1734 (O_1734,N_48980,N_45768);
nor UO_1735 (O_1735,N_45946,N_45223);
or UO_1736 (O_1736,N_49164,N_46453);
or UO_1737 (O_1737,N_45390,N_45819);
xor UO_1738 (O_1738,N_46576,N_48688);
or UO_1739 (O_1739,N_49169,N_47412);
or UO_1740 (O_1740,N_45540,N_48560);
or UO_1741 (O_1741,N_45123,N_49902);
and UO_1742 (O_1742,N_45860,N_48401);
nand UO_1743 (O_1743,N_48524,N_45217);
and UO_1744 (O_1744,N_47050,N_46772);
and UO_1745 (O_1745,N_49140,N_45093);
and UO_1746 (O_1746,N_47896,N_45894);
nand UO_1747 (O_1747,N_49021,N_46939);
or UO_1748 (O_1748,N_45221,N_46242);
and UO_1749 (O_1749,N_47528,N_48523);
xor UO_1750 (O_1750,N_46558,N_45476);
and UO_1751 (O_1751,N_49572,N_48119);
or UO_1752 (O_1752,N_45242,N_48189);
or UO_1753 (O_1753,N_47797,N_48979);
or UO_1754 (O_1754,N_48134,N_46892);
nand UO_1755 (O_1755,N_46855,N_45159);
nor UO_1756 (O_1756,N_47684,N_49675);
nand UO_1757 (O_1757,N_49303,N_45119);
or UO_1758 (O_1758,N_47794,N_46700);
and UO_1759 (O_1759,N_45538,N_47804);
and UO_1760 (O_1760,N_48201,N_48883);
nand UO_1761 (O_1761,N_47714,N_49700);
and UO_1762 (O_1762,N_46733,N_47671);
xor UO_1763 (O_1763,N_45857,N_48897);
xor UO_1764 (O_1764,N_49310,N_46626);
nand UO_1765 (O_1765,N_47676,N_49756);
and UO_1766 (O_1766,N_49351,N_48554);
nand UO_1767 (O_1767,N_45671,N_46153);
nor UO_1768 (O_1768,N_46384,N_45226);
or UO_1769 (O_1769,N_45930,N_47292);
xor UO_1770 (O_1770,N_49943,N_47206);
and UO_1771 (O_1771,N_45088,N_49274);
or UO_1772 (O_1772,N_47558,N_48299);
and UO_1773 (O_1773,N_48469,N_45374);
nand UO_1774 (O_1774,N_49014,N_49030);
and UO_1775 (O_1775,N_47503,N_49172);
or UO_1776 (O_1776,N_46610,N_46308);
or UO_1777 (O_1777,N_45491,N_47310);
xor UO_1778 (O_1778,N_46846,N_45634);
or UO_1779 (O_1779,N_47569,N_47306);
xor UO_1780 (O_1780,N_48593,N_47362);
nor UO_1781 (O_1781,N_49479,N_48325);
and UO_1782 (O_1782,N_46199,N_45786);
nand UO_1783 (O_1783,N_49835,N_48083);
nor UO_1784 (O_1784,N_48762,N_46571);
or UO_1785 (O_1785,N_49106,N_49329);
nor UO_1786 (O_1786,N_47117,N_49399);
nand UO_1787 (O_1787,N_46394,N_47838);
xnor UO_1788 (O_1788,N_49808,N_46170);
xnor UO_1789 (O_1789,N_46035,N_49909);
nor UO_1790 (O_1790,N_47322,N_49079);
xor UO_1791 (O_1791,N_49045,N_47424);
xor UO_1792 (O_1792,N_45275,N_47993);
or UO_1793 (O_1793,N_47013,N_46752);
and UO_1794 (O_1794,N_46230,N_46027);
or UO_1795 (O_1795,N_46761,N_49617);
nand UO_1796 (O_1796,N_47954,N_47330);
and UO_1797 (O_1797,N_45210,N_47934);
nor UO_1798 (O_1798,N_48440,N_45008);
or UO_1799 (O_1799,N_46487,N_48370);
and UO_1800 (O_1800,N_49893,N_46113);
and UO_1801 (O_1801,N_47230,N_47951);
nand UO_1802 (O_1802,N_49983,N_49218);
nor UO_1803 (O_1803,N_45069,N_48136);
and UO_1804 (O_1804,N_48484,N_46168);
and UO_1805 (O_1805,N_49593,N_45592);
nor UO_1806 (O_1806,N_46674,N_47631);
xnor UO_1807 (O_1807,N_49585,N_45186);
xor UO_1808 (O_1808,N_48887,N_48970);
nor UO_1809 (O_1809,N_49685,N_46935);
nor UO_1810 (O_1810,N_47658,N_46980);
and UO_1811 (O_1811,N_46311,N_47965);
or UO_1812 (O_1812,N_49789,N_49709);
and UO_1813 (O_1813,N_46208,N_45292);
nand UO_1814 (O_1814,N_45468,N_49622);
or UO_1815 (O_1815,N_47877,N_47618);
nor UO_1816 (O_1816,N_47522,N_49044);
and UO_1817 (O_1817,N_49933,N_47431);
or UO_1818 (O_1818,N_46098,N_49565);
and UO_1819 (O_1819,N_46423,N_49910);
or UO_1820 (O_1820,N_45963,N_45366);
nor UO_1821 (O_1821,N_47290,N_47473);
and UO_1822 (O_1822,N_48103,N_47280);
nor UO_1823 (O_1823,N_47187,N_47742);
xnor UO_1824 (O_1824,N_45791,N_48528);
nor UO_1825 (O_1825,N_45297,N_47165);
or UO_1826 (O_1826,N_47636,N_48510);
nor UO_1827 (O_1827,N_48658,N_46399);
and UO_1828 (O_1828,N_45713,N_46402);
or UO_1829 (O_1829,N_47022,N_47700);
nor UO_1830 (O_1830,N_48194,N_49842);
or UO_1831 (O_1831,N_47086,N_45607);
nor UO_1832 (O_1832,N_46375,N_45369);
nand UO_1833 (O_1833,N_46581,N_49482);
and UO_1834 (O_1834,N_49813,N_46387);
xnor UO_1835 (O_1835,N_47009,N_48967);
or UO_1836 (O_1836,N_48556,N_46062);
nand UO_1837 (O_1837,N_49848,N_48519);
nand UO_1838 (O_1838,N_47046,N_49023);
xnor UO_1839 (O_1839,N_46824,N_47736);
nand UO_1840 (O_1840,N_45075,N_47216);
and UO_1841 (O_1841,N_47240,N_46893);
nor UO_1842 (O_1842,N_48848,N_46718);
nand UO_1843 (O_1843,N_48939,N_47066);
nor UO_1844 (O_1844,N_46330,N_46017);
nand UO_1845 (O_1845,N_47683,N_48580);
xor UO_1846 (O_1846,N_45736,N_48940);
nand UO_1847 (O_1847,N_48585,N_45566);
nand UO_1848 (O_1848,N_48639,N_46439);
or UO_1849 (O_1849,N_46979,N_49717);
nor UO_1850 (O_1850,N_48002,N_45227);
nand UO_1851 (O_1851,N_49810,N_45001);
or UO_1852 (O_1852,N_45721,N_47513);
xnor UO_1853 (O_1853,N_49434,N_45927);
nor UO_1854 (O_1854,N_48133,N_49736);
xnor UO_1855 (O_1855,N_47653,N_47096);
nor UO_1856 (O_1856,N_49352,N_49892);
nor UO_1857 (O_1857,N_48721,N_48307);
and UO_1858 (O_1858,N_48543,N_45480);
nand UO_1859 (O_1859,N_47885,N_49661);
or UO_1860 (O_1860,N_48076,N_46458);
and UO_1861 (O_1861,N_49159,N_47444);
and UO_1862 (O_1862,N_49355,N_47378);
and UO_1863 (O_1863,N_45065,N_46001);
nor UO_1864 (O_1864,N_49415,N_48965);
and UO_1865 (O_1865,N_45268,N_47669);
nand UO_1866 (O_1866,N_48889,N_48990);
nand UO_1867 (O_1867,N_48918,N_46916);
nand UO_1868 (O_1868,N_46682,N_49542);
nand UO_1869 (O_1869,N_47309,N_46322);
nor UO_1870 (O_1870,N_46157,N_45980);
nor UO_1871 (O_1871,N_48872,N_46550);
and UO_1872 (O_1872,N_49616,N_45939);
nor UO_1873 (O_1873,N_47542,N_46142);
nor UO_1874 (O_1874,N_48410,N_46580);
xnor UO_1875 (O_1875,N_47945,N_45922);
nor UO_1876 (O_1876,N_47282,N_49210);
and UO_1877 (O_1877,N_48569,N_46503);
and UO_1878 (O_1878,N_48621,N_46919);
xor UO_1879 (O_1879,N_46336,N_46474);
xnor UO_1880 (O_1880,N_46964,N_46365);
and UO_1881 (O_1881,N_47049,N_45185);
nor UO_1882 (O_1882,N_46110,N_45304);
and UO_1883 (O_1883,N_45312,N_46796);
or UO_1884 (O_1884,N_49606,N_49651);
or UO_1885 (O_1885,N_46676,N_45762);
nor UO_1886 (O_1886,N_45886,N_47893);
or UO_1887 (O_1887,N_48210,N_46643);
and UO_1888 (O_1888,N_48596,N_48685);
nor UO_1889 (O_1889,N_46866,N_46143);
xor UO_1890 (O_1890,N_49284,N_49401);
nand UO_1891 (O_1891,N_49063,N_48262);
nor UO_1892 (O_1892,N_45195,N_47151);
or UO_1893 (O_1893,N_46152,N_49273);
and UO_1894 (O_1894,N_48110,N_46898);
xnor UO_1895 (O_1895,N_45112,N_47231);
nand UO_1896 (O_1896,N_46087,N_45365);
xor UO_1897 (O_1897,N_46212,N_49052);
nor UO_1898 (O_1898,N_45237,N_48946);
and UO_1899 (O_1899,N_45387,N_49189);
nand UO_1900 (O_1900,N_46652,N_46800);
nor UO_1901 (O_1901,N_46215,N_48697);
nor UO_1902 (O_1902,N_47160,N_49584);
xor UO_1903 (O_1903,N_48017,N_47343);
nand UO_1904 (O_1904,N_46993,N_48949);
nor UO_1905 (O_1905,N_47942,N_47866);
nor UO_1906 (O_1906,N_47722,N_45829);
and UO_1907 (O_1907,N_47697,N_45726);
nor UO_1908 (O_1908,N_45154,N_47996);
nor UO_1909 (O_1909,N_45681,N_49632);
nand UO_1910 (O_1910,N_45956,N_49521);
nand UO_1911 (O_1911,N_48793,N_47547);
nor UO_1912 (O_1912,N_47940,N_45436);
nor UO_1913 (O_1913,N_49450,N_47335);
and UO_1914 (O_1914,N_47340,N_46623);
nand UO_1915 (O_1915,N_45895,N_46269);
xnor UO_1916 (O_1916,N_45211,N_45635);
and UO_1917 (O_1917,N_46376,N_47061);
or UO_1918 (O_1918,N_46100,N_45804);
nand UO_1919 (O_1919,N_49002,N_49272);
nor UO_1920 (O_1920,N_46902,N_48473);
xor UO_1921 (O_1921,N_45457,N_48452);
nand UO_1922 (O_1922,N_47872,N_46480);
nor UO_1923 (O_1923,N_45847,N_49680);
or UO_1924 (O_1924,N_45502,N_46635);
nor UO_1925 (O_1925,N_45151,N_45919);
nand UO_1926 (O_1926,N_48820,N_49207);
and UO_1927 (O_1927,N_48051,N_48072);
or UO_1928 (O_1928,N_48571,N_48390);
nor UO_1929 (O_1929,N_45595,N_45115);
or UO_1930 (O_1930,N_48391,N_47598);
nand UO_1931 (O_1931,N_49997,N_45564);
and UO_1932 (O_1932,N_46930,N_45611);
nand UO_1933 (O_1933,N_47029,N_47732);
or UO_1934 (O_1934,N_45006,N_48729);
nor UO_1935 (O_1935,N_49426,N_48539);
nand UO_1936 (O_1936,N_46295,N_48491);
nor UO_1937 (O_1937,N_45906,N_49658);
xnor UO_1938 (O_1938,N_48365,N_49261);
or UO_1939 (O_1939,N_45830,N_46692);
and UO_1940 (O_1940,N_47301,N_47488);
or UO_1941 (O_1941,N_45329,N_45398);
and UO_1942 (O_1942,N_48495,N_45950);
or UO_1943 (O_1943,N_46894,N_45426);
and UO_1944 (O_1944,N_47699,N_47449);
and UO_1945 (O_1945,N_46259,N_47386);
or UO_1946 (O_1946,N_49368,N_49660);
nand UO_1947 (O_1947,N_49718,N_47018);
or UO_1948 (O_1948,N_46328,N_46319);
nor UO_1949 (O_1949,N_45059,N_47210);
nor UO_1950 (O_1950,N_46591,N_45624);
nand UO_1951 (O_1951,N_46467,N_45578);
nand UO_1952 (O_1952,N_49084,N_47173);
nor UO_1953 (O_1953,N_48929,N_47497);
nand UO_1954 (O_1954,N_49493,N_47632);
and UO_1955 (O_1955,N_49340,N_45483);
and UO_1956 (O_1956,N_45960,N_46430);
and UO_1957 (O_1957,N_48768,N_45852);
nor UO_1958 (O_1958,N_48316,N_48408);
nand UO_1959 (O_1959,N_47901,N_46835);
or UO_1960 (O_1960,N_49048,N_49775);
nand UO_1961 (O_1961,N_48416,N_48916);
and UO_1962 (O_1962,N_46134,N_49343);
nor UO_1963 (O_1963,N_49130,N_46207);
xor UO_1964 (O_1964,N_48343,N_48280);
xor UO_1965 (O_1965,N_49062,N_45576);
or UO_1966 (O_1966,N_49175,N_48490);
nand UO_1967 (O_1967,N_48324,N_49466);
or UO_1968 (O_1968,N_48197,N_46177);
and UO_1969 (O_1969,N_47882,N_47440);
or UO_1970 (O_1970,N_47902,N_47961);
and UO_1971 (O_1971,N_47215,N_48619);
and UO_1972 (O_1972,N_47194,N_47073);
or UO_1973 (O_1973,N_45060,N_48060);
nand UO_1974 (O_1974,N_48320,N_48315);
and UO_1975 (O_1975,N_47217,N_45944);
and UO_1976 (O_1976,N_47768,N_49491);
nand UO_1977 (O_1977,N_47303,N_49341);
and UO_1978 (O_1978,N_49506,N_45425);
xor UO_1979 (O_1979,N_48340,N_45889);
nand UO_1980 (O_1980,N_45926,N_46123);
nor UO_1981 (O_1981,N_45177,N_45140);
or UO_1982 (O_1982,N_48763,N_47426);
nand UO_1983 (O_1983,N_48806,N_48673);
and UO_1984 (O_1984,N_46822,N_46544);
nor UO_1985 (O_1985,N_45633,N_49690);
xnor UO_1986 (O_1986,N_46528,N_45845);
nand UO_1987 (O_1987,N_47517,N_46388);
and UO_1988 (O_1988,N_46442,N_49080);
and UO_1989 (O_1989,N_46284,N_49300);
nand UO_1990 (O_1990,N_49295,N_47403);
nand UO_1991 (O_1991,N_46041,N_46817);
and UO_1992 (O_1992,N_45458,N_45751);
nand UO_1993 (O_1993,N_48212,N_49444);
or UO_1994 (O_1994,N_47886,N_47275);
nor UO_1995 (O_1995,N_48288,N_46788);
nand UO_1996 (O_1996,N_47720,N_45479);
or UO_1997 (O_1997,N_45971,N_45505);
nor UO_1998 (O_1998,N_49528,N_47476);
or UO_1999 (O_1999,N_47316,N_45559);
or UO_2000 (O_2000,N_45338,N_45925);
xnor UO_2001 (O_2001,N_47041,N_49772);
nand UO_2002 (O_2002,N_47234,N_48764);
and UO_2003 (O_2003,N_45572,N_46239);
nand UO_2004 (O_2004,N_45172,N_49650);
nor UO_2005 (O_2005,N_49767,N_48642);
and UO_2006 (O_2006,N_45409,N_45849);
nor UO_2007 (O_2007,N_45731,N_46089);
and UO_2008 (O_2008,N_47447,N_45910);
or UO_2009 (O_2009,N_47438,N_46970);
and UO_2010 (O_2010,N_48252,N_49176);
nand UO_2011 (O_2011,N_46687,N_47818);
nor UO_2012 (O_2012,N_45330,N_46443);
and UO_2013 (O_2013,N_46067,N_48759);
nand UO_2014 (O_2014,N_46410,N_46262);
xor UO_2015 (O_2015,N_49498,N_48055);
or UO_2016 (O_2016,N_46229,N_45658);
nor UO_2017 (O_2017,N_48505,N_46661);
nand UO_2018 (O_2018,N_49908,N_47325);
nand UO_2019 (O_2019,N_48849,N_48037);
or UO_2020 (O_2020,N_47765,N_46464);
or UO_2021 (O_2021,N_48927,N_49502);
nand UO_2022 (O_2022,N_47339,N_46947);
nor UO_2023 (O_2023,N_47830,N_47894);
xor UO_2024 (O_2024,N_45775,N_48772);
xor UO_2025 (O_2025,N_47868,N_47181);
nand UO_2026 (O_2026,N_47997,N_46518);
and UO_2027 (O_2027,N_45994,N_48750);
or UO_2028 (O_2028,N_46526,N_45155);
or UO_2029 (O_2029,N_45160,N_48041);
and UO_2030 (O_2030,N_48962,N_46000);
and UO_2031 (O_2031,N_45427,N_47879);
nand UO_2032 (O_2032,N_47767,N_49451);
nor UO_2033 (O_2033,N_47615,N_48978);
xnor UO_2034 (O_2034,N_47180,N_45244);
nor UO_2035 (O_2035,N_45952,N_45437);
and UO_2036 (O_2036,N_48181,N_49781);
nand UO_2037 (O_2037,N_47441,N_46857);
and UO_2038 (O_2038,N_46174,N_49249);
nor UO_2039 (O_2039,N_47064,N_47474);
xnor UO_2040 (O_2040,N_48248,N_47775);
nor UO_2041 (O_2041,N_49553,N_47888);
and UO_2042 (O_2042,N_48160,N_47922);
or UO_2043 (O_2043,N_45690,N_45864);
and UO_2044 (O_2044,N_47745,N_47835);
nand UO_2045 (O_2045,N_47404,N_45656);
nor UO_2046 (O_2046,N_48249,N_48038);
or UO_2047 (O_2047,N_48738,N_45493);
nand UO_2048 (O_2048,N_47959,N_47691);
or UO_2049 (O_2049,N_48808,N_47287);
or UO_2050 (O_2050,N_47783,N_49915);
nor UO_2051 (O_2051,N_48409,N_46946);
and UO_2052 (O_2052,N_45367,N_49406);
nand UO_2053 (O_2053,N_45582,N_47734);
nand UO_2054 (O_2054,N_45837,N_47100);
and UO_2055 (O_2055,N_49982,N_47810);
or UO_2056 (O_2056,N_45976,N_45463);
nor UO_2057 (O_2057,N_45495,N_47402);
nor UO_2058 (O_2058,N_48847,N_46670);
nand UO_2059 (O_2059,N_47419,N_45623);
xnor UO_2060 (O_2060,N_46130,N_46933);
and UO_2061 (O_2061,N_48997,N_45914);
nand UO_2062 (O_2062,N_47107,N_48354);
nand UO_2063 (O_2063,N_48701,N_45053);
nand UO_2064 (O_2064,N_47147,N_45235);
and UO_2065 (O_2065,N_48001,N_49604);
nand UO_2066 (O_2066,N_45545,N_49008);
or UO_2067 (O_2067,N_47463,N_49361);
or UO_2068 (O_2068,N_49744,N_46522);
xnor UO_2069 (O_2069,N_48047,N_47020);
nor UO_2070 (O_2070,N_48521,N_48687);
nor UO_2071 (O_2071,N_48319,N_46805);
or UO_2072 (O_2072,N_48154,N_45149);
or UO_2073 (O_2073,N_46173,N_49917);
or UO_2074 (O_2074,N_48087,N_49679);
or UO_2075 (O_2075,N_47307,N_48950);
xnor UO_2076 (O_2076,N_47164,N_49803);
nor UO_2077 (O_2077,N_45156,N_49411);
or UO_2078 (O_2078,N_45609,N_48295);
and UO_2079 (O_2079,N_48234,N_48355);
xnor UO_2080 (O_2080,N_46773,N_47472);
nand UO_2081 (O_2081,N_48935,N_49941);
nand UO_2082 (O_2082,N_49275,N_49128);
and UO_2083 (O_2083,N_48865,N_47672);
and UO_2084 (O_2084,N_49071,N_48747);
or UO_2085 (O_2085,N_49376,N_48511);
nor UO_2086 (O_2086,N_49362,N_49786);
and UO_2087 (O_2087,N_45197,N_46118);
and UO_2088 (O_2088,N_48531,N_47958);
or UO_2089 (O_2089,N_48836,N_48333);
and UO_2090 (O_2090,N_46501,N_49869);
or UO_2091 (O_2091,N_49913,N_45062);
and UO_2092 (O_2092,N_47002,N_47892);
nand UO_2093 (O_2093,N_46548,N_48640);
nor UO_2094 (O_2094,N_47271,N_47650);
and UO_2095 (O_2095,N_48393,N_46044);
xor UO_2096 (O_2096,N_48805,N_48573);
nand UO_2097 (O_2097,N_49453,N_49610);
or UO_2098 (O_2098,N_47141,N_49203);
nand UO_2099 (O_2099,N_47494,N_46447);
or UO_2100 (O_2100,N_45184,N_47304);
and UO_2101 (O_2101,N_46596,N_45347);
nand UO_2102 (O_2102,N_47267,N_45639);
nor UO_2103 (O_2103,N_47565,N_49372);
and UO_2104 (O_2104,N_45076,N_48458);
nand UO_2105 (O_2105,N_47005,N_46702);
and UO_2106 (O_2106,N_48879,N_46053);
or UO_2107 (O_2107,N_46808,N_48536);
nand UO_2108 (O_2108,N_46525,N_46600);
nor UO_2109 (O_2109,N_48930,N_48021);
and UO_2110 (O_2110,N_49689,N_47651);
and UO_2111 (O_2111,N_46183,N_48668);
nor UO_2112 (O_2112,N_46218,N_46934);
or UO_2113 (O_2113,N_45752,N_49099);
and UO_2114 (O_2114,N_46749,N_49473);
nor UO_2115 (O_2115,N_45923,N_46381);
nor UO_2116 (O_2116,N_46848,N_48943);
or UO_2117 (O_2117,N_47247,N_47183);
nand UO_2118 (O_2118,N_47332,N_45589);
nand UO_2119 (O_2119,N_45709,N_47145);
nor UO_2120 (O_2120,N_48306,N_46002);
nand UO_2121 (O_2121,N_48641,N_47223);
nor UO_2122 (O_2122,N_47616,N_47033);
and UO_2123 (O_2123,N_46968,N_47459);
or UO_2124 (O_2124,N_46714,N_47860);
nand UO_2125 (O_2125,N_47805,N_45068);
nand UO_2126 (O_2126,N_49081,N_46961);
and UO_2127 (O_2127,N_48971,N_45080);
nand UO_2128 (O_2128,N_46553,N_47635);
or UO_2129 (O_2129,N_45662,N_47496);
nand UO_2130 (O_2130,N_49243,N_47701);
and UO_2131 (O_2131,N_49991,N_47482);
xnor UO_2132 (O_2132,N_47763,N_49639);
nand UO_2133 (O_2133,N_49377,N_45949);
nand UO_2134 (O_2134,N_46422,N_49922);
and UO_2135 (O_2135,N_48500,N_48202);
or UO_2136 (O_2136,N_45753,N_47090);
and UO_2137 (O_2137,N_47108,N_49322);
or UO_2138 (O_2138,N_46889,N_49104);
nor UO_2139 (O_2139,N_47119,N_49395);
and UO_2140 (O_2140,N_47244,N_45441);
or UO_2141 (O_2141,N_49316,N_46856);
nor UO_2142 (O_2142,N_49828,N_45805);
or UO_2143 (O_2143,N_49911,N_47366);
nand UO_2144 (O_2144,N_47586,N_47655);
and UO_2145 (O_2145,N_48256,N_49993);
nand UO_2146 (O_2146,N_48881,N_49315);
and UO_2147 (O_2147,N_48527,N_47749);
nand UO_2148 (O_2148,N_47410,N_45039);
nor UO_2149 (O_2149,N_49431,N_47859);
and UO_2150 (O_2150,N_46419,N_47500);
and UO_2151 (O_2151,N_47341,N_47848);
nor UO_2152 (O_2152,N_49026,N_45517);
or UO_2153 (O_2153,N_46994,N_46472);
or UO_2154 (O_2154,N_49171,N_47583);
and UO_2155 (O_2155,N_45542,N_47004);
or UO_2156 (O_2156,N_48253,N_46958);
nor UO_2157 (O_2157,N_47557,N_49746);
and UO_2158 (O_2158,N_49812,N_46962);
nor UO_2159 (O_2159,N_46271,N_49520);
nand UO_2160 (O_2160,N_48842,N_46829);
nor UO_2161 (O_2161,N_47428,N_48876);
xor UO_2162 (O_2162,N_49884,N_49497);
or UO_2163 (O_2163,N_47998,N_48782);
nor UO_2164 (O_2164,N_46669,N_48318);
and UO_2165 (O_2165,N_45727,N_45017);
or UO_2166 (O_2166,N_45434,N_46238);
nor UO_2167 (O_2167,N_48574,N_49695);
xor UO_2168 (O_2168,N_47416,N_47429);
nand UO_2169 (O_2169,N_49688,N_47570);
or UO_2170 (O_2170,N_49478,N_47670);
nand UO_2171 (O_2171,N_46463,N_49396);
or UO_2172 (O_2172,N_48481,N_48300);
xnor UO_2173 (O_2173,N_46706,N_47274);
or UO_2174 (O_2174,N_49942,N_49323);
nor UO_2175 (O_2175,N_47928,N_47326);
xor UO_2176 (O_2176,N_49150,N_49460);
nand UO_2177 (O_2177,N_49215,N_46960);
nor UO_2178 (O_2178,N_45579,N_45878);
nand UO_2179 (O_2179,N_46395,N_49359);
nor UO_2180 (O_2180,N_46046,N_47171);
xnor UO_2181 (O_2181,N_49098,N_46495);
nor UO_2182 (O_2182,N_45084,N_49600);
and UO_2183 (O_2183,N_49824,N_48853);
nand UO_2184 (O_2184,N_45959,N_45116);
or UO_2185 (O_2185,N_48448,N_49006);
or UO_2186 (O_2186,N_49664,N_46333);
and UO_2187 (O_2187,N_48689,N_48902);
or UO_2188 (O_2188,N_47169,N_48126);
nor UO_2189 (O_2189,N_49291,N_49845);
xnor UO_2190 (O_2190,N_47288,N_48559);
nor UO_2191 (O_2191,N_46374,N_48675);
or UO_2192 (O_2192,N_47370,N_46592);
and UO_2193 (O_2193,N_49536,N_47789);
nor UO_2194 (O_2194,N_45598,N_45459);
nand UO_2195 (O_2195,N_45420,N_46832);
or UO_2196 (O_2196,N_48330,N_48382);
and UO_2197 (O_2197,N_47045,N_47487);
xnor UO_2198 (O_2198,N_47016,N_49389);
nor UO_2199 (O_2199,N_49852,N_46575);
and UO_2200 (O_2200,N_46792,N_48618);
and UO_2201 (O_2201,N_46931,N_45005);
nand UO_2202 (O_2202,N_45932,N_48745);
nand UO_2203 (O_2203,N_48026,N_47380);
or UO_2204 (O_2204,N_48180,N_48609);
and UO_2205 (O_2205,N_46184,N_48142);
nand UO_2206 (O_2206,N_49177,N_47695);
nor UO_2207 (O_2207,N_49181,N_48577);
nor UO_2208 (O_2208,N_47852,N_47573);
and UO_2209 (O_2209,N_45229,N_48612);
and UO_2210 (O_2210,N_48686,N_48218);
and UO_2211 (O_2211,N_49900,N_47481);
or UO_2212 (O_2212,N_45122,N_45536);
or UO_2213 (O_2213,N_46562,N_45827);
and UO_2214 (O_2214,N_47546,N_49090);
nand UO_2215 (O_2215,N_48825,N_45290);
nand UO_2216 (O_2216,N_45419,N_46563);
or UO_2217 (O_2217,N_45601,N_46910);
nand UO_2218 (O_2218,N_49384,N_47981);
nor UO_2219 (O_2219,N_47687,N_49952);
xnor UO_2220 (O_2220,N_48616,N_49668);
nor UO_2221 (O_2221,N_48591,N_46435);
and UO_2222 (O_2222,N_49178,N_48818);
or UO_2223 (O_2223,N_49412,N_48392);
nor UO_2224 (O_2224,N_48513,N_45986);
nand UO_2225 (O_2225,N_48425,N_45620);
and UO_2226 (O_2226,N_45454,N_49889);
and UO_2227 (O_2227,N_47870,N_48799);
nand UO_2228 (O_2228,N_49698,N_48958);
xor UO_2229 (O_2229,N_46990,N_47559);
nand UO_2230 (O_2230,N_45413,N_47858);
or UO_2231 (O_2231,N_47399,N_48964);
or UO_2232 (O_2232,N_49241,N_48974);
nor UO_2233 (O_2233,N_48169,N_49202);
or UO_2234 (O_2234,N_48022,N_46014);
nor UO_2235 (O_2235,N_48766,N_48752);
nand UO_2236 (O_2236,N_49843,N_49405);
nor UO_2237 (O_2237,N_45045,N_46735);
and UO_2238 (O_2238,N_47813,N_46593);
nand UO_2239 (O_2239,N_45259,N_45521);
and UO_2240 (O_2240,N_47507,N_46343);
xor UO_2241 (O_2241,N_48813,N_45553);
xnor UO_2242 (O_2242,N_45165,N_45307);
and UO_2243 (O_2243,N_45550,N_49888);
xor UO_2244 (O_2244,N_47744,N_48402);
nand UO_2245 (O_2245,N_47091,N_46379);
nor UO_2246 (O_2246,N_46236,N_48450);
nand UO_2247 (O_2247,N_47458,N_45291);
xnor UO_2248 (O_2248,N_46246,N_49235);
xor UO_2249 (O_2249,N_47918,N_49187);
and UO_2250 (O_2250,N_49935,N_46689);
nor UO_2251 (O_2251,N_48869,N_46595);
nand UO_2252 (O_2252,N_48236,N_49569);
nor UO_2253 (O_2253,N_47204,N_49566);
nor UO_2254 (O_2254,N_45178,N_46586);
and UO_2255 (O_2255,N_48525,N_47905);
nor UO_2256 (O_2256,N_45513,N_46362);
and UO_2257 (O_2257,N_48749,N_46938);
xnor UO_2258 (O_2258,N_45755,N_49363);
or UO_2259 (O_2259,N_46079,N_46864);
nand UO_2260 (O_2260,N_48335,N_45009);
or UO_2261 (O_2261,N_48407,N_45296);
or UO_2262 (O_2262,N_49586,N_47388);
nand UO_2263 (O_2263,N_45761,N_48232);
nand UO_2264 (O_2264,N_47543,N_49311);
nor UO_2265 (O_2265,N_49495,N_46494);
nor UO_2266 (O_2266,N_49876,N_49649);
nor UO_2267 (O_2267,N_45862,N_45722);
and UO_2268 (O_2268,N_47588,N_45025);
nor UO_2269 (O_2269,N_45350,N_49925);
nand UO_2270 (O_2270,N_45405,N_48213);
nor UO_2271 (O_2271,N_49392,N_48710);
and UO_2272 (O_2272,N_48233,N_47784);
and UO_2273 (O_2273,N_49931,N_47728);
or UO_2274 (O_2274,N_48356,N_45511);
xnor UO_2275 (O_2275,N_45676,N_45246);
nor UO_2276 (O_2276,N_46057,N_49559);
nor UO_2277 (O_2277,N_45899,N_45067);
nor UO_2278 (O_2278,N_48018,N_46351);
or UO_2279 (O_2279,N_45640,N_47110);
and UO_2280 (O_2280,N_46158,N_47242);
and UO_2281 (O_2281,N_46871,N_48788);
and UO_2282 (O_2282,N_49928,N_47936);
and UO_2283 (O_2283,N_49857,N_47229);
and UO_2284 (O_2284,N_45082,N_48624);
or UO_2285 (O_2285,N_45407,N_49557);
nor UO_2286 (O_2286,N_47010,N_48214);
or UO_2287 (O_2287,N_47182,N_46819);
and UO_2288 (O_2288,N_46663,N_45379);
and UO_2289 (O_2289,N_46809,N_45496);
and UO_2290 (O_2290,N_49853,N_49147);
or UO_2291 (O_2291,N_46154,N_48586);
and UO_2292 (O_2292,N_47448,N_46830);
nand UO_2293 (O_2293,N_49637,N_45228);
or UO_2294 (O_2294,N_45030,N_48301);
or UO_2295 (O_2295,N_45238,N_45013);
or UO_2296 (O_2296,N_48033,N_47627);
nand UO_2297 (O_2297,N_46148,N_45810);
or UO_2298 (O_2298,N_47508,N_45586);
and UO_2299 (O_2299,N_48905,N_47063);
and UO_2300 (O_2300,N_46880,N_45957);
nand UO_2301 (O_2301,N_48851,N_49096);
nor UO_2302 (O_2302,N_46536,N_48061);
nor UO_2303 (O_2303,N_45516,N_48969);
or UO_2304 (O_2304,N_46037,N_46781);
and UO_2305 (O_2305,N_48841,N_47051);
nand UO_2306 (O_2306,N_46738,N_47948);
nor UO_2307 (O_2307,N_48581,N_48079);
and UO_2308 (O_2308,N_48599,N_49234);
or UO_2309 (O_2309,N_47647,N_47824);
and UO_2310 (O_2310,N_46599,N_47154);
or UO_2311 (O_2311,N_47032,N_48992);
nor UO_2312 (O_2312,N_47212,N_48696);
and UO_2313 (O_2313,N_46709,N_48777);
or UO_2314 (O_2314,N_48713,N_48564);
nand UO_2315 (O_2315,N_46288,N_49580);
and UO_2316 (O_2316,N_45216,N_49659);
and UO_2317 (O_2317,N_48414,N_47535);
or UO_2318 (O_2318,N_45260,N_46514);
xnor UO_2319 (O_2319,N_48127,N_48829);
xor UO_2320 (O_2320,N_49682,N_49755);
nand UO_2321 (O_2321,N_46568,N_48920);
nor UO_2322 (O_2322,N_46159,N_47690);
or UO_2323 (O_2323,N_47572,N_46957);
nor UO_2324 (O_2324,N_48802,N_45854);
nand UO_2325 (O_2325,N_45765,N_47512);
xor UO_2326 (O_2326,N_47779,N_49762);
and UO_2327 (O_2327,N_46743,N_49827);
and UO_2328 (O_2328,N_46603,N_45742);
and UO_2329 (O_2329,N_49965,N_46918);
and UO_2330 (O_2330,N_46360,N_49371);
or UO_2331 (O_2331,N_47693,N_48464);
and UO_2332 (O_2332,N_47593,N_48332);
nand UO_2333 (O_2333,N_46009,N_47490);
nand UO_2334 (O_2334,N_49783,N_49512);
or UO_2335 (O_2335,N_48558,N_47312);
and UO_2336 (O_2336,N_48957,N_46567);
nor UO_2337 (O_2337,N_49939,N_48737);
nor UO_2338 (O_2338,N_49879,N_45231);
and UO_2339 (O_2339,N_49850,N_48741);
or UO_2340 (O_2340,N_46047,N_48530);
or UO_2341 (O_2341,N_45225,N_48007);
nor UO_2342 (O_2342,N_48226,N_46190);
and UO_2343 (O_2343,N_49484,N_48506);
nand UO_2344 (O_2344,N_48837,N_46851);
xnor UO_2345 (O_2345,N_45079,N_46666);
and UO_2346 (O_2346,N_49807,N_45501);
and UO_2347 (O_2347,N_46924,N_48433);
and UO_2348 (O_2348,N_46403,N_46407);
or UO_2349 (O_2349,N_49703,N_47420);
nand UO_2350 (O_2350,N_46720,N_45710);
nor UO_2351 (O_2351,N_48800,N_46564);
and UO_2352 (O_2352,N_49950,N_49594);
or UO_2353 (O_2353,N_49220,N_48255);
xor UO_2354 (O_2354,N_46459,N_45780);
nand UO_2355 (O_2355,N_46776,N_49973);
nand UO_2356 (O_2356,N_46697,N_47943);
and UO_2357 (O_2357,N_47614,N_47823);
nand UO_2358 (O_2358,N_48429,N_45985);
xnor UO_2359 (O_2359,N_46713,N_48456);
and UO_2360 (O_2360,N_47457,N_45319);
xor UO_2361 (O_2361,N_45280,N_45264);
or UO_2362 (O_2362,N_49250,N_46755);
nor UO_2363 (O_2363,N_45529,N_46291);
and UO_2364 (O_2364,N_48694,N_49155);
or UO_2365 (O_2365,N_45308,N_48338);
or UO_2366 (O_2366,N_46481,N_46601);
nand UO_2367 (O_2367,N_49873,N_45630);
and UO_2368 (O_2368,N_49238,N_46341);
nand UO_2369 (O_2369,N_49954,N_46252);
nor UO_2370 (O_2370,N_46767,N_48540);
nor UO_2371 (O_2371,N_45596,N_48875);
nor UO_2372 (O_2372,N_47455,N_48283);
nand UO_2373 (O_2373,N_46574,N_47401);
nor UO_2374 (O_2374,N_47994,N_49138);
or UO_2375 (O_2375,N_49379,N_49457);
nand UO_2376 (O_2376,N_45381,N_47964);
and UO_2377 (O_2377,N_48819,N_48709);
nand UO_2378 (O_2378,N_49545,N_48955);
or UO_2379 (O_2379,N_47471,N_49118);
or UO_2380 (O_2380,N_46632,N_48563);
nand UO_2381 (O_2381,N_48653,N_46066);
or UO_2382 (O_2382,N_45898,N_48293);
or UO_2383 (O_2383,N_46261,N_48243);
nand UO_2384 (O_2384,N_46664,N_46325);
and UO_2385 (O_2385,N_46321,N_47833);
or UO_2386 (O_2386,N_49005,N_49535);
xnor UO_2387 (O_2387,N_47042,N_46837);
or UO_2388 (O_2388,N_47039,N_47989);
xor UO_2389 (O_2389,N_46329,N_46438);
and UO_2390 (O_2390,N_48312,N_47580);
or UO_2391 (O_2391,N_49504,N_48719);
or UO_2392 (O_2392,N_45683,N_48859);
and UO_2393 (O_2393,N_49387,N_49266);
or UO_2394 (O_2394,N_49656,N_46820);
nor UO_2395 (O_2395,N_49441,N_48904);
nor UO_2396 (O_2396,N_46234,N_45689);
nand UO_2397 (O_2397,N_47597,N_45871);
or UO_2398 (O_2398,N_49990,N_48680);
nand UO_2399 (O_2399,N_45486,N_47363);
or UO_2400 (O_2400,N_47556,N_47984);
nand UO_2401 (O_2401,N_47571,N_48375);
or UO_2402 (O_2402,N_48963,N_48742);
and UO_2403 (O_2403,N_48486,N_47192);
nand UO_2404 (O_2404,N_49354,N_47462);
nor UO_2405 (O_2405,N_46879,N_47023);
xor UO_2406 (O_2406,N_47397,N_46589);
nor UO_2407 (O_2407,N_47530,N_49115);
and UO_2408 (O_2408,N_48903,N_48466);
nand UO_2409 (O_2409,N_46969,N_45342);
nor UO_2410 (O_2410,N_47531,N_48831);
nand UO_2411 (O_2411,N_46136,N_47652);
xor UO_2412 (O_2412,N_47692,N_48331);
and UO_2413 (O_2413,N_47551,N_45414);
and UO_2414 (O_2414,N_49669,N_45142);
and UO_2415 (O_2415,N_46055,N_48812);
nand UO_2416 (O_2416,N_47291,N_45793);
or UO_2417 (O_2417,N_49251,N_49222);
and UO_2418 (O_2418,N_46768,N_45204);
nand UO_2419 (O_2419,N_46959,N_45750);
or UO_2420 (O_2420,N_48009,N_45215);
nor UO_2421 (O_2421,N_47178,N_47327);
and UO_2422 (O_2422,N_49349,N_47970);
and UO_2423 (O_2423,N_49242,N_47030);
or UO_2424 (O_2424,N_45797,N_49350);
nand UO_2425 (O_2425,N_47969,N_47235);
nand UO_2426 (O_2426,N_47347,N_49280);
or UO_2427 (O_2427,N_48094,N_45866);
or UO_2428 (O_2428,N_46324,N_46301);
xnor UO_2429 (O_2429,N_46200,N_45693);
nand UO_2430 (O_2430,N_46086,N_49180);
xor UO_2431 (O_2431,N_49296,N_47761);
and UO_2432 (O_2432,N_46163,N_49678);
nor UO_2433 (O_2433,N_46051,N_45617);
xnor UO_2434 (O_2434,N_46146,N_46685);
nand UO_2435 (O_2435,N_46160,N_47592);
or UO_2436 (O_2436,N_46470,N_48337);
nor UO_2437 (O_2437,N_45373,N_46390);
nand UO_2438 (O_2438,N_49634,N_47604);
nand UO_2439 (O_2439,N_45048,N_48221);
xnor UO_2440 (O_2440,N_45410,N_49060);
or UO_2441 (O_2441,N_47133,N_46195);
nor UO_2442 (O_2442,N_48660,N_48711);
and UO_2443 (O_2443,N_47908,N_48894);
xor UO_2444 (O_2444,N_48421,N_46280);
and UO_2445 (O_2445,N_48186,N_46327);
nand UO_2446 (O_2446,N_48864,N_45626);
nor UO_2447 (O_2447,N_47084,N_48867);
and UO_2448 (O_2448,N_49936,N_48896);
and UO_2449 (O_2449,N_49776,N_47871);
nand UO_2450 (O_2450,N_49277,N_49820);
nor UO_2451 (O_2451,N_46050,N_45445);
nor UO_2452 (O_2452,N_49714,N_47729);
and UO_2453 (O_2453,N_49711,N_47142);
and UO_2454 (O_2454,N_46845,N_47679);
or UO_2455 (O_2455,N_45947,N_45759);
nand UO_2456 (O_2456,N_46203,N_47509);
nand UO_2457 (O_2457,N_46539,N_46579);
nand UO_2458 (O_2458,N_49707,N_47179);
nand UO_2459 (O_2459,N_47130,N_47454);
nand UO_2460 (O_2460,N_46221,N_45723);
nand UO_2461 (O_2461,N_49432,N_49972);
and UO_2462 (O_2462,N_48933,N_47826);
and UO_2463 (O_2463,N_46411,N_45707);
and UO_2464 (O_2464,N_45734,N_47348);
nor UO_2465 (O_2465,N_49124,N_49778);
nor UO_2466 (O_2466,N_47665,N_46505);
nand UO_2467 (O_2467,N_47491,N_46683);
nand UO_2468 (O_2468,N_45256,N_45931);
nand UO_2469 (O_2469,N_45492,N_46424);
nand UO_2470 (O_2470,N_48855,N_48796);
and UO_2471 (O_2471,N_47293,N_48058);
or UO_2472 (O_2472,N_49838,N_45461);
nor UO_2473 (O_2473,N_48501,N_49477);
nand UO_2474 (O_2474,N_49818,N_45774);
nor UO_2475 (O_2475,N_46948,N_48743);
or UO_2476 (O_2476,N_45532,N_47921);
nor UO_2477 (O_2477,N_47365,N_49037);
nor UO_2478 (O_2478,N_46433,N_48069);
nor UO_2479 (O_2479,N_48611,N_45310);
nor UO_2480 (O_2480,N_48740,N_48479);
nor UO_2481 (O_2481,N_49875,N_48845);
nand UO_2482 (O_2482,N_46016,N_47207);
nand UO_2483 (O_2483,N_46923,N_46929);
and UO_2484 (O_2484,N_45125,N_46890);
xor UO_2485 (O_2485,N_47252,N_45037);
and UO_2486 (O_2486,N_46660,N_45047);
xor UO_2487 (O_2487,N_49855,N_46520);
and UO_2488 (O_2488,N_49225,N_46843);
nand UO_2489 (O_2489,N_46609,N_47382);
and UO_2490 (O_2490,N_48509,N_46936);
and UO_2491 (O_2491,N_48342,N_45772);
nor UO_2492 (O_2492,N_49770,N_49112);
nor UO_2493 (O_2493,N_45552,N_48553);
and UO_2494 (O_2494,N_47174,N_48419);
nand UO_2495 (O_2495,N_46149,N_48804);
or UO_2496 (O_2496,N_45612,N_49455);
nand UO_2497 (O_2497,N_45998,N_48483);
or UO_2498 (O_2498,N_47238,N_49959);
nand UO_2499 (O_2499,N_47369,N_48118);
nand UO_2500 (O_2500,N_48548,N_46068);
and UO_2501 (O_2501,N_46359,N_48604);
and UO_2502 (O_2502,N_46950,N_46120);
nand UO_2503 (O_2503,N_45935,N_48796);
nor UO_2504 (O_2504,N_49761,N_47875);
and UO_2505 (O_2505,N_49897,N_49610);
and UO_2506 (O_2506,N_45772,N_49537);
nor UO_2507 (O_2507,N_45362,N_46545);
and UO_2508 (O_2508,N_48866,N_47410);
and UO_2509 (O_2509,N_47072,N_48743);
nor UO_2510 (O_2510,N_45792,N_46874);
or UO_2511 (O_2511,N_49858,N_47545);
xor UO_2512 (O_2512,N_45288,N_47383);
nor UO_2513 (O_2513,N_47116,N_45135);
nor UO_2514 (O_2514,N_46381,N_45610);
nand UO_2515 (O_2515,N_49144,N_47871);
nand UO_2516 (O_2516,N_47124,N_48767);
nor UO_2517 (O_2517,N_48719,N_46810);
or UO_2518 (O_2518,N_49265,N_47774);
nor UO_2519 (O_2519,N_45232,N_47098);
nor UO_2520 (O_2520,N_49182,N_45881);
nand UO_2521 (O_2521,N_48929,N_46091);
nor UO_2522 (O_2522,N_46602,N_49331);
and UO_2523 (O_2523,N_47768,N_46091);
nand UO_2524 (O_2524,N_49143,N_48844);
and UO_2525 (O_2525,N_47556,N_46262);
nand UO_2526 (O_2526,N_47601,N_47029);
or UO_2527 (O_2527,N_49567,N_46196);
and UO_2528 (O_2528,N_45964,N_46869);
and UO_2529 (O_2529,N_46940,N_49546);
nand UO_2530 (O_2530,N_46808,N_47788);
nor UO_2531 (O_2531,N_46986,N_48143);
or UO_2532 (O_2532,N_48327,N_48681);
nand UO_2533 (O_2533,N_47671,N_46770);
nor UO_2534 (O_2534,N_47267,N_47189);
and UO_2535 (O_2535,N_48800,N_49000);
nand UO_2536 (O_2536,N_48031,N_49013);
or UO_2537 (O_2537,N_47258,N_45210);
nor UO_2538 (O_2538,N_45766,N_45410);
xor UO_2539 (O_2539,N_46516,N_45821);
and UO_2540 (O_2540,N_46407,N_48568);
and UO_2541 (O_2541,N_49250,N_48680);
nor UO_2542 (O_2542,N_49140,N_49525);
nand UO_2543 (O_2543,N_48164,N_47677);
or UO_2544 (O_2544,N_47821,N_46569);
or UO_2545 (O_2545,N_48279,N_47193);
nor UO_2546 (O_2546,N_48657,N_47535);
and UO_2547 (O_2547,N_49606,N_48788);
nor UO_2548 (O_2548,N_46758,N_46287);
nor UO_2549 (O_2549,N_46288,N_49394);
xnor UO_2550 (O_2550,N_49134,N_48906);
or UO_2551 (O_2551,N_48661,N_47146);
and UO_2552 (O_2552,N_49944,N_46296);
xor UO_2553 (O_2553,N_49152,N_46162);
nor UO_2554 (O_2554,N_48672,N_45319);
nand UO_2555 (O_2555,N_48267,N_47727);
or UO_2556 (O_2556,N_45318,N_48616);
nand UO_2557 (O_2557,N_46963,N_47895);
and UO_2558 (O_2558,N_49876,N_46623);
nor UO_2559 (O_2559,N_48808,N_48584);
nand UO_2560 (O_2560,N_48278,N_49936);
nor UO_2561 (O_2561,N_45859,N_47036);
nor UO_2562 (O_2562,N_48463,N_48879);
nand UO_2563 (O_2563,N_48192,N_48858);
and UO_2564 (O_2564,N_49888,N_49762);
xnor UO_2565 (O_2565,N_45113,N_46735);
nor UO_2566 (O_2566,N_48429,N_49856);
or UO_2567 (O_2567,N_48608,N_45064);
nor UO_2568 (O_2568,N_47363,N_45092);
or UO_2569 (O_2569,N_46528,N_49887);
and UO_2570 (O_2570,N_46429,N_49260);
and UO_2571 (O_2571,N_48885,N_45046);
nand UO_2572 (O_2572,N_46942,N_49317);
and UO_2573 (O_2573,N_49905,N_48189);
nand UO_2574 (O_2574,N_47411,N_45130);
nand UO_2575 (O_2575,N_45759,N_45958);
nand UO_2576 (O_2576,N_48405,N_47141);
nor UO_2577 (O_2577,N_49986,N_46032);
nor UO_2578 (O_2578,N_47802,N_47905);
nor UO_2579 (O_2579,N_46945,N_48029);
and UO_2580 (O_2580,N_49007,N_45434);
and UO_2581 (O_2581,N_45127,N_48763);
nor UO_2582 (O_2582,N_46437,N_46728);
nand UO_2583 (O_2583,N_46596,N_46077);
and UO_2584 (O_2584,N_47081,N_47183);
or UO_2585 (O_2585,N_49553,N_45422);
and UO_2586 (O_2586,N_49268,N_46128);
and UO_2587 (O_2587,N_47052,N_47593);
nand UO_2588 (O_2588,N_47924,N_47375);
or UO_2589 (O_2589,N_47883,N_48676);
nor UO_2590 (O_2590,N_47605,N_48760);
nand UO_2591 (O_2591,N_49353,N_49923);
nand UO_2592 (O_2592,N_47651,N_48340);
xor UO_2593 (O_2593,N_45427,N_45864);
nand UO_2594 (O_2594,N_49871,N_47633);
and UO_2595 (O_2595,N_46236,N_49013);
or UO_2596 (O_2596,N_47626,N_47443);
nand UO_2597 (O_2597,N_47078,N_46792);
nor UO_2598 (O_2598,N_46240,N_47810);
nand UO_2599 (O_2599,N_49677,N_45788);
nand UO_2600 (O_2600,N_45086,N_48829);
or UO_2601 (O_2601,N_49297,N_46257);
or UO_2602 (O_2602,N_48842,N_48681);
and UO_2603 (O_2603,N_49741,N_49623);
and UO_2604 (O_2604,N_49709,N_49347);
nand UO_2605 (O_2605,N_46813,N_48907);
nor UO_2606 (O_2606,N_46884,N_48273);
xnor UO_2607 (O_2607,N_49157,N_46542);
xnor UO_2608 (O_2608,N_45076,N_48932);
or UO_2609 (O_2609,N_46722,N_45983);
and UO_2610 (O_2610,N_47710,N_46901);
and UO_2611 (O_2611,N_48788,N_49965);
nor UO_2612 (O_2612,N_47648,N_49648);
or UO_2613 (O_2613,N_49830,N_45981);
or UO_2614 (O_2614,N_45681,N_46298);
xor UO_2615 (O_2615,N_45495,N_48257);
and UO_2616 (O_2616,N_49357,N_45272);
nor UO_2617 (O_2617,N_48236,N_48720);
or UO_2618 (O_2618,N_49463,N_47852);
xor UO_2619 (O_2619,N_46387,N_47029);
nand UO_2620 (O_2620,N_47496,N_45682);
nor UO_2621 (O_2621,N_49161,N_49073);
or UO_2622 (O_2622,N_45143,N_48596);
or UO_2623 (O_2623,N_48420,N_48339);
xnor UO_2624 (O_2624,N_46616,N_47235);
or UO_2625 (O_2625,N_48498,N_45382);
nand UO_2626 (O_2626,N_48458,N_45818);
nor UO_2627 (O_2627,N_47850,N_49186);
nand UO_2628 (O_2628,N_47734,N_45328);
nor UO_2629 (O_2629,N_45480,N_48556);
nor UO_2630 (O_2630,N_46674,N_48058);
or UO_2631 (O_2631,N_49470,N_49256);
nand UO_2632 (O_2632,N_47138,N_49044);
xor UO_2633 (O_2633,N_48883,N_47073);
and UO_2634 (O_2634,N_46366,N_47478);
nand UO_2635 (O_2635,N_47805,N_45555);
nor UO_2636 (O_2636,N_45213,N_49280);
nor UO_2637 (O_2637,N_46850,N_49683);
or UO_2638 (O_2638,N_48731,N_49207);
or UO_2639 (O_2639,N_45189,N_47680);
nand UO_2640 (O_2640,N_46028,N_45098);
or UO_2641 (O_2641,N_46775,N_48006);
nand UO_2642 (O_2642,N_48316,N_48594);
and UO_2643 (O_2643,N_45097,N_48556);
or UO_2644 (O_2644,N_48660,N_45728);
or UO_2645 (O_2645,N_49238,N_46135);
nand UO_2646 (O_2646,N_47316,N_48514);
nand UO_2647 (O_2647,N_46556,N_49589);
and UO_2648 (O_2648,N_49591,N_46917);
or UO_2649 (O_2649,N_47701,N_49406);
or UO_2650 (O_2650,N_48443,N_46291);
nand UO_2651 (O_2651,N_47972,N_47905);
nor UO_2652 (O_2652,N_46221,N_49072);
nor UO_2653 (O_2653,N_45590,N_48144);
and UO_2654 (O_2654,N_45104,N_45144);
or UO_2655 (O_2655,N_47616,N_48361);
nor UO_2656 (O_2656,N_47557,N_48272);
nand UO_2657 (O_2657,N_49961,N_45460);
nand UO_2658 (O_2658,N_45276,N_49306);
nor UO_2659 (O_2659,N_49159,N_47208);
xnor UO_2660 (O_2660,N_47188,N_47554);
xnor UO_2661 (O_2661,N_48384,N_48377);
or UO_2662 (O_2662,N_47201,N_46239);
nor UO_2663 (O_2663,N_45701,N_45916);
nor UO_2664 (O_2664,N_46705,N_48502);
or UO_2665 (O_2665,N_48640,N_45948);
or UO_2666 (O_2666,N_47214,N_45804);
nor UO_2667 (O_2667,N_45806,N_45711);
nor UO_2668 (O_2668,N_45291,N_45816);
or UO_2669 (O_2669,N_46578,N_45818);
nand UO_2670 (O_2670,N_45065,N_47225);
and UO_2671 (O_2671,N_48850,N_49660);
xor UO_2672 (O_2672,N_45248,N_47706);
nor UO_2673 (O_2673,N_48576,N_48173);
or UO_2674 (O_2674,N_48662,N_49902);
nor UO_2675 (O_2675,N_47398,N_48454);
and UO_2676 (O_2676,N_48605,N_45582);
nand UO_2677 (O_2677,N_45692,N_47770);
and UO_2678 (O_2678,N_49543,N_46389);
or UO_2679 (O_2679,N_49390,N_46630);
xnor UO_2680 (O_2680,N_46074,N_46267);
or UO_2681 (O_2681,N_45893,N_46133);
nor UO_2682 (O_2682,N_47559,N_46734);
or UO_2683 (O_2683,N_48178,N_49526);
nand UO_2684 (O_2684,N_45246,N_46044);
xor UO_2685 (O_2685,N_45257,N_46428);
nor UO_2686 (O_2686,N_45129,N_47328);
or UO_2687 (O_2687,N_49596,N_48824);
or UO_2688 (O_2688,N_49690,N_47884);
nor UO_2689 (O_2689,N_46193,N_45308);
nand UO_2690 (O_2690,N_49873,N_47776);
xnor UO_2691 (O_2691,N_48324,N_45241);
nor UO_2692 (O_2692,N_49645,N_49637);
and UO_2693 (O_2693,N_49317,N_46219);
or UO_2694 (O_2694,N_45711,N_48210);
nand UO_2695 (O_2695,N_48489,N_45215);
or UO_2696 (O_2696,N_47783,N_49888);
nand UO_2697 (O_2697,N_46679,N_45655);
or UO_2698 (O_2698,N_47549,N_47818);
xnor UO_2699 (O_2699,N_49326,N_45142);
and UO_2700 (O_2700,N_46925,N_47078);
nand UO_2701 (O_2701,N_47821,N_48505);
nand UO_2702 (O_2702,N_45256,N_48008);
nand UO_2703 (O_2703,N_48385,N_49289);
or UO_2704 (O_2704,N_48410,N_46448);
nand UO_2705 (O_2705,N_46999,N_46093);
and UO_2706 (O_2706,N_46093,N_47323);
nand UO_2707 (O_2707,N_45778,N_45698);
nor UO_2708 (O_2708,N_46964,N_49568);
or UO_2709 (O_2709,N_48187,N_49109);
xnor UO_2710 (O_2710,N_48301,N_45501);
xnor UO_2711 (O_2711,N_48929,N_47851);
or UO_2712 (O_2712,N_47682,N_48391);
and UO_2713 (O_2713,N_48754,N_49917);
or UO_2714 (O_2714,N_48422,N_47090);
nand UO_2715 (O_2715,N_48741,N_47580);
or UO_2716 (O_2716,N_46758,N_48539);
xnor UO_2717 (O_2717,N_46206,N_46884);
or UO_2718 (O_2718,N_49102,N_49636);
and UO_2719 (O_2719,N_45088,N_49739);
and UO_2720 (O_2720,N_47016,N_45019);
nand UO_2721 (O_2721,N_46870,N_47118);
and UO_2722 (O_2722,N_46477,N_45475);
nor UO_2723 (O_2723,N_46522,N_49860);
and UO_2724 (O_2724,N_48130,N_48728);
and UO_2725 (O_2725,N_49593,N_48241);
nor UO_2726 (O_2726,N_48326,N_46803);
or UO_2727 (O_2727,N_45088,N_46219);
nor UO_2728 (O_2728,N_47226,N_48057);
nand UO_2729 (O_2729,N_47832,N_47798);
xor UO_2730 (O_2730,N_49983,N_48015);
and UO_2731 (O_2731,N_46113,N_49768);
xor UO_2732 (O_2732,N_49630,N_49428);
or UO_2733 (O_2733,N_47285,N_47447);
or UO_2734 (O_2734,N_49911,N_49722);
or UO_2735 (O_2735,N_45598,N_45635);
and UO_2736 (O_2736,N_45194,N_47214);
xnor UO_2737 (O_2737,N_45602,N_49180);
xnor UO_2738 (O_2738,N_48506,N_49358);
nor UO_2739 (O_2739,N_47052,N_45084);
nor UO_2740 (O_2740,N_49657,N_47004);
nor UO_2741 (O_2741,N_46759,N_45552);
and UO_2742 (O_2742,N_47193,N_49942);
or UO_2743 (O_2743,N_49968,N_48114);
or UO_2744 (O_2744,N_47395,N_47845);
nand UO_2745 (O_2745,N_47885,N_47773);
or UO_2746 (O_2746,N_46533,N_45933);
nor UO_2747 (O_2747,N_46758,N_48810);
or UO_2748 (O_2748,N_49378,N_45349);
nand UO_2749 (O_2749,N_45633,N_49027);
nand UO_2750 (O_2750,N_47066,N_49282);
and UO_2751 (O_2751,N_46166,N_46566);
nor UO_2752 (O_2752,N_45993,N_46208);
or UO_2753 (O_2753,N_45529,N_47510);
nor UO_2754 (O_2754,N_45586,N_45838);
or UO_2755 (O_2755,N_46826,N_45833);
nor UO_2756 (O_2756,N_45781,N_48836);
nor UO_2757 (O_2757,N_49879,N_48496);
or UO_2758 (O_2758,N_46293,N_47565);
nand UO_2759 (O_2759,N_49305,N_48467);
and UO_2760 (O_2760,N_45517,N_46238);
xor UO_2761 (O_2761,N_49943,N_47468);
and UO_2762 (O_2762,N_45992,N_48709);
nand UO_2763 (O_2763,N_49208,N_46229);
and UO_2764 (O_2764,N_45934,N_48983);
nor UO_2765 (O_2765,N_46213,N_49987);
and UO_2766 (O_2766,N_47908,N_47979);
and UO_2767 (O_2767,N_45475,N_47943);
and UO_2768 (O_2768,N_49177,N_46702);
nand UO_2769 (O_2769,N_46813,N_46555);
and UO_2770 (O_2770,N_46858,N_49564);
and UO_2771 (O_2771,N_45392,N_49263);
nor UO_2772 (O_2772,N_45939,N_48670);
or UO_2773 (O_2773,N_47869,N_48057);
and UO_2774 (O_2774,N_48222,N_45096);
or UO_2775 (O_2775,N_47893,N_45266);
and UO_2776 (O_2776,N_47898,N_47885);
nand UO_2777 (O_2777,N_48554,N_46320);
and UO_2778 (O_2778,N_45369,N_48957);
nand UO_2779 (O_2779,N_47751,N_47705);
nor UO_2780 (O_2780,N_46013,N_45596);
nor UO_2781 (O_2781,N_45580,N_45965);
xor UO_2782 (O_2782,N_49440,N_46771);
or UO_2783 (O_2783,N_47094,N_48127);
and UO_2784 (O_2784,N_47622,N_49075);
and UO_2785 (O_2785,N_49402,N_48082);
nor UO_2786 (O_2786,N_47666,N_47935);
nor UO_2787 (O_2787,N_48064,N_45953);
nor UO_2788 (O_2788,N_47488,N_46365);
or UO_2789 (O_2789,N_45362,N_49862);
nand UO_2790 (O_2790,N_48897,N_45567);
nor UO_2791 (O_2791,N_46706,N_45902);
nor UO_2792 (O_2792,N_47336,N_49201);
and UO_2793 (O_2793,N_49259,N_48376);
xnor UO_2794 (O_2794,N_47329,N_48384);
nand UO_2795 (O_2795,N_49287,N_47449);
nand UO_2796 (O_2796,N_47984,N_49124);
or UO_2797 (O_2797,N_48298,N_48253);
nand UO_2798 (O_2798,N_48036,N_45814);
nand UO_2799 (O_2799,N_45528,N_48305);
or UO_2800 (O_2800,N_45765,N_45589);
and UO_2801 (O_2801,N_47820,N_46844);
nand UO_2802 (O_2802,N_45649,N_48174);
nor UO_2803 (O_2803,N_47883,N_49649);
and UO_2804 (O_2804,N_45397,N_46721);
and UO_2805 (O_2805,N_45493,N_45999);
or UO_2806 (O_2806,N_48334,N_48132);
nor UO_2807 (O_2807,N_49945,N_46551);
or UO_2808 (O_2808,N_48006,N_45072);
and UO_2809 (O_2809,N_48690,N_48857);
or UO_2810 (O_2810,N_47410,N_49045);
and UO_2811 (O_2811,N_49896,N_47734);
or UO_2812 (O_2812,N_47444,N_46788);
and UO_2813 (O_2813,N_49933,N_45352);
and UO_2814 (O_2814,N_48318,N_49589);
or UO_2815 (O_2815,N_46201,N_48663);
nand UO_2816 (O_2816,N_48613,N_47884);
nand UO_2817 (O_2817,N_48209,N_45329);
nor UO_2818 (O_2818,N_47563,N_48012);
xor UO_2819 (O_2819,N_48159,N_45232);
or UO_2820 (O_2820,N_45776,N_49448);
and UO_2821 (O_2821,N_46538,N_45931);
or UO_2822 (O_2822,N_47434,N_46979);
nand UO_2823 (O_2823,N_47493,N_46896);
and UO_2824 (O_2824,N_49704,N_47210);
and UO_2825 (O_2825,N_48685,N_47930);
nand UO_2826 (O_2826,N_48826,N_49053);
and UO_2827 (O_2827,N_46935,N_48628);
nand UO_2828 (O_2828,N_47009,N_49280);
xor UO_2829 (O_2829,N_46189,N_47739);
nand UO_2830 (O_2830,N_47185,N_47570);
and UO_2831 (O_2831,N_46772,N_46362);
nand UO_2832 (O_2832,N_45444,N_47966);
or UO_2833 (O_2833,N_48010,N_46138);
and UO_2834 (O_2834,N_46476,N_45849);
and UO_2835 (O_2835,N_48895,N_49895);
nor UO_2836 (O_2836,N_49877,N_46788);
nor UO_2837 (O_2837,N_47752,N_47740);
nand UO_2838 (O_2838,N_45145,N_46465);
or UO_2839 (O_2839,N_48863,N_49078);
nand UO_2840 (O_2840,N_47114,N_47609);
nor UO_2841 (O_2841,N_48837,N_49962);
nor UO_2842 (O_2842,N_45014,N_45651);
or UO_2843 (O_2843,N_45456,N_49126);
or UO_2844 (O_2844,N_46202,N_45462);
or UO_2845 (O_2845,N_45987,N_47902);
or UO_2846 (O_2846,N_48350,N_45738);
and UO_2847 (O_2847,N_46995,N_49083);
nand UO_2848 (O_2848,N_45376,N_46057);
and UO_2849 (O_2849,N_49311,N_47126);
nand UO_2850 (O_2850,N_48602,N_49669);
nand UO_2851 (O_2851,N_47781,N_46113);
nor UO_2852 (O_2852,N_46732,N_48721);
nand UO_2853 (O_2853,N_49289,N_47542);
or UO_2854 (O_2854,N_45148,N_48701);
and UO_2855 (O_2855,N_49779,N_46174);
and UO_2856 (O_2856,N_49778,N_49622);
nand UO_2857 (O_2857,N_49939,N_45598);
xnor UO_2858 (O_2858,N_46483,N_46098);
nor UO_2859 (O_2859,N_47944,N_45818);
nor UO_2860 (O_2860,N_46356,N_48670);
nor UO_2861 (O_2861,N_46577,N_47860);
and UO_2862 (O_2862,N_46651,N_45453);
and UO_2863 (O_2863,N_45775,N_49473);
and UO_2864 (O_2864,N_46514,N_48545);
xor UO_2865 (O_2865,N_47937,N_45375);
nand UO_2866 (O_2866,N_46160,N_49452);
or UO_2867 (O_2867,N_49506,N_49603);
and UO_2868 (O_2868,N_45381,N_49641);
xnor UO_2869 (O_2869,N_49897,N_46805);
and UO_2870 (O_2870,N_48677,N_47972);
nor UO_2871 (O_2871,N_48024,N_45616);
or UO_2872 (O_2872,N_45452,N_48255);
and UO_2873 (O_2873,N_49693,N_47262);
nor UO_2874 (O_2874,N_45030,N_48008);
or UO_2875 (O_2875,N_45820,N_45329);
and UO_2876 (O_2876,N_49887,N_49130);
xor UO_2877 (O_2877,N_45699,N_45738);
and UO_2878 (O_2878,N_48050,N_46994);
nor UO_2879 (O_2879,N_46541,N_48675);
and UO_2880 (O_2880,N_47586,N_45154);
nor UO_2881 (O_2881,N_45916,N_49792);
nand UO_2882 (O_2882,N_49010,N_45333);
and UO_2883 (O_2883,N_46590,N_48114);
and UO_2884 (O_2884,N_45275,N_47856);
and UO_2885 (O_2885,N_48048,N_45073);
or UO_2886 (O_2886,N_49843,N_47188);
xor UO_2887 (O_2887,N_48128,N_47124);
or UO_2888 (O_2888,N_49882,N_48843);
nand UO_2889 (O_2889,N_47189,N_46725);
nor UO_2890 (O_2890,N_49487,N_46744);
nand UO_2891 (O_2891,N_49923,N_45122);
nor UO_2892 (O_2892,N_49435,N_49959);
and UO_2893 (O_2893,N_45835,N_49530);
and UO_2894 (O_2894,N_46556,N_45329);
or UO_2895 (O_2895,N_49028,N_48077);
and UO_2896 (O_2896,N_45584,N_47396);
nand UO_2897 (O_2897,N_47133,N_49454);
nand UO_2898 (O_2898,N_49699,N_47311);
nor UO_2899 (O_2899,N_48157,N_46904);
nor UO_2900 (O_2900,N_46471,N_46066);
nor UO_2901 (O_2901,N_46885,N_45525);
nand UO_2902 (O_2902,N_46606,N_47760);
and UO_2903 (O_2903,N_48868,N_48282);
nor UO_2904 (O_2904,N_45834,N_47092);
and UO_2905 (O_2905,N_46549,N_45222);
nor UO_2906 (O_2906,N_48256,N_49568);
xnor UO_2907 (O_2907,N_46914,N_45306);
nand UO_2908 (O_2908,N_46272,N_49037);
nand UO_2909 (O_2909,N_45889,N_49798);
or UO_2910 (O_2910,N_48455,N_48135);
nand UO_2911 (O_2911,N_47955,N_45447);
nand UO_2912 (O_2912,N_48321,N_48616);
and UO_2913 (O_2913,N_48865,N_46239);
and UO_2914 (O_2914,N_46683,N_45026);
nand UO_2915 (O_2915,N_48958,N_46807);
or UO_2916 (O_2916,N_47804,N_48300);
nor UO_2917 (O_2917,N_45600,N_48412);
nand UO_2918 (O_2918,N_48582,N_45272);
nor UO_2919 (O_2919,N_48897,N_47867);
and UO_2920 (O_2920,N_49364,N_48860);
nor UO_2921 (O_2921,N_48501,N_46469);
nor UO_2922 (O_2922,N_46107,N_48303);
nor UO_2923 (O_2923,N_47328,N_46501);
and UO_2924 (O_2924,N_47180,N_45741);
and UO_2925 (O_2925,N_45772,N_45039);
xnor UO_2926 (O_2926,N_48449,N_49301);
nor UO_2927 (O_2927,N_45838,N_47827);
nand UO_2928 (O_2928,N_49201,N_47595);
nor UO_2929 (O_2929,N_46190,N_49160);
nand UO_2930 (O_2930,N_45738,N_47171);
nand UO_2931 (O_2931,N_47465,N_47612);
nand UO_2932 (O_2932,N_45318,N_45646);
and UO_2933 (O_2933,N_47941,N_46087);
nand UO_2934 (O_2934,N_46428,N_49946);
nor UO_2935 (O_2935,N_45528,N_49788);
nor UO_2936 (O_2936,N_49337,N_45020);
or UO_2937 (O_2937,N_46315,N_45506);
and UO_2938 (O_2938,N_46949,N_49921);
nor UO_2939 (O_2939,N_49722,N_48842);
or UO_2940 (O_2940,N_45336,N_48357);
nand UO_2941 (O_2941,N_48454,N_46780);
or UO_2942 (O_2942,N_48077,N_49394);
or UO_2943 (O_2943,N_47263,N_48419);
nor UO_2944 (O_2944,N_48439,N_48392);
xor UO_2945 (O_2945,N_49602,N_48453);
or UO_2946 (O_2946,N_45662,N_45303);
nor UO_2947 (O_2947,N_49844,N_46403);
nand UO_2948 (O_2948,N_46475,N_46298);
and UO_2949 (O_2949,N_48124,N_48352);
or UO_2950 (O_2950,N_47313,N_45819);
and UO_2951 (O_2951,N_45361,N_49939);
or UO_2952 (O_2952,N_46642,N_45317);
nand UO_2953 (O_2953,N_48099,N_48992);
and UO_2954 (O_2954,N_49837,N_49971);
and UO_2955 (O_2955,N_47558,N_48962);
nand UO_2956 (O_2956,N_46287,N_45823);
xor UO_2957 (O_2957,N_48296,N_47400);
nand UO_2958 (O_2958,N_46759,N_46872);
nand UO_2959 (O_2959,N_47162,N_46532);
or UO_2960 (O_2960,N_48825,N_47554);
nand UO_2961 (O_2961,N_45111,N_46366);
or UO_2962 (O_2962,N_47339,N_49204);
or UO_2963 (O_2963,N_49864,N_47953);
nor UO_2964 (O_2964,N_47651,N_48451);
nand UO_2965 (O_2965,N_46900,N_46776);
or UO_2966 (O_2966,N_47959,N_49845);
xor UO_2967 (O_2967,N_45218,N_49861);
nand UO_2968 (O_2968,N_49216,N_46439);
and UO_2969 (O_2969,N_45172,N_47251);
or UO_2970 (O_2970,N_49959,N_45183);
or UO_2971 (O_2971,N_45981,N_45059);
xnor UO_2972 (O_2972,N_46023,N_46089);
nand UO_2973 (O_2973,N_48750,N_46926);
or UO_2974 (O_2974,N_46730,N_47390);
nor UO_2975 (O_2975,N_49409,N_48493);
xor UO_2976 (O_2976,N_49667,N_49228);
and UO_2977 (O_2977,N_45140,N_48676);
and UO_2978 (O_2978,N_49803,N_46939);
and UO_2979 (O_2979,N_47883,N_45259);
or UO_2980 (O_2980,N_49475,N_47508);
nand UO_2981 (O_2981,N_46287,N_45563);
and UO_2982 (O_2982,N_49491,N_47462);
nand UO_2983 (O_2983,N_45004,N_46201);
nor UO_2984 (O_2984,N_49511,N_47896);
nor UO_2985 (O_2985,N_48761,N_45689);
or UO_2986 (O_2986,N_47057,N_45302);
and UO_2987 (O_2987,N_48930,N_46062);
or UO_2988 (O_2988,N_46386,N_45725);
or UO_2989 (O_2989,N_45807,N_47519);
and UO_2990 (O_2990,N_47720,N_45048);
nand UO_2991 (O_2991,N_45944,N_45706);
and UO_2992 (O_2992,N_46157,N_47908);
and UO_2993 (O_2993,N_45969,N_45856);
and UO_2994 (O_2994,N_49102,N_49634);
or UO_2995 (O_2995,N_47667,N_46515);
or UO_2996 (O_2996,N_47117,N_45228);
nor UO_2997 (O_2997,N_48695,N_47806);
nor UO_2998 (O_2998,N_46778,N_45784);
or UO_2999 (O_2999,N_49008,N_45403);
nand UO_3000 (O_3000,N_47958,N_48646);
or UO_3001 (O_3001,N_47841,N_45491);
nand UO_3002 (O_3002,N_48792,N_48612);
or UO_3003 (O_3003,N_45299,N_48173);
nand UO_3004 (O_3004,N_45567,N_47855);
or UO_3005 (O_3005,N_49568,N_48070);
nand UO_3006 (O_3006,N_45884,N_49448);
xnor UO_3007 (O_3007,N_49908,N_45600);
nor UO_3008 (O_3008,N_47202,N_49060);
xor UO_3009 (O_3009,N_49907,N_49676);
and UO_3010 (O_3010,N_47294,N_46911);
nor UO_3011 (O_3011,N_49190,N_45140);
or UO_3012 (O_3012,N_45216,N_45214);
xor UO_3013 (O_3013,N_49832,N_49111);
or UO_3014 (O_3014,N_49108,N_46305);
and UO_3015 (O_3015,N_47466,N_45973);
nor UO_3016 (O_3016,N_45257,N_49068);
or UO_3017 (O_3017,N_48005,N_49626);
xnor UO_3018 (O_3018,N_49315,N_45788);
nand UO_3019 (O_3019,N_46268,N_48671);
and UO_3020 (O_3020,N_45880,N_48367);
nand UO_3021 (O_3021,N_46168,N_46822);
and UO_3022 (O_3022,N_45398,N_47259);
nor UO_3023 (O_3023,N_48261,N_46251);
nand UO_3024 (O_3024,N_49173,N_48312);
nand UO_3025 (O_3025,N_49651,N_47313);
nor UO_3026 (O_3026,N_48122,N_46024);
nand UO_3027 (O_3027,N_45485,N_45186);
nor UO_3028 (O_3028,N_45859,N_48073);
nand UO_3029 (O_3029,N_47789,N_49809);
and UO_3030 (O_3030,N_48640,N_47366);
or UO_3031 (O_3031,N_46715,N_48519);
and UO_3032 (O_3032,N_45249,N_46708);
nor UO_3033 (O_3033,N_45907,N_46402);
xor UO_3034 (O_3034,N_48853,N_47179);
nor UO_3035 (O_3035,N_46915,N_47821);
or UO_3036 (O_3036,N_47791,N_46040);
or UO_3037 (O_3037,N_46467,N_48823);
xnor UO_3038 (O_3038,N_47814,N_48472);
and UO_3039 (O_3039,N_47867,N_48006);
xnor UO_3040 (O_3040,N_48145,N_47088);
and UO_3041 (O_3041,N_48911,N_49076);
nand UO_3042 (O_3042,N_45413,N_46557);
or UO_3043 (O_3043,N_48645,N_48670);
nor UO_3044 (O_3044,N_45357,N_49011);
nand UO_3045 (O_3045,N_45705,N_45231);
nand UO_3046 (O_3046,N_49145,N_45164);
or UO_3047 (O_3047,N_47385,N_47296);
and UO_3048 (O_3048,N_46467,N_47919);
and UO_3049 (O_3049,N_48738,N_46846);
nor UO_3050 (O_3050,N_47638,N_49686);
or UO_3051 (O_3051,N_47393,N_45144);
nand UO_3052 (O_3052,N_47824,N_48724);
or UO_3053 (O_3053,N_46162,N_49410);
nor UO_3054 (O_3054,N_49090,N_48202);
or UO_3055 (O_3055,N_49179,N_49298);
or UO_3056 (O_3056,N_45212,N_48524);
nand UO_3057 (O_3057,N_48135,N_48456);
and UO_3058 (O_3058,N_45680,N_48946);
xor UO_3059 (O_3059,N_47201,N_49047);
nand UO_3060 (O_3060,N_46729,N_48085);
or UO_3061 (O_3061,N_49461,N_48208);
nor UO_3062 (O_3062,N_47055,N_47676);
nand UO_3063 (O_3063,N_48565,N_48406);
nand UO_3064 (O_3064,N_45148,N_45602);
nor UO_3065 (O_3065,N_46723,N_49171);
and UO_3066 (O_3066,N_49775,N_49958);
nor UO_3067 (O_3067,N_49387,N_46499);
nand UO_3068 (O_3068,N_47594,N_46660);
or UO_3069 (O_3069,N_48251,N_49337);
nand UO_3070 (O_3070,N_47287,N_49704);
nand UO_3071 (O_3071,N_47566,N_45096);
or UO_3072 (O_3072,N_45784,N_46332);
xor UO_3073 (O_3073,N_48374,N_49135);
and UO_3074 (O_3074,N_46834,N_47811);
or UO_3075 (O_3075,N_46828,N_45939);
nor UO_3076 (O_3076,N_46314,N_45172);
nand UO_3077 (O_3077,N_46624,N_47769);
nor UO_3078 (O_3078,N_45941,N_45391);
nor UO_3079 (O_3079,N_48802,N_47869);
nand UO_3080 (O_3080,N_46801,N_47853);
nand UO_3081 (O_3081,N_45547,N_46367);
or UO_3082 (O_3082,N_48411,N_46890);
or UO_3083 (O_3083,N_49948,N_45352);
and UO_3084 (O_3084,N_45512,N_45267);
nand UO_3085 (O_3085,N_49396,N_49224);
nand UO_3086 (O_3086,N_49643,N_49308);
nand UO_3087 (O_3087,N_49483,N_46185);
xnor UO_3088 (O_3088,N_49706,N_47811);
nor UO_3089 (O_3089,N_49720,N_48548);
or UO_3090 (O_3090,N_48693,N_45301);
and UO_3091 (O_3091,N_47765,N_46362);
xnor UO_3092 (O_3092,N_47233,N_49603);
or UO_3093 (O_3093,N_45764,N_47924);
nand UO_3094 (O_3094,N_45575,N_48301);
nor UO_3095 (O_3095,N_48871,N_49878);
nand UO_3096 (O_3096,N_48930,N_49867);
nor UO_3097 (O_3097,N_49868,N_48220);
xnor UO_3098 (O_3098,N_47294,N_46204);
and UO_3099 (O_3099,N_46638,N_45775);
and UO_3100 (O_3100,N_45315,N_48329);
nor UO_3101 (O_3101,N_46566,N_46351);
or UO_3102 (O_3102,N_47450,N_45755);
and UO_3103 (O_3103,N_46429,N_46663);
nor UO_3104 (O_3104,N_48184,N_45036);
nor UO_3105 (O_3105,N_46361,N_49574);
nor UO_3106 (O_3106,N_46296,N_46148);
and UO_3107 (O_3107,N_49450,N_48833);
xnor UO_3108 (O_3108,N_47504,N_47219);
nor UO_3109 (O_3109,N_45837,N_46359);
nand UO_3110 (O_3110,N_45650,N_47765);
and UO_3111 (O_3111,N_48110,N_45351);
or UO_3112 (O_3112,N_48478,N_49751);
nand UO_3113 (O_3113,N_45422,N_47220);
nand UO_3114 (O_3114,N_46579,N_47965);
nor UO_3115 (O_3115,N_46391,N_45614);
nor UO_3116 (O_3116,N_46757,N_45841);
nor UO_3117 (O_3117,N_47089,N_47261);
or UO_3118 (O_3118,N_48449,N_45354);
nand UO_3119 (O_3119,N_45090,N_45419);
or UO_3120 (O_3120,N_46595,N_49434);
nand UO_3121 (O_3121,N_47953,N_48036);
and UO_3122 (O_3122,N_47185,N_45747);
nor UO_3123 (O_3123,N_48776,N_46769);
or UO_3124 (O_3124,N_45667,N_48864);
and UO_3125 (O_3125,N_45522,N_45899);
nor UO_3126 (O_3126,N_48844,N_45465);
nor UO_3127 (O_3127,N_45256,N_46971);
nand UO_3128 (O_3128,N_46121,N_46321);
or UO_3129 (O_3129,N_45091,N_48634);
and UO_3130 (O_3130,N_48516,N_45866);
and UO_3131 (O_3131,N_46124,N_49840);
nor UO_3132 (O_3132,N_45416,N_46843);
or UO_3133 (O_3133,N_47441,N_47995);
and UO_3134 (O_3134,N_47167,N_48441);
nor UO_3135 (O_3135,N_46565,N_45208);
nor UO_3136 (O_3136,N_48135,N_46908);
and UO_3137 (O_3137,N_49850,N_45932);
nor UO_3138 (O_3138,N_47138,N_46554);
nand UO_3139 (O_3139,N_47291,N_45628);
and UO_3140 (O_3140,N_45174,N_49917);
and UO_3141 (O_3141,N_45430,N_47533);
xnor UO_3142 (O_3142,N_47027,N_45419);
or UO_3143 (O_3143,N_49832,N_45707);
and UO_3144 (O_3144,N_49864,N_47319);
nand UO_3145 (O_3145,N_45890,N_49140);
and UO_3146 (O_3146,N_48366,N_45169);
nand UO_3147 (O_3147,N_45476,N_46450);
nand UO_3148 (O_3148,N_45462,N_49680);
nand UO_3149 (O_3149,N_48825,N_46421);
and UO_3150 (O_3150,N_47701,N_48512);
and UO_3151 (O_3151,N_48988,N_46200);
nand UO_3152 (O_3152,N_46490,N_48028);
nand UO_3153 (O_3153,N_49019,N_48530);
nor UO_3154 (O_3154,N_46687,N_47951);
and UO_3155 (O_3155,N_46567,N_45271);
xor UO_3156 (O_3156,N_46014,N_47551);
or UO_3157 (O_3157,N_49763,N_47624);
or UO_3158 (O_3158,N_48600,N_47624);
nor UO_3159 (O_3159,N_47848,N_46098);
xnor UO_3160 (O_3160,N_45427,N_46489);
nand UO_3161 (O_3161,N_48983,N_49743);
xnor UO_3162 (O_3162,N_47672,N_48203);
and UO_3163 (O_3163,N_46313,N_47648);
xor UO_3164 (O_3164,N_49103,N_49660);
nor UO_3165 (O_3165,N_49333,N_46223);
and UO_3166 (O_3166,N_47634,N_45102);
and UO_3167 (O_3167,N_46870,N_47439);
xor UO_3168 (O_3168,N_49881,N_46520);
and UO_3169 (O_3169,N_48919,N_48315);
nor UO_3170 (O_3170,N_46414,N_45197);
xnor UO_3171 (O_3171,N_46759,N_49133);
nor UO_3172 (O_3172,N_48060,N_46269);
nor UO_3173 (O_3173,N_47672,N_46729);
xor UO_3174 (O_3174,N_49987,N_48435);
or UO_3175 (O_3175,N_49382,N_46211);
nor UO_3176 (O_3176,N_46730,N_49471);
or UO_3177 (O_3177,N_49902,N_47515);
nand UO_3178 (O_3178,N_45195,N_45686);
nand UO_3179 (O_3179,N_46291,N_46979);
and UO_3180 (O_3180,N_46084,N_49088);
or UO_3181 (O_3181,N_48219,N_49802);
and UO_3182 (O_3182,N_46279,N_47020);
or UO_3183 (O_3183,N_48567,N_47108);
nand UO_3184 (O_3184,N_45110,N_48236);
and UO_3185 (O_3185,N_47574,N_49539);
xor UO_3186 (O_3186,N_45556,N_45541);
nand UO_3187 (O_3187,N_48344,N_46607);
nor UO_3188 (O_3188,N_46588,N_48332);
nand UO_3189 (O_3189,N_47148,N_46985);
nand UO_3190 (O_3190,N_46088,N_47015);
or UO_3191 (O_3191,N_49927,N_48788);
nor UO_3192 (O_3192,N_46726,N_46921);
nor UO_3193 (O_3193,N_45035,N_49963);
xnor UO_3194 (O_3194,N_48738,N_45118);
and UO_3195 (O_3195,N_46992,N_47480);
and UO_3196 (O_3196,N_49645,N_47734);
nand UO_3197 (O_3197,N_47267,N_49430);
nor UO_3198 (O_3198,N_47314,N_48600);
nand UO_3199 (O_3199,N_45824,N_47551);
nand UO_3200 (O_3200,N_49915,N_47421);
nor UO_3201 (O_3201,N_48729,N_46243);
or UO_3202 (O_3202,N_45098,N_49838);
nand UO_3203 (O_3203,N_46122,N_48534);
nor UO_3204 (O_3204,N_48283,N_46898);
nand UO_3205 (O_3205,N_47137,N_45796);
nor UO_3206 (O_3206,N_46304,N_46786);
and UO_3207 (O_3207,N_48810,N_46970);
xor UO_3208 (O_3208,N_46273,N_49335);
nand UO_3209 (O_3209,N_48412,N_46713);
and UO_3210 (O_3210,N_48892,N_46299);
nand UO_3211 (O_3211,N_48110,N_48053);
and UO_3212 (O_3212,N_47580,N_45653);
and UO_3213 (O_3213,N_45237,N_46241);
nor UO_3214 (O_3214,N_48629,N_48333);
or UO_3215 (O_3215,N_46515,N_47999);
and UO_3216 (O_3216,N_46607,N_49264);
or UO_3217 (O_3217,N_45754,N_49049);
nand UO_3218 (O_3218,N_49876,N_49503);
xnor UO_3219 (O_3219,N_47098,N_45859);
nor UO_3220 (O_3220,N_49815,N_46060);
or UO_3221 (O_3221,N_45365,N_48065);
and UO_3222 (O_3222,N_46770,N_48943);
and UO_3223 (O_3223,N_49871,N_45335);
nor UO_3224 (O_3224,N_49268,N_48553);
xor UO_3225 (O_3225,N_47965,N_47624);
and UO_3226 (O_3226,N_47019,N_49524);
nand UO_3227 (O_3227,N_47159,N_49700);
or UO_3228 (O_3228,N_47418,N_49002);
and UO_3229 (O_3229,N_47149,N_48126);
nor UO_3230 (O_3230,N_49633,N_48095);
nor UO_3231 (O_3231,N_46260,N_46828);
and UO_3232 (O_3232,N_49850,N_46406);
or UO_3233 (O_3233,N_49675,N_49769);
nor UO_3234 (O_3234,N_46893,N_48447);
and UO_3235 (O_3235,N_49814,N_45582);
and UO_3236 (O_3236,N_47390,N_49967);
nand UO_3237 (O_3237,N_49492,N_45955);
nor UO_3238 (O_3238,N_48655,N_49651);
and UO_3239 (O_3239,N_46109,N_49401);
nand UO_3240 (O_3240,N_48263,N_45056);
nand UO_3241 (O_3241,N_48427,N_47190);
nand UO_3242 (O_3242,N_47538,N_49576);
nor UO_3243 (O_3243,N_45759,N_47630);
or UO_3244 (O_3244,N_48616,N_48229);
nor UO_3245 (O_3245,N_45299,N_48594);
and UO_3246 (O_3246,N_47080,N_46243);
nor UO_3247 (O_3247,N_45772,N_45526);
nand UO_3248 (O_3248,N_46741,N_45940);
nand UO_3249 (O_3249,N_47491,N_49474);
nor UO_3250 (O_3250,N_47396,N_48010);
and UO_3251 (O_3251,N_48138,N_48698);
or UO_3252 (O_3252,N_48655,N_49381);
xnor UO_3253 (O_3253,N_46560,N_49471);
or UO_3254 (O_3254,N_47628,N_47070);
xnor UO_3255 (O_3255,N_48114,N_45146);
xnor UO_3256 (O_3256,N_46077,N_49583);
nor UO_3257 (O_3257,N_47711,N_49023);
nor UO_3258 (O_3258,N_46132,N_49770);
nor UO_3259 (O_3259,N_49125,N_47964);
xnor UO_3260 (O_3260,N_46263,N_49341);
and UO_3261 (O_3261,N_46326,N_48183);
nor UO_3262 (O_3262,N_46857,N_49878);
nand UO_3263 (O_3263,N_49699,N_48973);
xor UO_3264 (O_3264,N_49637,N_49567);
and UO_3265 (O_3265,N_45337,N_47358);
nor UO_3266 (O_3266,N_45162,N_45904);
or UO_3267 (O_3267,N_45482,N_47049);
or UO_3268 (O_3268,N_45794,N_48164);
or UO_3269 (O_3269,N_48749,N_45108);
or UO_3270 (O_3270,N_46043,N_48768);
or UO_3271 (O_3271,N_48421,N_46298);
or UO_3272 (O_3272,N_46676,N_49218);
nand UO_3273 (O_3273,N_45400,N_46993);
nand UO_3274 (O_3274,N_46596,N_48529);
or UO_3275 (O_3275,N_46088,N_48971);
nor UO_3276 (O_3276,N_47586,N_48946);
and UO_3277 (O_3277,N_45916,N_48596);
and UO_3278 (O_3278,N_47624,N_46408);
nand UO_3279 (O_3279,N_45121,N_46412);
nor UO_3280 (O_3280,N_47625,N_48340);
nand UO_3281 (O_3281,N_48084,N_47996);
nand UO_3282 (O_3282,N_47155,N_47567);
nand UO_3283 (O_3283,N_47094,N_49031);
or UO_3284 (O_3284,N_46408,N_48651);
nand UO_3285 (O_3285,N_48206,N_47118);
or UO_3286 (O_3286,N_48036,N_46312);
and UO_3287 (O_3287,N_45304,N_45203);
and UO_3288 (O_3288,N_46268,N_49199);
nand UO_3289 (O_3289,N_47558,N_49649);
and UO_3290 (O_3290,N_49521,N_49978);
nor UO_3291 (O_3291,N_47492,N_47939);
or UO_3292 (O_3292,N_46353,N_48201);
xnor UO_3293 (O_3293,N_49787,N_48202);
nand UO_3294 (O_3294,N_46242,N_47000);
nand UO_3295 (O_3295,N_49226,N_47092);
nand UO_3296 (O_3296,N_48104,N_48189);
nor UO_3297 (O_3297,N_49231,N_45133);
nand UO_3298 (O_3298,N_48255,N_48411);
nand UO_3299 (O_3299,N_48735,N_46467);
and UO_3300 (O_3300,N_46867,N_47033);
or UO_3301 (O_3301,N_49002,N_47221);
and UO_3302 (O_3302,N_46684,N_49159);
xor UO_3303 (O_3303,N_47434,N_46730);
nor UO_3304 (O_3304,N_45495,N_46423);
or UO_3305 (O_3305,N_45691,N_49208);
and UO_3306 (O_3306,N_46675,N_48350);
or UO_3307 (O_3307,N_45355,N_45812);
or UO_3308 (O_3308,N_48065,N_47945);
nand UO_3309 (O_3309,N_48120,N_46505);
nand UO_3310 (O_3310,N_46017,N_49532);
or UO_3311 (O_3311,N_48498,N_46542);
or UO_3312 (O_3312,N_48677,N_47539);
nand UO_3313 (O_3313,N_46569,N_47012);
nand UO_3314 (O_3314,N_47872,N_49281);
and UO_3315 (O_3315,N_46514,N_47700);
nand UO_3316 (O_3316,N_47831,N_45628);
nor UO_3317 (O_3317,N_45368,N_47686);
and UO_3318 (O_3318,N_46557,N_45774);
or UO_3319 (O_3319,N_46910,N_49103);
nand UO_3320 (O_3320,N_49630,N_46058);
and UO_3321 (O_3321,N_49546,N_48566);
and UO_3322 (O_3322,N_49043,N_45388);
nor UO_3323 (O_3323,N_49796,N_45923);
nand UO_3324 (O_3324,N_45986,N_45273);
xor UO_3325 (O_3325,N_47117,N_49485);
nand UO_3326 (O_3326,N_46800,N_49659);
nor UO_3327 (O_3327,N_49349,N_45599);
nor UO_3328 (O_3328,N_46605,N_48509);
nand UO_3329 (O_3329,N_47452,N_46789);
nor UO_3330 (O_3330,N_47043,N_45567);
and UO_3331 (O_3331,N_47419,N_46603);
nor UO_3332 (O_3332,N_47982,N_48802);
or UO_3333 (O_3333,N_46831,N_45066);
or UO_3334 (O_3334,N_45594,N_49505);
nor UO_3335 (O_3335,N_47517,N_49239);
xnor UO_3336 (O_3336,N_48947,N_48767);
and UO_3337 (O_3337,N_47588,N_46571);
and UO_3338 (O_3338,N_46435,N_49404);
nor UO_3339 (O_3339,N_48464,N_48648);
and UO_3340 (O_3340,N_47983,N_45442);
nand UO_3341 (O_3341,N_45838,N_48490);
nand UO_3342 (O_3342,N_47828,N_46964);
or UO_3343 (O_3343,N_46052,N_48297);
nor UO_3344 (O_3344,N_46255,N_45070);
and UO_3345 (O_3345,N_48125,N_49581);
nand UO_3346 (O_3346,N_45696,N_47324);
nor UO_3347 (O_3347,N_47671,N_49363);
xor UO_3348 (O_3348,N_47485,N_48371);
and UO_3349 (O_3349,N_47881,N_47808);
and UO_3350 (O_3350,N_47653,N_48385);
or UO_3351 (O_3351,N_45660,N_49734);
nor UO_3352 (O_3352,N_45656,N_45380);
nand UO_3353 (O_3353,N_49307,N_46324);
and UO_3354 (O_3354,N_45172,N_47863);
nor UO_3355 (O_3355,N_49794,N_45673);
nand UO_3356 (O_3356,N_45245,N_49617);
and UO_3357 (O_3357,N_46515,N_45171);
and UO_3358 (O_3358,N_45300,N_46160);
and UO_3359 (O_3359,N_46395,N_49261);
xnor UO_3360 (O_3360,N_47816,N_48829);
xnor UO_3361 (O_3361,N_49749,N_49617);
and UO_3362 (O_3362,N_49234,N_45832);
and UO_3363 (O_3363,N_45603,N_45424);
or UO_3364 (O_3364,N_46689,N_47546);
nand UO_3365 (O_3365,N_45203,N_45928);
nor UO_3366 (O_3366,N_47086,N_46668);
nand UO_3367 (O_3367,N_47764,N_47770);
nand UO_3368 (O_3368,N_47329,N_49971);
nand UO_3369 (O_3369,N_45438,N_46599);
nor UO_3370 (O_3370,N_49808,N_45372);
xor UO_3371 (O_3371,N_47331,N_49699);
nand UO_3372 (O_3372,N_49725,N_48109);
or UO_3373 (O_3373,N_48446,N_45518);
nand UO_3374 (O_3374,N_46393,N_48001);
nand UO_3375 (O_3375,N_48078,N_45622);
nand UO_3376 (O_3376,N_47594,N_47618);
nand UO_3377 (O_3377,N_48947,N_45770);
or UO_3378 (O_3378,N_45978,N_47388);
and UO_3379 (O_3379,N_47516,N_47569);
and UO_3380 (O_3380,N_48827,N_45289);
nor UO_3381 (O_3381,N_46091,N_47368);
xor UO_3382 (O_3382,N_48665,N_48070);
or UO_3383 (O_3383,N_49671,N_49166);
xnor UO_3384 (O_3384,N_46558,N_46700);
nand UO_3385 (O_3385,N_47997,N_48965);
and UO_3386 (O_3386,N_47497,N_48383);
and UO_3387 (O_3387,N_48598,N_46969);
and UO_3388 (O_3388,N_48308,N_48845);
nor UO_3389 (O_3389,N_48993,N_49649);
nand UO_3390 (O_3390,N_46423,N_48716);
xnor UO_3391 (O_3391,N_48013,N_49729);
nor UO_3392 (O_3392,N_46289,N_48902);
or UO_3393 (O_3393,N_48471,N_46246);
or UO_3394 (O_3394,N_45282,N_46302);
and UO_3395 (O_3395,N_46283,N_48586);
xor UO_3396 (O_3396,N_48836,N_45707);
nor UO_3397 (O_3397,N_49641,N_45992);
nor UO_3398 (O_3398,N_49839,N_47730);
nor UO_3399 (O_3399,N_48837,N_49227);
and UO_3400 (O_3400,N_48914,N_45293);
xor UO_3401 (O_3401,N_47337,N_45568);
and UO_3402 (O_3402,N_47453,N_47844);
nand UO_3403 (O_3403,N_45074,N_49568);
or UO_3404 (O_3404,N_49771,N_45685);
and UO_3405 (O_3405,N_48668,N_48319);
nor UO_3406 (O_3406,N_46113,N_46899);
nor UO_3407 (O_3407,N_45621,N_46835);
nor UO_3408 (O_3408,N_46722,N_47832);
or UO_3409 (O_3409,N_48257,N_46050);
nor UO_3410 (O_3410,N_46078,N_48946);
nor UO_3411 (O_3411,N_49441,N_45242);
and UO_3412 (O_3412,N_49279,N_46242);
nor UO_3413 (O_3413,N_47759,N_46110);
or UO_3414 (O_3414,N_49046,N_49625);
and UO_3415 (O_3415,N_46070,N_49003);
xor UO_3416 (O_3416,N_48448,N_46475);
or UO_3417 (O_3417,N_48522,N_45242);
and UO_3418 (O_3418,N_46189,N_45495);
xnor UO_3419 (O_3419,N_49061,N_48082);
and UO_3420 (O_3420,N_46556,N_45050);
and UO_3421 (O_3421,N_46818,N_49308);
nor UO_3422 (O_3422,N_47933,N_49525);
or UO_3423 (O_3423,N_47037,N_47188);
nand UO_3424 (O_3424,N_47126,N_49410);
xnor UO_3425 (O_3425,N_46393,N_47112);
nor UO_3426 (O_3426,N_45553,N_48573);
nand UO_3427 (O_3427,N_46476,N_48481);
xor UO_3428 (O_3428,N_46731,N_45563);
nand UO_3429 (O_3429,N_49406,N_49483);
xnor UO_3430 (O_3430,N_48057,N_47841);
and UO_3431 (O_3431,N_48286,N_48034);
and UO_3432 (O_3432,N_48022,N_49144);
nand UO_3433 (O_3433,N_45561,N_45189);
or UO_3434 (O_3434,N_46046,N_49792);
or UO_3435 (O_3435,N_48593,N_46852);
nor UO_3436 (O_3436,N_47809,N_49433);
and UO_3437 (O_3437,N_49645,N_48503);
xor UO_3438 (O_3438,N_45671,N_48034);
xor UO_3439 (O_3439,N_48596,N_45349);
or UO_3440 (O_3440,N_45545,N_47613);
or UO_3441 (O_3441,N_45697,N_45669);
xor UO_3442 (O_3442,N_46088,N_49147);
or UO_3443 (O_3443,N_47157,N_47031);
nor UO_3444 (O_3444,N_47789,N_47842);
nand UO_3445 (O_3445,N_47781,N_47526);
nand UO_3446 (O_3446,N_45878,N_45223);
nor UO_3447 (O_3447,N_47874,N_49864);
and UO_3448 (O_3448,N_49427,N_48709);
nor UO_3449 (O_3449,N_47663,N_46779);
or UO_3450 (O_3450,N_48499,N_48601);
nand UO_3451 (O_3451,N_49315,N_48415);
nor UO_3452 (O_3452,N_48545,N_46453);
nand UO_3453 (O_3453,N_45348,N_47003);
and UO_3454 (O_3454,N_45747,N_49887);
nand UO_3455 (O_3455,N_46098,N_46306);
nor UO_3456 (O_3456,N_46772,N_48731);
and UO_3457 (O_3457,N_48130,N_46708);
nor UO_3458 (O_3458,N_45581,N_47507);
or UO_3459 (O_3459,N_46021,N_47896);
and UO_3460 (O_3460,N_49501,N_46654);
nand UO_3461 (O_3461,N_47808,N_49750);
and UO_3462 (O_3462,N_48156,N_45457);
nand UO_3463 (O_3463,N_46352,N_48497);
or UO_3464 (O_3464,N_46946,N_45346);
and UO_3465 (O_3465,N_47762,N_46870);
nand UO_3466 (O_3466,N_45507,N_49431);
and UO_3467 (O_3467,N_46308,N_48840);
nand UO_3468 (O_3468,N_48472,N_49665);
and UO_3469 (O_3469,N_49917,N_45436);
or UO_3470 (O_3470,N_47012,N_45553);
and UO_3471 (O_3471,N_45267,N_45463);
or UO_3472 (O_3472,N_45888,N_46168);
nor UO_3473 (O_3473,N_49720,N_46143);
or UO_3474 (O_3474,N_45185,N_47409);
nand UO_3475 (O_3475,N_47277,N_46735);
nand UO_3476 (O_3476,N_46620,N_45781);
nand UO_3477 (O_3477,N_47006,N_48130);
or UO_3478 (O_3478,N_48615,N_45611);
nand UO_3479 (O_3479,N_47899,N_48628);
nand UO_3480 (O_3480,N_48795,N_45112);
xor UO_3481 (O_3481,N_45525,N_45984);
or UO_3482 (O_3482,N_48106,N_46726);
and UO_3483 (O_3483,N_46858,N_47363);
xnor UO_3484 (O_3484,N_48353,N_45290);
and UO_3485 (O_3485,N_45126,N_46716);
or UO_3486 (O_3486,N_45242,N_48947);
or UO_3487 (O_3487,N_48122,N_45278);
nand UO_3488 (O_3488,N_48007,N_45314);
nor UO_3489 (O_3489,N_45649,N_47073);
and UO_3490 (O_3490,N_46080,N_49717);
nand UO_3491 (O_3491,N_48598,N_45165);
xor UO_3492 (O_3492,N_48495,N_49633);
nand UO_3493 (O_3493,N_48300,N_47169);
and UO_3494 (O_3494,N_48501,N_48751);
nand UO_3495 (O_3495,N_48150,N_45151);
nand UO_3496 (O_3496,N_46192,N_46954);
nand UO_3497 (O_3497,N_45910,N_48620);
or UO_3498 (O_3498,N_48366,N_45606);
or UO_3499 (O_3499,N_45229,N_46868);
and UO_3500 (O_3500,N_46261,N_47403);
nand UO_3501 (O_3501,N_46887,N_46236);
or UO_3502 (O_3502,N_46099,N_49231);
nand UO_3503 (O_3503,N_45919,N_47870);
xnor UO_3504 (O_3504,N_45401,N_45479);
or UO_3505 (O_3505,N_49151,N_45017);
nor UO_3506 (O_3506,N_45131,N_46894);
or UO_3507 (O_3507,N_48397,N_45259);
or UO_3508 (O_3508,N_45206,N_46326);
nor UO_3509 (O_3509,N_48745,N_45790);
nand UO_3510 (O_3510,N_47410,N_48494);
nor UO_3511 (O_3511,N_48404,N_46726);
and UO_3512 (O_3512,N_46788,N_46454);
or UO_3513 (O_3513,N_45401,N_49641);
nor UO_3514 (O_3514,N_47171,N_49117);
nor UO_3515 (O_3515,N_47387,N_49068);
nand UO_3516 (O_3516,N_48042,N_47123);
or UO_3517 (O_3517,N_46270,N_48247);
nand UO_3518 (O_3518,N_46172,N_49569);
nor UO_3519 (O_3519,N_48613,N_48293);
and UO_3520 (O_3520,N_45781,N_46920);
nand UO_3521 (O_3521,N_47830,N_46532);
and UO_3522 (O_3522,N_46105,N_49882);
or UO_3523 (O_3523,N_48751,N_47626);
and UO_3524 (O_3524,N_46857,N_49279);
and UO_3525 (O_3525,N_48973,N_48761);
nor UO_3526 (O_3526,N_49863,N_46561);
and UO_3527 (O_3527,N_47330,N_45218);
nor UO_3528 (O_3528,N_48620,N_45737);
or UO_3529 (O_3529,N_45619,N_46769);
and UO_3530 (O_3530,N_48952,N_49342);
or UO_3531 (O_3531,N_45800,N_47581);
or UO_3532 (O_3532,N_48967,N_47446);
nand UO_3533 (O_3533,N_45357,N_46638);
or UO_3534 (O_3534,N_48298,N_49358);
xnor UO_3535 (O_3535,N_45012,N_47193);
nor UO_3536 (O_3536,N_49068,N_47975);
xor UO_3537 (O_3537,N_48434,N_49732);
nor UO_3538 (O_3538,N_45430,N_49935);
nor UO_3539 (O_3539,N_45809,N_49224);
or UO_3540 (O_3540,N_47447,N_47194);
and UO_3541 (O_3541,N_45884,N_48174);
and UO_3542 (O_3542,N_47445,N_48000);
nor UO_3543 (O_3543,N_46360,N_45954);
nor UO_3544 (O_3544,N_46647,N_45905);
xnor UO_3545 (O_3545,N_45192,N_45311);
or UO_3546 (O_3546,N_48686,N_45012);
nor UO_3547 (O_3547,N_46654,N_47181);
or UO_3548 (O_3548,N_49716,N_48629);
nor UO_3549 (O_3549,N_45697,N_48913);
nor UO_3550 (O_3550,N_46892,N_49172);
or UO_3551 (O_3551,N_47766,N_47774);
and UO_3552 (O_3552,N_47940,N_48465);
nand UO_3553 (O_3553,N_49289,N_45007);
nand UO_3554 (O_3554,N_48607,N_48480);
and UO_3555 (O_3555,N_47758,N_45735);
and UO_3556 (O_3556,N_49017,N_46789);
xor UO_3557 (O_3557,N_47202,N_47415);
or UO_3558 (O_3558,N_46274,N_45209);
and UO_3559 (O_3559,N_49363,N_46072);
and UO_3560 (O_3560,N_49649,N_46773);
or UO_3561 (O_3561,N_48284,N_45039);
xor UO_3562 (O_3562,N_48362,N_47170);
nand UO_3563 (O_3563,N_47445,N_47713);
or UO_3564 (O_3564,N_46350,N_45612);
nor UO_3565 (O_3565,N_45571,N_48622);
and UO_3566 (O_3566,N_48119,N_49455);
nand UO_3567 (O_3567,N_48575,N_48714);
nor UO_3568 (O_3568,N_48835,N_45551);
nand UO_3569 (O_3569,N_49426,N_47919);
nand UO_3570 (O_3570,N_49921,N_48142);
or UO_3571 (O_3571,N_45651,N_48788);
xor UO_3572 (O_3572,N_46949,N_45170);
or UO_3573 (O_3573,N_45186,N_45148);
and UO_3574 (O_3574,N_45679,N_47893);
nand UO_3575 (O_3575,N_48205,N_45012);
or UO_3576 (O_3576,N_45632,N_48922);
and UO_3577 (O_3577,N_48186,N_49281);
nor UO_3578 (O_3578,N_49704,N_47309);
nand UO_3579 (O_3579,N_45661,N_47940);
or UO_3580 (O_3580,N_48045,N_46417);
nand UO_3581 (O_3581,N_45806,N_45555);
and UO_3582 (O_3582,N_49859,N_47642);
nand UO_3583 (O_3583,N_49818,N_45958);
and UO_3584 (O_3584,N_47491,N_48002);
and UO_3585 (O_3585,N_48233,N_49159);
nand UO_3586 (O_3586,N_45438,N_45788);
or UO_3587 (O_3587,N_46475,N_45718);
nand UO_3588 (O_3588,N_49057,N_46665);
and UO_3589 (O_3589,N_46740,N_45217);
nand UO_3590 (O_3590,N_48443,N_45828);
and UO_3591 (O_3591,N_47157,N_48019);
nor UO_3592 (O_3592,N_45364,N_45241);
nor UO_3593 (O_3593,N_48413,N_45256);
nor UO_3594 (O_3594,N_49969,N_45313);
and UO_3595 (O_3595,N_47258,N_47441);
and UO_3596 (O_3596,N_46143,N_45124);
and UO_3597 (O_3597,N_45320,N_49576);
xor UO_3598 (O_3598,N_47999,N_48362);
and UO_3599 (O_3599,N_47980,N_46860);
nor UO_3600 (O_3600,N_48116,N_47908);
nand UO_3601 (O_3601,N_48046,N_48163);
nand UO_3602 (O_3602,N_47903,N_48653);
nor UO_3603 (O_3603,N_45864,N_46816);
or UO_3604 (O_3604,N_49115,N_49654);
and UO_3605 (O_3605,N_47346,N_49220);
nand UO_3606 (O_3606,N_47664,N_46814);
or UO_3607 (O_3607,N_48167,N_45084);
and UO_3608 (O_3608,N_49686,N_45163);
or UO_3609 (O_3609,N_49917,N_46999);
nor UO_3610 (O_3610,N_45467,N_48995);
or UO_3611 (O_3611,N_45122,N_48831);
and UO_3612 (O_3612,N_45624,N_45930);
nand UO_3613 (O_3613,N_45132,N_45023);
nor UO_3614 (O_3614,N_48298,N_46724);
nor UO_3615 (O_3615,N_45539,N_48731);
or UO_3616 (O_3616,N_45751,N_47019);
and UO_3617 (O_3617,N_47198,N_49562);
or UO_3618 (O_3618,N_47184,N_45385);
xnor UO_3619 (O_3619,N_49548,N_46327);
and UO_3620 (O_3620,N_49782,N_47772);
xor UO_3621 (O_3621,N_48665,N_49499);
xnor UO_3622 (O_3622,N_47449,N_48080);
xor UO_3623 (O_3623,N_45432,N_48028);
nor UO_3624 (O_3624,N_47867,N_48374);
nor UO_3625 (O_3625,N_49050,N_48789);
and UO_3626 (O_3626,N_46607,N_45342);
xor UO_3627 (O_3627,N_49445,N_48882);
and UO_3628 (O_3628,N_45191,N_49029);
nor UO_3629 (O_3629,N_46860,N_45203);
nor UO_3630 (O_3630,N_46888,N_45413);
and UO_3631 (O_3631,N_48476,N_45912);
or UO_3632 (O_3632,N_49081,N_47246);
nor UO_3633 (O_3633,N_46594,N_48202);
nor UO_3634 (O_3634,N_45317,N_46662);
nand UO_3635 (O_3635,N_45717,N_48832);
xor UO_3636 (O_3636,N_46875,N_49856);
or UO_3637 (O_3637,N_47746,N_46389);
or UO_3638 (O_3638,N_46017,N_49054);
xor UO_3639 (O_3639,N_46443,N_49477);
and UO_3640 (O_3640,N_49030,N_47646);
and UO_3641 (O_3641,N_45289,N_48246);
nor UO_3642 (O_3642,N_48215,N_46029);
nor UO_3643 (O_3643,N_46594,N_46619);
or UO_3644 (O_3644,N_47609,N_47981);
nor UO_3645 (O_3645,N_45587,N_49805);
xor UO_3646 (O_3646,N_49116,N_49945);
nand UO_3647 (O_3647,N_49724,N_45906);
and UO_3648 (O_3648,N_46591,N_46077);
nand UO_3649 (O_3649,N_48492,N_48283);
xnor UO_3650 (O_3650,N_47495,N_47567);
and UO_3651 (O_3651,N_45989,N_46735);
or UO_3652 (O_3652,N_48405,N_48315);
nand UO_3653 (O_3653,N_45725,N_48559);
and UO_3654 (O_3654,N_48980,N_48501);
nand UO_3655 (O_3655,N_47056,N_48947);
or UO_3656 (O_3656,N_48402,N_47338);
xor UO_3657 (O_3657,N_48104,N_46258);
or UO_3658 (O_3658,N_49469,N_49563);
xnor UO_3659 (O_3659,N_46461,N_48561);
or UO_3660 (O_3660,N_49653,N_48832);
nand UO_3661 (O_3661,N_46554,N_48915);
xor UO_3662 (O_3662,N_47579,N_47394);
xnor UO_3663 (O_3663,N_46890,N_45976);
nor UO_3664 (O_3664,N_46482,N_45770);
xnor UO_3665 (O_3665,N_47412,N_48400);
nand UO_3666 (O_3666,N_47450,N_47762);
and UO_3667 (O_3667,N_49151,N_48244);
or UO_3668 (O_3668,N_49988,N_47997);
nor UO_3669 (O_3669,N_47266,N_48525);
or UO_3670 (O_3670,N_49843,N_47624);
nor UO_3671 (O_3671,N_46848,N_48758);
nor UO_3672 (O_3672,N_47450,N_48937);
and UO_3673 (O_3673,N_49076,N_47554);
xnor UO_3674 (O_3674,N_45684,N_47979);
nor UO_3675 (O_3675,N_48679,N_47853);
xor UO_3676 (O_3676,N_46805,N_49768);
nor UO_3677 (O_3677,N_49251,N_49522);
or UO_3678 (O_3678,N_47874,N_45627);
nor UO_3679 (O_3679,N_49211,N_49907);
nor UO_3680 (O_3680,N_48625,N_48163);
nand UO_3681 (O_3681,N_47055,N_46749);
xnor UO_3682 (O_3682,N_48595,N_48537);
nand UO_3683 (O_3683,N_47477,N_45140);
nor UO_3684 (O_3684,N_46587,N_47765);
nor UO_3685 (O_3685,N_48726,N_48616);
nor UO_3686 (O_3686,N_48550,N_49762);
nor UO_3687 (O_3687,N_49903,N_47457);
and UO_3688 (O_3688,N_48249,N_49897);
or UO_3689 (O_3689,N_48926,N_48331);
nor UO_3690 (O_3690,N_45329,N_49251);
nor UO_3691 (O_3691,N_48282,N_46146);
or UO_3692 (O_3692,N_46482,N_49315);
xor UO_3693 (O_3693,N_47996,N_49184);
and UO_3694 (O_3694,N_48179,N_46035);
and UO_3695 (O_3695,N_48201,N_48475);
and UO_3696 (O_3696,N_45920,N_48955);
nand UO_3697 (O_3697,N_48724,N_47688);
and UO_3698 (O_3698,N_49353,N_45821);
and UO_3699 (O_3699,N_45107,N_47438);
nor UO_3700 (O_3700,N_49266,N_46783);
xnor UO_3701 (O_3701,N_49575,N_49654);
and UO_3702 (O_3702,N_49556,N_47672);
nand UO_3703 (O_3703,N_45665,N_49517);
xor UO_3704 (O_3704,N_46459,N_48711);
or UO_3705 (O_3705,N_46724,N_47242);
and UO_3706 (O_3706,N_47436,N_47618);
or UO_3707 (O_3707,N_47730,N_46480);
or UO_3708 (O_3708,N_49980,N_45368);
and UO_3709 (O_3709,N_49262,N_49172);
nor UO_3710 (O_3710,N_45975,N_45526);
xor UO_3711 (O_3711,N_45534,N_49129);
and UO_3712 (O_3712,N_45135,N_49231);
xnor UO_3713 (O_3713,N_47093,N_49080);
xor UO_3714 (O_3714,N_49144,N_45843);
nor UO_3715 (O_3715,N_49293,N_47180);
xnor UO_3716 (O_3716,N_45620,N_47355);
nand UO_3717 (O_3717,N_49344,N_46003);
or UO_3718 (O_3718,N_46480,N_48706);
nand UO_3719 (O_3719,N_47949,N_46923);
or UO_3720 (O_3720,N_48928,N_49292);
xnor UO_3721 (O_3721,N_45958,N_47727);
nor UO_3722 (O_3722,N_45437,N_45317);
nor UO_3723 (O_3723,N_49509,N_45440);
xor UO_3724 (O_3724,N_49350,N_45419);
and UO_3725 (O_3725,N_49860,N_47324);
or UO_3726 (O_3726,N_48461,N_48837);
or UO_3727 (O_3727,N_47664,N_46157);
or UO_3728 (O_3728,N_45751,N_47223);
nor UO_3729 (O_3729,N_45476,N_46324);
nand UO_3730 (O_3730,N_46602,N_45131);
nand UO_3731 (O_3731,N_45696,N_45797);
nand UO_3732 (O_3732,N_48835,N_49614);
and UO_3733 (O_3733,N_48655,N_45826);
xnor UO_3734 (O_3734,N_46602,N_47782);
nand UO_3735 (O_3735,N_47178,N_46084);
xnor UO_3736 (O_3736,N_48023,N_47869);
nor UO_3737 (O_3737,N_49892,N_46904);
nor UO_3738 (O_3738,N_47727,N_47367);
nor UO_3739 (O_3739,N_48101,N_49359);
or UO_3740 (O_3740,N_48889,N_49126);
and UO_3741 (O_3741,N_47534,N_45642);
nor UO_3742 (O_3742,N_48925,N_47611);
nand UO_3743 (O_3743,N_49636,N_49518);
and UO_3744 (O_3744,N_49270,N_48380);
and UO_3745 (O_3745,N_45621,N_45582);
nor UO_3746 (O_3746,N_47875,N_48449);
and UO_3747 (O_3747,N_48512,N_45559);
or UO_3748 (O_3748,N_48719,N_49325);
nand UO_3749 (O_3749,N_47062,N_46346);
nor UO_3750 (O_3750,N_46092,N_45176);
and UO_3751 (O_3751,N_49240,N_45469);
nor UO_3752 (O_3752,N_49063,N_45285);
nand UO_3753 (O_3753,N_46021,N_45321);
and UO_3754 (O_3754,N_47036,N_47100);
nand UO_3755 (O_3755,N_46162,N_48310);
nor UO_3756 (O_3756,N_47591,N_46425);
nor UO_3757 (O_3757,N_48892,N_45261);
nor UO_3758 (O_3758,N_46846,N_49196);
or UO_3759 (O_3759,N_48893,N_48389);
nand UO_3760 (O_3760,N_49041,N_49894);
xor UO_3761 (O_3761,N_47951,N_49579);
nor UO_3762 (O_3762,N_46708,N_49748);
nor UO_3763 (O_3763,N_48168,N_46412);
nand UO_3764 (O_3764,N_49871,N_48974);
nor UO_3765 (O_3765,N_46376,N_48178);
or UO_3766 (O_3766,N_48253,N_46622);
nand UO_3767 (O_3767,N_49221,N_47700);
or UO_3768 (O_3768,N_45486,N_46577);
nand UO_3769 (O_3769,N_48798,N_47954);
xor UO_3770 (O_3770,N_48280,N_47530);
xor UO_3771 (O_3771,N_45103,N_46018);
nor UO_3772 (O_3772,N_46955,N_49541);
or UO_3773 (O_3773,N_49802,N_47331);
nor UO_3774 (O_3774,N_45717,N_47800);
nor UO_3775 (O_3775,N_48042,N_46100);
and UO_3776 (O_3776,N_47920,N_45743);
xor UO_3777 (O_3777,N_48015,N_48827);
or UO_3778 (O_3778,N_49732,N_45638);
and UO_3779 (O_3779,N_46968,N_48355);
and UO_3780 (O_3780,N_45271,N_47886);
and UO_3781 (O_3781,N_46418,N_45696);
nor UO_3782 (O_3782,N_47841,N_48288);
nand UO_3783 (O_3783,N_47952,N_48651);
or UO_3784 (O_3784,N_47117,N_48496);
or UO_3785 (O_3785,N_47554,N_47954);
nor UO_3786 (O_3786,N_47509,N_48269);
nor UO_3787 (O_3787,N_47817,N_47569);
or UO_3788 (O_3788,N_47525,N_48504);
and UO_3789 (O_3789,N_47458,N_49092);
and UO_3790 (O_3790,N_45853,N_47685);
or UO_3791 (O_3791,N_46178,N_47035);
or UO_3792 (O_3792,N_49219,N_45061);
nand UO_3793 (O_3793,N_48218,N_49361);
xor UO_3794 (O_3794,N_48890,N_48320);
nor UO_3795 (O_3795,N_46856,N_48106);
or UO_3796 (O_3796,N_46976,N_47904);
nor UO_3797 (O_3797,N_48778,N_45267);
nor UO_3798 (O_3798,N_49817,N_49908);
nand UO_3799 (O_3799,N_46186,N_46169);
nor UO_3800 (O_3800,N_48128,N_49909);
and UO_3801 (O_3801,N_48812,N_48129);
nand UO_3802 (O_3802,N_45625,N_46690);
xor UO_3803 (O_3803,N_45839,N_47808);
xnor UO_3804 (O_3804,N_46876,N_48158);
or UO_3805 (O_3805,N_47100,N_49898);
or UO_3806 (O_3806,N_48528,N_49162);
xor UO_3807 (O_3807,N_49799,N_47598);
and UO_3808 (O_3808,N_46096,N_48042);
nor UO_3809 (O_3809,N_46770,N_48275);
xnor UO_3810 (O_3810,N_46378,N_49936);
and UO_3811 (O_3811,N_48318,N_48957);
nand UO_3812 (O_3812,N_49460,N_45495);
nor UO_3813 (O_3813,N_45316,N_48720);
nand UO_3814 (O_3814,N_46611,N_49124);
or UO_3815 (O_3815,N_47967,N_49460);
nor UO_3816 (O_3816,N_48637,N_45234);
nand UO_3817 (O_3817,N_46463,N_45123);
or UO_3818 (O_3818,N_46148,N_45643);
or UO_3819 (O_3819,N_45425,N_48894);
nor UO_3820 (O_3820,N_49240,N_47608);
or UO_3821 (O_3821,N_45391,N_48014);
nor UO_3822 (O_3822,N_45790,N_45021);
or UO_3823 (O_3823,N_49166,N_47677);
nor UO_3824 (O_3824,N_45296,N_46409);
nor UO_3825 (O_3825,N_45378,N_45410);
nand UO_3826 (O_3826,N_47759,N_46508);
nor UO_3827 (O_3827,N_48876,N_48767);
nand UO_3828 (O_3828,N_48369,N_46778);
nand UO_3829 (O_3829,N_48329,N_45683);
nand UO_3830 (O_3830,N_48178,N_45024);
and UO_3831 (O_3831,N_48431,N_45274);
nor UO_3832 (O_3832,N_47893,N_47832);
and UO_3833 (O_3833,N_47424,N_45735);
xor UO_3834 (O_3834,N_46577,N_49754);
or UO_3835 (O_3835,N_48827,N_48550);
nand UO_3836 (O_3836,N_49859,N_49897);
and UO_3837 (O_3837,N_47817,N_48975);
nand UO_3838 (O_3838,N_45242,N_48676);
nand UO_3839 (O_3839,N_45182,N_49520);
nor UO_3840 (O_3840,N_46428,N_46204);
nand UO_3841 (O_3841,N_47683,N_49290);
or UO_3842 (O_3842,N_49309,N_49997);
nor UO_3843 (O_3843,N_48021,N_45165);
and UO_3844 (O_3844,N_46786,N_46699);
and UO_3845 (O_3845,N_47541,N_48560);
nor UO_3846 (O_3846,N_45393,N_47208);
nand UO_3847 (O_3847,N_46807,N_48832);
nor UO_3848 (O_3848,N_49360,N_45802);
and UO_3849 (O_3849,N_45348,N_47294);
nand UO_3850 (O_3850,N_47211,N_49014);
and UO_3851 (O_3851,N_47753,N_49017);
and UO_3852 (O_3852,N_46649,N_48392);
or UO_3853 (O_3853,N_47221,N_49951);
and UO_3854 (O_3854,N_46136,N_46155);
or UO_3855 (O_3855,N_48451,N_47034);
and UO_3856 (O_3856,N_48054,N_48670);
nor UO_3857 (O_3857,N_45775,N_49450);
or UO_3858 (O_3858,N_48080,N_46854);
or UO_3859 (O_3859,N_46819,N_48484);
nor UO_3860 (O_3860,N_49025,N_49023);
xnor UO_3861 (O_3861,N_48287,N_45864);
nor UO_3862 (O_3862,N_46280,N_48105);
nand UO_3863 (O_3863,N_48934,N_45589);
and UO_3864 (O_3864,N_46125,N_46665);
or UO_3865 (O_3865,N_49503,N_47766);
and UO_3866 (O_3866,N_47272,N_46951);
nand UO_3867 (O_3867,N_46704,N_49825);
nor UO_3868 (O_3868,N_49641,N_45473);
xor UO_3869 (O_3869,N_47359,N_46780);
and UO_3870 (O_3870,N_45043,N_45216);
nand UO_3871 (O_3871,N_45681,N_47881);
and UO_3872 (O_3872,N_46015,N_45330);
and UO_3873 (O_3873,N_45820,N_49931);
nor UO_3874 (O_3874,N_47737,N_48729);
xor UO_3875 (O_3875,N_49153,N_48938);
and UO_3876 (O_3876,N_48647,N_46850);
and UO_3877 (O_3877,N_49738,N_49240);
xor UO_3878 (O_3878,N_48543,N_45936);
nand UO_3879 (O_3879,N_49075,N_47762);
nor UO_3880 (O_3880,N_45872,N_46874);
and UO_3881 (O_3881,N_47445,N_49654);
nor UO_3882 (O_3882,N_47836,N_45041);
nand UO_3883 (O_3883,N_48144,N_47322);
and UO_3884 (O_3884,N_48632,N_48765);
nor UO_3885 (O_3885,N_46040,N_45800);
nor UO_3886 (O_3886,N_49644,N_48822);
and UO_3887 (O_3887,N_48649,N_49407);
xor UO_3888 (O_3888,N_47162,N_45005);
and UO_3889 (O_3889,N_45943,N_48560);
nor UO_3890 (O_3890,N_48706,N_49053);
nor UO_3891 (O_3891,N_49642,N_46626);
and UO_3892 (O_3892,N_47507,N_46462);
and UO_3893 (O_3893,N_48728,N_46885);
and UO_3894 (O_3894,N_45352,N_47102);
and UO_3895 (O_3895,N_47749,N_46556);
or UO_3896 (O_3896,N_49671,N_46066);
and UO_3897 (O_3897,N_48914,N_45927);
and UO_3898 (O_3898,N_46349,N_47605);
nor UO_3899 (O_3899,N_46560,N_47722);
or UO_3900 (O_3900,N_45299,N_47576);
or UO_3901 (O_3901,N_49068,N_48891);
nand UO_3902 (O_3902,N_49129,N_49471);
and UO_3903 (O_3903,N_47043,N_49154);
and UO_3904 (O_3904,N_46364,N_48743);
or UO_3905 (O_3905,N_45008,N_49359);
and UO_3906 (O_3906,N_46181,N_49697);
nand UO_3907 (O_3907,N_46819,N_46594);
nor UO_3908 (O_3908,N_46092,N_49883);
xnor UO_3909 (O_3909,N_45061,N_49874);
and UO_3910 (O_3910,N_48488,N_45916);
nor UO_3911 (O_3911,N_48130,N_47687);
and UO_3912 (O_3912,N_48156,N_48337);
nand UO_3913 (O_3913,N_46007,N_47526);
nand UO_3914 (O_3914,N_46543,N_47772);
xnor UO_3915 (O_3915,N_48106,N_47935);
nand UO_3916 (O_3916,N_49217,N_47941);
and UO_3917 (O_3917,N_46585,N_45087);
xnor UO_3918 (O_3918,N_49159,N_48624);
nand UO_3919 (O_3919,N_45887,N_46555);
nor UO_3920 (O_3920,N_49596,N_45740);
nand UO_3921 (O_3921,N_46129,N_45266);
xnor UO_3922 (O_3922,N_46104,N_46271);
nor UO_3923 (O_3923,N_48317,N_45101);
and UO_3924 (O_3924,N_45998,N_49023);
or UO_3925 (O_3925,N_46843,N_46022);
nand UO_3926 (O_3926,N_47459,N_45680);
nand UO_3927 (O_3927,N_47690,N_45776);
xor UO_3928 (O_3928,N_47168,N_46647);
xor UO_3929 (O_3929,N_49940,N_48246);
nand UO_3930 (O_3930,N_47348,N_46193);
nand UO_3931 (O_3931,N_47321,N_48439);
and UO_3932 (O_3932,N_49330,N_45975);
or UO_3933 (O_3933,N_49433,N_47822);
and UO_3934 (O_3934,N_48331,N_45957);
or UO_3935 (O_3935,N_49276,N_49433);
nand UO_3936 (O_3936,N_46462,N_48414);
and UO_3937 (O_3937,N_46772,N_45361);
or UO_3938 (O_3938,N_48045,N_46921);
nor UO_3939 (O_3939,N_48860,N_48822);
or UO_3940 (O_3940,N_46577,N_46710);
and UO_3941 (O_3941,N_45031,N_45870);
nor UO_3942 (O_3942,N_46098,N_46198);
nand UO_3943 (O_3943,N_45845,N_48248);
or UO_3944 (O_3944,N_45472,N_47025);
and UO_3945 (O_3945,N_49926,N_47021);
or UO_3946 (O_3946,N_48831,N_45567);
nand UO_3947 (O_3947,N_48843,N_47781);
xor UO_3948 (O_3948,N_45067,N_46481);
and UO_3949 (O_3949,N_45199,N_48650);
and UO_3950 (O_3950,N_49692,N_47699);
and UO_3951 (O_3951,N_47494,N_47165);
nand UO_3952 (O_3952,N_47852,N_47598);
nor UO_3953 (O_3953,N_49197,N_45062);
nand UO_3954 (O_3954,N_45144,N_45488);
nand UO_3955 (O_3955,N_46012,N_47097);
and UO_3956 (O_3956,N_48927,N_47237);
or UO_3957 (O_3957,N_48913,N_49748);
nand UO_3958 (O_3958,N_49215,N_47798);
and UO_3959 (O_3959,N_45498,N_47925);
or UO_3960 (O_3960,N_47291,N_45557);
or UO_3961 (O_3961,N_48799,N_46130);
and UO_3962 (O_3962,N_45239,N_45892);
nor UO_3963 (O_3963,N_45358,N_46815);
xor UO_3964 (O_3964,N_45347,N_45419);
nand UO_3965 (O_3965,N_49750,N_47196);
or UO_3966 (O_3966,N_49636,N_45452);
nand UO_3967 (O_3967,N_45291,N_45589);
nor UO_3968 (O_3968,N_45356,N_45493);
or UO_3969 (O_3969,N_46790,N_47386);
nor UO_3970 (O_3970,N_49850,N_48268);
and UO_3971 (O_3971,N_47030,N_46421);
and UO_3972 (O_3972,N_45614,N_48890);
and UO_3973 (O_3973,N_48649,N_49456);
nand UO_3974 (O_3974,N_48221,N_48865);
nand UO_3975 (O_3975,N_47099,N_46311);
and UO_3976 (O_3976,N_48158,N_49257);
and UO_3977 (O_3977,N_45073,N_49234);
or UO_3978 (O_3978,N_46646,N_47117);
and UO_3979 (O_3979,N_45129,N_49483);
and UO_3980 (O_3980,N_49519,N_45371);
and UO_3981 (O_3981,N_48395,N_45812);
nand UO_3982 (O_3982,N_49011,N_48946);
xnor UO_3983 (O_3983,N_48769,N_47867);
nor UO_3984 (O_3984,N_47591,N_48259);
or UO_3985 (O_3985,N_45640,N_47073);
nor UO_3986 (O_3986,N_47418,N_49732);
nor UO_3987 (O_3987,N_45073,N_49219);
nor UO_3988 (O_3988,N_49585,N_46739);
or UO_3989 (O_3989,N_45664,N_45835);
nor UO_3990 (O_3990,N_47842,N_45225);
nor UO_3991 (O_3991,N_46380,N_49720);
nor UO_3992 (O_3992,N_45882,N_45899);
nor UO_3993 (O_3993,N_48691,N_48431);
nand UO_3994 (O_3994,N_49772,N_45205);
or UO_3995 (O_3995,N_45997,N_48268);
nand UO_3996 (O_3996,N_49575,N_49095);
or UO_3997 (O_3997,N_47650,N_45328);
or UO_3998 (O_3998,N_46534,N_49711);
nand UO_3999 (O_3999,N_47912,N_49556);
nor UO_4000 (O_4000,N_45354,N_47272);
nand UO_4001 (O_4001,N_47132,N_45713);
and UO_4002 (O_4002,N_47721,N_47737);
nor UO_4003 (O_4003,N_45125,N_46868);
nand UO_4004 (O_4004,N_49933,N_45618);
nand UO_4005 (O_4005,N_47232,N_46195);
and UO_4006 (O_4006,N_45662,N_46617);
nand UO_4007 (O_4007,N_45318,N_49416);
xor UO_4008 (O_4008,N_49957,N_47850);
and UO_4009 (O_4009,N_48337,N_47288);
and UO_4010 (O_4010,N_49822,N_45779);
nand UO_4011 (O_4011,N_46268,N_48418);
or UO_4012 (O_4012,N_46442,N_48804);
nor UO_4013 (O_4013,N_46626,N_45067);
nand UO_4014 (O_4014,N_49025,N_49629);
or UO_4015 (O_4015,N_49670,N_47416);
xnor UO_4016 (O_4016,N_48230,N_46875);
nand UO_4017 (O_4017,N_48435,N_46639);
nor UO_4018 (O_4018,N_46376,N_49369);
or UO_4019 (O_4019,N_49514,N_47196);
nor UO_4020 (O_4020,N_45816,N_48819);
and UO_4021 (O_4021,N_45893,N_48742);
nand UO_4022 (O_4022,N_45995,N_45888);
nor UO_4023 (O_4023,N_47046,N_49408);
nor UO_4024 (O_4024,N_46431,N_45476);
and UO_4025 (O_4025,N_47265,N_47857);
and UO_4026 (O_4026,N_48547,N_45471);
and UO_4027 (O_4027,N_47487,N_47011);
nand UO_4028 (O_4028,N_48330,N_48105);
and UO_4029 (O_4029,N_48441,N_46576);
nor UO_4030 (O_4030,N_47491,N_46545);
nand UO_4031 (O_4031,N_49390,N_46922);
and UO_4032 (O_4032,N_49865,N_49016);
nor UO_4033 (O_4033,N_47460,N_49436);
xor UO_4034 (O_4034,N_48292,N_49166);
xnor UO_4035 (O_4035,N_49189,N_47471);
nor UO_4036 (O_4036,N_45150,N_48484);
or UO_4037 (O_4037,N_45248,N_47585);
xor UO_4038 (O_4038,N_46420,N_47546);
nand UO_4039 (O_4039,N_47130,N_47581);
and UO_4040 (O_4040,N_47932,N_46639);
nand UO_4041 (O_4041,N_48775,N_49745);
nor UO_4042 (O_4042,N_46320,N_45119);
and UO_4043 (O_4043,N_46535,N_47935);
or UO_4044 (O_4044,N_47306,N_45662);
and UO_4045 (O_4045,N_47901,N_45940);
nor UO_4046 (O_4046,N_46312,N_45600);
nand UO_4047 (O_4047,N_46606,N_45425);
nand UO_4048 (O_4048,N_45651,N_49683);
nor UO_4049 (O_4049,N_45870,N_49453);
nor UO_4050 (O_4050,N_46622,N_49446);
nor UO_4051 (O_4051,N_47718,N_47004);
nor UO_4052 (O_4052,N_47735,N_45737);
nand UO_4053 (O_4053,N_49500,N_47522);
nand UO_4054 (O_4054,N_47235,N_47027);
and UO_4055 (O_4055,N_49730,N_49935);
or UO_4056 (O_4056,N_48109,N_48778);
or UO_4057 (O_4057,N_46719,N_48036);
nor UO_4058 (O_4058,N_47917,N_47118);
or UO_4059 (O_4059,N_45759,N_48086);
nor UO_4060 (O_4060,N_47007,N_45736);
and UO_4061 (O_4061,N_46455,N_47132);
nand UO_4062 (O_4062,N_49541,N_49471);
nand UO_4063 (O_4063,N_48929,N_49230);
nand UO_4064 (O_4064,N_47359,N_49824);
and UO_4065 (O_4065,N_48723,N_48590);
or UO_4066 (O_4066,N_48273,N_45065);
or UO_4067 (O_4067,N_47076,N_48899);
and UO_4068 (O_4068,N_49025,N_46189);
nand UO_4069 (O_4069,N_45724,N_49455);
or UO_4070 (O_4070,N_47049,N_47550);
and UO_4071 (O_4071,N_48296,N_47326);
nor UO_4072 (O_4072,N_47891,N_46785);
nor UO_4073 (O_4073,N_45465,N_46586);
nand UO_4074 (O_4074,N_49302,N_49683);
nor UO_4075 (O_4075,N_46230,N_46655);
or UO_4076 (O_4076,N_45796,N_47698);
xor UO_4077 (O_4077,N_49283,N_46150);
nand UO_4078 (O_4078,N_45234,N_47028);
nor UO_4079 (O_4079,N_45393,N_47248);
and UO_4080 (O_4080,N_48382,N_49644);
and UO_4081 (O_4081,N_45992,N_46008);
and UO_4082 (O_4082,N_48447,N_45830);
nand UO_4083 (O_4083,N_45437,N_46709);
nand UO_4084 (O_4084,N_49795,N_49135);
nand UO_4085 (O_4085,N_48960,N_46887);
nor UO_4086 (O_4086,N_46334,N_45657);
and UO_4087 (O_4087,N_46296,N_48164);
nor UO_4088 (O_4088,N_48245,N_48479);
and UO_4089 (O_4089,N_47363,N_49586);
nor UO_4090 (O_4090,N_45265,N_45541);
nor UO_4091 (O_4091,N_49005,N_45645);
and UO_4092 (O_4092,N_45424,N_46906);
and UO_4093 (O_4093,N_45716,N_47885);
nand UO_4094 (O_4094,N_45108,N_48036);
or UO_4095 (O_4095,N_45238,N_48156);
or UO_4096 (O_4096,N_48162,N_49576);
xnor UO_4097 (O_4097,N_49486,N_45149);
xor UO_4098 (O_4098,N_49711,N_49129);
xor UO_4099 (O_4099,N_46511,N_47724);
xnor UO_4100 (O_4100,N_49666,N_49482);
nand UO_4101 (O_4101,N_45982,N_45791);
and UO_4102 (O_4102,N_48329,N_48540);
xnor UO_4103 (O_4103,N_46421,N_47201);
and UO_4104 (O_4104,N_47564,N_46553);
nand UO_4105 (O_4105,N_49175,N_48533);
xor UO_4106 (O_4106,N_48833,N_45492);
or UO_4107 (O_4107,N_45166,N_45883);
or UO_4108 (O_4108,N_47449,N_45472);
nor UO_4109 (O_4109,N_48124,N_49786);
and UO_4110 (O_4110,N_47613,N_46826);
nor UO_4111 (O_4111,N_47012,N_46421);
nor UO_4112 (O_4112,N_48690,N_46426);
nor UO_4113 (O_4113,N_46707,N_46112);
nand UO_4114 (O_4114,N_49210,N_49474);
or UO_4115 (O_4115,N_48147,N_45109);
xor UO_4116 (O_4116,N_46161,N_49580);
xnor UO_4117 (O_4117,N_45348,N_46715);
nor UO_4118 (O_4118,N_46478,N_47291);
nor UO_4119 (O_4119,N_45008,N_47048);
nand UO_4120 (O_4120,N_45452,N_46407);
or UO_4121 (O_4121,N_45746,N_46720);
nor UO_4122 (O_4122,N_45029,N_48212);
or UO_4123 (O_4123,N_49924,N_48753);
nor UO_4124 (O_4124,N_48464,N_48865);
and UO_4125 (O_4125,N_47394,N_47639);
xor UO_4126 (O_4126,N_49596,N_47914);
and UO_4127 (O_4127,N_49343,N_47512);
and UO_4128 (O_4128,N_48826,N_47228);
nand UO_4129 (O_4129,N_45946,N_49343);
nor UO_4130 (O_4130,N_47417,N_48382);
nand UO_4131 (O_4131,N_46528,N_46687);
nand UO_4132 (O_4132,N_46829,N_46742);
nand UO_4133 (O_4133,N_48146,N_46960);
xor UO_4134 (O_4134,N_49116,N_45038);
and UO_4135 (O_4135,N_46417,N_46736);
and UO_4136 (O_4136,N_49263,N_46400);
nor UO_4137 (O_4137,N_45246,N_49168);
xnor UO_4138 (O_4138,N_45813,N_49574);
and UO_4139 (O_4139,N_49193,N_46891);
nand UO_4140 (O_4140,N_45580,N_45844);
or UO_4141 (O_4141,N_46487,N_49960);
or UO_4142 (O_4142,N_46405,N_46829);
nor UO_4143 (O_4143,N_49173,N_46443);
or UO_4144 (O_4144,N_46582,N_47179);
nand UO_4145 (O_4145,N_47785,N_48349);
or UO_4146 (O_4146,N_48585,N_46150);
or UO_4147 (O_4147,N_46127,N_48660);
nand UO_4148 (O_4148,N_46598,N_47931);
nand UO_4149 (O_4149,N_47496,N_49369);
or UO_4150 (O_4150,N_49509,N_49978);
and UO_4151 (O_4151,N_45257,N_48157);
xor UO_4152 (O_4152,N_47670,N_47135);
nor UO_4153 (O_4153,N_49720,N_46274);
nand UO_4154 (O_4154,N_47771,N_47641);
and UO_4155 (O_4155,N_49221,N_45122);
xnor UO_4156 (O_4156,N_45881,N_45394);
nand UO_4157 (O_4157,N_48667,N_49352);
or UO_4158 (O_4158,N_46368,N_45712);
and UO_4159 (O_4159,N_48953,N_49368);
nand UO_4160 (O_4160,N_49539,N_46409);
and UO_4161 (O_4161,N_45770,N_46076);
nand UO_4162 (O_4162,N_49982,N_47700);
nor UO_4163 (O_4163,N_49747,N_49203);
and UO_4164 (O_4164,N_47879,N_48340);
nor UO_4165 (O_4165,N_49546,N_47879);
or UO_4166 (O_4166,N_45680,N_49408);
and UO_4167 (O_4167,N_48329,N_48642);
nor UO_4168 (O_4168,N_47104,N_45322);
nor UO_4169 (O_4169,N_47982,N_47948);
nor UO_4170 (O_4170,N_45973,N_49455);
and UO_4171 (O_4171,N_47820,N_47144);
xor UO_4172 (O_4172,N_49950,N_47155);
nor UO_4173 (O_4173,N_47129,N_45140);
nor UO_4174 (O_4174,N_48251,N_46717);
and UO_4175 (O_4175,N_48524,N_49473);
or UO_4176 (O_4176,N_47017,N_47008);
nand UO_4177 (O_4177,N_45709,N_48576);
nor UO_4178 (O_4178,N_45974,N_45049);
or UO_4179 (O_4179,N_48062,N_48815);
or UO_4180 (O_4180,N_45180,N_48730);
xnor UO_4181 (O_4181,N_48431,N_47200);
xnor UO_4182 (O_4182,N_47615,N_46654);
or UO_4183 (O_4183,N_49940,N_49023);
and UO_4184 (O_4184,N_46432,N_46247);
xor UO_4185 (O_4185,N_45922,N_48856);
xor UO_4186 (O_4186,N_47578,N_46953);
nor UO_4187 (O_4187,N_48711,N_48135);
nand UO_4188 (O_4188,N_45523,N_47323);
or UO_4189 (O_4189,N_48302,N_47679);
and UO_4190 (O_4190,N_47919,N_49553);
or UO_4191 (O_4191,N_48473,N_46137);
or UO_4192 (O_4192,N_45221,N_47076);
xnor UO_4193 (O_4193,N_49895,N_46130);
nor UO_4194 (O_4194,N_45440,N_49601);
and UO_4195 (O_4195,N_48293,N_49593);
and UO_4196 (O_4196,N_49923,N_49403);
nor UO_4197 (O_4197,N_46572,N_46325);
xnor UO_4198 (O_4198,N_49604,N_49027);
nand UO_4199 (O_4199,N_47325,N_47999);
and UO_4200 (O_4200,N_47839,N_49909);
nand UO_4201 (O_4201,N_48290,N_46750);
xnor UO_4202 (O_4202,N_49049,N_47572);
nor UO_4203 (O_4203,N_47466,N_47363);
nand UO_4204 (O_4204,N_45474,N_48246);
and UO_4205 (O_4205,N_46933,N_48362);
nand UO_4206 (O_4206,N_48201,N_48227);
or UO_4207 (O_4207,N_45535,N_48879);
nor UO_4208 (O_4208,N_46518,N_49189);
nand UO_4209 (O_4209,N_46393,N_47180);
nor UO_4210 (O_4210,N_46987,N_49830);
nand UO_4211 (O_4211,N_46494,N_45335);
xor UO_4212 (O_4212,N_46725,N_46495);
nor UO_4213 (O_4213,N_49323,N_46355);
or UO_4214 (O_4214,N_47188,N_49170);
nand UO_4215 (O_4215,N_47091,N_48205);
nor UO_4216 (O_4216,N_46720,N_49281);
nand UO_4217 (O_4217,N_45699,N_48187);
and UO_4218 (O_4218,N_48921,N_49759);
or UO_4219 (O_4219,N_47989,N_48652);
and UO_4220 (O_4220,N_49503,N_48464);
nand UO_4221 (O_4221,N_46620,N_46707);
nand UO_4222 (O_4222,N_48799,N_47868);
or UO_4223 (O_4223,N_46214,N_49386);
nand UO_4224 (O_4224,N_48800,N_45117);
nor UO_4225 (O_4225,N_45121,N_46304);
or UO_4226 (O_4226,N_45072,N_47431);
xnor UO_4227 (O_4227,N_46144,N_49940);
or UO_4228 (O_4228,N_46165,N_45881);
or UO_4229 (O_4229,N_49256,N_46758);
nor UO_4230 (O_4230,N_48396,N_49138);
nand UO_4231 (O_4231,N_49967,N_47531);
nand UO_4232 (O_4232,N_45084,N_49927);
nor UO_4233 (O_4233,N_49460,N_49738);
and UO_4234 (O_4234,N_45914,N_48598);
or UO_4235 (O_4235,N_49237,N_46262);
and UO_4236 (O_4236,N_47957,N_49416);
nor UO_4237 (O_4237,N_49780,N_46215);
nand UO_4238 (O_4238,N_48168,N_48621);
and UO_4239 (O_4239,N_48272,N_46904);
nand UO_4240 (O_4240,N_45383,N_47647);
nand UO_4241 (O_4241,N_47808,N_46044);
nand UO_4242 (O_4242,N_48954,N_47633);
nand UO_4243 (O_4243,N_46897,N_47244);
nor UO_4244 (O_4244,N_48136,N_49384);
and UO_4245 (O_4245,N_48848,N_45368);
and UO_4246 (O_4246,N_47328,N_48485);
and UO_4247 (O_4247,N_45756,N_48648);
or UO_4248 (O_4248,N_47623,N_47280);
or UO_4249 (O_4249,N_45839,N_49236);
nor UO_4250 (O_4250,N_49128,N_45968);
xor UO_4251 (O_4251,N_47809,N_46765);
nand UO_4252 (O_4252,N_47498,N_49584);
xnor UO_4253 (O_4253,N_47147,N_47320);
nor UO_4254 (O_4254,N_48289,N_47759);
or UO_4255 (O_4255,N_47173,N_48623);
or UO_4256 (O_4256,N_49823,N_45408);
xnor UO_4257 (O_4257,N_48795,N_48557);
or UO_4258 (O_4258,N_48537,N_49422);
or UO_4259 (O_4259,N_46541,N_48367);
or UO_4260 (O_4260,N_47224,N_46824);
nor UO_4261 (O_4261,N_46049,N_45170);
nor UO_4262 (O_4262,N_47632,N_48933);
nor UO_4263 (O_4263,N_46146,N_45570);
or UO_4264 (O_4264,N_49837,N_46967);
or UO_4265 (O_4265,N_45846,N_45448);
or UO_4266 (O_4266,N_46302,N_46547);
nand UO_4267 (O_4267,N_47897,N_47594);
nand UO_4268 (O_4268,N_49569,N_48064);
nor UO_4269 (O_4269,N_47217,N_46418);
and UO_4270 (O_4270,N_49597,N_47697);
or UO_4271 (O_4271,N_47581,N_48969);
nor UO_4272 (O_4272,N_47619,N_47597);
and UO_4273 (O_4273,N_48331,N_48636);
or UO_4274 (O_4274,N_46071,N_48886);
nand UO_4275 (O_4275,N_48831,N_46352);
nor UO_4276 (O_4276,N_47071,N_45817);
and UO_4277 (O_4277,N_48448,N_46850);
or UO_4278 (O_4278,N_48215,N_49370);
and UO_4279 (O_4279,N_48972,N_48106);
and UO_4280 (O_4280,N_48642,N_48396);
and UO_4281 (O_4281,N_49012,N_49955);
nor UO_4282 (O_4282,N_49266,N_45583);
nand UO_4283 (O_4283,N_46104,N_45083);
nand UO_4284 (O_4284,N_45754,N_49176);
xor UO_4285 (O_4285,N_47973,N_47201);
or UO_4286 (O_4286,N_47069,N_48753);
nor UO_4287 (O_4287,N_49641,N_47351);
or UO_4288 (O_4288,N_46224,N_46911);
xnor UO_4289 (O_4289,N_46475,N_47884);
or UO_4290 (O_4290,N_47864,N_48454);
nor UO_4291 (O_4291,N_49777,N_48594);
and UO_4292 (O_4292,N_49238,N_45704);
and UO_4293 (O_4293,N_47958,N_47108);
and UO_4294 (O_4294,N_45420,N_47180);
nand UO_4295 (O_4295,N_45409,N_48300);
nand UO_4296 (O_4296,N_45150,N_48939);
xor UO_4297 (O_4297,N_49201,N_47486);
nor UO_4298 (O_4298,N_45211,N_48137);
or UO_4299 (O_4299,N_49362,N_49873);
nand UO_4300 (O_4300,N_48655,N_47909);
and UO_4301 (O_4301,N_47552,N_47392);
or UO_4302 (O_4302,N_46849,N_47262);
nor UO_4303 (O_4303,N_48304,N_45511);
and UO_4304 (O_4304,N_45313,N_48751);
and UO_4305 (O_4305,N_46262,N_48263);
nor UO_4306 (O_4306,N_46087,N_48343);
and UO_4307 (O_4307,N_49011,N_47339);
and UO_4308 (O_4308,N_48796,N_45898);
and UO_4309 (O_4309,N_46617,N_45151);
nor UO_4310 (O_4310,N_49113,N_48683);
nor UO_4311 (O_4311,N_48250,N_47371);
nand UO_4312 (O_4312,N_45530,N_47404);
and UO_4313 (O_4313,N_45792,N_45700);
nand UO_4314 (O_4314,N_47476,N_47309);
and UO_4315 (O_4315,N_47750,N_48824);
or UO_4316 (O_4316,N_49752,N_46796);
or UO_4317 (O_4317,N_45503,N_46856);
or UO_4318 (O_4318,N_45657,N_45418);
nand UO_4319 (O_4319,N_45157,N_48072);
and UO_4320 (O_4320,N_48038,N_47087);
nor UO_4321 (O_4321,N_47007,N_46472);
or UO_4322 (O_4322,N_49797,N_48192);
nor UO_4323 (O_4323,N_46516,N_47130);
nor UO_4324 (O_4324,N_45850,N_45371);
and UO_4325 (O_4325,N_48489,N_47340);
nand UO_4326 (O_4326,N_47988,N_47502);
or UO_4327 (O_4327,N_49232,N_49536);
or UO_4328 (O_4328,N_49665,N_46171);
nand UO_4329 (O_4329,N_48553,N_49285);
and UO_4330 (O_4330,N_49846,N_46536);
xnor UO_4331 (O_4331,N_45792,N_45600);
or UO_4332 (O_4332,N_47120,N_46968);
nand UO_4333 (O_4333,N_45828,N_48100);
nand UO_4334 (O_4334,N_48519,N_46806);
or UO_4335 (O_4335,N_48887,N_46128);
and UO_4336 (O_4336,N_45460,N_46799);
nor UO_4337 (O_4337,N_48396,N_47061);
nor UO_4338 (O_4338,N_48123,N_48812);
and UO_4339 (O_4339,N_48779,N_45662);
xor UO_4340 (O_4340,N_49204,N_47439);
and UO_4341 (O_4341,N_49080,N_47111);
nor UO_4342 (O_4342,N_46254,N_48975);
or UO_4343 (O_4343,N_45490,N_46358);
nor UO_4344 (O_4344,N_45756,N_45482);
and UO_4345 (O_4345,N_49859,N_45355);
and UO_4346 (O_4346,N_48501,N_45021);
or UO_4347 (O_4347,N_45177,N_49246);
nor UO_4348 (O_4348,N_46674,N_46523);
and UO_4349 (O_4349,N_47305,N_47001);
nor UO_4350 (O_4350,N_49243,N_45729);
and UO_4351 (O_4351,N_45010,N_48583);
and UO_4352 (O_4352,N_47741,N_49577);
nor UO_4353 (O_4353,N_47703,N_47883);
or UO_4354 (O_4354,N_46946,N_46205);
xor UO_4355 (O_4355,N_48272,N_46279);
and UO_4356 (O_4356,N_49371,N_46848);
xor UO_4357 (O_4357,N_47713,N_49147);
nand UO_4358 (O_4358,N_47124,N_48678);
or UO_4359 (O_4359,N_45952,N_49128);
nor UO_4360 (O_4360,N_45097,N_45791);
and UO_4361 (O_4361,N_46541,N_48593);
nor UO_4362 (O_4362,N_45463,N_46565);
nand UO_4363 (O_4363,N_47913,N_46910);
and UO_4364 (O_4364,N_45712,N_48311);
nand UO_4365 (O_4365,N_47372,N_47930);
or UO_4366 (O_4366,N_48815,N_47295);
nand UO_4367 (O_4367,N_47257,N_46846);
nand UO_4368 (O_4368,N_48745,N_48599);
nand UO_4369 (O_4369,N_47020,N_49719);
nor UO_4370 (O_4370,N_45987,N_48978);
and UO_4371 (O_4371,N_48967,N_48624);
xor UO_4372 (O_4372,N_48883,N_46282);
and UO_4373 (O_4373,N_47632,N_49070);
or UO_4374 (O_4374,N_46593,N_49561);
xnor UO_4375 (O_4375,N_48463,N_49263);
nand UO_4376 (O_4376,N_45118,N_49506);
and UO_4377 (O_4377,N_49679,N_47685);
nor UO_4378 (O_4378,N_47505,N_48961);
or UO_4379 (O_4379,N_48115,N_47096);
nand UO_4380 (O_4380,N_48384,N_46244);
and UO_4381 (O_4381,N_45571,N_48627);
xor UO_4382 (O_4382,N_48128,N_47653);
or UO_4383 (O_4383,N_48888,N_47200);
nand UO_4384 (O_4384,N_45318,N_49591);
and UO_4385 (O_4385,N_47500,N_48620);
and UO_4386 (O_4386,N_48130,N_45891);
and UO_4387 (O_4387,N_49018,N_45652);
and UO_4388 (O_4388,N_49701,N_48348);
and UO_4389 (O_4389,N_45497,N_49747);
xor UO_4390 (O_4390,N_46536,N_45109);
and UO_4391 (O_4391,N_47962,N_49739);
and UO_4392 (O_4392,N_48968,N_48737);
and UO_4393 (O_4393,N_45282,N_45069);
xor UO_4394 (O_4394,N_46779,N_45622);
and UO_4395 (O_4395,N_49273,N_47259);
nor UO_4396 (O_4396,N_49266,N_48977);
nand UO_4397 (O_4397,N_45004,N_47950);
nor UO_4398 (O_4398,N_46626,N_46113);
nand UO_4399 (O_4399,N_45570,N_49806);
and UO_4400 (O_4400,N_46748,N_46706);
xor UO_4401 (O_4401,N_46237,N_48852);
nand UO_4402 (O_4402,N_45703,N_46916);
xnor UO_4403 (O_4403,N_47540,N_46026);
nor UO_4404 (O_4404,N_45642,N_47076);
or UO_4405 (O_4405,N_49016,N_46637);
xnor UO_4406 (O_4406,N_45985,N_49327);
and UO_4407 (O_4407,N_49012,N_45904);
nor UO_4408 (O_4408,N_48387,N_46796);
nand UO_4409 (O_4409,N_45306,N_48362);
or UO_4410 (O_4410,N_49325,N_49096);
nand UO_4411 (O_4411,N_47035,N_45271);
nor UO_4412 (O_4412,N_49056,N_48080);
nand UO_4413 (O_4413,N_46299,N_47357);
nand UO_4414 (O_4414,N_47787,N_46224);
nand UO_4415 (O_4415,N_46141,N_48707);
nor UO_4416 (O_4416,N_48824,N_46580);
nand UO_4417 (O_4417,N_49666,N_45941);
and UO_4418 (O_4418,N_45836,N_45075);
nand UO_4419 (O_4419,N_49051,N_49044);
xnor UO_4420 (O_4420,N_46144,N_49232);
nand UO_4421 (O_4421,N_48802,N_45035);
and UO_4422 (O_4422,N_45268,N_49079);
nor UO_4423 (O_4423,N_47537,N_49520);
or UO_4424 (O_4424,N_48203,N_45827);
nor UO_4425 (O_4425,N_47009,N_49026);
nand UO_4426 (O_4426,N_48300,N_48144);
nor UO_4427 (O_4427,N_46798,N_47493);
nand UO_4428 (O_4428,N_49926,N_46167);
nor UO_4429 (O_4429,N_47669,N_48447);
or UO_4430 (O_4430,N_48677,N_47112);
or UO_4431 (O_4431,N_48201,N_49942);
and UO_4432 (O_4432,N_46816,N_49257);
nand UO_4433 (O_4433,N_46823,N_45272);
nor UO_4434 (O_4434,N_49302,N_48449);
or UO_4435 (O_4435,N_48431,N_49000);
or UO_4436 (O_4436,N_46779,N_48851);
or UO_4437 (O_4437,N_48690,N_48917);
nor UO_4438 (O_4438,N_47719,N_49145);
nand UO_4439 (O_4439,N_48265,N_46587);
or UO_4440 (O_4440,N_45261,N_48245);
nand UO_4441 (O_4441,N_45951,N_49443);
and UO_4442 (O_4442,N_46696,N_49160);
and UO_4443 (O_4443,N_48072,N_47977);
nand UO_4444 (O_4444,N_47570,N_49135);
and UO_4445 (O_4445,N_48847,N_46064);
and UO_4446 (O_4446,N_46441,N_48534);
nand UO_4447 (O_4447,N_48506,N_49510);
and UO_4448 (O_4448,N_45215,N_45253);
xnor UO_4449 (O_4449,N_46361,N_45942);
or UO_4450 (O_4450,N_45997,N_46285);
or UO_4451 (O_4451,N_46720,N_46443);
or UO_4452 (O_4452,N_45949,N_49039);
xor UO_4453 (O_4453,N_49511,N_48996);
and UO_4454 (O_4454,N_45577,N_48506);
or UO_4455 (O_4455,N_46016,N_45724);
and UO_4456 (O_4456,N_46532,N_46518);
and UO_4457 (O_4457,N_48299,N_46864);
or UO_4458 (O_4458,N_47746,N_48802);
and UO_4459 (O_4459,N_48501,N_49143);
nand UO_4460 (O_4460,N_48505,N_46344);
and UO_4461 (O_4461,N_48741,N_45801);
nand UO_4462 (O_4462,N_46632,N_46382);
nand UO_4463 (O_4463,N_46028,N_49706);
nand UO_4464 (O_4464,N_48472,N_47094);
and UO_4465 (O_4465,N_45158,N_49719);
or UO_4466 (O_4466,N_45580,N_46174);
or UO_4467 (O_4467,N_46728,N_48025);
nand UO_4468 (O_4468,N_49057,N_47840);
nand UO_4469 (O_4469,N_49207,N_48036);
nor UO_4470 (O_4470,N_46446,N_46550);
nor UO_4471 (O_4471,N_46070,N_48177);
and UO_4472 (O_4472,N_47574,N_49528);
and UO_4473 (O_4473,N_47768,N_46108);
or UO_4474 (O_4474,N_47646,N_46120);
nor UO_4475 (O_4475,N_45089,N_45229);
or UO_4476 (O_4476,N_48463,N_48064);
nand UO_4477 (O_4477,N_46670,N_49003);
and UO_4478 (O_4478,N_46100,N_49910);
nor UO_4479 (O_4479,N_49356,N_49504);
nor UO_4480 (O_4480,N_45019,N_49961);
or UO_4481 (O_4481,N_45667,N_46353);
nand UO_4482 (O_4482,N_47740,N_48425);
nor UO_4483 (O_4483,N_49503,N_46300);
and UO_4484 (O_4484,N_45840,N_45253);
nand UO_4485 (O_4485,N_47236,N_49431);
and UO_4486 (O_4486,N_45032,N_49757);
and UO_4487 (O_4487,N_45739,N_48644);
and UO_4488 (O_4488,N_45973,N_46927);
or UO_4489 (O_4489,N_45600,N_45314);
or UO_4490 (O_4490,N_45550,N_47637);
and UO_4491 (O_4491,N_45721,N_48012);
or UO_4492 (O_4492,N_48960,N_49474);
and UO_4493 (O_4493,N_49856,N_45193);
and UO_4494 (O_4494,N_46306,N_46968);
or UO_4495 (O_4495,N_47197,N_48314);
or UO_4496 (O_4496,N_45881,N_49269);
nand UO_4497 (O_4497,N_48543,N_47590);
nor UO_4498 (O_4498,N_47270,N_49280);
nor UO_4499 (O_4499,N_45441,N_47170);
nand UO_4500 (O_4500,N_46139,N_48966);
nor UO_4501 (O_4501,N_48230,N_47737);
and UO_4502 (O_4502,N_46052,N_45947);
nor UO_4503 (O_4503,N_46630,N_45175);
and UO_4504 (O_4504,N_48269,N_49146);
or UO_4505 (O_4505,N_45140,N_45633);
and UO_4506 (O_4506,N_49386,N_47929);
nor UO_4507 (O_4507,N_45330,N_49959);
nor UO_4508 (O_4508,N_46105,N_46779);
nand UO_4509 (O_4509,N_45419,N_45195);
and UO_4510 (O_4510,N_45075,N_47644);
nor UO_4511 (O_4511,N_47021,N_45831);
or UO_4512 (O_4512,N_49337,N_45163);
and UO_4513 (O_4513,N_45823,N_48236);
nor UO_4514 (O_4514,N_48877,N_49217);
xnor UO_4515 (O_4515,N_49725,N_47680);
or UO_4516 (O_4516,N_46628,N_47601);
and UO_4517 (O_4517,N_47735,N_45142);
or UO_4518 (O_4518,N_47551,N_49636);
nand UO_4519 (O_4519,N_47422,N_47709);
nor UO_4520 (O_4520,N_46937,N_46128);
nor UO_4521 (O_4521,N_49195,N_48491);
or UO_4522 (O_4522,N_46298,N_47747);
and UO_4523 (O_4523,N_47666,N_48445);
and UO_4524 (O_4524,N_47066,N_45172);
or UO_4525 (O_4525,N_45763,N_49324);
or UO_4526 (O_4526,N_46788,N_48905);
or UO_4527 (O_4527,N_49076,N_48140);
or UO_4528 (O_4528,N_48157,N_49268);
or UO_4529 (O_4529,N_48924,N_47793);
and UO_4530 (O_4530,N_47786,N_45355);
nor UO_4531 (O_4531,N_48065,N_48296);
or UO_4532 (O_4532,N_49503,N_45652);
nor UO_4533 (O_4533,N_45545,N_48043);
xnor UO_4534 (O_4534,N_46323,N_48806);
or UO_4535 (O_4535,N_47834,N_47657);
xor UO_4536 (O_4536,N_49859,N_47391);
nand UO_4537 (O_4537,N_47138,N_49136);
or UO_4538 (O_4538,N_49450,N_47306);
and UO_4539 (O_4539,N_46075,N_49383);
or UO_4540 (O_4540,N_49357,N_48255);
xnor UO_4541 (O_4541,N_45744,N_45394);
or UO_4542 (O_4542,N_49797,N_47409);
xnor UO_4543 (O_4543,N_47944,N_47735);
and UO_4544 (O_4544,N_49719,N_49314);
or UO_4545 (O_4545,N_46007,N_45766);
and UO_4546 (O_4546,N_49815,N_48503);
nand UO_4547 (O_4547,N_46082,N_48178);
and UO_4548 (O_4548,N_47125,N_47254);
nor UO_4549 (O_4549,N_49081,N_45505);
xnor UO_4550 (O_4550,N_46768,N_45581);
nand UO_4551 (O_4551,N_49102,N_48334);
nand UO_4552 (O_4552,N_46622,N_49629);
or UO_4553 (O_4553,N_45338,N_49431);
nor UO_4554 (O_4554,N_45110,N_45797);
nor UO_4555 (O_4555,N_45720,N_45597);
or UO_4556 (O_4556,N_48713,N_49757);
or UO_4557 (O_4557,N_48486,N_47782);
nor UO_4558 (O_4558,N_48255,N_45487);
xor UO_4559 (O_4559,N_48384,N_48828);
xnor UO_4560 (O_4560,N_49260,N_47515);
xnor UO_4561 (O_4561,N_47683,N_46305);
or UO_4562 (O_4562,N_47969,N_45259);
nand UO_4563 (O_4563,N_46212,N_47057);
or UO_4564 (O_4564,N_47377,N_45726);
nand UO_4565 (O_4565,N_46422,N_49672);
or UO_4566 (O_4566,N_47522,N_47055);
and UO_4567 (O_4567,N_48206,N_46730);
nand UO_4568 (O_4568,N_49168,N_49566);
nor UO_4569 (O_4569,N_49475,N_45038);
or UO_4570 (O_4570,N_45154,N_45584);
nand UO_4571 (O_4571,N_49081,N_45176);
nor UO_4572 (O_4572,N_49211,N_46617);
nor UO_4573 (O_4573,N_49374,N_49204);
nor UO_4574 (O_4574,N_49517,N_46861);
nand UO_4575 (O_4575,N_45942,N_45238);
nand UO_4576 (O_4576,N_48611,N_46383);
xnor UO_4577 (O_4577,N_46574,N_45402);
nand UO_4578 (O_4578,N_46194,N_49394);
nand UO_4579 (O_4579,N_49601,N_45765);
or UO_4580 (O_4580,N_48752,N_49525);
or UO_4581 (O_4581,N_47818,N_49745);
or UO_4582 (O_4582,N_45762,N_48128);
nand UO_4583 (O_4583,N_49831,N_46445);
nand UO_4584 (O_4584,N_46750,N_45128);
or UO_4585 (O_4585,N_45079,N_48606);
and UO_4586 (O_4586,N_47565,N_49058);
nand UO_4587 (O_4587,N_45419,N_47503);
nor UO_4588 (O_4588,N_46657,N_48951);
nand UO_4589 (O_4589,N_47319,N_48782);
nand UO_4590 (O_4590,N_49481,N_48421);
nand UO_4591 (O_4591,N_46582,N_46663);
xnor UO_4592 (O_4592,N_49592,N_49469);
nor UO_4593 (O_4593,N_49132,N_48031);
nand UO_4594 (O_4594,N_49851,N_49780);
xnor UO_4595 (O_4595,N_47777,N_49183);
and UO_4596 (O_4596,N_45884,N_48098);
or UO_4597 (O_4597,N_48457,N_49187);
nor UO_4598 (O_4598,N_45014,N_48115);
nor UO_4599 (O_4599,N_48745,N_49666);
or UO_4600 (O_4600,N_48298,N_49541);
and UO_4601 (O_4601,N_47881,N_47949);
nand UO_4602 (O_4602,N_48216,N_48115);
nor UO_4603 (O_4603,N_49276,N_47916);
or UO_4604 (O_4604,N_46615,N_45824);
and UO_4605 (O_4605,N_49757,N_48940);
nor UO_4606 (O_4606,N_45049,N_49843);
and UO_4607 (O_4607,N_45957,N_47812);
nand UO_4608 (O_4608,N_45832,N_48061);
nand UO_4609 (O_4609,N_47254,N_48769);
and UO_4610 (O_4610,N_47846,N_46109);
or UO_4611 (O_4611,N_47813,N_46159);
nand UO_4612 (O_4612,N_47481,N_45295);
nor UO_4613 (O_4613,N_48699,N_47769);
nor UO_4614 (O_4614,N_48906,N_47284);
and UO_4615 (O_4615,N_47599,N_48811);
and UO_4616 (O_4616,N_49715,N_49157);
and UO_4617 (O_4617,N_48755,N_48057);
nor UO_4618 (O_4618,N_46408,N_47553);
nand UO_4619 (O_4619,N_49262,N_48296);
and UO_4620 (O_4620,N_48107,N_46428);
and UO_4621 (O_4621,N_48042,N_49223);
or UO_4622 (O_4622,N_48455,N_46606);
and UO_4623 (O_4623,N_49225,N_45905);
and UO_4624 (O_4624,N_47068,N_47918);
and UO_4625 (O_4625,N_46233,N_48805);
nor UO_4626 (O_4626,N_49259,N_45264);
or UO_4627 (O_4627,N_48323,N_49486);
or UO_4628 (O_4628,N_47703,N_47917);
nand UO_4629 (O_4629,N_49771,N_49147);
and UO_4630 (O_4630,N_48714,N_46036);
or UO_4631 (O_4631,N_46285,N_47676);
nand UO_4632 (O_4632,N_49820,N_46144);
xor UO_4633 (O_4633,N_45969,N_46038);
and UO_4634 (O_4634,N_45480,N_48287);
xor UO_4635 (O_4635,N_48514,N_47632);
nor UO_4636 (O_4636,N_48680,N_49972);
or UO_4637 (O_4637,N_46241,N_47848);
and UO_4638 (O_4638,N_45839,N_49934);
nor UO_4639 (O_4639,N_45938,N_45045);
or UO_4640 (O_4640,N_47044,N_46567);
or UO_4641 (O_4641,N_47899,N_45637);
nand UO_4642 (O_4642,N_45180,N_49035);
and UO_4643 (O_4643,N_47882,N_46404);
nor UO_4644 (O_4644,N_47415,N_47604);
and UO_4645 (O_4645,N_49300,N_48558);
or UO_4646 (O_4646,N_47704,N_46542);
xnor UO_4647 (O_4647,N_47201,N_49712);
nand UO_4648 (O_4648,N_45489,N_45201);
or UO_4649 (O_4649,N_47608,N_47611);
or UO_4650 (O_4650,N_47294,N_48798);
and UO_4651 (O_4651,N_45910,N_49379);
nor UO_4652 (O_4652,N_48518,N_47005);
and UO_4653 (O_4653,N_49031,N_49061);
or UO_4654 (O_4654,N_46949,N_48392);
and UO_4655 (O_4655,N_47503,N_45122);
xnor UO_4656 (O_4656,N_47592,N_49934);
and UO_4657 (O_4657,N_49516,N_45797);
nand UO_4658 (O_4658,N_48458,N_49708);
or UO_4659 (O_4659,N_48263,N_49673);
and UO_4660 (O_4660,N_49784,N_47773);
and UO_4661 (O_4661,N_49291,N_48472);
nand UO_4662 (O_4662,N_48684,N_46233);
nor UO_4663 (O_4663,N_49284,N_46490);
nor UO_4664 (O_4664,N_48899,N_47979);
nand UO_4665 (O_4665,N_47569,N_45683);
nand UO_4666 (O_4666,N_47544,N_47332);
nor UO_4667 (O_4667,N_46387,N_48198);
nand UO_4668 (O_4668,N_48554,N_48066);
or UO_4669 (O_4669,N_49364,N_47559);
or UO_4670 (O_4670,N_46422,N_46941);
nand UO_4671 (O_4671,N_49337,N_48164);
and UO_4672 (O_4672,N_48106,N_46876);
or UO_4673 (O_4673,N_48754,N_47152);
nor UO_4674 (O_4674,N_49387,N_49113);
and UO_4675 (O_4675,N_46704,N_45127);
and UO_4676 (O_4676,N_47273,N_47727);
and UO_4677 (O_4677,N_46079,N_46413);
nor UO_4678 (O_4678,N_46682,N_48583);
nand UO_4679 (O_4679,N_49943,N_49349);
and UO_4680 (O_4680,N_45743,N_46728);
nand UO_4681 (O_4681,N_49250,N_45755);
nand UO_4682 (O_4682,N_47443,N_48920);
nor UO_4683 (O_4683,N_48283,N_47477);
or UO_4684 (O_4684,N_45360,N_46521);
or UO_4685 (O_4685,N_47306,N_48922);
and UO_4686 (O_4686,N_48988,N_47870);
and UO_4687 (O_4687,N_49216,N_49294);
and UO_4688 (O_4688,N_49198,N_48412);
nor UO_4689 (O_4689,N_47280,N_48844);
nand UO_4690 (O_4690,N_49272,N_48446);
and UO_4691 (O_4691,N_45062,N_47712);
or UO_4692 (O_4692,N_48245,N_45524);
nand UO_4693 (O_4693,N_45982,N_47086);
nor UO_4694 (O_4694,N_47582,N_49760);
and UO_4695 (O_4695,N_48358,N_47655);
nor UO_4696 (O_4696,N_48123,N_47932);
nand UO_4697 (O_4697,N_48126,N_46833);
nand UO_4698 (O_4698,N_47531,N_45823);
nor UO_4699 (O_4699,N_45705,N_49520);
xnor UO_4700 (O_4700,N_48245,N_48953);
nor UO_4701 (O_4701,N_45827,N_46029);
and UO_4702 (O_4702,N_49507,N_47974);
nor UO_4703 (O_4703,N_49995,N_46070);
nor UO_4704 (O_4704,N_47189,N_48535);
and UO_4705 (O_4705,N_47596,N_46117);
nor UO_4706 (O_4706,N_47497,N_49481);
xnor UO_4707 (O_4707,N_48975,N_46729);
nor UO_4708 (O_4708,N_49894,N_49419);
or UO_4709 (O_4709,N_49152,N_47801);
nor UO_4710 (O_4710,N_45019,N_49416);
nor UO_4711 (O_4711,N_46003,N_49285);
and UO_4712 (O_4712,N_45433,N_49250);
and UO_4713 (O_4713,N_48900,N_45432);
nor UO_4714 (O_4714,N_47802,N_45015);
nand UO_4715 (O_4715,N_48387,N_45415);
nand UO_4716 (O_4716,N_46306,N_46137);
or UO_4717 (O_4717,N_46395,N_47844);
nand UO_4718 (O_4718,N_46726,N_48446);
or UO_4719 (O_4719,N_49729,N_46872);
xor UO_4720 (O_4720,N_49098,N_47377);
or UO_4721 (O_4721,N_45355,N_48702);
nor UO_4722 (O_4722,N_49592,N_45350);
xnor UO_4723 (O_4723,N_45808,N_48829);
or UO_4724 (O_4724,N_47522,N_47384);
and UO_4725 (O_4725,N_48389,N_48291);
and UO_4726 (O_4726,N_49950,N_49972);
nand UO_4727 (O_4727,N_47287,N_45346);
nor UO_4728 (O_4728,N_48790,N_48142);
and UO_4729 (O_4729,N_49629,N_49498);
and UO_4730 (O_4730,N_48711,N_47365);
and UO_4731 (O_4731,N_47535,N_46183);
or UO_4732 (O_4732,N_46027,N_48597);
nor UO_4733 (O_4733,N_49927,N_47006);
nand UO_4734 (O_4734,N_47022,N_46381);
and UO_4735 (O_4735,N_48084,N_47602);
and UO_4736 (O_4736,N_45756,N_48197);
xor UO_4737 (O_4737,N_48768,N_45851);
and UO_4738 (O_4738,N_46349,N_47531);
and UO_4739 (O_4739,N_47101,N_49396);
nand UO_4740 (O_4740,N_49514,N_46584);
and UO_4741 (O_4741,N_45374,N_49543);
nor UO_4742 (O_4742,N_48521,N_48660);
nor UO_4743 (O_4743,N_49879,N_48862);
nor UO_4744 (O_4744,N_48707,N_45436);
xor UO_4745 (O_4745,N_47373,N_49586);
nor UO_4746 (O_4746,N_48338,N_48278);
nor UO_4747 (O_4747,N_46075,N_48897);
or UO_4748 (O_4748,N_47861,N_49784);
nor UO_4749 (O_4749,N_46677,N_49522);
nor UO_4750 (O_4750,N_49313,N_49507);
or UO_4751 (O_4751,N_48531,N_46919);
and UO_4752 (O_4752,N_47489,N_45116);
and UO_4753 (O_4753,N_48649,N_46943);
nor UO_4754 (O_4754,N_48554,N_46350);
or UO_4755 (O_4755,N_45377,N_45648);
or UO_4756 (O_4756,N_48417,N_46585);
nand UO_4757 (O_4757,N_46751,N_47830);
or UO_4758 (O_4758,N_45612,N_45447);
and UO_4759 (O_4759,N_49333,N_45368);
nor UO_4760 (O_4760,N_47179,N_49583);
or UO_4761 (O_4761,N_48495,N_48582);
or UO_4762 (O_4762,N_49133,N_48750);
and UO_4763 (O_4763,N_45180,N_48773);
xor UO_4764 (O_4764,N_46713,N_47561);
nand UO_4765 (O_4765,N_45293,N_49038);
nor UO_4766 (O_4766,N_49898,N_46028);
and UO_4767 (O_4767,N_46841,N_47898);
and UO_4768 (O_4768,N_48955,N_49606);
xnor UO_4769 (O_4769,N_45531,N_46861);
nand UO_4770 (O_4770,N_45770,N_47730);
nor UO_4771 (O_4771,N_49849,N_46675);
nor UO_4772 (O_4772,N_49779,N_46477);
or UO_4773 (O_4773,N_49505,N_47432);
xor UO_4774 (O_4774,N_47117,N_46637);
or UO_4775 (O_4775,N_49528,N_46080);
and UO_4776 (O_4776,N_47951,N_49161);
nand UO_4777 (O_4777,N_46311,N_46956);
or UO_4778 (O_4778,N_46641,N_47076);
or UO_4779 (O_4779,N_46669,N_45725);
nand UO_4780 (O_4780,N_45423,N_45078);
and UO_4781 (O_4781,N_47045,N_45466);
nor UO_4782 (O_4782,N_45299,N_49754);
or UO_4783 (O_4783,N_47730,N_45160);
and UO_4784 (O_4784,N_49694,N_46699);
nand UO_4785 (O_4785,N_49243,N_46817);
nor UO_4786 (O_4786,N_45785,N_49250);
and UO_4787 (O_4787,N_46909,N_49748);
nand UO_4788 (O_4788,N_46364,N_48604);
or UO_4789 (O_4789,N_45252,N_48754);
nand UO_4790 (O_4790,N_49155,N_45567);
and UO_4791 (O_4791,N_45020,N_47947);
nor UO_4792 (O_4792,N_49916,N_49576);
nor UO_4793 (O_4793,N_45278,N_48517);
nand UO_4794 (O_4794,N_46428,N_49173);
and UO_4795 (O_4795,N_48333,N_45007);
and UO_4796 (O_4796,N_45849,N_45715);
nand UO_4797 (O_4797,N_46273,N_49252);
nand UO_4798 (O_4798,N_49510,N_48843);
nand UO_4799 (O_4799,N_48839,N_45547);
and UO_4800 (O_4800,N_48282,N_49871);
and UO_4801 (O_4801,N_48866,N_46076);
nand UO_4802 (O_4802,N_49210,N_48827);
nand UO_4803 (O_4803,N_45534,N_46318);
and UO_4804 (O_4804,N_48130,N_47702);
nand UO_4805 (O_4805,N_47371,N_49520);
nor UO_4806 (O_4806,N_45121,N_46135);
or UO_4807 (O_4807,N_48433,N_45234);
nand UO_4808 (O_4808,N_45525,N_47006);
or UO_4809 (O_4809,N_49966,N_49822);
or UO_4810 (O_4810,N_45914,N_49145);
nand UO_4811 (O_4811,N_46180,N_45783);
nor UO_4812 (O_4812,N_49766,N_49689);
or UO_4813 (O_4813,N_46284,N_47953);
xnor UO_4814 (O_4814,N_48363,N_49843);
xnor UO_4815 (O_4815,N_46118,N_45782);
nor UO_4816 (O_4816,N_48151,N_49026);
nand UO_4817 (O_4817,N_46944,N_45442);
nand UO_4818 (O_4818,N_47305,N_45274);
nor UO_4819 (O_4819,N_49362,N_45473);
xnor UO_4820 (O_4820,N_47285,N_49806);
xnor UO_4821 (O_4821,N_46816,N_46055);
nand UO_4822 (O_4822,N_46380,N_47337);
xor UO_4823 (O_4823,N_46463,N_46077);
nor UO_4824 (O_4824,N_45628,N_45206);
nand UO_4825 (O_4825,N_46855,N_49861);
and UO_4826 (O_4826,N_45420,N_46309);
and UO_4827 (O_4827,N_46426,N_48171);
nand UO_4828 (O_4828,N_45622,N_49259);
or UO_4829 (O_4829,N_47485,N_46040);
nand UO_4830 (O_4830,N_47983,N_47109);
and UO_4831 (O_4831,N_45890,N_45458);
and UO_4832 (O_4832,N_46580,N_45196);
nand UO_4833 (O_4833,N_48980,N_48841);
xnor UO_4834 (O_4834,N_48973,N_49019);
and UO_4835 (O_4835,N_47447,N_45987);
or UO_4836 (O_4836,N_45312,N_47419);
or UO_4837 (O_4837,N_47385,N_46737);
xnor UO_4838 (O_4838,N_45563,N_46445);
nand UO_4839 (O_4839,N_45696,N_45978);
and UO_4840 (O_4840,N_47428,N_47301);
nor UO_4841 (O_4841,N_49549,N_47080);
nand UO_4842 (O_4842,N_45046,N_46603);
and UO_4843 (O_4843,N_47538,N_49712);
or UO_4844 (O_4844,N_46637,N_49060);
and UO_4845 (O_4845,N_47815,N_45458);
and UO_4846 (O_4846,N_48018,N_46588);
nand UO_4847 (O_4847,N_47390,N_47965);
nor UO_4848 (O_4848,N_45413,N_47583);
nor UO_4849 (O_4849,N_46304,N_48051);
and UO_4850 (O_4850,N_47140,N_45875);
nand UO_4851 (O_4851,N_46051,N_46785);
nand UO_4852 (O_4852,N_48851,N_46359);
nor UO_4853 (O_4853,N_47446,N_45670);
and UO_4854 (O_4854,N_45427,N_46026);
nand UO_4855 (O_4855,N_45284,N_45651);
nand UO_4856 (O_4856,N_47993,N_45020);
nand UO_4857 (O_4857,N_47369,N_47777);
and UO_4858 (O_4858,N_49410,N_46249);
nand UO_4859 (O_4859,N_49171,N_46840);
nor UO_4860 (O_4860,N_45303,N_46515);
nand UO_4861 (O_4861,N_47575,N_47123);
xnor UO_4862 (O_4862,N_46900,N_49919);
nand UO_4863 (O_4863,N_47951,N_49207);
nor UO_4864 (O_4864,N_49426,N_48284);
and UO_4865 (O_4865,N_49474,N_47980);
nor UO_4866 (O_4866,N_49114,N_48890);
and UO_4867 (O_4867,N_46081,N_49689);
and UO_4868 (O_4868,N_45457,N_46549);
or UO_4869 (O_4869,N_49990,N_45103);
or UO_4870 (O_4870,N_45678,N_48424);
or UO_4871 (O_4871,N_45504,N_47495);
nand UO_4872 (O_4872,N_49355,N_46736);
nor UO_4873 (O_4873,N_49534,N_49465);
and UO_4874 (O_4874,N_49543,N_48760);
or UO_4875 (O_4875,N_46301,N_47202);
and UO_4876 (O_4876,N_49203,N_47429);
or UO_4877 (O_4877,N_48312,N_45618);
and UO_4878 (O_4878,N_47826,N_47677);
and UO_4879 (O_4879,N_47585,N_45689);
and UO_4880 (O_4880,N_46243,N_49994);
nand UO_4881 (O_4881,N_47477,N_49678);
xor UO_4882 (O_4882,N_46769,N_46122);
or UO_4883 (O_4883,N_45484,N_47287);
nor UO_4884 (O_4884,N_49143,N_47471);
nor UO_4885 (O_4885,N_47299,N_49816);
nand UO_4886 (O_4886,N_45229,N_49098);
xor UO_4887 (O_4887,N_46598,N_46146);
nand UO_4888 (O_4888,N_49904,N_45241);
and UO_4889 (O_4889,N_47273,N_48878);
or UO_4890 (O_4890,N_45274,N_47976);
nor UO_4891 (O_4891,N_49716,N_46628);
nand UO_4892 (O_4892,N_47766,N_48078);
nand UO_4893 (O_4893,N_46414,N_47010);
nand UO_4894 (O_4894,N_49129,N_46448);
nand UO_4895 (O_4895,N_47724,N_49903);
and UO_4896 (O_4896,N_46671,N_49936);
or UO_4897 (O_4897,N_46141,N_49504);
xnor UO_4898 (O_4898,N_46415,N_47356);
nor UO_4899 (O_4899,N_47338,N_48840);
nand UO_4900 (O_4900,N_49203,N_46308);
and UO_4901 (O_4901,N_48722,N_47447);
nand UO_4902 (O_4902,N_47589,N_46929);
nand UO_4903 (O_4903,N_46481,N_47326);
nor UO_4904 (O_4904,N_46311,N_48606);
and UO_4905 (O_4905,N_49882,N_48952);
and UO_4906 (O_4906,N_46570,N_46683);
and UO_4907 (O_4907,N_49071,N_47840);
xor UO_4908 (O_4908,N_48304,N_45224);
and UO_4909 (O_4909,N_45693,N_45616);
xnor UO_4910 (O_4910,N_45646,N_47750);
or UO_4911 (O_4911,N_47037,N_47927);
and UO_4912 (O_4912,N_49118,N_49840);
or UO_4913 (O_4913,N_45172,N_49076);
nand UO_4914 (O_4914,N_45481,N_48928);
nand UO_4915 (O_4915,N_46194,N_46773);
nand UO_4916 (O_4916,N_46518,N_49860);
nand UO_4917 (O_4917,N_48965,N_49354);
nor UO_4918 (O_4918,N_48258,N_49439);
nand UO_4919 (O_4919,N_48937,N_46345);
or UO_4920 (O_4920,N_49737,N_47703);
and UO_4921 (O_4921,N_48128,N_47046);
and UO_4922 (O_4922,N_48904,N_47326);
nor UO_4923 (O_4923,N_49869,N_49479);
nor UO_4924 (O_4924,N_46328,N_47291);
nand UO_4925 (O_4925,N_47785,N_46608);
nand UO_4926 (O_4926,N_45912,N_49328);
or UO_4927 (O_4927,N_47022,N_45183);
nor UO_4928 (O_4928,N_46204,N_46780);
and UO_4929 (O_4929,N_47445,N_45702);
nand UO_4930 (O_4930,N_46935,N_47838);
or UO_4931 (O_4931,N_48022,N_45344);
and UO_4932 (O_4932,N_47151,N_45104);
and UO_4933 (O_4933,N_45440,N_47338);
nor UO_4934 (O_4934,N_48137,N_48575);
nand UO_4935 (O_4935,N_49319,N_48834);
or UO_4936 (O_4936,N_45859,N_49166);
or UO_4937 (O_4937,N_48053,N_49805);
or UO_4938 (O_4938,N_48361,N_46272);
and UO_4939 (O_4939,N_46687,N_45162);
and UO_4940 (O_4940,N_48666,N_45400);
nor UO_4941 (O_4941,N_46743,N_48669);
or UO_4942 (O_4942,N_47021,N_47337);
nand UO_4943 (O_4943,N_49505,N_49967);
nor UO_4944 (O_4944,N_48544,N_48229);
nand UO_4945 (O_4945,N_47375,N_49749);
or UO_4946 (O_4946,N_46315,N_46189);
xnor UO_4947 (O_4947,N_47242,N_47073);
nand UO_4948 (O_4948,N_47840,N_46137);
nor UO_4949 (O_4949,N_48649,N_46211);
or UO_4950 (O_4950,N_48987,N_45499);
nor UO_4951 (O_4951,N_48600,N_48781);
or UO_4952 (O_4952,N_47703,N_46092);
and UO_4953 (O_4953,N_48812,N_49366);
nand UO_4954 (O_4954,N_49565,N_46898);
nor UO_4955 (O_4955,N_47274,N_48476);
or UO_4956 (O_4956,N_47230,N_48101);
xor UO_4957 (O_4957,N_45441,N_46629);
or UO_4958 (O_4958,N_49007,N_49901);
nor UO_4959 (O_4959,N_48072,N_45303);
or UO_4960 (O_4960,N_45139,N_49775);
nor UO_4961 (O_4961,N_46310,N_45948);
or UO_4962 (O_4962,N_46387,N_49493);
nand UO_4963 (O_4963,N_48393,N_49934);
nor UO_4964 (O_4964,N_45496,N_45465);
nor UO_4965 (O_4965,N_47781,N_47049);
and UO_4966 (O_4966,N_45495,N_49383);
nor UO_4967 (O_4967,N_47170,N_46668);
nor UO_4968 (O_4968,N_46391,N_45933);
or UO_4969 (O_4969,N_48629,N_49616);
or UO_4970 (O_4970,N_48824,N_47639);
nand UO_4971 (O_4971,N_48190,N_45399);
nor UO_4972 (O_4972,N_47874,N_47208);
and UO_4973 (O_4973,N_48508,N_45260);
nor UO_4974 (O_4974,N_49968,N_46513);
and UO_4975 (O_4975,N_45357,N_49323);
nor UO_4976 (O_4976,N_45624,N_46601);
nand UO_4977 (O_4977,N_49361,N_49418);
nor UO_4978 (O_4978,N_45917,N_45966);
or UO_4979 (O_4979,N_46713,N_47397);
or UO_4980 (O_4980,N_46236,N_48885);
or UO_4981 (O_4981,N_46578,N_49705);
nor UO_4982 (O_4982,N_48781,N_47199);
nand UO_4983 (O_4983,N_45989,N_47968);
and UO_4984 (O_4984,N_48376,N_48034);
nor UO_4985 (O_4985,N_48623,N_47680);
nor UO_4986 (O_4986,N_48905,N_47035);
and UO_4987 (O_4987,N_49013,N_46798);
nor UO_4988 (O_4988,N_49051,N_46271);
or UO_4989 (O_4989,N_48134,N_45749);
or UO_4990 (O_4990,N_49557,N_49169);
or UO_4991 (O_4991,N_48037,N_49637);
and UO_4992 (O_4992,N_46709,N_47735);
and UO_4993 (O_4993,N_45325,N_46260);
nand UO_4994 (O_4994,N_45943,N_45685);
nor UO_4995 (O_4995,N_48269,N_46407);
and UO_4996 (O_4996,N_48661,N_47283);
and UO_4997 (O_4997,N_49721,N_49458);
nand UO_4998 (O_4998,N_48379,N_45671);
nor UO_4999 (O_4999,N_47019,N_45117);
endmodule