module basic_500_3000_500_30_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_260,In_368);
or U1 (N_1,In_402,In_9);
or U2 (N_2,In_297,In_41);
nand U3 (N_3,In_334,In_296);
and U4 (N_4,In_97,In_219);
and U5 (N_5,In_477,In_206);
nand U6 (N_6,In_32,In_484);
nor U7 (N_7,In_249,In_110);
nand U8 (N_8,In_475,In_486);
nor U9 (N_9,In_418,In_374);
and U10 (N_10,In_258,In_191);
nand U11 (N_11,In_422,In_287);
and U12 (N_12,In_198,In_90);
or U13 (N_13,In_330,In_454);
nand U14 (N_14,In_417,In_464);
and U15 (N_15,In_423,In_226);
or U16 (N_16,In_107,In_393);
nor U17 (N_17,In_326,In_58);
or U18 (N_18,In_201,In_295);
and U19 (N_19,In_491,In_432);
and U20 (N_20,In_92,In_139);
nor U21 (N_21,In_203,In_461);
and U22 (N_22,In_310,In_37);
nor U23 (N_23,In_140,In_291);
or U24 (N_24,In_98,In_100);
nand U25 (N_25,In_298,In_439);
and U26 (N_26,In_50,In_425);
nor U27 (N_27,In_487,In_19);
nand U28 (N_28,In_150,In_343);
and U29 (N_29,In_300,In_273);
and U30 (N_30,In_324,In_220);
nor U31 (N_31,In_337,In_333);
or U32 (N_32,In_102,In_153);
nor U33 (N_33,In_174,In_444);
or U34 (N_34,In_363,In_332);
nor U35 (N_35,In_14,In_134);
or U36 (N_36,In_69,In_453);
or U37 (N_37,In_240,In_474);
nor U38 (N_38,In_128,In_395);
nor U39 (N_39,In_307,In_212);
and U40 (N_40,In_391,In_105);
or U41 (N_41,In_106,In_168);
nand U42 (N_42,In_305,In_170);
nor U43 (N_43,In_381,In_5);
and U44 (N_44,In_25,In_377);
nor U45 (N_45,In_103,In_489);
nor U46 (N_46,In_4,In_1);
nor U47 (N_47,In_427,In_158);
nor U48 (N_48,In_421,In_341);
or U49 (N_49,In_118,In_59);
nor U50 (N_50,In_53,In_0);
and U51 (N_51,In_472,In_160);
nor U52 (N_52,In_397,In_48);
nor U53 (N_53,In_179,In_87);
and U54 (N_54,In_216,In_451);
or U55 (N_55,In_325,In_496);
and U56 (N_56,In_483,In_346);
or U57 (N_57,In_161,In_457);
and U58 (N_58,In_121,In_141);
or U59 (N_59,In_351,In_406);
or U60 (N_60,In_135,In_403);
nand U61 (N_61,In_31,In_211);
nor U62 (N_62,In_30,In_469);
nor U63 (N_63,In_71,In_154);
or U64 (N_64,In_450,In_312);
or U65 (N_65,In_88,In_43);
nand U66 (N_66,In_83,In_336);
and U67 (N_67,In_183,In_431);
and U68 (N_68,In_367,In_455);
nand U69 (N_69,In_15,In_338);
nand U70 (N_70,In_282,In_271);
and U71 (N_71,In_224,In_490);
nand U72 (N_72,In_319,In_120);
and U73 (N_73,In_364,In_241);
or U74 (N_74,In_236,In_6);
and U75 (N_75,In_429,In_152);
nor U76 (N_76,In_399,In_452);
and U77 (N_77,In_144,In_498);
nand U78 (N_78,In_189,In_348);
and U79 (N_79,In_199,In_447);
and U80 (N_80,In_167,In_331);
and U81 (N_81,In_221,In_178);
nand U82 (N_82,In_380,In_479);
or U83 (N_83,In_250,In_45);
or U84 (N_84,In_210,In_392);
nand U85 (N_85,In_163,In_378);
xor U86 (N_86,In_232,In_294);
nand U87 (N_87,In_394,In_443);
and U88 (N_88,In_123,In_438);
nand U89 (N_89,In_497,In_99);
and U90 (N_90,In_230,In_366);
and U91 (N_91,In_116,In_54);
and U92 (N_92,In_360,In_376);
nand U93 (N_93,In_459,In_27);
nand U94 (N_94,In_34,In_449);
nor U95 (N_95,In_57,In_290);
and U96 (N_96,In_318,In_493);
nor U97 (N_97,In_205,In_492);
nor U98 (N_98,In_130,In_186);
and U99 (N_99,In_75,In_372);
and U100 (N_100,In_478,In_96);
and U101 (N_101,In_315,In_227);
nand U102 (N_102,In_164,N_2);
or U103 (N_103,In_414,In_286);
and U104 (N_104,In_237,In_355);
and U105 (N_105,N_27,In_238);
and U106 (N_106,In_488,In_404);
or U107 (N_107,In_95,In_146);
and U108 (N_108,In_137,In_2);
nand U109 (N_109,In_47,In_76);
nand U110 (N_110,In_33,In_101);
and U111 (N_111,N_51,In_149);
nor U112 (N_112,N_7,In_356);
or U113 (N_113,In_384,In_229);
nand U114 (N_114,In_410,In_359);
or U115 (N_115,In_151,In_280);
or U116 (N_116,In_223,In_18);
nand U117 (N_117,In_354,N_77);
nand U118 (N_118,In_214,In_306);
nor U119 (N_119,N_36,In_382);
nand U120 (N_120,In_188,In_39);
or U121 (N_121,N_9,In_292);
nand U122 (N_122,In_499,In_344);
and U123 (N_123,In_166,In_316);
xnor U124 (N_124,In_284,In_481);
nand U125 (N_125,N_13,In_379);
and U126 (N_126,N_23,In_52);
nand U127 (N_127,In_259,In_430);
and U128 (N_128,In_10,In_86);
xnor U129 (N_129,N_12,In_63);
nor U130 (N_130,In_353,In_339);
nor U131 (N_131,In_79,N_60);
xnor U132 (N_132,In_187,In_435);
or U133 (N_133,In_28,In_108);
nor U134 (N_134,In_147,In_126);
or U135 (N_135,In_114,In_327);
nor U136 (N_136,In_24,In_207);
or U137 (N_137,In_46,N_49);
nor U138 (N_138,N_44,In_218);
nand U139 (N_139,In_131,In_244);
or U140 (N_140,In_78,In_442);
or U141 (N_141,In_361,N_91);
and U142 (N_142,In_350,In_60);
nand U143 (N_143,In_66,In_390);
nand U144 (N_144,In_279,In_313);
nor U145 (N_145,In_234,In_177);
or U146 (N_146,In_62,N_68);
or U147 (N_147,In_433,In_458);
or U148 (N_148,In_460,In_272);
or U149 (N_149,N_73,In_373);
and U150 (N_150,N_74,In_270);
nand U151 (N_151,In_387,In_20);
nor U152 (N_152,In_358,In_70);
or U153 (N_153,In_266,In_371);
nand U154 (N_154,N_50,In_12);
nand U155 (N_155,In_252,In_405);
or U156 (N_156,In_246,N_54);
or U157 (N_157,In_415,N_11);
nand U158 (N_158,In_85,In_445);
or U159 (N_159,In_276,N_5);
nand U160 (N_160,In_217,In_196);
or U161 (N_161,In_243,N_81);
or U162 (N_162,In_49,In_193);
nor U163 (N_163,In_148,In_145);
nand U164 (N_164,In_328,In_302);
nand U165 (N_165,N_14,N_16);
or U166 (N_166,In_357,In_200);
nor U167 (N_167,N_55,In_420);
and U168 (N_168,N_41,In_225);
or U169 (N_169,In_35,In_335);
nand U170 (N_170,In_94,In_262);
and U171 (N_171,In_485,In_281);
and U172 (N_172,In_265,N_65);
nor U173 (N_173,N_76,N_29);
and U174 (N_174,In_285,N_15);
nand U175 (N_175,In_180,In_93);
and U176 (N_176,In_400,In_195);
nand U177 (N_177,In_209,N_53);
or U178 (N_178,N_86,In_77);
and U179 (N_179,In_197,In_303);
or U180 (N_180,In_16,In_329);
or U181 (N_181,N_69,N_80);
and U182 (N_182,In_267,In_182);
or U183 (N_183,In_288,In_320);
nand U184 (N_184,In_428,In_213);
and U185 (N_185,In_143,In_263);
or U186 (N_186,In_342,In_375);
or U187 (N_187,In_426,N_84);
or U188 (N_188,In_89,N_99);
nor U189 (N_189,In_67,In_22);
and U190 (N_190,N_85,N_47);
xor U191 (N_191,N_90,N_57);
or U192 (N_192,In_301,In_122);
nand U193 (N_193,N_20,In_293);
or U194 (N_194,In_44,N_43);
or U195 (N_195,N_78,In_463);
nand U196 (N_196,In_247,In_13);
and U197 (N_197,N_42,In_471);
or U198 (N_198,In_446,N_26);
or U199 (N_199,N_1,In_456);
nor U200 (N_200,N_169,N_189);
nand U201 (N_201,In_314,In_132);
nand U202 (N_202,N_95,In_419);
or U203 (N_203,In_157,N_70);
nor U204 (N_204,N_157,In_261);
nor U205 (N_205,N_132,In_115);
or U206 (N_206,N_195,N_79);
or U207 (N_207,In_466,In_185);
or U208 (N_208,In_278,N_104);
or U209 (N_209,In_119,In_127);
or U210 (N_210,In_388,N_185);
or U211 (N_211,N_3,In_416);
or U212 (N_212,N_172,N_66);
nand U213 (N_213,In_190,N_147);
nor U214 (N_214,N_107,N_154);
or U215 (N_215,N_196,N_178);
and U216 (N_216,N_146,N_133);
nor U217 (N_217,In_72,In_65);
and U218 (N_218,In_253,N_30);
nor U219 (N_219,In_80,N_100);
nand U220 (N_220,N_163,N_75);
and U221 (N_221,N_59,N_125);
or U222 (N_222,In_169,In_42);
or U223 (N_223,In_245,In_248);
and U224 (N_224,In_277,N_38);
nand U225 (N_225,N_149,N_24);
and U226 (N_226,N_130,In_215);
and U227 (N_227,In_228,N_32);
or U228 (N_228,N_4,In_36);
nor U229 (N_229,In_274,In_321);
nand U230 (N_230,In_311,N_93);
nor U231 (N_231,In_268,In_142);
nand U232 (N_232,N_48,In_437);
nor U233 (N_233,N_22,In_124);
and U234 (N_234,In_441,N_88);
and U235 (N_235,N_39,In_204);
or U236 (N_236,In_370,In_476);
nor U237 (N_237,N_102,N_67);
nand U238 (N_238,In_411,In_138);
and U239 (N_239,In_465,In_64);
and U240 (N_240,N_158,N_153);
and U241 (N_241,In_283,N_89);
nor U242 (N_242,In_264,In_40);
or U243 (N_243,In_494,N_109);
nand U244 (N_244,N_46,N_199);
or U245 (N_245,N_171,N_96);
or U246 (N_246,In_7,N_33);
nor U247 (N_247,In_173,In_184);
nor U248 (N_248,N_31,N_160);
or U249 (N_249,In_467,In_73);
nand U250 (N_250,N_113,In_255);
or U251 (N_251,In_408,In_176);
or U252 (N_252,In_117,N_111);
and U253 (N_253,In_317,N_143);
and U254 (N_254,In_68,N_167);
nor U255 (N_255,N_181,In_308);
nand U256 (N_256,N_148,N_123);
or U257 (N_257,N_0,N_128);
or U258 (N_258,In_257,In_91);
nand U259 (N_259,In_55,In_175);
nand U260 (N_260,In_424,N_162);
and U261 (N_261,N_144,N_71);
and U262 (N_262,N_142,N_135);
nand U263 (N_263,In_256,N_186);
or U264 (N_264,N_176,N_175);
or U265 (N_265,In_275,In_362);
nor U266 (N_266,In_462,In_113);
nor U267 (N_267,In_309,In_129);
nand U268 (N_268,In_136,In_347);
nor U269 (N_269,N_62,N_87);
nand U270 (N_270,N_105,N_97);
and U271 (N_271,In_412,In_17);
or U272 (N_272,In_26,N_197);
nand U273 (N_273,N_139,In_133);
nand U274 (N_274,N_131,In_396);
or U275 (N_275,In_409,N_98);
nand U276 (N_276,In_51,In_233);
or U277 (N_277,In_125,N_191);
or U278 (N_278,N_117,In_345);
nand U279 (N_279,N_37,In_192);
nor U280 (N_280,N_198,N_179);
nor U281 (N_281,N_25,N_168);
and U282 (N_282,N_166,In_208);
and U283 (N_283,N_159,N_155);
nor U284 (N_284,In_470,N_19);
nor U285 (N_285,N_116,In_3);
nor U286 (N_286,N_56,N_40);
or U287 (N_287,N_126,N_183);
nand U288 (N_288,N_34,N_45);
nand U289 (N_289,N_108,In_239);
nor U290 (N_290,N_61,In_81);
and U291 (N_291,N_192,N_184);
nand U292 (N_292,In_74,N_180);
nor U293 (N_293,N_138,In_473);
or U294 (N_294,In_242,In_352);
and U295 (N_295,In_8,N_120);
and U296 (N_296,N_145,In_159);
or U297 (N_297,In_155,In_202);
or U298 (N_298,In_269,N_118);
and U299 (N_299,N_165,N_17);
or U300 (N_300,N_92,In_11);
and U301 (N_301,N_234,N_101);
nand U302 (N_302,In_111,N_262);
nor U303 (N_303,N_263,N_218);
nand U304 (N_304,N_151,In_84);
nor U305 (N_305,N_205,N_211);
and U306 (N_306,N_201,N_203);
and U307 (N_307,N_229,N_28);
nor U308 (N_308,N_240,In_289);
nand U309 (N_309,N_182,In_61);
nor U310 (N_310,N_119,N_82);
or U311 (N_311,N_278,N_279);
nor U312 (N_312,N_209,N_283);
and U313 (N_313,N_190,N_288);
nand U314 (N_314,In_251,N_194);
and U315 (N_315,In_38,In_56);
and U316 (N_316,N_295,N_63);
or U317 (N_317,N_140,In_171);
nor U318 (N_318,N_276,N_266);
and U319 (N_319,N_231,N_248);
nor U320 (N_320,N_251,In_440);
nand U321 (N_321,N_246,N_204);
xor U322 (N_322,In_401,N_290);
or U323 (N_323,N_294,N_232);
and U324 (N_324,N_259,N_241);
nand U325 (N_325,In_436,In_480);
nor U326 (N_326,N_21,N_292);
nand U327 (N_327,In_162,In_389);
nor U328 (N_328,In_448,N_280);
or U329 (N_329,N_272,N_223);
and U330 (N_330,N_110,In_165);
and U331 (N_331,N_112,N_156);
nor U332 (N_332,N_267,N_237);
and U333 (N_333,In_109,N_253);
or U334 (N_334,N_216,N_296);
and U335 (N_335,In_365,N_215);
nor U336 (N_336,In_235,N_122);
nand U337 (N_337,N_270,N_299);
or U338 (N_338,N_208,N_212);
or U339 (N_339,N_271,N_224);
or U340 (N_340,In_222,N_177);
nor U341 (N_341,N_291,N_258);
nand U342 (N_342,N_35,N_217);
and U343 (N_343,N_6,N_282);
nand U344 (N_344,N_273,In_468);
nor U345 (N_345,N_83,N_121);
and U346 (N_346,In_340,N_161);
nand U347 (N_347,In_21,N_150);
or U348 (N_348,N_239,In_112);
and U349 (N_349,N_114,N_227);
nand U350 (N_350,N_298,N_286);
nand U351 (N_351,N_225,N_213);
nor U352 (N_352,N_141,N_228);
and U353 (N_353,N_136,N_285);
nor U354 (N_354,N_72,N_103);
and U355 (N_355,In_322,N_137);
and U356 (N_356,In_434,N_220);
and U357 (N_357,N_233,N_252);
nor U358 (N_358,N_235,N_265);
nand U359 (N_359,N_250,N_275);
nor U360 (N_360,N_254,N_256);
and U361 (N_361,N_260,N_174);
nand U362 (N_362,N_202,In_304);
and U363 (N_363,In_194,N_257);
nand U364 (N_364,In_172,N_10);
nor U365 (N_365,N_249,N_238);
nand U366 (N_366,In_23,N_222);
or U367 (N_367,N_247,N_124);
nand U368 (N_368,N_274,N_268);
nand U369 (N_369,N_214,N_261);
and U370 (N_370,In_413,N_244);
and U371 (N_371,In_383,In_385);
or U372 (N_372,N_206,In_369);
xnor U373 (N_373,N_129,N_230);
nand U374 (N_374,In_323,N_269);
nand U375 (N_375,N_187,In_82);
nor U376 (N_376,N_134,N_221);
or U377 (N_377,N_200,N_58);
nand U378 (N_378,In_299,N_293);
nor U379 (N_379,N_173,N_170);
nand U380 (N_380,N_188,N_193);
nand U381 (N_381,N_152,N_255);
nor U382 (N_382,N_289,In_156);
nand U383 (N_383,In_398,In_29);
xor U384 (N_384,N_264,N_8);
nor U385 (N_385,N_94,In_104);
nor U386 (N_386,N_207,N_245);
nor U387 (N_387,In_254,N_115);
nor U388 (N_388,N_64,N_297);
nor U389 (N_389,N_106,N_287);
nand U390 (N_390,In_407,N_277);
nor U391 (N_391,N_219,In_495);
and U392 (N_392,In_482,N_210);
and U393 (N_393,N_284,N_164);
or U394 (N_394,In_181,N_226);
nand U395 (N_395,In_231,In_386);
nand U396 (N_396,N_242,N_52);
nand U397 (N_397,N_127,N_281);
and U398 (N_398,N_18,N_236);
nor U399 (N_399,In_349,N_243);
nand U400 (N_400,N_330,N_346);
nand U401 (N_401,N_314,N_385);
or U402 (N_402,N_381,N_394);
or U403 (N_403,N_341,N_317);
or U404 (N_404,N_366,N_310);
and U405 (N_405,N_359,N_320);
or U406 (N_406,N_342,N_362);
or U407 (N_407,N_304,N_311);
nand U408 (N_408,N_328,N_389);
nor U409 (N_409,N_395,N_355);
nand U410 (N_410,N_367,N_344);
nor U411 (N_411,N_368,N_354);
or U412 (N_412,N_343,N_369);
nor U413 (N_413,N_332,N_315);
and U414 (N_414,N_336,N_326);
or U415 (N_415,N_388,N_397);
and U416 (N_416,N_374,N_383);
nor U417 (N_417,N_338,N_387);
nand U418 (N_418,N_324,N_305);
or U419 (N_419,N_363,N_357);
and U420 (N_420,N_337,N_301);
or U421 (N_421,N_360,N_375);
or U422 (N_422,N_365,N_396);
nand U423 (N_423,N_384,N_303);
nand U424 (N_424,N_370,N_345);
or U425 (N_425,N_372,N_316);
nor U426 (N_426,N_358,N_349);
nand U427 (N_427,N_340,N_390);
and U428 (N_428,N_334,N_373);
nor U429 (N_429,N_352,N_356);
or U430 (N_430,N_319,N_302);
nand U431 (N_431,N_307,N_308);
or U432 (N_432,N_347,N_393);
nor U433 (N_433,N_378,N_306);
nand U434 (N_434,N_379,N_392);
or U435 (N_435,N_376,N_377);
and U436 (N_436,N_331,N_309);
nor U437 (N_437,N_361,N_313);
nand U438 (N_438,N_323,N_386);
or U439 (N_439,N_348,N_353);
and U440 (N_440,N_399,N_321);
or U441 (N_441,N_364,N_322);
and U442 (N_442,N_300,N_329);
or U443 (N_443,N_351,N_380);
nor U444 (N_444,N_339,N_391);
nor U445 (N_445,N_318,N_335);
or U446 (N_446,N_312,N_327);
nand U447 (N_447,N_350,N_325);
nor U448 (N_448,N_333,N_398);
nor U449 (N_449,N_371,N_382);
and U450 (N_450,N_352,N_319);
and U451 (N_451,N_361,N_381);
or U452 (N_452,N_304,N_302);
and U453 (N_453,N_386,N_381);
nor U454 (N_454,N_334,N_367);
nand U455 (N_455,N_375,N_390);
or U456 (N_456,N_314,N_331);
nor U457 (N_457,N_375,N_331);
nor U458 (N_458,N_371,N_385);
nor U459 (N_459,N_386,N_358);
nor U460 (N_460,N_365,N_307);
or U461 (N_461,N_384,N_314);
or U462 (N_462,N_336,N_349);
nand U463 (N_463,N_351,N_394);
and U464 (N_464,N_305,N_365);
xor U465 (N_465,N_338,N_362);
nand U466 (N_466,N_366,N_368);
and U467 (N_467,N_388,N_392);
and U468 (N_468,N_313,N_393);
and U469 (N_469,N_359,N_300);
nand U470 (N_470,N_358,N_327);
and U471 (N_471,N_354,N_343);
nand U472 (N_472,N_348,N_314);
nand U473 (N_473,N_346,N_339);
nand U474 (N_474,N_392,N_313);
nand U475 (N_475,N_346,N_362);
or U476 (N_476,N_336,N_322);
nand U477 (N_477,N_384,N_301);
xnor U478 (N_478,N_388,N_382);
and U479 (N_479,N_385,N_328);
nand U480 (N_480,N_351,N_323);
and U481 (N_481,N_341,N_304);
nand U482 (N_482,N_374,N_399);
nand U483 (N_483,N_372,N_354);
or U484 (N_484,N_342,N_337);
nand U485 (N_485,N_326,N_303);
nor U486 (N_486,N_333,N_337);
and U487 (N_487,N_383,N_373);
nor U488 (N_488,N_350,N_340);
and U489 (N_489,N_337,N_322);
or U490 (N_490,N_368,N_391);
or U491 (N_491,N_357,N_334);
or U492 (N_492,N_345,N_356);
and U493 (N_493,N_350,N_392);
or U494 (N_494,N_351,N_347);
nand U495 (N_495,N_307,N_324);
nor U496 (N_496,N_378,N_345);
or U497 (N_497,N_347,N_370);
and U498 (N_498,N_355,N_349);
nand U499 (N_499,N_313,N_307);
nor U500 (N_500,N_439,N_457);
or U501 (N_501,N_433,N_489);
nand U502 (N_502,N_487,N_412);
or U503 (N_503,N_473,N_430);
and U504 (N_504,N_498,N_422);
nor U505 (N_505,N_438,N_475);
xnor U506 (N_506,N_435,N_474);
and U507 (N_507,N_417,N_429);
and U508 (N_508,N_491,N_471);
and U509 (N_509,N_463,N_407);
nor U510 (N_510,N_446,N_458);
and U511 (N_511,N_424,N_468);
nor U512 (N_512,N_479,N_493);
or U513 (N_513,N_443,N_414);
or U514 (N_514,N_478,N_431);
nor U515 (N_515,N_403,N_425);
nor U516 (N_516,N_482,N_404);
and U517 (N_517,N_405,N_445);
nand U518 (N_518,N_467,N_413);
nor U519 (N_519,N_495,N_426);
nor U520 (N_520,N_428,N_454);
nor U521 (N_521,N_436,N_420);
and U522 (N_522,N_469,N_437);
or U523 (N_523,N_434,N_410);
or U524 (N_524,N_406,N_462);
and U525 (N_525,N_401,N_416);
or U526 (N_526,N_460,N_448);
nor U527 (N_527,N_411,N_464);
nor U528 (N_528,N_470,N_496);
and U529 (N_529,N_499,N_402);
nor U530 (N_530,N_441,N_408);
nor U531 (N_531,N_451,N_418);
nand U532 (N_532,N_423,N_409);
nor U533 (N_533,N_483,N_447);
nor U534 (N_534,N_472,N_461);
nand U535 (N_535,N_490,N_494);
or U536 (N_536,N_427,N_449);
and U537 (N_537,N_453,N_450);
and U538 (N_538,N_415,N_459);
nand U539 (N_539,N_465,N_485);
and U540 (N_540,N_484,N_452);
or U541 (N_541,N_440,N_400);
and U542 (N_542,N_444,N_481);
and U543 (N_543,N_432,N_419);
and U544 (N_544,N_497,N_442);
nand U545 (N_545,N_455,N_421);
nand U546 (N_546,N_466,N_476);
nor U547 (N_547,N_456,N_486);
xnor U548 (N_548,N_477,N_488);
nor U549 (N_549,N_480,N_492);
and U550 (N_550,N_427,N_419);
or U551 (N_551,N_422,N_455);
and U552 (N_552,N_425,N_440);
nor U553 (N_553,N_494,N_424);
nor U554 (N_554,N_464,N_426);
nand U555 (N_555,N_418,N_405);
nand U556 (N_556,N_485,N_428);
nand U557 (N_557,N_456,N_419);
and U558 (N_558,N_453,N_444);
and U559 (N_559,N_446,N_408);
and U560 (N_560,N_440,N_472);
nand U561 (N_561,N_453,N_465);
nand U562 (N_562,N_453,N_425);
or U563 (N_563,N_417,N_499);
nand U564 (N_564,N_431,N_452);
and U565 (N_565,N_476,N_487);
nor U566 (N_566,N_492,N_473);
and U567 (N_567,N_418,N_468);
nor U568 (N_568,N_405,N_413);
nand U569 (N_569,N_458,N_419);
xnor U570 (N_570,N_419,N_423);
xnor U571 (N_571,N_426,N_484);
nand U572 (N_572,N_490,N_488);
nand U573 (N_573,N_404,N_445);
and U574 (N_574,N_468,N_457);
and U575 (N_575,N_405,N_426);
nor U576 (N_576,N_415,N_478);
nand U577 (N_577,N_497,N_459);
nor U578 (N_578,N_459,N_477);
and U579 (N_579,N_474,N_473);
nor U580 (N_580,N_437,N_436);
nor U581 (N_581,N_429,N_449);
and U582 (N_582,N_421,N_477);
nand U583 (N_583,N_430,N_412);
and U584 (N_584,N_477,N_490);
nor U585 (N_585,N_497,N_414);
nand U586 (N_586,N_442,N_432);
nor U587 (N_587,N_417,N_413);
nand U588 (N_588,N_488,N_434);
nand U589 (N_589,N_408,N_486);
and U590 (N_590,N_400,N_485);
nand U591 (N_591,N_442,N_405);
or U592 (N_592,N_456,N_434);
nor U593 (N_593,N_404,N_442);
and U594 (N_594,N_472,N_432);
or U595 (N_595,N_429,N_442);
nor U596 (N_596,N_456,N_478);
nand U597 (N_597,N_401,N_444);
and U598 (N_598,N_495,N_422);
or U599 (N_599,N_407,N_444);
and U600 (N_600,N_531,N_504);
nor U601 (N_601,N_517,N_582);
and U602 (N_602,N_551,N_577);
or U603 (N_603,N_564,N_575);
nand U604 (N_604,N_533,N_562);
and U605 (N_605,N_572,N_509);
or U606 (N_606,N_569,N_502);
nand U607 (N_607,N_599,N_546);
or U608 (N_608,N_567,N_574);
or U609 (N_609,N_587,N_571);
and U610 (N_610,N_512,N_561);
nand U611 (N_611,N_588,N_583);
nor U612 (N_612,N_523,N_506);
and U613 (N_613,N_536,N_578);
nor U614 (N_614,N_503,N_552);
nor U615 (N_615,N_508,N_550);
nor U616 (N_616,N_511,N_521);
and U617 (N_617,N_522,N_535);
nor U618 (N_618,N_539,N_501);
nand U619 (N_619,N_515,N_544);
nand U620 (N_620,N_518,N_547);
nand U621 (N_621,N_557,N_568);
nand U622 (N_622,N_542,N_520);
or U623 (N_623,N_580,N_594);
nor U624 (N_624,N_526,N_591);
and U625 (N_625,N_585,N_528);
nand U626 (N_626,N_589,N_541);
and U627 (N_627,N_576,N_534);
or U628 (N_628,N_556,N_597);
or U629 (N_629,N_514,N_593);
and U630 (N_630,N_505,N_581);
nand U631 (N_631,N_570,N_553);
nand U632 (N_632,N_513,N_532);
and U633 (N_633,N_586,N_543);
nand U634 (N_634,N_530,N_598);
or U635 (N_635,N_549,N_558);
or U636 (N_636,N_563,N_525);
and U637 (N_637,N_510,N_555);
xnor U638 (N_638,N_559,N_596);
and U639 (N_639,N_500,N_565);
and U640 (N_640,N_590,N_554);
and U641 (N_641,N_519,N_560);
or U642 (N_642,N_507,N_524);
nor U643 (N_643,N_545,N_529);
or U644 (N_644,N_540,N_548);
nand U645 (N_645,N_527,N_537);
nand U646 (N_646,N_584,N_595);
nand U647 (N_647,N_579,N_573);
and U648 (N_648,N_592,N_516);
nor U649 (N_649,N_566,N_538);
and U650 (N_650,N_534,N_593);
nor U651 (N_651,N_529,N_534);
and U652 (N_652,N_599,N_572);
or U653 (N_653,N_515,N_533);
nand U654 (N_654,N_590,N_504);
and U655 (N_655,N_517,N_553);
or U656 (N_656,N_575,N_546);
or U657 (N_657,N_549,N_552);
or U658 (N_658,N_561,N_578);
or U659 (N_659,N_577,N_548);
nor U660 (N_660,N_517,N_552);
nand U661 (N_661,N_587,N_508);
nor U662 (N_662,N_593,N_589);
or U663 (N_663,N_585,N_525);
or U664 (N_664,N_599,N_511);
nand U665 (N_665,N_591,N_598);
nor U666 (N_666,N_503,N_517);
nand U667 (N_667,N_550,N_572);
nand U668 (N_668,N_533,N_544);
or U669 (N_669,N_542,N_540);
nor U670 (N_670,N_589,N_537);
xnor U671 (N_671,N_597,N_504);
or U672 (N_672,N_583,N_515);
or U673 (N_673,N_594,N_519);
nand U674 (N_674,N_549,N_535);
nor U675 (N_675,N_523,N_534);
and U676 (N_676,N_591,N_581);
and U677 (N_677,N_537,N_587);
or U678 (N_678,N_545,N_588);
or U679 (N_679,N_588,N_507);
nand U680 (N_680,N_514,N_511);
nand U681 (N_681,N_587,N_544);
nor U682 (N_682,N_517,N_546);
xnor U683 (N_683,N_554,N_593);
nor U684 (N_684,N_562,N_549);
and U685 (N_685,N_540,N_545);
or U686 (N_686,N_560,N_515);
nand U687 (N_687,N_508,N_502);
nor U688 (N_688,N_525,N_586);
or U689 (N_689,N_538,N_540);
and U690 (N_690,N_539,N_515);
nand U691 (N_691,N_518,N_587);
or U692 (N_692,N_573,N_531);
nor U693 (N_693,N_513,N_510);
nand U694 (N_694,N_588,N_590);
and U695 (N_695,N_579,N_565);
nand U696 (N_696,N_525,N_584);
nand U697 (N_697,N_599,N_549);
nand U698 (N_698,N_561,N_567);
or U699 (N_699,N_511,N_523);
nor U700 (N_700,N_669,N_619);
or U701 (N_701,N_629,N_672);
nor U702 (N_702,N_618,N_637);
nand U703 (N_703,N_646,N_684);
nand U704 (N_704,N_687,N_692);
nor U705 (N_705,N_647,N_658);
nor U706 (N_706,N_657,N_636);
or U707 (N_707,N_662,N_641);
and U708 (N_708,N_661,N_638);
and U709 (N_709,N_697,N_622);
nor U710 (N_710,N_627,N_664);
nor U711 (N_711,N_604,N_611);
or U712 (N_712,N_630,N_617);
nor U713 (N_713,N_624,N_612);
or U714 (N_714,N_674,N_600);
or U715 (N_715,N_660,N_693);
nor U716 (N_716,N_691,N_665);
or U717 (N_717,N_663,N_654);
and U718 (N_718,N_602,N_613);
and U719 (N_719,N_689,N_688);
or U720 (N_720,N_643,N_675);
and U721 (N_721,N_652,N_607);
nor U722 (N_722,N_606,N_685);
nand U723 (N_723,N_695,N_651);
nand U724 (N_724,N_620,N_655);
nor U725 (N_725,N_610,N_682);
and U726 (N_726,N_632,N_680);
and U727 (N_727,N_667,N_668);
and U728 (N_728,N_666,N_648);
nand U729 (N_729,N_642,N_681);
or U730 (N_730,N_694,N_656);
nand U731 (N_731,N_659,N_690);
nor U732 (N_732,N_678,N_616);
or U733 (N_733,N_614,N_609);
nand U734 (N_734,N_631,N_603);
xor U735 (N_735,N_605,N_679);
nor U736 (N_736,N_698,N_671);
or U737 (N_737,N_673,N_633);
or U738 (N_738,N_699,N_634);
nor U739 (N_739,N_608,N_644);
or U740 (N_740,N_626,N_615);
and U741 (N_741,N_621,N_635);
or U742 (N_742,N_686,N_625);
and U743 (N_743,N_601,N_683);
nor U744 (N_744,N_696,N_649);
or U745 (N_745,N_645,N_650);
nor U746 (N_746,N_677,N_640);
nand U747 (N_747,N_639,N_628);
or U748 (N_748,N_623,N_676);
nor U749 (N_749,N_670,N_653);
nor U750 (N_750,N_619,N_696);
and U751 (N_751,N_656,N_652);
and U752 (N_752,N_653,N_605);
nand U753 (N_753,N_640,N_649);
nor U754 (N_754,N_661,N_619);
nor U755 (N_755,N_643,N_657);
nand U756 (N_756,N_639,N_605);
nand U757 (N_757,N_670,N_688);
and U758 (N_758,N_609,N_674);
nor U759 (N_759,N_665,N_676);
and U760 (N_760,N_649,N_655);
and U761 (N_761,N_681,N_617);
nand U762 (N_762,N_603,N_649);
and U763 (N_763,N_630,N_640);
nor U764 (N_764,N_629,N_650);
or U765 (N_765,N_694,N_620);
and U766 (N_766,N_611,N_614);
nand U767 (N_767,N_655,N_619);
or U768 (N_768,N_693,N_607);
nor U769 (N_769,N_625,N_692);
and U770 (N_770,N_691,N_618);
nand U771 (N_771,N_610,N_695);
and U772 (N_772,N_677,N_655);
or U773 (N_773,N_683,N_691);
and U774 (N_774,N_673,N_651);
or U775 (N_775,N_612,N_677);
xor U776 (N_776,N_607,N_699);
or U777 (N_777,N_645,N_669);
nand U778 (N_778,N_617,N_687);
and U779 (N_779,N_696,N_607);
or U780 (N_780,N_663,N_638);
and U781 (N_781,N_682,N_654);
nor U782 (N_782,N_604,N_642);
nor U783 (N_783,N_690,N_652);
nand U784 (N_784,N_630,N_623);
nor U785 (N_785,N_698,N_611);
nand U786 (N_786,N_685,N_607);
nor U787 (N_787,N_675,N_618);
and U788 (N_788,N_693,N_623);
or U789 (N_789,N_600,N_669);
nor U790 (N_790,N_605,N_641);
or U791 (N_791,N_641,N_606);
nor U792 (N_792,N_641,N_686);
nand U793 (N_793,N_617,N_623);
nor U794 (N_794,N_632,N_618);
and U795 (N_795,N_691,N_627);
or U796 (N_796,N_657,N_616);
or U797 (N_797,N_631,N_691);
nand U798 (N_798,N_654,N_659);
and U799 (N_799,N_620,N_621);
or U800 (N_800,N_792,N_722);
and U801 (N_801,N_707,N_747);
and U802 (N_802,N_795,N_751);
and U803 (N_803,N_708,N_717);
or U804 (N_804,N_735,N_783);
nor U805 (N_805,N_720,N_742);
or U806 (N_806,N_715,N_701);
nor U807 (N_807,N_781,N_797);
and U808 (N_808,N_782,N_749);
nand U809 (N_809,N_787,N_765);
and U810 (N_810,N_790,N_719);
nor U811 (N_811,N_773,N_743);
or U812 (N_812,N_777,N_785);
nand U813 (N_813,N_744,N_703);
nor U814 (N_814,N_752,N_767);
or U815 (N_815,N_728,N_704);
nor U816 (N_816,N_753,N_726);
nor U817 (N_817,N_713,N_736);
nor U818 (N_818,N_725,N_706);
and U819 (N_819,N_780,N_796);
and U820 (N_820,N_770,N_724);
or U821 (N_821,N_764,N_779);
nand U822 (N_822,N_702,N_716);
nand U823 (N_823,N_729,N_798);
nand U824 (N_824,N_740,N_794);
and U825 (N_825,N_714,N_786);
nand U826 (N_826,N_756,N_776);
nand U827 (N_827,N_775,N_737);
and U828 (N_828,N_700,N_778);
nand U829 (N_829,N_799,N_754);
nor U830 (N_830,N_761,N_746);
and U831 (N_831,N_757,N_769);
nor U832 (N_832,N_738,N_709);
or U833 (N_833,N_759,N_727);
or U834 (N_834,N_788,N_748);
and U835 (N_835,N_741,N_721);
or U836 (N_836,N_745,N_784);
and U837 (N_837,N_772,N_730);
and U838 (N_838,N_731,N_750);
nor U839 (N_839,N_733,N_768);
and U840 (N_840,N_771,N_723);
and U841 (N_841,N_774,N_732);
and U842 (N_842,N_793,N_705);
or U843 (N_843,N_718,N_758);
nor U844 (N_844,N_739,N_755);
nand U845 (N_845,N_789,N_763);
nand U846 (N_846,N_760,N_791);
and U847 (N_847,N_710,N_734);
nor U848 (N_848,N_712,N_762);
nor U849 (N_849,N_766,N_711);
or U850 (N_850,N_702,N_785);
xor U851 (N_851,N_765,N_785);
or U852 (N_852,N_790,N_721);
or U853 (N_853,N_781,N_790);
nand U854 (N_854,N_755,N_701);
and U855 (N_855,N_754,N_779);
and U856 (N_856,N_790,N_740);
or U857 (N_857,N_790,N_770);
and U858 (N_858,N_700,N_740);
and U859 (N_859,N_777,N_760);
and U860 (N_860,N_703,N_771);
nand U861 (N_861,N_715,N_786);
or U862 (N_862,N_724,N_752);
nand U863 (N_863,N_731,N_723);
or U864 (N_864,N_716,N_728);
or U865 (N_865,N_739,N_737);
nor U866 (N_866,N_762,N_795);
nand U867 (N_867,N_772,N_799);
or U868 (N_868,N_738,N_733);
or U869 (N_869,N_700,N_705);
or U870 (N_870,N_717,N_753);
nor U871 (N_871,N_786,N_765);
or U872 (N_872,N_724,N_731);
and U873 (N_873,N_724,N_748);
nor U874 (N_874,N_716,N_727);
nor U875 (N_875,N_708,N_765);
or U876 (N_876,N_761,N_728);
nand U877 (N_877,N_705,N_786);
and U878 (N_878,N_759,N_715);
nor U879 (N_879,N_754,N_718);
nor U880 (N_880,N_726,N_789);
or U881 (N_881,N_720,N_758);
nand U882 (N_882,N_769,N_724);
and U883 (N_883,N_705,N_701);
and U884 (N_884,N_706,N_783);
nand U885 (N_885,N_717,N_723);
and U886 (N_886,N_714,N_709);
nand U887 (N_887,N_733,N_739);
nand U888 (N_888,N_757,N_747);
nand U889 (N_889,N_748,N_760);
or U890 (N_890,N_744,N_726);
nor U891 (N_891,N_727,N_784);
and U892 (N_892,N_765,N_799);
nor U893 (N_893,N_799,N_750);
nor U894 (N_894,N_792,N_720);
and U895 (N_895,N_713,N_751);
or U896 (N_896,N_770,N_710);
and U897 (N_897,N_776,N_784);
and U898 (N_898,N_713,N_777);
nand U899 (N_899,N_711,N_797);
or U900 (N_900,N_833,N_897);
nor U901 (N_901,N_812,N_860);
nand U902 (N_902,N_802,N_863);
and U903 (N_903,N_844,N_820);
and U904 (N_904,N_801,N_896);
nand U905 (N_905,N_835,N_865);
nand U906 (N_906,N_883,N_831);
nor U907 (N_907,N_858,N_848);
nand U908 (N_908,N_877,N_881);
nand U909 (N_909,N_888,N_815);
nand U910 (N_910,N_866,N_817);
or U911 (N_911,N_819,N_845);
and U912 (N_912,N_880,N_869);
nor U913 (N_913,N_895,N_874);
nand U914 (N_914,N_837,N_800);
and U915 (N_915,N_868,N_898);
nand U916 (N_916,N_856,N_809);
and U917 (N_917,N_829,N_867);
or U918 (N_918,N_872,N_825);
nor U919 (N_919,N_832,N_859);
nand U920 (N_920,N_852,N_854);
and U921 (N_921,N_830,N_839);
nand U922 (N_922,N_841,N_840);
or U923 (N_923,N_828,N_816);
and U924 (N_924,N_882,N_875);
and U925 (N_925,N_824,N_884);
and U926 (N_926,N_807,N_870);
and U927 (N_927,N_894,N_899);
or U928 (N_928,N_849,N_846);
nand U929 (N_929,N_803,N_842);
and U930 (N_930,N_822,N_864);
nor U931 (N_931,N_804,N_811);
nand U932 (N_932,N_827,N_889);
or U933 (N_933,N_826,N_850);
and U934 (N_934,N_810,N_893);
and U935 (N_935,N_885,N_806);
nor U936 (N_936,N_823,N_876);
nor U937 (N_937,N_879,N_890);
nand U938 (N_938,N_873,N_862);
nand U939 (N_939,N_857,N_834);
or U940 (N_940,N_813,N_808);
and U941 (N_941,N_892,N_838);
nor U942 (N_942,N_821,N_886);
and U943 (N_943,N_891,N_861);
or U944 (N_944,N_878,N_847);
nand U945 (N_945,N_851,N_887);
or U946 (N_946,N_805,N_814);
nand U947 (N_947,N_855,N_853);
or U948 (N_948,N_818,N_836);
and U949 (N_949,N_871,N_843);
and U950 (N_950,N_843,N_866);
nor U951 (N_951,N_813,N_817);
nand U952 (N_952,N_851,N_812);
or U953 (N_953,N_877,N_859);
or U954 (N_954,N_815,N_898);
nor U955 (N_955,N_821,N_842);
and U956 (N_956,N_868,N_862);
nor U957 (N_957,N_817,N_820);
and U958 (N_958,N_856,N_818);
nor U959 (N_959,N_856,N_814);
nand U960 (N_960,N_829,N_860);
and U961 (N_961,N_883,N_899);
nor U962 (N_962,N_865,N_849);
and U963 (N_963,N_806,N_812);
nor U964 (N_964,N_820,N_894);
and U965 (N_965,N_854,N_820);
nor U966 (N_966,N_829,N_834);
nand U967 (N_967,N_862,N_866);
and U968 (N_968,N_850,N_827);
nand U969 (N_969,N_817,N_850);
and U970 (N_970,N_843,N_816);
xor U971 (N_971,N_878,N_809);
or U972 (N_972,N_898,N_888);
nor U973 (N_973,N_857,N_831);
or U974 (N_974,N_891,N_800);
and U975 (N_975,N_847,N_857);
and U976 (N_976,N_805,N_815);
and U977 (N_977,N_846,N_831);
nand U978 (N_978,N_879,N_871);
and U979 (N_979,N_834,N_846);
and U980 (N_980,N_864,N_854);
nand U981 (N_981,N_821,N_826);
or U982 (N_982,N_863,N_850);
nand U983 (N_983,N_824,N_808);
nor U984 (N_984,N_810,N_860);
nor U985 (N_985,N_835,N_890);
nor U986 (N_986,N_839,N_863);
nand U987 (N_987,N_843,N_837);
nand U988 (N_988,N_837,N_824);
and U989 (N_989,N_819,N_878);
and U990 (N_990,N_873,N_861);
nand U991 (N_991,N_883,N_869);
nor U992 (N_992,N_882,N_831);
nor U993 (N_993,N_893,N_818);
nand U994 (N_994,N_861,N_894);
or U995 (N_995,N_879,N_806);
nand U996 (N_996,N_891,N_867);
and U997 (N_997,N_867,N_857);
nor U998 (N_998,N_825,N_804);
nor U999 (N_999,N_824,N_889);
nor U1000 (N_1000,N_929,N_997);
and U1001 (N_1001,N_947,N_918);
or U1002 (N_1002,N_914,N_967);
and U1003 (N_1003,N_973,N_946);
or U1004 (N_1004,N_976,N_992);
and U1005 (N_1005,N_954,N_987);
or U1006 (N_1006,N_906,N_931);
or U1007 (N_1007,N_936,N_960);
or U1008 (N_1008,N_958,N_905);
and U1009 (N_1009,N_942,N_979);
nand U1010 (N_1010,N_900,N_941);
nor U1011 (N_1011,N_911,N_993);
nand U1012 (N_1012,N_991,N_915);
nand U1013 (N_1013,N_933,N_969);
nand U1014 (N_1014,N_961,N_930);
nand U1015 (N_1015,N_998,N_980);
nor U1016 (N_1016,N_952,N_927);
nor U1017 (N_1017,N_925,N_985);
nor U1018 (N_1018,N_981,N_978);
nand U1019 (N_1019,N_943,N_913);
nand U1020 (N_1020,N_984,N_966);
and U1021 (N_1021,N_994,N_951);
and U1022 (N_1022,N_944,N_963);
and U1023 (N_1023,N_945,N_995);
or U1024 (N_1024,N_977,N_972);
xnor U1025 (N_1025,N_912,N_975);
nand U1026 (N_1026,N_937,N_970);
nor U1027 (N_1027,N_938,N_986);
and U1028 (N_1028,N_959,N_950);
nor U1029 (N_1029,N_955,N_919);
nor U1030 (N_1030,N_902,N_910);
or U1031 (N_1031,N_968,N_999);
or U1032 (N_1032,N_988,N_962);
and U1033 (N_1033,N_932,N_957);
or U1034 (N_1034,N_908,N_964);
and U1035 (N_1035,N_920,N_909);
and U1036 (N_1036,N_990,N_901);
or U1037 (N_1037,N_953,N_956);
and U1038 (N_1038,N_948,N_940);
nand U1039 (N_1039,N_917,N_949);
or U1040 (N_1040,N_974,N_926);
or U1041 (N_1041,N_907,N_928);
nor U1042 (N_1042,N_982,N_934);
nand U1043 (N_1043,N_923,N_916);
nor U1044 (N_1044,N_903,N_939);
nor U1045 (N_1045,N_989,N_922);
nand U1046 (N_1046,N_983,N_904);
nor U1047 (N_1047,N_924,N_921);
nor U1048 (N_1048,N_971,N_996);
nand U1049 (N_1049,N_935,N_965);
nor U1050 (N_1050,N_908,N_907);
and U1051 (N_1051,N_964,N_950);
or U1052 (N_1052,N_995,N_959);
nor U1053 (N_1053,N_917,N_996);
or U1054 (N_1054,N_918,N_964);
or U1055 (N_1055,N_993,N_961);
nor U1056 (N_1056,N_903,N_988);
and U1057 (N_1057,N_946,N_901);
nand U1058 (N_1058,N_972,N_920);
and U1059 (N_1059,N_904,N_930);
or U1060 (N_1060,N_935,N_970);
nand U1061 (N_1061,N_927,N_924);
nor U1062 (N_1062,N_945,N_971);
or U1063 (N_1063,N_926,N_965);
or U1064 (N_1064,N_979,N_912);
or U1065 (N_1065,N_930,N_991);
or U1066 (N_1066,N_997,N_902);
nor U1067 (N_1067,N_931,N_901);
and U1068 (N_1068,N_958,N_992);
nor U1069 (N_1069,N_995,N_935);
or U1070 (N_1070,N_946,N_986);
nand U1071 (N_1071,N_923,N_924);
or U1072 (N_1072,N_927,N_935);
nor U1073 (N_1073,N_973,N_965);
and U1074 (N_1074,N_965,N_987);
and U1075 (N_1075,N_925,N_900);
nor U1076 (N_1076,N_941,N_916);
nand U1077 (N_1077,N_971,N_974);
or U1078 (N_1078,N_925,N_981);
nand U1079 (N_1079,N_925,N_972);
or U1080 (N_1080,N_948,N_961);
nor U1081 (N_1081,N_995,N_920);
or U1082 (N_1082,N_916,N_938);
nand U1083 (N_1083,N_945,N_926);
nand U1084 (N_1084,N_926,N_942);
nand U1085 (N_1085,N_963,N_969);
and U1086 (N_1086,N_999,N_971);
nand U1087 (N_1087,N_999,N_946);
and U1088 (N_1088,N_903,N_975);
and U1089 (N_1089,N_979,N_972);
and U1090 (N_1090,N_952,N_901);
or U1091 (N_1091,N_907,N_964);
nand U1092 (N_1092,N_950,N_909);
and U1093 (N_1093,N_930,N_978);
and U1094 (N_1094,N_922,N_956);
nand U1095 (N_1095,N_958,N_910);
nor U1096 (N_1096,N_922,N_970);
nor U1097 (N_1097,N_928,N_910);
or U1098 (N_1098,N_935,N_953);
nor U1099 (N_1099,N_969,N_962);
xnor U1100 (N_1100,N_1064,N_1058);
nand U1101 (N_1101,N_1031,N_1057);
nor U1102 (N_1102,N_1024,N_1063);
nand U1103 (N_1103,N_1079,N_1048);
or U1104 (N_1104,N_1046,N_1001);
and U1105 (N_1105,N_1092,N_1081);
nand U1106 (N_1106,N_1020,N_1065);
nor U1107 (N_1107,N_1089,N_1072);
nand U1108 (N_1108,N_1038,N_1044);
and U1109 (N_1109,N_1022,N_1097);
and U1110 (N_1110,N_1066,N_1070);
or U1111 (N_1111,N_1034,N_1054);
or U1112 (N_1112,N_1042,N_1084);
and U1113 (N_1113,N_1026,N_1099);
nor U1114 (N_1114,N_1052,N_1069);
or U1115 (N_1115,N_1039,N_1027);
and U1116 (N_1116,N_1041,N_1021);
nand U1117 (N_1117,N_1028,N_1003);
nor U1118 (N_1118,N_1023,N_1004);
nand U1119 (N_1119,N_1088,N_1007);
or U1120 (N_1120,N_1029,N_1078);
nand U1121 (N_1121,N_1050,N_1037);
xnor U1122 (N_1122,N_1030,N_1040);
and U1123 (N_1123,N_1015,N_1091);
and U1124 (N_1124,N_1077,N_1080);
nand U1125 (N_1125,N_1036,N_1047);
nand U1126 (N_1126,N_1083,N_1045);
nor U1127 (N_1127,N_1060,N_1067);
and U1128 (N_1128,N_1017,N_1000);
or U1129 (N_1129,N_1082,N_1049);
nand U1130 (N_1130,N_1059,N_1014);
nor U1131 (N_1131,N_1053,N_1009);
and U1132 (N_1132,N_1035,N_1068);
nor U1133 (N_1133,N_1013,N_1086);
and U1134 (N_1134,N_1005,N_1096);
or U1135 (N_1135,N_1012,N_1095);
and U1136 (N_1136,N_1093,N_1032);
and U1137 (N_1137,N_1025,N_1051);
or U1138 (N_1138,N_1074,N_1016);
nand U1139 (N_1139,N_1055,N_1019);
or U1140 (N_1140,N_1056,N_1071);
nand U1141 (N_1141,N_1076,N_1010);
nand U1142 (N_1142,N_1011,N_1085);
nor U1143 (N_1143,N_1098,N_1008);
and U1144 (N_1144,N_1090,N_1006);
nor U1145 (N_1145,N_1062,N_1002);
or U1146 (N_1146,N_1018,N_1087);
or U1147 (N_1147,N_1094,N_1033);
and U1148 (N_1148,N_1073,N_1075);
nand U1149 (N_1149,N_1043,N_1061);
or U1150 (N_1150,N_1066,N_1078);
and U1151 (N_1151,N_1095,N_1032);
nand U1152 (N_1152,N_1030,N_1099);
nand U1153 (N_1153,N_1074,N_1053);
nand U1154 (N_1154,N_1094,N_1051);
nor U1155 (N_1155,N_1025,N_1003);
and U1156 (N_1156,N_1043,N_1007);
nand U1157 (N_1157,N_1062,N_1014);
nand U1158 (N_1158,N_1006,N_1017);
nand U1159 (N_1159,N_1057,N_1055);
nand U1160 (N_1160,N_1002,N_1026);
or U1161 (N_1161,N_1068,N_1078);
nor U1162 (N_1162,N_1050,N_1076);
or U1163 (N_1163,N_1065,N_1034);
nand U1164 (N_1164,N_1008,N_1051);
nor U1165 (N_1165,N_1066,N_1042);
and U1166 (N_1166,N_1038,N_1056);
nand U1167 (N_1167,N_1082,N_1074);
or U1168 (N_1168,N_1045,N_1033);
nor U1169 (N_1169,N_1034,N_1041);
nor U1170 (N_1170,N_1080,N_1051);
nand U1171 (N_1171,N_1020,N_1077);
and U1172 (N_1172,N_1013,N_1045);
nor U1173 (N_1173,N_1018,N_1003);
xnor U1174 (N_1174,N_1065,N_1009);
and U1175 (N_1175,N_1026,N_1009);
or U1176 (N_1176,N_1000,N_1030);
nor U1177 (N_1177,N_1002,N_1000);
nor U1178 (N_1178,N_1067,N_1061);
nand U1179 (N_1179,N_1052,N_1087);
nor U1180 (N_1180,N_1055,N_1017);
nand U1181 (N_1181,N_1054,N_1064);
nand U1182 (N_1182,N_1096,N_1058);
nor U1183 (N_1183,N_1086,N_1095);
and U1184 (N_1184,N_1054,N_1075);
or U1185 (N_1185,N_1037,N_1071);
nand U1186 (N_1186,N_1019,N_1062);
nor U1187 (N_1187,N_1023,N_1096);
or U1188 (N_1188,N_1039,N_1031);
nor U1189 (N_1189,N_1016,N_1034);
or U1190 (N_1190,N_1039,N_1086);
and U1191 (N_1191,N_1088,N_1016);
and U1192 (N_1192,N_1083,N_1054);
or U1193 (N_1193,N_1032,N_1068);
and U1194 (N_1194,N_1013,N_1020);
nand U1195 (N_1195,N_1056,N_1089);
or U1196 (N_1196,N_1006,N_1035);
or U1197 (N_1197,N_1072,N_1085);
nor U1198 (N_1198,N_1095,N_1034);
or U1199 (N_1199,N_1036,N_1033);
and U1200 (N_1200,N_1197,N_1178);
nor U1201 (N_1201,N_1103,N_1107);
nor U1202 (N_1202,N_1102,N_1146);
and U1203 (N_1203,N_1144,N_1169);
nor U1204 (N_1204,N_1176,N_1151);
and U1205 (N_1205,N_1118,N_1177);
and U1206 (N_1206,N_1181,N_1150);
and U1207 (N_1207,N_1171,N_1163);
xor U1208 (N_1208,N_1152,N_1175);
xor U1209 (N_1209,N_1128,N_1140);
or U1210 (N_1210,N_1159,N_1120);
nor U1211 (N_1211,N_1192,N_1122);
and U1212 (N_1212,N_1195,N_1139);
nand U1213 (N_1213,N_1137,N_1138);
or U1214 (N_1214,N_1148,N_1183);
or U1215 (N_1215,N_1133,N_1145);
and U1216 (N_1216,N_1104,N_1130);
nand U1217 (N_1217,N_1124,N_1131);
and U1218 (N_1218,N_1185,N_1114);
or U1219 (N_1219,N_1147,N_1193);
nor U1220 (N_1220,N_1165,N_1108);
nand U1221 (N_1221,N_1172,N_1100);
nor U1222 (N_1222,N_1123,N_1167);
or U1223 (N_1223,N_1153,N_1142);
nand U1224 (N_1224,N_1127,N_1141);
nand U1225 (N_1225,N_1154,N_1184);
and U1226 (N_1226,N_1164,N_1129);
or U1227 (N_1227,N_1199,N_1156);
or U1228 (N_1228,N_1143,N_1160);
or U1229 (N_1229,N_1187,N_1106);
nand U1230 (N_1230,N_1162,N_1136);
nor U1231 (N_1231,N_1119,N_1112);
and U1232 (N_1232,N_1135,N_1121);
nand U1233 (N_1233,N_1198,N_1173);
and U1234 (N_1234,N_1188,N_1157);
or U1235 (N_1235,N_1132,N_1125);
and U1236 (N_1236,N_1166,N_1179);
nand U1237 (N_1237,N_1101,N_1180);
or U1238 (N_1238,N_1168,N_1182);
and U1239 (N_1239,N_1134,N_1161);
or U1240 (N_1240,N_1109,N_1126);
nand U1241 (N_1241,N_1155,N_1190);
nor U1242 (N_1242,N_1196,N_1105);
and U1243 (N_1243,N_1186,N_1158);
and U1244 (N_1244,N_1116,N_1189);
or U1245 (N_1245,N_1170,N_1117);
or U1246 (N_1246,N_1194,N_1115);
or U1247 (N_1247,N_1191,N_1110);
nor U1248 (N_1248,N_1174,N_1149);
or U1249 (N_1249,N_1111,N_1113);
and U1250 (N_1250,N_1179,N_1150);
nand U1251 (N_1251,N_1141,N_1120);
xor U1252 (N_1252,N_1111,N_1161);
nand U1253 (N_1253,N_1189,N_1187);
nand U1254 (N_1254,N_1116,N_1147);
and U1255 (N_1255,N_1163,N_1109);
nand U1256 (N_1256,N_1100,N_1177);
nand U1257 (N_1257,N_1168,N_1170);
nor U1258 (N_1258,N_1174,N_1175);
nor U1259 (N_1259,N_1190,N_1123);
and U1260 (N_1260,N_1158,N_1126);
nand U1261 (N_1261,N_1128,N_1196);
nor U1262 (N_1262,N_1194,N_1191);
nor U1263 (N_1263,N_1145,N_1187);
and U1264 (N_1264,N_1120,N_1189);
nand U1265 (N_1265,N_1188,N_1116);
and U1266 (N_1266,N_1182,N_1112);
and U1267 (N_1267,N_1133,N_1157);
nor U1268 (N_1268,N_1184,N_1157);
or U1269 (N_1269,N_1196,N_1102);
nand U1270 (N_1270,N_1183,N_1130);
or U1271 (N_1271,N_1157,N_1123);
nor U1272 (N_1272,N_1185,N_1183);
and U1273 (N_1273,N_1158,N_1185);
nand U1274 (N_1274,N_1117,N_1164);
or U1275 (N_1275,N_1105,N_1134);
nor U1276 (N_1276,N_1104,N_1147);
and U1277 (N_1277,N_1150,N_1142);
or U1278 (N_1278,N_1140,N_1153);
nand U1279 (N_1279,N_1138,N_1160);
and U1280 (N_1280,N_1117,N_1100);
or U1281 (N_1281,N_1153,N_1143);
and U1282 (N_1282,N_1106,N_1112);
or U1283 (N_1283,N_1135,N_1167);
nor U1284 (N_1284,N_1105,N_1189);
or U1285 (N_1285,N_1101,N_1107);
and U1286 (N_1286,N_1182,N_1115);
and U1287 (N_1287,N_1187,N_1100);
nand U1288 (N_1288,N_1194,N_1143);
and U1289 (N_1289,N_1136,N_1132);
nand U1290 (N_1290,N_1125,N_1192);
nand U1291 (N_1291,N_1148,N_1124);
nor U1292 (N_1292,N_1132,N_1186);
nor U1293 (N_1293,N_1103,N_1129);
nor U1294 (N_1294,N_1190,N_1104);
and U1295 (N_1295,N_1194,N_1134);
nor U1296 (N_1296,N_1181,N_1183);
nor U1297 (N_1297,N_1103,N_1197);
or U1298 (N_1298,N_1127,N_1177);
and U1299 (N_1299,N_1101,N_1126);
or U1300 (N_1300,N_1231,N_1254);
nand U1301 (N_1301,N_1251,N_1269);
nor U1302 (N_1302,N_1236,N_1293);
nor U1303 (N_1303,N_1228,N_1256);
nor U1304 (N_1304,N_1289,N_1237);
nand U1305 (N_1305,N_1245,N_1259);
or U1306 (N_1306,N_1225,N_1285);
nor U1307 (N_1307,N_1253,N_1246);
or U1308 (N_1308,N_1276,N_1243);
nand U1309 (N_1309,N_1207,N_1217);
and U1310 (N_1310,N_1248,N_1252);
nor U1311 (N_1311,N_1263,N_1211);
or U1312 (N_1312,N_1216,N_1279);
nand U1313 (N_1313,N_1299,N_1203);
nand U1314 (N_1314,N_1204,N_1235);
or U1315 (N_1315,N_1264,N_1219);
and U1316 (N_1316,N_1233,N_1277);
nand U1317 (N_1317,N_1290,N_1273);
or U1318 (N_1318,N_1280,N_1242);
and U1319 (N_1319,N_1268,N_1260);
nand U1320 (N_1320,N_1227,N_1287);
nor U1321 (N_1321,N_1267,N_1257);
or U1322 (N_1322,N_1230,N_1292);
and U1323 (N_1323,N_1281,N_1229);
nor U1324 (N_1324,N_1221,N_1223);
nand U1325 (N_1325,N_1296,N_1206);
nand U1326 (N_1326,N_1222,N_1266);
or U1327 (N_1327,N_1265,N_1202);
or U1328 (N_1328,N_1294,N_1226);
or U1329 (N_1329,N_1271,N_1270);
or U1330 (N_1330,N_1232,N_1244);
and U1331 (N_1331,N_1241,N_1284);
and U1332 (N_1332,N_1297,N_1215);
and U1333 (N_1333,N_1238,N_1288);
nand U1334 (N_1334,N_1255,N_1298);
or U1335 (N_1335,N_1249,N_1261);
nand U1336 (N_1336,N_1201,N_1205);
nor U1337 (N_1337,N_1210,N_1200);
and U1338 (N_1338,N_1286,N_1220);
or U1339 (N_1339,N_1283,N_1282);
nor U1340 (N_1340,N_1240,N_1212);
nand U1341 (N_1341,N_1272,N_1208);
and U1342 (N_1342,N_1213,N_1275);
nor U1343 (N_1343,N_1262,N_1239);
nor U1344 (N_1344,N_1258,N_1291);
nor U1345 (N_1345,N_1209,N_1214);
and U1346 (N_1346,N_1250,N_1247);
and U1347 (N_1347,N_1234,N_1274);
and U1348 (N_1348,N_1295,N_1218);
nor U1349 (N_1349,N_1278,N_1224);
nand U1350 (N_1350,N_1211,N_1245);
nor U1351 (N_1351,N_1236,N_1204);
and U1352 (N_1352,N_1266,N_1251);
nor U1353 (N_1353,N_1262,N_1297);
and U1354 (N_1354,N_1212,N_1253);
nand U1355 (N_1355,N_1295,N_1219);
nand U1356 (N_1356,N_1228,N_1227);
nand U1357 (N_1357,N_1274,N_1291);
and U1358 (N_1358,N_1262,N_1220);
or U1359 (N_1359,N_1259,N_1295);
or U1360 (N_1360,N_1252,N_1274);
nor U1361 (N_1361,N_1293,N_1216);
nand U1362 (N_1362,N_1241,N_1263);
or U1363 (N_1363,N_1235,N_1269);
or U1364 (N_1364,N_1267,N_1223);
nor U1365 (N_1365,N_1291,N_1229);
and U1366 (N_1366,N_1234,N_1271);
nor U1367 (N_1367,N_1236,N_1273);
nor U1368 (N_1368,N_1236,N_1296);
nor U1369 (N_1369,N_1291,N_1250);
or U1370 (N_1370,N_1241,N_1267);
nand U1371 (N_1371,N_1224,N_1233);
nand U1372 (N_1372,N_1250,N_1239);
or U1373 (N_1373,N_1214,N_1217);
nor U1374 (N_1374,N_1264,N_1226);
and U1375 (N_1375,N_1299,N_1297);
nor U1376 (N_1376,N_1277,N_1211);
and U1377 (N_1377,N_1255,N_1273);
nand U1378 (N_1378,N_1279,N_1224);
and U1379 (N_1379,N_1298,N_1293);
nand U1380 (N_1380,N_1259,N_1235);
nor U1381 (N_1381,N_1221,N_1226);
or U1382 (N_1382,N_1267,N_1299);
nand U1383 (N_1383,N_1273,N_1221);
or U1384 (N_1384,N_1259,N_1282);
nand U1385 (N_1385,N_1254,N_1276);
nand U1386 (N_1386,N_1214,N_1263);
or U1387 (N_1387,N_1206,N_1282);
nor U1388 (N_1388,N_1235,N_1287);
and U1389 (N_1389,N_1250,N_1243);
and U1390 (N_1390,N_1261,N_1267);
and U1391 (N_1391,N_1299,N_1253);
or U1392 (N_1392,N_1288,N_1285);
nand U1393 (N_1393,N_1281,N_1221);
or U1394 (N_1394,N_1200,N_1279);
or U1395 (N_1395,N_1200,N_1288);
nor U1396 (N_1396,N_1207,N_1242);
nand U1397 (N_1397,N_1226,N_1268);
nand U1398 (N_1398,N_1207,N_1268);
nor U1399 (N_1399,N_1229,N_1286);
or U1400 (N_1400,N_1385,N_1349);
nand U1401 (N_1401,N_1342,N_1378);
or U1402 (N_1402,N_1303,N_1320);
or U1403 (N_1403,N_1368,N_1355);
and U1404 (N_1404,N_1361,N_1330);
nor U1405 (N_1405,N_1352,N_1309);
and U1406 (N_1406,N_1334,N_1381);
nor U1407 (N_1407,N_1371,N_1347);
nor U1408 (N_1408,N_1379,N_1364);
or U1409 (N_1409,N_1363,N_1338);
and U1410 (N_1410,N_1351,N_1344);
and U1411 (N_1411,N_1398,N_1380);
and U1412 (N_1412,N_1369,N_1337);
nand U1413 (N_1413,N_1393,N_1331);
nand U1414 (N_1414,N_1365,N_1374);
nor U1415 (N_1415,N_1373,N_1315);
or U1416 (N_1416,N_1307,N_1392);
or U1417 (N_1417,N_1383,N_1394);
and U1418 (N_1418,N_1318,N_1314);
nand U1419 (N_1419,N_1333,N_1335);
xor U1420 (N_1420,N_1304,N_1332);
and U1421 (N_1421,N_1395,N_1313);
nand U1422 (N_1422,N_1386,N_1327);
and U1423 (N_1423,N_1345,N_1359);
nor U1424 (N_1424,N_1343,N_1350);
nor U1425 (N_1425,N_1390,N_1356);
nor U1426 (N_1426,N_1375,N_1376);
nand U1427 (N_1427,N_1324,N_1340);
nor U1428 (N_1428,N_1366,N_1308);
nor U1429 (N_1429,N_1377,N_1310);
nand U1430 (N_1430,N_1321,N_1354);
nand U1431 (N_1431,N_1360,N_1382);
or U1432 (N_1432,N_1329,N_1312);
or U1433 (N_1433,N_1391,N_1325);
nor U1434 (N_1434,N_1399,N_1306);
and U1435 (N_1435,N_1370,N_1300);
nand U1436 (N_1436,N_1372,N_1316);
and U1437 (N_1437,N_1388,N_1302);
or U1438 (N_1438,N_1339,N_1384);
and U1439 (N_1439,N_1328,N_1358);
or U1440 (N_1440,N_1357,N_1305);
and U1441 (N_1441,N_1348,N_1396);
nand U1442 (N_1442,N_1346,N_1397);
or U1443 (N_1443,N_1336,N_1389);
nor U1444 (N_1444,N_1362,N_1326);
nor U1445 (N_1445,N_1311,N_1353);
nand U1446 (N_1446,N_1387,N_1323);
and U1447 (N_1447,N_1301,N_1341);
or U1448 (N_1448,N_1322,N_1367);
and U1449 (N_1449,N_1319,N_1317);
nor U1450 (N_1450,N_1362,N_1364);
nor U1451 (N_1451,N_1337,N_1345);
and U1452 (N_1452,N_1307,N_1395);
and U1453 (N_1453,N_1381,N_1339);
nand U1454 (N_1454,N_1313,N_1345);
and U1455 (N_1455,N_1391,N_1321);
nor U1456 (N_1456,N_1325,N_1398);
nor U1457 (N_1457,N_1315,N_1395);
or U1458 (N_1458,N_1382,N_1397);
nor U1459 (N_1459,N_1365,N_1345);
and U1460 (N_1460,N_1375,N_1328);
or U1461 (N_1461,N_1358,N_1341);
nand U1462 (N_1462,N_1303,N_1355);
and U1463 (N_1463,N_1309,N_1328);
nor U1464 (N_1464,N_1385,N_1381);
nand U1465 (N_1465,N_1315,N_1369);
nand U1466 (N_1466,N_1363,N_1396);
and U1467 (N_1467,N_1313,N_1364);
nor U1468 (N_1468,N_1308,N_1355);
nor U1469 (N_1469,N_1371,N_1360);
or U1470 (N_1470,N_1309,N_1332);
nand U1471 (N_1471,N_1378,N_1341);
or U1472 (N_1472,N_1396,N_1399);
or U1473 (N_1473,N_1310,N_1321);
and U1474 (N_1474,N_1308,N_1383);
nand U1475 (N_1475,N_1314,N_1358);
and U1476 (N_1476,N_1307,N_1310);
or U1477 (N_1477,N_1302,N_1308);
and U1478 (N_1478,N_1374,N_1361);
and U1479 (N_1479,N_1334,N_1343);
nand U1480 (N_1480,N_1320,N_1392);
and U1481 (N_1481,N_1310,N_1388);
or U1482 (N_1482,N_1371,N_1325);
nor U1483 (N_1483,N_1336,N_1395);
nand U1484 (N_1484,N_1343,N_1378);
nand U1485 (N_1485,N_1313,N_1352);
or U1486 (N_1486,N_1371,N_1312);
nor U1487 (N_1487,N_1333,N_1300);
nand U1488 (N_1488,N_1322,N_1352);
or U1489 (N_1489,N_1391,N_1300);
or U1490 (N_1490,N_1353,N_1360);
or U1491 (N_1491,N_1365,N_1321);
nor U1492 (N_1492,N_1330,N_1397);
nand U1493 (N_1493,N_1318,N_1338);
or U1494 (N_1494,N_1345,N_1321);
nor U1495 (N_1495,N_1376,N_1391);
or U1496 (N_1496,N_1370,N_1344);
nand U1497 (N_1497,N_1324,N_1314);
and U1498 (N_1498,N_1394,N_1339);
nand U1499 (N_1499,N_1348,N_1302);
or U1500 (N_1500,N_1422,N_1409);
or U1501 (N_1501,N_1431,N_1438);
nand U1502 (N_1502,N_1416,N_1419);
or U1503 (N_1503,N_1492,N_1487);
or U1504 (N_1504,N_1439,N_1453);
nor U1505 (N_1505,N_1496,N_1404);
nor U1506 (N_1506,N_1420,N_1459);
nor U1507 (N_1507,N_1433,N_1466);
nand U1508 (N_1508,N_1470,N_1418);
or U1509 (N_1509,N_1449,N_1405);
and U1510 (N_1510,N_1456,N_1414);
or U1511 (N_1511,N_1475,N_1445);
and U1512 (N_1512,N_1469,N_1442);
nor U1513 (N_1513,N_1450,N_1401);
nand U1514 (N_1514,N_1423,N_1421);
nand U1515 (N_1515,N_1479,N_1461);
nor U1516 (N_1516,N_1489,N_1432);
or U1517 (N_1517,N_1494,N_1463);
nor U1518 (N_1518,N_1444,N_1457);
nor U1519 (N_1519,N_1435,N_1478);
nor U1520 (N_1520,N_1408,N_1468);
nand U1521 (N_1521,N_1467,N_1499);
or U1522 (N_1522,N_1452,N_1437);
and U1523 (N_1523,N_1484,N_1415);
and U1524 (N_1524,N_1441,N_1460);
nand U1525 (N_1525,N_1491,N_1424);
and U1526 (N_1526,N_1473,N_1486);
nand U1527 (N_1527,N_1417,N_1498);
or U1528 (N_1528,N_1447,N_1476);
and U1529 (N_1529,N_1481,N_1471);
or U1530 (N_1530,N_1497,N_1426);
nor U1531 (N_1531,N_1406,N_1482);
nand U1532 (N_1532,N_1402,N_1410);
nor U1533 (N_1533,N_1464,N_1472);
nor U1534 (N_1534,N_1436,N_1493);
or U1535 (N_1535,N_1407,N_1425);
and U1536 (N_1536,N_1400,N_1451);
and U1537 (N_1537,N_1490,N_1495);
or U1538 (N_1538,N_1448,N_1465);
or U1539 (N_1539,N_1413,N_1412);
nor U1540 (N_1540,N_1411,N_1474);
nor U1541 (N_1541,N_1427,N_1428);
nand U1542 (N_1542,N_1434,N_1454);
or U1543 (N_1543,N_1440,N_1430);
and U1544 (N_1544,N_1462,N_1488);
and U1545 (N_1545,N_1485,N_1446);
or U1546 (N_1546,N_1480,N_1477);
nor U1547 (N_1547,N_1429,N_1443);
nor U1548 (N_1548,N_1455,N_1483);
nand U1549 (N_1549,N_1403,N_1458);
nor U1550 (N_1550,N_1424,N_1492);
nand U1551 (N_1551,N_1427,N_1417);
nor U1552 (N_1552,N_1493,N_1496);
and U1553 (N_1553,N_1447,N_1494);
and U1554 (N_1554,N_1425,N_1442);
nor U1555 (N_1555,N_1466,N_1491);
nor U1556 (N_1556,N_1406,N_1484);
or U1557 (N_1557,N_1411,N_1480);
and U1558 (N_1558,N_1467,N_1489);
nand U1559 (N_1559,N_1459,N_1433);
nor U1560 (N_1560,N_1446,N_1409);
nand U1561 (N_1561,N_1413,N_1482);
nand U1562 (N_1562,N_1434,N_1411);
nand U1563 (N_1563,N_1465,N_1423);
nand U1564 (N_1564,N_1419,N_1444);
and U1565 (N_1565,N_1487,N_1414);
xor U1566 (N_1566,N_1440,N_1446);
nand U1567 (N_1567,N_1465,N_1441);
nor U1568 (N_1568,N_1412,N_1431);
nand U1569 (N_1569,N_1443,N_1422);
and U1570 (N_1570,N_1444,N_1451);
and U1571 (N_1571,N_1407,N_1439);
nand U1572 (N_1572,N_1452,N_1453);
nor U1573 (N_1573,N_1482,N_1446);
or U1574 (N_1574,N_1454,N_1493);
and U1575 (N_1575,N_1455,N_1435);
nand U1576 (N_1576,N_1402,N_1407);
or U1577 (N_1577,N_1415,N_1452);
nor U1578 (N_1578,N_1403,N_1432);
nor U1579 (N_1579,N_1485,N_1475);
nor U1580 (N_1580,N_1415,N_1495);
and U1581 (N_1581,N_1466,N_1413);
nor U1582 (N_1582,N_1416,N_1472);
nand U1583 (N_1583,N_1424,N_1494);
nor U1584 (N_1584,N_1450,N_1490);
or U1585 (N_1585,N_1486,N_1401);
or U1586 (N_1586,N_1412,N_1445);
and U1587 (N_1587,N_1489,N_1479);
nand U1588 (N_1588,N_1470,N_1438);
nor U1589 (N_1589,N_1455,N_1401);
or U1590 (N_1590,N_1455,N_1460);
nor U1591 (N_1591,N_1472,N_1483);
or U1592 (N_1592,N_1407,N_1421);
and U1593 (N_1593,N_1487,N_1439);
or U1594 (N_1594,N_1483,N_1429);
or U1595 (N_1595,N_1459,N_1476);
nor U1596 (N_1596,N_1436,N_1401);
and U1597 (N_1597,N_1423,N_1457);
nand U1598 (N_1598,N_1431,N_1450);
nor U1599 (N_1599,N_1464,N_1479);
or U1600 (N_1600,N_1528,N_1504);
nor U1601 (N_1601,N_1578,N_1502);
nand U1602 (N_1602,N_1590,N_1539);
nor U1603 (N_1603,N_1547,N_1533);
and U1604 (N_1604,N_1513,N_1545);
and U1605 (N_1605,N_1520,N_1549);
nand U1606 (N_1606,N_1562,N_1551);
and U1607 (N_1607,N_1577,N_1574);
and U1608 (N_1608,N_1530,N_1519);
nand U1609 (N_1609,N_1514,N_1521);
nand U1610 (N_1610,N_1567,N_1535);
and U1611 (N_1611,N_1525,N_1589);
or U1612 (N_1612,N_1587,N_1524);
xnor U1613 (N_1613,N_1522,N_1536);
nor U1614 (N_1614,N_1596,N_1531);
nor U1615 (N_1615,N_1565,N_1512);
nor U1616 (N_1616,N_1588,N_1599);
or U1617 (N_1617,N_1540,N_1532);
nor U1618 (N_1618,N_1523,N_1576);
nand U1619 (N_1619,N_1557,N_1564);
nand U1620 (N_1620,N_1548,N_1580);
nand U1621 (N_1621,N_1500,N_1529);
or U1622 (N_1622,N_1586,N_1582);
or U1623 (N_1623,N_1591,N_1534);
xnor U1624 (N_1624,N_1595,N_1505);
or U1625 (N_1625,N_1509,N_1542);
or U1626 (N_1626,N_1511,N_1556);
or U1627 (N_1627,N_1526,N_1563);
nor U1628 (N_1628,N_1516,N_1553);
nor U1629 (N_1629,N_1570,N_1518);
or U1630 (N_1630,N_1543,N_1552);
or U1631 (N_1631,N_1503,N_1550);
or U1632 (N_1632,N_1544,N_1597);
and U1633 (N_1633,N_1555,N_1538);
nand U1634 (N_1634,N_1546,N_1584);
nand U1635 (N_1635,N_1537,N_1527);
nor U1636 (N_1636,N_1561,N_1581);
nand U1637 (N_1637,N_1585,N_1566);
nor U1638 (N_1638,N_1517,N_1593);
and U1639 (N_1639,N_1541,N_1575);
and U1640 (N_1640,N_1559,N_1560);
nor U1641 (N_1641,N_1507,N_1515);
nand U1642 (N_1642,N_1510,N_1508);
or U1643 (N_1643,N_1583,N_1594);
and U1644 (N_1644,N_1501,N_1558);
nand U1645 (N_1645,N_1592,N_1506);
and U1646 (N_1646,N_1579,N_1569);
nor U1647 (N_1647,N_1571,N_1554);
or U1648 (N_1648,N_1573,N_1598);
nor U1649 (N_1649,N_1572,N_1568);
or U1650 (N_1650,N_1537,N_1569);
and U1651 (N_1651,N_1584,N_1594);
or U1652 (N_1652,N_1545,N_1593);
or U1653 (N_1653,N_1555,N_1574);
and U1654 (N_1654,N_1532,N_1522);
and U1655 (N_1655,N_1566,N_1563);
and U1656 (N_1656,N_1597,N_1545);
or U1657 (N_1657,N_1509,N_1545);
and U1658 (N_1658,N_1526,N_1533);
nor U1659 (N_1659,N_1578,N_1511);
nand U1660 (N_1660,N_1586,N_1521);
and U1661 (N_1661,N_1589,N_1598);
nor U1662 (N_1662,N_1546,N_1531);
nand U1663 (N_1663,N_1547,N_1541);
and U1664 (N_1664,N_1552,N_1597);
and U1665 (N_1665,N_1561,N_1522);
and U1666 (N_1666,N_1571,N_1563);
nand U1667 (N_1667,N_1505,N_1560);
or U1668 (N_1668,N_1545,N_1563);
nand U1669 (N_1669,N_1530,N_1554);
and U1670 (N_1670,N_1549,N_1596);
nor U1671 (N_1671,N_1521,N_1565);
and U1672 (N_1672,N_1561,N_1589);
and U1673 (N_1673,N_1509,N_1511);
nor U1674 (N_1674,N_1553,N_1523);
and U1675 (N_1675,N_1545,N_1579);
nor U1676 (N_1676,N_1516,N_1513);
nor U1677 (N_1677,N_1529,N_1559);
nor U1678 (N_1678,N_1560,N_1520);
or U1679 (N_1679,N_1517,N_1557);
nor U1680 (N_1680,N_1534,N_1587);
or U1681 (N_1681,N_1531,N_1586);
nand U1682 (N_1682,N_1524,N_1527);
xor U1683 (N_1683,N_1569,N_1556);
nor U1684 (N_1684,N_1580,N_1571);
nor U1685 (N_1685,N_1500,N_1566);
and U1686 (N_1686,N_1591,N_1505);
or U1687 (N_1687,N_1544,N_1550);
nand U1688 (N_1688,N_1528,N_1553);
and U1689 (N_1689,N_1527,N_1581);
or U1690 (N_1690,N_1562,N_1573);
nand U1691 (N_1691,N_1596,N_1593);
nand U1692 (N_1692,N_1550,N_1522);
and U1693 (N_1693,N_1511,N_1535);
nor U1694 (N_1694,N_1566,N_1512);
nand U1695 (N_1695,N_1593,N_1535);
and U1696 (N_1696,N_1553,N_1562);
nand U1697 (N_1697,N_1520,N_1535);
nand U1698 (N_1698,N_1556,N_1565);
nor U1699 (N_1699,N_1502,N_1561);
nand U1700 (N_1700,N_1666,N_1668);
or U1701 (N_1701,N_1663,N_1657);
nor U1702 (N_1702,N_1670,N_1682);
and U1703 (N_1703,N_1676,N_1605);
and U1704 (N_1704,N_1631,N_1613);
and U1705 (N_1705,N_1677,N_1646);
nand U1706 (N_1706,N_1658,N_1681);
or U1707 (N_1707,N_1699,N_1632);
nor U1708 (N_1708,N_1662,N_1629);
nor U1709 (N_1709,N_1690,N_1624);
or U1710 (N_1710,N_1640,N_1698);
or U1711 (N_1711,N_1610,N_1696);
nor U1712 (N_1712,N_1679,N_1626);
or U1713 (N_1713,N_1619,N_1689);
nand U1714 (N_1714,N_1622,N_1636);
or U1715 (N_1715,N_1612,N_1683);
or U1716 (N_1716,N_1680,N_1604);
and U1717 (N_1717,N_1635,N_1606);
or U1718 (N_1718,N_1660,N_1695);
or U1719 (N_1719,N_1672,N_1625);
and U1720 (N_1720,N_1694,N_1639);
nand U1721 (N_1721,N_1609,N_1651);
and U1722 (N_1722,N_1652,N_1615);
or U1723 (N_1723,N_1684,N_1603);
or U1724 (N_1724,N_1618,N_1687);
nor U1725 (N_1725,N_1608,N_1616);
and U1726 (N_1726,N_1664,N_1621);
nand U1727 (N_1727,N_1661,N_1673);
nor U1728 (N_1728,N_1647,N_1678);
nor U1729 (N_1729,N_1685,N_1617);
or U1730 (N_1730,N_1637,N_1601);
nand U1731 (N_1731,N_1634,N_1697);
and U1732 (N_1732,N_1620,N_1686);
and U1733 (N_1733,N_1655,N_1674);
nor U1734 (N_1734,N_1671,N_1688);
nand U1735 (N_1735,N_1649,N_1669);
and U1736 (N_1736,N_1602,N_1656);
nand U1737 (N_1737,N_1693,N_1665);
nand U1738 (N_1738,N_1600,N_1653);
or U1739 (N_1739,N_1675,N_1614);
or U1740 (N_1740,N_1650,N_1667);
and U1741 (N_1741,N_1630,N_1642);
and U1742 (N_1742,N_1644,N_1638);
nor U1743 (N_1743,N_1654,N_1607);
and U1744 (N_1744,N_1691,N_1628);
nand U1745 (N_1745,N_1692,N_1633);
or U1746 (N_1746,N_1648,N_1643);
nand U1747 (N_1747,N_1659,N_1645);
or U1748 (N_1748,N_1623,N_1641);
or U1749 (N_1749,N_1611,N_1627);
and U1750 (N_1750,N_1625,N_1689);
and U1751 (N_1751,N_1629,N_1625);
nor U1752 (N_1752,N_1641,N_1620);
and U1753 (N_1753,N_1642,N_1659);
or U1754 (N_1754,N_1600,N_1679);
nand U1755 (N_1755,N_1686,N_1647);
nor U1756 (N_1756,N_1646,N_1611);
nand U1757 (N_1757,N_1637,N_1659);
and U1758 (N_1758,N_1642,N_1664);
or U1759 (N_1759,N_1693,N_1689);
nand U1760 (N_1760,N_1688,N_1657);
and U1761 (N_1761,N_1630,N_1699);
xnor U1762 (N_1762,N_1642,N_1683);
and U1763 (N_1763,N_1688,N_1624);
nor U1764 (N_1764,N_1695,N_1622);
nor U1765 (N_1765,N_1610,N_1692);
nor U1766 (N_1766,N_1608,N_1646);
nand U1767 (N_1767,N_1654,N_1688);
or U1768 (N_1768,N_1693,N_1637);
or U1769 (N_1769,N_1675,N_1688);
nand U1770 (N_1770,N_1620,N_1651);
nor U1771 (N_1771,N_1663,N_1610);
and U1772 (N_1772,N_1605,N_1691);
nand U1773 (N_1773,N_1600,N_1615);
and U1774 (N_1774,N_1623,N_1669);
nand U1775 (N_1775,N_1607,N_1652);
nor U1776 (N_1776,N_1612,N_1671);
nor U1777 (N_1777,N_1693,N_1615);
or U1778 (N_1778,N_1641,N_1687);
nor U1779 (N_1779,N_1697,N_1671);
or U1780 (N_1780,N_1654,N_1615);
nor U1781 (N_1781,N_1673,N_1694);
nand U1782 (N_1782,N_1608,N_1672);
or U1783 (N_1783,N_1695,N_1684);
nand U1784 (N_1784,N_1635,N_1600);
nor U1785 (N_1785,N_1600,N_1650);
and U1786 (N_1786,N_1626,N_1695);
nand U1787 (N_1787,N_1684,N_1685);
nand U1788 (N_1788,N_1681,N_1657);
or U1789 (N_1789,N_1651,N_1688);
nand U1790 (N_1790,N_1664,N_1657);
and U1791 (N_1791,N_1669,N_1655);
nor U1792 (N_1792,N_1617,N_1635);
or U1793 (N_1793,N_1669,N_1615);
nor U1794 (N_1794,N_1684,N_1676);
and U1795 (N_1795,N_1637,N_1688);
nand U1796 (N_1796,N_1639,N_1613);
nand U1797 (N_1797,N_1698,N_1643);
nand U1798 (N_1798,N_1653,N_1637);
and U1799 (N_1799,N_1670,N_1611);
and U1800 (N_1800,N_1756,N_1764);
nor U1801 (N_1801,N_1702,N_1735);
nor U1802 (N_1802,N_1758,N_1722);
nor U1803 (N_1803,N_1727,N_1723);
and U1804 (N_1804,N_1761,N_1798);
nor U1805 (N_1805,N_1714,N_1717);
nand U1806 (N_1806,N_1784,N_1705);
nand U1807 (N_1807,N_1730,N_1787);
nor U1808 (N_1808,N_1765,N_1703);
and U1809 (N_1809,N_1791,N_1708);
and U1810 (N_1810,N_1748,N_1778);
or U1811 (N_1811,N_1720,N_1795);
and U1812 (N_1812,N_1750,N_1709);
or U1813 (N_1813,N_1721,N_1736);
nand U1814 (N_1814,N_1719,N_1728);
nor U1815 (N_1815,N_1771,N_1785);
or U1816 (N_1816,N_1793,N_1700);
nand U1817 (N_1817,N_1743,N_1767);
nand U1818 (N_1818,N_1755,N_1786);
nor U1819 (N_1819,N_1760,N_1790);
and U1820 (N_1820,N_1742,N_1751);
and U1821 (N_1821,N_1770,N_1759);
nor U1822 (N_1822,N_1746,N_1763);
and U1823 (N_1823,N_1716,N_1773);
and U1824 (N_1824,N_1741,N_1766);
nand U1825 (N_1825,N_1725,N_1729);
nand U1826 (N_1826,N_1737,N_1779);
nor U1827 (N_1827,N_1749,N_1744);
nor U1828 (N_1828,N_1788,N_1774);
and U1829 (N_1829,N_1734,N_1776);
nor U1830 (N_1830,N_1738,N_1796);
nand U1831 (N_1831,N_1732,N_1733);
and U1832 (N_1832,N_1710,N_1726);
or U1833 (N_1833,N_1718,N_1794);
and U1834 (N_1834,N_1731,N_1711);
or U1835 (N_1835,N_1724,N_1740);
nor U1836 (N_1836,N_1792,N_1747);
nor U1837 (N_1837,N_1783,N_1715);
or U1838 (N_1838,N_1799,N_1701);
nand U1839 (N_1839,N_1789,N_1706);
nand U1840 (N_1840,N_1745,N_1752);
or U1841 (N_1841,N_1762,N_1768);
or U1842 (N_1842,N_1797,N_1707);
or U1843 (N_1843,N_1782,N_1739);
nand U1844 (N_1844,N_1712,N_1775);
and U1845 (N_1845,N_1757,N_1754);
or U1846 (N_1846,N_1704,N_1780);
nor U1847 (N_1847,N_1772,N_1777);
nor U1848 (N_1848,N_1753,N_1781);
or U1849 (N_1849,N_1769,N_1713);
or U1850 (N_1850,N_1759,N_1769);
nand U1851 (N_1851,N_1751,N_1761);
or U1852 (N_1852,N_1709,N_1746);
or U1853 (N_1853,N_1783,N_1756);
and U1854 (N_1854,N_1759,N_1765);
or U1855 (N_1855,N_1711,N_1704);
and U1856 (N_1856,N_1738,N_1761);
nand U1857 (N_1857,N_1731,N_1780);
nand U1858 (N_1858,N_1743,N_1719);
nand U1859 (N_1859,N_1705,N_1769);
and U1860 (N_1860,N_1756,N_1744);
nand U1861 (N_1861,N_1767,N_1718);
and U1862 (N_1862,N_1730,N_1739);
nor U1863 (N_1863,N_1703,N_1725);
or U1864 (N_1864,N_1763,N_1750);
or U1865 (N_1865,N_1734,N_1770);
and U1866 (N_1866,N_1725,N_1716);
nand U1867 (N_1867,N_1754,N_1718);
and U1868 (N_1868,N_1795,N_1737);
or U1869 (N_1869,N_1776,N_1708);
and U1870 (N_1870,N_1742,N_1710);
and U1871 (N_1871,N_1700,N_1779);
or U1872 (N_1872,N_1782,N_1783);
nand U1873 (N_1873,N_1707,N_1781);
and U1874 (N_1874,N_1783,N_1790);
nand U1875 (N_1875,N_1776,N_1709);
nand U1876 (N_1876,N_1791,N_1712);
and U1877 (N_1877,N_1723,N_1780);
nor U1878 (N_1878,N_1786,N_1734);
nor U1879 (N_1879,N_1711,N_1762);
xnor U1880 (N_1880,N_1775,N_1724);
nor U1881 (N_1881,N_1752,N_1737);
nand U1882 (N_1882,N_1797,N_1706);
nor U1883 (N_1883,N_1700,N_1797);
and U1884 (N_1884,N_1741,N_1731);
nand U1885 (N_1885,N_1732,N_1722);
nor U1886 (N_1886,N_1757,N_1738);
or U1887 (N_1887,N_1710,N_1727);
or U1888 (N_1888,N_1741,N_1757);
nand U1889 (N_1889,N_1763,N_1751);
nor U1890 (N_1890,N_1758,N_1754);
or U1891 (N_1891,N_1712,N_1772);
and U1892 (N_1892,N_1714,N_1796);
nand U1893 (N_1893,N_1788,N_1732);
nand U1894 (N_1894,N_1705,N_1793);
or U1895 (N_1895,N_1775,N_1748);
or U1896 (N_1896,N_1723,N_1729);
or U1897 (N_1897,N_1741,N_1745);
nand U1898 (N_1898,N_1739,N_1732);
nor U1899 (N_1899,N_1775,N_1788);
nand U1900 (N_1900,N_1879,N_1806);
or U1901 (N_1901,N_1812,N_1845);
and U1902 (N_1902,N_1853,N_1881);
or U1903 (N_1903,N_1895,N_1876);
nand U1904 (N_1904,N_1893,N_1805);
nor U1905 (N_1905,N_1835,N_1869);
nor U1906 (N_1906,N_1885,N_1852);
or U1907 (N_1907,N_1865,N_1892);
nor U1908 (N_1908,N_1886,N_1858);
and U1909 (N_1909,N_1841,N_1877);
or U1910 (N_1910,N_1833,N_1800);
or U1911 (N_1911,N_1888,N_1813);
and U1912 (N_1912,N_1820,N_1831);
or U1913 (N_1913,N_1856,N_1815);
nor U1914 (N_1914,N_1836,N_1880);
and U1915 (N_1915,N_1819,N_1842);
nor U1916 (N_1916,N_1882,N_1840);
nor U1917 (N_1917,N_1898,N_1871);
or U1918 (N_1918,N_1837,N_1846);
or U1919 (N_1919,N_1897,N_1811);
nand U1920 (N_1920,N_1807,N_1821);
and U1921 (N_1921,N_1875,N_1823);
nand U1922 (N_1922,N_1867,N_1894);
nand U1923 (N_1923,N_1822,N_1872);
or U1924 (N_1924,N_1851,N_1863);
and U1925 (N_1925,N_1816,N_1818);
nor U1926 (N_1926,N_1839,N_1884);
nor U1927 (N_1927,N_1817,N_1808);
or U1928 (N_1928,N_1868,N_1809);
or U1929 (N_1929,N_1825,N_1843);
nand U1930 (N_1930,N_1828,N_1878);
or U1931 (N_1931,N_1826,N_1857);
and U1932 (N_1932,N_1861,N_1896);
and U1933 (N_1933,N_1803,N_1870);
nor U1934 (N_1934,N_1889,N_1848);
nor U1935 (N_1935,N_1847,N_1834);
and U1936 (N_1936,N_1802,N_1859);
or U1937 (N_1937,N_1873,N_1860);
or U1938 (N_1938,N_1824,N_1887);
nand U1939 (N_1939,N_1829,N_1899);
and U1940 (N_1940,N_1814,N_1810);
or U1941 (N_1941,N_1844,N_1874);
or U1942 (N_1942,N_1801,N_1850);
and U1943 (N_1943,N_1804,N_1838);
or U1944 (N_1944,N_1891,N_1855);
or U1945 (N_1945,N_1827,N_1890);
and U1946 (N_1946,N_1862,N_1849);
and U1947 (N_1947,N_1883,N_1864);
and U1948 (N_1948,N_1866,N_1832);
or U1949 (N_1949,N_1854,N_1830);
or U1950 (N_1950,N_1810,N_1809);
nor U1951 (N_1951,N_1877,N_1804);
nand U1952 (N_1952,N_1810,N_1887);
and U1953 (N_1953,N_1819,N_1801);
nand U1954 (N_1954,N_1848,N_1845);
or U1955 (N_1955,N_1869,N_1880);
or U1956 (N_1956,N_1872,N_1884);
nor U1957 (N_1957,N_1868,N_1871);
xnor U1958 (N_1958,N_1821,N_1875);
nor U1959 (N_1959,N_1810,N_1846);
nor U1960 (N_1960,N_1873,N_1856);
and U1961 (N_1961,N_1896,N_1821);
nand U1962 (N_1962,N_1824,N_1823);
nor U1963 (N_1963,N_1874,N_1851);
and U1964 (N_1964,N_1852,N_1861);
nand U1965 (N_1965,N_1848,N_1870);
or U1966 (N_1966,N_1858,N_1891);
nand U1967 (N_1967,N_1851,N_1894);
and U1968 (N_1968,N_1877,N_1874);
nor U1969 (N_1969,N_1816,N_1810);
and U1970 (N_1970,N_1818,N_1810);
xnor U1971 (N_1971,N_1866,N_1804);
nor U1972 (N_1972,N_1885,N_1828);
nand U1973 (N_1973,N_1848,N_1823);
nor U1974 (N_1974,N_1892,N_1874);
nand U1975 (N_1975,N_1873,N_1880);
or U1976 (N_1976,N_1867,N_1896);
nor U1977 (N_1977,N_1866,N_1893);
or U1978 (N_1978,N_1853,N_1852);
nand U1979 (N_1979,N_1820,N_1850);
and U1980 (N_1980,N_1825,N_1820);
nor U1981 (N_1981,N_1879,N_1807);
and U1982 (N_1982,N_1843,N_1846);
and U1983 (N_1983,N_1808,N_1872);
nor U1984 (N_1984,N_1857,N_1849);
and U1985 (N_1985,N_1810,N_1839);
and U1986 (N_1986,N_1899,N_1889);
xor U1987 (N_1987,N_1807,N_1874);
nor U1988 (N_1988,N_1839,N_1850);
nor U1989 (N_1989,N_1870,N_1826);
nor U1990 (N_1990,N_1889,N_1857);
or U1991 (N_1991,N_1888,N_1859);
nor U1992 (N_1992,N_1899,N_1834);
nand U1993 (N_1993,N_1877,N_1839);
nor U1994 (N_1994,N_1833,N_1843);
nand U1995 (N_1995,N_1801,N_1892);
nand U1996 (N_1996,N_1807,N_1800);
nand U1997 (N_1997,N_1854,N_1836);
and U1998 (N_1998,N_1830,N_1804);
nand U1999 (N_1999,N_1877,N_1855);
and U2000 (N_2000,N_1952,N_1906);
nor U2001 (N_2001,N_1992,N_1981);
and U2002 (N_2002,N_1909,N_1922);
nand U2003 (N_2003,N_1964,N_1965);
nor U2004 (N_2004,N_1950,N_1969);
nand U2005 (N_2005,N_1963,N_1998);
nand U2006 (N_2006,N_1928,N_1924);
and U2007 (N_2007,N_1959,N_1915);
nor U2008 (N_2008,N_1962,N_1957);
and U2009 (N_2009,N_1900,N_1983);
and U2010 (N_2010,N_1933,N_1989);
nand U2011 (N_2011,N_1990,N_1901);
nand U2012 (N_2012,N_1960,N_1947);
nand U2013 (N_2013,N_1925,N_1934);
nor U2014 (N_2014,N_1910,N_1991);
nand U2015 (N_2015,N_1911,N_1953);
and U2016 (N_2016,N_1980,N_1971);
or U2017 (N_2017,N_1918,N_1919);
or U2018 (N_2018,N_1905,N_1994);
or U2019 (N_2019,N_1916,N_1967);
nand U2020 (N_2020,N_1974,N_1927);
or U2021 (N_2021,N_1939,N_1944);
and U2022 (N_2022,N_1943,N_1908);
nor U2023 (N_2023,N_1951,N_1940);
nor U2024 (N_2024,N_1945,N_1999);
or U2025 (N_2025,N_1904,N_1949);
and U2026 (N_2026,N_1946,N_1923);
and U2027 (N_2027,N_1937,N_1935);
and U2028 (N_2028,N_1987,N_1932);
nand U2029 (N_2029,N_1941,N_1982);
nand U2030 (N_2030,N_1931,N_1977);
and U2031 (N_2031,N_1917,N_1984);
nor U2032 (N_2032,N_1968,N_1948);
or U2033 (N_2033,N_1956,N_1976);
nor U2034 (N_2034,N_1929,N_1926);
and U2035 (N_2035,N_1970,N_1921);
nor U2036 (N_2036,N_1978,N_1954);
and U2037 (N_2037,N_1966,N_1930);
nand U2038 (N_2038,N_1936,N_1913);
and U2039 (N_2039,N_1942,N_1985);
or U2040 (N_2040,N_1958,N_1975);
and U2041 (N_2041,N_1920,N_1996);
and U2042 (N_2042,N_1972,N_1907);
or U2043 (N_2043,N_1997,N_1993);
or U2044 (N_2044,N_1902,N_1955);
nor U2045 (N_2045,N_1979,N_1973);
nor U2046 (N_2046,N_1914,N_1903);
nand U2047 (N_2047,N_1912,N_1995);
nand U2048 (N_2048,N_1988,N_1986);
nand U2049 (N_2049,N_1961,N_1938);
and U2050 (N_2050,N_1944,N_1925);
nand U2051 (N_2051,N_1931,N_1935);
nor U2052 (N_2052,N_1937,N_1981);
nand U2053 (N_2053,N_1968,N_1924);
nor U2054 (N_2054,N_1947,N_1984);
nor U2055 (N_2055,N_1915,N_1981);
nor U2056 (N_2056,N_1932,N_1902);
nor U2057 (N_2057,N_1953,N_1939);
or U2058 (N_2058,N_1944,N_1919);
nor U2059 (N_2059,N_1967,N_1996);
or U2060 (N_2060,N_1945,N_1962);
nor U2061 (N_2061,N_1920,N_1967);
and U2062 (N_2062,N_1967,N_1998);
nand U2063 (N_2063,N_1912,N_1996);
and U2064 (N_2064,N_1946,N_1901);
or U2065 (N_2065,N_1986,N_1968);
and U2066 (N_2066,N_1920,N_1926);
or U2067 (N_2067,N_1902,N_1900);
nand U2068 (N_2068,N_1954,N_1947);
or U2069 (N_2069,N_1909,N_1911);
and U2070 (N_2070,N_1918,N_1915);
and U2071 (N_2071,N_1981,N_1939);
or U2072 (N_2072,N_1928,N_1980);
nand U2073 (N_2073,N_1978,N_1902);
xnor U2074 (N_2074,N_1909,N_1961);
or U2075 (N_2075,N_1930,N_1943);
and U2076 (N_2076,N_1982,N_1951);
and U2077 (N_2077,N_1938,N_1958);
or U2078 (N_2078,N_1937,N_1900);
and U2079 (N_2079,N_1924,N_1927);
nor U2080 (N_2080,N_1989,N_1998);
or U2081 (N_2081,N_1972,N_1939);
and U2082 (N_2082,N_1969,N_1934);
nand U2083 (N_2083,N_1980,N_1908);
or U2084 (N_2084,N_1936,N_1945);
or U2085 (N_2085,N_1906,N_1911);
nor U2086 (N_2086,N_1906,N_1939);
nand U2087 (N_2087,N_1967,N_1993);
or U2088 (N_2088,N_1948,N_1993);
or U2089 (N_2089,N_1927,N_1930);
and U2090 (N_2090,N_1905,N_1960);
or U2091 (N_2091,N_1900,N_1913);
or U2092 (N_2092,N_1969,N_1911);
or U2093 (N_2093,N_1974,N_1948);
and U2094 (N_2094,N_1957,N_1979);
and U2095 (N_2095,N_1977,N_1904);
nand U2096 (N_2096,N_1900,N_1922);
nor U2097 (N_2097,N_1973,N_1990);
and U2098 (N_2098,N_1900,N_1979);
and U2099 (N_2099,N_1937,N_1902);
nand U2100 (N_2100,N_2084,N_2060);
or U2101 (N_2101,N_2017,N_2058);
or U2102 (N_2102,N_2015,N_2031);
nand U2103 (N_2103,N_2074,N_2081);
nand U2104 (N_2104,N_2048,N_2095);
and U2105 (N_2105,N_2042,N_2028);
and U2106 (N_2106,N_2008,N_2009);
nor U2107 (N_2107,N_2072,N_2023);
nor U2108 (N_2108,N_2027,N_2085);
nor U2109 (N_2109,N_2054,N_2014);
nor U2110 (N_2110,N_2099,N_2080);
and U2111 (N_2111,N_2030,N_2034);
nor U2112 (N_2112,N_2013,N_2019);
and U2113 (N_2113,N_2029,N_2063);
nor U2114 (N_2114,N_2018,N_2082);
nand U2115 (N_2115,N_2077,N_2020);
nor U2116 (N_2116,N_2079,N_2087);
nor U2117 (N_2117,N_2000,N_2024);
or U2118 (N_2118,N_2040,N_2075);
and U2119 (N_2119,N_2059,N_2002);
nor U2120 (N_2120,N_2041,N_2065);
nand U2121 (N_2121,N_2003,N_2096);
and U2122 (N_2122,N_2053,N_2061);
or U2123 (N_2123,N_2076,N_2064);
nand U2124 (N_2124,N_2055,N_2046);
and U2125 (N_2125,N_2078,N_2051);
nand U2126 (N_2126,N_2033,N_2089);
or U2127 (N_2127,N_2067,N_2032);
and U2128 (N_2128,N_2021,N_2049);
nor U2129 (N_2129,N_2069,N_2011);
nor U2130 (N_2130,N_2088,N_2037);
nor U2131 (N_2131,N_2025,N_2062);
and U2132 (N_2132,N_2004,N_2086);
or U2133 (N_2133,N_2038,N_2006);
nor U2134 (N_2134,N_2093,N_2098);
nor U2135 (N_2135,N_2012,N_2052);
and U2136 (N_2136,N_2094,N_2097);
and U2137 (N_2137,N_2083,N_2044);
and U2138 (N_2138,N_2092,N_2056);
or U2139 (N_2139,N_2001,N_2016);
and U2140 (N_2140,N_2071,N_2022);
nand U2141 (N_2141,N_2039,N_2007);
nor U2142 (N_2142,N_2035,N_2036);
nor U2143 (N_2143,N_2068,N_2091);
or U2144 (N_2144,N_2010,N_2045);
or U2145 (N_2145,N_2026,N_2090);
nand U2146 (N_2146,N_2057,N_2066);
and U2147 (N_2147,N_2050,N_2073);
nor U2148 (N_2148,N_2070,N_2047);
nand U2149 (N_2149,N_2043,N_2005);
nor U2150 (N_2150,N_2053,N_2045);
nor U2151 (N_2151,N_2085,N_2071);
and U2152 (N_2152,N_2057,N_2049);
or U2153 (N_2153,N_2060,N_2004);
or U2154 (N_2154,N_2017,N_2059);
nor U2155 (N_2155,N_2075,N_2021);
nand U2156 (N_2156,N_2005,N_2069);
nand U2157 (N_2157,N_2035,N_2043);
or U2158 (N_2158,N_2037,N_2036);
or U2159 (N_2159,N_2099,N_2073);
nand U2160 (N_2160,N_2096,N_2097);
nand U2161 (N_2161,N_2005,N_2062);
and U2162 (N_2162,N_2088,N_2047);
and U2163 (N_2163,N_2023,N_2056);
or U2164 (N_2164,N_2002,N_2076);
or U2165 (N_2165,N_2048,N_2063);
or U2166 (N_2166,N_2036,N_2044);
nand U2167 (N_2167,N_2060,N_2095);
and U2168 (N_2168,N_2044,N_2009);
nand U2169 (N_2169,N_2047,N_2010);
or U2170 (N_2170,N_2007,N_2079);
and U2171 (N_2171,N_2048,N_2046);
or U2172 (N_2172,N_2083,N_2088);
and U2173 (N_2173,N_2033,N_2031);
and U2174 (N_2174,N_2093,N_2002);
and U2175 (N_2175,N_2098,N_2072);
or U2176 (N_2176,N_2064,N_2085);
nand U2177 (N_2177,N_2063,N_2060);
and U2178 (N_2178,N_2046,N_2097);
or U2179 (N_2179,N_2068,N_2094);
nor U2180 (N_2180,N_2071,N_2003);
nand U2181 (N_2181,N_2033,N_2082);
nor U2182 (N_2182,N_2003,N_2069);
nor U2183 (N_2183,N_2064,N_2095);
or U2184 (N_2184,N_2080,N_2097);
nor U2185 (N_2185,N_2066,N_2019);
nor U2186 (N_2186,N_2022,N_2017);
nor U2187 (N_2187,N_2057,N_2074);
nor U2188 (N_2188,N_2062,N_2046);
nand U2189 (N_2189,N_2047,N_2063);
nand U2190 (N_2190,N_2012,N_2004);
nor U2191 (N_2191,N_2041,N_2016);
nand U2192 (N_2192,N_2029,N_2000);
nand U2193 (N_2193,N_2021,N_2040);
or U2194 (N_2194,N_2092,N_2018);
nor U2195 (N_2195,N_2091,N_2014);
nand U2196 (N_2196,N_2011,N_2092);
nor U2197 (N_2197,N_2088,N_2001);
nand U2198 (N_2198,N_2071,N_2014);
nor U2199 (N_2199,N_2067,N_2049);
nor U2200 (N_2200,N_2166,N_2131);
nand U2201 (N_2201,N_2102,N_2157);
or U2202 (N_2202,N_2187,N_2103);
or U2203 (N_2203,N_2156,N_2197);
nor U2204 (N_2204,N_2107,N_2120);
nor U2205 (N_2205,N_2100,N_2148);
nor U2206 (N_2206,N_2108,N_2167);
nor U2207 (N_2207,N_2149,N_2128);
or U2208 (N_2208,N_2199,N_2143);
or U2209 (N_2209,N_2147,N_2198);
and U2210 (N_2210,N_2171,N_2188);
nor U2211 (N_2211,N_2192,N_2181);
or U2212 (N_2212,N_2174,N_2165);
nand U2213 (N_2213,N_2138,N_2196);
nand U2214 (N_2214,N_2150,N_2112);
nor U2215 (N_2215,N_2104,N_2164);
and U2216 (N_2216,N_2117,N_2179);
nor U2217 (N_2217,N_2134,N_2124);
or U2218 (N_2218,N_2145,N_2175);
and U2219 (N_2219,N_2111,N_2189);
nand U2220 (N_2220,N_2169,N_2172);
and U2221 (N_2221,N_2126,N_2130);
nor U2222 (N_2222,N_2193,N_2144);
or U2223 (N_2223,N_2123,N_2159);
nor U2224 (N_2224,N_2125,N_2162);
and U2225 (N_2225,N_2121,N_2146);
nor U2226 (N_2226,N_2163,N_2106);
nand U2227 (N_2227,N_2113,N_2176);
or U2228 (N_2228,N_2151,N_2180);
nor U2229 (N_2229,N_2178,N_2119);
nand U2230 (N_2230,N_2141,N_2127);
nand U2231 (N_2231,N_2153,N_2190);
or U2232 (N_2232,N_2139,N_2168);
nor U2233 (N_2233,N_2105,N_2194);
and U2234 (N_2234,N_2155,N_2137);
and U2235 (N_2235,N_2132,N_2136);
or U2236 (N_2236,N_2140,N_2115);
nor U2237 (N_2237,N_2110,N_2184);
nor U2238 (N_2238,N_2195,N_2185);
and U2239 (N_2239,N_2161,N_2118);
nand U2240 (N_2240,N_2170,N_2191);
or U2241 (N_2241,N_2177,N_2183);
or U2242 (N_2242,N_2152,N_2160);
nand U2243 (N_2243,N_2182,N_2114);
and U2244 (N_2244,N_2186,N_2135);
and U2245 (N_2245,N_2122,N_2173);
nand U2246 (N_2246,N_2142,N_2116);
or U2247 (N_2247,N_2129,N_2158);
nand U2248 (N_2248,N_2109,N_2133);
or U2249 (N_2249,N_2101,N_2154);
nand U2250 (N_2250,N_2151,N_2110);
nand U2251 (N_2251,N_2149,N_2165);
and U2252 (N_2252,N_2124,N_2163);
or U2253 (N_2253,N_2112,N_2188);
nor U2254 (N_2254,N_2178,N_2128);
xnor U2255 (N_2255,N_2159,N_2167);
or U2256 (N_2256,N_2165,N_2180);
nor U2257 (N_2257,N_2115,N_2135);
or U2258 (N_2258,N_2179,N_2125);
or U2259 (N_2259,N_2157,N_2183);
or U2260 (N_2260,N_2170,N_2147);
or U2261 (N_2261,N_2147,N_2146);
or U2262 (N_2262,N_2191,N_2163);
nand U2263 (N_2263,N_2103,N_2162);
or U2264 (N_2264,N_2193,N_2109);
nand U2265 (N_2265,N_2198,N_2182);
nand U2266 (N_2266,N_2145,N_2136);
nor U2267 (N_2267,N_2190,N_2150);
and U2268 (N_2268,N_2178,N_2180);
and U2269 (N_2269,N_2104,N_2161);
or U2270 (N_2270,N_2181,N_2126);
nor U2271 (N_2271,N_2156,N_2159);
or U2272 (N_2272,N_2155,N_2166);
nor U2273 (N_2273,N_2151,N_2191);
nor U2274 (N_2274,N_2102,N_2194);
nand U2275 (N_2275,N_2186,N_2121);
or U2276 (N_2276,N_2195,N_2111);
and U2277 (N_2277,N_2185,N_2172);
nand U2278 (N_2278,N_2130,N_2136);
nand U2279 (N_2279,N_2173,N_2124);
or U2280 (N_2280,N_2179,N_2148);
nand U2281 (N_2281,N_2169,N_2189);
and U2282 (N_2282,N_2199,N_2174);
and U2283 (N_2283,N_2191,N_2139);
or U2284 (N_2284,N_2110,N_2176);
nor U2285 (N_2285,N_2145,N_2160);
or U2286 (N_2286,N_2120,N_2183);
nand U2287 (N_2287,N_2136,N_2171);
and U2288 (N_2288,N_2189,N_2155);
nor U2289 (N_2289,N_2150,N_2188);
or U2290 (N_2290,N_2178,N_2106);
and U2291 (N_2291,N_2106,N_2138);
or U2292 (N_2292,N_2194,N_2169);
or U2293 (N_2293,N_2176,N_2182);
and U2294 (N_2294,N_2184,N_2173);
and U2295 (N_2295,N_2124,N_2192);
nand U2296 (N_2296,N_2126,N_2170);
nor U2297 (N_2297,N_2169,N_2184);
and U2298 (N_2298,N_2196,N_2162);
or U2299 (N_2299,N_2134,N_2179);
nand U2300 (N_2300,N_2268,N_2204);
or U2301 (N_2301,N_2273,N_2210);
nor U2302 (N_2302,N_2242,N_2276);
nand U2303 (N_2303,N_2201,N_2226);
or U2304 (N_2304,N_2296,N_2209);
or U2305 (N_2305,N_2294,N_2272);
nor U2306 (N_2306,N_2257,N_2252);
nor U2307 (N_2307,N_2230,N_2298);
and U2308 (N_2308,N_2234,N_2216);
nor U2309 (N_2309,N_2241,N_2289);
and U2310 (N_2310,N_2202,N_2225);
and U2311 (N_2311,N_2227,N_2214);
or U2312 (N_2312,N_2215,N_2228);
xor U2313 (N_2313,N_2287,N_2278);
nand U2314 (N_2314,N_2208,N_2207);
nor U2315 (N_2315,N_2211,N_2256);
nand U2316 (N_2316,N_2229,N_2219);
and U2317 (N_2317,N_2212,N_2250);
nor U2318 (N_2318,N_2246,N_2240);
nand U2319 (N_2319,N_2275,N_2281);
nor U2320 (N_2320,N_2200,N_2279);
nor U2321 (N_2321,N_2249,N_2218);
nor U2322 (N_2322,N_2248,N_2264);
nor U2323 (N_2323,N_2295,N_2277);
or U2324 (N_2324,N_2221,N_2299);
nand U2325 (N_2325,N_2260,N_2203);
xor U2326 (N_2326,N_2238,N_2220);
nor U2327 (N_2327,N_2283,N_2266);
or U2328 (N_2328,N_2236,N_2244);
or U2329 (N_2329,N_2217,N_2269);
nor U2330 (N_2330,N_2274,N_2251);
and U2331 (N_2331,N_2286,N_2280);
or U2332 (N_2332,N_2245,N_2205);
nor U2333 (N_2333,N_2297,N_2290);
nor U2334 (N_2334,N_2265,N_2292);
nand U2335 (N_2335,N_2271,N_2243);
nand U2336 (N_2336,N_2284,N_2263);
nand U2337 (N_2337,N_2267,N_2288);
or U2338 (N_2338,N_2247,N_2255);
nor U2339 (N_2339,N_2239,N_2232);
nand U2340 (N_2340,N_2206,N_2222);
or U2341 (N_2341,N_2293,N_2213);
or U2342 (N_2342,N_2254,N_2258);
and U2343 (N_2343,N_2235,N_2224);
nor U2344 (N_2344,N_2285,N_2291);
nor U2345 (N_2345,N_2262,N_2282);
or U2346 (N_2346,N_2261,N_2253);
or U2347 (N_2347,N_2233,N_2237);
or U2348 (N_2348,N_2231,N_2259);
nor U2349 (N_2349,N_2270,N_2223);
or U2350 (N_2350,N_2232,N_2212);
xor U2351 (N_2351,N_2216,N_2256);
nor U2352 (N_2352,N_2292,N_2263);
and U2353 (N_2353,N_2288,N_2205);
or U2354 (N_2354,N_2269,N_2262);
and U2355 (N_2355,N_2257,N_2232);
or U2356 (N_2356,N_2252,N_2238);
nand U2357 (N_2357,N_2211,N_2247);
nand U2358 (N_2358,N_2217,N_2280);
nor U2359 (N_2359,N_2244,N_2251);
nor U2360 (N_2360,N_2210,N_2220);
or U2361 (N_2361,N_2203,N_2242);
nor U2362 (N_2362,N_2280,N_2223);
nor U2363 (N_2363,N_2285,N_2232);
nor U2364 (N_2364,N_2272,N_2230);
and U2365 (N_2365,N_2219,N_2248);
nand U2366 (N_2366,N_2217,N_2207);
or U2367 (N_2367,N_2237,N_2224);
nor U2368 (N_2368,N_2218,N_2242);
nand U2369 (N_2369,N_2297,N_2260);
or U2370 (N_2370,N_2291,N_2230);
nand U2371 (N_2371,N_2226,N_2292);
nand U2372 (N_2372,N_2216,N_2263);
nor U2373 (N_2373,N_2212,N_2267);
and U2374 (N_2374,N_2292,N_2202);
nand U2375 (N_2375,N_2267,N_2268);
nor U2376 (N_2376,N_2266,N_2236);
or U2377 (N_2377,N_2203,N_2209);
and U2378 (N_2378,N_2256,N_2282);
and U2379 (N_2379,N_2226,N_2286);
or U2380 (N_2380,N_2251,N_2252);
nor U2381 (N_2381,N_2206,N_2262);
nor U2382 (N_2382,N_2293,N_2237);
and U2383 (N_2383,N_2293,N_2219);
nand U2384 (N_2384,N_2267,N_2270);
nor U2385 (N_2385,N_2270,N_2241);
nor U2386 (N_2386,N_2215,N_2224);
and U2387 (N_2387,N_2209,N_2201);
nand U2388 (N_2388,N_2228,N_2207);
nand U2389 (N_2389,N_2207,N_2235);
and U2390 (N_2390,N_2247,N_2259);
or U2391 (N_2391,N_2213,N_2240);
or U2392 (N_2392,N_2222,N_2226);
nor U2393 (N_2393,N_2201,N_2294);
or U2394 (N_2394,N_2246,N_2291);
or U2395 (N_2395,N_2243,N_2250);
and U2396 (N_2396,N_2245,N_2280);
nor U2397 (N_2397,N_2254,N_2289);
nor U2398 (N_2398,N_2229,N_2224);
nor U2399 (N_2399,N_2225,N_2270);
nand U2400 (N_2400,N_2366,N_2364);
or U2401 (N_2401,N_2392,N_2372);
nor U2402 (N_2402,N_2397,N_2367);
and U2403 (N_2403,N_2342,N_2386);
nor U2404 (N_2404,N_2324,N_2321);
nor U2405 (N_2405,N_2334,N_2351);
nor U2406 (N_2406,N_2368,N_2359);
or U2407 (N_2407,N_2385,N_2379);
and U2408 (N_2408,N_2356,N_2352);
and U2409 (N_2409,N_2340,N_2345);
nand U2410 (N_2410,N_2317,N_2396);
and U2411 (N_2411,N_2312,N_2353);
and U2412 (N_2412,N_2399,N_2314);
or U2413 (N_2413,N_2393,N_2354);
nor U2414 (N_2414,N_2341,N_2388);
nor U2415 (N_2415,N_2311,N_2308);
and U2416 (N_2416,N_2316,N_2337);
nor U2417 (N_2417,N_2380,N_2306);
and U2418 (N_2418,N_2329,N_2344);
nor U2419 (N_2419,N_2384,N_2303);
xnor U2420 (N_2420,N_2326,N_2309);
and U2421 (N_2421,N_2325,N_2391);
nand U2422 (N_2422,N_2374,N_2383);
and U2423 (N_2423,N_2362,N_2347);
nand U2424 (N_2424,N_2377,N_2376);
nor U2425 (N_2425,N_2333,N_2373);
or U2426 (N_2426,N_2335,N_2305);
nor U2427 (N_2427,N_2328,N_2322);
nand U2428 (N_2428,N_2330,N_2360);
and U2429 (N_2429,N_2304,N_2361);
nor U2430 (N_2430,N_2338,N_2323);
and U2431 (N_2431,N_2319,N_2331);
or U2432 (N_2432,N_2355,N_2332);
or U2433 (N_2433,N_2395,N_2371);
nand U2434 (N_2434,N_2318,N_2349);
and U2435 (N_2435,N_2313,N_2394);
nor U2436 (N_2436,N_2302,N_2307);
nor U2437 (N_2437,N_2358,N_2369);
and U2438 (N_2438,N_2363,N_2390);
nand U2439 (N_2439,N_2320,N_2382);
and U2440 (N_2440,N_2339,N_2370);
and U2441 (N_2441,N_2315,N_2381);
or U2442 (N_2442,N_2389,N_2300);
nand U2443 (N_2443,N_2348,N_2336);
or U2444 (N_2444,N_2378,N_2398);
nand U2445 (N_2445,N_2346,N_2350);
or U2446 (N_2446,N_2387,N_2375);
nor U2447 (N_2447,N_2343,N_2365);
or U2448 (N_2448,N_2310,N_2301);
and U2449 (N_2449,N_2357,N_2327);
nor U2450 (N_2450,N_2352,N_2324);
and U2451 (N_2451,N_2333,N_2346);
or U2452 (N_2452,N_2371,N_2356);
or U2453 (N_2453,N_2374,N_2346);
nor U2454 (N_2454,N_2373,N_2371);
or U2455 (N_2455,N_2330,N_2307);
nor U2456 (N_2456,N_2357,N_2318);
nand U2457 (N_2457,N_2344,N_2350);
and U2458 (N_2458,N_2304,N_2391);
nor U2459 (N_2459,N_2387,N_2390);
or U2460 (N_2460,N_2322,N_2338);
xnor U2461 (N_2461,N_2394,N_2356);
nand U2462 (N_2462,N_2350,N_2327);
and U2463 (N_2463,N_2322,N_2350);
or U2464 (N_2464,N_2337,N_2360);
nor U2465 (N_2465,N_2306,N_2333);
nor U2466 (N_2466,N_2355,N_2329);
nand U2467 (N_2467,N_2325,N_2339);
or U2468 (N_2468,N_2358,N_2325);
nor U2469 (N_2469,N_2390,N_2344);
nand U2470 (N_2470,N_2369,N_2376);
or U2471 (N_2471,N_2345,N_2336);
nand U2472 (N_2472,N_2351,N_2320);
or U2473 (N_2473,N_2325,N_2324);
and U2474 (N_2474,N_2368,N_2305);
nand U2475 (N_2475,N_2313,N_2308);
and U2476 (N_2476,N_2377,N_2317);
and U2477 (N_2477,N_2341,N_2321);
nand U2478 (N_2478,N_2353,N_2317);
or U2479 (N_2479,N_2370,N_2391);
nand U2480 (N_2480,N_2359,N_2336);
nand U2481 (N_2481,N_2334,N_2324);
xnor U2482 (N_2482,N_2301,N_2340);
and U2483 (N_2483,N_2380,N_2394);
and U2484 (N_2484,N_2376,N_2386);
nand U2485 (N_2485,N_2312,N_2392);
or U2486 (N_2486,N_2345,N_2330);
nor U2487 (N_2487,N_2351,N_2341);
or U2488 (N_2488,N_2301,N_2372);
nand U2489 (N_2489,N_2310,N_2318);
and U2490 (N_2490,N_2322,N_2341);
nand U2491 (N_2491,N_2309,N_2308);
and U2492 (N_2492,N_2355,N_2363);
nor U2493 (N_2493,N_2341,N_2352);
nor U2494 (N_2494,N_2332,N_2340);
nor U2495 (N_2495,N_2357,N_2387);
and U2496 (N_2496,N_2330,N_2380);
and U2497 (N_2497,N_2351,N_2382);
or U2498 (N_2498,N_2344,N_2382);
or U2499 (N_2499,N_2333,N_2312);
and U2500 (N_2500,N_2432,N_2480);
or U2501 (N_2501,N_2461,N_2475);
nor U2502 (N_2502,N_2456,N_2429);
and U2503 (N_2503,N_2491,N_2498);
or U2504 (N_2504,N_2448,N_2420);
or U2505 (N_2505,N_2426,N_2441);
nand U2506 (N_2506,N_2451,N_2492);
nor U2507 (N_2507,N_2495,N_2442);
or U2508 (N_2508,N_2499,N_2427);
nand U2509 (N_2509,N_2490,N_2484);
or U2510 (N_2510,N_2488,N_2440);
nor U2511 (N_2511,N_2467,N_2469);
or U2512 (N_2512,N_2485,N_2411);
nor U2513 (N_2513,N_2470,N_2452);
or U2514 (N_2514,N_2455,N_2446);
and U2515 (N_2515,N_2439,N_2430);
nand U2516 (N_2516,N_2450,N_2415);
and U2517 (N_2517,N_2459,N_2412);
nor U2518 (N_2518,N_2425,N_2418);
and U2519 (N_2519,N_2458,N_2493);
nor U2520 (N_2520,N_2483,N_2403);
and U2521 (N_2521,N_2428,N_2416);
or U2522 (N_2522,N_2419,N_2486);
and U2523 (N_2523,N_2474,N_2407);
nor U2524 (N_2524,N_2404,N_2494);
nand U2525 (N_2525,N_2482,N_2472);
nor U2526 (N_2526,N_2460,N_2464);
nand U2527 (N_2527,N_2497,N_2479);
xnor U2528 (N_2528,N_2433,N_2405);
nand U2529 (N_2529,N_2487,N_2447);
nor U2530 (N_2530,N_2410,N_2465);
nand U2531 (N_2531,N_2434,N_2468);
or U2532 (N_2532,N_2424,N_2436);
nand U2533 (N_2533,N_2423,N_2496);
nand U2534 (N_2534,N_2402,N_2473);
nand U2535 (N_2535,N_2401,N_2462);
or U2536 (N_2536,N_2476,N_2422);
nor U2537 (N_2537,N_2463,N_2408);
nand U2538 (N_2538,N_2466,N_2431);
nor U2539 (N_2539,N_2437,N_2477);
and U2540 (N_2540,N_2443,N_2414);
nor U2541 (N_2541,N_2453,N_2471);
or U2542 (N_2542,N_2417,N_2435);
and U2543 (N_2543,N_2413,N_2489);
and U2544 (N_2544,N_2478,N_2449);
nor U2545 (N_2545,N_2421,N_2400);
or U2546 (N_2546,N_2444,N_2445);
or U2547 (N_2547,N_2454,N_2457);
nor U2548 (N_2548,N_2409,N_2438);
nand U2549 (N_2549,N_2481,N_2406);
and U2550 (N_2550,N_2424,N_2419);
nor U2551 (N_2551,N_2471,N_2434);
nand U2552 (N_2552,N_2490,N_2424);
nor U2553 (N_2553,N_2455,N_2415);
and U2554 (N_2554,N_2472,N_2442);
nand U2555 (N_2555,N_2426,N_2465);
and U2556 (N_2556,N_2484,N_2441);
or U2557 (N_2557,N_2444,N_2436);
nor U2558 (N_2558,N_2439,N_2429);
or U2559 (N_2559,N_2460,N_2407);
or U2560 (N_2560,N_2405,N_2469);
or U2561 (N_2561,N_2478,N_2495);
nor U2562 (N_2562,N_2410,N_2434);
and U2563 (N_2563,N_2498,N_2475);
and U2564 (N_2564,N_2421,N_2483);
nor U2565 (N_2565,N_2407,N_2487);
nor U2566 (N_2566,N_2430,N_2459);
or U2567 (N_2567,N_2417,N_2463);
nand U2568 (N_2568,N_2432,N_2406);
nor U2569 (N_2569,N_2455,N_2497);
nand U2570 (N_2570,N_2465,N_2424);
nor U2571 (N_2571,N_2459,N_2494);
xor U2572 (N_2572,N_2422,N_2430);
nor U2573 (N_2573,N_2434,N_2478);
nand U2574 (N_2574,N_2456,N_2487);
nand U2575 (N_2575,N_2447,N_2463);
nand U2576 (N_2576,N_2403,N_2406);
nor U2577 (N_2577,N_2441,N_2462);
or U2578 (N_2578,N_2409,N_2421);
and U2579 (N_2579,N_2491,N_2458);
nor U2580 (N_2580,N_2410,N_2472);
or U2581 (N_2581,N_2450,N_2433);
and U2582 (N_2582,N_2484,N_2440);
nand U2583 (N_2583,N_2480,N_2403);
or U2584 (N_2584,N_2495,N_2411);
and U2585 (N_2585,N_2417,N_2495);
and U2586 (N_2586,N_2481,N_2433);
nor U2587 (N_2587,N_2452,N_2456);
nand U2588 (N_2588,N_2413,N_2492);
and U2589 (N_2589,N_2424,N_2440);
and U2590 (N_2590,N_2420,N_2416);
nand U2591 (N_2591,N_2464,N_2456);
and U2592 (N_2592,N_2456,N_2415);
nand U2593 (N_2593,N_2488,N_2422);
and U2594 (N_2594,N_2406,N_2404);
nand U2595 (N_2595,N_2420,N_2485);
nand U2596 (N_2596,N_2446,N_2421);
nor U2597 (N_2597,N_2494,N_2421);
nand U2598 (N_2598,N_2418,N_2475);
and U2599 (N_2599,N_2463,N_2444);
or U2600 (N_2600,N_2578,N_2563);
nor U2601 (N_2601,N_2579,N_2559);
nand U2602 (N_2602,N_2523,N_2582);
or U2603 (N_2603,N_2521,N_2581);
nand U2604 (N_2604,N_2584,N_2537);
nor U2605 (N_2605,N_2575,N_2553);
nand U2606 (N_2606,N_2561,N_2535);
nor U2607 (N_2607,N_2515,N_2543);
nand U2608 (N_2608,N_2550,N_2549);
or U2609 (N_2609,N_2599,N_2597);
nor U2610 (N_2610,N_2539,N_2518);
and U2611 (N_2611,N_2514,N_2510);
nand U2612 (N_2612,N_2538,N_2595);
or U2613 (N_2613,N_2557,N_2560);
nand U2614 (N_2614,N_2577,N_2574);
and U2615 (N_2615,N_2567,N_2590);
nand U2616 (N_2616,N_2511,N_2500);
or U2617 (N_2617,N_2513,N_2516);
and U2618 (N_2618,N_2570,N_2585);
and U2619 (N_2619,N_2540,N_2503);
nor U2620 (N_2620,N_2542,N_2565);
and U2621 (N_2621,N_2576,N_2517);
and U2622 (N_2622,N_2558,N_2530);
and U2623 (N_2623,N_2527,N_2572);
or U2624 (N_2624,N_2544,N_2545);
or U2625 (N_2625,N_2522,N_2534);
or U2626 (N_2626,N_2508,N_2568);
and U2627 (N_2627,N_2592,N_2533);
or U2628 (N_2628,N_2598,N_2507);
and U2629 (N_2629,N_2509,N_2525);
nor U2630 (N_2630,N_2593,N_2512);
nand U2631 (N_2631,N_2588,N_2531);
nand U2632 (N_2632,N_2564,N_2562);
nand U2633 (N_2633,N_2519,N_2555);
nand U2634 (N_2634,N_2548,N_2583);
nor U2635 (N_2635,N_2524,N_2589);
nand U2636 (N_2636,N_2502,N_2591);
and U2637 (N_2637,N_2587,N_2554);
nor U2638 (N_2638,N_2596,N_2536);
and U2639 (N_2639,N_2552,N_2541);
nand U2640 (N_2640,N_2520,N_2551);
and U2641 (N_2641,N_2506,N_2569);
or U2642 (N_2642,N_2547,N_2501);
or U2643 (N_2643,N_2586,N_2594);
or U2644 (N_2644,N_2566,N_2505);
or U2645 (N_2645,N_2532,N_2504);
nor U2646 (N_2646,N_2529,N_2573);
nand U2647 (N_2647,N_2580,N_2526);
or U2648 (N_2648,N_2556,N_2546);
or U2649 (N_2649,N_2528,N_2571);
and U2650 (N_2650,N_2560,N_2561);
nand U2651 (N_2651,N_2543,N_2577);
nand U2652 (N_2652,N_2595,N_2554);
nand U2653 (N_2653,N_2585,N_2539);
or U2654 (N_2654,N_2512,N_2508);
and U2655 (N_2655,N_2556,N_2509);
or U2656 (N_2656,N_2564,N_2560);
nor U2657 (N_2657,N_2548,N_2584);
nor U2658 (N_2658,N_2558,N_2550);
nor U2659 (N_2659,N_2528,N_2562);
nor U2660 (N_2660,N_2514,N_2528);
and U2661 (N_2661,N_2500,N_2536);
and U2662 (N_2662,N_2578,N_2522);
nand U2663 (N_2663,N_2556,N_2582);
and U2664 (N_2664,N_2557,N_2587);
and U2665 (N_2665,N_2559,N_2569);
and U2666 (N_2666,N_2556,N_2592);
or U2667 (N_2667,N_2581,N_2503);
nor U2668 (N_2668,N_2565,N_2564);
nand U2669 (N_2669,N_2550,N_2561);
nor U2670 (N_2670,N_2553,N_2545);
and U2671 (N_2671,N_2509,N_2595);
nand U2672 (N_2672,N_2514,N_2540);
nand U2673 (N_2673,N_2560,N_2555);
nand U2674 (N_2674,N_2508,N_2555);
or U2675 (N_2675,N_2523,N_2552);
nand U2676 (N_2676,N_2541,N_2595);
nor U2677 (N_2677,N_2557,N_2532);
nand U2678 (N_2678,N_2532,N_2566);
nor U2679 (N_2679,N_2549,N_2519);
or U2680 (N_2680,N_2519,N_2569);
nor U2681 (N_2681,N_2524,N_2567);
nor U2682 (N_2682,N_2513,N_2567);
or U2683 (N_2683,N_2519,N_2502);
nand U2684 (N_2684,N_2576,N_2570);
or U2685 (N_2685,N_2547,N_2570);
nand U2686 (N_2686,N_2552,N_2562);
and U2687 (N_2687,N_2538,N_2557);
nand U2688 (N_2688,N_2566,N_2502);
nor U2689 (N_2689,N_2575,N_2510);
nor U2690 (N_2690,N_2559,N_2597);
nand U2691 (N_2691,N_2554,N_2506);
and U2692 (N_2692,N_2584,N_2594);
nand U2693 (N_2693,N_2558,N_2595);
and U2694 (N_2694,N_2541,N_2559);
and U2695 (N_2695,N_2533,N_2570);
nor U2696 (N_2696,N_2595,N_2533);
and U2697 (N_2697,N_2520,N_2534);
nand U2698 (N_2698,N_2571,N_2529);
and U2699 (N_2699,N_2545,N_2501);
or U2700 (N_2700,N_2606,N_2627);
or U2701 (N_2701,N_2671,N_2696);
nor U2702 (N_2702,N_2681,N_2624);
or U2703 (N_2703,N_2699,N_2648);
nand U2704 (N_2704,N_2677,N_2611);
or U2705 (N_2705,N_2662,N_2658);
or U2706 (N_2706,N_2687,N_2641);
nand U2707 (N_2707,N_2632,N_2666);
or U2708 (N_2708,N_2676,N_2689);
nor U2709 (N_2709,N_2633,N_2649);
or U2710 (N_2710,N_2665,N_2603);
nor U2711 (N_2711,N_2605,N_2613);
and U2712 (N_2712,N_2652,N_2634);
or U2713 (N_2713,N_2655,N_2646);
nand U2714 (N_2714,N_2674,N_2617);
and U2715 (N_2715,N_2683,N_2673);
and U2716 (N_2716,N_2610,N_2675);
nor U2717 (N_2717,N_2668,N_2688);
and U2718 (N_2718,N_2621,N_2615);
nor U2719 (N_2719,N_2691,N_2639);
and U2720 (N_2720,N_2653,N_2623);
nor U2721 (N_2721,N_2663,N_2670);
or U2722 (N_2722,N_2626,N_2614);
nor U2723 (N_2723,N_2612,N_2622);
nand U2724 (N_2724,N_2659,N_2651);
nor U2725 (N_2725,N_2620,N_2682);
nand U2726 (N_2726,N_2625,N_2660);
nor U2727 (N_2727,N_2604,N_2644);
or U2728 (N_2728,N_2616,N_2630);
nor U2729 (N_2729,N_2685,N_2654);
nand U2730 (N_2730,N_2647,N_2609);
nand U2731 (N_2731,N_2608,N_2631);
or U2732 (N_2732,N_2694,N_2680);
nand U2733 (N_2733,N_2645,N_2637);
nor U2734 (N_2734,N_2664,N_2635);
or U2735 (N_2735,N_2656,N_2693);
or U2736 (N_2736,N_2679,N_2686);
nor U2737 (N_2737,N_2643,N_2600);
or U2738 (N_2738,N_2661,N_2690);
nor U2739 (N_2739,N_2697,N_2692);
nand U2740 (N_2740,N_2669,N_2667);
or U2741 (N_2741,N_2602,N_2607);
and U2742 (N_2742,N_2636,N_2628);
nor U2743 (N_2743,N_2672,N_2601);
nand U2744 (N_2744,N_2629,N_2684);
or U2745 (N_2745,N_2698,N_2650);
and U2746 (N_2746,N_2618,N_2678);
and U2747 (N_2747,N_2642,N_2619);
nand U2748 (N_2748,N_2638,N_2657);
nor U2749 (N_2749,N_2695,N_2640);
nand U2750 (N_2750,N_2678,N_2621);
nand U2751 (N_2751,N_2690,N_2605);
or U2752 (N_2752,N_2672,N_2609);
nor U2753 (N_2753,N_2637,N_2609);
nand U2754 (N_2754,N_2629,N_2606);
and U2755 (N_2755,N_2614,N_2608);
or U2756 (N_2756,N_2644,N_2610);
or U2757 (N_2757,N_2666,N_2681);
and U2758 (N_2758,N_2635,N_2623);
or U2759 (N_2759,N_2618,N_2635);
nand U2760 (N_2760,N_2656,N_2610);
nor U2761 (N_2761,N_2680,N_2675);
nor U2762 (N_2762,N_2659,N_2686);
nor U2763 (N_2763,N_2624,N_2634);
or U2764 (N_2764,N_2613,N_2662);
and U2765 (N_2765,N_2622,N_2613);
nand U2766 (N_2766,N_2645,N_2651);
or U2767 (N_2767,N_2693,N_2688);
nor U2768 (N_2768,N_2601,N_2645);
and U2769 (N_2769,N_2603,N_2683);
nand U2770 (N_2770,N_2660,N_2662);
or U2771 (N_2771,N_2673,N_2691);
nor U2772 (N_2772,N_2634,N_2641);
or U2773 (N_2773,N_2618,N_2624);
or U2774 (N_2774,N_2640,N_2639);
nand U2775 (N_2775,N_2643,N_2695);
nand U2776 (N_2776,N_2634,N_2680);
and U2777 (N_2777,N_2666,N_2609);
and U2778 (N_2778,N_2668,N_2660);
nand U2779 (N_2779,N_2653,N_2612);
nor U2780 (N_2780,N_2654,N_2628);
and U2781 (N_2781,N_2640,N_2638);
nand U2782 (N_2782,N_2693,N_2623);
or U2783 (N_2783,N_2651,N_2663);
nand U2784 (N_2784,N_2654,N_2693);
nor U2785 (N_2785,N_2655,N_2680);
and U2786 (N_2786,N_2679,N_2611);
nand U2787 (N_2787,N_2673,N_2639);
nor U2788 (N_2788,N_2633,N_2627);
nand U2789 (N_2789,N_2638,N_2662);
nor U2790 (N_2790,N_2630,N_2646);
or U2791 (N_2791,N_2617,N_2653);
nand U2792 (N_2792,N_2629,N_2654);
and U2793 (N_2793,N_2693,N_2682);
and U2794 (N_2794,N_2657,N_2639);
nand U2795 (N_2795,N_2625,N_2627);
nand U2796 (N_2796,N_2609,N_2602);
nand U2797 (N_2797,N_2639,N_2698);
or U2798 (N_2798,N_2671,N_2650);
nand U2799 (N_2799,N_2684,N_2675);
nor U2800 (N_2800,N_2712,N_2749);
and U2801 (N_2801,N_2733,N_2780);
and U2802 (N_2802,N_2783,N_2796);
nand U2803 (N_2803,N_2767,N_2700);
or U2804 (N_2804,N_2707,N_2764);
or U2805 (N_2805,N_2770,N_2742);
nor U2806 (N_2806,N_2731,N_2797);
nor U2807 (N_2807,N_2761,N_2702);
nand U2808 (N_2808,N_2743,N_2759);
nor U2809 (N_2809,N_2762,N_2735);
and U2810 (N_2810,N_2785,N_2757);
nand U2811 (N_2811,N_2772,N_2737);
nand U2812 (N_2812,N_2798,N_2708);
or U2813 (N_2813,N_2769,N_2746);
or U2814 (N_2814,N_2787,N_2722);
nand U2815 (N_2815,N_2745,N_2738);
or U2816 (N_2816,N_2703,N_2747);
nand U2817 (N_2817,N_2799,N_2718);
nand U2818 (N_2818,N_2768,N_2732);
nand U2819 (N_2819,N_2771,N_2740);
or U2820 (N_2820,N_2776,N_2766);
or U2821 (N_2821,N_2778,N_2790);
or U2822 (N_2822,N_2713,N_2777);
or U2823 (N_2823,N_2717,N_2793);
and U2824 (N_2824,N_2788,N_2774);
nor U2825 (N_2825,N_2705,N_2724);
nand U2826 (N_2826,N_2752,N_2792);
and U2827 (N_2827,N_2781,N_2786);
and U2828 (N_2828,N_2789,N_2736);
nand U2829 (N_2829,N_2754,N_2760);
or U2830 (N_2830,N_2750,N_2701);
and U2831 (N_2831,N_2727,N_2711);
or U2832 (N_2832,N_2758,N_2773);
or U2833 (N_2833,N_2744,N_2706);
or U2834 (N_2834,N_2791,N_2728);
and U2835 (N_2835,N_2723,N_2714);
and U2836 (N_2836,N_2765,N_2710);
or U2837 (N_2837,N_2720,N_2734);
and U2838 (N_2838,N_2715,N_2741);
nor U2839 (N_2839,N_2755,N_2779);
nor U2840 (N_2840,N_2704,N_2794);
and U2841 (N_2841,N_2763,N_2748);
or U2842 (N_2842,N_2726,N_2721);
nand U2843 (N_2843,N_2716,N_2719);
and U2844 (N_2844,N_2753,N_2782);
or U2845 (N_2845,N_2729,N_2730);
nor U2846 (N_2846,N_2709,N_2725);
nor U2847 (N_2847,N_2775,N_2795);
and U2848 (N_2848,N_2784,N_2739);
or U2849 (N_2849,N_2751,N_2756);
nor U2850 (N_2850,N_2765,N_2759);
and U2851 (N_2851,N_2760,N_2776);
nand U2852 (N_2852,N_2764,N_2783);
or U2853 (N_2853,N_2741,N_2797);
or U2854 (N_2854,N_2714,N_2782);
or U2855 (N_2855,N_2798,N_2749);
xor U2856 (N_2856,N_2762,N_2755);
or U2857 (N_2857,N_2728,N_2757);
nand U2858 (N_2858,N_2791,N_2703);
nand U2859 (N_2859,N_2750,N_2779);
nand U2860 (N_2860,N_2795,N_2726);
nand U2861 (N_2861,N_2755,N_2719);
and U2862 (N_2862,N_2734,N_2728);
nor U2863 (N_2863,N_2720,N_2712);
or U2864 (N_2864,N_2715,N_2763);
and U2865 (N_2865,N_2790,N_2763);
nor U2866 (N_2866,N_2710,N_2719);
nand U2867 (N_2867,N_2760,N_2766);
nand U2868 (N_2868,N_2754,N_2775);
or U2869 (N_2869,N_2758,N_2742);
and U2870 (N_2870,N_2744,N_2704);
nand U2871 (N_2871,N_2704,N_2706);
and U2872 (N_2872,N_2786,N_2716);
and U2873 (N_2873,N_2720,N_2713);
nand U2874 (N_2874,N_2787,N_2783);
or U2875 (N_2875,N_2781,N_2713);
xnor U2876 (N_2876,N_2752,N_2762);
nor U2877 (N_2877,N_2765,N_2769);
or U2878 (N_2878,N_2781,N_2741);
and U2879 (N_2879,N_2789,N_2758);
nor U2880 (N_2880,N_2729,N_2702);
or U2881 (N_2881,N_2794,N_2701);
or U2882 (N_2882,N_2728,N_2720);
or U2883 (N_2883,N_2761,N_2726);
or U2884 (N_2884,N_2775,N_2794);
nand U2885 (N_2885,N_2742,N_2725);
and U2886 (N_2886,N_2711,N_2734);
or U2887 (N_2887,N_2755,N_2788);
nand U2888 (N_2888,N_2760,N_2785);
and U2889 (N_2889,N_2716,N_2736);
nand U2890 (N_2890,N_2748,N_2711);
nand U2891 (N_2891,N_2745,N_2721);
xnor U2892 (N_2892,N_2735,N_2738);
or U2893 (N_2893,N_2770,N_2794);
or U2894 (N_2894,N_2759,N_2796);
or U2895 (N_2895,N_2700,N_2728);
or U2896 (N_2896,N_2709,N_2769);
nand U2897 (N_2897,N_2795,N_2754);
or U2898 (N_2898,N_2719,N_2703);
xor U2899 (N_2899,N_2775,N_2728);
and U2900 (N_2900,N_2827,N_2807);
nand U2901 (N_2901,N_2853,N_2898);
nor U2902 (N_2902,N_2835,N_2842);
nor U2903 (N_2903,N_2830,N_2886);
nand U2904 (N_2904,N_2848,N_2809);
or U2905 (N_2905,N_2802,N_2892);
nor U2906 (N_2906,N_2836,N_2808);
nand U2907 (N_2907,N_2803,N_2881);
nor U2908 (N_2908,N_2871,N_2819);
nor U2909 (N_2909,N_2899,N_2846);
and U2910 (N_2910,N_2818,N_2862);
and U2911 (N_2911,N_2888,N_2890);
nor U2912 (N_2912,N_2882,N_2864);
or U2913 (N_2913,N_2851,N_2816);
and U2914 (N_2914,N_2840,N_2884);
or U2915 (N_2915,N_2875,N_2887);
nand U2916 (N_2916,N_2863,N_2852);
and U2917 (N_2917,N_2877,N_2831);
and U2918 (N_2918,N_2815,N_2820);
nor U2919 (N_2919,N_2874,N_2883);
nand U2920 (N_2920,N_2872,N_2861);
or U2921 (N_2921,N_2858,N_2814);
and U2922 (N_2922,N_2829,N_2839);
nor U2923 (N_2923,N_2873,N_2832);
or U2924 (N_2924,N_2879,N_2843);
or U2925 (N_2925,N_2868,N_2896);
nor U2926 (N_2926,N_2893,N_2854);
nand U2927 (N_2927,N_2833,N_2876);
nand U2928 (N_2928,N_2878,N_2824);
or U2929 (N_2929,N_2822,N_2817);
nor U2930 (N_2930,N_2823,N_2804);
and U2931 (N_2931,N_2845,N_2850);
or U2932 (N_2932,N_2880,N_2821);
and U2933 (N_2933,N_2811,N_2800);
nand U2934 (N_2934,N_2891,N_2885);
or U2935 (N_2935,N_2834,N_2870);
or U2936 (N_2936,N_2865,N_2844);
nor U2937 (N_2937,N_2856,N_2805);
or U2938 (N_2938,N_2860,N_2857);
nand U2939 (N_2939,N_2869,N_2866);
or U2940 (N_2940,N_2810,N_2889);
or U2941 (N_2941,N_2813,N_2855);
nand U2942 (N_2942,N_2849,N_2837);
nand U2943 (N_2943,N_2826,N_2806);
and U2944 (N_2944,N_2841,N_2897);
nor U2945 (N_2945,N_2812,N_2828);
or U2946 (N_2946,N_2895,N_2847);
and U2947 (N_2947,N_2894,N_2859);
nor U2948 (N_2948,N_2801,N_2825);
and U2949 (N_2949,N_2838,N_2867);
nor U2950 (N_2950,N_2868,N_2846);
nand U2951 (N_2951,N_2846,N_2839);
nand U2952 (N_2952,N_2846,N_2876);
nand U2953 (N_2953,N_2884,N_2821);
nor U2954 (N_2954,N_2817,N_2804);
and U2955 (N_2955,N_2887,N_2829);
nand U2956 (N_2956,N_2860,N_2815);
or U2957 (N_2957,N_2818,N_2853);
nor U2958 (N_2958,N_2861,N_2865);
and U2959 (N_2959,N_2822,N_2890);
or U2960 (N_2960,N_2859,N_2830);
or U2961 (N_2961,N_2833,N_2886);
or U2962 (N_2962,N_2820,N_2834);
nor U2963 (N_2963,N_2801,N_2832);
or U2964 (N_2964,N_2875,N_2885);
and U2965 (N_2965,N_2858,N_2868);
or U2966 (N_2966,N_2858,N_2801);
or U2967 (N_2967,N_2833,N_2832);
or U2968 (N_2968,N_2831,N_2879);
or U2969 (N_2969,N_2829,N_2827);
and U2970 (N_2970,N_2826,N_2861);
nor U2971 (N_2971,N_2816,N_2855);
or U2972 (N_2972,N_2848,N_2840);
nand U2973 (N_2973,N_2848,N_2825);
nand U2974 (N_2974,N_2868,N_2854);
and U2975 (N_2975,N_2846,N_2892);
or U2976 (N_2976,N_2853,N_2800);
nor U2977 (N_2977,N_2818,N_2816);
nand U2978 (N_2978,N_2890,N_2840);
or U2979 (N_2979,N_2882,N_2818);
nand U2980 (N_2980,N_2857,N_2895);
nand U2981 (N_2981,N_2822,N_2805);
and U2982 (N_2982,N_2892,N_2828);
or U2983 (N_2983,N_2885,N_2812);
or U2984 (N_2984,N_2858,N_2849);
nor U2985 (N_2985,N_2814,N_2816);
or U2986 (N_2986,N_2895,N_2894);
and U2987 (N_2987,N_2880,N_2833);
nand U2988 (N_2988,N_2866,N_2855);
or U2989 (N_2989,N_2824,N_2801);
or U2990 (N_2990,N_2813,N_2854);
or U2991 (N_2991,N_2802,N_2812);
and U2992 (N_2992,N_2824,N_2850);
nor U2993 (N_2993,N_2898,N_2836);
nand U2994 (N_2994,N_2884,N_2839);
and U2995 (N_2995,N_2891,N_2808);
nand U2996 (N_2996,N_2827,N_2839);
nand U2997 (N_2997,N_2892,N_2849);
or U2998 (N_2998,N_2834,N_2880);
nor U2999 (N_2999,N_2856,N_2895);
nand UO_0 (O_0,N_2920,N_2913);
xor UO_1 (O_1,N_2944,N_2963);
and UO_2 (O_2,N_2960,N_2950);
and UO_3 (O_3,N_2982,N_2974);
nor UO_4 (O_4,N_2917,N_2957);
or UO_5 (O_5,N_2969,N_2933);
nand UO_6 (O_6,N_2901,N_2915);
and UO_7 (O_7,N_2996,N_2945);
nor UO_8 (O_8,N_2967,N_2987);
and UO_9 (O_9,N_2977,N_2991);
and UO_10 (O_10,N_2946,N_2995);
or UO_11 (O_11,N_2981,N_2926);
and UO_12 (O_12,N_2904,N_2902);
and UO_13 (O_13,N_2951,N_2999);
and UO_14 (O_14,N_2972,N_2927);
or UO_15 (O_15,N_2984,N_2923);
or UO_16 (O_16,N_2906,N_2964);
and UO_17 (O_17,N_2986,N_2905);
nand UO_18 (O_18,N_2962,N_2966);
nor UO_19 (O_19,N_2975,N_2997);
and UO_20 (O_20,N_2956,N_2983);
nand UO_21 (O_21,N_2958,N_2989);
and UO_22 (O_22,N_2925,N_2919);
nand UO_23 (O_23,N_2914,N_2993);
and UO_24 (O_24,N_2911,N_2968);
nand UO_25 (O_25,N_2943,N_2955);
and UO_26 (O_26,N_2979,N_2978);
nor UO_27 (O_27,N_2922,N_2932);
nand UO_28 (O_28,N_2970,N_2907);
or UO_29 (O_29,N_2936,N_2998);
and UO_30 (O_30,N_2934,N_2908);
or UO_31 (O_31,N_2994,N_2924);
nand UO_32 (O_32,N_2961,N_2935);
nand UO_33 (O_33,N_2985,N_2941);
and UO_34 (O_34,N_2988,N_2939);
nor UO_35 (O_35,N_2949,N_2990);
or UO_36 (O_36,N_2948,N_2959);
and UO_37 (O_37,N_2930,N_2929);
nand UO_38 (O_38,N_2910,N_2980);
or UO_39 (O_39,N_2909,N_2903);
or UO_40 (O_40,N_2942,N_2953);
nor UO_41 (O_41,N_2916,N_2992);
or UO_42 (O_42,N_2940,N_2900);
or UO_43 (O_43,N_2921,N_2938);
and UO_44 (O_44,N_2965,N_2976);
or UO_45 (O_45,N_2931,N_2918);
nor UO_46 (O_46,N_2928,N_2971);
and UO_47 (O_47,N_2947,N_2954);
nor UO_48 (O_48,N_2952,N_2973);
or UO_49 (O_49,N_2937,N_2912);
nor UO_50 (O_50,N_2935,N_2937);
and UO_51 (O_51,N_2957,N_2990);
nand UO_52 (O_52,N_2912,N_2982);
and UO_53 (O_53,N_2910,N_2913);
and UO_54 (O_54,N_2918,N_2955);
nand UO_55 (O_55,N_2925,N_2997);
nand UO_56 (O_56,N_2945,N_2907);
nor UO_57 (O_57,N_2920,N_2959);
nor UO_58 (O_58,N_2910,N_2937);
or UO_59 (O_59,N_2989,N_2929);
nand UO_60 (O_60,N_2913,N_2918);
nand UO_61 (O_61,N_2926,N_2911);
nand UO_62 (O_62,N_2911,N_2988);
and UO_63 (O_63,N_2925,N_2972);
and UO_64 (O_64,N_2989,N_2942);
and UO_65 (O_65,N_2916,N_2926);
or UO_66 (O_66,N_2998,N_2983);
and UO_67 (O_67,N_2936,N_2938);
and UO_68 (O_68,N_2966,N_2919);
and UO_69 (O_69,N_2988,N_2915);
nor UO_70 (O_70,N_2921,N_2918);
nand UO_71 (O_71,N_2957,N_2954);
nor UO_72 (O_72,N_2973,N_2969);
or UO_73 (O_73,N_2966,N_2975);
nand UO_74 (O_74,N_2941,N_2983);
nand UO_75 (O_75,N_2970,N_2904);
nor UO_76 (O_76,N_2928,N_2958);
nand UO_77 (O_77,N_2923,N_2909);
nor UO_78 (O_78,N_2905,N_2962);
or UO_79 (O_79,N_2916,N_2981);
and UO_80 (O_80,N_2964,N_2913);
nand UO_81 (O_81,N_2948,N_2937);
xor UO_82 (O_82,N_2949,N_2984);
or UO_83 (O_83,N_2967,N_2980);
and UO_84 (O_84,N_2911,N_2987);
nor UO_85 (O_85,N_2995,N_2953);
or UO_86 (O_86,N_2961,N_2951);
nand UO_87 (O_87,N_2960,N_2935);
nor UO_88 (O_88,N_2909,N_2911);
and UO_89 (O_89,N_2993,N_2952);
or UO_90 (O_90,N_2921,N_2983);
or UO_91 (O_91,N_2950,N_2981);
nand UO_92 (O_92,N_2919,N_2961);
nor UO_93 (O_93,N_2981,N_2955);
nor UO_94 (O_94,N_2996,N_2963);
nor UO_95 (O_95,N_2911,N_2947);
or UO_96 (O_96,N_2999,N_2919);
nand UO_97 (O_97,N_2984,N_2973);
or UO_98 (O_98,N_2933,N_2985);
nand UO_99 (O_99,N_2965,N_2973);
and UO_100 (O_100,N_2959,N_2934);
or UO_101 (O_101,N_2905,N_2983);
nor UO_102 (O_102,N_2990,N_2906);
nor UO_103 (O_103,N_2972,N_2930);
and UO_104 (O_104,N_2981,N_2973);
and UO_105 (O_105,N_2953,N_2970);
nor UO_106 (O_106,N_2970,N_2913);
nand UO_107 (O_107,N_2987,N_2962);
or UO_108 (O_108,N_2938,N_2906);
nor UO_109 (O_109,N_2962,N_2994);
nor UO_110 (O_110,N_2930,N_2961);
nor UO_111 (O_111,N_2916,N_2948);
nor UO_112 (O_112,N_2948,N_2983);
nand UO_113 (O_113,N_2908,N_2910);
nor UO_114 (O_114,N_2975,N_2986);
nor UO_115 (O_115,N_2963,N_2995);
nor UO_116 (O_116,N_2971,N_2968);
or UO_117 (O_117,N_2994,N_2940);
nor UO_118 (O_118,N_2903,N_2911);
nand UO_119 (O_119,N_2906,N_2903);
or UO_120 (O_120,N_2913,N_2936);
or UO_121 (O_121,N_2933,N_2928);
nor UO_122 (O_122,N_2903,N_2967);
or UO_123 (O_123,N_2952,N_2935);
and UO_124 (O_124,N_2946,N_2967);
nand UO_125 (O_125,N_2988,N_2966);
or UO_126 (O_126,N_2997,N_2965);
or UO_127 (O_127,N_2917,N_2982);
and UO_128 (O_128,N_2975,N_2915);
and UO_129 (O_129,N_2917,N_2972);
and UO_130 (O_130,N_2966,N_2985);
or UO_131 (O_131,N_2979,N_2995);
nor UO_132 (O_132,N_2984,N_2953);
nand UO_133 (O_133,N_2916,N_2970);
and UO_134 (O_134,N_2906,N_2908);
or UO_135 (O_135,N_2918,N_2950);
nand UO_136 (O_136,N_2994,N_2910);
nand UO_137 (O_137,N_2958,N_2955);
nor UO_138 (O_138,N_2968,N_2925);
and UO_139 (O_139,N_2926,N_2923);
nand UO_140 (O_140,N_2955,N_2936);
or UO_141 (O_141,N_2942,N_2984);
nand UO_142 (O_142,N_2942,N_2921);
nand UO_143 (O_143,N_2931,N_2949);
nor UO_144 (O_144,N_2959,N_2958);
nor UO_145 (O_145,N_2993,N_2967);
or UO_146 (O_146,N_2963,N_2948);
xor UO_147 (O_147,N_2982,N_2981);
nor UO_148 (O_148,N_2939,N_2982);
nor UO_149 (O_149,N_2968,N_2913);
or UO_150 (O_150,N_2963,N_2983);
and UO_151 (O_151,N_2971,N_2930);
nor UO_152 (O_152,N_2916,N_2961);
nand UO_153 (O_153,N_2942,N_2928);
and UO_154 (O_154,N_2911,N_2994);
nor UO_155 (O_155,N_2910,N_2903);
or UO_156 (O_156,N_2910,N_2965);
and UO_157 (O_157,N_2985,N_2996);
or UO_158 (O_158,N_2993,N_2946);
nor UO_159 (O_159,N_2941,N_2923);
nand UO_160 (O_160,N_2950,N_2973);
and UO_161 (O_161,N_2946,N_2917);
nor UO_162 (O_162,N_2905,N_2931);
nor UO_163 (O_163,N_2942,N_2994);
nand UO_164 (O_164,N_2964,N_2932);
and UO_165 (O_165,N_2991,N_2932);
nor UO_166 (O_166,N_2945,N_2967);
nand UO_167 (O_167,N_2942,N_2974);
nor UO_168 (O_168,N_2977,N_2941);
or UO_169 (O_169,N_2969,N_2906);
nand UO_170 (O_170,N_2996,N_2998);
and UO_171 (O_171,N_2903,N_2954);
nor UO_172 (O_172,N_2901,N_2922);
nand UO_173 (O_173,N_2960,N_2994);
and UO_174 (O_174,N_2971,N_2990);
and UO_175 (O_175,N_2945,N_2970);
nand UO_176 (O_176,N_2926,N_2934);
or UO_177 (O_177,N_2960,N_2977);
nor UO_178 (O_178,N_2940,N_2956);
and UO_179 (O_179,N_2981,N_2930);
nand UO_180 (O_180,N_2944,N_2990);
or UO_181 (O_181,N_2924,N_2999);
and UO_182 (O_182,N_2965,N_2907);
nor UO_183 (O_183,N_2946,N_2900);
and UO_184 (O_184,N_2977,N_2996);
nor UO_185 (O_185,N_2976,N_2913);
nand UO_186 (O_186,N_2997,N_2938);
or UO_187 (O_187,N_2950,N_2929);
nor UO_188 (O_188,N_2966,N_2999);
and UO_189 (O_189,N_2958,N_2979);
nand UO_190 (O_190,N_2942,N_2986);
or UO_191 (O_191,N_2965,N_2963);
and UO_192 (O_192,N_2955,N_2951);
nor UO_193 (O_193,N_2921,N_2937);
or UO_194 (O_194,N_2977,N_2955);
nor UO_195 (O_195,N_2921,N_2900);
nor UO_196 (O_196,N_2986,N_2983);
and UO_197 (O_197,N_2946,N_2991);
or UO_198 (O_198,N_2950,N_2958);
or UO_199 (O_199,N_2912,N_2908);
or UO_200 (O_200,N_2922,N_2935);
and UO_201 (O_201,N_2913,N_2989);
or UO_202 (O_202,N_2946,N_2976);
nand UO_203 (O_203,N_2967,N_2914);
or UO_204 (O_204,N_2924,N_2944);
and UO_205 (O_205,N_2980,N_2937);
and UO_206 (O_206,N_2987,N_2925);
and UO_207 (O_207,N_2985,N_2940);
and UO_208 (O_208,N_2959,N_2975);
nand UO_209 (O_209,N_2986,N_2915);
nor UO_210 (O_210,N_2968,N_2900);
nand UO_211 (O_211,N_2901,N_2918);
nand UO_212 (O_212,N_2987,N_2965);
xnor UO_213 (O_213,N_2993,N_2925);
nand UO_214 (O_214,N_2963,N_2979);
or UO_215 (O_215,N_2902,N_2995);
and UO_216 (O_216,N_2918,N_2936);
nor UO_217 (O_217,N_2945,N_2986);
nand UO_218 (O_218,N_2905,N_2943);
nand UO_219 (O_219,N_2960,N_2996);
or UO_220 (O_220,N_2997,N_2976);
nand UO_221 (O_221,N_2984,N_2910);
and UO_222 (O_222,N_2929,N_2976);
or UO_223 (O_223,N_2942,N_2980);
and UO_224 (O_224,N_2931,N_2922);
or UO_225 (O_225,N_2943,N_2906);
or UO_226 (O_226,N_2961,N_2948);
nor UO_227 (O_227,N_2949,N_2933);
nand UO_228 (O_228,N_2961,N_2924);
or UO_229 (O_229,N_2910,N_2905);
nand UO_230 (O_230,N_2965,N_2958);
and UO_231 (O_231,N_2920,N_2950);
nor UO_232 (O_232,N_2959,N_2950);
nand UO_233 (O_233,N_2986,N_2935);
nor UO_234 (O_234,N_2992,N_2923);
and UO_235 (O_235,N_2995,N_2923);
nor UO_236 (O_236,N_2970,N_2949);
nor UO_237 (O_237,N_2939,N_2911);
nor UO_238 (O_238,N_2911,N_2995);
nor UO_239 (O_239,N_2939,N_2985);
nor UO_240 (O_240,N_2937,N_2930);
or UO_241 (O_241,N_2995,N_2965);
and UO_242 (O_242,N_2979,N_2936);
and UO_243 (O_243,N_2949,N_2973);
and UO_244 (O_244,N_2925,N_2996);
nand UO_245 (O_245,N_2963,N_2931);
nor UO_246 (O_246,N_2996,N_2915);
nor UO_247 (O_247,N_2963,N_2908);
nor UO_248 (O_248,N_2969,N_2996);
and UO_249 (O_249,N_2939,N_2992);
nand UO_250 (O_250,N_2956,N_2967);
nor UO_251 (O_251,N_2992,N_2951);
or UO_252 (O_252,N_2945,N_2998);
or UO_253 (O_253,N_2901,N_2986);
or UO_254 (O_254,N_2920,N_2960);
nand UO_255 (O_255,N_2926,N_2989);
xor UO_256 (O_256,N_2934,N_2916);
or UO_257 (O_257,N_2986,N_2981);
nor UO_258 (O_258,N_2949,N_2928);
or UO_259 (O_259,N_2919,N_2946);
nor UO_260 (O_260,N_2987,N_2904);
nor UO_261 (O_261,N_2900,N_2994);
and UO_262 (O_262,N_2908,N_2970);
nor UO_263 (O_263,N_2925,N_2914);
nand UO_264 (O_264,N_2922,N_2957);
and UO_265 (O_265,N_2962,N_2992);
nand UO_266 (O_266,N_2907,N_2995);
nand UO_267 (O_267,N_2984,N_2994);
and UO_268 (O_268,N_2942,N_2937);
or UO_269 (O_269,N_2972,N_2910);
or UO_270 (O_270,N_2938,N_2983);
nand UO_271 (O_271,N_2953,N_2922);
and UO_272 (O_272,N_2916,N_2985);
or UO_273 (O_273,N_2932,N_2982);
and UO_274 (O_274,N_2916,N_2959);
nor UO_275 (O_275,N_2941,N_2900);
or UO_276 (O_276,N_2986,N_2963);
or UO_277 (O_277,N_2923,N_2920);
or UO_278 (O_278,N_2984,N_2902);
nor UO_279 (O_279,N_2967,N_2971);
nor UO_280 (O_280,N_2926,N_2996);
or UO_281 (O_281,N_2924,N_2933);
nor UO_282 (O_282,N_2923,N_2966);
and UO_283 (O_283,N_2972,N_2911);
nor UO_284 (O_284,N_2908,N_2983);
and UO_285 (O_285,N_2935,N_2964);
nor UO_286 (O_286,N_2958,N_2993);
nand UO_287 (O_287,N_2956,N_2932);
nand UO_288 (O_288,N_2978,N_2999);
or UO_289 (O_289,N_2952,N_2909);
nor UO_290 (O_290,N_2962,N_2969);
or UO_291 (O_291,N_2966,N_2935);
and UO_292 (O_292,N_2923,N_2980);
and UO_293 (O_293,N_2946,N_2908);
nand UO_294 (O_294,N_2925,N_2966);
and UO_295 (O_295,N_2948,N_2953);
nor UO_296 (O_296,N_2949,N_2996);
nor UO_297 (O_297,N_2903,N_2966);
or UO_298 (O_298,N_2954,N_2965);
and UO_299 (O_299,N_2922,N_2992);
nand UO_300 (O_300,N_2951,N_2981);
nor UO_301 (O_301,N_2907,N_2912);
and UO_302 (O_302,N_2935,N_2942);
nor UO_303 (O_303,N_2936,N_2914);
and UO_304 (O_304,N_2931,N_2986);
nand UO_305 (O_305,N_2980,N_2915);
nand UO_306 (O_306,N_2911,N_2922);
nand UO_307 (O_307,N_2909,N_2904);
nor UO_308 (O_308,N_2911,N_2963);
nor UO_309 (O_309,N_2906,N_2992);
or UO_310 (O_310,N_2988,N_2974);
or UO_311 (O_311,N_2904,N_2999);
or UO_312 (O_312,N_2968,N_2944);
and UO_313 (O_313,N_2994,N_2958);
and UO_314 (O_314,N_2988,N_2926);
or UO_315 (O_315,N_2926,N_2985);
and UO_316 (O_316,N_2991,N_2929);
nand UO_317 (O_317,N_2970,N_2940);
nand UO_318 (O_318,N_2907,N_2923);
or UO_319 (O_319,N_2975,N_2958);
or UO_320 (O_320,N_2980,N_2963);
nand UO_321 (O_321,N_2993,N_2919);
nor UO_322 (O_322,N_2988,N_2975);
nand UO_323 (O_323,N_2948,N_2942);
nor UO_324 (O_324,N_2911,N_2927);
nor UO_325 (O_325,N_2982,N_2905);
or UO_326 (O_326,N_2985,N_2956);
and UO_327 (O_327,N_2987,N_2900);
and UO_328 (O_328,N_2969,N_2905);
and UO_329 (O_329,N_2901,N_2970);
nand UO_330 (O_330,N_2935,N_2981);
nand UO_331 (O_331,N_2913,N_2954);
nand UO_332 (O_332,N_2936,N_2929);
nand UO_333 (O_333,N_2979,N_2975);
and UO_334 (O_334,N_2923,N_2902);
nand UO_335 (O_335,N_2999,N_2930);
nand UO_336 (O_336,N_2963,N_2990);
nor UO_337 (O_337,N_2900,N_2924);
and UO_338 (O_338,N_2994,N_2978);
or UO_339 (O_339,N_2977,N_2911);
or UO_340 (O_340,N_2918,N_2978);
and UO_341 (O_341,N_2903,N_2992);
and UO_342 (O_342,N_2920,N_2956);
nor UO_343 (O_343,N_2900,N_2955);
and UO_344 (O_344,N_2992,N_2934);
and UO_345 (O_345,N_2984,N_2914);
and UO_346 (O_346,N_2976,N_2957);
or UO_347 (O_347,N_2993,N_2992);
nand UO_348 (O_348,N_2944,N_2994);
and UO_349 (O_349,N_2986,N_2923);
nor UO_350 (O_350,N_2924,N_2936);
nand UO_351 (O_351,N_2982,N_2979);
nand UO_352 (O_352,N_2936,N_2920);
nor UO_353 (O_353,N_2957,N_2964);
nand UO_354 (O_354,N_2949,N_2995);
nand UO_355 (O_355,N_2965,N_2906);
nand UO_356 (O_356,N_2908,N_2915);
or UO_357 (O_357,N_2919,N_2944);
and UO_358 (O_358,N_2946,N_2944);
nand UO_359 (O_359,N_2986,N_2967);
and UO_360 (O_360,N_2940,N_2972);
nand UO_361 (O_361,N_2948,N_2920);
nor UO_362 (O_362,N_2929,N_2965);
nand UO_363 (O_363,N_2948,N_2976);
or UO_364 (O_364,N_2914,N_2986);
nor UO_365 (O_365,N_2991,N_2944);
nand UO_366 (O_366,N_2934,N_2917);
and UO_367 (O_367,N_2951,N_2931);
or UO_368 (O_368,N_2906,N_2913);
and UO_369 (O_369,N_2915,N_2921);
or UO_370 (O_370,N_2952,N_2939);
nand UO_371 (O_371,N_2955,N_2960);
nor UO_372 (O_372,N_2975,N_2945);
or UO_373 (O_373,N_2967,N_2952);
nand UO_374 (O_374,N_2920,N_2910);
and UO_375 (O_375,N_2946,N_2952);
and UO_376 (O_376,N_2953,N_2918);
or UO_377 (O_377,N_2913,N_2974);
or UO_378 (O_378,N_2932,N_2901);
or UO_379 (O_379,N_2975,N_2929);
xor UO_380 (O_380,N_2993,N_2905);
nand UO_381 (O_381,N_2928,N_2973);
or UO_382 (O_382,N_2915,N_2981);
or UO_383 (O_383,N_2908,N_2913);
nor UO_384 (O_384,N_2954,N_2979);
or UO_385 (O_385,N_2993,N_2910);
and UO_386 (O_386,N_2900,N_2951);
or UO_387 (O_387,N_2972,N_2959);
nand UO_388 (O_388,N_2998,N_2964);
and UO_389 (O_389,N_2966,N_2905);
or UO_390 (O_390,N_2973,N_2985);
and UO_391 (O_391,N_2970,N_2931);
and UO_392 (O_392,N_2951,N_2909);
nand UO_393 (O_393,N_2936,N_2990);
nor UO_394 (O_394,N_2933,N_2982);
and UO_395 (O_395,N_2925,N_2991);
nor UO_396 (O_396,N_2945,N_2994);
nand UO_397 (O_397,N_2959,N_2909);
and UO_398 (O_398,N_2983,N_2920);
or UO_399 (O_399,N_2921,N_2998);
nand UO_400 (O_400,N_2944,N_2975);
nor UO_401 (O_401,N_2925,N_2977);
or UO_402 (O_402,N_2999,N_2957);
nand UO_403 (O_403,N_2908,N_2924);
and UO_404 (O_404,N_2999,N_2992);
nor UO_405 (O_405,N_2945,N_2969);
and UO_406 (O_406,N_2904,N_2989);
or UO_407 (O_407,N_2945,N_2902);
nand UO_408 (O_408,N_2965,N_2966);
nand UO_409 (O_409,N_2963,N_2985);
or UO_410 (O_410,N_2963,N_2956);
nor UO_411 (O_411,N_2981,N_2972);
nand UO_412 (O_412,N_2902,N_2901);
or UO_413 (O_413,N_2936,N_2991);
and UO_414 (O_414,N_2993,N_2991);
nor UO_415 (O_415,N_2959,N_2917);
or UO_416 (O_416,N_2976,N_2935);
or UO_417 (O_417,N_2900,N_2914);
or UO_418 (O_418,N_2988,N_2936);
or UO_419 (O_419,N_2927,N_2926);
or UO_420 (O_420,N_2956,N_2914);
or UO_421 (O_421,N_2978,N_2915);
nand UO_422 (O_422,N_2916,N_2942);
and UO_423 (O_423,N_2918,N_2928);
nand UO_424 (O_424,N_2916,N_2903);
nor UO_425 (O_425,N_2972,N_2914);
nor UO_426 (O_426,N_2992,N_2928);
nand UO_427 (O_427,N_2925,N_2943);
or UO_428 (O_428,N_2962,N_2964);
and UO_429 (O_429,N_2955,N_2948);
nand UO_430 (O_430,N_2993,N_2961);
or UO_431 (O_431,N_2945,N_2993);
nand UO_432 (O_432,N_2988,N_2991);
and UO_433 (O_433,N_2919,N_2994);
nor UO_434 (O_434,N_2907,N_2946);
nand UO_435 (O_435,N_2961,N_2970);
and UO_436 (O_436,N_2912,N_2936);
nand UO_437 (O_437,N_2905,N_2938);
nor UO_438 (O_438,N_2989,N_2915);
or UO_439 (O_439,N_2937,N_2905);
or UO_440 (O_440,N_2960,N_2903);
and UO_441 (O_441,N_2908,N_2916);
and UO_442 (O_442,N_2922,N_2981);
nand UO_443 (O_443,N_2931,N_2936);
nand UO_444 (O_444,N_2927,N_2913);
nand UO_445 (O_445,N_2944,N_2949);
or UO_446 (O_446,N_2976,N_2988);
or UO_447 (O_447,N_2922,N_2909);
and UO_448 (O_448,N_2947,N_2997);
nand UO_449 (O_449,N_2998,N_2941);
and UO_450 (O_450,N_2969,N_2953);
nor UO_451 (O_451,N_2933,N_2911);
nor UO_452 (O_452,N_2959,N_2973);
and UO_453 (O_453,N_2967,N_2932);
and UO_454 (O_454,N_2912,N_2987);
or UO_455 (O_455,N_2994,N_2931);
and UO_456 (O_456,N_2959,N_2904);
or UO_457 (O_457,N_2929,N_2908);
and UO_458 (O_458,N_2968,N_2931);
nor UO_459 (O_459,N_2996,N_2939);
nor UO_460 (O_460,N_2937,N_2958);
or UO_461 (O_461,N_2940,N_2935);
nor UO_462 (O_462,N_2976,N_2911);
nor UO_463 (O_463,N_2954,N_2971);
and UO_464 (O_464,N_2998,N_2938);
and UO_465 (O_465,N_2906,N_2934);
and UO_466 (O_466,N_2914,N_2932);
and UO_467 (O_467,N_2922,N_2942);
and UO_468 (O_468,N_2909,N_2965);
or UO_469 (O_469,N_2991,N_2935);
nor UO_470 (O_470,N_2966,N_2955);
and UO_471 (O_471,N_2953,N_2939);
nand UO_472 (O_472,N_2927,N_2986);
nand UO_473 (O_473,N_2996,N_2991);
and UO_474 (O_474,N_2940,N_2962);
and UO_475 (O_475,N_2933,N_2905);
nand UO_476 (O_476,N_2961,N_2979);
nand UO_477 (O_477,N_2972,N_2993);
or UO_478 (O_478,N_2930,N_2940);
and UO_479 (O_479,N_2974,N_2983);
and UO_480 (O_480,N_2938,N_2954);
nor UO_481 (O_481,N_2970,N_2980);
or UO_482 (O_482,N_2915,N_2927);
nor UO_483 (O_483,N_2950,N_2968);
nand UO_484 (O_484,N_2987,N_2910);
nor UO_485 (O_485,N_2968,N_2958);
or UO_486 (O_486,N_2975,N_2957);
and UO_487 (O_487,N_2930,N_2928);
nand UO_488 (O_488,N_2929,N_2903);
or UO_489 (O_489,N_2984,N_2936);
and UO_490 (O_490,N_2997,N_2951);
nand UO_491 (O_491,N_2927,N_2996);
nand UO_492 (O_492,N_2915,N_2964);
and UO_493 (O_493,N_2916,N_2977);
or UO_494 (O_494,N_2969,N_2975);
and UO_495 (O_495,N_2935,N_2992);
or UO_496 (O_496,N_2932,N_2990);
nand UO_497 (O_497,N_2967,N_2985);
nor UO_498 (O_498,N_2927,N_2969);
nand UO_499 (O_499,N_2980,N_2904);
endmodule