module basic_1000_10000_1500_20_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
xor U0 (N_0,In_294,In_937);
and U1 (N_1,In_703,In_874);
xor U2 (N_2,In_879,In_163);
nand U3 (N_3,In_953,In_389);
and U4 (N_4,In_911,In_566);
nand U5 (N_5,In_268,In_834);
or U6 (N_6,In_319,In_84);
xor U7 (N_7,In_688,In_460);
nor U8 (N_8,In_348,In_423);
nor U9 (N_9,In_510,In_773);
or U10 (N_10,In_624,In_190);
and U11 (N_11,In_941,In_264);
nand U12 (N_12,In_998,In_237);
nor U13 (N_13,In_211,In_44);
nand U14 (N_14,In_945,In_247);
or U15 (N_15,In_584,In_801);
and U16 (N_16,In_298,In_628);
xor U17 (N_17,In_990,In_931);
nand U18 (N_18,In_783,In_743);
and U19 (N_19,In_497,In_305);
and U20 (N_20,In_77,In_607);
nor U21 (N_21,In_713,In_453);
or U22 (N_22,In_704,In_507);
nand U23 (N_23,In_295,In_822);
nor U24 (N_24,In_153,In_860);
nor U25 (N_25,In_936,In_477);
nor U26 (N_26,In_340,In_616);
nand U27 (N_27,In_577,In_666);
xnor U28 (N_28,In_925,In_414);
and U29 (N_29,In_260,In_406);
or U30 (N_30,In_641,In_304);
or U31 (N_31,In_357,In_228);
and U32 (N_32,In_330,In_287);
nand U33 (N_33,In_90,In_642);
xnor U34 (N_34,In_904,In_184);
nor U35 (N_35,In_848,In_473);
or U36 (N_36,In_574,In_645);
xnor U37 (N_37,In_440,In_336);
nor U38 (N_38,In_632,In_189);
xor U39 (N_39,In_684,In_432);
and U40 (N_40,In_402,In_382);
nor U41 (N_41,In_66,In_977);
xnor U42 (N_42,In_138,In_139);
nor U43 (N_43,In_907,In_255);
or U44 (N_44,In_608,In_15);
or U45 (N_45,In_444,In_31);
and U46 (N_46,In_101,In_325);
nor U47 (N_47,In_568,In_621);
or U48 (N_48,In_929,In_697);
xnor U49 (N_49,In_622,In_331);
nor U50 (N_50,In_58,In_209);
xor U51 (N_51,In_226,In_395);
nor U52 (N_52,In_290,In_479);
and U53 (N_53,In_531,In_837);
nand U54 (N_54,In_129,In_286);
nor U55 (N_55,In_698,In_321);
or U56 (N_56,In_564,In_455);
nor U57 (N_57,In_445,In_427);
xor U58 (N_58,In_823,In_639);
and U59 (N_59,In_465,In_814);
nand U60 (N_60,In_441,In_875);
nor U61 (N_61,In_862,In_757);
xor U62 (N_62,In_40,In_905);
nand U63 (N_63,In_384,In_575);
and U64 (N_64,In_85,In_764);
or U65 (N_65,In_393,In_789);
and U66 (N_66,In_722,In_399);
xnor U67 (N_67,In_147,In_779);
and U68 (N_68,In_483,In_988);
nand U69 (N_69,In_508,In_644);
nand U70 (N_70,In_685,In_106);
nor U71 (N_71,In_513,In_748);
or U72 (N_72,In_454,In_191);
or U73 (N_73,In_711,In_766);
xnor U74 (N_74,In_344,In_571);
or U75 (N_75,In_123,In_281);
or U76 (N_76,In_0,In_463);
xor U77 (N_77,In_299,In_475);
nor U78 (N_78,In_989,In_643);
nand U79 (N_79,In_241,In_657);
nand U80 (N_80,In_57,In_912);
xor U81 (N_81,In_485,In_278);
and U82 (N_82,In_864,In_438);
nand U83 (N_83,In_873,In_595);
nand U84 (N_84,In_313,In_366);
nand U85 (N_85,In_638,In_346);
nand U86 (N_86,In_846,In_21);
and U87 (N_87,In_746,In_503);
xnor U88 (N_88,In_60,In_474);
nand U89 (N_89,In_901,In_887);
xor U90 (N_90,In_899,In_649);
nand U91 (N_91,In_322,In_968);
nand U92 (N_92,In_620,In_733);
or U93 (N_93,In_387,In_419);
or U94 (N_94,In_315,In_256);
and U95 (N_95,In_464,In_374);
and U96 (N_96,In_702,In_556);
xor U97 (N_97,In_426,In_650);
nand U98 (N_98,In_248,In_780);
nand U99 (N_99,In_240,In_122);
nor U100 (N_100,In_902,In_200);
nor U101 (N_101,In_108,In_560);
nor U102 (N_102,In_561,In_536);
nor U103 (N_103,In_198,In_527);
and U104 (N_104,In_232,In_30);
and U105 (N_105,In_647,In_415);
or U106 (N_106,In_222,In_665);
or U107 (N_107,In_64,In_553);
or U108 (N_108,In_776,In_699);
or U109 (N_109,In_442,In_431);
nor U110 (N_110,In_859,In_107);
xnor U111 (N_111,In_709,In_732);
or U112 (N_112,In_784,In_932);
nand U113 (N_113,In_367,In_158);
xor U114 (N_114,In_48,In_243);
nor U115 (N_115,In_663,In_750);
nor U116 (N_116,In_920,In_249);
nor U117 (N_117,In_996,In_132);
and U118 (N_118,In_46,In_22);
nand U119 (N_119,In_323,In_917);
or U120 (N_120,In_832,In_514);
xor U121 (N_121,In_809,In_654);
nand U122 (N_122,In_839,In_959);
and U123 (N_123,In_919,In_565);
xnor U124 (N_124,In_457,In_712);
or U125 (N_125,In_962,In_117);
nand U126 (N_126,In_221,In_254);
xor U127 (N_127,In_401,In_80);
or U128 (N_128,In_913,In_715);
nand U129 (N_129,In_597,In_771);
and U130 (N_130,In_334,In_606);
nor U131 (N_131,In_602,In_24);
nor U132 (N_132,In_731,In_522);
nor U133 (N_133,In_615,In_377);
nand U134 (N_134,In_960,In_817);
or U135 (N_135,In_850,In_852);
and U136 (N_136,In_276,In_56);
xor U137 (N_137,In_829,In_429);
and U138 (N_138,In_942,In_300);
or U139 (N_139,In_133,In_686);
xnor U140 (N_140,In_493,In_231);
or U141 (N_141,In_235,In_782);
nand U142 (N_142,In_74,In_131);
nor U143 (N_143,In_705,In_469);
nand U144 (N_144,In_885,In_370);
xnor U145 (N_145,In_926,In_121);
or U146 (N_146,In_633,In_843);
xor U147 (N_147,In_86,In_856);
xor U148 (N_148,In_140,In_659);
or U149 (N_149,In_589,In_634);
nand U150 (N_150,In_542,In_603);
and U151 (N_151,In_605,In_204);
or U152 (N_152,In_283,In_736);
nor U153 (N_153,In_687,In_800);
and U154 (N_154,In_799,In_417);
or U155 (N_155,In_528,In_857);
nand U156 (N_156,In_552,In_26);
nand U157 (N_157,In_328,In_915);
and U158 (N_158,In_17,In_157);
or U159 (N_159,In_179,In_821);
and U160 (N_160,In_950,In_738);
nand U161 (N_161,In_381,In_554);
and U162 (N_162,In_368,In_934);
nor U163 (N_163,In_316,In_866);
or U164 (N_164,In_827,In_38);
nand U165 (N_165,In_103,In_413);
and U166 (N_166,In_892,In_403);
and U167 (N_167,In_626,In_50);
or U168 (N_168,In_270,In_807);
or U169 (N_169,In_535,In_867);
xnor U170 (N_170,In_753,In_233);
xor U171 (N_171,In_742,In_311);
and U172 (N_172,In_45,In_113);
xor U173 (N_173,In_302,In_694);
nor U174 (N_174,In_7,In_193);
or U175 (N_175,In_65,In_420);
nand U176 (N_176,In_187,In_338);
nand U177 (N_177,In_450,In_617);
xnor U178 (N_178,In_98,In_136);
nand U179 (N_179,In_745,In_923);
nand U180 (N_180,In_358,In_559);
xor U181 (N_181,In_635,In_545);
or U182 (N_182,In_886,In_692);
xor U183 (N_183,In_869,In_227);
xor U184 (N_184,In_379,In_109);
nand U185 (N_185,In_79,In_161);
xnor U186 (N_186,In_640,In_218);
xor U187 (N_187,In_562,In_333);
and U188 (N_188,In_672,In_239);
and U189 (N_189,In_760,In_914);
nand U190 (N_190,In_585,In_288);
xnor U191 (N_191,In_747,In_938);
nor U192 (N_192,In_55,In_360);
xnor U193 (N_193,In_115,In_412);
xnor U194 (N_194,In_487,In_482);
or U195 (N_195,In_973,In_655);
or U196 (N_196,In_156,In_196);
xnor U197 (N_197,In_981,In_70);
nor U198 (N_198,In_439,In_97);
or U199 (N_199,In_20,In_598);
nand U200 (N_200,In_754,In_335);
xnor U201 (N_201,In_957,In_73);
and U202 (N_202,In_94,In_159);
or U203 (N_203,In_437,In_434);
xor U204 (N_204,In_588,In_212);
nand U205 (N_205,In_601,In_756);
xor U206 (N_206,In_435,In_296);
and U207 (N_207,In_840,In_262);
and U208 (N_208,In_517,In_490);
or U209 (N_209,In_2,In_930);
xnor U210 (N_210,In_819,In_274);
or U211 (N_211,In_682,In_112);
and U212 (N_212,In_365,In_660);
and U213 (N_213,In_969,In_383);
nand U214 (N_214,In_521,In_266);
or U215 (N_215,In_767,In_261);
or U216 (N_216,In_408,In_975);
nor U217 (N_217,In_125,In_223);
xor U218 (N_218,In_951,In_965);
or U219 (N_219,In_691,In_803);
nand U220 (N_220,In_145,In_735);
or U221 (N_221,In_689,In_794);
nand U222 (N_222,In_897,In_908);
nor U223 (N_223,In_155,In_105);
nand U224 (N_224,In_199,In_708);
nor U225 (N_225,In_349,In_786);
and U226 (N_226,In_549,In_669);
nor U227 (N_227,In_728,In_512);
or U228 (N_228,In_301,In_253);
xor U229 (N_229,In_587,In_967);
nor U230 (N_230,In_308,In_385);
or U231 (N_231,In_41,In_250);
xnor U232 (N_232,In_785,In_197);
xor U233 (N_233,In_206,In_831);
and U234 (N_234,In_798,In_54);
nand U235 (N_235,In_216,In_581);
xor U236 (N_236,In_148,In_592);
or U237 (N_237,In_502,In_933);
or U238 (N_238,In_667,In_416);
nand U239 (N_239,In_543,In_893);
xnor U240 (N_240,In_882,In_623);
nand U241 (N_241,In_579,In_119);
nor U242 (N_242,In_195,In_166);
or U243 (N_243,In_171,In_533);
nand U244 (N_244,In_979,In_976);
and U245 (N_245,In_927,In_854);
nand U246 (N_246,In_356,In_152);
or U247 (N_247,In_394,In_570);
or U248 (N_248,In_982,In_978);
nand U249 (N_249,In_991,In_353);
nand U250 (N_250,In_863,In_948);
nor U251 (N_251,In_214,In_110);
xor U252 (N_252,In_997,In_12);
nand U253 (N_253,In_128,In_371);
nand U254 (N_254,In_940,In_741);
nor U255 (N_255,In_826,In_81);
nor U256 (N_256,In_815,In_208);
or U257 (N_257,In_631,In_878);
nand U258 (N_258,In_397,In_600);
nand U259 (N_259,In_451,In_718);
or U260 (N_260,In_806,In_462);
nor U261 (N_261,In_114,In_398);
nor U262 (N_262,In_309,In_386);
or U263 (N_263,In_966,In_154);
nand U264 (N_264,In_530,In_791);
nand U265 (N_265,In_599,In_185);
or U266 (N_266,In_787,In_245);
xor U267 (N_267,In_749,In_13);
and U268 (N_268,In_781,In_96);
xnor U269 (N_269,In_774,In_519);
or U270 (N_270,In_611,In_267);
or U271 (N_271,In_244,In_345);
xor U272 (N_272,In_47,In_471);
xor U273 (N_273,In_961,In_470);
nor U274 (N_274,In_160,In_14);
nor U275 (N_275,In_636,In_424);
or U276 (N_276,In_486,In_546);
or U277 (N_277,In_271,In_538);
xnor U278 (N_278,In_572,In_25);
and U279 (N_279,In_143,In_721);
xor U280 (N_280,In_795,In_452);
xor U281 (N_281,In_10,In_164);
nor U282 (N_282,In_591,In_376);
and U283 (N_283,In_590,In_99);
nor U284 (N_284,In_762,In_759);
nor U285 (N_285,In_52,In_668);
nand U286 (N_286,In_596,In_625);
xnor U287 (N_287,In_956,In_236);
nand U288 (N_288,In_326,In_207);
and U289 (N_289,In_242,In_884);
nand U290 (N_290,In_284,In_534);
or U291 (N_291,In_529,In_693);
xor U292 (N_292,In_987,In_303);
nand U293 (N_293,In_280,In_11);
nand U294 (N_294,In_312,In_263);
nor U295 (N_295,In_777,In_39);
nand U296 (N_296,In_37,In_355);
nand U297 (N_297,In_855,In_4);
and U298 (N_298,In_496,In_847);
nand U299 (N_299,In_16,In_730);
nor U300 (N_300,In_307,In_29);
nor U301 (N_301,In_540,In_828);
nor U302 (N_302,In_726,In_719);
xnor U303 (N_303,In_364,In_755);
or U304 (N_304,In_944,In_3);
nor U305 (N_305,In_224,In_734);
or U306 (N_306,In_898,In_310);
nor U307 (N_307,In_896,In_964);
nand U308 (N_308,In_468,In_467);
or U309 (N_309,In_405,In_42);
xor U310 (N_310,In_443,In_993);
xor U311 (N_311,In_238,In_142);
and U312 (N_312,In_895,In_230);
and U313 (N_313,In_146,In_740);
or U314 (N_314,In_797,In_49);
xnor U315 (N_315,In_62,In_729);
or U316 (N_316,In_317,In_111);
xor U317 (N_317,In_272,In_448);
or U318 (N_318,In_201,In_396);
or U319 (N_319,In_215,In_182);
and U320 (N_320,In_63,In_82);
nand U321 (N_321,In_717,In_681);
xnor U322 (N_322,In_351,In_943);
nand U323 (N_323,In_835,In_618);
and U324 (N_324,In_935,In_130);
xnor U325 (N_325,In_768,In_812);
nand U326 (N_326,In_980,In_924);
nor U327 (N_327,In_656,In_499);
xor U328 (N_328,In_788,In_576);
nand U329 (N_329,In_770,In_868);
and U330 (N_330,In_76,In_18);
nand U331 (N_331,In_43,In_891);
or U332 (N_332,In_761,In_796);
xor U333 (N_333,In_498,In_375);
nor U334 (N_334,In_362,In_578);
nand U335 (N_335,In_292,In_151);
and U336 (N_336,In_277,In_820);
nand U337 (N_337,In_359,In_752);
nor U338 (N_338,In_583,In_410);
or U339 (N_339,In_739,In_985);
and U340 (N_340,In_104,In_339);
xnor U341 (N_341,In_167,In_174);
and U342 (N_342,In_378,In_72);
and U343 (N_343,In_337,In_352);
nand U344 (N_344,In_994,In_461);
and U345 (N_345,In_524,In_793);
and U346 (N_346,In_293,In_246);
or U347 (N_347,In_888,In_180);
or U348 (N_348,In_818,In_68);
or U349 (N_349,In_509,In_202);
and U350 (N_350,In_217,In_314);
xor U351 (N_351,In_102,In_478);
xnor U352 (N_352,In_404,In_910);
nor U353 (N_353,In_203,In_983);
nand U354 (N_354,In_918,In_342);
nand U355 (N_355,In_78,In_134);
xnor U356 (N_356,In_939,In_594);
and U357 (N_357,In_723,In_995);
xnor U358 (N_358,In_518,In_664);
or U359 (N_359,In_537,In_34);
xnor U360 (N_360,In_33,In_329);
and U361 (N_361,In_548,In_804);
xor U362 (N_362,In_257,In_484);
and U363 (N_363,In_630,In_372);
xnor U364 (N_364,In_551,In_433);
xnor U365 (N_365,In_137,In_289);
or U366 (N_366,In_285,In_544);
nor U367 (N_367,In_674,In_954);
nor U368 (N_368,In_418,In_306);
nand U369 (N_369,In_258,In_838);
xor U370 (N_370,In_168,In_347);
and U371 (N_371,In_83,In_833);
nor U372 (N_372,In_9,In_841);
and U373 (N_373,In_422,In_380);
or U374 (N_374,In_186,In_569);
xor U375 (N_375,In_646,In_150);
or U376 (N_376,In_567,In_523);
nand U377 (N_377,In_350,In_903);
nand U378 (N_378,In_5,In_28);
nor U379 (N_379,In_593,In_890);
nor U380 (N_380,In_547,In_676);
or U381 (N_381,In_495,In_853);
or U382 (N_382,In_273,In_662);
nor U383 (N_383,In_727,In_805);
nor U384 (N_384,In_972,In_19);
and U385 (N_385,In_744,In_671);
xnor U386 (N_386,In_751,In_459);
nand U387 (N_387,In_872,In_71);
nor U388 (N_388,In_558,In_225);
and U389 (N_389,In_341,In_928);
nand U390 (N_390,In_36,In_291);
or U391 (N_391,In_614,In_178);
or U392 (N_392,In_955,In_53);
nand U393 (N_393,In_765,In_844);
nand U394 (N_394,In_458,In_165);
and U395 (N_395,In_706,In_192);
nor U396 (N_396,In_75,In_619);
nand U397 (N_397,In_210,In_332);
nor U398 (N_398,In_170,In_69);
nor U399 (N_399,In_637,In_87);
xor U400 (N_400,In_970,In_586);
nand U401 (N_401,In_627,In_851);
nand U402 (N_402,In_737,In_947);
nor U403 (N_403,In_871,In_532);
and U404 (N_404,In_778,In_842);
nor U405 (N_405,In_61,In_67);
nor U406 (N_406,In_318,In_999);
nor U407 (N_407,In_769,In_836);
and U408 (N_408,In_511,In_390);
nor U409 (N_409,In_648,In_909);
nand U410 (N_410,In_491,In_501);
and U411 (N_411,In_725,In_881);
nand U412 (N_412,In_279,In_849);
nor U413 (N_413,In_506,In_188);
or U414 (N_414,In_696,In_428);
nor U415 (N_415,In_51,In_388);
or U416 (N_416,In_494,In_652);
and U417 (N_417,In_880,In_526);
or U418 (N_418,In_27,In_557);
and U419 (N_419,In_141,In_610);
xnor U420 (N_420,In_758,In_673);
xnor U421 (N_421,In_126,In_612);
nor U422 (N_422,In_775,In_516);
xnor U423 (N_423,In_720,In_6);
nand U424 (N_424,In_1,In_992);
and U425 (N_425,In_275,In_489);
nor U426 (N_426,In_100,In_220);
nor U427 (N_427,In_89,In_714);
or U428 (N_428,In_407,In_555);
or U429 (N_429,In_701,In_824);
or U430 (N_430,In_916,In_525);
or U431 (N_431,In_144,In_700);
and U432 (N_432,In_172,In_361);
nand U433 (N_433,In_481,In_392);
and U434 (N_434,In_845,In_716);
xnor U435 (N_435,In_176,In_124);
xnor U436 (N_436,In_825,In_472);
or U437 (N_437,In_678,In_679);
or U438 (N_438,In_320,In_421);
nand U439 (N_439,In_906,In_447);
nand U440 (N_440,In_282,In_658);
nor U441 (N_441,In_889,In_883);
and U442 (N_442,In_573,In_861);
nand U443 (N_443,In_194,In_476);
or U444 (N_444,In_480,In_870);
nand U445 (N_445,In_369,In_466);
or U446 (N_446,In_974,In_149);
xor U447 (N_447,In_651,In_492);
or U448 (N_448,In_265,In_91);
or U449 (N_449,In_790,In_922);
and U450 (N_450,In_175,In_446);
and U451 (N_451,In_436,In_986);
or U452 (N_452,In_8,In_865);
or U453 (N_453,In_373,In_425);
nor U454 (N_454,In_504,In_604);
nor U455 (N_455,In_116,In_259);
nand U456 (N_456,In_269,In_813);
nor U457 (N_457,In_695,In_792);
nor U458 (N_458,In_670,In_456);
and U459 (N_459,In_580,In_181);
nor U460 (N_460,In_710,In_127);
or U461 (N_461,In_539,In_411);
or U462 (N_462,In_324,In_877);
nor U463 (N_463,In_653,In_858);
and U464 (N_464,In_830,In_120);
nor U465 (N_465,In_680,In_582);
or U466 (N_466,In_449,In_391);
or U467 (N_467,In_500,In_505);
and U468 (N_468,In_88,In_354);
and U469 (N_469,In_430,In_93);
nand U470 (N_470,In_177,In_251);
nor U471 (N_471,In_95,In_675);
or U472 (N_472,In_327,In_609);
or U473 (N_473,In_550,In_297);
nand U474 (N_474,In_724,In_205);
xor U475 (N_475,In_183,In_213);
or U476 (N_476,In_946,In_135);
or U477 (N_477,In_363,In_629);
and U478 (N_478,In_23,In_677);
nand U479 (N_479,In_900,In_162);
xor U480 (N_480,In_219,In_894);
or U481 (N_481,In_707,In_984);
or U482 (N_482,In_763,In_690);
nor U483 (N_483,In_810,In_963);
xor U484 (N_484,In_488,In_59);
nor U485 (N_485,In_541,In_952);
nand U486 (N_486,In_563,In_613);
xor U487 (N_487,In_921,In_816);
nor U488 (N_488,In_169,In_400);
or U489 (N_489,In_520,In_811);
and U490 (N_490,In_876,In_661);
or U491 (N_491,In_234,In_343);
or U492 (N_492,In_971,In_515);
xnor U493 (N_493,In_118,In_802);
xnor U494 (N_494,In_683,In_32);
nand U495 (N_495,In_808,In_252);
nor U496 (N_496,In_949,In_229);
or U497 (N_497,In_173,In_35);
xor U498 (N_498,In_92,In_958);
or U499 (N_499,In_772,In_409);
and U500 (N_500,N_91,N_389);
and U501 (N_501,N_405,N_356);
xnor U502 (N_502,N_298,N_273);
nand U503 (N_503,N_425,N_40);
or U504 (N_504,N_155,N_317);
and U505 (N_505,N_357,N_131);
xor U506 (N_506,N_485,N_351);
nor U507 (N_507,N_461,N_483);
nand U508 (N_508,N_120,N_364);
or U509 (N_509,N_375,N_417);
or U510 (N_510,N_304,N_388);
nand U511 (N_511,N_428,N_161);
and U512 (N_512,N_238,N_419);
nor U513 (N_513,N_194,N_224);
nor U514 (N_514,N_463,N_430);
nor U515 (N_515,N_191,N_151);
xor U516 (N_516,N_133,N_324);
xor U517 (N_517,N_482,N_452);
xor U518 (N_518,N_380,N_29);
nand U519 (N_519,N_175,N_255);
nand U520 (N_520,N_221,N_148);
and U521 (N_521,N_289,N_164);
and U522 (N_522,N_59,N_159);
nor U523 (N_523,N_200,N_81);
nand U524 (N_524,N_270,N_400);
nor U525 (N_525,N_15,N_451);
xor U526 (N_526,N_25,N_19);
nand U527 (N_527,N_440,N_297);
nor U528 (N_528,N_471,N_17);
xor U529 (N_529,N_416,N_193);
xor U530 (N_530,N_113,N_363);
nor U531 (N_531,N_267,N_207);
and U532 (N_532,N_382,N_127);
and U533 (N_533,N_61,N_185);
xor U534 (N_534,N_182,N_147);
xnor U535 (N_535,N_467,N_299);
or U536 (N_536,N_248,N_307);
nor U537 (N_537,N_88,N_287);
and U538 (N_538,N_285,N_160);
nand U539 (N_539,N_208,N_145);
xnor U540 (N_540,N_239,N_42);
or U541 (N_541,N_371,N_404);
nor U542 (N_542,N_46,N_190);
or U543 (N_543,N_432,N_16);
xor U544 (N_544,N_349,N_170);
nand U545 (N_545,N_308,N_309);
nor U546 (N_546,N_453,N_86);
nor U547 (N_547,N_408,N_251);
or U548 (N_548,N_481,N_369);
and U549 (N_549,N_266,N_384);
or U550 (N_550,N_424,N_7);
or U551 (N_551,N_499,N_354);
and U552 (N_552,N_105,N_288);
xnor U553 (N_553,N_275,N_77);
nor U554 (N_554,N_90,N_82);
and U555 (N_555,N_395,N_387);
nand U556 (N_556,N_486,N_296);
nand U557 (N_557,N_262,N_236);
or U558 (N_558,N_187,N_129);
and U559 (N_559,N_427,N_496);
nor U560 (N_560,N_277,N_237);
nor U561 (N_561,N_258,N_123);
xor U562 (N_562,N_246,N_318);
or U563 (N_563,N_128,N_210);
or U564 (N_564,N_286,N_144);
and U565 (N_565,N_319,N_337);
or U566 (N_566,N_150,N_149);
or U567 (N_567,N_274,N_102);
nor U568 (N_568,N_117,N_179);
or U569 (N_569,N_203,N_98);
and U570 (N_570,N_21,N_323);
and U571 (N_571,N_344,N_279);
and U572 (N_572,N_28,N_233);
nand U573 (N_573,N_85,N_80);
xor U574 (N_574,N_60,N_108);
nand U575 (N_575,N_495,N_465);
and U576 (N_576,N_435,N_54);
nor U577 (N_577,N_243,N_249);
and U578 (N_578,N_36,N_83);
nor U579 (N_579,N_184,N_459);
nand U580 (N_580,N_346,N_26);
nand U581 (N_581,N_163,N_263);
and U582 (N_582,N_10,N_392);
or U583 (N_583,N_97,N_413);
xnor U584 (N_584,N_23,N_283);
xnor U585 (N_585,N_366,N_368);
xor U586 (N_586,N_22,N_295);
xnor U587 (N_587,N_256,N_330);
or U588 (N_588,N_429,N_100);
or U589 (N_589,N_409,N_18);
and U590 (N_590,N_312,N_332);
nand U591 (N_591,N_55,N_403);
nand U592 (N_592,N_230,N_104);
nand U593 (N_593,N_301,N_172);
nor U594 (N_594,N_306,N_34);
nor U595 (N_595,N_213,N_245);
and U596 (N_596,N_342,N_347);
nor U597 (N_597,N_303,N_30);
nor U598 (N_598,N_2,N_116);
or U599 (N_599,N_410,N_247);
xnor U600 (N_600,N_444,N_271);
and U601 (N_601,N_242,N_56);
xnor U602 (N_602,N_231,N_462);
nor U603 (N_603,N_69,N_436);
or U604 (N_604,N_215,N_51);
nand U605 (N_605,N_45,N_216);
nor U606 (N_606,N_446,N_195);
nand U607 (N_607,N_438,N_33);
or U608 (N_608,N_268,N_406);
nor U609 (N_609,N_326,N_442);
nor U610 (N_610,N_365,N_196);
nor U611 (N_611,N_95,N_358);
xnor U612 (N_612,N_259,N_367);
nor U613 (N_613,N_139,N_261);
nor U614 (N_614,N_449,N_126);
and U615 (N_615,N_464,N_254);
nand U616 (N_616,N_204,N_205);
nand U617 (N_617,N_362,N_333);
nand U618 (N_618,N_73,N_250);
or U619 (N_619,N_209,N_479);
nor U620 (N_620,N_78,N_186);
and U621 (N_621,N_350,N_386);
or U622 (N_622,N_477,N_99);
and U623 (N_623,N_361,N_206);
and U624 (N_624,N_327,N_52);
and U625 (N_625,N_112,N_293);
nand U626 (N_626,N_378,N_79);
and U627 (N_627,N_89,N_13);
nor U628 (N_628,N_498,N_92);
or U629 (N_629,N_157,N_125);
nand U630 (N_630,N_457,N_93);
xnor U631 (N_631,N_325,N_494);
nand U632 (N_632,N_320,N_39);
or U633 (N_633,N_488,N_192);
xor U634 (N_634,N_158,N_87);
or U635 (N_635,N_136,N_35);
xor U636 (N_636,N_257,N_228);
nor U637 (N_637,N_497,N_244);
and U638 (N_638,N_458,N_162);
or U639 (N_639,N_478,N_314);
xor U640 (N_640,N_402,N_454);
and U641 (N_641,N_252,N_154);
and U642 (N_642,N_171,N_352);
or U643 (N_643,N_422,N_281);
nand U644 (N_644,N_360,N_290);
nor U645 (N_645,N_101,N_441);
or U646 (N_646,N_165,N_343);
nor U647 (N_647,N_241,N_394);
and U648 (N_648,N_493,N_472);
or U649 (N_649,N_188,N_9);
nand U650 (N_650,N_1,N_381);
nor U651 (N_651,N_37,N_146);
nand U652 (N_652,N_311,N_130);
nand U653 (N_653,N_359,N_225);
nand U654 (N_654,N_132,N_466);
or U655 (N_655,N_313,N_14);
or U656 (N_656,N_321,N_393);
and U657 (N_657,N_374,N_302);
nor U658 (N_658,N_44,N_71);
nor U659 (N_659,N_11,N_24);
and U660 (N_660,N_67,N_338);
xor U661 (N_661,N_121,N_212);
nand U662 (N_662,N_235,N_229);
or U663 (N_663,N_201,N_473);
xor U664 (N_664,N_57,N_469);
and U665 (N_665,N_234,N_423);
and U666 (N_666,N_48,N_339);
xnor U667 (N_667,N_345,N_8);
and U668 (N_668,N_41,N_178);
and U669 (N_669,N_468,N_109);
xnor U670 (N_670,N_448,N_110);
and U671 (N_671,N_300,N_174);
nand U672 (N_672,N_43,N_445);
nor U673 (N_673,N_226,N_272);
nor U674 (N_674,N_376,N_334);
or U675 (N_675,N_426,N_32);
and U676 (N_676,N_460,N_167);
and U677 (N_677,N_27,N_421);
xor U678 (N_678,N_218,N_183);
xnor U679 (N_679,N_168,N_3);
nand U680 (N_680,N_118,N_370);
xor U681 (N_681,N_456,N_373);
nand U682 (N_682,N_142,N_198);
nand U683 (N_683,N_401,N_119);
nand U684 (N_684,N_407,N_280);
nand U685 (N_685,N_396,N_140);
nand U686 (N_686,N_138,N_227);
nand U687 (N_687,N_180,N_199);
nand U688 (N_688,N_12,N_222);
nor U689 (N_689,N_348,N_276);
nand U690 (N_690,N_177,N_447);
or U691 (N_691,N_476,N_437);
nand U692 (N_692,N_6,N_336);
xnor U693 (N_693,N_291,N_390);
nor U694 (N_694,N_107,N_372);
nand U695 (N_695,N_265,N_64);
xnor U696 (N_696,N_106,N_63);
nand U697 (N_697,N_124,N_260);
nor U698 (N_698,N_399,N_315);
nand U699 (N_699,N_156,N_487);
nor U700 (N_700,N_450,N_316);
nand U701 (N_701,N_31,N_340);
nand U702 (N_702,N_341,N_96);
xnor U703 (N_703,N_103,N_53);
or U704 (N_704,N_489,N_115);
nor U705 (N_705,N_49,N_68);
nor U706 (N_706,N_418,N_217);
nor U707 (N_707,N_282,N_50);
and U708 (N_708,N_111,N_253);
and U709 (N_709,N_211,N_329);
nor U710 (N_710,N_66,N_202);
nor U711 (N_711,N_398,N_411);
nor U712 (N_712,N_433,N_443);
and U713 (N_713,N_70,N_474);
nand U714 (N_714,N_62,N_264);
and U715 (N_715,N_292,N_122);
xnor U716 (N_716,N_38,N_377);
nor U717 (N_717,N_72,N_47);
or U718 (N_718,N_434,N_135);
nor U719 (N_719,N_322,N_84);
xnor U720 (N_720,N_328,N_137);
nand U721 (N_721,N_491,N_153);
nand U722 (N_722,N_232,N_197);
nor U723 (N_723,N_415,N_490);
nor U724 (N_724,N_412,N_220);
and U725 (N_725,N_74,N_5);
and U726 (N_726,N_141,N_214);
xnor U727 (N_727,N_152,N_414);
or U728 (N_728,N_470,N_475);
nor U729 (N_729,N_76,N_94);
nor U730 (N_730,N_114,N_173);
nand U731 (N_731,N_166,N_189);
or U732 (N_732,N_492,N_391);
or U733 (N_733,N_65,N_480);
or U734 (N_734,N_379,N_284);
xor U735 (N_735,N_331,N_439);
xnor U736 (N_736,N_305,N_455);
and U737 (N_737,N_169,N_240);
or U738 (N_738,N_397,N_294);
nor U739 (N_739,N_310,N_4);
and U740 (N_740,N_219,N_335);
nor U741 (N_741,N_383,N_269);
nand U742 (N_742,N_58,N_0);
nor U743 (N_743,N_223,N_181);
or U744 (N_744,N_484,N_278);
or U745 (N_745,N_134,N_385);
nand U746 (N_746,N_353,N_20);
or U747 (N_747,N_355,N_431);
or U748 (N_748,N_143,N_420);
xor U749 (N_749,N_176,N_75);
nor U750 (N_750,N_323,N_334);
or U751 (N_751,N_86,N_398);
xnor U752 (N_752,N_214,N_51);
and U753 (N_753,N_496,N_351);
xnor U754 (N_754,N_174,N_176);
xnor U755 (N_755,N_12,N_118);
or U756 (N_756,N_406,N_486);
nand U757 (N_757,N_213,N_60);
nand U758 (N_758,N_210,N_468);
xor U759 (N_759,N_392,N_165);
or U760 (N_760,N_303,N_67);
or U761 (N_761,N_82,N_194);
or U762 (N_762,N_493,N_289);
and U763 (N_763,N_313,N_213);
nor U764 (N_764,N_97,N_64);
xor U765 (N_765,N_400,N_123);
xor U766 (N_766,N_63,N_283);
nand U767 (N_767,N_229,N_450);
nor U768 (N_768,N_336,N_182);
nor U769 (N_769,N_320,N_143);
nor U770 (N_770,N_413,N_132);
xnor U771 (N_771,N_342,N_148);
and U772 (N_772,N_452,N_469);
nor U773 (N_773,N_54,N_270);
xnor U774 (N_774,N_258,N_482);
or U775 (N_775,N_177,N_239);
xor U776 (N_776,N_21,N_243);
nor U777 (N_777,N_58,N_426);
nor U778 (N_778,N_351,N_120);
or U779 (N_779,N_256,N_93);
and U780 (N_780,N_184,N_231);
xnor U781 (N_781,N_133,N_22);
or U782 (N_782,N_442,N_126);
nand U783 (N_783,N_47,N_488);
or U784 (N_784,N_64,N_145);
and U785 (N_785,N_181,N_431);
and U786 (N_786,N_219,N_175);
or U787 (N_787,N_365,N_86);
nor U788 (N_788,N_170,N_488);
xnor U789 (N_789,N_267,N_170);
or U790 (N_790,N_237,N_195);
nand U791 (N_791,N_468,N_94);
xnor U792 (N_792,N_301,N_71);
xnor U793 (N_793,N_176,N_483);
and U794 (N_794,N_14,N_225);
xor U795 (N_795,N_273,N_418);
and U796 (N_796,N_331,N_252);
xor U797 (N_797,N_471,N_60);
or U798 (N_798,N_274,N_434);
or U799 (N_799,N_365,N_124);
and U800 (N_800,N_118,N_381);
nor U801 (N_801,N_275,N_374);
nor U802 (N_802,N_432,N_81);
xnor U803 (N_803,N_322,N_17);
xor U804 (N_804,N_278,N_472);
xnor U805 (N_805,N_264,N_10);
nand U806 (N_806,N_433,N_246);
or U807 (N_807,N_380,N_362);
xnor U808 (N_808,N_230,N_157);
nand U809 (N_809,N_248,N_176);
nand U810 (N_810,N_277,N_128);
nor U811 (N_811,N_200,N_134);
or U812 (N_812,N_259,N_113);
nor U813 (N_813,N_292,N_118);
or U814 (N_814,N_109,N_168);
xnor U815 (N_815,N_191,N_168);
and U816 (N_816,N_278,N_80);
or U817 (N_817,N_53,N_253);
xnor U818 (N_818,N_300,N_201);
or U819 (N_819,N_243,N_154);
or U820 (N_820,N_128,N_281);
and U821 (N_821,N_277,N_304);
or U822 (N_822,N_64,N_469);
and U823 (N_823,N_425,N_485);
nand U824 (N_824,N_419,N_460);
xnor U825 (N_825,N_110,N_166);
or U826 (N_826,N_243,N_5);
and U827 (N_827,N_39,N_446);
or U828 (N_828,N_95,N_446);
and U829 (N_829,N_216,N_327);
nand U830 (N_830,N_419,N_399);
nor U831 (N_831,N_255,N_497);
xor U832 (N_832,N_437,N_332);
and U833 (N_833,N_253,N_278);
and U834 (N_834,N_242,N_27);
nand U835 (N_835,N_406,N_452);
xor U836 (N_836,N_41,N_405);
and U837 (N_837,N_352,N_433);
and U838 (N_838,N_215,N_27);
xnor U839 (N_839,N_317,N_481);
nor U840 (N_840,N_107,N_467);
and U841 (N_841,N_174,N_349);
or U842 (N_842,N_185,N_178);
nor U843 (N_843,N_477,N_488);
nor U844 (N_844,N_368,N_2);
nor U845 (N_845,N_485,N_444);
and U846 (N_846,N_345,N_375);
nor U847 (N_847,N_484,N_197);
and U848 (N_848,N_288,N_364);
and U849 (N_849,N_434,N_104);
or U850 (N_850,N_314,N_313);
xnor U851 (N_851,N_324,N_168);
and U852 (N_852,N_286,N_142);
nor U853 (N_853,N_287,N_466);
nand U854 (N_854,N_115,N_364);
nand U855 (N_855,N_19,N_68);
nand U856 (N_856,N_371,N_158);
and U857 (N_857,N_319,N_153);
xnor U858 (N_858,N_241,N_285);
nor U859 (N_859,N_123,N_82);
and U860 (N_860,N_351,N_33);
or U861 (N_861,N_219,N_163);
and U862 (N_862,N_41,N_227);
or U863 (N_863,N_153,N_106);
nand U864 (N_864,N_94,N_8);
xnor U865 (N_865,N_313,N_367);
and U866 (N_866,N_67,N_64);
and U867 (N_867,N_363,N_6);
xnor U868 (N_868,N_371,N_40);
and U869 (N_869,N_148,N_23);
nor U870 (N_870,N_173,N_152);
nor U871 (N_871,N_325,N_59);
xor U872 (N_872,N_346,N_462);
nor U873 (N_873,N_84,N_297);
or U874 (N_874,N_226,N_460);
nor U875 (N_875,N_326,N_161);
xnor U876 (N_876,N_256,N_472);
or U877 (N_877,N_198,N_497);
or U878 (N_878,N_262,N_96);
xnor U879 (N_879,N_94,N_75);
or U880 (N_880,N_285,N_257);
xor U881 (N_881,N_348,N_293);
or U882 (N_882,N_176,N_430);
and U883 (N_883,N_47,N_25);
nor U884 (N_884,N_468,N_313);
nor U885 (N_885,N_476,N_327);
xnor U886 (N_886,N_419,N_341);
or U887 (N_887,N_485,N_335);
xor U888 (N_888,N_316,N_391);
nor U889 (N_889,N_324,N_255);
nor U890 (N_890,N_261,N_205);
xor U891 (N_891,N_94,N_220);
or U892 (N_892,N_347,N_203);
and U893 (N_893,N_202,N_162);
and U894 (N_894,N_479,N_214);
and U895 (N_895,N_81,N_470);
or U896 (N_896,N_152,N_30);
xnor U897 (N_897,N_294,N_82);
or U898 (N_898,N_438,N_207);
nand U899 (N_899,N_96,N_278);
or U900 (N_900,N_350,N_275);
and U901 (N_901,N_45,N_103);
or U902 (N_902,N_302,N_43);
and U903 (N_903,N_249,N_311);
nand U904 (N_904,N_380,N_402);
xnor U905 (N_905,N_133,N_360);
xor U906 (N_906,N_421,N_66);
nand U907 (N_907,N_279,N_213);
or U908 (N_908,N_368,N_265);
nand U909 (N_909,N_151,N_43);
or U910 (N_910,N_68,N_175);
nor U911 (N_911,N_151,N_93);
and U912 (N_912,N_157,N_249);
nor U913 (N_913,N_440,N_268);
and U914 (N_914,N_235,N_351);
or U915 (N_915,N_187,N_379);
nand U916 (N_916,N_219,N_73);
nor U917 (N_917,N_339,N_86);
xnor U918 (N_918,N_403,N_476);
nor U919 (N_919,N_469,N_363);
nand U920 (N_920,N_163,N_307);
nand U921 (N_921,N_19,N_93);
and U922 (N_922,N_133,N_450);
nand U923 (N_923,N_206,N_9);
nand U924 (N_924,N_143,N_86);
xnor U925 (N_925,N_43,N_157);
nor U926 (N_926,N_265,N_58);
or U927 (N_927,N_396,N_384);
xnor U928 (N_928,N_489,N_330);
or U929 (N_929,N_373,N_236);
nand U930 (N_930,N_399,N_417);
or U931 (N_931,N_309,N_69);
or U932 (N_932,N_319,N_321);
and U933 (N_933,N_129,N_218);
or U934 (N_934,N_178,N_104);
xnor U935 (N_935,N_311,N_284);
nor U936 (N_936,N_308,N_210);
xor U937 (N_937,N_145,N_315);
nand U938 (N_938,N_46,N_499);
and U939 (N_939,N_141,N_3);
xnor U940 (N_940,N_209,N_415);
nor U941 (N_941,N_351,N_408);
xnor U942 (N_942,N_100,N_472);
nor U943 (N_943,N_410,N_281);
nor U944 (N_944,N_30,N_313);
xor U945 (N_945,N_422,N_69);
or U946 (N_946,N_29,N_478);
nor U947 (N_947,N_285,N_128);
xnor U948 (N_948,N_111,N_225);
xnor U949 (N_949,N_368,N_162);
nor U950 (N_950,N_448,N_248);
xnor U951 (N_951,N_432,N_249);
or U952 (N_952,N_209,N_491);
xor U953 (N_953,N_115,N_259);
and U954 (N_954,N_430,N_226);
nor U955 (N_955,N_373,N_218);
and U956 (N_956,N_387,N_114);
xor U957 (N_957,N_493,N_15);
and U958 (N_958,N_92,N_448);
nor U959 (N_959,N_91,N_223);
and U960 (N_960,N_114,N_17);
and U961 (N_961,N_432,N_342);
and U962 (N_962,N_142,N_365);
and U963 (N_963,N_311,N_14);
nand U964 (N_964,N_299,N_75);
nand U965 (N_965,N_344,N_165);
and U966 (N_966,N_77,N_180);
or U967 (N_967,N_413,N_37);
nand U968 (N_968,N_143,N_90);
xor U969 (N_969,N_250,N_413);
and U970 (N_970,N_324,N_394);
nor U971 (N_971,N_403,N_144);
or U972 (N_972,N_321,N_249);
and U973 (N_973,N_247,N_412);
nand U974 (N_974,N_2,N_233);
and U975 (N_975,N_248,N_153);
nor U976 (N_976,N_409,N_211);
and U977 (N_977,N_6,N_231);
nand U978 (N_978,N_74,N_273);
or U979 (N_979,N_14,N_282);
nand U980 (N_980,N_284,N_481);
xnor U981 (N_981,N_469,N_89);
or U982 (N_982,N_175,N_377);
and U983 (N_983,N_195,N_162);
nor U984 (N_984,N_451,N_156);
or U985 (N_985,N_104,N_158);
or U986 (N_986,N_135,N_255);
and U987 (N_987,N_371,N_122);
nand U988 (N_988,N_271,N_337);
nand U989 (N_989,N_485,N_0);
xor U990 (N_990,N_332,N_122);
or U991 (N_991,N_374,N_414);
xor U992 (N_992,N_328,N_385);
nor U993 (N_993,N_364,N_52);
or U994 (N_994,N_434,N_158);
and U995 (N_995,N_66,N_45);
or U996 (N_996,N_228,N_379);
nand U997 (N_997,N_63,N_56);
and U998 (N_998,N_14,N_262);
and U999 (N_999,N_263,N_0);
or U1000 (N_1000,N_534,N_942);
nand U1001 (N_1001,N_711,N_606);
nand U1002 (N_1002,N_652,N_974);
nor U1003 (N_1003,N_776,N_687);
and U1004 (N_1004,N_768,N_596);
nor U1005 (N_1005,N_678,N_516);
or U1006 (N_1006,N_803,N_869);
xor U1007 (N_1007,N_787,N_580);
nor U1008 (N_1008,N_985,N_524);
or U1009 (N_1009,N_877,N_635);
nand U1010 (N_1010,N_912,N_639);
nand U1011 (N_1011,N_710,N_892);
or U1012 (N_1012,N_653,N_626);
and U1013 (N_1013,N_781,N_889);
nand U1014 (N_1014,N_778,N_631);
or U1015 (N_1015,N_574,N_988);
and U1016 (N_1016,N_713,N_663);
nand U1017 (N_1017,N_566,N_940);
nor U1018 (N_1018,N_730,N_794);
or U1019 (N_1019,N_885,N_982);
and U1020 (N_1020,N_608,N_856);
nand U1021 (N_1021,N_640,N_643);
or U1022 (N_1022,N_503,N_792);
xor U1023 (N_1023,N_948,N_757);
and U1024 (N_1024,N_604,N_677);
and U1025 (N_1025,N_984,N_804);
nand U1026 (N_1026,N_660,N_509);
or U1027 (N_1027,N_665,N_676);
nor U1028 (N_1028,N_759,N_650);
and U1029 (N_1029,N_707,N_598);
xor U1030 (N_1030,N_599,N_949);
and U1031 (N_1031,N_783,N_797);
nand U1032 (N_1032,N_751,N_893);
and U1033 (N_1033,N_884,N_709);
xnor U1034 (N_1034,N_541,N_867);
or U1035 (N_1035,N_934,N_664);
or U1036 (N_1036,N_573,N_789);
and U1037 (N_1037,N_531,N_915);
or U1038 (N_1038,N_829,N_822);
nor U1039 (N_1039,N_696,N_763);
nand U1040 (N_1040,N_718,N_769);
or U1041 (N_1041,N_507,N_513);
or U1042 (N_1042,N_966,N_960);
or U1043 (N_1043,N_755,N_998);
nand U1044 (N_1044,N_540,N_762);
nand U1045 (N_1045,N_786,N_584);
and U1046 (N_1046,N_932,N_758);
nor U1047 (N_1047,N_728,N_590);
and U1048 (N_1048,N_914,N_878);
nand U1049 (N_1049,N_920,N_801);
nor U1050 (N_1050,N_629,N_883);
and U1051 (N_1051,N_815,N_777);
or U1052 (N_1052,N_656,N_539);
nor U1053 (N_1053,N_902,N_634);
nand U1054 (N_1054,N_968,N_738);
xor U1055 (N_1055,N_575,N_649);
nor U1056 (N_1056,N_957,N_847);
xnor U1057 (N_1057,N_838,N_805);
and U1058 (N_1058,N_866,N_908);
nor U1059 (N_1059,N_522,N_773);
nor U1060 (N_1060,N_938,N_673);
nand U1061 (N_1061,N_705,N_567);
or U1062 (N_1062,N_833,N_546);
and U1063 (N_1063,N_700,N_973);
nor U1064 (N_1064,N_782,N_548);
nor U1065 (N_1065,N_645,N_824);
xor U1066 (N_1066,N_670,N_625);
xor U1067 (N_1067,N_875,N_736);
and U1068 (N_1068,N_680,N_962);
nand U1069 (N_1069,N_981,N_734);
nand U1070 (N_1070,N_505,N_809);
or U1071 (N_1071,N_860,N_658);
nand U1072 (N_1072,N_870,N_853);
nand U1073 (N_1073,N_514,N_836);
nand U1074 (N_1074,N_578,N_935);
nand U1075 (N_1075,N_615,N_894);
or U1076 (N_1076,N_739,N_717);
or U1077 (N_1077,N_544,N_963);
nand U1078 (N_1078,N_504,N_729);
nor U1079 (N_1079,N_770,N_852);
nand U1080 (N_1080,N_810,N_979);
xnor U1081 (N_1081,N_909,N_535);
nor U1082 (N_1082,N_901,N_565);
or U1083 (N_1083,N_771,N_987);
and U1084 (N_1084,N_951,N_719);
and U1085 (N_1085,N_742,N_550);
and U1086 (N_1086,N_986,N_701);
or U1087 (N_1087,N_931,N_947);
nor U1088 (N_1088,N_841,N_882);
nor U1089 (N_1089,N_927,N_807);
or U1090 (N_1090,N_814,N_501);
and U1091 (N_1091,N_821,N_843);
or U1092 (N_1092,N_732,N_679);
xor U1093 (N_1093,N_582,N_648);
and U1094 (N_1094,N_971,N_588);
nor U1095 (N_1095,N_695,N_594);
nor U1096 (N_1096,N_846,N_502);
xor U1097 (N_1097,N_785,N_952);
nor U1098 (N_1098,N_965,N_720);
nand U1099 (N_1099,N_969,N_537);
nand U1100 (N_1100,N_826,N_560);
or U1101 (N_1101,N_918,N_623);
and U1102 (N_1102,N_570,N_610);
xnor U1103 (N_1103,N_989,N_585);
or U1104 (N_1104,N_735,N_970);
nor U1105 (N_1105,N_808,N_800);
xnor U1106 (N_1106,N_558,N_572);
or U1107 (N_1107,N_812,N_609);
xor U1108 (N_1108,N_708,N_681);
nor U1109 (N_1109,N_529,N_992);
xnor U1110 (N_1110,N_896,N_749);
nand U1111 (N_1111,N_830,N_748);
xor U1112 (N_1112,N_933,N_586);
xnor U1113 (N_1113,N_863,N_555);
or U1114 (N_1114,N_684,N_876);
and U1115 (N_1115,N_691,N_930);
and U1116 (N_1116,N_618,N_557);
nand U1117 (N_1117,N_593,N_724);
xnor U1118 (N_1118,N_500,N_521);
xnor U1119 (N_1119,N_644,N_581);
nor U1120 (N_1120,N_811,N_577);
nand U1121 (N_1121,N_905,N_651);
nor U1122 (N_1122,N_628,N_512);
xor U1123 (N_1123,N_904,N_697);
and U1124 (N_1124,N_997,N_611);
or U1125 (N_1125,N_520,N_726);
nand U1126 (N_1126,N_667,N_858);
or U1127 (N_1127,N_690,N_636);
xor U1128 (N_1128,N_674,N_552);
xnor U1129 (N_1129,N_793,N_890);
xnor U1130 (N_1130,N_672,N_551);
xor U1131 (N_1131,N_756,N_953);
nand U1132 (N_1132,N_819,N_659);
nand U1133 (N_1133,N_706,N_842);
xnor U1134 (N_1134,N_929,N_950);
or U1135 (N_1135,N_845,N_903);
nor U1136 (N_1136,N_996,N_620);
xor U1137 (N_1137,N_641,N_775);
nor U1138 (N_1138,N_703,N_579);
or U1139 (N_1139,N_595,N_871);
or U1140 (N_1140,N_817,N_831);
nand U1141 (N_1141,N_796,N_741);
or U1142 (N_1142,N_798,N_693);
xor U1143 (N_1143,N_954,N_995);
xor U1144 (N_1144,N_937,N_622);
or U1145 (N_1145,N_760,N_848);
and U1146 (N_1146,N_964,N_538);
nor U1147 (N_1147,N_559,N_666);
nand U1148 (N_1148,N_563,N_941);
or U1149 (N_1149,N_916,N_511);
nand U1150 (N_1150,N_880,N_857);
xnor U1151 (N_1151,N_621,N_823);
and U1152 (N_1152,N_784,N_632);
or U1153 (N_1153,N_955,N_849);
xnor U1154 (N_1154,N_617,N_881);
or U1155 (N_1155,N_515,N_865);
and U1156 (N_1156,N_692,N_619);
nor U1157 (N_1157,N_961,N_510);
or U1158 (N_1158,N_714,N_767);
nand U1159 (N_1159,N_806,N_688);
xnor U1160 (N_1160,N_872,N_716);
nand U1161 (N_1161,N_980,N_698);
and U1162 (N_1162,N_939,N_723);
nand U1163 (N_1163,N_855,N_655);
nand U1164 (N_1164,N_879,N_603);
nand U1165 (N_1165,N_589,N_788);
xnor U1166 (N_1166,N_922,N_820);
nor U1167 (N_1167,N_854,N_910);
and U1168 (N_1168,N_576,N_545);
nand U1169 (N_1169,N_859,N_633);
nor U1170 (N_1170,N_600,N_850);
and U1171 (N_1171,N_840,N_704);
xnor U1172 (N_1172,N_747,N_553);
or U1173 (N_1173,N_668,N_991);
xor U1174 (N_1174,N_977,N_592);
or U1175 (N_1175,N_921,N_740);
xor U1176 (N_1176,N_669,N_612);
xor U1177 (N_1177,N_518,N_627);
nor U1178 (N_1178,N_616,N_542);
nor U1179 (N_1179,N_924,N_946);
and U1180 (N_1180,N_897,N_891);
or U1181 (N_1181,N_699,N_795);
and U1182 (N_1182,N_779,N_813);
xor U1183 (N_1183,N_862,N_834);
and U1184 (N_1184,N_630,N_899);
and U1185 (N_1185,N_959,N_868);
and U1186 (N_1186,N_554,N_683);
and U1187 (N_1187,N_525,N_752);
and U1188 (N_1188,N_682,N_712);
and U1189 (N_1189,N_564,N_765);
or U1190 (N_1190,N_568,N_675);
and U1191 (N_1191,N_972,N_825);
nand U1192 (N_1192,N_907,N_888);
nor U1193 (N_1193,N_647,N_591);
or U1194 (N_1194,N_605,N_967);
or U1195 (N_1195,N_999,N_895);
nor U1196 (N_1196,N_835,N_753);
nor U1197 (N_1197,N_642,N_956);
or U1198 (N_1198,N_519,N_827);
and U1199 (N_1199,N_983,N_750);
or U1200 (N_1200,N_597,N_958);
and U1201 (N_1201,N_613,N_527);
xor U1202 (N_1202,N_780,N_837);
xor U1203 (N_1203,N_828,N_913);
xor U1204 (N_1204,N_614,N_994);
xor U1205 (N_1205,N_601,N_976);
nor U1206 (N_1206,N_900,N_602);
nand U1207 (N_1207,N_873,N_764);
and U1208 (N_1208,N_790,N_844);
nor U1209 (N_1209,N_689,N_911);
nand U1210 (N_1210,N_654,N_766);
nor U1211 (N_1211,N_945,N_936);
and U1212 (N_1212,N_919,N_925);
and U1213 (N_1213,N_508,N_832);
nor U1214 (N_1214,N_562,N_506);
xor U1215 (N_1215,N_536,N_923);
or U1216 (N_1216,N_928,N_721);
xnor U1217 (N_1217,N_737,N_887);
or U1218 (N_1218,N_526,N_607);
xnor U1219 (N_1219,N_772,N_532);
or U1220 (N_1220,N_523,N_637);
xnor U1221 (N_1221,N_851,N_561);
or U1222 (N_1222,N_906,N_799);
nor U1223 (N_1223,N_746,N_733);
and U1224 (N_1224,N_556,N_990);
nand U1225 (N_1225,N_774,N_818);
and U1226 (N_1226,N_543,N_926);
or U1227 (N_1227,N_685,N_569);
nand U1228 (N_1228,N_694,N_743);
nand U1229 (N_1229,N_646,N_686);
nand U1230 (N_1230,N_861,N_583);
xnor U1231 (N_1231,N_917,N_662);
or U1232 (N_1232,N_731,N_874);
or U1233 (N_1233,N_993,N_715);
xnor U1234 (N_1234,N_528,N_886);
nand U1235 (N_1235,N_671,N_549);
nor U1236 (N_1236,N_745,N_638);
xor U1237 (N_1237,N_744,N_761);
nand U1238 (N_1238,N_754,N_943);
xor U1239 (N_1239,N_533,N_587);
xor U1240 (N_1240,N_944,N_547);
nand U1241 (N_1241,N_661,N_816);
nor U1242 (N_1242,N_839,N_727);
xnor U1243 (N_1243,N_725,N_571);
nor U1244 (N_1244,N_975,N_517);
xnor U1245 (N_1245,N_624,N_791);
nor U1246 (N_1246,N_978,N_702);
nor U1247 (N_1247,N_802,N_898);
nand U1248 (N_1248,N_864,N_722);
and U1249 (N_1249,N_530,N_657);
and U1250 (N_1250,N_747,N_956);
xnor U1251 (N_1251,N_519,N_987);
nor U1252 (N_1252,N_892,N_779);
or U1253 (N_1253,N_957,N_703);
xor U1254 (N_1254,N_905,N_754);
nand U1255 (N_1255,N_513,N_876);
and U1256 (N_1256,N_650,N_960);
and U1257 (N_1257,N_645,N_687);
and U1258 (N_1258,N_605,N_839);
or U1259 (N_1259,N_757,N_975);
and U1260 (N_1260,N_849,N_798);
xor U1261 (N_1261,N_913,N_841);
xor U1262 (N_1262,N_689,N_646);
and U1263 (N_1263,N_734,N_945);
or U1264 (N_1264,N_940,N_504);
nand U1265 (N_1265,N_938,N_811);
and U1266 (N_1266,N_950,N_902);
or U1267 (N_1267,N_725,N_946);
xnor U1268 (N_1268,N_959,N_966);
and U1269 (N_1269,N_904,N_882);
or U1270 (N_1270,N_870,N_685);
nor U1271 (N_1271,N_769,N_738);
and U1272 (N_1272,N_702,N_937);
nand U1273 (N_1273,N_563,N_710);
and U1274 (N_1274,N_762,N_856);
nand U1275 (N_1275,N_523,N_629);
and U1276 (N_1276,N_839,N_972);
nand U1277 (N_1277,N_989,N_890);
xnor U1278 (N_1278,N_740,N_680);
nand U1279 (N_1279,N_648,N_653);
xor U1280 (N_1280,N_781,N_610);
nor U1281 (N_1281,N_823,N_862);
xnor U1282 (N_1282,N_610,N_953);
xnor U1283 (N_1283,N_568,N_896);
nor U1284 (N_1284,N_617,N_816);
nor U1285 (N_1285,N_877,N_894);
and U1286 (N_1286,N_979,N_544);
or U1287 (N_1287,N_707,N_860);
or U1288 (N_1288,N_500,N_962);
xnor U1289 (N_1289,N_611,N_694);
and U1290 (N_1290,N_618,N_944);
or U1291 (N_1291,N_869,N_728);
and U1292 (N_1292,N_908,N_666);
xor U1293 (N_1293,N_880,N_580);
or U1294 (N_1294,N_569,N_718);
or U1295 (N_1295,N_848,N_734);
nor U1296 (N_1296,N_563,N_547);
or U1297 (N_1297,N_932,N_987);
nor U1298 (N_1298,N_992,N_629);
nand U1299 (N_1299,N_516,N_743);
xnor U1300 (N_1300,N_950,N_755);
or U1301 (N_1301,N_588,N_512);
or U1302 (N_1302,N_809,N_805);
nor U1303 (N_1303,N_726,N_605);
nor U1304 (N_1304,N_905,N_642);
nand U1305 (N_1305,N_966,N_870);
xnor U1306 (N_1306,N_652,N_715);
nand U1307 (N_1307,N_539,N_511);
and U1308 (N_1308,N_605,N_806);
and U1309 (N_1309,N_712,N_578);
and U1310 (N_1310,N_826,N_647);
and U1311 (N_1311,N_762,N_546);
nor U1312 (N_1312,N_895,N_529);
or U1313 (N_1313,N_815,N_939);
xor U1314 (N_1314,N_608,N_801);
nor U1315 (N_1315,N_924,N_736);
xnor U1316 (N_1316,N_563,N_606);
xor U1317 (N_1317,N_694,N_830);
nand U1318 (N_1318,N_999,N_537);
nor U1319 (N_1319,N_709,N_768);
nor U1320 (N_1320,N_875,N_614);
or U1321 (N_1321,N_633,N_949);
nor U1322 (N_1322,N_976,N_825);
or U1323 (N_1323,N_581,N_548);
and U1324 (N_1324,N_862,N_968);
and U1325 (N_1325,N_808,N_824);
nand U1326 (N_1326,N_760,N_930);
or U1327 (N_1327,N_890,N_560);
nand U1328 (N_1328,N_550,N_954);
and U1329 (N_1329,N_715,N_987);
nand U1330 (N_1330,N_883,N_758);
and U1331 (N_1331,N_868,N_742);
nor U1332 (N_1332,N_949,N_930);
and U1333 (N_1333,N_726,N_849);
and U1334 (N_1334,N_572,N_593);
and U1335 (N_1335,N_652,N_676);
nand U1336 (N_1336,N_636,N_961);
and U1337 (N_1337,N_884,N_565);
nand U1338 (N_1338,N_713,N_817);
or U1339 (N_1339,N_811,N_664);
or U1340 (N_1340,N_800,N_873);
xor U1341 (N_1341,N_687,N_975);
and U1342 (N_1342,N_852,N_859);
and U1343 (N_1343,N_565,N_737);
or U1344 (N_1344,N_936,N_584);
nor U1345 (N_1345,N_819,N_957);
nor U1346 (N_1346,N_654,N_681);
nor U1347 (N_1347,N_638,N_835);
xor U1348 (N_1348,N_630,N_969);
or U1349 (N_1349,N_590,N_501);
nor U1350 (N_1350,N_729,N_765);
or U1351 (N_1351,N_661,N_986);
xnor U1352 (N_1352,N_751,N_880);
or U1353 (N_1353,N_672,N_554);
and U1354 (N_1354,N_572,N_536);
nor U1355 (N_1355,N_695,N_574);
nand U1356 (N_1356,N_969,N_893);
xnor U1357 (N_1357,N_599,N_658);
xor U1358 (N_1358,N_961,N_573);
nor U1359 (N_1359,N_550,N_951);
nand U1360 (N_1360,N_815,N_503);
or U1361 (N_1361,N_633,N_895);
xnor U1362 (N_1362,N_661,N_923);
nor U1363 (N_1363,N_795,N_707);
xnor U1364 (N_1364,N_534,N_542);
nor U1365 (N_1365,N_659,N_674);
and U1366 (N_1366,N_951,N_984);
nor U1367 (N_1367,N_773,N_610);
nor U1368 (N_1368,N_881,N_755);
nand U1369 (N_1369,N_556,N_588);
nand U1370 (N_1370,N_904,N_893);
or U1371 (N_1371,N_687,N_999);
and U1372 (N_1372,N_956,N_659);
xnor U1373 (N_1373,N_943,N_692);
xnor U1374 (N_1374,N_585,N_791);
or U1375 (N_1375,N_619,N_779);
nor U1376 (N_1376,N_646,N_764);
nand U1377 (N_1377,N_521,N_968);
nor U1378 (N_1378,N_953,N_644);
nor U1379 (N_1379,N_830,N_965);
or U1380 (N_1380,N_996,N_568);
xnor U1381 (N_1381,N_930,N_785);
nand U1382 (N_1382,N_714,N_783);
xnor U1383 (N_1383,N_546,N_968);
nor U1384 (N_1384,N_937,N_824);
xnor U1385 (N_1385,N_805,N_503);
or U1386 (N_1386,N_674,N_843);
nand U1387 (N_1387,N_769,N_683);
or U1388 (N_1388,N_818,N_950);
nand U1389 (N_1389,N_624,N_568);
and U1390 (N_1390,N_934,N_971);
nor U1391 (N_1391,N_845,N_988);
or U1392 (N_1392,N_951,N_906);
nor U1393 (N_1393,N_725,N_842);
and U1394 (N_1394,N_500,N_608);
nand U1395 (N_1395,N_614,N_851);
and U1396 (N_1396,N_936,N_512);
nor U1397 (N_1397,N_938,N_779);
nand U1398 (N_1398,N_785,N_615);
xor U1399 (N_1399,N_547,N_733);
nor U1400 (N_1400,N_500,N_620);
or U1401 (N_1401,N_547,N_766);
nand U1402 (N_1402,N_851,N_701);
and U1403 (N_1403,N_905,N_853);
nor U1404 (N_1404,N_711,N_551);
and U1405 (N_1405,N_583,N_990);
nand U1406 (N_1406,N_696,N_626);
xnor U1407 (N_1407,N_669,N_802);
xor U1408 (N_1408,N_816,N_571);
nand U1409 (N_1409,N_521,N_979);
and U1410 (N_1410,N_740,N_881);
nor U1411 (N_1411,N_781,N_751);
xor U1412 (N_1412,N_637,N_559);
xor U1413 (N_1413,N_671,N_650);
and U1414 (N_1414,N_504,N_875);
and U1415 (N_1415,N_914,N_517);
xor U1416 (N_1416,N_765,N_843);
nor U1417 (N_1417,N_550,N_580);
xnor U1418 (N_1418,N_826,N_544);
and U1419 (N_1419,N_957,N_573);
and U1420 (N_1420,N_874,N_934);
and U1421 (N_1421,N_676,N_540);
xor U1422 (N_1422,N_956,N_580);
and U1423 (N_1423,N_810,N_583);
and U1424 (N_1424,N_737,N_848);
nand U1425 (N_1425,N_549,N_594);
nand U1426 (N_1426,N_604,N_816);
or U1427 (N_1427,N_747,N_931);
and U1428 (N_1428,N_573,N_625);
and U1429 (N_1429,N_713,N_807);
and U1430 (N_1430,N_972,N_641);
xnor U1431 (N_1431,N_912,N_505);
and U1432 (N_1432,N_577,N_672);
nor U1433 (N_1433,N_781,N_614);
xor U1434 (N_1434,N_685,N_853);
nand U1435 (N_1435,N_733,N_878);
nand U1436 (N_1436,N_524,N_949);
nor U1437 (N_1437,N_590,N_559);
and U1438 (N_1438,N_724,N_664);
or U1439 (N_1439,N_534,N_779);
and U1440 (N_1440,N_782,N_816);
nand U1441 (N_1441,N_549,N_830);
nand U1442 (N_1442,N_754,N_526);
or U1443 (N_1443,N_557,N_781);
xnor U1444 (N_1444,N_621,N_779);
nor U1445 (N_1445,N_823,N_900);
or U1446 (N_1446,N_718,N_683);
nand U1447 (N_1447,N_912,N_667);
xor U1448 (N_1448,N_984,N_860);
or U1449 (N_1449,N_631,N_854);
nor U1450 (N_1450,N_991,N_951);
nor U1451 (N_1451,N_991,N_885);
or U1452 (N_1452,N_528,N_594);
xor U1453 (N_1453,N_929,N_826);
nor U1454 (N_1454,N_632,N_955);
nand U1455 (N_1455,N_751,N_761);
and U1456 (N_1456,N_941,N_525);
or U1457 (N_1457,N_616,N_507);
or U1458 (N_1458,N_541,N_636);
xor U1459 (N_1459,N_575,N_841);
or U1460 (N_1460,N_742,N_726);
nor U1461 (N_1461,N_950,N_787);
xor U1462 (N_1462,N_822,N_602);
nor U1463 (N_1463,N_524,N_572);
or U1464 (N_1464,N_657,N_799);
nand U1465 (N_1465,N_692,N_505);
nand U1466 (N_1466,N_586,N_553);
nor U1467 (N_1467,N_584,N_665);
or U1468 (N_1468,N_738,N_890);
or U1469 (N_1469,N_653,N_996);
and U1470 (N_1470,N_590,N_869);
nand U1471 (N_1471,N_599,N_998);
xor U1472 (N_1472,N_971,N_718);
or U1473 (N_1473,N_689,N_600);
and U1474 (N_1474,N_691,N_734);
nand U1475 (N_1475,N_709,N_856);
and U1476 (N_1476,N_768,N_804);
xnor U1477 (N_1477,N_985,N_706);
or U1478 (N_1478,N_530,N_762);
xor U1479 (N_1479,N_868,N_755);
nand U1480 (N_1480,N_842,N_678);
nand U1481 (N_1481,N_555,N_942);
nor U1482 (N_1482,N_921,N_501);
nor U1483 (N_1483,N_628,N_667);
or U1484 (N_1484,N_871,N_642);
or U1485 (N_1485,N_852,N_829);
or U1486 (N_1486,N_671,N_883);
nor U1487 (N_1487,N_621,N_613);
or U1488 (N_1488,N_606,N_695);
or U1489 (N_1489,N_521,N_908);
nand U1490 (N_1490,N_560,N_803);
or U1491 (N_1491,N_804,N_998);
xor U1492 (N_1492,N_716,N_541);
nand U1493 (N_1493,N_751,N_732);
or U1494 (N_1494,N_915,N_688);
xor U1495 (N_1495,N_611,N_613);
or U1496 (N_1496,N_519,N_515);
or U1497 (N_1497,N_539,N_634);
or U1498 (N_1498,N_716,N_764);
nand U1499 (N_1499,N_889,N_576);
nand U1500 (N_1500,N_1242,N_1164);
or U1501 (N_1501,N_1347,N_1104);
and U1502 (N_1502,N_1379,N_1223);
nor U1503 (N_1503,N_1381,N_1322);
xor U1504 (N_1504,N_1324,N_1253);
or U1505 (N_1505,N_1076,N_1110);
nor U1506 (N_1506,N_1252,N_1276);
or U1507 (N_1507,N_1405,N_1101);
xor U1508 (N_1508,N_1154,N_1304);
or U1509 (N_1509,N_1266,N_1409);
nand U1510 (N_1510,N_1335,N_1007);
nand U1511 (N_1511,N_1378,N_1091);
or U1512 (N_1512,N_1058,N_1486);
nor U1513 (N_1513,N_1408,N_1180);
and U1514 (N_1514,N_1174,N_1410);
or U1515 (N_1515,N_1213,N_1466);
xnor U1516 (N_1516,N_1018,N_1418);
and U1517 (N_1517,N_1022,N_1470);
or U1518 (N_1518,N_1032,N_1207);
xnor U1519 (N_1519,N_1234,N_1107);
and U1520 (N_1520,N_1493,N_1231);
and U1521 (N_1521,N_1286,N_1222);
and U1522 (N_1522,N_1126,N_1212);
and U1523 (N_1523,N_1219,N_1145);
or U1524 (N_1524,N_1436,N_1461);
nand U1525 (N_1525,N_1331,N_1224);
and U1526 (N_1526,N_1415,N_1259);
nand U1527 (N_1527,N_1281,N_1293);
xor U1528 (N_1528,N_1351,N_1098);
xor U1529 (N_1529,N_1177,N_1463);
and U1530 (N_1530,N_1425,N_1414);
and U1531 (N_1531,N_1271,N_1416);
nor U1532 (N_1532,N_1201,N_1264);
nand U1533 (N_1533,N_1348,N_1480);
xor U1534 (N_1534,N_1065,N_1204);
nor U1535 (N_1535,N_1393,N_1021);
xor U1536 (N_1536,N_1319,N_1491);
xor U1537 (N_1537,N_1469,N_1360);
and U1538 (N_1538,N_1310,N_1163);
xor U1539 (N_1539,N_1254,N_1394);
nand U1540 (N_1540,N_1453,N_1141);
and U1541 (N_1541,N_1395,N_1419);
or U1542 (N_1542,N_1217,N_1454);
or U1543 (N_1543,N_1450,N_1376);
nor U1544 (N_1544,N_1250,N_1489);
xnor U1545 (N_1545,N_1066,N_1037);
xnor U1546 (N_1546,N_1485,N_1333);
nor U1547 (N_1547,N_1270,N_1236);
nor U1548 (N_1548,N_1129,N_1183);
nand U1549 (N_1549,N_1467,N_1239);
nor U1550 (N_1550,N_1495,N_1114);
and U1551 (N_1551,N_1195,N_1245);
xor U1552 (N_1552,N_1434,N_1136);
nand U1553 (N_1553,N_1274,N_1277);
and U1554 (N_1554,N_1159,N_1339);
nor U1555 (N_1555,N_1228,N_1216);
and U1556 (N_1556,N_1144,N_1040);
and U1557 (N_1557,N_1192,N_1374);
nor U1558 (N_1558,N_1413,N_1388);
nand U1559 (N_1559,N_1084,N_1299);
nor U1560 (N_1560,N_1465,N_1090);
xnor U1561 (N_1561,N_1093,N_1048);
and U1562 (N_1562,N_1170,N_1105);
xnor U1563 (N_1563,N_1317,N_1297);
or U1564 (N_1564,N_1043,N_1165);
nand U1565 (N_1565,N_1312,N_1314);
nand U1566 (N_1566,N_1191,N_1382);
nor U1567 (N_1567,N_1392,N_1205);
or U1568 (N_1568,N_1143,N_1490);
or U1569 (N_1569,N_1196,N_1108);
nor U1570 (N_1570,N_1285,N_1328);
xor U1571 (N_1571,N_1476,N_1346);
and U1572 (N_1572,N_1435,N_1063);
nand U1573 (N_1573,N_1462,N_1255);
or U1574 (N_1574,N_1341,N_1122);
nand U1575 (N_1575,N_1306,N_1471);
and U1576 (N_1576,N_1373,N_1363);
and U1577 (N_1577,N_1316,N_1083);
xnor U1578 (N_1578,N_1268,N_1315);
and U1579 (N_1579,N_1189,N_1181);
nor U1580 (N_1580,N_1280,N_1230);
nor U1581 (N_1581,N_1370,N_1087);
or U1582 (N_1582,N_1368,N_1155);
or U1583 (N_1583,N_1355,N_1133);
or U1584 (N_1584,N_1118,N_1215);
or U1585 (N_1585,N_1404,N_1138);
nand U1586 (N_1586,N_1477,N_1421);
nand U1587 (N_1587,N_1160,N_1439);
and U1588 (N_1588,N_1068,N_1369);
nand U1589 (N_1589,N_1012,N_1289);
nand U1590 (N_1590,N_1171,N_1102);
xnor U1591 (N_1591,N_1124,N_1218);
and U1592 (N_1592,N_1292,N_1377);
or U1593 (N_1593,N_1197,N_1326);
or U1594 (N_1594,N_1238,N_1246);
or U1595 (N_1595,N_1130,N_1194);
or U1596 (N_1596,N_1095,N_1406);
nand U1597 (N_1597,N_1287,N_1361);
nor U1598 (N_1598,N_1142,N_1092);
xnor U1599 (N_1599,N_1120,N_1082);
nor U1600 (N_1600,N_1041,N_1232);
and U1601 (N_1601,N_1423,N_1320);
nor U1602 (N_1602,N_1015,N_1496);
or U1603 (N_1603,N_1175,N_1064);
xnor U1604 (N_1604,N_1146,N_1352);
xnor U1605 (N_1605,N_1483,N_1031);
nor U1606 (N_1606,N_1047,N_1332);
or U1607 (N_1607,N_1460,N_1256);
xor U1608 (N_1608,N_1446,N_1283);
and U1609 (N_1609,N_1096,N_1052);
and U1610 (N_1610,N_1073,N_1455);
and U1611 (N_1611,N_1221,N_1407);
xnor U1612 (N_1612,N_1176,N_1449);
or U1613 (N_1613,N_1071,N_1305);
xor U1614 (N_1614,N_1167,N_1023);
nand U1615 (N_1615,N_1033,N_1327);
or U1616 (N_1616,N_1457,N_1028);
xor U1617 (N_1617,N_1235,N_1123);
nor U1618 (N_1618,N_1488,N_1301);
nand U1619 (N_1619,N_1440,N_1429);
nor U1620 (N_1620,N_1099,N_1448);
and U1621 (N_1621,N_1147,N_1267);
nor U1622 (N_1622,N_1148,N_1337);
xnor U1623 (N_1623,N_1070,N_1121);
or U1624 (N_1624,N_1088,N_1038);
or U1625 (N_1625,N_1002,N_1139);
nand U1626 (N_1626,N_1029,N_1077);
and U1627 (N_1627,N_1056,N_1311);
xor U1628 (N_1628,N_1003,N_1251);
xor U1629 (N_1629,N_1135,N_1074);
or U1630 (N_1630,N_1132,N_1479);
or U1631 (N_1631,N_1019,N_1062);
xnor U1632 (N_1632,N_1389,N_1349);
nand U1633 (N_1633,N_1000,N_1458);
nand U1634 (N_1634,N_1203,N_1150);
xnor U1635 (N_1635,N_1225,N_1334);
nor U1636 (N_1636,N_1278,N_1067);
nand U1637 (N_1637,N_1072,N_1206);
xor U1638 (N_1638,N_1004,N_1290);
xor U1639 (N_1639,N_1411,N_1166);
and U1640 (N_1640,N_1119,N_1447);
and U1641 (N_1641,N_1309,N_1249);
nor U1642 (N_1642,N_1050,N_1010);
or U1643 (N_1643,N_1430,N_1039);
nor U1644 (N_1644,N_1350,N_1162);
nor U1645 (N_1645,N_1198,N_1433);
xor U1646 (N_1646,N_1432,N_1403);
xor U1647 (N_1647,N_1342,N_1288);
nor U1648 (N_1648,N_1226,N_1086);
nor U1649 (N_1649,N_1353,N_1422);
nor U1650 (N_1650,N_1325,N_1079);
xor U1651 (N_1651,N_1487,N_1127);
nand U1652 (N_1652,N_1030,N_1112);
or U1653 (N_1653,N_1420,N_1321);
nor U1654 (N_1654,N_1296,N_1398);
nor U1655 (N_1655,N_1359,N_1013);
xor U1656 (N_1656,N_1412,N_1386);
nor U1657 (N_1657,N_1494,N_1024);
and U1658 (N_1658,N_1243,N_1391);
or U1659 (N_1659,N_1202,N_1291);
or U1660 (N_1660,N_1459,N_1340);
and U1661 (N_1661,N_1140,N_1044);
nor U1662 (N_1662,N_1472,N_1046);
nor U1663 (N_1663,N_1061,N_1179);
nand U1664 (N_1664,N_1116,N_1153);
and U1665 (N_1665,N_1345,N_1258);
and U1666 (N_1666,N_1016,N_1357);
nor U1667 (N_1667,N_1053,N_1168);
nor U1668 (N_1668,N_1025,N_1380);
nor U1669 (N_1669,N_1428,N_1443);
nor U1670 (N_1670,N_1027,N_1478);
or U1671 (N_1671,N_1452,N_1426);
nand U1672 (N_1672,N_1307,N_1158);
or U1673 (N_1673,N_1302,N_1051);
and U1674 (N_1674,N_1329,N_1308);
xor U1675 (N_1675,N_1275,N_1375);
xnor U1676 (N_1676,N_1244,N_1397);
nand U1677 (N_1677,N_1385,N_1109);
and U1678 (N_1678,N_1240,N_1437);
nand U1679 (N_1679,N_1248,N_1001);
or U1680 (N_1680,N_1282,N_1257);
and U1681 (N_1681,N_1190,N_1134);
xor U1682 (N_1682,N_1366,N_1473);
nand U1683 (N_1683,N_1399,N_1354);
or U1684 (N_1684,N_1492,N_1484);
xnor U1685 (N_1685,N_1272,N_1300);
nand U1686 (N_1686,N_1094,N_1263);
nor U1687 (N_1687,N_1036,N_1006);
or U1688 (N_1688,N_1152,N_1057);
or U1689 (N_1689,N_1227,N_1273);
nor U1690 (N_1690,N_1424,N_1161);
nand U1691 (N_1691,N_1210,N_1438);
nor U1692 (N_1692,N_1372,N_1008);
xnor U1693 (N_1693,N_1451,N_1295);
xnor U1694 (N_1694,N_1365,N_1497);
or U1695 (N_1695,N_1384,N_1303);
or U1696 (N_1696,N_1208,N_1009);
xnor U1697 (N_1697,N_1468,N_1131);
or U1698 (N_1698,N_1279,N_1034);
nand U1699 (N_1699,N_1338,N_1020);
xnor U1700 (N_1700,N_1185,N_1362);
xnor U1701 (N_1701,N_1026,N_1209);
nor U1702 (N_1702,N_1214,N_1401);
and U1703 (N_1703,N_1117,N_1233);
nor U1704 (N_1704,N_1237,N_1184);
xnor U1705 (N_1705,N_1330,N_1417);
xnor U1706 (N_1706,N_1344,N_1113);
nand U1707 (N_1707,N_1474,N_1178);
or U1708 (N_1708,N_1156,N_1481);
or U1709 (N_1709,N_1157,N_1475);
or U1710 (N_1710,N_1464,N_1049);
or U1711 (N_1711,N_1014,N_1294);
and U1712 (N_1712,N_1358,N_1103);
xor U1713 (N_1713,N_1017,N_1269);
nand U1714 (N_1714,N_1364,N_1396);
nand U1715 (N_1715,N_1035,N_1137);
or U1716 (N_1716,N_1445,N_1149);
nand U1717 (N_1717,N_1111,N_1172);
nor U1718 (N_1718,N_1151,N_1241);
xnor U1719 (N_1719,N_1097,N_1284);
nand U1720 (N_1720,N_1211,N_1128);
xor U1721 (N_1721,N_1106,N_1182);
nor U1722 (N_1722,N_1060,N_1059);
nor U1723 (N_1723,N_1005,N_1383);
xor U1724 (N_1724,N_1261,N_1442);
xnor U1725 (N_1725,N_1427,N_1343);
xor U1726 (N_1726,N_1456,N_1011);
nor U1727 (N_1727,N_1247,N_1173);
nor U1728 (N_1728,N_1260,N_1356);
and U1729 (N_1729,N_1265,N_1229);
and U1730 (N_1730,N_1441,N_1100);
xnor U1731 (N_1731,N_1187,N_1075);
xnor U1732 (N_1732,N_1042,N_1371);
nor U1733 (N_1733,N_1089,N_1313);
nand U1734 (N_1734,N_1045,N_1080);
nor U1735 (N_1735,N_1444,N_1125);
and U1736 (N_1736,N_1262,N_1402);
nand U1737 (N_1737,N_1482,N_1431);
nor U1738 (N_1738,N_1055,N_1188);
and U1739 (N_1739,N_1400,N_1498);
xnor U1740 (N_1740,N_1298,N_1085);
xor U1741 (N_1741,N_1078,N_1069);
and U1742 (N_1742,N_1199,N_1054);
xnor U1743 (N_1743,N_1318,N_1323);
xor U1744 (N_1744,N_1336,N_1081);
nor U1745 (N_1745,N_1390,N_1186);
or U1746 (N_1746,N_1387,N_1367);
xnor U1747 (N_1747,N_1169,N_1220);
nor U1748 (N_1748,N_1499,N_1193);
nand U1749 (N_1749,N_1115,N_1200);
and U1750 (N_1750,N_1138,N_1240);
or U1751 (N_1751,N_1494,N_1059);
nand U1752 (N_1752,N_1133,N_1167);
nand U1753 (N_1753,N_1011,N_1104);
and U1754 (N_1754,N_1201,N_1186);
nand U1755 (N_1755,N_1307,N_1203);
or U1756 (N_1756,N_1445,N_1062);
xor U1757 (N_1757,N_1424,N_1155);
nand U1758 (N_1758,N_1170,N_1456);
nand U1759 (N_1759,N_1058,N_1004);
nor U1760 (N_1760,N_1260,N_1110);
or U1761 (N_1761,N_1012,N_1409);
or U1762 (N_1762,N_1379,N_1067);
and U1763 (N_1763,N_1326,N_1219);
xor U1764 (N_1764,N_1465,N_1348);
or U1765 (N_1765,N_1076,N_1211);
xnor U1766 (N_1766,N_1342,N_1102);
or U1767 (N_1767,N_1016,N_1128);
xnor U1768 (N_1768,N_1311,N_1317);
xnor U1769 (N_1769,N_1248,N_1242);
nand U1770 (N_1770,N_1319,N_1108);
nand U1771 (N_1771,N_1225,N_1165);
nor U1772 (N_1772,N_1117,N_1158);
xnor U1773 (N_1773,N_1001,N_1190);
or U1774 (N_1774,N_1339,N_1305);
nor U1775 (N_1775,N_1142,N_1288);
nand U1776 (N_1776,N_1071,N_1324);
nand U1777 (N_1777,N_1088,N_1110);
or U1778 (N_1778,N_1439,N_1198);
nor U1779 (N_1779,N_1263,N_1031);
nand U1780 (N_1780,N_1109,N_1100);
nor U1781 (N_1781,N_1382,N_1365);
or U1782 (N_1782,N_1224,N_1357);
and U1783 (N_1783,N_1083,N_1192);
and U1784 (N_1784,N_1397,N_1020);
nor U1785 (N_1785,N_1000,N_1208);
nand U1786 (N_1786,N_1133,N_1435);
nor U1787 (N_1787,N_1284,N_1024);
xor U1788 (N_1788,N_1228,N_1271);
xor U1789 (N_1789,N_1114,N_1104);
nor U1790 (N_1790,N_1311,N_1384);
nor U1791 (N_1791,N_1136,N_1103);
xor U1792 (N_1792,N_1154,N_1309);
xnor U1793 (N_1793,N_1295,N_1423);
or U1794 (N_1794,N_1226,N_1437);
or U1795 (N_1795,N_1029,N_1014);
nor U1796 (N_1796,N_1170,N_1484);
and U1797 (N_1797,N_1154,N_1039);
xnor U1798 (N_1798,N_1008,N_1480);
and U1799 (N_1799,N_1010,N_1401);
nand U1800 (N_1800,N_1000,N_1155);
nor U1801 (N_1801,N_1342,N_1207);
xor U1802 (N_1802,N_1253,N_1484);
nand U1803 (N_1803,N_1099,N_1145);
and U1804 (N_1804,N_1337,N_1003);
xor U1805 (N_1805,N_1223,N_1321);
or U1806 (N_1806,N_1120,N_1131);
nor U1807 (N_1807,N_1434,N_1452);
nand U1808 (N_1808,N_1436,N_1371);
or U1809 (N_1809,N_1043,N_1382);
nand U1810 (N_1810,N_1229,N_1051);
nor U1811 (N_1811,N_1305,N_1196);
nand U1812 (N_1812,N_1193,N_1005);
nand U1813 (N_1813,N_1208,N_1443);
nand U1814 (N_1814,N_1077,N_1423);
and U1815 (N_1815,N_1401,N_1380);
xor U1816 (N_1816,N_1110,N_1252);
nor U1817 (N_1817,N_1263,N_1131);
nor U1818 (N_1818,N_1406,N_1394);
xnor U1819 (N_1819,N_1107,N_1435);
xor U1820 (N_1820,N_1136,N_1453);
or U1821 (N_1821,N_1028,N_1279);
or U1822 (N_1822,N_1066,N_1491);
or U1823 (N_1823,N_1378,N_1262);
xor U1824 (N_1824,N_1246,N_1187);
nand U1825 (N_1825,N_1034,N_1373);
xnor U1826 (N_1826,N_1403,N_1271);
or U1827 (N_1827,N_1427,N_1019);
and U1828 (N_1828,N_1087,N_1337);
or U1829 (N_1829,N_1113,N_1235);
or U1830 (N_1830,N_1147,N_1360);
nand U1831 (N_1831,N_1234,N_1176);
and U1832 (N_1832,N_1247,N_1232);
xor U1833 (N_1833,N_1163,N_1000);
nand U1834 (N_1834,N_1206,N_1455);
nand U1835 (N_1835,N_1087,N_1259);
nor U1836 (N_1836,N_1184,N_1178);
or U1837 (N_1837,N_1230,N_1089);
nor U1838 (N_1838,N_1429,N_1003);
nand U1839 (N_1839,N_1018,N_1412);
nor U1840 (N_1840,N_1145,N_1021);
and U1841 (N_1841,N_1325,N_1197);
and U1842 (N_1842,N_1005,N_1176);
or U1843 (N_1843,N_1347,N_1446);
nand U1844 (N_1844,N_1462,N_1148);
nand U1845 (N_1845,N_1324,N_1049);
nor U1846 (N_1846,N_1237,N_1378);
xor U1847 (N_1847,N_1298,N_1485);
nor U1848 (N_1848,N_1243,N_1258);
nand U1849 (N_1849,N_1469,N_1283);
nand U1850 (N_1850,N_1167,N_1055);
xor U1851 (N_1851,N_1339,N_1073);
nand U1852 (N_1852,N_1251,N_1134);
nand U1853 (N_1853,N_1315,N_1227);
and U1854 (N_1854,N_1280,N_1324);
and U1855 (N_1855,N_1082,N_1026);
nor U1856 (N_1856,N_1220,N_1053);
and U1857 (N_1857,N_1118,N_1308);
nor U1858 (N_1858,N_1087,N_1132);
and U1859 (N_1859,N_1403,N_1053);
nor U1860 (N_1860,N_1480,N_1060);
nand U1861 (N_1861,N_1293,N_1140);
nor U1862 (N_1862,N_1267,N_1156);
and U1863 (N_1863,N_1068,N_1050);
and U1864 (N_1864,N_1278,N_1277);
xnor U1865 (N_1865,N_1249,N_1366);
nand U1866 (N_1866,N_1032,N_1458);
or U1867 (N_1867,N_1395,N_1104);
xor U1868 (N_1868,N_1026,N_1277);
nand U1869 (N_1869,N_1118,N_1198);
xnor U1870 (N_1870,N_1339,N_1117);
xor U1871 (N_1871,N_1137,N_1377);
or U1872 (N_1872,N_1045,N_1002);
xor U1873 (N_1873,N_1161,N_1174);
nand U1874 (N_1874,N_1255,N_1315);
nand U1875 (N_1875,N_1077,N_1258);
xor U1876 (N_1876,N_1275,N_1059);
nand U1877 (N_1877,N_1435,N_1389);
and U1878 (N_1878,N_1492,N_1406);
and U1879 (N_1879,N_1232,N_1241);
nor U1880 (N_1880,N_1387,N_1099);
xor U1881 (N_1881,N_1068,N_1211);
or U1882 (N_1882,N_1403,N_1383);
nand U1883 (N_1883,N_1357,N_1372);
nand U1884 (N_1884,N_1168,N_1440);
xnor U1885 (N_1885,N_1474,N_1327);
and U1886 (N_1886,N_1264,N_1105);
nand U1887 (N_1887,N_1063,N_1294);
xor U1888 (N_1888,N_1142,N_1119);
nor U1889 (N_1889,N_1258,N_1118);
nor U1890 (N_1890,N_1314,N_1480);
and U1891 (N_1891,N_1423,N_1269);
nand U1892 (N_1892,N_1396,N_1012);
nand U1893 (N_1893,N_1375,N_1406);
nor U1894 (N_1894,N_1241,N_1466);
or U1895 (N_1895,N_1337,N_1357);
nor U1896 (N_1896,N_1463,N_1285);
and U1897 (N_1897,N_1342,N_1456);
nand U1898 (N_1898,N_1046,N_1383);
and U1899 (N_1899,N_1353,N_1073);
xor U1900 (N_1900,N_1115,N_1120);
and U1901 (N_1901,N_1130,N_1216);
or U1902 (N_1902,N_1023,N_1030);
xor U1903 (N_1903,N_1454,N_1429);
or U1904 (N_1904,N_1085,N_1017);
nand U1905 (N_1905,N_1233,N_1000);
and U1906 (N_1906,N_1402,N_1244);
or U1907 (N_1907,N_1013,N_1458);
or U1908 (N_1908,N_1200,N_1367);
or U1909 (N_1909,N_1432,N_1420);
xor U1910 (N_1910,N_1058,N_1124);
or U1911 (N_1911,N_1032,N_1416);
xnor U1912 (N_1912,N_1357,N_1441);
xor U1913 (N_1913,N_1120,N_1418);
or U1914 (N_1914,N_1026,N_1190);
or U1915 (N_1915,N_1335,N_1031);
xor U1916 (N_1916,N_1233,N_1331);
nand U1917 (N_1917,N_1162,N_1146);
nand U1918 (N_1918,N_1266,N_1174);
nand U1919 (N_1919,N_1306,N_1472);
xor U1920 (N_1920,N_1498,N_1005);
nor U1921 (N_1921,N_1197,N_1043);
nand U1922 (N_1922,N_1273,N_1313);
xnor U1923 (N_1923,N_1444,N_1424);
nor U1924 (N_1924,N_1294,N_1400);
nor U1925 (N_1925,N_1004,N_1390);
nor U1926 (N_1926,N_1455,N_1401);
xnor U1927 (N_1927,N_1264,N_1372);
and U1928 (N_1928,N_1361,N_1109);
nor U1929 (N_1929,N_1444,N_1174);
nor U1930 (N_1930,N_1458,N_1018);
nand U1931 (N_1931,N_1244,N_1329);
and U1932 (N_1932,N_1379,N_1243);
nor U1933 (N_1933,N_1187,N_1346);
and U1934 (N_1934,N_1422,N_1193);
xnor U1935 (N_1935,N_1124,N_1232);
nor U1936 (N_1936,N_1362,N_1198);
nor U1937 (N_1937,N_1466,N_1492);
nor U1938 (N_1938,N_1376,N_1092);
xor U1939 (N_1939,N_1317,N_1352);
xnor U1940 (N_1940,N_1303,N_1420);
or U1941 (N_1941,N_1091,N_1236);
nor U1942 (N_1942,N_1321,N_1000);
nand U1943 (N_1943,N_1359,N_1236);
nand U1944 (N_1944,N_1266,N_1419);
or U1945 (N_1945,N_1001,N_1305);
xnor U1946 (N_1946,N_1290,N_1448);
or U1947 (N_1947,N_1237,N_1059);
or U1948 (N_1948,N_1466,N_1351);
and U1949 (N_1949,N_1256,N_1461);
or U1950 (N_1950,N_1386,N_1122);
nor U1951 (N_1951,N_1350,N_1209);
xnor U1952 (N_1952,N_1169,N_1135);
nor U1953 (N_1953,N_1371,N_1087);
and U1954 (N_1954,N_1198,N_1430);
and U1955 (N_1955,N_1493,N_1191);
nand U1956 (N_1956,N_1432,N_1178);
and U1957 (N_1957,N_1015,N_1493);
and U1958 (N_1958,N_1058,N_1279);
nand U1959 (N_1959,N_1045,N_1054);
xor U1960 (N_1960,N_1456,N_1203);
and U1961 (N_1961,N_1495,N_1198);
xor U1962 (N_1962,N_1266,N_1235);
and U1963 (N_1963,N_1240,N_1450);
xnor U1964 (N_1964,N_1299,N_1452);
or U1965 (N_1965,N_1354,N_1152);
nand U1966 (N_1966,N_1412,N_1236);
xor U1967 (N_1967,N_1360,N_1024);
nand U1968 (N_1968,N_1001,N_1126);
and U1969 (N_1969,N_1373,N_1377);
nand U1970 (N_1970,N_1195,N_1127);
nand U1971 (N_1971,N_1112,N_1419);
nand U1972 (N_1972,N_1315,N_1272);
nand U1973 (N_1973,N_1122,N_1242);
nand U1974 (N_1974,N_1287,N_1402);
nand U1975 (N_1975,N_1459,N_1219);
and U1976 (N_1976,N_1413,N_1050);
nand U1977 (N_1977,N_1416,N_1194);
nor U1978 (N_1978,N_1390,N_1402);
xnor U1979 (N_1979,N_1322,N_1428);
or U1980 (N_1980,N_1064,N_1244);
or U1981 (N_1981,N_1076,N_1118);
and U1982 (N_1982,N_1434,N_1039);
nand U1983 (N_1983,N_1119,N_1055);
nand U1984 (N_1984,N_1453,N_1158);
nand U1985 (N_1985,N_1342,N_1096);
nor U1986 (N_1986,N_1176,N_1137);
or U1987 (N_1987,N_1455,N_1014);
and U1988 (N_1988,N_1004,N_1393);
xor U1989 (N_1989,N_1112,N_1025);
and U1990 (N_1990,N_1166,N_1320);
xor U1991 (N_1991,N_1138,N_1424);
or U1992 (N_1992,N_1393,N_1276);
and U1993 (N_1993,N_1309,N_1075);
nor U1994 (N_1994,N_1033,N_1446);
nand U1995 (N_1995,N_1086,N_1169);
nor U1996 (N_1996,N_1347,N_1480);
xor U1997 (N_1997,N_1492,N_1242);
xnor U1998 (N_1998,N_1268,N_1434);
nand U1999 (N_1999,N_1150,N_1253);
xor U2000 (N_2000,N_1638,N_1879);
and U2001 (N_2001,N_1713,N_1597);
xnor U2002 (N_2002,N_1580,N_1570);
nor U2003 (N_2003,N_1553,N_1880);
nor U2004 (N_2004,N_1962,N_1610);
and U2005 (N_2005,N_1500,N_1598);
or U2006 (N_2006,N_1948,N_1842);
and U2007 (N_2007,N_1536,N_1994);
and U2008 (N_2008,N_1819,N_1967);
and U2009 (N_2009,N_1956,N_1796);
nand U2010 (N_2010,N_1798,N_1832);
and U2011 (N_2011,N_1606,N_1579);
and U2012 (N_2012,N_1601,N_1679);
xnor U2013 (N_2013,N_1671,N_1916);
xnor U2014 (N_2014,N_1603,N_1735);
nor U2015 (N_2015,N_1985,N_1787);
and U2016 (N_2016,N_1673,N_1803);
nand U2017 (N_2017,N_1582,N_1546);
nor U2018 (N_2018,N_1693,N_1890);
nand U2019 (N_2019,N_1760,N_1745);
and U2020 (N_2020,N_1641,N_1504);
nand U2021 (N_2021,N_1812,N_1823);
and U2022 (N_2022,N_1992,N_1799);
or U2023 (N_2023,N_1868,N_1981);
and U2024 (N_2024,N_1851,N_1505);
or U2025 (N_2025,N_1840,N_1839);
nor U2026 (N_2026,N_1651,N_1913);
nand U2027 (N_2027,N_1650,N_1736);
nor U2028 (N_2028,N_1747,N_1810);
nand U2029 (N_2029,N_1847,N_1562);
nand U2030 (N_2030,N_1827,N_1881);
nand U2031 (N_2031,N_1507,N_1518);
nand U2032 (N_2032,N_1521,N_1894);
nand U2033 (N_2033,N_1949,N_1891);
nor U2034 (N_2034,N_1593,N_1777);
nor U2035 (N_2035,N_1738,N_1729);
xor U2036 (N_2036,N_1857,N_1677);
nor U2037 (N_2037,N_1618,N_1841);
and U2038 (N_2038,N_1969,N_1686);
and U2039 (N_2039,N_1733,N_1631);
xor U2040 (N_2040,N_1608,N_1990);
or U2041 (N_2041,N_1587,N_1634);
nand U2042 (N_2042,N_1542,N_1909);
or U2043 (N_2043,N_1946,N_1706);
or U2044 (N_2044,N_1635,N_1600);
or U2045 (N_2045,N_1555,N_1554);
xor U2046 (N_2046,N_1757,N_1972);
xor U2047 (N_2047,N_1649,N_1674);
nand U2048 (N_2048,N_1765,N_1564);
or U2049 (N_2049,N_1940,N_1699);
nand U2050 (N_2050,N_1814,N_1843);
xnor U2051 (N_2051,N_1973,N_1933);
nor U2052 (N_2052,N_1742,N_1975);
xnor U2053 (N_2053,N_1636,N_1987);
xnor U2054 (N_2054,N_1860,N_1807);
or U2055 (N_2055,N_1774,N_1947);
nor U2056 (N_2056,N_1691,N_1567);
nand U2057 (N_2057,N_1853,N_1805);
or U2058 (N_2058,N_1936,N_1758);
or U2059 (N_2059,N_1914,N_1833);
nand U2060 (N_2060,N_1563,N_1731);
xnor U2061 (N_2061,N_1604,N_1503);
and U2062 (N_2062,N_1859,N_1535);
nand U2063 (N_2063,N_1957,N_1509);
nand U2064 (N_2064,N_1617,N_1780);
nor U2065 (N_2065,N_1937,N_1676);
or U2066 (N_2066,N_1788,N_1565);
nor U2067 (N_2067,N_1640,N_1690);
xor U2068 (N_2068,N_1872,N_1613);
nor U2069 (N_2069,N_1854,N_1719);
and U2070 (N_2070,N_1718,N_1510);
and U2071 (N_2071,N_1547,N_1566);
nor U2072 (N_2072,N_1659,N_1801);
xnor U2073 (N_2073,N_1834,N_1688);
or U2074 (N_2074,N_1978,N_1974);
nand U2075 (N_2075,N_1938,N_1895);
nand U2076 (N_2076,N_1870,N_1715);
and U2077 (N_2077,N_1685,N_1941);
and U2078 (N_2078,N_1825,N_1701);
xor U2079 (N_2079,N_1885,N_1928);
xor U2080 (N_2080,N_1900,N_1664);
nand U2081 (N_2081,N_1951,N_1931);
nor U2082 (N_2082,N_1714,N_1906);
xor U2083 (N_2083,N_1668,N_1995);
or U2084 (N_2084,N_1539,N_1532);
or U2085 (N_2085,N_1945,N_1764);
and U2086 (N_2086,N_1771,N_1616);
and U2087 (N_2087,N_1520,N_1929);
nand U2088 (N_2088,N_1922,N_1911);
nor U2089 (N_2089,N_1915,N_1522);
xnor U2090 (N_2090,N_1590,N_1980);
nand U2091 (N_2091,N_1519,N_1727);
or U2092 (N_2092,N_1923,N_1892);
and U2093 (N_2093,N_1768,N_1611);
xor U2094 (N_2094,N_1815,N_1556);
nor U2095 (N_2095,N_1658,N_1512);
nand U2096 (N_2096,N_1935,N_1537);
nor U2097 (N_2097,N_1529,N_1550);
nor U2098 (N_2098,N_1501,N_1950);
or U2099 (N_2099,N_1836,N_1667);
and U2100 (N_2100,N_1577,N_1762);
and U2101 (N_2101,N_1934,N_1709);
and U2102 (N_2102,N_1811,N_1878);
and U2103 (N_2103,N_1795,N_1644);
and U2104 (N_2104,N_1919,N_1769);
xor U2105 (N_2105,N_1741,N_1898);
or U2106 (N_2106,N_1921,N_1605);
nor U2107 (N_2107,N_1983,N_1952);
and U2108 (N_2108,N_1508,N_1607);
nor U2109 (N_2109,N_1904,N_1568);
and U2110 (N_2110,N_1794,N_1646);
nor U2111 (N_2111,N_1991,N_1797);
nor U2112 (N_2112,N_1920,N_1767);
and U2113 (N_2113,N_1573,N_1902);
nand U2114 (N_2114,N_1627,N_1986);
xnor U2115 (N_2115,N_1903,N_1557);
nand U2116 (N_2116,N_1831,N_1943);
nand U2117 (N_2117,N_1687,N_1866);
xnor U2118 (N_2118,N_1953,N_1785);
nand U2119 (N_2119,N_1846,N_1707);
nor U2120 (N_2120,N_1591,N_1726);
nand U2121 (N_2121,N_1786,N_1822);
nand U2122 (N_2122,N_1622,N_1761);
nand U2123 (N_2123,N_1800,N_1632);
and U2124 (N_2124,N_1540,N_1855);
and U2125 (N_2125,N_1963,N_1506);
nor U2126 (N_2126,N_1924,N_1663);
nand U2127 (N_2127,N_1932,N_1524);
nor U2128 (N_2128,N_1625,N_1558);
xnor U2129 (N_2129,N_1999,N_1721);
nand U2130 (N_2130,N_1865,N_1645);
or U2131 (N_2131,N_1525,N_1643);
xnor U2132 (N_2132,N_1626,N_1630);
nor U2133 (N_2133,N_1702,N_1844);
or U2134 (N_2134,N_1551,N_1887);
xnor U2135 (N_2135,N_1901,N_1817);
nor U2136 (N_2136,N_1837,N_1942);
xor U2137 (N_2137,N_1628,N_1516);
or U2138 (N_2138,N_1633,N_1620);
and U2139 (N_2139,N_1862,N_1700);
nor U2140 (N_2140,N_1778,N_1734);
nand U2141 (N_2141,N_1623,N_1873);
nand U2142 (N_2142,N_1581,N_1907);
nand U2143 (N_2143,N_1681,N_1569);
nand U2144 (N_2144,N_1875,N_1548);
xnor U2145 (N_2145,N_1694,N_1530);
nor U2146 (N_2146,N_1829,N_1653);
and U2147 (N_2147,N_1806,N_1559);
and U2148 (N_2148,N_1711,N_1514);
nand U2149 (N_2149,N_1808,N_1656);
or U2150 (N_2150,N_1680,N_1899);
xor U2151 (N_2151,N_1657,N_1982);
or U2152 (N_2152,N_1752,N_1861);
xor U2153 (N_2153,N_1589,N_1867);
or U2154 (N_2154,N_1908,N_1670);
nand U2155 (N_2155,N_1882,N_1748);
xnor U2156 (N_2156,N_1523,N_1665);
or U2157 (N_2157,N_1594,N_1662);
and U2158 (N_2158,N_1884,N_1669);
or U2159 (N_2159,N_1609,N_1998);
and U2160 (N_2160,N_1820,N_1918);
and U2161 (N_2161,N_1858,N_1716);
and U2162 (N_2162,N_1912,N_1615);
and U2163 (N_2163,N_1578,N_1544);
or U2164 (N_2164,N_1743,N_1776);
or U2165 (N_2165,N_1592,N_1792);
or U2166 (N_2166,N_1538,N_1960);
and U2167 (N_2167,N_1804,N_1828);
and U2168 (N_2168,N_1897,N_1583);
nand U2169 (N_2169,N_1958,N_1939);
and U2170 (N_2170,N_1964,N_1730);
nor U2171 (N_2171,N_1988,N_1955);
or U2172 (N_2172,N_1545,N_1655);
xnor U2173 (N_2173,N_1838,N_1809);
nor U2174 (N_2174,N_1612,N_1692);
nand U2175 (N_2175,N_1585,N_1888);
xnor U2176 (N_2176,N_1886,N_1511);
nor U2177 (N_2177,N_1763,N_1750);
nand U2178 (N_2178,N_1528,N_1639);
and U2179 (N_2179,N_1652,N_1813);
xnor U2180 (N_2180,N_1683,N_1560);
xnor U2181 (N_2181,N_1977,N_1779);
nand U2182 (N_2182,N_1997,N_1527);
nor U2183 (N_2183,N_1648,N_1791);
xnor U2184 (N_2184,N_1818,N_1584);
xnor U2185 (N_2185,N_1697,N_1624);
nor U2186 (N_2186,N_1678,N_1789);
nand U2187 (N_2187,N_1874,N_1712);
or U2188 (N_2188,N_1826,N_1954);
and U2189 (N_2189,N_1864,N_1526);
or U2190 (N_2190,N_1925,N_1850);
or U2191 (N_2191,N_1596,N_1513);
xnor U2192 (N_2192,N_1703,N_1749);
and U2193 (N_2193,N_1739,N_1572);
xnor U2194 (N_2194,N_1772,N_1517);
and U2195 (N_2195,N_1737,N_1732);
xnor U2196 (N_2196,N_1848,N_1927);
and U2197 (N_2197,N_1984,N_1599);
xnor U2198 (N_2198,N_1849,N_1724);
and U2199 (N_2199,N_1710,N_1821);
nor U2200 (N_2200,N_1852,N_1696);
nand U2201 (N_2201,N_1770,N_1723);
nand U2202 (N_2202,N_1830,N_1744);
and U2203 (N_2203,N_1753,N_1588);
or U2204 (N_2204,N_1602,N_1595);
or U2205 (N_2205,N_1534,N_1845);
nand U2206 (N_2206,N_1773,N_1754);
or U2207 (N_2207,N_1802,N_1619);
and U2208 (N_2208,N_1698,N_1684);
nand U2209 (N_2209,N_1647,N_1728);
nor U2210 (N_2210,N_1725,N_1660);
nand U2211 (N_2211,N_1782,N_1863);
nand U2212 (N_2212,N_1549,N_1968);
xnor U2213 (N_2213,N_1871,N_1695);
or U2214 (N_2214,N_1746,N_1893);
or U2215 (N_2215,N_1989,N_1944);
nand U2216 (N_2216,N_1876,N_1642);
nand U2217 (N_2217,N_1543,N_1961);
xor U2218 (N_2218,N_1751,N_1971);
nand U2219 (N_2219,N_1552,N_1629);
and U2220 (N_2220,N_1720,N_1905);
and U2221 (N_2221,N_1970,N_1883);
and U2222 (N_2222,N_1571,N_1869);
nor U2223 (N_2223,N_1816,N_1689);
and U2224 (N_2224,N_1910,N_1637);
or U2225 (N_2225,N_1666,N_1704);
or U2226 (N_2226,N_1759,N_1775);
nand U2227 (N_2227,N_1515,N_1966);
nor U2228 (N_2228,N_1784,N_1783);
xnor U2229 (N_2229,N_1889,N_1576);
nand U2230 (N_2230,N_1722,N_1976);
nor U2231 (N_2231,N_1755,N_1672);
nor U2232 (N_2232,N_1835,N_1766);
nand U2233 (N_2233,N_1824,N_1682);
and U2234 (N_2234,N_1705,N_1926);
xor U2235 (N_2235,N_1531,N_1917);
xnor U2236 (N_2236,N_1790,N_1856);
or U2237 (N_2237,N_1740,N_1574);
xor U2238 (N_2238,N_1781,N_1661);
or U2239 (N_2239,N_1996,N_1675);
nor U2240 (N_2240,N_1793,N_1614);
nand U2241 (N_2241,N_1896,N_1654);
xnor U2242 (N_2242,N_1877,N_1502);
and U2243 (N_2243,N_1979,N_1717);
nand U2244 (N_2244,N_1965,N_1708);
and U2245 (N_2245,N_1541,N_1575);
nand U2246 (N_2246,N_1586,N_1930);
or U2247 (N_2247,N_1959,N_1993);
nand U2248 (N_2248,N_1561,N_1533);
or U2249 (N_2249,N_1756,N_1621);
nor U2250 (N_2250,N_1831,N_1751);
or U2251 (N_2251,N_1527,N_1626);
nand U2252 (N_2252,N_1795,N_1729);
and U2253 (N_2253,N_1608,N_1582);
and U2254 (N_2254,N_1895,N_1676);
and U2255 (N_2255,N_1711,N_1755);
nor U2256 (N_2256,N_1539,N_1564);
nor U2257 (N_2257,N_1982,N_1624);
or U2258 (N_2258,N_1823,N_1619);
nor U2259 (N_2259,N_1969,N_1869);
and U2260 (N_2260,N_1883,N_1772);
or U2261 (N_2261,N_1855,N_1764);
nor U2262 (N_2262,N_1505,N_1818);
nor U2263 (N_2263,N_1817,N_1573);
nand U2264 (N_2264,N_1849,N_1706);
nand U2265 (N_2265,N_1788,N_1657);
or U2266 (N_2266,N_1627,N_1768);
or U2267 (N_2267,N_1602,N_1572);
nor U2268 (N_2268,N_1951,N_1994);
xnor U2269 (N_2269,N_1961,N_1730);
nand U2270 (N_2270,N_1926,N_1856);
and U2271 (N_2271,N_1567,N_1976);
nor U2272 (N_2272,N_1553,N_1592);
nand U2273 (N_2273,N_1580,N_1923);
nor U2274 (N_2274,N_1737,N_1803);
xor U2275 (N_2275,N_1729,N_1973);
xor U2276 (N_2276,N_1502,N_1604);
nand U2277 (N_2277,N_1788,N_1824);
or U2278 (N_2278,N_1537,N_1960);
nand U2279 (N_2279,N_1930,N_1864);
and U2280 (N_2280,N_1554,N_1561);
nor U2281 (N_2281,N_1843,N_1853);
nor U2282 (N_2282,N_1908,N_1620);
or U2283 (N_2283,N_1519,N_1762);
nor U2284 (N_2284,N_1820,N_1914);
nor U2285 (N_2285,N_1544,N_1714);
or U2286 (N_2286,N_1978,N_1897);
nand U2287 (N_2287,N_1767,N_1771);
and U2288 (N_2288,N_1591,N_1581);
and U2289 (N_2289,N_1698,N_1535);
nor U2290 (N_2290,N_1693,N_1519);
or U2291 (N_2291,N_1632,N_1534);
nor U2292 (N_2292,N_1608,N_1782);
nor U2293 (N_2293,N_1674,N_1986);
and U2294 (N_2294,N_1727,N_1799);
nand U2295 (N_2295,N_1588,N_1889);
xnor U2296 (N_2296,N_1757,N_1794);
and U2297 (N_2297,N_1686,N_1679);
nor U2298 (N_2298,N_1700,N_1856);
nor U2299 (N_2299,N_1532,N_1705);
or U2300 (N_2300,N_1946,N_1851);
or U2301 (N_2301,N_1755,N_1825);
nand U2302 (N_2302,N_1685,N_1691);
nor U2303 (N_2303,N_1599,N_1760);
xnor U2304 (N_2304,N_1714,N_1765);
nor U2305 (N_2305,N_1984,N_1973);
nand U2306 (N_2306,N_1528,N_1757);
or U2307 (N_2307,N_1820,N_1892);
and U2308 (N_2308,N_1559,N_1609);
and U2309 (N_2309,N_1797,N_1864);
nand U2310 (N_2310,N_1799,N_1938);
nor U2311 (N_2311,N_1934,N_1985);
nand U2312 (N_2312,N_1690,N_1642);
nand U2313 (N_2313,N_1957,N_1833);
xnor U2314 (N_2314,N_1947,N_1552);
and U2315 (N_2315,N_1883,N_1695);
and U2316 (N_2316,N_1901,N_1782);
xnor U2317 (N_2317,N_1730,N_1524);
nor U2318 (N_2318,N_1575,N_1667);
nor U2319 (N_2319,N_1954,N_1883);
xor U2320 (N_2320,N_1692,N_1801);
nand U2321 (N_2321,N_1719,N_1932);
xor U2322 (N_2322,N_1951,N_1799);
xnor U2323 (N_2323,N_1580,N_1789);
nand U2324 (N_2324,N_1590,N_1762);
xor U2325 (N_2325,N_1799,N_1889);
nor U2326 (N_2326,N_1507,N_1634);
xnor U2327 (N_2327,N_1676,N_1703);
and U2328 (N_2328,N_1869,N_1825);
xnor U2329 (N_2329,N_1961,N_1562);
xor U2330 (N_2330,N_1867,N_1996);
nand U2331 (N_2331,N_1747,N_1862);
or U2332 (N_2332,N_1906,N_1806);
and U2333 (N_2333,N_1502,N_1835);
or U2334 (N_2334,N_1914,N_1855);
nor U2335 (N_2335,N_1845,N_1875);
xor U2336 (N_2336,N_1535,N_1935);
and U2337 (N_2337,N_1942,N_1662);
or U2338 (N_2338,N_1770,N_1906);
or U2339 (N_2339,N_1745,N_1581);
nand U2340 (N_2340,N_1686,N_1881);
nand U2341 (N_2341,N_1788,N_1874);
xnor U2342 (N_2342,N_1714,N_1502);
nor U2343 (N_2343,N_1611,N_1574);
or U2344 (N_2344,N_1839,N_1580);
nand U2345 (N_2345,N_1511,N_1554);
nor U2346 (N_2346,N_1624,N_1839);
xor U2347 (N_2347,N_1634,N_1793);
nor U2348 (N_2348,N_1509,N_1639);
or U2349 (N_2349,N_1751,N_1998);
nor U2350 (N_2350,N_1787,N_1561);
xor U2351 (N_2351,N_1828,N_1896);
xor U2352 (N_2352,N_1848,N_1693);
nand U2353 (N_2353,N_1849,N_1841);
and U2354 (N_2354,N_1546,N_1937);
and U2355 (N_2355,N_1901,N_1768);
xnor U2356 (N_2356,N_1598,N_1533);
and U2357 (N_2357,N_1664,N_1799);
nand U2358 (N_2358,N_1765,N_1800);
or U2359 (N_2359,N_1686,N_1802);
xor U2360 (N_2360,N_1970,N_1835);
and U2361 (N_2361,N_1783,N_1941);
nand U2362 (N_2362,N_1897,N_1518);
or U2363 (N_2363,N_1842,N_1721);
nor U2364 (N_2364,N_1713,N_1893);
nand U2365 (N_2365,N_1761,N_1922);
xnor U2366 (N_2366,N_1845,N_1607);
and U2367 (N_2367,N_1870,N_1614);
or U2368 (N_2368,N_1512,N_1567);
nand U2369 (N_2369,N_1871,N_1530);
nor U2370 (N_2370,N_1773,N_1570);
and U2371 (N_2371,N_1931,N_1596);
and U2372 (N_2372,N_1772,N_1627);
nor U2373 (N_2373,N_1924,N_1715);
or U2374 (N_2374,N_1939,N_1998);
and U2375 (N_2375,N_1561,N_1943);
xor U2376 (N_2376,N_1792,N_1793);
and U2377 (N_2377,N_1757,N_1857);
nor U2378 (N_2378,N_1638,N_1823);
nor U2379 (N_2379,N_1616,N_1777);
or U2380 (N_2380,N_1835,N_1874);
and U2381 (N_2381,N_1891,N_1604);
nor U2382 (N_2382,N_1693,N_1790);
and U2383 (N_2383,N_1921,N_1579);
or U2384 (N_2384,N_1699,N_1707);
xor U2385 (N_2385,N_1579,N_1944);
xor U2386 (N_2386,N_1697,N_1507);
nor U2387 (N_2387,N_1674,N_1697);
nand U2388 (N_2388,N_1734,N_1664);
and U2389 (N_2389,N_1840,N_1740);
or U2390 (N_2390,N_1681,N_1741);
or U2391 (N_2391,N_1972,N_1781);
or U2392 (N_2392,N_1984,N_1810);
or U2393 (N_2393,N_1971,N_1707);
nand U2394 (N_2394,N_1661,N_1922);
nand U2395 (N_2395,N_1792,N_1827);
xnor U2396 (N_2396,N_1929,N_1685);
xor U2397 (N_2397,N_1838,N_1672);
nand U2398 (N_2398,N_1726,N_1859);
nand U2399 (N_2399,N_1659,N_1500);
xor U2400 (N_2400,N_1632,N_1975);
xor U2401 (N_2401,N_1906,N_1720);
xor U2402 (N_2402,N_1987,N_1741);
and U2403 (N_2403,N_1757,N_1739);
nor U2404 (N_2404,N_1982,N_1728);
or U2405 (N_2405,N_1576,N_1902);
or U2406 (N_2406,N_1789,N_1741);
nor U2407 (N_2407,N_1785,N_1566);
nand U2408 (N_2408,N_1511,N_1805);
xor U2409 (N_2409,N_1965,N_1810);
xor U2410 (N_2410,N_1945,N_1746);
and U2411 (N_2411,N_1837,N_1758);
and U2412 (N_2412,N_1564,N_1660);
nor U2413 (N_2413,N_1622,N_1727);
or U2414 (N_2414,N_1661,N_1815);
and U2415 (N_2415,N_1803,N_1723);
nor U2416 (N_2416,N_1549,N_1612);
nand U2417 (N_2417,N_1747,N_1968);
and U2418 (N_2418,N_1748,N_1926);
or U2419 (N_2419,N_1870,N_1562);
xor U2420 (N_2420,N_1688,N_1806);
xnor U2421 (N_2421,N_1774,N_1704);
nor U2422 (N_2422,N_1556,N_1512);
or U2423 (N_2423,N_1933,N_1530);
nor U2424 (N_2424,N_1849,N_1804);
and U2425 (N_2425,N_1884,N_1823);
xor U2426 (N_2426,N_1510,N_1532);
and U2427 (N_2427,N_1531,N_1741);
or U2428 (N_2428,N_1732,N_1571);
nor U2429 (N_2429,N_1913,N_1930);
nand U2430 (N_2430,N_1715,N_1520);
xor U2431 (N_2431,N_1925,N_1890);
nor U2432 (N_2432,N_1633,N_1836);
and U2433 (N_2433,N_1884,N_1558);
or U2434 (N_2434,N_1792,N_1505);
xnor U2435 (N_2435,N_1676,N_1967);
xor U2436 (N_2436,N_1720,N_1777);
xnor U2437 (N_2437,N_1988,N_1964);
xor U2438 (N_2438,N_1723,N_1663);
nor U2439 (N_2439,N_1854,N_1541);
xor U2440 (N_2440,N_1758,N_1995);
nand U2441 (N_2441,N_1859,N_1735);
xnor U2442 (N_2442,N_1549,N_1690);
nand U2443 (N_2443,N_1699,N_1709);
nand U2444 (N_2444,N_1633,N_1674);
or U2445 (N_2445,N_1773,N_1664);
xor U2446 (N_2446,N_1877,N_1646);
xnor U2447 (N_2447,N_1764,N_1799);
and U2448 (N_2448,N_1976,N_1899);
and U2449 (N_2449,N_1832,N_1748);
xnor U2450 (N_2450,N_1687,N_1656);
nor U2451 (N_2451,N_1968,N_1836);
xor U2452 (N_2452,N_1554,N_1587);
nor U2453 (N_2453,N_1550,N_1931);
or U2454 (N_2454,N_1796,N_1663);
nor U2455 (N_2455,N_1816,N_1646);
or U2456 (N_2456,N_1566,N_1889);
nand U2457 (N_2457,N_1842,N_1707);
nor U2458 (N_2458,N_1627,N_1710);
xor U2459 (N_2459,N_1834,N_1691);
nand U2460 (N_2460,N_1668,N_1765);
nand U2461 (N_2461,N_1538,N_1859);
or U2462 (N_2462,N_1883,N_1847);
nand U2463 (N_2463,N_1586,N_1636);
xnor U2464 (N_2464,N_1527,N_1613);
nor U2465 (N_2465,N_1580,N_1849);
nand U2466 (N_2466,N_1589,N_1954);
nor U2467 (N_2467,N_1792,N_1894);
xor U2468 (N_2468,N_1757,N_1749);
nand U2469 (N_2469,N_1618,N_1960);
xnor U2470 (N_2470,N_1790,N_1750);
and U2471 (N_2471,N_1962,N_1911);
and U2472 (N_2472,N_1587,N_1507);
nand U2473 (N_2473,N_1895,N_1500);
nand U2474 (N_2474,N_1918,N_1815);
nand U2475 (N_2475,N_1837,N_1874);
and U2476 (N_2476,N_1874,N_1545);
nand U2477 (N_2477,N_1678,N_1829);
and U2478 (N_2478,N_1818,N_1737);
and U2479 (N_2479,N_1662,N_1976);
or U2480 (N_2480,N_1932,N_1564);
xnor U2481 (N_2481,N_1757,N_1879);
or U2482 (N_2482,N_1776,N_1788);
nand U2483 (N_2483,N_1574,N_1938);
nand U2484 (N_2484,N_1911,N_1725);
xor U2485 (N_2485,N_1685,N_1536);
xor U2486 (N_2486,N_1882,N_1868);
and U2487 (N_2487,N_1617,N_1934);
nor U2488 (N_2488,N_1985,N_1594);
nor U2489 (N_2489,N_1514,N_1865);
nor U2490 (N_2490,N_1982,N_1541);
xor U2491 (N_2491,N_1529,N_1586);
xor U2492 (N_2492,N_1835,N_1679);
and U2493 (N_2493,N_1664,N_1988);
xnor U2494 (N_2494,N_1569,N_1654);
xor U2495 (N_2495,N_1536,N_1821);
or U2496 (N_2496,N_1720,N_1746);
or U2497 (N_2497,N_1796,N_1975);
xor U2498 (N_2498,N_1821,N_1627);
nor U2499 (N_2499,N_1505,N_1580);
or U2500 (N_2500,N_2002,N_2076);
and U2501 (N_2501,N_2177,N_2173);
or U2502 (N_2502,N_2244,N_2105);
xor U2503 (N_2503,N_2292,N_2263);
or U2504 (N_2504,N_2127,N_2289);
xor U2505 (N_2505,N_2125,N_2174);
xor U2506 (N_2506,N_2410,N_2024);
and U2507 (N_2507,N_2334,N_2182);
or U2508 (N_2508,N_2286,N_2219);
and U2509 (N_2509,N_2402,N_2029);
nor U2510 (N_2510,N_2128,N_2456);
xor U2511 (N_2511,N_2232,N_2435);
xnor U2512 (N_2512,N_2101,N_2179);
and U2513 (N_2513,N_2248,N_2097);
nor U2514 (N_2514,N_2006,N_2160);
xor U2515 (N_2515,N_2418,N_2276);
nand U2516 (N_2516,N_2324,N_2480);
xor U2517 (N_2517,N_2359,N_2090);
nor U2518 (N_2518,N_2197,N_2004);
or U2519 (N_2519,N_2208,N_2371);
or U2520 (N_2520,N_2149,N_2466);
or U2521 (N_2521,N_2467,N_2134);
and U2522 (N_2522,N_2448,N_2071);
xnor U2523 (N_2523,N_2189,N_2463);
nand U2524 (N_2524,N_2027,N_2056);
nor U2525 (N_2525,N_2477,N_2345);
or U2526 (N_2526,N_2238,N_2034);
nand U2527 (N_2527,N_2469,N_2307);
nor U2528 (N_2528,N_2319,N_2057);
nand U2529 (N_2529,N_2042,N_2183);
xnor U2530 (N_2530,N_2385,N_2171);
nor U2531 (N_2531,N_2404,N_2329);
nor U2532 (N_2532,N_2100,N_2495);
and U2533 (N_2533,N_2356,N_2077);
and U2534 (N_2534,N_2227,N_2479);
or U2535 (N_2535,N_2215,N_2114);
nand U2536 (N_2536,N_2428,N_2031);
or U2537 (N_2537,N_2360,N_2164);
nand U2538 (N_2538,N_2204,N_2451);
nor U2539 (N_2539,N_2054,N_2152);
nor U2540 (N_2540,N_2303,N_2066);
nor U2541 (N_2541,N_2080,N_2383);
and U2542 (N_2542,N_2187,N_2492);
nand U2543 (N_2543,N_2353,N_2295);
or U2544 (N_2544,N_2421,N_2009);
nor U2545 (N_2545,N_2382,N_2355);
or U2546 (N_2546,N_2417,N_2321);
and U2547 (N_2547,N_2255,N_2157);
nand U2548 (N_2548,N_2102,N_2343);
nand U2549 (N_2549,N_2362,N_2335);
or U2550 (N_2550,N_2283,N_2357);
nand U2551 (N_2551,N_2078,N_2339);
nor U2552 (N_2552,N_2482,N_2239);
xor U2553 (N_2553,N_2203,N_2142);
or U2554 (N_2554,N_2414,N_2316);
nor U2555 (N_2555,N_2144,N_2206);
and U2556 (N_2556,N_2400,N_2279);
nor U2557 (N_2557,N_2023,N_2322);
xor U2558 (N_2558,N_2106,N_2044);
or U2559 (N_2559,N_2475,N_2222);
nor U2560 (N_2560,N_2099,N_2061);
xor U2561 (N_2561,N_2005,N_2202);
nand U2562 (N_2562,N_2424,N_2312);
and U2563 (N_2563,N_2167,N_2046);
xor U2564 (N_2564,N_2209,N_2342);
nor U2565 (N_2565,N_2432,N_2070);
xnor U2566 (N_2566,N_2120,N_2459);
nor U2567 (N_2567,N_2272,N_2301);
xor U2568 (N_2568,N_2180,N_2347);
xnor U2569 (N_2569,N_2490,N_2007);
xor U2570 (N_2570,N_2373,N_2069);
xnor U2571 (N_2571,N_2384,N_2083);
or U2572 (N_2572,N_2141,N_2025);
nand U2573 (N_2573,N_2089,N_2415);
or U2574 (N_2574,N_2454,N_2457);
nor U2575 (N_2575,N_2496,N_2228);
or U2576 (N_2576,N_2434,N_2299);
and U2577 (N_2577,N_2165,N_2472);
nand U2578 (N_2578,N_2484,N_2168);
nand U2579 (N_2579,N_2131,N_2133);
nand U2580 (N_2580,N_2224,N_2052);
nand U2581 (N_2581,N_2358,N_2267);
nor U2582 (N_2582,N_2470,N_2039);
nor U2583 (N_2583,N_2391,N_2241);
and U2584 (N_2584,N_2060,N_2218);
nand U2585 (N_2585,N_2422,N_2104);
and U2586 (N_2586,N_2092,N_2344);
and U2587 (N_2587,N_2113,N_2211);
or U2588 (N_2588,N_2491,N_2455);
or U2589 (N_2589,N_2116,N_2230);
xor U2590 (N_2590,N_2291,N_2259);
or U2591 (N_2591,N_2161,N_2201);
xor U2592 (N_2592,N_2348,N_2137);
nand U2593 (N_2593,N_2226,N_2341);
nand U2594 (N_2594,N_2266,N_2285);
xor U2595 (N_2595,N_2254,N_2364);
nand U2596 (N_2596,N_2370,N_2433);
nor U2597 (N_2597,N_2000,N_2409);
or U2598 (N_2598,N_2170,N_2444);
or U2599 (N_2599,N_2058,N_2423);
xnor U2600 (N_2600,N_2465,N_2441);
nand U2601 (N_2601,N_2265,N_2041);
and U2602 (N_2602,N_2368,N_2452);
xor U2603 (N_2603,N_2458,N_2297);
or U2604 (N_2604,N_2158,N_2437);
nor U2605 (N_2605,N_2013,N_2003);
and U2606 (N_2606,N_2126,N_2253);
nand U2607 (N_2607,N_2446,N_2185);
nand U2608 (N_2608,N_2225,N_2354);
and U2609 (N_2609,N_2124,N_2050);
nand U2610 (N_2610,N_2175,N_2079);
xnor U2611 (N_2611,N_2350,N_2110);
xor U2612 (N_2612,N_2181,N_2481);
nand U2613 (N_2613,N_2284,N_2489);
xor U2614 (N_2614,N_2453,N_2325);
and U2615 (N_2615,N_2240,N_2396);
nand U2616 (N_2616,N_2351,N_2067);
nor U2617 (N_2617,N_2352,N_2443);
and U2618 (N_2618,N_2498,N_2176);
xnor U2619 (N_2619,N_2395,N_2375);
nand U2620 (N_2620,N_2073,N_2086);
nor U2621 (N_2621,N_2115,N_2411);
nor U2622 (N_2622,N_2336,N_2143);
and U2623 (N_2623,N_2059,N_2327);
or U2624 (N_2624,N_2111,N_2403);
nor U2625 (N_2625,N_2381,N_2091);
nor U2626 (N_2626,N_2030,N_2166);
or U2627 (N_2627,N_2365,N_2314);
nand U2628 (N_2628,N_2223,N_2107);
nor U2629 (N_2629,N_2326,N_2213);
or U2630 (N_2630,N_2026,N_2081);
nor U2631 (N_2631,N_2135,N_2407);
or U2632 (N_2632,N_2497,N_2011);
or U2633 (N_2633,N_2264,N_2393);
nand U2634 (N_2634,N_2191,N_2450);
nor U2635 (N_2635,N_2427,N_2320);
nor U2636 (N_2636,N_2290,N_2129);
or U2637 (N_2637,N_2035,N_2261);
or U2638 (N_2638,N_2460,N_2374);
nor U2639 (N_2639,N_2499,N_2010);
or U2640 (N_2640,N_2132,N_2159);
nand U2641 (N_2641,N_2186,N_2436);
or U2642 (N_2642,N_2055,N_2274);
and U2643 (N_2643,N_2449,N_2094);
xor U2644 (N_2644,N_2269,N_2075);
nand U2645 (N_2645,N_2147,N_2318);
or U2646 (N_2646,N_2298,N_2461);
nand U2647 (N_2647,N_2193,N_2406);
or U2648 (N_2648,N_2262,N_2445);
xor U2649 (N_2649,N_2118,N_2233);
nand U2650 (N_2650,N_2257,N_2172);
or U2651 (N_2651,N_2315,N_2040);
nand U2652 (N_2652,N_2212,N_2271);
or U2653 (N_2653,N_2088,N_2369);
xor U2654 (N_2654,N_2018,N_2333);
nor U2655 (N_2655,N_2287,N_2416);
xnor U2656 (N_2656,N_2156,N_2022);
and U2657 (N_2657,N_2098,N_2273);
nor U2658 (N_2658,N_2379,N_2464);
nand U2659 (N_2659,N_2296,N_2093);
nand U2660 (N_2660,N_2305,N_2425);
xor U2661 (N_2661,N_2085,N_2234);
and U2662 (N_2662,N_2270,N_2012);
nand U2663 (N_2663,N_2317,N_2488);
xnor U2664 (N_2664,N_2447,N_2140);
or U2665 (N_2665,N_2340,N_2471);
nand U2666 (N_2666,N_2431,N_2309);
and U2667 (N_2667,N_2426,N_2268);
nand U2668 (N_2668,N_2275,N_2237);
xnor U2669 (N_2669,N_2281,N_2151);
or U2670 (N_2670,N_2214,N_2439);
nand U2671 (N_2671,N_2243,N_2096);
nor U2672 (N_2672,N_2108,N_2401);
or U2673 (N_2673,N_2020,N_2062);
nand U2674 (N_2674,N_2119,N_2138);
nor U2675 (N_2675,N_2280,N_2200);
or U2676 (N_2676,N_2277,N_2372);
or U2677 (N_2677,N_2331,N_2494);
and U2678 (N_2678,N_2493,N_2256);
and U2679 (N_2679,N_2074,N_2468);
xnor U2680 (N_2680,N_2246,N_2420);
and U2681 (N_2681,N_2178,N_2084);
nor U2682 (N_2682,N_2103,N_2051);
nand U2683 (N_2683,N_2412,N_2288);
or U2684 (N_2684,N_2260,N_2019);
nor U2685 (N_2685,N_2473,N_2389);
nor U2686 (N_2686,N_2386,N_2242);
nor U2687 (N_2687,N_2229,N_2036);
nor U2688 (N_2688,N_2117,N_2235);
nor U2689 (N_2689,N_2419,N_2068);
or U2690 (N_2690,N_2109,N_2462);
nand U2691 (N_2691,N_2049,N_2377);
xor U2692 (N_2692,N_2053,N_2048);
nand U2693 (N_2693,N_2387,N_2408);
xnor U2694 (N_2694,N_2217,N_2205);
xnor U2695 (N_2695,N_2130,N_2349);
or U2696 (N_2696,N_2065,N_2394);
xnor U2697 (N_2697,N_2249,N_2148);
nand U2698 (N_2698,N_2278,N_2430);
and U2699 (N_2699,N_2399,N_2380);
nand U2700 (N_2700,N_2037,N_2438);
nor U2701 (N_2701,N_2304,N_2008);
and U2702 (N_2702,N_2258,N_2442);
or U2703 (N_2703,N_2332,N_2184);
nand U2704 (N_2704,N_2440,N_2043);
nor U2705 (N_2705,N_2478,N_2150);
and U2706 (N_2706,N_2330,N_2014);
nor U2707 (N_2707,N_2038,N_2308);
xor U2708 (N_2708,N_2337,N_2021);
or U2709 (N_2709,N_2282,N_2221);
nand U2710 (N_2710,N_2210,N_2476);
or U2711 (N_2711,N_2346,N_2064);
xor U2712 (N_2712,N_2155,N_2095);
nor U2713 (N_2713,N_2220,N_2047);
nand U2714 (N_2714,N_2028,N_2486);
and U2715 (N_2715,N_2300,N_2194);
or U2716 (N_2716,N_2207,N_2216);
and U2717 (N_2717,N_2121,N_2293);
nor U2718 (N_2718,N_2112,N_2413);
nor U2719 (N_2719,N_2376,N_2323);
and U2720 (N_2720,N_2328,N_2032);
xnor U2721 (N_2721,N_2001,N_2146);
nor U2722 (N_2722,N_2196,N_2072);
nor U2723 (N_2723,N_2154,N_2123);
and U2724 (N_2724,N_2252,N_2153);
nand U2725 (N_2725,N_2145,N_2169);
nand U2726 (N_2726,N_2247,N_2311);
xnor U2727 (N_2727,N_2122,N_2045);
and U2728 (N_2728,N_2136,N_2250);
xnor U2729 (N_2729,N_2017,N_2378);
nand U2730 (N_2730,N_2483,N_2195);
nor U2731 (N_2731,N_2015,N_2236);
nor U2732 (N_2732,N_2474,N_2082);
or U2733 (N_2733,N_2313,N_2429);
xor U2734 (N_2734,N_2485,N_2392);
or U2735 (N_2735,N_2405,N_2361);
nor U2736 (N_2736,N_2363,N_2198);
nor U2737 (N_2737,N_2163,N_2016);
nor U2738 (N_2738,N_2306,N_2398);
nand U2739 (N_2739,N_2397,N_2188);
and U2740 (N_2740,N_2139,N_2033);
xor U2741 (N_2741,N_2087,N_2390);
nand U2742 (N_2742,N_2231,N_2199);
nand U2743 (N_2743,N_2063,N_2366);
or U2744 (N_2744,N_2190,N_2162);
and U2745 (N_2745,N_2367,N_2310);
nand U2746 (N_2746,N_2294,N_2388);
or U2747 (N_2747,N_2251,N_2487);
nand U2748 (N_2748,N_2192,N_2302);
or U2749 (N_2749,N_2338,N_2245);
nand U2750 (N_2750,N_2152,N_2055);
nand U2751 (N_2751,N_2371,N_2306);
xnor U2752 (N_2752,N_2015,N_2104);
nor U2753 (N_2753,N_2291,N_2476);
nand U2754 (N_2754,N_2392,N_2125);
nor U2755 (N_2755,N_2075,N_2438);
nand U2756 (N_2756,N_2127,N_2362);
nand U2757 (N_2757,N_2365,N_2185);
and U2758 (N_2758,N_2354,N_2272);
nor U2759 (N_2759,N_2420,N_2261);
or U2760 (N_2760,N_2049,N_2480);
xor U2761 (N_2761,N_2396,N_2493);
xor U2762 (N_2762,N_2473,N_2333);
or U2763 (N_2763,N_2067,N_2176);
nand U2764 (N_2764,N_2128,N_2075);
or U2765 (N_2765,N_2421,N_2190);
or U2766 (N_2766,N_2266,N_2295);
xnor U2767 (N_2767,N_2076,N_2015);
or U2768 (N_2768,N_2214,N_2404);
nand U2769 (N_2769,N_2241,N_2143);
and U2770 (N_2770,N_2482,N_2407);
nand U2771 (N_2771,N_2218,N_2470);
or U2772 (N_2772,N_2344,N_2094);
xor U2773 (N_2773,N_2374,N_2307);
or U2774 (N_2774,N_2150,N_2402);
xor U2775 (N_2775,N_2279,N_2025);
nor U2776 (N_2776,N_2365,N_2148);
and U2777 (N_2777,N_2384,N_2386);
nor U2778 (N_2778,N_2189,N_2059);
or U2779 (N_2779,N_2209,N_2211);
nor U2780 (N_2780,N_2025,N_2036);
nand U2781 (N_2781,N_2142,N_2215);
nand U2782 (N_2782,N_2078,N_2421);
or U2783 (N_2783,N_2092,N_2212);
xor U2784 (N_2784,N_2458,N_2320);
xor U2785 (N_2785,N_2193,N_2367);
and U2786 (N_2786,N_2249,N_2083);
xnor U2787 (N_2787,N_2361,N_2209);
nand U2788 (N_2788,N_2225,N_2334);
nor U2789 (N_2789,N_2083,N_2345);
or U2790 (N_2790,N_2140,N_2058);
nor U2791 (N_2791,N_2161,N_2335);
nand U2792 (N_2792,N_2021,N_2092);
and U2793 (N_2793,N_2466,N_2026);
xor U2794 (N_2794,N_2420,N_2028);
nor U2795 (N_2795,N_2268,N_2151);
xnor U2796 (N_2796,N_2318,N_2437);
or U2797 (N_2797,N_2281,N_2275);
and U2798 (N_2798,N_2414,N_2447);
nor U2799 (N_2799,N_2407,N_2393);
xnor U2800 (N_2800,N_2304,N_2094);
and U2801 (N_2801,N_2320,N_2254);
nand U2802 (N_2802,N_2252,N_2067);
nor U2803 (N_2803,N_2180,N_2072);
or U2804 (N_2804,N_2453,N_2378);
and U2805 (N_2805,N_2393,N_2421);
or U2806 (N_2806,N_2055,N_2016);
nor U2807 (N_2807,N_2243,N_2301);
and U2808 (N_2808,N_2410,N_2018);
nor U2809 (N_2809,N_2123,N_2465);
xnor U2810 (N_2810,N_2002,N_2006);
nor U2811 (N_2811,N_2112,N_2113);
nand U2812 (N_2812,N_2044,N_2438);
and U2813 (N_2813,N_2405,N_2206);
nor U2814 (N_2814,N_2438,N_2188);
nand U2815 (N_2815,N_2157,N_2047);
nor U2816 (N_2816,N_2268,N_2469);
nand U2817 (N_2817,N_2137,N_2202);
nor U2818 (N_2818,N_2308,N_2193);
nand U2819 (N_2819,N_2233,N_2029);
or U2820 (N_2820,N_2267,N_2466);
or U2821 (N_2821,N_2429,N_2361);
and U2822 (N_2822,N_2445,N_2052);
nand U2823 (N_2823,N_2362,N_2123);
and U2824 (N_2824,N_2473,N_2468);
nor U2825 (N_2825,N_2126,N_2380);
nor U2826 (N_2826,N_2054,N_2194);
or U2827 (N_2827,N_2219,N_2247);
xnor U2828 (N_2828,N_2193,N_2305);
and U2829 (N_2829,N_2231,N_2073);
nor U2830 (N_2830,N_2491,N_2359);
nand U2831 (N_2831,N_2022,N_2470);
nor U2832 (N_2832,N_2379,N_2271);
and U2833 (N_2833,N_2439,N_2279);
nor U2834 (N_2834,N_2194,N_2362);
or U2835 (N_2835,N_2069,N_2473);
or U2836 (N_2836,N_2134,N_2063);
nand U2837 (N_2837,N_2380,N_2362);
and U2838 (N_2838,N_2029,N_2393);
nor U2839 (N_2839,N_2112,N_2471);
or U2840 (N_2840,N_2068,N_2267);
and U2841 (N_2841,N_2172,N_2443);
and U2842 (N_2842,N_2036,N_2348);
or U2843 (N_2843,N_2224,N_2353);
nand U2844 (N_2844,N_2015,N_2344);
or U2845 (N_2845,N_2246,N_2241);
xnor U2846 (N_2846,N_2186,N_2391);
or U2847 (N_2847,N_2409,N_2162);
nor U2848 (N_2848,N_2369,N_2311);
nand U2849 (N_2849,N_2420,N_2328);
nand U2850 (N_2850,N_2115,N_2475);
xor U2851 (N_2851,N_2014,N_2056);
nor U2852 (N_2852,N_2406,N_2414);
or U2853 (N_2853,N_2022,N_2319);
nor U2854 (N_2854,N_2175,N_2463);
or U2855 (N_2855,N_2476,N_2286);
nand U2856 (N_2856,N_2467,N_2328);
nor U2857 (N_2857,N_2046,N_2186);
nand U2858 (N_2858,N_2163,N_2494);
xor U2859 (N_2859,N_2026,N_2266);
xor U2860 (N_2860,N_2331,N_2068);
nand U2861 (N_2861,N_2305,N_2261);
xnor U2862 (N_2862,N_2056,N_2111);
or U2863 (N_2863,N_2148,N_2404);
xnor U2864 (N_2864,N_2452,N_2270);
nor U2865 (N_2865,N_2352,N_2300);
nor U2866 (N_2866,N_2437,N_2238);
or U2867 (N_2867,N_2118,N_2191);
and U2868 (N_2868,N_2194,N_2260);
nor U2869 (N_2869,N_2385,N_2209);
xnor U2870 (N_2870,N_2114,N_2079);
or U2871 (N_2871,N_2321,N_2183);
xor U2872 (N_2872,N_2405,N_2305);
nor U2873 (N_2873,N_2492,N_2347);
or U2874 (N_2874,N_2442,N_2041);
nand U2875 (N_2875,N_2368,N_2420);
and U2876 (N_2876,N_2160,N_2484);
xnor U2877 (N_2877,N_2023,N_2096);
xor U2878 (N_2878,N_2243,N_2394);
nor U2879 (N_2879,N_2238,N_2467);
nor U2880 (N_2880,N_2242,N_2432);
and U2881 (N_2881,N_2446,N_2168);
xor U2882 (N_2882,N_2427,N_2355);
xnor U2883 (N_2883,N_2272,N_2059);
xnor U2884 (N_2884,N_2141,N_2269);
or U2885 (N_2885,N_2382,N_2380);
xor U2886 (N_2886,N_2233,N_2069);
or U2887 (N_2887,N_2146,N_2226);
or U2888 (N_2888,N_2497,N_2352);
nor U2889 (N_2889,N_2272,N_2297);
nand U2890 (N_2890,N_2060,N_2259);
or U2891 (N_2891,N_2320,N_2315);
or U2892 (N_2892,N_2291,N_2300);
or U2893 (N_2893,N_2258,N_2055);
xnor U2894 (N_2894,N_2145,N_2299);
xor U2895 (N_2895,N_2269,N_2000);
and U2896 (N_2896,N_2381,N_2292);
nor U2897 (N_2897,N_2354,N_2416);
nor U2898 (N_2898,N_2403,N_2421);
nand U2899 (N_2899,N_2045,N_2334);
xnor U2900 (N_2900,N_2170,N_2329);
nand U2901 (N_2901,N_2371,N_2112);
nand U2902 (N_2902,N_2228,N_2482);
xor U2903 (N_2903,N_2063,N_2078);
xor U2904 (N_2904,N_2246,N_2012);
or U2905 (N_2905,N_2433,N_2495);
nand U2906 (N_2906,N_2449,N_2378);
or U2907 (N_2907,N_2139,N_2367);
nand U2908 (N_2908,N_2499,N_2196);
xor U2909 (N_2909,N_2126,N_2130);
nor U2910 (N_2910,N_2008,N_2341);
or U2911 (N_2911,N_2354,N_2153);
nand U2912 (N_2912,N_2121,N_2328);
nand U2913 (N_2913,N_2347,N_2292);
and U2914 (N_2914,N_2371,N_2068);
or U2915 (N_2915,N_2430,N_2355);
and U2916 (N_2916,N_2320,N_2243);
xor U2917 (N_2917,N_2043,N_2435);
nor U2918 (N_2918,N_2079,N_2045);
xor U2919 (N_2919,N_2389,N_2114);
xnor U2920 (N_2920,N_2349,N_2362);
xnor U2921 (N_2921,N_2390,N_2494);
nor U2922 (N_2922,N_2466,N_2422);
nand U2923 (N_2923,N_2463,N_2248);
xnor U2924 (N_2924,N_2297,N_2476);
nor U2925 (N_2925,N_2112,N_2149);
xor U2926 (N_2926,N_2331,N_2442);
nor U2927 (N_2927,N_2311,N_2207);
and U2928 (N_2928,N_2088,N_2380);
nand U2929 (N_2929,N_2012,N_2303);
xnor U2930 (N_2930,N_2413,N_2276);
nor U2931 (N_2931,N_2072,N_2232);
nor U2932 (N_2932,N_2127,N_2139);
and U2933 (N_2933,N_2159,N_2215);
and U2934 (N_2934,N_2099,N_2165);
or U2935 (N_2935,N_2128,N_2400);
xor U2936 (N_2936,N_2237,N_2460);
nor U2937 (N_2937,N_2277,N_2338);
xnor U2938 (N_2938,N_2205,N_2227);
nor U2939 (N_2939,N_2237,N_2088);
or U2940 (N_2940,N_2118,N_2262);
nor U2941 (N_2941,N_2086,N_2248);
and U2942 (N_2942,N_2347,N_2384);
and U2943 (N_2943,N_2427,N_2273);
and U2944 (N_2944,N_2209,N_2230);
xor U2945 (N_2945,N_2416,N_2104);
nor U2946 (N_2946,N_2287,N_2146);
nand U2947 (N_2947,N_2039,N_2107);
nand U2948 (N_2948,N_2367,N_2243);
xor U2949 (N_2949,N_2492,N_2260);
and U2950 (N_2950,N_2448,N_2449);
and U2951 (N_2951,N_2083,N_2225);
xor U2952 (N_2952,N_2374,N_2442);
xnor U2953 (N_2953,N_2281,N_2096);
and U2954 (N_2954,N_2463,N_2027);
nand U2955 (N_2955,N_2327,N_2072);
nor U2956 (N_2956,N_2349,N_2087);
xnor U2957 (N_2957,N_2227,N_2368);
xor U2958 (N_2958,N_2292,N_2121);
and U2959 (N_2959,N_2031,N_2332);
nand U2960 (N_2960,N_2386,N_2025);
or U2961 (N_2961,N_2063,N_2032);
or U2962 (N_2962,N_2466,N_2003);
nand U2963 (N_2963,N_2070,N_2328);
nor U2964 (N_2964,N_2485,N_2096);
and U2965 (N_2965,N_2062,N_2014);
and U2966 (N_2966,N_2424,N_2333);
nand U2967 (N_2967,N_2112,N_2467);
xor U2968 (N_2968,N_2082,N_2247);
and U2969 (N_2969,N_2236,N_2314);
nand U2970 (N_2970,N_2135,N_2475);
nand U2971 (N_2971,N_2405,N_2431);
or U2972 (N_2972,N_2146,N_2176);
and U2973 (N_2973,N_2452,N_2493);
nor U2974 (N_2974,N_2419,N_2466);
nor U2975 (N_2975,N_2005,N_2189);
nor U2976 (N_2976,N_2260,N_2127);
xnor U2977 (N_2977,N_2406,N_2429);
or U2978 (N_2978,N_2485,N_2100);
nand U2979 (N_2979,N_2353,N_2350);
nor U2980 (N_2980,N_2424,N_2392);
nand U2981 (N_2981,N_2212,N_2039);
xor U2982 (N_2982,N_2234,N_2369);
or U2983 (N_2983,N_2199,N_2150);
xnor U2984 (N_2984,N_2263,N_2415);
xnor U2985 (N_2985,N_2122,N_2107);
and U2986 (N_2986,N_2423,N_2413);
xor U2987 (N_2987,N_2036,N_2359);
and U2988 (N_2988,N_2109,N_2291);
nor U2989 (N_2989,N_2087,N_2345);
nand U2990 (N_2990,N_2001,N_2275);
nand U2991 (N_2991,N_2320,N_2437);
and U2992 (N_2992,N_2179,N_2030);
or U2993 (N_2993,N_2095,N_2125);
nor U2994 (N_2994,N_2189,N_2092);
and U2995 (N_2995,N_2371,N_2485);
nand U2996 (N_2996,N_2315,N_2252);
and U2997 (N_2997,N_2134,N_2064);
xor U2998 (N_2998,N_2138,N_2025);
and U2999 (N_2999,N_2285,N_2374);
or U3000 (N_3000,N_2586,N_2740);
nor U3001 (N_3001,N_2862,N_2625);
or U3002 (N_3002,N_2764,N_2706);
nand U3003 (N_3003,N_2923,N_2572);
or U3004 (N_3004,N_2555,N_2747);
or U3005 (N_3005,N_2629,N_2989);
nor U3006 (N_3006,N_2860,N_2615);
and U3007 (N_3007,N_2893,N_2504);
nor U3008 (N_3008,N_2818,N_2717);
or U3009 (N_3009,N_2633,N_2506);
nand U3010 (N_3010,N_2929,N_2795);
nand U3011 (N_3011,N_2531,N_2578);
or U3012 (N_3012,N_2925,N_2708);
or U3013 (N_3013,N_2593,N_2533);
xor U3014 (N_3014,N_2933,N_2928);
nor U3015 (N_3015,N_2857,N_2820);
nand U3016 (N_3016,N_2843,N_2725);
or U3017 (N_3017,N_2694,N_2605);
nand U3018 (N_3018,N_2731,N_2516);
xnor U3019 (N_3019,N_2544,N_2879);
xnor U3020 (N_3020,N_2695,N_2597);
and U3021 (N_3021,N_2556,N_2618);
and U3022 (N_3022,N_2664,N_2906);
and U3023 (N_3023,N_2545,N_2554);
and U3024 (N_3024,N_2676,N_2981);
and U3025 (N_3025,N_2998,N_2596);
and U3026 (N_3026,N_2643,N_2965);
or U3027 (N_3027,N_2953,N_2610);
nand U3028 (N_3028,N_2524,N_2546);
or U3029 (N_3029,N_2598,N_2808);
or U3030 (N_3030,N_2767,N_2744);
xor U3031 (N_3031,N_2587,N_2940);
and U3032 (N_3032,N_2541,N_2713);
and U3033 (N_3033,N_2776,N_2865);
xor U3034 (N_3034,N_2873,N_2805);
nor U3035 (N_3035,N_2759,N_2811);
nor U3036 (N_3036,N_2913,N_2992);
nand U3037 (N_3037,N_2727,N_2660);
nand U3038 (N_3038,N_2617,N_2883);
or U3039 (N_3039,N_2966,N_2967);
nor U3040 (N_3040,N_2803,N_2773);
nand U3041 (N_3041,N_2648,N_2963);
xor U3042 (N_3042,N_2716,N_2909);
and U3043 (N_3043,N_2874,N_2737);
nor U3044 (N_3044,N_2920,N_2601);
and U3045 (N_3045,N_2858,N_2631);
xor U3046 (N_3046,N_2709,N_2707);
nor U3047 (N_3047,N_2526,N_2916);
xor U3048 (N_3048,N_2634,N_2749);
nor U3049 (N_3049,N_2688,N_2842);
xor U3050 (N_3050,N_2885,N_2936);
and U3051 (N_3051,N_2964,N_2557);
xor U3052 (N_3052,N_2856,N_2897);
nand U3053 (N_3053,N_2500,N_2658);
and U3054 (N_3054,N_2907,N_2792);
xnor U3055 (N_3055,N_2612,N_2765);
or U3056 (N_3056,N_2525,N_2815);
nand U3057 (N_3057,N_2974,N_2917);
nor U3058 (N_3058,N_2642,N_2594);
nor U3059 (N_3059,N_2637,N_2548);
or U3060 (N_3060,N_2960,N_2774);
or U3061 (N_3061,N_2882,N_2821);
xor U3062 (N_3062,N_2589,N_2576);
xor U3063 (N_3063,N_2997,N_2715);
and U3064 (N_3064,N_2949,N_2881);
or U3065 (N_3065,N_2793,N_2761);
or U3066 (N_3066,N_2835,N_2538);
nor U3067 (N_3067,N_2507,N_2990);
and U3068 (N_3068,N_2509,N_2653);
xnor U3069 (N_3069,N_2654,N_2791);
nand U3070 (N_3070,N_2668,N_2646);
xnor U3071 (N_3071,N_2922,N_2978);
and U3072 (N_3072,N_2914,N_2743);
and U3073 (N_3073,N_2899,N_2769);
nor U3074 (N_3074,N_2732,N_2563);
xnor U3075 (N_3075,N_2638,N_2799);
xor U3076 (N_3076,N_2956,N_2512);
nand U3077 (N_3077,N_2838,N_2673);
and U3078 (N_3078,N_2867,N_2996);
or U3079 (N_3079,N_2816,N_2937);
nor U3080 (N_3080,N_2574,N_2700);
and U3081 (N_3081,N_2891,N_2861);
xor U3082 (N_3082,N_2809,N_2942);
and U3083 (N_3083,N_2698,N_2851);
or U3084 (N_3084,N_2840,N_2918);
or U3085 (N_3085,N_2896,N_2846);
or U3086 (N_3086,N_2505,N_2943);
nand U3087 (N_3087,N_2566,N_2845);
nand U3088 (N_3088,N_2650,N_2611);
or U3089 (N_3089,N_2961,N_2588);
and U3090 (N_3090,N_2626,N_2827);
nor U3091 (N_3091,N_2868,N_2542);
or U3092 (N_3092,N_2549,N_2983);
nor U3093 (N_3093,N_2718,N_2995);
nand U3094 (N_3094,N_2518,N_2550);
and U3095 (N_3095,N_2647,N_2508);
xnor U3096 (N_3096,N_2817,N_2705);
or U3097 (N_3097,N_2592,N_2780);
or U3098 (N_3098,N_2620,N_2609);
or U3099 (N_3099,N_2924,N_2517);
xor U3100 (N_3100,N_2781,N_2575);
nor U3101 (N_3101,N_2750,N_2675);
or U3102 (N_3102,N_2639,N_2704);
or U3103 (N_3103,N_2947,N_2714);
and U3104 (N_3104,N_2567,N_2502);
and U3105 (N_3105,N_2934,N_2655);
nor U3106 (N_3106,N_2553,N_2685);
nor U3107 (N_3107,N_2739,N_2969);
or U3108 (N_3108,N_2600,N_2682);
xnor U3109 (N_3109,N_2959,N_2813);
and U3110 (N_3110,N_2733,N_2863);
nor U3111 (N_3111,N_2900,N_2772);
xnor U3112 (N_3112,N_2841,N_2683);
or U3113 (N_3113,N_2726,N_2958);
nor U3114 (N_3114,N_2875,N_2738);
and U3115 (N_3115,N_2910,N_2833);
nor U3116 (N_3116,N_2831,N_2926);
xor U3117 (N_3117,N_2822,N_2890);
nand U3118 (N_3118,N_2614,N_2754);
xor U3119 (N_3119,N_2748,N_2537);
or U3120 (N_3120,N_2692,N_2806);
or U3121 (N_3121,N_2849,N_2939);
nor U3122 (N_3122,N_2884,N_2919);
and U3123 (N_3123,N_2562,N_2573);
and U3124 (N_3124,N_2880,N_2606);
xor U3125 (N_3125,N_2693,N_2935);
and U3126 (N_3126,N_2689,N_2886);
and U3127 (N_3127,N_2973,N_2657);
xor U3128 (N_3128,N_2632,N_2972);
nand U3129 (N_3129,N_2641,N_2870);
or U3130 (N_3130,N_2510,N_2666);
or U3131 (N_3131,N_2837,N_2665);
nor U3132 (N_3132,N_2786,N_2762);
and U3133 (N_3133,N_2911,N_2902);
and U3134 (N_3134,N_2898,N_2591);
nand U3135 (N_3135,N_2640,N_2677);
and U3136 (N_3136,N_2814,N_2832);
xnor U3137 (N_3137,N_2853,N_2932);
nand U3138 (N_3138,N_2830,N_2607);
or U3139 (N_3139,N_2741,N_2703);
nor U3140 (N_3140,N_2825,N_2687);
or U3141 (N_3141,N_2946,N_2904);
nand U3142 (N_3142,N_2968,N_2728);
or U3143 (N_3143,N_2812,N_2515);
nor U3144 (N_3144,N_2790,N_2794);
nand U3145 (N_3145,N_2590,N_2871);
or U3146 (N_3146,N_2941,N_2608);
nand U3147 (N_3147,N_2690,N_2752);
nand U3148 (N_3148,N_2905,N_2771);
nand U3149 (N_3149,N_2604,N_2571);
nor U3150 (N_3150,N_2945,N_2635);
and U3151 (N_3151,N_2735,N_2944);
and U3152 (N_3152,N_2672,N_2568);
nand U3153 (N_3153,N_2669,N_2696);
or U3154 (N_3154,N_2957,N_2616);
nor U3155 (N_3155,N_2684,N_2595);
nor U3156 (N_3156,N_2511,N_2852);
nor U3157 (N_3157,N_2577,N_2745);
and U3158 (N_3158,N_2987,N_2921);
nand U3159 (N_3159,N_2547,N_2603);
nand U3160 (N_3160,N_2864,N_2982);
nor U3161 (N_3161,N_2519,N_2746);
xnor U3162 (N_3162,N_2915,N_2804);
and U3163 (N_3163,N_2580,N_2686);
nor U3164 (N_3164,N_2829,N_2532);
nand U3165 (N_3165,N_2661,N_2892);
nand U3166 (N_3166,N_2579,N_2520);
xor U3167 (N_3167,N_2513,N_2758);
and U3168 (N_3168,N_2994,N_2980);
and U3169 (N_3169,N_2866,N_2583);
nand U3170 (N_3170,N_2938,N_2670);
xnor U3171 (N_3171,N_2988,N_2766);
nand U3172 (N_3172,N_2659,N_2539);
or U3173 (N_3173,N_2736,N_2662);
nor U3174 (N_3174,N_2787,N_2819);
xnor U3175 (N_3175,N_2889,N_2826);
or U3176 (N_3176,N_2619,N_2798);
and U3177 (N_3177,N_2878,N_2775);
or U3178 (N_3178,N_2564,N_2777);
and U3179 (N_3179,N_2763,N_2561);
xor U3180 (N_3180,N_2622,N_2970);
xnor U3181 (N_3181,N_2742,N_2651);
nand U3182 (N_3182,N_2894,N_2710);
nor U3183 (N_3183,N_2801,N_2636);
and U3184 (N_3184,N_2644,N_2678);
xor U3185 (N_3185,N_2971,N_2521);
nand U3186 (N_3186,N_2663,N_2950);
xnor U3187 (N_3187,N_2999,N_2702);
xnor U3188 (N_3188,N_2697,N_2681);
and U3189 (N_3189,N_2755,N_2584);
xnor U3190 (N_3190,N_2789,N_2784);
xor U3191 (N_3191,N_2797,N_2802);
xor U3192 (N_3192,N_2530,N_2711);
nor U3193 (N_3193,N_2975,N_2523);
nand U3194 (N_3194,N_2770,N_2854);
nand U3195 (N_3195,N_2788,N_2514);
or U3196 (N_3196,N_2667,N_2834);
or U3197 (N_3197,N_2585,N_2800);
nor U3198 (N_3198,N_2543,N_2985);
nor U3199 (N_3199,N_2501,N_2536);
nor U3200 (N_3200,N_2552,N_2721);
or U3201 (N_3201,N_2720,N_2551);
xor U3202 (N_3202,N_2522,N_2701);
nand U3203 (N_3203,N_2903,N_2569);
xor U3204 (N_3204,N_2652,N_2691);
or U3205 (N_3205,N_2824,N_2602);
nand U3206 (N_3206,N_2850,N_2570);
xnor U3207 (N_3207,N_2984,N_2847);
and U3208 (N_3208,N_2869,N_2779);
nor U3209 (N_3209,N_2722,N_2699);
xor U3210 (N_3210,N_2859,N_2581);
nand U3211 (N_3211,N_2529,N_2734);
nor U3212 (N_3212,N_2599,N_2778);
nor U3213 (N_3213,N_2855,N_2623);
nor U3214 (N_3214,N_2872,N_2807);
xor U3215 (N_3215,N_2844,N_2785);
or U3216 (N_3216,N_2558,N_2559);
xnor U3217 (N_3217,N_2680,N_2931);
nor U3218 (N_3218,N_2712,N_2540);
and U3219 (N_3219,N_2565,N_2671);
or U3220 (N_3220,N_2991,N_2630);
or U3221 (N_3221,N_2534,N_2848);
and U3222 (N_3222,N_2979,N_2901);
xor U3223 (N_3223,N_2757,N_2783);
nand U3224 (N_3224,N_2962,N_2503);
nor U3225 (N_3225,N_2954,N_2895);
and U3226 (N_3226,N_2823,N_2912);
and U3227 (N_3227,N_2977,N_2723);
or U3228 (N_3228,N_2951,N_2887);
nand U3229 (N_3229,N_2724,N_2753);
nand U3230 (N_3230,N_2927,N_2930);
or U3231 (N_3231,N_2955,N_2876);
or U3232 (N_3232,N_2810,N_2952);
xor U3233 (N_3233,N_2624,N_2760);
nand U3234 (N_3234,N_2679,N_2782);
and U3235 (N_3235,N_2751,N_2986);
and U3236 (N_3236,N_2674,N_2527);
xnor U3237 (N_3237,N_2976,N_2993);
nor U3238 (N_3238,N_2560,N_2828);
and U3239 (N_3239,N_2730,N_2908);
nand U3240 (N_3240,N_2796,N_2582);
xor U3241 (N_3241,N_2768,N_2888);
nor U3242 (N_3242,N_2948,N_2621);
and U3243 (N_3243,N_2627,N_2839);
or U3244 (N_3244,N_2649,N_2613);
nor U3245 (N_3245,N_2656,N_2756);
or U3246 (N_3246,N_2628,N_2528);
nor U3247 (N_3247,N_2836,N_2729);
xor U3248 (N_3248,N_2877,N_2535);
nand U3249 (N_3249,N_2645,N_2719);
nand U3250 (N_3250,N_2605,N_2765);
xnor U3251 (N_3251,N_2513,N_2695);
or U3252 (N_3252,N_2581,N_2564);
nand U3253 (N_3253,N_2907,N_2611);
nand U3254 (N_3254,N_2690,N_2786);
nand U3255 (N_3255,N_2742,N_2519);
nor U3256 (N_3256,N_2517,N_2992);
xor U3257 (N_3257,N_2595,N_2993);
or U3258 (N_3258,N_2835,N_2522);
and U3259 (N_3259,N_2523,N_2599);
nor U3260 (N_3260,N_2696,N_2661);
xnor U3261 (N_3261,N_2741,N_2679);
xnor U3262 (N_3262,N_2816,N_2558);
nand U3263 (N_3263,N_2645,N_2794);
nand U3264 (N_3264,N_2944,N_2910);
xor U3265 (N_3265,N_2970,N_2828);
nand U3266 (N_3266,N_2596,N_2875);
nor U3267 (N_3267,N_2820,N_2543);
and U3268 (N_3268,N_2569,N_2728);
and U3269 (N_3269,N_2952,N_2702);
or U3270 (N_3270,N_2720,N_2666);
nor U3271 (N_3271,N_2617,N_2793);
or U3272 (N_3272,N_2829,N_2558);
nand U3273 (N_3273,N_2744,N_2935);
and U3274 (N_3274,N_2813,N_2628);
or U3275 (N_3275,N_2748,N_2659);
nand U3276 (N_3276,N_2735,N_2701);
and U3277 (N_3277,N_2852,N_2831);
xor U3278 (N_3278,N_2951,N_2681);
nor U3279 (N_3279,N_2966,N_2535);
nor U3280 (N_3280,N_2705,N_2620);
and U3281 (N_3281,N_2913,N_2806);
nor U3282 (N_3282,N_2695,N_2632);
and U3283 (N_3283,N_2562,N_2695);
and U3284 (N_3284,N_2795,N_2810);
nand U3285 (N_3285,N_2805,N_2863);
or U3286 (N_3286,N_2608,N_2528);
xor U3287 (N_3287,N_2790,N_2600);
nor U3288 (N_3288,N_2615,N_2600);
or U3289 (N_3289,N_2980,N_2662);
nand U3290 (N_3290,N_2842,N_2738);
nand U3291 (N_3291,N_2992,N_2745);
or U3292 (N_3292,N_2580,N_2955);
nand U3293 (N_3293,N_2692,N_2830);
nand U3294 (N_3294,N_2675,N_2509);
xor U3295 (N_3295,N_2903,N_2619);
xor U3296 (N_3296,N_2770,N_2896);
or U3297 (N_3297,N_2507,N_2806);
or U3298 (N_3298,N_2984,N_2747);
or U3299 (N_3299,N_2926,N_2951);
and U3300 (N_3300,N_2589,N_2725);
or U3301 (N_3301,N_2615,N_2653);
or U3302 (N_3302,N_2565,N_2632);
nor U3303 (N_3303,N_2624,N_2931);
xor U3304 (N_3304,N_2775,N_2614);
nand U3305 (N_3305,N_2786,N_2511);
nand U3306 (N_3306,N_2610,N_2829);
xor U3307 (N_3307,N_2859,N_2914);
xnor U3308 (N_3308,N_2670,N_2787);
and U3309 (N_3309,N_2968,N_2567);
or U3310 (N_3310,N_2848,N_2556);
xnor U3311 (N_3311,N_2704,N_2742);
xnor U3312 (N_3312,N_2614,N_2780);
or U3313 (N_3313,N_2824,N_2702);
nor U3314 (N_3314,N_2604,N_2594);
nand U3315 (N_3315,N_2688,N_2548);
nand U3316 (N_3316,N_2536,N_2650);
nand U3317 (N_3317,N_2667,N_2848);
xnor U3318 (N_3318,N_2794,N_2682);
nand U3319 (N_3319,N_2750,N_2819);
xnor U3320 (N_3320,N_2772,N_2790);
and U3321 (N_3321,N_2532,N_2508);
nand U3322 (N_3322,N_2885,N_2577);
nand U3323 (N_3323,N_2925,N_2513);
nor U3324 (N_3324,N_2504,N_2859);
or U3325 (N_3325,N_2961,N_2977);
nor U3326 (N_3326,N_2783,N_2500);
nor U3327 (N_3327,N_2720,N_2898);
and U3328 (N_3328,N_2618,N_2538);
nand U3329 (N_3329,N_2620,N_2702);
and U3330 (N_3330,N_2742,N_2555);
and U3331 (N_3331,N_2836,N_2811);
xor U3332 (N_3332,N_2809,N_2981);
nor U3333 (N_3333,N_2690,N_2771);
nand U3334 (N_3334,N_2719,N_2631);
or U3335 (N_3335,N_2767,N_2676);
nor U3336 (N_3336,N_2750,N_2656);
nor U3337 (N_3337,N_2718,N_2997);
or U3338 (N_3338,N_2660,N_2910);
xor U3339 (N_3339,N_2569,N_2584);
or U3340 (N_3340,N_2739,N_2560);
nor U3341 (N_3341,N_2837,N_2780);
xor U3342 (N_3342,N_2934,N_2710);
and U3343 (N_3343,N_2908,N_2651);
nand U3344 (N_3344,N_2601,N_2562);
and U3345 (N_3345,N_2587,N_2523);
or U3346 (N_3346,N_2554,N_2581);
xor U3347 (N_3347,N_2886,N_2990);
nor U3348 (N_3348,N_2521,N_2894);
nor U3349 (N_3349,N_2890,N_2971);
xor U3350 (N_3350,N_2642,N_2529);
nand U3351 (N_3351,N_2916,N_2724);
and U3352 (N_3352,N_2594,N_2600);
nor U3353 (N_3353,N_2738,N_2853);
nand U3354 (N_3354,N_2728,N_2578);
and U3355 (N_3355,N_2958,N_2725);
nor U3356 (N_3356,N_2870,N_2884);
nor U3357 (N_3357,N_2706,N_2538);
and U3358 (N_3358,N_2552,N_2642);
or U3359 (N_3359,N_2675,N_2555);
nand U3360 (N_3360,N_2988,N_2943);
and U3361 (N_3361,N_2965,N_2713);
or U3362 (N_3362,N_2605,N_2592);
nand U3363 (N_3363,N_2902,N_2869);
nor U3364 (N_3364,N_2598,N_2561);
nor U3365 (N_3365,N_2860,N_2637);
xnor U3366 (N_3366,N_2830,N_2962);
nand U3367 (N_3367,N_2534,N_2931);
nand U3368 (N_3368,N_2583,N_2765);
nor U3369 (N_3369,N_2883,N_2650);
or U3370 (N_3370,N_2521,N_2582);
xor U3371 (N_3371,N_2524,N_2613);
or U3372 (N_3372,N_2976,N_2908);
nand U3373 (N_3373,N_2705,N_2720);
nand U3374 (N_3374,N_2953,N_2895);
and U3375 (N_3375,N_2713,N_2740);
or U3376 (N_3376,N_2603,N_2717);
nor U3377 (N_3377,N_2823,N_2870);
xor U3378 (N_3378,N_2699,N_2620);
and U3379 (N_3379,N_2876,N_2644);
nor U3380 (N_3380,N_2648,N_2851);
nand U3381 (N_3381,N_2535,N_2612);
xnor U3382 (N_3382,N_2502,N_2528);
nor U3383 (N_3383,N_2986,N_2649);
and U3384 (N_3384,N_2964,N_2620);
and U3385 (N_3385,N_2958,N_2786);
and U3386 (N_3386,N_2997,N_2714);
or U3387 (N_3387,N_2727,N_2693);
nor U3388 (N_3388,N_2990,N_2986);
xor U3389 (N_3389,N_2879,N_2792);
nor U3390 (N_3390,N_2912,N_2861);
nor U3391 (N_3391,N_2598,N_2984);
and U3392 (N_3392,N_2724,N_2679);
xnor U3393 (N_3393,N_2915,N_2916);
or U3394 (N_3394,N_2893,N_2723);
nor U3395 (N_3395,N_2756,N_2543);
nand U3396 (N_3396,N_2951,N_2925);
and U3397 (N_3397,N_2572,N_2790);
xor U3398 (N_3398,N_2929,N_2607);
xnor U3399 (N_3399,N_2610,N_2653);
nor U3400 (N_3400,N_2668,N_2731);
and U3401 (N_3401,N_2807,N_2567);
xor U3402 (N_3402,N_2564,N_2654);
xor U3403 (N_3403,N_2829,N_2504);
or U3404 (N_3404,N_2508,N_2863);
nor U3405 (N_3405,N_2960,N_2742);
or U3406 (N_3406,N_2620,N_2565);
nand U3407 (N_3407,N_2580,N_2930);
nand U3408 (N_3408,N_2877,N_2686);
and U3409 (N_3409,N_2632,N_2591);
xnor U3410 (N_3410,N_2827,N_2532);
nand U3411 (N_3411,N_2886,N_2641);
or U3412 (N_3412,N_2738,N_2921);
nand U3413 (N_3413,N_2719,N_2941);
or U3414 (N_3414,N_2544,N_2981);
or U3415 (N_3415,N_2885,N_2723);
nor U3416 (N_3416,N_2798,N_2713);
nand U3417 (N_3417,N_2536,N_2775);
and U3418 (N_3418,N_2636,N_2682);
and U3419 (N_3419,N_2825,N_2933);
xnor U3420 (N_3420,N_2606,N_2923);
xor U3421 (N_3421,N_2800,N_2983);
or U3422 (N_3422,N_2561,N_2647);
nor U3423 (N_3423,N_2596,N_2558);
nand U3424 (N_3424,N_2631,N_2630);
and U3425 (N_3425,N_2586,N_2541);
nor U3426 (N_3426,N_2649,N_2980);
xnor U3427 (N_3427,N_2885,N_2654);
nor U3428 (N_3428,N_2566,N_2814);
nor U3429 (N_3429,N_2881,N_2781);
and U3430 (N_3430,N_2555,N_2922);
nor U3431 (N_3431,N_2726,N_2545);
or U3432 (N_3432,N_2652,N_2702);
and U3433 (N_3433,N_2812,N_2974);
or U3434 (N_3434,N_2717,N_2963);
and U3435 (N_3435,N_2600,N_2533);
or U3436 (N_3436,N_2991,N_2542);
and U3437 (N_3437,N_2732,N_2753);
nor U3438 (N_3438,N_2751,N_2725);
xor U3439 (N_3439,N_2519,N_2723);
nand U3440 (N_3440,N_2751,N_2684);
and U3441 (N_3441,N_2830,N_2533);
nand U3442 (N_3442,N_2514,N_2970);
or U3443 (N_3443,N_2581,N_2660);
nor U3444 (N_3444,N_2660,N_2563);
and U3445 (N_3445,N_2651,N_2841);
nor U3446 (N_3446,N_2657,N_2735);
xnor U3447 (N_3447,N_2849,N_2846);
and U3448 (N_3448,N_2527,N_2868);
or U3449 (N_3449,N_2545,N_2977);
nand U3450 (N_3450,N_2844,N_2575);
and U3451 (N_3451,N_2809,N_2819);
nor U3452 (N_3452,N_2877,N_2523);
nor U3453 (N_3453,N_2588,N_2558);
nor U3454 (N_3454,N_2516,N_2528);
and U3455 (N_3455,N_2765,N_2696);
nand U3456 (N_3456,N_2518,N_2622);
nor U3457 (N_3457,N_2767,N_2701);
nor U3458 (N_3458,N_2780,N_2713);
and U3459 (N_3459,N_2931,N_2516);
or U3460 (N_3460,N_2640,N_2631);
nand U3461 (N_3461,N_2765,N_2592);
nand U3462 (N_3462,N_2522,N_2774);
xor U3463 (N_3463,N_2737,N_2844);
nor U3464 (N_3464,N_2914,N_2603);
nor U3465 (N_3465,N_2698,N_2819);
xnor U3466 (N_3466,N_2742,N_2845);
nor U3467 (N_3467,N_2928,N_2609);
and U3468 (N_3468,N_2786,N_2917);
nor U3469 (N_3469,N_2789,N_2991);
and U3470 (N_3470,N_2928,N_2611);
and U3471 (N_3471,N_2664,N_2781);
and U3472 (N_3472,N_2507,N_2587);
or U3473 (N_3473,N_2755,N_2564);
nor U3474 (N_3474,N_2666,N_2531);
and U3475 (N_3475,N_2557,N_2613);
and U3476 (N_3476,N_2785,N_2819);
and U3477 (N_3477,N_2770,N_2735);
or U3478 (N_3478,N_2977,N_2935);
nor U3479 (N_3479,N_2638,N_2649);
xnor U3480 (N_3480,N_2555,N_2519);
nor U3481 (N_3481,N_2783,N_2646);
nand U3482 (N_3482,N_2977,N_2531);
xor U3483 (N_3483,N_2935,N_2900);
xnor U3484 (N_3484,N_2900,N_2742);
xor U3485 (N_3485,N_2851,N_2700);
and U3486 (N_3486,N_2577,N_2762);
xnor U3487 (N_3487,N_2733,N_2728);
or U3488 (N_3488,N_2627,N_2864);
nand U3489 (N_3489,N_2919,N_2846);
nand U3490 (N_3490,N_2819,N_2649);
nand U3491 (N_3491,N_2760,N_2752);
xor U3492 (N_3492,N_2909,N_2867);
or U3493 (N_3493,N_2796,N_2671);
or U3494 (N_3494,N_2799,N_2947);
and U3495 (N_3495,N_2644,N_2672);
nor U3496 (N_3496,N_2707,N_2548);
xor U3497 (N_3497,N_2510,N_2934);
or U3498 (N_3498,N_2814,N_2766);
and U3499 (N_3499,N_2946,N_2783);
nand U3500 (N_3500,N_3437,N_3238);
and U3501 (N_3501,N_3129,N_3454);
nor U3502 (N_3502,N_3003,N_3269);
xnor U3503 (N_3503,N_3015,N_3205);
or U3504 (N_3504,N_3194,N_3117);
xnor U3505 (N_3505,N_3250,N_3039);
nor U3506 (N_3506,N_3209,N_3315);
xnor U3507 (N_3507,N_3064,N_3285);
and U3508 (N_3508,N_3466,N_3057);
or U3509 (N_3509,N_3183,N_3195);
and U3510 (N_3510,N_3027,N_3332);
xnor U3511 (N_3511,N_3000,N_3331);
xor U3512 (N_3512,N_3424,N_3125);
nor U3513 (N_3513,N_3002,N_3499);
xor U3514 (N_3514,N_3381,N_3029);
nor U3515 (N_3515,N_3407,N_3274);
xor U3516 (N_3516,N_3028,N_3386);
nor U3517 (N_3517,N_3107,N_3410);
nor U3518 (N_3518,N_3305,N_3357);
nand U3519 (N_3519,N_3334,N_3236);
xnor U3520 (N_3520,N_3151,N_3382);
nor U3521 (N_3521,N_3435,N_3438);
or U3522 (N_3522,N_3323,N_3110);
xor U3523 (N_3523,N_3477,N_3088);
and U3524 (N_3524,N_3380,N_3019);
or U3525 (N_3525,N_3047,N_3384);
nand U3526 (N_3526,N_3218,N_3358);
xor U3527 (N_3527,N_3145,N_3493);
nand U3528 (N_3528,N_3237,N_3496);
and U3529 (N_3529,N_3230,N_3364);
nor U3530 (N_3530,N_3257,N_3051);
and U3531 (N_3531,N_3127,N_3313);
and U3532 (N_3532,N_3378,N_3228);
and U3533 (N_3533,N_3263,N_3174);
xnor U3534 (N_3534,N_3076,N_3402);
nor U3535 (N_3535,N_3337,N_3389);
nand U3536 (N_3536,N_3494,N_3373);
nand U3537 (N_3537,N_3128,N_3404);
nand U3538 (N_3538,N_3137,N_3460);
or U3539 (N_3539,N_3343,N_3231);
nor U3540 (N_3540,N_3401,N_3159);
nor U3541 (N_3541,N_3246,N_3254);
nor U3542 (N_3542,N_3295,N_3397);
and U3543 (N_3543,N_3054,N_3310);
nand U3544 (N_3544,N_3041,N_3249);
nor U3545 (N_3545,N_3006,N_3255);
nor U3546 (N_3546,N_3468,N_3045);
and U3547 (N_3547,N_3324,N_3072);
nor U3548 (N_3548,N_3363,N_3316);
or U3549 (N_3549,N_3105,N_3393);
or U3550 (N_3550,N_3467,N_3166);
and U3551 (N_3551,N_3241,N_3154);
xor U3552 (N_3552,N_3396,N_3068);
and U3553 (N_3553,N_3414,N_3175);
nand U3554 (N_3554,N_3208,N_3232);
xnor U3555 (N_3555,N_3244,N_3248);
nor U3556 (N_3556,N_3115,N_3116);
nand U3557 (N_3557,N_3239,N_3063);
xor U3558 (N_3558,N_3060,N_3318);
and U3559 (N_3559,N_3187,N_3261);
nor U3560 (N_3560,N_3355,N_3066);
nor U3561 (N_3561,N_3476,N_3018);
xor U3562 (N_3562,N_3158,N_3283);
nor U3563 (N_3563,N_3044,N_3413);
or U3564 (N_3564,N_3480,N_3036);
or U3565 (N_3565,N_3356,N_3299);
nand U3566 (N_3566,N_3368,N_3472);
or U3567 (N_3567,N_3266,N_3059);
or U3568 (N_3568,N_3056,N_3233);
nor U3569 (N_3569,N_3433,N_3012);
nor U3570 (N_3570,N_3383,N_3312);
nand U3571 (N_3571,N_3021,N_3138);
xnor U3572 (N_3572,N_3052,N_3459);
xor U3573 (N_3573,N_3284,N_3037);
nand U3574 (N_3574,N_3446,N_3449);
nand U3575 (N_3575,N_3270,N_3394);
nand U3576 (N_3576,N_3227,N_3286);
xor U3577 (N_3577,N_3014,N_3023);
or U3578 (N_3578,N_3176,N_3149);
nor U3579 (N_3579,N_3418,N_3069);
nand U3580 (N_3580,N_3217,N_3490);
xnor U3581 (N_3581,N_3092,N_3247);
xor U3582 (N_3582,N_3017,N_3173);
nand U3583 (N_3583,N_3294,N_3349);
nand U3584 (N_3584,N_3055,N_3091);
nand U3585 (N_3585,N_3366,N_3111);
and U3586 (N_3586,N_3053,N_3262);
or U3587 (N_3587,N_3361,N_3048);
or U3588 (N_3588,N_3197,N_3081);
nand U3589 (N_3589,N_3234,N_3156);
xnor U3590 (N_3590,N_3367,N_3279);
nor U3591 (N_3591,N_3082,N_3181);
or U3592 (N_3592,N_3010,N_3399);
or U3593 (N_3593,N_3497,N_3296);
or U3594 (N_3594,N_3353,N_3415);
xnor U3595 (N_3595,N_3009,N_3345);
or U3596 (N_3596,N_3034,N_3202);
nor U3597 (N_3597,N_3222,N_3350);
xnor U3598 (N_3598,N_3152,N_3462);
nand U3599 (N_3599,N_3346,N_3097);
or U3600 (N_3600,N_3013,N_3276);
nand U3601 (N_3601,N_3142,N_3405);
nor U3602 (N_3602,N_3471,N_3201);
nand U3603 (N_3603,N_3083,N_3409);
and U3604 (N_3604,N_3292,N_3336);
nor U3605 (N_3605,N_3426,N_3192);
and U3606 (N_3606,N_3443,N_3163);
or U3607 (N_3607,N_3133,N_3180);
xnor U3608 (N_3608,N_3224,N_3320);
nand U3609 (N_3609,N_3379,N_3431);
nand U3610 (N_3610,N_3008,N_3385);
and U3611 (N_3611,N_3134,N_3422);
or U3612 (N_3612,N_3483,N_3432);
and U3613 (N_3613,N_3419,N_3155);
nand U3614 (N_3614,N_3141,N_3165);
xnor U3615 (N_3615,N_3297,N_3425);
and U3616 (N_3616,N_3475,N_3179);
nor U3617 (N_3617,N_3440,N_3289);
nor U3618 (N_3618,N_3136,N_3408);
xnor U3619 (N_3619,N_3147,N_3428);
and U3620 (N_3620,N_3188,N_3022);
nand U3621 (N_3621,N_3321,N_3311);
xor U3622 (N_3622,N_3120,N_3464);
xnor U3623 (N_3623,N_3333,N_3168);
and U3624 (N_3624,N_3280,N_3093);
nand U3625 (N_3625,N_3338,N_3293);
or U3626 (N_3626,N_3245,N_3445);
nand U3627 (N_3627,N_3075,N_3342);
nand U3628 (N_3628,N_3043,N_3328);
nor U3629 (N_3629,N_3112,N_3096);
or U3630 (N_3630,N_3287,N_3359);
nor U3631 (N_3631,N_3164,N_3114);
xnor U3632 (N_3632,N_3388,N_3146);
and U3633 (N_3633,N_3077,N_3211);
or U3634 (N_3634,N_3061,N_3278);
xor U3635 (N_3635,N_3025,N_3203);
or U3636 (N_3636,N_3453,N_3186);
xor U3637 (N_3637,N_3212,N_3090);
nor U3638 (N_3638,N_3423,N_3348);
xnor U3639 (N_3639,N_3360,N_3122);
xnor U3640 (N_3640,N_3387,N_3371);
xnor U3641 (N_3641,N_3220,N_3032);
or U3642 (N_3642,N_3492,N_3160);
nand U3643 (N_3643,N_3272,N_3302);
nor U3644 (N_3644,N_3079,N_3474);
nor U3645 (N_3645,N_3420,N_3121);
nand U3646 (N_3646,N_3307,N_3259);
xor U3647 (N_3647,N_3215,N_3298);
nand U3648 (N_3648,N_3450,N_3461);
nand U3649 (N_3649,N_3268,N_3135);
xnor U3650 (N_3650,N_3304,N_3495);
and U3651 (N_3651,N_3240,N_3369);
or U3652 (N_3652,N_3339,N_3126);
xor U3653 (N_3653,N_3016,N_3065);
nand U3654 (N_3654,N_3265,N_3277);
xor U3655 (N_3655,N_3235,N_3098);
and U3656 (N_3656,N_3322,N_3223);
nand U3657 (N_3657,N_3103,N_3275);
nor U3658 (N_3658,N_3335,N_3319);
xor U3659 (N_3659,N_3071,N_3119);
or U3660 (N_3660,N_3398,N_3001);
or U3661 (N_3661,N_3300,N_3271);
and U3662 (N_3662,N_3131,N_3007);
and U3663 (N_3663,N_3229,N_3221);
or U3664 (N_3664,N_3099,N_3441);
nand U3665 (N_3665,N_3049,N_3282);
and U3666 (N_3666,N_3153,N_3078);
xnor U3667 (N_3667,N_3488,N_3258);
nand U3668 (N_3668,N_3487,N_3354);
or U3669 (N_3669,N_3470,N_3340);
xnor U3670 (N_3670,N_3108,N_3171);
nor U3671 (N_3671,N_3486,N_3370);
nor U3672 (N_3672,N_3484,N_3144);
and U3673 (N_3673,N_3252,N_3291);
and U3674 (N_3674,N_3411,N_3273);
and U3675 (N_3675,N_3498,N_3113);
xnor U3676 (N_3676,N_3463,N_3458);
nand U3677 (N_3677,N_3004,N_3362);
and U3678 (N_3678,N_3478,N_3104);
xor U3679 (N_3679,N_3086,N_3465);
nor U3680 (N_3680,N_3352,N_3177);
and U3681 (N_3681,N_3200,N_3281);
nor U3682 (N_3682,N_3301,N_3434);
nand U3683 (N_3683,N_3395,N_3406);
nor U3684 (N_3684,N_3011,N_3143);
or U3685 (N_3685,N_3344,N_3062);
and U3686 (N_3686,N_3172,N_3020);
xor U3687 (N_3687,N_3429,N_3267);
and U3688 (N_3688,N_3089,N_3288);
nor U3689 (N_3689,N_3306,N_3489);
xor U3690 (N_3690,N_3417,N_3167);
and U3691 (N_3691,N_3225,N_3102);
nor U3692 (N_3692,N_3412,N_3216);
or U3693 (N_3693,N_3095,N_3341);
nor U3694 (N_3694,N_3376,N_3226);
nand U3695 (N_3695,N_3193,N_3213);
or U3696 (N_3696,N_3189,N_3132);
and U3697 (N_3697,N_3005,N_3150);
nor U3698 (N_3698,N_3094,N_3198);
xor U3699 (N_3699,N_3439,N_3100);
or U3700 (N_3700,N_3067,N_3325);
nor U3701 (N_3701,N_3253,N_3469);
xor U3702 (N_3702,N_3491,N_3451);
nand U3703 (N_3703,N_3481,N_3196);
and U3704 (N_3704,N_3400,N_3442);
and U3705 (N_3705,N_3214,N_3184);
and U3706 (N_3706,N_3421,N_3485);
or U3707 (N_3707,N_3042,N_3087);
or U3708 (N_3708,N_3124,N_3084);
and U3709 (N_3709,N_3207,N_3085);
xor U3710 (N_3710,N_3264,N_3448);
xor U3711 (N_3711,N_3427,N_3130);
nor U3712 (N_3712,N_3219,N_3375);
and U3713 (N_3713,N_3330,N_3243);
or U3714 (N_3714,N_3482,N_3457);
xnor U3715 (N_3715,N_3351,N_3372);
xor U3716 (N_3716,N_3473,N_3050);
xnor U3717 (N_3717,N_3178,N_3317);
and U3718 (N_3718,N_3191,N_3073);
and U3719 (N_3719,N_3308,N_3392);
or U3720 (N_3720,N_3455,N_3026);
and U3721 (N_3721,N_3190,N_3242);
and U3722 (N_3722,N_3080,N_3038);
nor U3723 (N_3723,N_3260,N_3140);
and U3724 (N_3724,N_3040,N_3290);
xor U3725 (N_3725,N_3447,N_3403);
xnor U3726 (N_3726,N_3101,N_3327);
nand U3727 (N_3727,N_3162,N_3416);
and U3728 (N_3728,N_3148,N_3479);
nor U3729 (N_3729,N_3206,N_3185);
nand U3730 (N_3730,N_3374,N_3182);
xor U3731 (N_3731,N_3430,N_3161);
or U3732 (N_3732,N_3070,N_3391);
xnor U3733 (N_3733,N_3390,N_3118);
or U3734 (N_3734,N_3139,N_3030);
xnor U3735 (N_3735,N_3106,N_3074);
or U3736 (N_3736,N_3347,N_3309);
or U3737 (N_3737,N_3251,N_3436);
xor U3738 (N_3738,N_3199,N_3326);
nor U3739 (N_3739,N_3444,N_3329);
and U3740 (N_3740,N_3314,N_3169);
nand U3741 (N_3741,N_3031,N_3256);
or U3742 (N_3742,N_3123,N_3204);
and U3743 (N_3743,N_3210,N_3303);
and U3744 (N_3744,N_3024,N_3170);
xor U3745 (N_3745,N_3157,N_3377);
or U3746 (N_3746,N_3109,N_3033);
xor U3747 (N_3747,N_3058,N_3035);
nand U3748 (N_3748,N_3452,N_3365);
nor U3749 (N_3749,N_3456,N_3046);
xnor U3750 (N_3750,N_3119,N_3035);
and U3751 (N_3751,N_3417,N_3232);
nand U3752 (N_3752,N_3486,N_3440);
xnor U3753 (N_3753,N_3117,N_3115);
nor U3754 (N_3754,N_3403,N_3268);
nand U3755 (N_3755,N_3279,N_3335);
or U3756 (N_3756,N_3081,N_3259);
nand U3757 (N_3757,N_3413,N_3333);
nor U3758 (N_3758,N_3400,N_3444);
nor U3759 (N_3759,N_3407,N_3442);
or U3760 (N_3760,N_3420,N_3070);
or U3761 (N_3761,N_3117,N_3060);
nor U3762 (N_3762,N_3047,N_3203);
nand U3763 (N_3763,N_3324,N_3435);
xnor U3764 (N_3764,N_3167,N_3155);
xor U3765 (N_3765,N_3094,N_3484);
nand U3766 (N_3766,N_3061,N_3024);
and U3767 (N_3767,N_3310,N_3227);
and U3768 (N_3768,N_3136,N_3433);
nor U3769 (N_3769,N_3214,N_3362);
nor U3770 (N_3770,N_3008,N_3232);
nand U3771 (N_3771,N_3181,N_3136);
nand U3772 (N_3772,N_3449,N_3189);
nand U3773 (N_3773,N_3463,N_3416);
or U3774 (N_3774,N_3252,N_3212);
xnor U3775 (N_3775,N_3137,N_3255);
or U3776 (N_3776,N_3186,N_3098);
nor U3777 (N_3777,N_3331,N_3214);
or U3778 (N_3778,N_3127,N_3475);
xor U3779 (N_3779,N_3105,N_3404);
or U3780 (N_3780,N_3016,N_3337);
or U3781 (N_3781,N_3073,N_3093);
or U3782 (N_3782,N_3361,N_3430);
and U3783 (N_3783,N_3479,N_3333);
and U3784 (N_3784,N_3072,N_3197);
and U3785 (N_3785,N_3060,N_3215);
and U3786 (N_3786,N_3365,N_3352);
xnor U3787 (N_3787,N_3156,N_3327);
xor U3788 (N_3788,N_3270,N_3482);
nand U3789 (N_3789,N_3016,N_3116);
or U3790 (N_3790,N_3238,N_3287);
xor U3791 (N_3791,N_3352,N_3208);
nand U3792 (N_3792,N_3214,N_3175);
and U3793 (N_3793,N_3073,N_3454);
and U3794 (N_3794,N_3117,N_3292);
xnor U3795 (N_3795,N_3171,N_3283);
and U3796 (N_3796,N_3118,N_3329);
xor U3797 (N_3797,N_3485,N_3321);
or U3798 (N_3798,N_3165,N_3091);
or U3799 (N_3799,N_3300,N_3463);
or U3800 (N_3800,N_3061,N_3377);
xor U3801 (N_3801,N_3359,N_3185);
or U3802 (N_3802,N_3059,N_3103);
and U3803 (N_3803,N_3123,N_3000);
nor U3804 (N_3804,N_3192,N_3305);
nand U3805 (N_3805,N_3126,N_3276);
xor U3806 (N_3806,N_3345,N_3266);
or U3807 (N_3807,N_3177,N_3244);
nor U3808 (N_3808,N_3165,N_3458);
and U3809 (N_3809,N_3404,N_3354);
nor U3810 (N_3810,N_3309,N_3279);
nor U3811 (N_3811,N_3099,N_3276);
and U3812 (N_3812,N_3071,N_3384);
nor U3813 (N_3813,N_3023,N_3219);
nor U3814 (N_3814,N_3174,N_3115);
and U3815 (N_3815,N_3098,N_3032);
and U3816 (N_3816,N_3387,N_3017);
nor U3817 (N_3817,N_3438,N_3280);
nor U3818 (N_3818,N_3010,N_3126);
nor U3819 (N_3819,N_3486,N_3476);
nand U3820 (N_3820,N_3307,N_3269);
nor U3821 (N_3821,N_3200,N_3187);
or U3822 (N_3822,N_3402,N_3174);
nand U3823 (N_3823,N_3274,N_3469);
nor U3824 (N_3824,N_3261,N_3025);
xor U3825 (N_3825,N_3124,N_3129);
and U3826 (N_3826,N_3393,N_3187);
xor U3827 (N_3827,N_3396,N_3373);
nor U3828 (N_3828,N_3069,N_3491);
nor U3829 (N_3829,N_3370,N_3329);
nand U3830 (N_3830,N_3197,N_3135);
nand U3831 (N_3831,N_3108,N_3413);
and U3832 (N_3832,N_3276,N_3263);
nor U3833 (N_3833,N_3349,N_3005);
xor U3834 (N_3834,N_3266,N_3242);
and U3835 (N_3835,N_3019,N_3472);
xor U3836 (N_3836,N_3431,N_3149);
or U3837 (N_3837,N_3341,N_3000);
xor U3838 (N_3838,N_3119,N_3425);
and U3839 (N_3839,N_3006,N_3438);
or U3840 (N_3840,N_3380,N_3212);
and U3841 (N_3841,N_3380,N_3162);
or U3842 (N_3842,N_3067,N_3373);
xor U3843 (N_3843,N_3230,N_3333);
nand U3844 (N_3844,N_3384,N_3278);
and U3845 (N_3845,N_3080,N_3007);
and U3846 (N_3846,N_3100,N_3026);
nand U3847 (N_3847,N_3401,N_3000);
and U3848 (N_3848,N_3421,N_3198);
and U3849 (N_3849,N_3167,N_3177);
nand U3850 (N_3850,N_3493,N_3034);
nand U3851 (N_3851,N_3001,N_3241);
and U3852 (N_3852,N_3450,N_3267);
or U3853 (N_3853,N_3358,N_3122);
or U3854 (N_3854,N_3039,N_3355);
nand U3855 (N_3855,N_3249,N_3438);
nor U3856 (N_3856,N_3131,N_3382);
or U3857 (N_3857,N_3364,N_3481);
nor U3858 (N_3858,N_3183,N_3317);
and U3859 (N_3859,N_3254,N_3088);
nand U3860 (N_3860,N_3202,N_3261);
nand U3861 (N_3861,N_3084,N_3310);
nand U3862 (N_3862,N_3371,N_3460);
xnor U3863 (N_3863,N_3276,N_3249);
nor U3864 (N_3864,N_3474,N_3471);
and U3865 (N_3865,N_3071,N_3131);
or U3866 (N_3866,N_3256,N_3070);
and U3867 (N_3867,N_3101,N_3185);
xnor U3868 (N_3868,N_3290,N_3410);
or U3869 (N_3869,N_3305,N_3042);
nor U3870 (N_3870,N_3265,N_3337);
nand U3871 (N_3871,N_3451,N_3042);
and U3872 (N_3872,N_3247,N_3165);
nor U3873 (N_3873,N_3278,N_3093);
xnor U3874 (N_3874,N_3480,N_3013);
and U3875 (N_3875,N_3439,N_3151);
xor U3876 (N_3876,N_3284,N_3351);
or U3877 (N_3877,N_3320,N_3116);
nand U3878 (N_3878,N_3252,N_3287);
and U3879 (N_3879,N_3368,N_3270);
or U3880 (N_3880,N_3123,N_3245);
nor U3881 (N_3881,N_3149,N_3225);
nor U3882 (N_3882,N_3266,N_3308);
or U3883 (N_3883,N_3045,N_3025);
nand U3884 (N_3884,N_3170,N_3195);
and U3885 (N_3885,N_3406,N_3418);
nand U3886 (N_3886,N_3452,N_3189);
or U3887 (N_3887,N_3062,N_3054);
nand U3888 (N_3888,N_3163,N_3149);
or U3889 (N_3889,N_3134,N_3116);
nor U3890 (N_3890,N_3262,N_3122);
and U3891 (N_3891,N_3020,N_3347);
or U3892 (N_3892,N_3055,N_3311);
or U3893 (N_3893,N_3309,N_3144);
xor U3894 (N_3894,N_3166,N_3365);
or U3895 (N_3895,N_3131,N_3362);
nand U3896 (N_3896,N_3094,N_3017);
xor U3897 (N_3897,N_3074,N_3038);
nand U3898 (N_3898,N_3365,N_3312);
nand U3899 (N_3899,N_3338,N_3084);
nor U3900 (N_3900,N_3371,N_3152);
or U3901 (N_3901,N_3431,N_3483);
nand U3902 (N_3902,N_3375,N_3389);
xor U3903 (N_3903,N_3070,N_3122);
nor U3904 (N_3904,N_3425,N_3106);
nor U3905 (N_3905,N_3373,N_3044);
nand U3906 (N_3906,N_3394,N_3213);
xnor U3907 (N_3907,N_3445,N_3135);
and U3908 (N_3908,N_3273,N_3356);
nand U3909 (N_3909,N_3146,N_3123);
and U3910 (N_3910,N_3022,N_3078);
or U3911 (N_3911,N_3425,N_3096);
and U3912 (N_3912,N_3389,N_3045);
xor U3913 (N_3913,N_3488,N_3459);
or U3914 (N_3914,N_3154,N_3191);
and U3915 (N_3915,N_3416,N_3168);
nor U3916 (N_3916,N_3007,N_3479);
or U3917 (N_3917,N_3198,N_3372);
and U3918 (N_3918,N_3013,N_3397);
or U3919 (N_3919,N_3158,N_3439);
nor U3920 (N_3920,N_3001,N_3441);
or U3921 (N_3921,N_3354,N_3158);
nand U3922 (N_3922,N_3196,N_3472);
or U3923 (N_3923,N_3438,N_3109);
xor U3924 (N_3924,N_3436,N_3481);
and U3925 (N_3925,N_3478,N_3248);
nand U3926 (N_3926,N_3309,N_3245);
and U3927 (N_3927,N_3066,N_3140);
or U3928 (N_3928,N_3360,N_3182);
and U3929 (N_3929,N_3389,N_3124);
nor U3930 (N_3930,N_3299,N_3481);
nand U3931 (N_3931,N_3165,N_3308);
nand U3932 (N_3932,N_3178,N_3125);
nand U3933 (N_3933,N_3078,N_3027);
and U3934 (N_3934,N_3000,N_3023);
xor U3935 (N_3935,N_3365,N_3369);
and U3936 (N_3936,N_3488,N_3388);
nand U3937 (N_3937,N_3336,N_3082);
or U3938 (N_3938,N_3087,N_3226);
and U3939 (N_3939,N_3032,N_3472);
xnor U3940 (N_3940,N_3127,N_3067);
nand U3941 (N_3941,N_3174,N_3342);
or U3942 (N_3942,N_3341,N_3035);
xor U3943 (N_3943,N_3000,N_3004);
nor U3944 (N_3944,N_3434,N_3249);
or U3945 (N_3945,N_3305,N_3472);
xor U3946 (N_3946,N_3015,N_3233);
nor U3947 (N_3947,N_3226,N_3496);
or U3948 (N_3948,N_3254,N_3104);
or U3949 (N_3949,N_3153,N_3312);
or U3950 (N_3950,N_3008,N_3015);
or U3951 (N_3951,N_3387,N_3031);
nand U3952 (N_3952,N_3201,N_3374);
nor U3953 (N_3953,N_3470,N_3473);
xor U3954 (N_3954,N_3119,N_3432);
and U3955 (N_3955,N_3210,N_3491);
or U3956 (N_3956,N_3466,N_3079);
nor U3957 (N_3957,N_3344,N_3127);
and U3958 (N_3958,N_3201,N_3308);
xor U3959 (N_3959,N_3409,N_3263);
nand U3960 (N_3960,N_3154,N_3326);
and U3961 (N_3961,N_3188,N_3181);
nor U3962 (N_3962,N_3152,N_3085);
xor U3963 (N_3963,N_3125,N_3071);
nor U3964 (N_3964,N_3285,N_3268);
nor U3965 (N_3965,N_3358,N_3091);
nor U3966 (N_3966,N_3031,N_3428);
and U3967 (N_3967,N_3005,N_3296);
and U3968 (N_3968,N_3130,N_3485);
or U3969 (N_3969,N_3271,N_3245);
or U3970 (N_3970,N_3268,N_3023);
nand U3971 (N_3971,N_3235,N_3490);
and U3972 (N_3972,N_3333,N_3119);
or U3973 (N_3973,N_3195,N_3161);
and U3974 (N_3974,N_3142,N_3198);
nor U3975 (N_3975,N_3321,N_3223);
and U3976 (N_3976,N_3228,N_3184);
and U3977 (N_3977,N_3125,N_3404);
nor U3978 (N_3978,N_3035,N_3001);
and U3979 (N_3979,N_3415,N_3093);
nand U3980 (N_3980,N_3461,N_3225);
or U3981 (N_3981,N_3121,N_3313);
and U3982 (N_3982,N_3429,N_3417);
nand U3983 (N_3983,N_3257,N_3080);
nand U3984 (N_3984,N_3245,N_3436);
or U3985 (N_3985,N_3089,N_3079);
nor U3986 (N_3986,N_3268,N_3161);
nand U3987 (N_3987,N_3442,N_3061);
nor U3988 (N_3988,N_3326,N_3318);
and U3989 (N_3989,N_3031,N_3349);
nand U3990 (N_3990,N_3405,N_3010);
xnor U3991 (N_3991,N_3317,N_3198);
and U3992 (N_3992,N_3193,N_3377);
or U3993 (N_3993,N_3003,N_3407);
and U3994 (N_3994,N_3130,N_3309);
nand U3995 (N_3995,N_3318,N_3270);
or U3996 (N_3996,N_3174,N_3233);
xor U3997 (N_3997,N_3166,N_3111);
nor U3998 (N_3998,N_3179,N_3329);
and U3999 (N_3999,N_3209,N_3069);
nand U4000 (N_4000,N_3794,N_3762);
or U4001 (N_4001,N_3609,N_3728);
nor U4002 (N_4002,N_3770,N_3937);
nand U4003 (N_4003,N_3997,N_3556);
xnor U4004 (N_4004,N_3536,N_3540);
xor U4005 (N_4005,N_3827,N_3961);
nand U4006 (N_4006,N_3968,N_3605);
xnor U4007 (N_4007,N_3682,N_3923);
nand U4008 (N_4008,N_3644,N_3700);
or U4009 (N_4009,N_3980,N_3962);
nor U4010 (N_4010,N_3763,N_3843);
xnor U4011 (N_4011,N_3876,N_3552);
xor U4012 (N_4012,N_3965,N_3883);
nand U4013 (N_4013,N_3721,N_3732);
xor U4014 (N_4014,N_3621,N_3839);
nor U4015 (N_4015,N_3982,N_3510);
nand U4016 (N_4016,N_3956,N_3767);
nor U4017 (N_4017,N_3882,N_3852);
or U4018 (N_4018,N_3888,N_3511);
nor U4019 (N_4019,N_3822,N_3769);
xnor U4020 (N_4020,N_3850,N_3869);
nor U4021 (N_4021,N_3713,N_3719);
or U4022 (N_4022,N_3651,N_3655);
and U4023 (N_4023,N_3571,N_3683);
nand U4024 (N_4024,N_3572,N_3625);
or U4025 (N_4025,N_3542,N_3668);
xnor U4026 (N_4026,N_3570,N_3630);
and U4027 (N_4027,N_3771,N_3518);
or U4028 (N_4028,N_3674,N_3875);
xor U4029 (N_4029,N_3847,N_3975);
and U4030 (N_4030,N_3910,N_3684);
xor U4031 (N_4031,N_3949,N_3753);
and U4032 (N_4032,N_3596,N_3972);
nand U4033 (N_4033,N_3585,N_3877);
nor U4034 (N_4034,N_3659,N_3969);
nand U4035 (N_4035,N_3742,N_3614);
nand U4036 (N_4036,N_3941,N_3787);
nand U4037 (N_4037,N_3564,N_3685);
or U4038 (N_4038,N_3523,N_3879);
or U4039 (N_4039,N_3546,N_3608);
nor U4040 (N_4040,N_3835,N_3681);
nand U4041 (N_4041,N_3884,N_3782);
xnor U4042 (N_4042,N_3637,N_3958);
nand U4043 (N_4043,N_3559,N_3967);
and U4044 (N_4044,N_3749,N_3993);
or U4045 (N_4045,N_3801,N_3901);
nand U4046 (N_4046,N_3873,N_3976);
xnor U4047 (N_4047,N_3567,N_3579);
nor U4048 (N_4048,N_3663,N_3952);
and U4049 (N_4049,N_3508,N_3823);
and U4050 (N_4050,N_3887,N_3768);
or U4051 (N_4051,N_3588,N_3754);
nor U4052 (N_4052,N_3954,N_3560);
and U4053 (N_4053,N_3731,N_3670);
or U4054 (N_4054,N_3631,N_3791);
xnor U4055 (N_4055,N_3589,N_3955);
or U4056 (N_4056,N_3927,N_3701);
and U4057 (N_4057,N_3706,N_3551);
nor U4058 (N_4058,N_3680,N_3624);
or U4059 (N_4059,N_3851,N_3730);
nor U4060 (N_4060,N_3999,N_3601);
or U4061 (N_4061,N_3964,N_3756);
nor U4062 (N_4062,N_3722,N_3909);
nor U4063 (N_4063,N_3626,N_3963);
nor U4064 (N_4064,N_3897,N_3533);
xnor U4065 (N_4065,N_3598,N_3603);
and U4066 (N_4066,N_3988,N_3917);
and U4067 (N_4067,N_3618,N_3842);
xnor U4068 (N_4068,N_3830,N_3765);
or U4069 (N_4069,N_3583,N_3678);
xnor U4070 (N_4070,N_3566,N_3720);
nand U4071 (N_4071,N_3779,N_3959);
xnor U4072 (N_4072,N_3613,N_3513);
xnor U4073 (N_4073,N_3845,N_3520);
and U4074 (N_4074,N_3790,N_3703);
xnor U4075 (N_4075,N_3857,N_3783);
or U4076 (N_4076,N_3718,N_3544);
nor U4077 (N_4077,N_3899,N_3619);
nor U4078 (N_4078,N_3848,N_3858);
or U4079 (N_4079,N_3810,N_3643);
and U4080 (N_4080,N_3995,N_3724);
or U4081 (N_4081,N_3911,N_3886);
nand U4082 (N_4082,N_3504,N_3778);
nor U4083 (N_4083,N_3951,N_3555);
nand U4084 (N_4084,N_3506,N_3737);
xnor U4085 (N_4085,N_3657,N_3940);
nor U4086 (N_4086,N_3890,N_3781);
and U4087 (N_4087,N_3814,N_3934);
or U4088 (N_4088,N_3872,N_3931);
xor U4089 (N_4089,N_3758,N_3832);
nand U4090 (N_4090,N_3634,N_3977);
and U4091 (N_4091,N_3824,N_3880);
nor U4092 (N_4092,N_3574,N_3831);
nor U4093 (N_4093,N_3776,N_3948);
and U4094 (N_4094,N_3528,N_3697);
xor U4095 (N_4095,N_3562,N_3970);
and U4096 (N_4096,N_3541,N_3777);
xnor U4097 (N_4097,N_3966,N_3727);
and U4098 (N_4098,N_3930,N_3702);
xor U4099 (N_4099,N_3519,N_3517);
or U4100 (N_4100,N_3532,N_3622);
nand U4101 (N_4101,N_3645,N_3512);
nor U4102 (N_4102,N_3994,N_3535);
or U4103 (N_4103,N_3616,N_3531);
xnor U4104 (N_4104,N_3925,N_3591);
nand U4105 (N_4105,N_3628,N_3974);
nor U4106 (N_4106,N_3792,N_3525);
and U4107 (N_4107,N_3597,N_3677);
nand U4108 (N_4108,N_3904,N_3650);
and U4109 (N_4109,N_3807,N_3895);
nor U4110 (N_4110,N_3748,N_3602);
nor U4111 (N_4111,N_3840,N_3635);
and U4112 (N_4112,N_3632,N_3662);
or U4113 (N_4113,N_3775,N_3979);
and U4114 (N_4114,N_3928,N_3543);
xnor U4115 (N_4115,N_3660,N_3836);
xor U4116 (N_4116,N_3906,N_3735);
or U4117 (N_4117,N_3766,N_3759);
and U4118 (N_4118,N_3921,N_3607);
xor U4119 (N_4119,N_3793,N_3649);
or U4120 (N_4120,N_3696,N_3726);
nand U4121 (N_4121,N_3889,N_3675);
or U4122 (N_4122,N_3561,N_3798);
nor U4123 (N_4123,N_3739,N_3648);
and U4124 (N_4124,N_3711,N_3529);
nor U4125 (N_4125,N_3623,N_3576);
nand U4126 (N_4126,N_3557,N_3580);
xor U4127 (N_4127,N_3745,N_3933);
xor U4128 (N_4128,N_3755,N_3802);
and U4129 (N_4129,N_3865,N_3587);
xnor U4130 (N_4130,N_3757,N_3919);
nor U4131 (N_4131,N_3834,N_3859);
or U4132 (N_4132,N_3803,N_3673);
or U4133 (N_4133,N_3825,N_3907);
and U4134 (N_4134,N_3939,N_3725);
or U4135 (N_4135,N_3584,N_3945);
nor U4136 (N_4136,N_3938,N_3554);
and U4137 (N_4137,N_3600,N_3691);
or U4138 (N_4138,N_3690,N_3590);
nand U4139 (N_4139,N_3699,N_3837);
xnor U4140 (N_4140,N_3985,N_3669);
nor U4141 (N_4141,N_3741,N_3522);
nor U4142 (N_4142,N_3990,N_3687);
or U4143 (N_4143,N_3971,N_3764);
or U4144 (N_4144,N_3599,N_3550);
xor U4145 (N_4145,N_3606,N_3861);
nor U4146 (N_4146,N_3563,N_3582);
nand U4147 (N_4147,N_3944,N_3878);
nor U4148 (N_4148,N_3929,N_3874);
nor U4149 (N_4149,N_3553,N_3558);
nor U4150 (N_4150,N_3548,N_3900);
or U4151 (N_4151,N_3867,N_3996);
nand U4152 (N_4152,N_3604,N_3885);
nor U4153 (N_4153,N_3908,N_3960);
nand U4154 (N_4154,N_3549,N_3692);
nor U4155 (N_4155,N_3534,N_3545);
nor U4156 (N_4156,N_3918,N_3978);
or U4157 (N_4157,N_3914,N_3983);
xor U4158 (N_4158,N_3710,N_3615);
or U4159 (N_4159,N_3640,N_3734);
xnor U4160 (N_4160,N_3676,N_3866);
nor U4161 (N_4161,N_3672,N_3568);
xor U4162 (N_4162,N_3515,N_3503);
or U4163 (N_4163,N_3594,N_3661);
nor U4164 (N_4164,N_3821,N_3805);
and U4165 (N_4165,N_3828,N_3986);
or U4166 (N_4166,N_3786,N_3813);
nor U4167 (N_4167,N_3653,N_3569);
nor U4168 (N_4168,N_3577,N_3844);
nand U4169 (N_4169,N_3505,N_3863);
or U4170 (N_4170,N_3774,N_3947);
xor U4171 (N_4171,N_3811,N_3855);
nor U4172 (N_4172,N_3924,N_3829);
nor U4173 (N_4173,N_3707,N_3521);
or U4174 (N_4174,N_3809,N_3633);
xor U4175 (N_4175,N_3526,N_3723);
nor U4176 (N_4176,N_3665,N_3989);
and U4177 (N_4177,N_3629,N_3679);
nor U4178 (N_4178,N_3627,N_3815);
nor U4179 (N_4179,N_3750,N_3743);
nor U4180 (N_4180,N_3800,N_3816);
nor U4181 (N_4181,N_3581,N_3573);
nand U4182 (N_4182,N_3870,N_3729);
xnor U4183 (N_4183,N_3751,N_3705);
nor U4184 (N_4184,N_3891,N_3981);
and U4185 (N_4185,N_3991,N_3746);
and U4186 (N_4186,N_3666,N_3507);
and U4187 (N_4187,N_3892,N_3785);
xor U4188 (N_4188,N_3654,N_3538);
nor U4189 (N_4189,N_3853,N_3820);
nor U4190 (N_4190,N_3826,N_3760);
xnor U4191 (N_4191,N_3698,N_3838);
nand U4192 (N_4192,N_3943,N_3902);
xnor U4193 (N_4193,N_3922,N_3856);
xnor U4194 (N_4194,N_3799,N_3935);
xnor U4195 (N_4195,N_3846,N_3854);
xnor U4196 (N_4196,N_3733,N_3984);
xnor U4197 (N_4197,N_3514,N_3689);
nand U4198 (N_4198,N_3841,N_3936);
nor U4199 (N_4199,N_3987,N_3860);
and U4200 (N_4200,N_3780,N_3772);
xnor U4201 (N_4201,N_3740,N_3881);
xnor U4202 (N_4202,N_3957,N_3864);
and U4203 (N_4203,N_3804,N_3736);
nor U4204 (N_4204,N_3942,N_3915);
or U4205 (N_4205,N_3788,N_3642);
xor U4206 (N_4206,N_3905,N_3638);
or U4207 (N_4207,N_3752,N_3586);
or U4208 (N_4208,N_3671,N_3695);
and U4209 (N_4209,N_3647,N_3524);
nor U4210 (N_4210,N_3694,N_3639);
nor U4211 (N_4211,N_3819,N_3620);
or U4212 (N_4212,N_3652,N_3871);
or U4213 (N_4213,N_3537,N_3656);
nor U4214 (N_4214,N_3950,N_3527);
nor U4215 (N_4215,N_3516,N_3708);
and U4216 (N_4216,N_3797,N_3808);
nand U4217 (N_4217,N_3578,N_3973);
xor U4218 (N_4218,N_3913,N_3611);
xor U4219 (N_4219,N_3920,N_3693);
nand U4220 (N_4220,N_3773,N_3500);
nor U4221 (N_4221,N_3501,N_3946);
xor U4222 (N_4222,N_3894,N_3789);
xor U4223 (N_4223,N_3761,N_3916);
or U4224 (N_4224,N_3714,N_3998);
nand U4225 (N_4225,N_3646,N_3795);
xor U4226 (N_4226,N_3738,N_3992);
nand U4227 (N_4227,N_3784,N_3747);
xnor U4228 (N_4228,N_3565,N_3593);
and U4229 (N_4229,N_3664,N_3658);
and U4230 (N_4230,N_3812,N_3641);
nor U4231 (N_4231,N_3817,N_3667);
or U4232 (N_4232,N_3893,N_3539);
nand U4233 (N_4233,N_3862,N_3712);
or U4234 (N_4234,N_3688,N_3595);
nor U4235 (N_4235,N_3704,N_3868);
or U4236 (N_4236,N_3898,N_3592);
and U4237 (N_4237,N_3806,N_3575);
and U4238 (N_4238,N_3715,N_3612);
nand U4239 (N_4239,N_3932,N_3953);
xnor U4240 (N_4240,N_3716,N_3547);
or U4241 (N_4241,N_3896,N_3849);
or U4242 (N_4242,N_3530,N_3912);
xor U4243 (N_4243,N_3833,N_3796);
xnor U4244 (N_4244,N_3926,N_3903);
nor U4245 (N_4245,N_3617,N_3717);
and U4246 (N_4246,N_3818,N_3744);
xnor U4247 (N_4247,N_3509,N_3686);
nand U4248 (N_4248,N_3636,N_3610);
xnor U4249 (N_4249,N_3502,N_3709);
nand U4250 (N_4250,N_3961,N_3720);
nor U4251 (N_4251,N_3876,N_3778);
xnor U4252 (N_4252,N_3812,N_3620);
nand U4253 (N_4253,N_3830,N_3600);
xor U4254 (N_4254,N_3576,N_3625);
nand U4255 (N_4255,N_3543,N_3583);
xor U4256 (N_4256,N_3776,N_3500);
nor U4257 (N_4257,N_3520,N_3868);
and U4258 (N_4258,N_3784,N_3998);
and U4259 (N_4259,N_3575,N_3785);
nor U4260 (N_4260,N_3763,N_3717);
and U4261 (N_4261,N_3992,N_3683);
nor U4262 (N_4262,N_3936,N_3993);
or U4263 (N_4263,N_3812,N_3957);
nor U4264 (N_4264,N_3995,N_3645);
and U4265 (N_4265,N_3766,N_3675);
nand U4266 (N_4266,N_3707,N_3919);
nand U4267 (N_4267,N_3621,N_3790);
nand U4268 (N_4268,N_3923,N_3509);
nor U4269 (N_4269,N_3641,N_3961);
xor U4270 (N_4270,N_3696,N_3693);
nand U4271 (N_4271,N_3696,N_3671);
or U4272 (N_4272,N_3952,N_3628);
nor U4273 (N_4273,N_3588,N_3928);
and U4274 (N_4274,N_3722,N_3966);
and U4275 (N_4275,N_3504,N_3673);
nand U4276 (N_4276,N_3673,N_3669);
and U4277 (N_4277,N_3553,N_3755);
or U4278 (N_4278,N_3975,N_3923);
nand U4279 (N_4279,N_3656,N_3979);
and U4280 (N_4280,N_3614,N_3683);
nor U4281 (N_4281,N_3500,N_3816);
xor U4282 (N_4282,N_3594,N_3552);
nor U4283 (N_4283,N_3613,N_3587);
nand U4284 (N_4284,N_3892,N_3805);
and U4285 (N_4285,N_3696,N_3674);
and U4286 (N_4286,N_3630,N_3998);
and U4287 (N_4287,N_3529,N_3584);
and U4288 (N_4288,N_3881,N_3914);
xor U4289 (N_4289,N_3773,N_3545);
or U4290 (N_4290,N_3959,N_3575);
nor U4291 (N_4291,N_3587,N_3606);
or U4292 (N_4292,N_3799,N_3841);
and U4293 (N_4293,N_3865,N_3533);
nand U4294 (N_4294,N_3886,N_3664);
xor U4295 (N_4295,N_3840,N_3581);
xor U4296 (N_4296,N_3574,N_3930);
nor U4297 (N_4297,N_3557,N_3739);
nor U4298 (N_4298,N_3834,N_3713);
nor U4299 (N_4299,N_3573,N_3709);
nand U4300 (N_4300,N_3604,N_3587);
nand U4301 (N_4301,N_3973,N_3591);
nor U4302 (N_4302,N_3975,N_3636);
and U4303 (N_4303,N_3703,N_3903);
nand U4304 (N_4304,N_3604,N_3869);
and U4305 (N_4305,N_3680,N_3736);
or U4306 (N_4306,N_3649,N_3822);
nand U4307 (N_4307,N_3884,N_3579);
nand U4308 (N_4308,N_3524,N_3755);
nor U4309 (N_4309,N_3855,N_3655);
nand U4310 (N_4310,N_3544,N_3571);
nand U4311 (N_4311,N_3505,N_3585);
and U4312 (N_4312,N_3630,N_3857);
or U4313 (N_4313,N_3707,N_3827);
xor U4314 (N_4314,N_3536,N_3524);
xnor U4315 (N_4315,N_3727,N_3811);
and U4316 (N_4316,N_3608,N_3670);
nand U4317 (N_4317,N_3712,N_3692);
xnor U4318 (N_4318,N_3513,N_3741);
nor U4319 (N_4319,N_3815,N_3908);
nand U4320 (N_4320,N_3631,N_3567);
or U4321 (N_4321,N_3765,N_3806);
nor U4322 (N_4322,N_3850,N_3727);
xnor U4323 (N_4323,N_3659,N_3996);
or U4324 (N_4324,N_3913,N_3716);
nor U4325 (N_4325,N_3661,N_3917);
or U4326 (N_4326,N_3646,N_3820);
nor U4327 (N_4327,N_3855,N_3821);
nand U4328 (N_4328,N_3552,N_3589);
nand U4329 (N_4329,N_3649,N_3510);
and U4330 (N_4330,N_3710,N_3619);
nand U4331 (N_4331,N_3774,N_3698);
or U4332 (N_4332,N_3542,N_3984);
xnor U4333 (N_4333,N_3870,N_3894);
xor U4334 (N_4334,N_3880,N_3603);
nor U4335 (N_4335,N_3586,N_3709);
nor U4336 (N_4336,N_3852,N_3996);
nand U4337 (N_4337,N_3995,N_3673);
nor U4338 (N_4338,N_3537,N_3651);
nand U4339 (N_4339,N_3610,N_3564);
or U4340 (N_4340,N_3784,N_3767);
and U4341 (N_4341,N_3936,N_3843);
and U4342 (N_4342,N_3679,N_3667);
nand U4343 (N_4343,N_3860,N_3854);
or U4344 (N_4344,N_3694,N_3813);
or U4345 (N_4345,N_3853,N_3861);
nand U4346 (N_4346,N_3507,N_3696);
nor U4347 (N_4347,N_3874,N_3583);
and U4348 (N_4348,N_3827,N_3960);
and U4349 (N_4349,N_3679,N_3572);
xor U4350 (N_4350,N_3831,N_3805);
nor U4351 (N_4351,N_3833,N_3802);
nand U4352 (N_4352,N_3987,N_3800);
nor U4353 (N_4353,N_3551,N_3924);
xor U4354 (N_4354,N_3867,N_3760);
and U4355 (N_4355,N_3526,N_3753);
nand U4356 (N_4356,N_3653,N_3897);
nand U4357 (N_4357,N_3598,N_3626);
and U4358 (N_4358,N_3913,N_3692);
nand U4359 (N_4359,N_3902,N_3971);
nor U4360 (N_4360,N_3589,N_3997);
xnor U4361 (N_4361,N_3636,N_3564);
nor U4362 (N_4362,N_3737,N_3631);
or U4363 (N_4363,N_3843,N_3686);
nor U4364 (N_4364,N_3977,N_3697);
nor U4365 (N_4365,N_3792,N_3835);
or U4366 (N_4366,N_3798,N_3706);
nand U4367 (N_4367,N_3871,N_3804);
xor U4368 (N_4368,N_3876,N_3655);
nand U4369 (N_4369,N_3573,N_3506);
nor U4370 (N_4370,N_3569,N_3587);
nor U4371 (N_4371,N_3617,N_3710);
xor U4372 (N_4372,N_3515,N_3851);
or U4373 (N_4373,N_3831,N_3847);
nand U4374 (N_4374,N_3863,N_3975);
xnor U4375 (N_4375,N_3669,N_3829);
and U4376 (N_4376,N_3699,N_3643);
xor U4377 (N_4377,N_3597,N_3515);
or U4378 (N_4378,N_3509,N_3770);
or U4379 (N_4379,N_3542,N_3726);
nand U4380 (N_4380,N_3786,N_3939);
nand U4381 (N_4381,N_3724,N_3747);
nor U4382 (N_4382,N_3942,N_3881);
nand U4383 (N_4383,N_3712,N_3500);
nand U4384 (N_4384,N_3994,N_3937);
and U4385 (N_4385,N_3602,N_3506);
and U4386 (N_4386,N_3628,N_3998);
nand U4387 (N_4387,N_3691,N_3760);
nor U4388 (N_4388,N_3665,N_3831);
nand U4389 (N_4389,N_3654,N_3591);
nand U4390 (N_4390,N_3559,N_3772);
and U4391 (N_4391,N_3540,N_3792);
and U4392 (N_4392,N_3505,N_3847);
or U4393 (N_4393,N_3881,N_3822);
xnor U4394 (N_4394,N_3961,N_3749);
and U4395 (N_4395,N_3554,N_3598);
nand U4396 (N_4396,N_3656,N_3605);
or U4397 (N_4397,N_3536,N_3756);
and U4398 (N_4398,N_3952,N_3619);
nand U4399 (N_4399,N_3626,N_3530);
nor U4400 (N_4400,N_3597,N_3553);
nor U4401 (N_4401,N_3841,N_3501);
nand U4402 (N_4402,N_3595,N_3954);
and U4403 (N_4403,N_3960,N_3681);
and U4404 (N_4404,N_3660,N_3640);
or U4405 (N_4405,N_3564,N_3932);
xor U4406 (N_4406,N_3701,N_3602);
nor U4407 (N_4407,N_3615,N_3996);
and U4408 (N_4408,N_3506,N_3699);
nor U4409 (N_4409,N_3891,N_3708);
and U4410 (N_4410,N_3870,N_3665);
xnor U4411 (N_4411,N_3714,N_3919);
and U4412 (N_4412,N_3921,N_3901);
xnor U4413 (N_4413,N_3754,N_3827);
and U4414 (N_4414,N_3573,N_3788);
and U4415 (N_4415,N_3875,N_3682);
and U4416 (N_4416,N_3960,N_3856);
xnor U4417 (N_4417,N_3946,N_3502);
nor U4418 (N_4418,N_3757,N_3708);
and U4419 (N_4419,N_3836,N_3757);
or U4420 (N_4420,N_3697,N_3547);
and U4421 (N_4421,N_3743,N_3850);
or U4422 (N_4422,N_3874,N_3906);
and U4423 (N_4423,N_3986,N_3512);
or U4424 (N_4424,N_3829,N_3551);
or U4425 (N_4425,N_3531,N_3885);
or U4426 (N_4426,N_3893,N_3918);
nor U4427 (N_4427,N_3682,N_3560);
nand U4428 (N_4428,N_3578,N_3623);
or U4429 (N_4429,N_3934,N_3764);
nor U4430 (N_4430,N_3613,N_3783);
xor U4431 (N_4431,N_3556,N_3983);
or U4432 (N_4432,N_3876,N_3961);
and U4433 (N_4433,N_3545,N_3968);
nor U4434 (N_4434,N_3842,N_3682);
and U4435 (N_4435,N_3728,N_3666);
nand U4436 (N_4436,N_3702,N_3723);
and U4437 (N_4437,N_3986,N_3698);
or U4438 (N_4438,N_3805,N_3859);
xnor U4439 (N_4439,N_3735,N_3925);
nor U4440 (N_4440,N_3838,N_3949);
xnor U4441 (N_4441,N_3678,N_3832);
and U4442 (N_4442,N_3900,N_3714);
nor U4443 (N_4443,N_3519,N_3901);
xnor U4444 (N_4444,N_3807,N_3868);
nor U4445 (N_4445,N_3656,N_3901);
xor U4446 (N_4446,N_3701,N_3787);
nand U4447 (N_4447,N_3907,N_3977);
nor U4448 (N_4448,N_3633,N_3973);
or U4449 (N_4449,N_3633,N_3518);
xor U4450 (N_4450,N_3577,N_3554);
and U4451 (N_4451,N_3993,N_3812);
or U4452 (N_4452,N_3790,N_3925);
or U4453 (N_4453,N_3624,N_3818);
or U4454 (N_4454,N_3980,N_3863);
nor U4455 (N_4455,N_3694,N_3916);
nor U4456 (N_4456,N_3627,N_3673);
and U4457 (N_4457,N_3817,N_3543);
nor U4458 (N_4458,N_3880,N_3738);
or U4459 (N_4459,N_3629,N_3872);
and U4460 (N_4460,N_3811,N_3955);
or U4461 (N_4461,N_3529,N_3573);
nand U4462 (N_4462,N_3582,N_3854);
and U4463 (N_4463,N_3840,N_3884);
nand U4464 (N_4464,N_3571,N_3700);
nand U4465 (N_4465,N_3824,N_3670);
or U4466 (N_4466,N_3953,N_3599);
or U4467 (N_4467,N_3733,N_3983);
nand U4468 (N_4468,N_3865,N_3526);
or U4469 (N_4469,N_3581,N_3855);
and U4470 (N_4470,N_3563,N_3926);
nand U4471 (N_4471,N_3755,N_3588);
xor U4472 (N_4472,N_3738,N_3741);
xnor U4473 (N_4473,N_3724,N_3702);
nand U4474 (N_4474,N_3844,N_3591);
xnor U4475 (N_4475,N_3930,N_3834);
nand U4476 (N_4476,N_3842,N_3758);
or U4477 (N_4477,N_3923,N_3558);
nor U4478 (N_4478,N_3687,N_3856);
or U4479 (N_4479,N_3506,N_3897);
and U4480 (N_4480,N_3770,N_3549);
xor U4481 (N_4481,N_3980,N_3501);
nor U4482 (N_4482,N_3864,N_3571);
or U4483 (N_4483,N_3956,N_3632);
nand U4484 (N_4484,N_3548,N_3965);
and U4485 (N_4485,N_3794,N_3549);
nor U4486 (N_4486,N_3584,N_3848);
xnor U4487 (N_4487,N_3786,N_3571);
or U4488 (N_4488,N_3766,N_3883);
or U4489 (N_4489,N_3764,N_3978);
or U4490 (N_4490,N_3675,N_3960);
xor U4491 (N_4491,N_3765,N_3694);
or U4492 (N_4492,N_3611,N_3999);
or U4493 (N_4493,N_3767,N_3595);
xor U4494 (N_4494,N_3787,N_3801);
xnor U4495 (N_4495,N_3521,N_3578);
and U4496 (N_4496,N_3537,N_3881);
nor U4497 (N_4497,N_3889,N_3752);
nand U4498 (N_4498,N_3946,N_3558);
nor U4499 (N_4499,N_3560,N_3730);
and U4500 (N_4500,N_4376,N_4474);
nand U4501 (N_4501,N_4081,N_4115);
nand U4502 (N_4502,N_4235,N_4187);
or U4503 (N_4503,N_4327,N_4247);
nand U4504 (N_4504,N_4328,N_4244);
or U4505 (N_4505,N_4489,N_4453);
and U4506 (N_4506,N_4041,N_4363);
and U4507 (N_4507,N_4050,N_4248);
and U4508 (N_4508,N_4373,N_4031);
nor U4509 (N_4509,N_4083,N_4001);
xnor U4510 (N_4510,N_4285,N_4215);
nor U4511 (N_4511,N_4319,N_4243);
nand U4512 (N_4512,N_4411,N_4483);
and U4513 (N_4513,N_4256,N_4185);
xor U4514 (N_4514,N_4389,N_4498);
xnor U4515 (N_4515,N_4109,N_4023);
or U4516 (N_4516,N_4129,N_4125);
nand U4517 (N_4517,N_4232,N_4422);
xor U4518 (N_4518,N_4291,N_4469);
nand U4519 (N_4519,N_4142,N_4384);
or U4520 (N_4520,N_4266,N_4211);
nand U4521 (N_4521,N_4107,N_4466);
and U4522 (N_4522,N_4245,N_4095);
nand U4523 (N_4523,N_4153,N_4370);
nand U4524 (N_4524,N_4262,N_4352);
and U4525 (N_4525,N_4089,N_4061);
xnor U4526 (N_4526,N_4416,N_4191);
xor U4527 (N_4527,N_4015,N_4400);
nor U4528 (N_4528,N_4003,N_4482);
xor U4529 (N_4529,N_4124,N_4274);
or U4530 (N_4530,N_4077,N_4417);
nand U4531 (N_4531,N_4216,N_4258);
and U4532 (N_4532,N_4340,N_4280);
xnor U4533 (N_4533,N_4074,N_4423);
xnor U4534 (N_4534,N_4009,N_4217);
xnor U4535 (N_4535,N_4073,N_4487);
and U4536 (N_4536,N_4457,N_4080);
nor U4537 (N_4537,N_4158,N_4257);
nor U4538 (N_4538,N_4007,N_4242);
and U4539 (N_4539,N_4306,N_4252);
and U4540 (N_4540,N_4298,N_4198);
and U4541 (N_4541,N_4193,N_4227);
nor U4542 (N_4542,N_4047,N_4288);
and U4543 (N_4543,N_4320,N_4163);
nand U4544 (N_4544,N_4428,N_4143);
or U4545 (N_4545,N_4412,N_4338);
and U4546 (N_4546,N_4255,N_4325);
nor U4547 (N_4547,N_4046,N_4164);
and U4548 (N_4548,N_4394,N_4408);
and U4549 (N_4549,N_4410,N_4100);
nand U4550 (N_4550,N_4155,N_4108);
or U4551 (N_4551,N_4149,N_4273);
nor U4552 (N_4552,N_4289,N_4383);
nand U4553 (N_4553,N_4287,N_4345);
xnor U4554 (N_4554,N_4126,N_4159);
nor U4555 (N_4555,N_4194,N_4203);
and U4556 (N_4556,N_4082,N_4398);
nor U4557 (N_4557,N_4069,N_4278);
nor U4558 (N_4558,N_4393,N_4018);
and U4559 (N_4559,N_4399,N_4059);
xnor U4560 (N_4560,N_4035,N_4296);
nor U4561 (N_4561,N_4360,N_4213);
nand U4562 (N_4562,N_4418,N_4254);
xnor U4563 (N_4563,N_4459,N_4406);
nor U4564 (N_4564,N_4478,N_4425);
xor U4565 (N_4565,N_4025,N_4043);
nor U4566 (N_4566,N_4378,N_4166);
nand U4567 (N_4567,N_4094,N_4314);
nor U4568 (N_4568,N_4356,N_4337);
xnor U4569 (N_4569,N_4004,N_4456);
xor U4570 (N_4570,N_4065,N_4174);
or U4571 (N_4571,N_4008,N_4091);
nand U4572 (N_4572,N_4171,N_4202);
nand U4573 (N_4573,N_4496,N_4409);
xor U4574 (N_4574,N_4177,N_4060);
nand U4575 (N_4575,N_4448,N_4246);
and U4576 (N_4576,N_4147,N_4068);
nand U4577 (N_4577,N_4434,N_4075);
nor U4578 (N_4578,N_4057,N_4197);
xor U4579 (N_4579,N_4313,N_4051);
xor U4580 (N_4580,N_4486,N_4386);
xor U4581 (N_4581,N_4052,N_4032);
xnor U4582 (N_4582,N_4214,N_4120);
xor U4583 (N_4583,N_4477,N_4200);
xnor U4584 (N_4584,N_4316,N_4268);
xor U4585 (N_4585,N_4377,N_4136);
xor U4586 (N_4586,N_4240,N_4414);
nor U4587 (N_4587,N_4455,N_4461);
nor U4588 (N_4588,N_4016,N_4460);
nor U4589 (N_4589,N_4267,N_4019);
xnor U4590 (N_4590,N_4467,N_4303);
nor U4591 (N_4591,N_4013,N_4105);
nand U4592 (N_4592,N_4076,N_4321);
xnor U4593 (N_4593,N_4465,N_4072);
nor U4594 (N_4594,N_4139,N_4223);
nand U4595 (N_4595,N_4006,N_4301);
xor U4596 (N_4596,N_4330,N_4495);
and U4597 (N_4597,N_4450,N_4055);
or U4598 (N_4598,N_4437,N_4140);
nand U4599 (N_4599,N_4010,N_4344);
nor U4600 (N_4600,N_4388,N_4172);
xor U4601 (N_4601,N_4146,N_4118);
nor U4602 (N_4602,N_4182,N_4403);
nand U4603 (N_4603,N_4259,N_4021);
or U4604 (N_4604,N_4475,N_4430);
nor U4605 (N_4605,N_4445,N_4440);
nor U4606 (N_4606,N_4219,N_4310);
and U4607 (N_4607,N_4331,N_4294);
nand U4608 (N_4608,N_4335,N_4098);
and U4609 (N_4609,N_4367,N_4020);
nand U4610 (N_4610,N_4375,N_4110);
nand U4611 (N_4611,N_4066,N_4229);
or U4612 (N_4612,N_4379,N_4368);
or U4613 (N_4613,N_4421,N_4299);
and U4614 (N_4614,N_4293,N_4261);
xnor U4615 (N_4615,N_4387,N_4024);
or U4616 (N_4616,N_4134,N_4183);
or U4617 (N_4617,N_4225,N_4271);
nand U4618 (N_4618,N_4151,N_4341);
or U4619 (N_4619,N_4405,N_4099);
and U4620 (N_4620,N_4300,N_4042);
and U4621 (N_4621,N_4471,N_4002);
nor U4622 (N_4622,N_4226,N_4438);
or U4623 (N_4623,N_4462,N_4053);
or U4624 (N_4624,N_4154,N_4106);
nor U4625 (N_4625,N_4000,N_4432);
and U4626 (N_4626,N_4112,N_4355);
nor U4627 (N_4627,N_4396,N_4169);
nand U4628 (N_4628,N_4179,N_4429);
xor U4629 (N_4629,N_4084,N_4307);
xnor U4630 (N_4630,N_4103,N_4427);
or U4631 (N_4631,N_4479,N_4208);
or U4632 (N_4632,N_4260,N_4284);
nor U4633 (N_4633,N_4443,N_4322);
or U4634 (N_4634,N_4184,N_4323);
and U4635 (N_4635,N_4404,N_4264);
and U4636 (N_4636,N_4144,N_4366);
or U4637 (N_4637,N_4026,N_4263);
nor U4638 (N_4638,N_4326,N_4119);
nand U4639 (N_4639,N_4117,N_4339);
or U4640 (N_4640,N_4464,N_4236);
nand U4641 (N_4641,N_4485,N_4090);
xor U4642 (N_4642,N_4148,N_4251);
and U4643 (N_4643,N_4454,N_4114);
and U4644 (N_4644,N_4441,N_4491);
nor U4645 (N_4645,N_4141,N_4093);
xnor U4646 (N_4646,N_4336,N_4249);
or U4647 (N_4647,N_4292,N_4311);
nor U4648 (N_4648,N_4038,N_4239);
and U4649 (N_4649,N_4354,N_4175);
and U4650 (N_4650,N_4269,N_4221);
xnor U4651 (N_4651,N_4064,N_4342);
and U4652 (N_4652,N_4401,N_4150);
and U4653 (N_4653,N_4241,N_4230);
xnor U4654 (N_4654,N_4343,N_4395);
nor U4655 (N_4655,N_4017,N_4011);
nor U4656 (N_4656,N_4022,N_4458);
nor U4657 (N_4657,N_4044,N_4176);
or U4658 (N_4658,N_4131,N_4380);
nand U4659 (N_4659,N_4062,N_4056);
or U4660 (N_4660,N_4447,N_4442);
nand U4661 (N_4661,N_4279,N_4283);
or U4662 (N_4662,N_4167,N_4204);
xnor U4663 (N_4663,N_4130,N_4029);
and U4664 (N_4664,N_4392,N_4036);
and U4665 (N_4665,N_4092,N_4282);
nor U4666 (N_4666,N_4222,N_4156);
or U4667 (N_4667,N_4196,N_4049);
xnor U4668 (N_4668,N_4201,N_4087);
nor U4669 (N_4669,N_4497,N_4250);
and U4670 (N_4670,N_4220,N_4039);
nor U4671 (N_4671,N_4365,N_4138);
and U4672 (N_4672,N_4488,N_4111);
nand U4673 (N_4673,N_4173,N_4494);
xor U4674 (N_4674,N_4332,N_4116);
nand U4675 (N_4675,N_4123,N_4424);
nor U4676 (N_4676,N_4195,N_4309);
nor U4677 (N_4677,N_4439,N_4228);
and U4678 (N_4678,N_4357,N_4463);
nand U4679 (N_4679,N_4484,N_4348);
or U4680 (N_4680,N_4048,N_4063);
nor U4681 (N_4681,N_4317,N_4234);
nand U4682 (N_4682,N_4426,N_4451);
nor U4683 (N_4683,N_4157,N_4444);
nor U4684 (N_4684,N_4290,N_4132);
and U4685 (N_4685,N_4402,N_4351);
xnor U4686 (N_4686,N_4034,N_4499);
xnor U4687 (N_4687,N_4372,N_4128);
and U4688 (N_4688,N_4127,N_4190);
nand U4689 (N_4689,N_4295,N_4079);
nand U4690 (N_4690,N_4033,N_4481);
or U4691 (N_4691,N_4407,N_4028);
xor U4692 (N_4692,N_4086,N_4361);
and U4693 (N_4693,N_4037,N_4358);
and U4694 (N_4694,N_4413,N_4420);
and U4695 (N_4695,N_4318,N_4433);
nor U4696 (N_4696,N_4473,N_4302);
and U4697 (N_4697,N_4178,N_4085);
nand U4698 (N_4698,N_4180,N_4027);
nand U4699 (N_4699,N_4212,N_4277);
and U4700 (N_4700,N_4121,N_4209);
or U4701 (N_4701,N_4371,N_4161);
or U4702 (N_4702,N_4346,N_4308);
nor U4703 (N_4703,N_4286,N_4054);
xnor U4704 (N_4704,N_4030,N_4186);
or U4705 (N_4705,N_4189,N_4382);
and U4706 (N_4706,N_4122,N_4233);
nand U4707 (N_4707,N_4133,N_4436);
and U4708 (N_4708,N_4012,N_4058);
and U4709 (N_4709,N_4472,N_4005);
and U4710 (N_4710,N_4096,N_4101);
nor U4711 (N_4711,N_4192,N_4419);
or U4712 (N_4712,N_4067,N_4170);
and U4713 (N_4713,N_4270,N_4364);
xnor U4714 (N_4714,N_4493,N_4480);
nand U4715 (N_4715,N_4353,N_4381);
nand U4716 (N_4716,N_4490,N_4468);
nand U4717 (N_4717,N_4359,N_4231);
nor U4718 (N_4718,N_4446,N_4304);
xnor U4719 (N_4719,N_4207,N_4102);
nand U4720 (N_4720,N_4181,N_4078);
nand U4721 (N_4721,N_4071,N_4168);
and U4722 (N_4722,N_4415,N_4275);
nand U4723 (N_4723,N_4206,N_4334);
nor U4724 (N_4724,N_4014,N_4135);
or U4725 (N_4725,N_4391,N_4276);
nor U4726 (N_4726,N_4435,N_4113);
and U4727 (N_4727,N_4362,N_4088);
or U4728 (N_4728,N_4165,N_4224);
nor U4729 (N_4729,N_4397,N_4152);
or U4730 (N_4730,N_4238,N_4272);
nor U4731 (N_4731,N_4324,N_4218);
and U4732 (N_4732,N_4385,N_4431);
or U4733 (N_4733,N_4374,N_4329);
and U4734 (N_4734,N_4470,N_4369);
nor U4735 (N_4735,N_4162,N_4188);
nor U4736 (N_4736,N_4312,N_4265);
xor U4737 (N_4737,N_4070,N_4160);
or U4738 (N_4738,N_4315,N_4476);
nand U4739 (N_4739,N_4137,N_4333);
nand U4740 (N_4740,N_4297,N_4390);
xor U4741 (N_4741,N_4045,N_4040);
xor U4742 (N_4742,N_4104,N_4199);
xnor U4743 (N_4743,N_4237,N_4253);
nand U4744 (N_4744,N_4347,N_4097);
nor U4745 (N_4745,N_4210,N_4205);
or U4746 (N_4746,N_4350,N_4305);
or U4747 (N_4747,N_4145,N_4449);
nor U4748 (N_4748,N_4281,N_4492);
xnor U4749 (N_4749,N_4349,N_4452);
nand U4750 (N_4750,N_4473,N_4058);
nor U4751 (N_4751,N_4035,N_4281);
xor U4752 (N_4752,N_4427,N_4335);
nand U4753 (N_4753,N_4197,N_4300);
xnor U4754 (N_4754,N_4487,N_4083);
xnor U4755 (N_4755,N_4317,N_4144);
nand U4756 (N_4756,N_4179,N_4488);
and U4757 (N_4757,N_4318,N_4159);
xor U4758 (N_4758,N_4350,N_4307);
and U4759 (N_4759,N_4192,N_4294);
and U4760 (N_4760,N_4345,N_4356);
xnor U4761 (N_4761,N_4095,N_4108);
nand U4762 (N_4762,N_4399,N_4276);
nor U4763 (N_4763,N_4032,N_4236);
nor U4764 (N_4764,N_4417,N_4301);
xor U4765 (N_4765,N_4406,N_4052);
xor U4766 (N_4766,N_4421,N_4126);
xnor U4767 (N_4767,N_4439,N_4338);
xor U4768 (N_4768,N_4433,N_4167);
or U4769 (N_4769,N_4174,N_4155);
nand U4770 (N_4770,N_4211,N_4344);
xnor U4771 (N_4771,N_4210,N_4113);
xor U4772 (N_4772,N_4134,N_4434);
xnor U4773 (N_4773,N_4271,N_4142);
xnor U4774 (N_4774,N_4111,N_4073);
nor U4775 (N_4775,N_4141,N_4492);
or U4776 (N_4776,N_4099,N_4281);
nand U4777 (N_4777,N_4164,N_4219);
or U4778 (N_4778,N_4122,N_4212);
and U4779 (N_4779,N_4226,N_4255);
xnor U4780 (N_4780,N_4115,N_4317);
and U4781 (N_4781,N_4209,N_4094);
and U4782 (N_4782,N_4370,N_4110);
nand U4783 (N_4783,N_4031,N_4114);
nor U4784 (N_4784,N_4317,N_4435);
xor U4785 (N_4785,N_4074,N_4273);
nor U4786 (N_4786,N_4294,N_4468);
nand U4787 (N_4787,N_4317,N_4289);
or U4788 (N_4788,N_4201,N_4223);
nand U4789 (N_4789,N_4443,N_4145);
or U4790 (N_4790,N_4472,N_4374);
and U4791 (N_4791,N_4147,N_4032);
or U4792 (N_4792,N_4088,N_4170);
or U4793 (N_4793,N_4032,N_4100);
and U4794 (N_4794,N_4054,N_4441);
nand U4795 (N_4795,N_4134,N_4357);
nor U4796 (N_4796,N_4336,N_4024);
and U4797 (N_4797,N_4262,N_4372);
xor U4798 (N_4798,N_4009,N_4392);
or U4799 (N_4799,N_4209,N_4383);
or U4800 (N_4800,N_4047,N_4120);
or U4801 (N_4801,N_4216,N_4062);
and U4802 (N_4802,N_4133,N_4109);
and U4803 (N_4803,N_4189,N_4038);
or U4804 (N_4804,N_4367,N_4098);
nor U4805 (N_4805,N_4049,N_4218);
or U4806 (N_4806,N_4046,N_4330);
xor U4807 (N_4807,N_4254,N_4247);
nand U4808 (N_4808,N_4018,N_4252);
or U4809 (N_4809,N_4489,N_4297);
nand U4810 (N_4810,N_4064,N_4387);
nand U4811 (N_4811,N_4156,N_4240);
nand U4812 (N_4812,N_4309,N_4172);
xor U4813 (N_4813,N_4370,N_4022);
or U4814 (N_4814,N_4313,N_4496);
or U4815 (N_4815,N_4257,N_4317);
nand U4816 (N_4816,N_4138,N_4250);
nand U4817 (N_4817,N_4475,N_4030);
and U4818 (N_4818,N_4220,N_4056);
or U4819 (N_4819,N_4443,N_4302);
nor U4820 (N_4820,N_4266,N_4116);
or U4821 (N_4821,N_4488,N_4362);
and U4822 (N_4822,N_4061,N_4399);
and U4823 (N_4823,N_4343,N_4362);
xnor U4824 (N_4824,N_4252,N_4237);
nand U4825 (N_4825,N_4498,N_4473);
and U4826 (N_4826,N_4274,N_4141);
xor U4827 (N_4827,N_4032,N_4215);
or U4828 (N_4828,N_4324,N_4358);
nand U4829 (N_4829,N_4066,N_4308);
nand U4830 (N_4830,N_4385,N_4082);
and U4831 (N_4831,N_4062,N_4428);
or U4832 (N_4832,N_4473,N_4011);
nor U4833 (N_4833,N_4104,N_4012);
xnor U4834 (N_4834,N_4336,N_4232);
xor U4835 (N_4835,N_4355,N_4330);
and U4836 (N_4836,N_4164,N_4021);
and U4837 (N_4837,N_4157,N_4385);
nand U4838 (N_4838,N_4267,N_4472);
xnor U4839 (N_4839,N_4372,N_4145);
nor U4840 (N_4840,N_4054,N_4035);
nand U4841 (N_4841,N_4276,N_4179);
nand U4842 (N_4842,N_4148,N_4054);
xor U4843 (N_4843,N_4181,N_4161);
nand U4844 (N_4844,N_4268,N_4136);
nor U4845 (N_4845,N_4016,N_4336);
nand U4846 (N_4846,N_4327,N_4178);
nand U4847 (N_4847,N_4387,N_4043);
and U4848 (N_4848,N_4462,N_4488);
or U4849 (N_4849,N_4385,N_4270);
nand U4850 (N_4850,N_4429,N_4376);
nand U4851 (N_4851,N_4280,N_4108);
nand U4852 (N_4852,N_4471,N_4242);
and U4853 (N_4853,N_4052,N_4453);
or U4854 (N_4854,N_4189,N_4424);
xnor U4855 (N_4855,N_4426,N_4372);
nand U4856 (N_4856,N_4271,N_4379);
and U4857 (N_4857,N_4078,N_4192);
nor U4858 (N_4858,N_4304,N_4419);
nor U4859 (N_4859,N_4362,N_4158);
or U4860 (N_4860,N_4452,N_4331);
nand U4861 (N_4861,N_4009,N_4154);
and U4862 (N_4862,N_4337,N_4322);
and U4863 (N_4863,N_4161,N_4122);
nor U4864 (N_4864,N_4305,N_4459);
nor U4865 (N_4865,N_4480,N_4038);
nor U4866 (N_4866,N_4186,N_4281);
xor U4867 (N_4867,N_4217,N_4260);
or U4868 (N_4868,N_4227,N_4158);
or U4869 (N_4869,N_4357,N_4426);
or U4870 (N_4870,N_4213,N_4145);
nand U4871 (N_4871,N_4224,N_4484);
and U4872 (N_4872,N_4313,N_4003);
nand U4873 (N_4873,N_4396,N_4301);
or U4874 (N_4874,N_4091,N_4122);
nor U4875 (N_4875,N_4253,N_4409);
nor U4876 (N_4876,N_4298,N_4244);
xnor U4877 (N_4877,N_4239,N_4048);
nand U4878 (N_4878,N_4442,N_4198);
nand U4879 (N_4879,N_4198,N_4114);
nor U4880 (N_4880,N_4245,N_4076);
or U4881 (N_4881,N_4367,N_4257);
and U4882 (N_4882,N_4066,N_4248);
nor U4883 (N_4883,N_4348,N_4227);
and U4884 (N_4884,N_4457,N_4133);
and U4885 (N_4885,N_4493,N_4454);
and U4886 (N_4886,N_4195,N_4409);
nor U4887 (N_4887,N_4070,N_4439);
and U4888 (N_4888,N_4133,N_4235);
nor U4889 (N_4889,N_4370,N_4302);
or U4890 (N_4890,N_4425,N_4358);
nand U4891 (N_4891,N_4452,N_4461);
nor U4892 (N_4892,N_4218,N_4400);
and U4893 (N_4893,N_4384,N_4175);
and U4894 (N_4894,N_4019,N_4304);
or U4895 (N_4895,N_4249,N_4152);
and U4896 (N_4896,N_4020,N_4265);
and U4897 (N_4897,N_4028,N_4467);
nand U4898 (N_4898,N_4094,N_4333);
xnor U4899 (N_4899,N_4290,N_4025);
nor U4900 (N_4900,N_4138,N_4222);
xnor U4901 (N_4901,N_4071,N_4163);
xnor U4902 (N_4902,N_4475,N_4225);
and U4903 (N_4903,N_4465,N_4372);
and U4904 (N_4904,N_4495,N_4175);
and U4905 (N_4905,N_4094,N_4250);
or U4906 (N_4906,N_4482,N_4144);
nand U4907 (N_4907,N_4373,N_4403);
or U4908 (N_4908,N_4264,N_4290);
or U4909 (N_4909,N_4275,N_4002);
nor U4910 (N_4910,N_4319,N_4066);
nor U4911 (N_4911,N_4347,N_4165);
nor U4912 (N_4912,N_4149,N_4021);
or U4913 (N_4913,N_4338,N_4362);
nor U4914 (N_4914,N_4031,N_4480);
nor U4915 (N_4915,N_4154,N_4012);
xnor U4916 (N_4916,N_4054,N_4195);
and U4917 (N_4917,N_4271,N_4085);
nor U4918 (N_4918,N_4459,N_4175);
nor U4919 (N_4919,N_4013,N_4384);
nor U4920 (N_4920,N_4476,N_4355);
or U4921 (N_4921,N_4446,N_4089);
xor U4922 (N_4922,N_4149,N_4454);
nand U4923 (N_4923,N_4444,N_4085);
nand U4924 (N_4924,N_4049,N_4475);
and U4925 (N_4925,N_4380,N_4341);
nand U4926 (N_4926,N_4368,N_4106);
nor U4927 (N_4927,N_4410,N_4341);
or U4928 (N_4928,N_4210,N_4475);
xnor U4929 (N_4929,N_4285,N_4477);
xnor U4930 (N_4930,N_4370,N_4242);
and U4931 (N_4931,N_4200,N_4239);
and U4932 (N_4932,N_4116,N_4063);
xor U4933 (N_4933,N_4052,N_4320);
nor U4934 (N_4934,N_4251,N_4436);
nor U4935 (N_4935,N_4150,N_4004);
nor U4936 (N_4936,N_4372,N_4412);
and U4937 (N_4937,N_4327,N_4146);
xor U4938 (N_4938,N_4473,N_4447);
and U4939 (N_4939,N_4453,N_4493);
nand U4940 (N_4940,N_4050,N_4465);
and U4941 (N_4941,N_4208,N_4195);
nand U4942 (N_4942,N_4367,N_4049);
nor U4943 (N_4943,N_4202,N_4448);
nand U4944 (N_4944,N_4451,N_4312);
or U4945 (N_4945,N_4035,N_4328);
or U4946 (N_4946,N_4408,N_4028);
nor U4947 (N_4947,N_4238,N_4139);
nor U4948 (N_4948,N_4441,N_4094);
nor U4949 (N_4949,N_4181,N_4267);
and U4950 (N_4950,N_4078,N_4234);
nand U4951 (N_4951,N_4200,N_4245);
xnor U4952 (N_4952,N_4485,N_4149);
xnor U4953 (N_4953,N_4286,N_4053);
xor U4954 (N_4954,N_4017,N_4471);
nor U4955 (N_4955,N_4189,N_4270);
xor U4956 (N_4956,N_4440,N_4136);
xnor U4957 (N_4957,N_4206,N_4186);
and U4958 (N_4958,N_4459,N_4280);
xnor U4959 (N_4959,N_4004,N_4155);
and U4960 (N_4960,N_4379,N_4043);
or U4961 (N_4961,N_4469,N_4142);
and U4962 (N_4962,N_4245,N_4106);
and U4963 (N_4963,N_4349,N_4085);
xnor U4964 (N_4964,N_4201,N_4434);
nor U4965 (N_4965,N_4035,N_4242);
or U4966 (N_4966,N_4138,N_4363);
xnor U4967 (N_4967,N_4336,N_4372);
and U4968 (N_4968,N_4257,N_4384);
and U4969 (N_4969,N_4342,N_4328);
or U4970 (N_4970,N_4338,N_4228);
or U4971 (N_4971,N_4460,N_4168);
and U4972 (N_4972,N_4330,N_4202);
xor U4973 (N_4973,N_4038,N_4455);
and U4974 (N_4974,N_4014,N_4018);
or U4975 (N_4975,N_4312,N_4380);
and U4976 (N_4976,N_4000,N_4325);
and U4977 (N_4977,N_4070,N_4434);
or U4978 (N_4978,N_4429,N_4366);
nand U4979 (N_4979,N_4318,N_4359);
nand U4980 (N_4980,N_4182,N_4406);
xnor U4981 (N_4981,N_4107,N_4364);
and U4982 (N_4982,N_4052,N_4351);
xor U4983 (N_4983,N_4228,N_4089);
or U4984 (N_4984,N_4309,N_4438);
and U4985 (N_4985,N_4115,N_4092);
xor U4986 (N_4986,N_4374,N_4088);
nor U4987 (N_4987,N_4160,N_4230);
or U4988 (N_4988,N_4449,N_4179);
and U4989 (N_4989,N_4212,N_4369);
xor U4990 (N_4990,N_4486,N_4320);
nor U4991 (N_4991,N_4096,N_4209);
or U4992 (N_4992,N_4349,N_4309);
nand U4993 (N_4993,N_4345,N_4009);
nand U4994 (N_4994,N_4297,N_4290);
xor U4995 (N_4995,N_4119,N_4374);
nand U4996 (N_4996,N_4318,N_4345);
xor U4997 (N_4997,N_4038,N_4240);
xnor U4998 (N_4998,N_4338,N_4194);
nand U4999 (N_4999,N_4225,N_4260);
nand U5000 (N_5000,N_4732,N_4939);
and U5001 (N_5001,N_4552,N_4865);
xnor U5002 (N_5002,N_4974,N_4760);
nand U5003 (N_5003,N_4557,N_4862);
nand U5004 (N_5004,N_4843,N_4813);
and U5005 (N_5005,N_4507,N_4540);
nor U5006 (N_5006,N_4863,N_4743);
and U5007 (N_5007,N_4703,N_4527);
and U5008 (N_5008,N_4963,N_4751);
and U5009 (N_5009,N_4806,N_4500);
or U5010 (N_5010,N_4822,N_4689);
or U5011 (N_5011,N_4807,N_4940);
nand U5012 (N_5012,N_4979,N_4699);
nor U5013 (N_5013,N_4891,N_4784);
or U5014 (N_5014,N_4578,N_4906);
and U5015 (N_5015,N_4568,N_4551);
xor U5016 (N_5016,N_4716,N_4966);
nor U5017 (N_5017,N_4772,N_4810);
nor U5018 (N_5018,N_4782,N_4528);
and U5019 (N_5019,N_4977,N_4763);
xor U5020 (N_5020,N_4580,N_4781);
xnor U5021 (N_5021,N_4741,N_4773);
nor U5022 (N_5022,N_4915,N_4944);
or U5023 (N_5023,N_4725,N_4561);
nand U5024 (N_5024,N_4892,N_4925);
xor U5025 (N_5025,N_4942,N_4984);
xnor U5026 (N_5026,N_4590,N_4541);
or U5027 (N_5027,N_4790,N_4860);
and U5028 (N_5028,N_4964,N_4625);
and U5029 (N_5029,N_4611,N_4785);
nand U5030 (N_5030,N_4727,N_4951);
nor U5031 (N_5031,N_4645,N_4890);
nor U5032 (N_5032,N_4538,N_4635);
nand U5033 (N_5033,N_4833,N_4735);
or U5034 (N_5034,N_4912,N_4986);
and U5035 (N_5035,N_4570,N_4564);
xnor U5036 (N_5036,N_4934,N_4852);
or U5037 (N_5037,N_4879,N_4644);
or U5038 (N_5038,N_4989,N_4731);
nor U5039 (N_5039,N_4853,N_4764);
xnor U5040 (N_5040,N_4624,N_4658);
and U5041 (N_5041,N_4796,N_4519);
or U5042 (N_5042,N_4893,N_4820);
and U5043 (N_5043,N_4631,N_4740);
or U5044 (N_5044,N_4677,N_4622);
nor U5045 (N_5045,N_4596,N_4530);
and U5046 (N_5046,N_4664,N_4577);
nor U5047 (N_5047,N_4554,N_4821);
or U5048 (N_5048,N_4562,N_4539);
nor U5049 (N_5049,N_4777,N_4526);
xor U5050 (N_5050,N_4723,N_4774);
and U5051 (N_5051,N_4982,N_4592);
nor U5052 (N_5052,N_4895,N_4824);
nand U5053 (N_5053,N_4585,N_4768);
nand U5054 (N_5054,N_4762,N_4867);
nor U5055 (N_5055,N_4767,N_4579);
and U5056 (N_5056,N_4722,N_4812);
nand U5057 (N_5057,N_4649,N_4945);
nand U5058 (N_5058,N_4943,N_4537);
nor U5059 (N_5059,N_4651,N_4887);
xnor U5060 (N_5060,N_4896,N_4965);
nand U5061 (N_5061,N_4673,N_4968);
and U5062 (N_5062,N_4769,N_4818);
or U5063 (N_5063,N_4758,N_4718);
or U5064 (N_5064,N_4829,N_4755);
xnor U5065 (N_5065,N_4857,N_4707);
and U5066 (N_5066,N_4819,N_4676);
nor U5067 (N_5067,N_4987,N_4503);
and U5068 (N_5068,N_4599,N_4612);
nand U5069 (N_5069,N_4981,N_4757);
nand U5070 (N_5070,N_4908,N_4931);
nor U5071 (N_5071,N_4911,N_4717);
and U5072 (N_5072,N_4949,N_4960);
nor U5073 (N_5073,N_4910,N_4980);
and U5074 (N_5074,N_4501,N_4505);
nor U5075 (N_5075,N_4745,N_4898);
nand U5076 (N_5076,N_4927,N_4525);
or U5077 (N_5077,N_4854,N_4826);
nor U5078 (N_5078,N_4866,N_4650);
or U5079 (N_5079,N_4555,N_4929);
xor U5080 (N_5080,N_4692,N_4778);
nor U5081 (N_5081,N_4665,N_4815);
or U5082 (N_5082,N_4514,N_4654);
nor U5083 (N_5083,N_4957,N_4695);
or U5084 (N_5084,N_4997,N_4633);
xor U5085 (N_5085,N_4720,N_4930);
nor U5086 (N_5086,N_4524,N_4582);
and U5087 (N_5087,N_4705,N_4656);
or U5088 (N_5088,N_4687,N_4846);
nor U5089 (N_5089,N_4688,N_4883);
nor U5090 (N_5090,N_4973,N_4531);
and U5091 (N_5091,N_4694,N_4598);
or U5092 (N_5092,N_4861,N_4825);
nand U5093 (N_5093,N_4588,N_4573);
xor U5094 (N_5094,N_4742,N_4954);
nor U5095 (N_5095,N_4840,N_4872);
and U5096 (N_5096,N_4881,N_4632);
and U5097 (N_5097,N_4606,N_4886);
xor U5098 (N_5098,N_4572,N_4765);
nand U5099 (N_5099,N_4549,N_4734);
nor U5100 (N_5100,N_4834,N_4907);
nand U5101 (N_5101,N_4961,N_4516);
and U5102 (N_5102,N_4704,N_4638);
nand U5103 (N_5103,N_4587,N_4926);
nand U5104 (N_5104,N_4506,N_4753);
nand U5105 (N_5105,N_4794,N_4999);
nor U5106 (N_5106,N_4534,N_4948);
xnor U5107 (N_5107,N_4803,N_4900);
or U5108 (N_5108,N_4680,N_4715);
nand U5109 (N_5109,N_4775,N_4706);
nand U5110 (N_5110,N_4848,N_4513);
xnor U5111 (N_5111,N_4604,N_4532);
and U5112 (N_5112,N_4750,N_4571);
nand U5113 (N_5113,N_4952,N_4621);
nor U5114 (N_5114,N_4574,N_4880);
and U5115 (N_5115,N_4522,N_4546);
or U5116 (N_5116,N_4874,N_4655);
and U5117 (N_5117,N_4657,N_4709);
nor U5118 (N_5118,N_4958,N_4730);
xnor U5119 (N_5119,N_4800,N_4601);
nor U5120 (N_5120,N_4941,N_4508);
xnor U5121 (N_5121,N_4913,N_4682);
xor U5122 (N_5122,N_4663,N_4988);
xor U5123 (N_5123,N_4842,N_4996);
and U5124 (N_5124,N_4623,N_4928);
nand U5125 (N_5125,N_4544,N_4661);
and U5126 (N_5126,N_4761,N_4643);
and U5127 (N_5127,N_4788,N_4637);
nand U5128 (N_5128,N_4569,N_4771);
xnor U5129 (N_5129,N_4798,N_4738);
nand U5130 (N_5130,N_4918,N_4509);
and U5131 (N_5131,N_4700,N_4754);
nor U5132 (N_5132,N_4858,N_4844);
nor U5133 (N_5133,N_4711,N_4809);
or U5134 (N_5134,N_4882,N_4737);
nor U5135 (N_5135,N_4991,N_4801);
nand U5136 (N_5136,N_4828,N_4972);
xor U5137 (N_5137,N_4576,N_4518);
and U5138 (N_5138,N_4831,N_4548);
and U5139 (N_5139,N_4628,N_4563);
or U5140 (N_5140,N_4618,N_4609);
and U5141 (N_5141,N_4967,N_4690);
nand U5142 (N_5142,N_4970,N_4935);
xor U5143 (N_5143,N_4708,N_4591);
nor U5144 (N_5144,N_4797,N_4841);
and U5145 (N_5145,N_4837,N_4593);
and U5146 (N_5146,N_4793,N_4947);
and U5147 (N_5147,N_4558,N_4904);
nor U5148 (N_5148,N_4630,N_4617);
and U5149 (N_5149,N_4678,N_4674);
nand U5150 (N_5150,N_4639,N_4681);
or U5151 (N_5151,N_4726,N_4671);
xnor U5152 (N_5152,N_4855,N_4971);
xor U5153 (N_5153,N_4502,N_4749);
xnor U5154 (N_5154,N_4567,N_4804);
nor U5155 (N_5155,N_4752,N_4993);
xnor U5156 (N_5156,N_4595,N_4652);
xnor U5157 (N_5157,N_4897,N_4786);
nor U5158 (N_5158,N_4924,N_4811);
nand U5159 (N_5159,N_4613,N_4602);
xnor U5160 (N_5160,N_4600,N_4620);
or U5161 (N_5161,N_4728,N_4698);
xor U5162 (N_5162,N_4545,N_4693);
nor U5163 (N_5163,N_4823,N_4504);
xor U5164 (N_5164,N_4744,N_4641);
and U5165 (N_5165,N_4510,N_4830);
or U5166 (N_5166,N_4556,N_4983);
or U5167 (N_5167,N_4878,N_4916);
nor U5168 (N_5168,N_4691,N_4871);
and U5169 (N_5169,N_4851,N_4873);
or U5170 (N_5170,N_4543,N_4901);
nor U5171 (N_5171,N_4648,N_4515);
nor U5172 (N_5172,N_4542,N_4583);
nor U5173 (N_5173,N_4608,N_4714);
nand U5174 (N_5174,N_4850,N_4697);
and U5175 (N_5175,N_4827,N_4729);
nand U5176 (N_5176,N_4683,N_4647);
and U5177 (N_5177,N_4759,N_4653);
or U5178 (N_5178,N_4845,N_4553);
or U5179 (N_5179,N_4933,N_4701);
xnor U5180 (N_5180,N_4962,N_4659);
or U5181 (N_5181,N_4710,N_4995);
nand U5182 (N_5182,N_4783,N_4616);
nand U5183 (N_5183,N_4584,N_4629);
or U5184 (N_5184,N_4521,N_4619);
nand U5185 (N_5185,N_4669,N_4789);
and U5186 (N_5186,N_4835,N_4791);
nand U5187 (N_5187,N_4594,N_4724);
xnor U5188 (N_5188,N_4956,N_4909);
nor U5189 (N_5189,N_4511,N_4646);
or U5190 (N_5190,N_4959,N_4627);
nor U5191 (N_5191,N_4859,N_4856);
or U5192 (N_5192,N_4696,N_4739);
xor U5193 (N_5193,N_4614,N_4756);
or U5194 (N_5194,N_4808,N_4953);
xnor U5195 (N_5195,N_4869,N_4955);
nor U5196 (N_5196,N_4899,N_4713);
nor U5197 (N_5197,N_4603,N_4805);
nor U5198 (N_5198,N_4839,N_4950);
nor U5199 (N_5199,N_4919,N_4792);
nand U5200 (N_5200,N_4679,N_4684);
nand U5201 (N_5201,N_4634,N_4636);
and U5202 (N_5202,N_4733,N_4990);
or U5203 (N_5203,N_4936,N_4816);
or U5204 (N_5204,N_4903,N_4660);
xor U5205 (N_5205,N_4884,N_4667);
and U5206 (N_5206,N_4994,N_4914);
xor U5207 (N_5207,N_4836,N_4668);
nor U5208 (N_5208,N_4640,N_4586);
nand U5209 (N_5209,N_4672,N_4921);
and U5210 (N_5210,N_4932,N_4870);
nand U5211 (N_5211,N_4675,N_4770);
and U5212 (N_5212,N_4766,N_4589);
nand U5213 (N_5213,N_4922,N_4559);
nor U5214 (N_5214,N_4795,N_4666);
and U5215 (N_5215,N_4747,N_4610);
or U5216 (N_5216,N_4523,N_4868);
xor U5217 (N_5217,N_4547,N_4702);
xor U5218 (N_5218,N_4565,N_4814);
nand U5219 (N_5219,N_4905,N_4992);
and U5220 (N_5220,N_4533,N_4923);
nor U5221 (N_5221,N_4712,N_4969);
or U5222 (N_5222,N_4560,N_4605);
nor U5223 (N_5223,N_4917,N_4566);
xnor U5224 (N_5224,N_4642,N_4877);
nor U5225 (N_5225,N_4597,N_4894);
or U5226 (N_5226,N_4517,N_4847);
and U5227 (N_5227,N_4885,N_4938);
or U5228 (N_5228,N_4736,N_4746);
xor U5229 (N_5229,N_4802,N_4626);
nor U5230 (N_5230,N_4888,N_4817);
and U5231 (N_5231,N_4685,N_4520);
and U5232 (N_5232,N_4838,N_4832);
xor U5233 (N_5233,N_4581,N_4976);
nand U5234 (N_5234,N_4529,N_4998);
or U5235 (N_5235,N_4849,N_4748);
xnor U5236 (N_5236,N_4512,N_4876);
xnor U5237 (N_5237,N_4575,N_4978);
xor U5238 (N_5238,N_4550,N_4902);
xor U5239 (N_5239,N_4889,N_4780);
and U5240 (N_5240,N_4799,N_4536);
nor U5241 (N_5241,N_4920,N_4615);
or U5242 (N_5242,N_4535,N_4776);
nor U5243 (N_5243,N_4670,N_4787);
or U5244 (N_5244,N_4686,N_4864);
nor U5245 (N_5245,N_4985,N_4975);
nand U5246 (N_5246,N_4721,N_4937);
and U5247 (N_5247,N_4719,N_4662);
nand U5248 (N_5248,N_4779,N_4875);
xor U5249 (N_5249,N_4946,N_4607);
xnor U5250 (N_5250,N_4710,N_4679);
nand U5251 (N_5251,N_4873,N_4918);
or U5252 (N_5252,N_4956,N_4878);
and U5253 (N_5253,N_4753,N_4646);
nand U5254 (N_5254,N_4706,N_4744);
nor U5255 (N_5255,N_4991,N_4921);
nand U5256 (N_5256,N_4626,N_4992);
nand U5257 (N_5257,N_4677,N_4806);
xnor U5258 (N_5258,N_4569,N_4650);
and U5259 (N_5259,N_4547,N_4735);
and U5260 (N_5260,N_4536,N_4569);
nor U5261 (N_5261,N_4994,N_4805);
nor U5262 (N_5262,N_4724,N_4706);
xor U5263 (N_5263,N_4651,N_4985);
or U5264 (N_5264,N_4775,N_4947);
nor U5265 (N_5265,N_4590,N_4572);
nand U5266 (N_5266,N_4601,N_4625);
nor U5267 (N_5267,N_4506,N_4598);
nand U5268 (N_5268,N_4794,N_4681);
or U5269 (N_5269,N_4690,N_4681);
xor U5270 (N_5270,N_4647,N_4949);
xnor U5271 (N_5271,N_4724,N_4792);
nand U5272 (N_5272,N_4773,N_4995);
or U5273 (N_5273,N_4648,N_4606);
and U5274 (N_5274,N_4747,N_4887);
and U5275 (N_5275,N_4526,N_4805);
xnor U5276 (N_5276,N_4924,N_4965);
and U5277 (N_5277,N_4786,N_4716);
nand U5278 (N_5278,N_4668,N_4636);
or U5279 (N_5279,N_4554,N_4551);
nand U5280 (N_5280,N_4777,N_4772);
and U5281 (N_5281,N_4877,N_4757);
and U5282 (N_5282,N_4912,N_4765);
xnor U5283 (N_5283,N_4602,N_4745);
xnor U5284 (N_5284,N_4671,N_4511);
xnor U5285 (N_5285,N_4614,N_4905);
nand U5286 (N_5286,N_4678,N_4739);
nand U5287 (N_5287,N_4760,N_4822);
xnor U5288 (N_5288,N_4949,N_4602);
xnor U5289 (N_5289,N_4786,N_4638);
and U5290 (N_5290,N_4651,N_4898);
or U5291 (N_5291,N_4803,N_4688);
nand U5292 (N_5292,N_4903,N_4605);
nand U5293 (N_5293,N_4689,N_4793);
nand U5294 (N_5294,N_4962,N_4596);
and U5295 (N_5295,N_4778,N_4841);
xor U5296 (N_5296,N_4620,N_4836);
xor U5297 (N_5297,N_4986,N_4643);
xor U5298 (N_5298,N_4550,N_4820);
nand U5299 (N_5299,N_4778,N_4601);
nand U5300 (N_5300,N_4731,N_4656);
and U5301 (N_5301,N_4680,N_4892);
nand U5302 (N_5302,N_4804,N_4812);
xnor U5303 (N_5303,N_4556,N_4503);
nand U5304 (N_5304,N_4648,N_4940);
xnor U5305 (N_5305,N_4975,N_4956);
xnor U5306 (N_5306,N_4841,N_4783);
nand U5307 (N_5307,N_4577,N_4603);
nand U5308 (N_5308,N_4890,N_4718);
nand U5309 (N_5309,N_4824,N_4777);
or U5310 (N_5310,N_4906,N_4915);
and U5311 (N_5311,N_4732,N_4972);
and U5312 (N_5312,N_4624,N_4670);
or U5313 (N_5313,N_4696,N_4600);
nand U5314 (N_5314,N_4665,N_4798);
and U5315 (N_5315,N_4787,N_4646);
xor U5316 (N_5316,N_4752,N_4847);
nor U5317 (N_5317,N_4541,N_4806);
nand U5318 (N_5318,N_4719,N_4834);
nor U5319 (N_5319,N_4780,N_4784);
xor U5320 (N_5320,N_4954,N_4606);
and U5321 (N_5321,N_4547,N_4711);
nor U5322 (N_5322,N_4817,N_4826);
or U5323 (N_5323,N_4754,N_4505);
nor U5324 (N_5324,N_4792,N_4628);
xor U5325 (N_5325,N_4676,N_4834);
or U5326 (N_5326,N_4557,N_4533);
nor U5327 (N_5327,N_4804,N_4646);
nand U5328 (N_5328,N_4974,N_4894);
xor U5329 (N_5329,N_4782,N_4628);
nand U5330 (N_5330,N_4648,N_4636);
nor U5331 (N_5331,N_4744,N_4614);
and U5332 (N_5332,N_4672,N_4782);
and U5333 (N_5333,N_4817,N_4640);
or U5334 (N_5334,N_4782,N_4664);
nor U5335 (N_5335,N_4969,N_4519);
or U5336 (N_5336,N_4588,N_4671);
or U5337 (N_5337,N_4655,N_4900);
nor U5338 (N_5338,N_4768,N_4704);
xor U5339 (N_5339,N_4756,N_4811);
or U5340 (N_5340,N_4691,N_4758);
xnor U5341 (N_5341,N_4776,N_4942);
nand U5342 (N_5342,N_4578,N_4776);
or U5343 (N_5343,N_4895,N_4572);
nand U5344 (N_5344,N_4857,N_4717);
xor U5345 (N_5345,N_4585,N_4733);
xnor U5346 (N_5346,N_4965,N_4520);
nand U5347 (N_5347,N_4969,N_4804);
or U5348 (N_5348,N_4587,N_4901);
or U5349 (N_5349,N_4724,N_4684);
and U5350 (N_5350,N_4593,N_4852);
or U5351 (N_5351,N_4869,N_4777);
and U5352 (N_5352,N_4968,N_4690);
or U5353 (N_5353,N_4506,N_4605);
nor U5354 (N_5354,N_4917,N_4641);
and U5355 (N_5355,N_4742,N_4541);
nor U5356 (N_5356,N_4557,N_4954);
and U5357 (N_5357,N_4781,N_4910);
and U5358 (N_5358,N_4729,N_4640);
nand U5359 (N_5359,N_4807,N_4858);
or U5360 (N_5360,N_4836,N_4800);
xor U5361 (N_5361,N_4907,N_4523);
xnor U5362 (N_5362,N_4869,N_4774);
and U5363 (N_5363,N_4832,N_4780);
nand U5364 (N_5364,N_4954,N_4528);
and U5365 (N_5365,N_4982,N_4892);
nor U5366 (N_5366,N_4930,N_4694);
and U5367 (N_5367,N_4661,N_4982);
nand U5368 (N_5368,N_4575,N_4659);
nor U5369 (N_5369,N_4689,N_4948);
xnor U5370 (N_5370,N_4765,N_4650);
nor U5371 (N_5371,N_4936,N_4812);
or U5372 (N_5372,N_4533,N_4639);
nor U5373 (N_5373,N_4630,N_4509);
or U5374 (N_5374,N_4683,N_4664);
nor U5375 (N_5375,N_4861,N_4754);
xnor U5376 (N_5376,N_4835,N_4908);
or U5377 (N_5377,N_4814,N_4656);
nand U5378 (N_5378,N_4596,N_4934);
nor U5379 (N_5379,N_4800,N_4622);
nand U5380 (N_5380,N_4505,N_4810);
nand U5381 (N_5381,N_4904,N_4949);
nand U5382 (N_5382,N_4801,N_4715);
or U5383 (N_5383,N_4889,N_4670);
nand U5384 (N_5384,N_4635,N_4547);
nor U5385 (N_5385,N_4872,N_4873);
nand U5386 (N_5386,N_4790,N_4743);
and U5387 (N_5387,N_4528,N_4684);
or U5388 (N_5388,N_4842,N_4754);
and U5389 (N_5389,N_4956,N_4794);
nor U5390 (N_5390,N_4702,N_4724);
nand U5391 (N_5391,N_4639,N_4894);
xor U5392 (N_5392,N_4892,N_4764);
or U5393 (N_5393,N_4753,N_4631);
xor U5394 (N_5394,N_4635,N_4525);
nand U5395 (N_5395,N_4604,N_4588);
or U5396 (N_5396,N_4662,N_4622);
nor U5397 (N_5397,N_4635,N_4913);
xor U5398 (N_5398,N_4840,N_4884);
xnor U5399 (N_5399,N_4606,N_4575);
nand U5400 (N_5400,N_4943,N_4650);
nand U5401 (N_5401,N_4534,N_4907);
and U5402 (N_5402,N_4960,N_4865);
nor U5403 (N_5403,N_4928,N_4593);
and U5404 (N_5404,N_4832,N_4894);
nand U5405 (N_5405,N_4500,N_4701);
nor U5406 (N_5406,N_4602,N_4941);
and U5407 (N_5407,N_4879,N_4850);
or U5408 (N_5408,N_4660,N_4577);
or U5409 (N_5409,N_4588,N_4643);
nor U5410 (N_5410,N_4535,N_4676);
or U5411 (N_5411,N_4827,N_4660);
or U5412 (N_5412,N_4979,N_4513);
nor U5413 (N_5413,N_4887,N_4618);
nor U5414 (N_5414,N_4562,N_4780);
and U5415 (N_5415,N_4856,N_4993);
nor U5416 (N_5416,N_4533,N_4581);
nand U5417 (N_5417,N_4811,N_4748);
and U5418 (N_5418,N_4904,N_4895);
nor U5419 (N_5419,N_4650,N_4745);
or U5420 (N_5420,N_4563,N_4923);
or U5421 (N_5421,N_4754,N_4880);
nand U5422 (N_5422,N_4789,N_4916);
nor U5423 (N_5423,N_4885,N_4631);
xnor U5424 (N_5424,N_4799,N_4917);
nor U5425 (N_5425,N_4861,N_4649);
nor U5426 (N_5426,N_4832,N_4979);
nand U5427 (N_5427,N_4972,N_4871);
and U5428 (N_5428,N_4561,N_4849);
and U5429 (N_5429,N_4523,N_4962);
and U5430 (N_5430,N_4574,N_4605);
or U5431 (N_5431,N_4965,N_4921);
or U5432 (N_5432,N_4674,N_4757);
nor U5433 (N_5433,N_4962,N_4812);
and U5434 (N_5434,N_4532,N_4661);
nand U5435 (N_5435,N_4778,N_4774);
or U5436 (N_5436,N_4545,N_4819);
nor U5437 (N_5437,N_4821,N_4655);
xor U5438 (N_5438,N_4698,N_4730);
or U5439 (N_5439,N_4797,N_4571);
or U5440 (N_5440,N_4853,N_4761);
or U5441 (N_5441,N_4502,N_4824);
and U5442 (N_5442,N_4509,N_4762);
and U5443 (N_5443,N_4903,N_4765);
nand U5444 (N_5444,N_4567,N_4575);
and U5445 (N_5445,N_4945,N_4662);
or U5446 (N_5446,N_4673,N_4993);
and U5447 (N_5447,N_4862,N_4666);
xnor U5448 (N_5448,N_4618,N_4870);
nor U5449 (N_5449,N_4763,N_4649);
and U5450 (N_5450,N_4719,N_4803);
nor U5451 (N_5451,N_4749,N_4764);
or U5452 (N_5452,N_4745,N_4943);
nor U5453 (N_5453,N_4579,N_4582);
nor U5454 (N_5454,N_4965,N_4525);
or U5455 (N_5455,N_4774,N_4588);
and U5456 (N_5456,N_4744,N_4604);
nand U5457 (N_5457,N_4796,N_4782);
or U5458 (N_5458,N_4710,N_4546);
nor U5459 (N_5459,N_4923,N_4787);
nor U5460 (N_5460,N_4937,N_4897);
xor U5461 (N_5461,N_4630,N_4743);
or U5462 (N_5462,N_4809,N_4572);
nand U5463 (N_5463,N_4989,N_4736);
and U5464 (N_5464,N_4572,N_4969);
xor U5465 (N_5465,N_4703,N_4543);
and U5466 (N_5466,N_4794,N_4722);
nor U5467 (N_5467,N_4797,N_4735);
xnor U5468 (N_5468,N_4603,N_4684);
xnor U5469 (N_5469,N_4586,N_4618);
and U5470 (N_5470,N_4878,N_4989);
nor U5471 (N_5471,N_4957,N_4747);
and U5472 (N_5472,N_4672,N_4816);
or U5473 (N_5473,N_4845,N_4870);
nor U5474 (N_5474,N_4633,N_4585);
nor U5475 (N_5475,N_4981,N_4881);
or U5476 (N_5476,N_4968,N_4822);
nor U5477 (N_5477,N_4910,N_4558);
or U5478 (N_5478,N_4627,N_4982);
and U5479 (N_5479,N_4757,N_4632);
nor U5480 (N_5480,N_4614,N_4561);
nor U5481 (N_5481,N_4922,N_4897);
nor U5482 (N_5482,N_4960,N_4607);
nor U5483 (N_5483,N_4814,N_4589);
nand U5484 (N_5484,N_4917,N_4894);
xor U5485 (N_5485,N_4747,N_4902);
or U5486 (N_5486,N_4559,N_4968);
nand U5487 (N_5487,N_4881,N_4856);
nand U5488 (N_5488,N_4535,N_4878);
and U5489 (N_5489,N_4621,N_4987);
nand U5490 (N_5490,N_4885,N_4886);
xor U5491 (N_5491,N_4598,N_4923);
and U5492 (N_5492,N_4939,N_4604);
or U5493 (N_5493,N_4579,N_4847);
or U5494 (N_5494,N_4770,N_4696);
nand U5495 (N_5495,N_4699,N_4645);
nand U5496 (N_5496,N_4985,N_4885);
and U5497 (N_5497,N_4834,N_4780);
or U5498 (N_5498,N_4573,N_4595);
or U5499 (N_5499,N_4596,N_4675);
xor U5500 (N_5500,N_5304,N_5406);
and U5501 (N_5501,N_5374,N_5072);
xnor U5502 (N_5502,N_5273,N_5239);
nand U5503 (N_5503,N_5266,N_5367);
or U5504 (N_5504,N_5372,N_5308);
nor U5505 (N_5505,N_5431,N_5134);
and U5506 (N_5506,N_5340,N_5172);
nand U5507 (N_5507,N_5133,N_5456);
xor U5508 (N_5508,N_5307,N_5389);
nor U5509 (N_5509,N_5339,N_5489);
and U5510 (N_5510,N_5199,N_5334);
nand U5511 (N_5511,N_5320,N_5143);
and U5512 (N_5512,N_5426,N_5032);
xnor U5513 (N_5513,N_5238,N_5263);
and U5514 (N_5514,N_5162,N_5355);
nor U5515 (N_5515,N_5121,N_5182);
xor U5516 (N_5516,N_5354,N_5081);
or U5517 (N_5517,N_5341,N_5042);
nand U5518 (N_5518,N_5119,N_5325);
nor U5519 (N_5519,N_5045,N_5030);
xnor U5520 (N_5520,N_5436,N_5262);
nand U5521 (N_5521,N_5327,N_5402);
and U5522 (N_5522,N_5346,N_5074);
nand U5523 (N_5523,N_5382,N_5094);
and U5524 (N_5524,N_5107,N_5386);
xor U5525 (N_5525,N_5015,N_5190);
nor U5526 (N_5526,N_5328,N_5314);
nand U5527 (N_5527,N_5113,N_5069);
or U5528 (N_5528,N_5318,N_5139);
and U5529 (N_5529,N_5211,N_5446);
and U5530 (N_5530,N_5159,N_5366);
xnor U5531 (N_5531,N_5203,N_5135);
nor U5532 (N_5532,N_5451,N_5319);
nor U5533 (N_5533,N_5153,N_5175);
xor U5534 (N_5534,N_5118,N_5324);
and U5535 (N_5535,N_5050,N_5394);
nor U5536 (N_5536,N_5057,N_5039);
xor U5537 (N_5537,N_5380,N_5112);
xor U5538 (N_5538,N_5071,N_5195);
nand U5539 (N_5539,N_5412,N_5260);
and U5540 (N_5540,N_5067,N_5192);
xnor U5541 (N_5541,N_5427,N_5458);
and U5542 (N_5542,N_5053,N_5255);
and U5543 (N_5543,N_5157,N_5124);
nand U5544 (N_5544,N_5205,N_5493);
nor U5545 (N_5545,N_5230,N_5087);
and U5546 (N_5546,N_5197,N_5289);
nand U5547 (N_5547,N_5046,N_5261);
nor U5548 (N_5548,N_5010,N_5496);
nand U5549 (N_5549,N_5006,N_5200);
nor U5550 (N_5550,N_5132,N_5165);
xor U5551 (N_5551,N_5375,N_5299);
and U5552 (N_5552,N_5467,N_5477);
xnor U5553 (N_5553,N_5189,N_5114);
or U5554 (N_5554,N_5193,N_5158);
xnor U5555 (N_5555,N_5103,N_5061);
xor U5556 (N_5556,N_5237,N_5288);
nand U5557 (N_5557,N_5123,N_5129);
and U5558 (N_5558,N_5098,N_5450);
nand U5559 (N_5559,N_5198,N_5399);
and U5560 (N_5560,N_5387,N_5208);
xnor U5561 (N_5561,N_5350,N_5429);
or U5562 (N_5562,N_5176,N_5016);
nor U5563 (N_5563,N_5309,N_5358);
or U5564 (N_5564,N_5316,N_5178);
and U5565 (N_5565,N_5290,N_5240);
and U5566 (N_5566,N_5023,N_5228);
and U5567 (N_5567,N_5322,N_5014);
or U5568 (N_5568,N_5302,N_5227);
nand U5569 (N_5569,N_5131,N_5225);
and U5570 (N_5570,N_5416,N_5461);
and U5571 (N_5571,N_5156,N_5422);
and U5572 (N_5572,N_5330,N_5108);
nor U5573 (N_5573,N_5438,N_5149);
nor U5574 (N_5574,N_5365,N_5086);
nand U5575 (N_5575,N_5463,N_5278);
nor U5576 (N_5576,N_5002,N_5017);
nand U5577 (N_5577,N_5277,N_5167);
or U5578 (N_5578,N_5281,N_5472);
or U5579 (N_5579,N_5474,N_5210);
and U5580 (N_5580,N_5020,N_5441);
or U5581 (N_5581,N_5353,N_5130);
and U5582 (N_5582,N_5024,N_5483);
or U5583 (N_5583,N_5233,N_5056);
nor U5584 (N_5584,N_5494,N_5226);
and U5585 (N_5585,N_5116,N_5005);
nand U5586 (N_5586,N_5095,N_5469);
nand U5587 (N_5587,N_5491,N_5012);
nor U5588 (N_5588,N_5435,N_5070);
nor U5589 (N_5589,N_5419,N_5151);
nand U5590 (N_5590,N_5055,N_5004);
or U5591 (N_5591,N_5425,N_5078);
xnor U5592 (N_5592,N_5183,N_5311);
nand U5593 (N_5593,N_5241,N_5079);
or U5594 (N_5594,N_5455,N_5284);
or U5595 (N_5595,N_5082,N_5404);
and U5596 (N_5596,N_5246,N_5342);
xor U5597 (N_5597,N_5044,N_5499);
nor U5598 (N_5598,N_5091,N_5173);
nand U5599 (N_5599,N_5076,N_5373);
nand U5600 (N_5600,N_5000,N_5329);
and U5601 (N_5601,N_5344,N_5312);
and U5602 (N_5602,N_5393,N_5473);
nor U5603 (N_5603,N_5080,N_5388);
nand U5604 (N_5604,N_5191,N_5092);
nand U5605 (N_5605,N_5279,N_5047);
nor U5606 (N_5606,N_5084,N_5478);
xor U5607 (N_5607,N_5206,N_5457);
xnor U5608 (N_5608,N_5338,N_5267);
nand U5609 (N_5609,N_5317,N_5185);
nor U5610 (N_5610,N_5378,N_5126);
and U5611 (N_5611,N_5180,N_5110);
nor U5612 (N_5612,N_5171,N_5048);
xor U5613 (N_5613,N_5009,N_5440);
nor U5614 (N_5614,N_5088,N_5271);
or U5615 (N_5615,N_5144,N_5305);
and U5616 (N_5616,N_5482,N_5270);
xor U5617 (N_5617,N_5101,N_5383);
xor U5618 (N_5618,N_5407,N_5424);
or U5619 (N_5619,N_5213,N_5253);
nand U5620 (N_5620,N_5054,N_5259);
xnor U5621 (N_5621,N_5034,N_5306);
nor U5622 (N_5622,N_5298,N_5218);
nor U5623 (N_5623,N_5196,N_5036);
nor U5624 (N_5624,N_5276,N_5128);
nand U5625 (N_5625,N_5408,N_5075);
nor U5626 (N_5626,N_5498,N_5220);
or U5627 (N_5627,N_5038,N_5186);
nor U5628 (N_5628,N_5377,N_5332);
or U5629 (N_5629,N_5464,N_5035);
xnor U5630 (N_5630,N_5179,N_5235);
nor U5631 (N_5631,N_5013,N_5359);
xnor U5632 (N_5632,N_5083,N_5452);
nor U5633 (N_5633,N_5480,N_5462);
and U5634 (N_5634,N_5117,N_5115);
xnor U5635 (N_5635,N_5364,N_5466);
xnor U5636 (N_5636,N_5140,N_5242);
nor U5637 (N_5637,N_5150,N_5100);
and U5638 (N_5638,N_5428,N_5099);
and U5639 (N_5639,N_5247,N_5037);
or U5640 (N_5640,N_5202,N_5174);
xor U5641 (N_5641,N_5326,N_5421);
xnor U5642 (N_5642,N_5357,N_5252);
nand U5643 (N_5643,N_5184,N_5043);
and U5644 (N_5644,N_5137,N_5291);
and U5645 (N_5645,N_5019,N_5488);
or U5646 (N_5646,N_5219,N_5418);
and U5647 (N_5647,N_5315,N_5122);
nor U5648 (N_5648,N_5430,N_5410);
nand U5649 (N_5649,N_5348,N_5077);
or U5650 (N_5650,N_5105,N_5396);
and U5651 (N_5651,N_5148,N_5433);
or U5652 (N_5652,N_5345,N_5217);
nor U5653 (N_5653,N_5347,N_5155);
and U5654 (N_5654,N_5363,N_5296);
and U5655 (N_5655,N_5468,N_5286);
nand U5656 (N_5656,N_5106,N_5384);
or U5657 (N_5657,N_5160,N_5275);
xnor U5658 (N_5658,N_5025,N_5381);
or U5659 (N_5659,N_5147,N_5164);
or U5660 (N_5660,N_5360,N_5026);
or U5661 (N_5661,N_5411,N_5254);
nor U5662 (N_5662,N_5104,N_5244);
or U5663 (N_5663,N_5051,N_5215);
or U5664 (N_5664,N_5371,N_5204);
nand U5665 (N_5665,N_5449,N_5181);
nand U5666 (N_5666,N_5370,N_5479);
nor U5667 (N_5667,N_5362,N_5231);
and U5668 (N_5668,N_5052,N_5064);
and U5669 (N_5669,N_5194,N_5287);
xnor U5670 (N_5670,N_5249,N_5391);
nand U5671 (N_5671,N_5187,N_5397);
xnor U5672 (N_5672,N_5297,N_5285);
and U5673 (N_5673,N_5403,N_5090);
nor U5674 (N_5674,N_5434,N_5352);
nand U5675 (N_5675,N_5018,N_5413);
and U5676 (N_5676,N_5001,N_5487);
nor U5677 (N_5677,N_5414,N_5216);
nor U5678 (N_5678,N_5447,N_5368);
nand U5679 (N_5679,N_5432,N_5400);
xor U5680 (N_5680,N_5321,N_5398);
nor U5681 (N_5681,N_5258,N_5243);
nand U5682 (N_5682,N_5136,N_5283);
nor U5683 (N_5683,N_5027,N_5093);
nand U5684 (N_5684,N_5442,N_5395);
nor U5685 (N_5685,N_5207,N_5303);
or U5686 (N_5686,N_5439,N_5146);
and U5687 (N_5687,N_5265,N_5420);
and U5688 (N_5688,N_5059,N_5465);
nor U5689 (N_5689,N_5484,N_5021);
nor U5690 (N_5690,N_5120,N_5063);
xor U5691 (N_5691,N_5471,N_5229);
nand U5692 (N_5692,N_5470,N_5343);
xnor U5693 (N_5693,N_5268,N_5029);
or U5694 (N_5694,N_5379,N_5356);
nor U5695 (N_5695,N_5476,N_5138);
nor U5696 (N_5696,N_5385,N_5066);
xnor U5697 (N_5697,N_5111,N_5096);
and U5698 (N_5698,N_5481,N_5495);
and U5699 (N_5699,N_5392,N_5033);
or U5700 (N_5700,N_5448,N_5443);
and U5701 (N_5701,N_5201,N_5269);
nand U5702 (N_5702,N_5444,N_5336);
nor U5703 (N_5703,N_5323,N_5351);
or U5704 (N_5704,N_5089,N_5486);
nand U5705 (N_5705,N_5460,N_5065);
nand U5706 (N_5706,N_5223,N_5068);
nor U5707 (N_5707,N_5141,N_5282);
or U5708 (N_5708,N_5154,N_5011);
xnor U5709 (N_5709,N_5295,N_5166);
or U5710 (N_5710,N_5280,N_5453);
and U5711 (N_5711,N_5293,N_5369);
xnor U5712 (N_5712,N_5177,N_5008);
xor U5713 (N_5713,N_5337,N_5170);
xor U5714 (N_5714,N_5142,N_5248);
nand U5715 (N_5715,N_5349,N_5445);
nand U5716 (N_5716,N_5292,N_5188);
nand U5717 (N_5717,N_5245,N_5028);
and U5718 (N_5718,N_5301,N_5485);
and U5719 (N_5719,N_5007,N_5003);
xor U5720 (N_5720,N_5361,N_5221);
or U5721 (N_5721,N_5073,N_5031);
and U5722 (N_5722,N_5168,N_5209);
nor U5723 (N_5723,N_5475,N_5152);
or U5724 (N_5724,N_5390,N_5423);
nor U5725 (N_5725,N_5294,N_5212);
nor U5726 (N_5726,N_5145,N_5163);
and U5727 (N_5727,N_5049,N_5125);
and U5728 (N_5728,N_5331,N_5401);
nand U5729 (N_5729,N_5251,N_5097);
nor U5730 (N_5730,N_5060,N_5256);
nand U5731 (N_5731,N_5300,N_5333);
nand U5732 (N_5732,N_5415,N_5127);
xor U5733 (N_5733,N_5214,N_5222);
or U5734 (N_5734,N_5161,N_5459);
or U5735 (N_5735,N_5041,N_5058);
nor U5736 (N_5736,N_5272,N_5062);
nand U5737 (N_5737,N_5274,N_5313);
and U5738 (N_5738,N_5490,N_5169);
and U5739 (N_5739,N_5376,N_5022);
xor U5740 (N_5740,N_5085,N_5409);
and U5741 (N_5741,N_5109,N_5405);
xnor U5742 (N_5742,N_5234,N_5102);
xor U5743 (N_5743,N_5492,N_5224);
and U5744 (N_5744,N_5250,N_5497);
nor U5745 (N_5745,N_5236,N_5454);
and U5746 (N_5746,N_5417,N_5335);
or U5747 (N_5747,N_5040,N_5310);
and U5748 (N_5748,N_5257,N_5232);
xor U5749 (N_5749,N_5437,N_5264);
and U5750 (N_5750,N_5298,N_5482);
nand U5751 (N_5751,N_5233,N_5379);
or U5752 (N_5752,N_5244,N_5049);
or U5753 (N_5753,N_5071,N_5426);
xor U5754 (N_5754,N_5045,N_5192);
nor U5755 (N_5755,N_5314,N_5085);
or U5756 (N_5756,N_5141,N_5387);
xor U5757 (N_5757,N_5397,N_5273);
nor U5758 (N_5758,N_5484,N_5094);
nand U5759 (N_5759,N_5061,N_5002);
xor U5760 (N_5760,N_5162,N_5405);
xor U5761 (N_5761,N_5158,N_5426);
or U5762 (N_5762,N_5058,N_5421);
xor U5763 (N_5763,N_5494,N_5343);
and U5764 (N_5764,N_5099,N_5289);
nor U5765 (N_5765,N_5305,N_5435);
xnor U5766 (N_5766,N_5194,N_5488);
nor U5767 (N_5767,N_5016,N_5216);
and U5768 (N_5768,N_5197,N_5285);
nand U5769 (N_5769,N_5477,N_5213);
and U5770 (N_5770,N_5461,N_5264);
nor U5771 (N_5771,N_5183,N_5019);
nor U5772 (N_5772,N_5361,N_5051);
nor U5773 (N_5773,N_5239,N_5164);
or U5774 (N_5774,N_5294,N_5388);
or U5775 (N_5775,N_5462,N_5319);
and U5776 (N_5776,N_5481,N_5244);
nand U5777 (N_5777,N_5345,N_5288);
or U5778 (N_5778,N_5492,N_5238);
and U5779 (N_5779,N_5045,N_5054);
or U5780 (N_5780,N_5208,N_5321);
or U5781 (N_5781,N_5172,N_5147);
nor U5782 (N_5782,N_5131,N_5401);
or U5783 (N_5783,N_5208,N_5246);
or U5784 (N_5784,N_5311,N_5367);
and U5785 (N_5785,N_5168,N_5179);
xor U5786 (N_5786,N_5485,N_5424);
and U5787 (N_5787,N_5067,N_5019);
or U5788 (N_5788,N_5384,N_5162);
nand U5789 (N_5789,N_5150,N_5445);
xnor U5790 (N_5790,N_5282,N_5166);
nand U5791 (N_5791,N_5163,N_5196);
nor U5792 (N_5792,N_5120,N_5219);
and U5793 (N_5793,N_5476,N_5260);
nor U5794 (N_5794,N_5098,N_5499);
and U5795 (N_5795,N_5380,N_5276);
nand U5796 (N_5796,N_5247,N_5133);
and U5797 (N_5797,N_5064,N_5372);
or U5798 (N_5798,N_5390,N_5229);
or U5799 (N_5799,N_5293,N_5365);
nor U5800 (N_5800,N_5022,N_5131);
nor U5801 (N_5801,N_5415,N_5215);
nand U5802 (N_5802,N_5049,N_5144);
and U5803 (N_5803,N_5439,N_5350);
xor U5804 (N_5804,N_5109,N_5428);
xor U5805 (N_5805,N_5241,N_5499);
nor U5806 (N_5806,N_5260,N_5219);
and U5807 (N_5807,N_5006,N_5487);
or U5808 (N_5808,N_5399,N_5248);
xor U5809 (N_5809,N_5180,N_5055);
or U5810 (N_5810,N_5487,N_5206);
xor U5811 (N_5811,N_5314,N_5143);
xor U5812 (N_5812,N_5078,N_5284);
nand U5813 (N_5813,N_5289,N_5294);
and U5814 (N_5814,N_5172,N_5294);
and U5815 (N_5815,N_5086,N_5284);
nor U5816 (N_5816,N_5075,N_5453);
and U5817 (N_5817,N_5175,N_5412);
nor U5818 (N_5818,N_5393,N_5183);
nor U5819 (N_5819,N_5015,N_5298);
nand U5820 (N_5820,N_5083,N_5466);
nand U5821 (N_5821,N_5102,N_5459);
or U5822 (N_5822,N_5172,N_5010);
and U5823 (N_5823,N_5441,N_5088);
and U5824 (N_5824,N_5115,N_5335);
and U5825 (N_5825,N_5135,N_5098);
nor U5826 (N_5826,N_5333,N_5491);
nor U5827 (N_5827,N_5351,N_5372);
nand U5828 (N_5828,N_5409,N_5255);
xor U5829 (N_5829,N_5270,N_5074);
xor U5830 (N_5830,N_5140,N_5039);
or U5831 (N_5831,N_5066,N_5256);
or U5832 (N_5832,N_5252,N_5496);
nor U5833 (N_5833,N_5393,N_5016);
xnor U5834 (N_5834,N_5065,N_5416);
nand U5835 (N_5835,N_5034,N_5448);
or U5836 (N_5836,N_5482,N_5124);
xnor U5837 (N_5837,N_5478,N_5228);
or U5838 (N_5838,N_5038,N_5276);
xor U5839 (N_5839,N_5456,N_5120);
xor U5840 (N_5840,N_5308,N_5176);
xnor U5841 (N_5841,N_5061,N_5269);
nand U5842 (N_5842,N_5065,N_5303);
or U5843 (N_5843,N_5186,N_5277);
xor U5844 (N_5844,N_5420,N_5360);
nor U5845 (N_5845,N_5408,N_5341);
xnor U5846 (N_5846,N_5339,N_5174);
or U5847 (N_5847,N_5477,N_5424);
nor U5848 (N_5848,N_5005,N_5136);
xnor U5849 (N_5849,N_5184,N_5185);
nor U5850 (N_5850,N_5380,N_5279);
nor U5851 (N_5851,N_5495,N_5461);
or U5852 (N_5852,N_5224,N_5435);
and U5853 (N_5853,N_5219,N_5331);
nand U5854 (N_5854,N_5015,N_5496);
and U5855 (N_5855,N_5137,N_5104);
or U5856 (N_5856,N_5137,N_5226);
and U5857 (N_5857,N_5360,N_5175);
nor U5858 (N_5858,N_5499,N_5475);
nor U5859 (N_5859,N_5479,N_5198);
or U5860 (N_5860,N_5391,N_5493);
xor U5861 (N_5861,N_5479,N_5030);
or U5862 (N_5862,N_5131,N_5292);
nor U5863 (N_5863,N_5386,N_5192);
or U5864 (N_5864,N_5114,N_5037);
nor U5865 (N_5865,N_5294,N_5267);
nor U5866 (N_5866,N_5384,N_5309);
nand U5867 (N_5867,N_5025,N_5450);
or U5868 (N_5868,N_5139,N_5065);
or U5869 (N_5869,N_5001,N_5209);
nand U5870 (N_5870,N_5482,N_5479);
nor U5871 (N_5871,N_5469,N_5416);
nand U5872 (N_5872,N_5453,N_5459);
xor U5873 (N_5873,N_5477,N_5280);
nand U5874 (N_5874,N_5205,N_5175);
and U5875 (N_5875,N_5391,N_5121);
xor U5876 (N_5876,N_5412,N_5135);
and U5877 (N_5877,N_5024,N_5091);
and U5878 (N_5878,N_5226,N_5236);
nor U5879 (N_5879,N_5210,N_5439);
or U5880 (N_5880,N_5458,N_5045);
nand U5881 (N_5881,N_5497,N_5323);
and U5882 (N_5882,N_5325,N_5230);
nand U5883 (N_5883,N_5405,N_5477);
xnor U5884 (N_5884,N_5370,N_5407);
nand U5885 (N_5885,N_5271,N_5172);
nand U5886 (N_5886,N_5181,N_5107);
nand U5887 (N_5887,N_5088,N_5282);
nor U5888 (N_5888,N_5248,N_5071);
nor U5889 (N_5889,N_5032,N_5427);
or U5890 (N_5890,N_5284,N_5178);
xor U5891 (N_5891,N_5319,N_5277);
nand U5892 (N_5892,N_5032,N_5174);
and U5893 (N_5893,N_5357,N_5062);
nand U5894 (N_5894,N_5021,N_5007);
and U5895 (N_5895,N_5318,N_5160);
xor U5896 (N_5896,N_5202,N_5229);
xor U5897 (N_5897,N_5208,N_5414);
nand U5898 (N_5898,N_5127,N_5347);
xor U5899 (N_5899,N_5009,N_5154);
nand U5900 (N_5900,N_5344,N_5337);
nor U5901 (N_5901,N_5444,N_5021);
nand U5902 (N_5902,N_5023,N_5377);
nand U5903 (N_5903,N_5323,N_5314);
nor U5904 (N_5904,N_5163,N_5081);
nor U5905 (N_5905,N_5288,N_5348);
nand U5906 (N_5906,N_5400,N_5334);
and U5907 (N_5907,N_5411,N_5070);
and U5908 (N_5908,N_5161,N_5141);
and U5909 (N_5909,N_5456,N_5443);
xnor U5910 (N_5910,N_5261,N_5060);
xnor U5911 (N_5911,N_5487,N_5397);
and U5912 (N_5912,N_5291,N_5062);
nand U5913 (N_5913,N_5078,N_5143);
and U5914 (N_5914,N_5168,N_5313);
xor U5915 (N_5915,N_5315,N_5435);
and U5916 (N_5916,N_5428,N_5410);
nor U5917 (N_5917,N_5461,N_5447);
and U5918 (N_5918,N_5115,N_5237);
xor U5919 (N_5919,N_5248,N_5037);
and U5920 (N_5920,N_5132,N_5335);
xnor U5921 (N_5921,N_5186,N_5346);
xnor U5922 (N_5922,N_5145,N_5406);
and U5923 (N_5923,N_5379,N_5327);
nor U5924 (N_5924,N_5130,N_5144);
xor U5925 (N_5925,N_5289,N_5356);
or U5926 (N_5926,N_5020,N_5254);
or U5927 (N_5927,N_5373,N_5353);
and U5928 (N_5928,N_5375,N_5326);
nor U5929 (N_5929,N_5327,N_5089);
or U5930 (N_5930,N_5269,N_5124);
nand U5931 (N_5931,N_5208,N_5301);
nand U5932 (N_5932,N_5406,N_5140);
nand U5933 (N_5933,N_5294,N_5044);
or U5934 (N_5934,N_5499,N_5075);
nor U5935 (N_5935,N_5065,N_5332);
and U5936 (N_5936,N_5300,N_5356);
and U5937 (N_5937,N_5390,N_5323);
xnor U5938 (N_5938,N_5365,N_5404);
nor U5939 (N_5939,N_5278,N_5110);
nor U5940 (N_5940,N_5402,N_5102);
nand U5941 (N_5941,N_5238,N_5135);
and U5942 (N_5942,N_5061,N_5496);
nor U5943 (N_5943,N_5213,N_5472);
nor U5944 (N_5944,N_5047,N_5119);
and U5945 (N_5945,N_5154,N_5437);
xnor U5946 (N_5946,N_5146,N_5297);
nand U5947 (N_5947,N_5077,N_5040);
or U5948 (N_5948,N_5279,N_5002);
xnor U5949 (N_5949,N_5435,N_5266);
and U5950 (N_5950,N_5288,N_5292);
nand U5951 (N_5951,N_5113,N_5260);
nor U5952 (N_5952,N_5210,N_5059);
nand U5953 (N_5953,N_5492,N_5061);
xnor U5954 (N_5954,N_5215,N_5135);
xor U5955 (N_5955,N_5481,N_5045);
nor U5956 (N_5956,N_5075,N_5188);
and U5957 (N_5957,N_5124,N_5259);
and U5958 (N_5958,N_5234,N_5056);
nor U5959 (N_5959,N_5493,N_5432);
and U5960 (N_5960,N_5263,N_5218);
and U5961 (N_5961,N_5404,N_5017);
and U5962 (N_5962,N_5360,N_5088);
and U5963 (N_5963,N_5297,N_5218);
nor U5964 (N_5964,N_5495,N_5110);
and U5965 (N_5965,N_5029,N_5321);
nand U5966 (N_5966,N_5496,N_5403);
or U5967 (N_5967,N_5377,N_5259);
nand U5968 (N_5968,N_5340,N_5094);
nand U5969 (N_5969,N_5298,N_5364);
nand U5970 (N_5970,N_5091,N_5462);
nand U5971 (N_5971,N_5475,N_5339);
and U5972 (N_5972,N_5373,N_5192);
nor U5973 (N_5973,N_5409,N_5118);
nand U5974 (N_5974,N_5177,N_5312);
nor U5975 (N_5975,N_5444,N_5280);
and U5976 (N_5976,N_5155,N_5424);
and U5977 (N_5977,N_5256,N_5360);
nor U5978 (N_5978,N_5283,N_5341);
nor U5979 (N_5979,N_5107,N_5281);
or U5980 (N_5980,N_5377,N_5499);
nand U5981 (N_5981,N_5240,N_5168);
nor U5982 (N_5982,N_5308,N_5452);
and U5983 (N_5983,N_5471,N_5299);
xor U5984 (N_5984,N_5049,N_5078);
or U5985 (N_5985,N_5420,N_5086);
xor U5986 (N_5986,N_5204,N_5101);
nand U5987 (N_5987,N_5047,N_5461);
nand U5988 (N_5988,N_5317,N_5495);
xor U5989 (N_5989,N_5489,N_5428);
or U5990 (N_5990,N_5485,N_5372);
and U5991 (N_5991,N_5035,N_5477);
or U5992 (N_5992,N_5483,N_5440);
nand U5993 (N_5993,N_5018,N_5073);
nand U5994 (N_5994,N_5421,N_5002);
and U5995 (N_5995,N_5420,N_5213);
nor U5996 (N_5996,N_5044,N_5200);
and U5997 (N_5997,N_5404,N_5241);
and U5998 (N_5998,N_5242,N_5441);
nand U5999 (N_5999,N_5032,N_5144);
or U6000 (N_6000,N_5811,N_5998);
nor U6001 (N_6001,N_5749,N_5560);
xor U6002 (N_6002,N_5692,N_5685);
or U6003 (N_6003,N_5697,N_5588);
xnor U6004 (N_6004,N_5923,N_5873);
nand U6005 (N_6005,N_5942,N_5769);
nand U6006 (N_6006,N_5841,N_5883);
and U6007 (N_6007,N_5765,N_5583);
nor U6008 (N_6008,N_5845,N_5870);
xnor U6009 (N_6009,N_5605,N_5686);
xor U6010 (N_6010,N_5719,N_5834);
nor U6011 (N_6011,N_5553,N_5791);
nand U6012 (N_6012,N_5664,N_5879);
nor U6013 (N_6013,N_5996,N_5562);
or U6014 (N_6014,N_5801,N_5533);
nor U6015 (N_6015,N_5954,N_5946);
or U6016 (N_6016,N_5542,N_5958);
xor U6017 (N_6017,N_5750,N_5520);
and U6018 (N_6018,N_5717,N_5930);
or U6019 (N_6019,N_5940,N_5854);
or U6020 (N_6020,N_5529,N_5613);
nor U6021 (N_6021,N_5943,N_5890);
and U6022 (N_6022,N_5563,N_5985);
and U6023 (N_6023,N_5671,N_5628);
nand U6024 (N_6024,N_5661,N_5868);
nor U6025 (N_6025,N_5986,N_5784);
and U6026 (N_6026,N_5687,N_5997);
nor U6027 (N_6027,N_5739,N_5939);
nor U6028 (N_6028,N_5781,N_5508);
nor U6029 (N_6029,N_5876,N_5531);
or U6030 (N_6030,N_5540,N_5523);
nor U6031 (N_6031,N_5695,N_5742);
and U6032 (N_6032,N_5838,N_5917);
nor U6033 (N_6033,N_5682,N_5753);
nand U6034 (N_6034,N_5855,N_5975);
nand U6035 (N_6035,N_5904,N_5952);
and U6036 (N_6036,N_5909,N_5751);
nor U6037 (N_6037,N_5595,N_5830);
nor U6038 (N_6038,N_5945,N_5568);
and U6039 (N_6039,N_5893,N_5672);
and U6040 (N_6040,N_5927,N_5994);
xor U6041 (N_6041,N_5561,N_5502);
nand U6042 (N_6042,N_5677,N_5813);
nand U6043 (N_6043,N_5809,N_5575);
and U6044 (N_6044,N_5715,N_5828);
nand U6045 (N_6045,N_5860,N_5853);
nor U6046 (N_6046,N_5983,N_5734);
or U6047 (N_6047,N_5735,N_5903);
and U6048 (N_6048,N_5888,N_5780);
nor U6049 (N_6049,N_5732,N_5698);
and U6050 (N_6050,N_5691,N_5637);
nor U6051 (N_6051,N_5777,N_5878);
xor U6052 (N_6052,N_5977,N_5793);
or U6053 (N_6053,N_5815,N_5938);
xor U6054 (N_6054,N_5999,N_5709);
nor U6055 (N_6055,N_5567,N_5901);
and U6056 (N_6056,N_5933,N_5899);
and U6057 (N_6057,N_5914,N_5882);
and U6058 (N_6058,N_5675,N_5960);
xor U6059 (N_6059,N_5645,N_5846);
or U6060 (N_6060,N_5835,N_5844);
or U6061 (N_6061,N_5574,N_5707);
nand U6062 (N_6062,N_5822,N_5987);
or U6063 (N_6063,N_5514,N_5956);
and U6064 (N_6064,N_5626,N_5569);
or U6065 (N_6065,N_5968,N_5738);
or U6066 (N_6066,N_5795,N_5849);
and U6067 (N_6067,N_5741,N_5979);
or U6068 (N_6068,N_5915,N_5772);
nand U6069 (N_6069,N_5866,N_5621);
xnor U6070 (N_6070,N_5537,N_5875);
nor U6071 (N_6071,N_5957,N_5897);
nor U6072 (N_6072,N_5526,N_5803);
or U6073 (N_6073,N_5551,N_5612);
xor U6074 (N_6074,N_5948,N_5907);
and U6075 (N_6075,N_5790,N_5874);
nand U6076 (N_6076,N_5651,N_5779);
nor U6077 (N_6077,N_5653,N_5951);
nand U6078 (N_6078,N_5949,N_5743);
nand U6079 (N_6079,N_5723,N_5934);
and U6080 (N_6080,N_5810,N_5762);
nor U6081 (N_6081,N_5729,N_5725);
nor U6082 (N_6082,N_5867,N_5877);
or U6083 (N_6083,N_5926,N_5991);
and U6084 (N_6084,N_5850,N_5688);
nand U6085 (N_6085,N_5722,N_5961);
xor U6086 (N_6086,N_5861,N_5929);
and U6087 (N_6087,N_5674,N_5716);
or U6088 (N_6088,N_5884,N_5837);
xnor U6089 (N_6089,N_5696,N_5895);
nand U6090 (N_6090,N_5840,N_5978);
and U6091 (N_6091,N_5988,N_5922);
or U6092 (N_6092,N_5591,N_5679);
nor U6093 (N_6093,N_5941,N_5746);
nor U6094 (N_6094,N_5599,N_5980);
nor U6095 (N_6095,N_5759,N_5507);
or U6096 (N_6096,N_5851,N_5964);
or U6097 (N_6097,N_5812,N_5789);
nand U6098 (N_6098,N_5639,N_5885);
nor U6099 (N_6099,N_5965,N_5608);
nor U6100 (N_6100,N_5549,N_5908);
xor U6101 (N_6101,N_5976,N_5635);
xnor U6102 (N_6102,N_5763,N_5678);
nor U6103 (N_6103,N_5902,N_5654);
xor U6104 (N_6104,N_5761,N_5842);
xnor U6105 (N_6105,N_5513,N_5871);
and U6106 (N_6106,N_5826,N_5816);
nand U6107 (N_6107,N_5831,N_5768);
or U6108 (N_6108,N_5788,N_5745);
nor U6109 (N_6109,N_5546,N_5623);
nand U6110 (N_6110,N_5571,N_5969);
nand U6111 (N_6111,N_5995,N_5510);
and U6112 (N_6112,N_5604,N_5598);
xnor U6113 (N_6113,N_5858,N_5548);
and U6114 (N_6114,N_5665,N_5913);
and U6115 (N_6115,N_5823,N_5869);
nand U6116 (N_6116,N_5924,N_5953);
and U6117 (N_6117,N_5655,N_5618);
nand U6118 (N_6118,N_5517,N_5754);
xor U6119 (N_6119,N_5606,N_5536);
nand U6120 (N_6120,N_5629,N_5936);
and U6121 (N_6121,N_5572,N_5865);
nor U6122 (N_6122,N_5689,N_5962);
xnor U6123 (N_6123,N_5658,N_5900);
xor U6124 (N_6124,N_5898,N_5556);
nor U6125 (N_6125,N_5555,N_5796);
and U6126 (N_6126,N_5594,N_5839);
or U6127 (N_6127,N_5764,N_5808);
or U6128 (N_6128,N_5974,N_5802);
nor U6129 (N_6129,N_5638,N_5760);
and U6130 (N_6130,N_5864,N_5600);
xor U6131 (N_6131,N_5557,N_5603);
nor U6132 (N_6132,N_5712,N_5984);
xnor U6133 (N_6133,N_5829,N_5950);
or U6134 (N_6134,N_5634,N_5543);
nand U6135 (N_6135,N_5578,N_5511);
or U6136 (N_6136,N_5972,N_5798);
xnor U6137 (N_6137,N_5642,N_5524);
nor U6138 (N_6138,N_5967,N_5630);
nand U6139 (N_6139,N_5805,N_5740);
nor U6140 (N_6140,N_5714,N_5683);
and U6141 (N_6141,N_5584,N_5652);
and U6142 (N_6142,N_5932,N_5710);
nand U6143 (N_6143,N_5947,N_5773);
nand U6144 (N_6144,N_5617,N_5503);
nor U6145 (N_6145,N_5771,N_5538);
nand U6146 (N_6146,N_5545,N_5752);
or U6147 (N_6147,N_5767,N_5582);
xnor U6148 (N_6148,N_5819,N_5919);
nor U6149 (N_6149,N_5570,N_5647);
or U6150 (N_6150,N_5731,N_5559);
nand U6151 (N_6151,N_5643,N_5676);
or U6152 (N_6152,N_5515,N_5766);
or U6153 (N_6153,N_5521,N_5579);
and U6154 (N_6154,N_5534,N_5859);
or U6155 (N_6155,N_5797,N_5663);
and U6156 (N_6156,N_5609,N_5852);
or U6157 (N_6157,N_5818,N_5680);
nand U6158 (N_6158,N_5916,N_5547);
nor U6159 (N_6159,N_5711,N_5586);
xnor U6160 (N_6160,N_5610,N_5641);
or U6161 (N_6161,N_5705,N_5959);
or U6162 (N_6162,N_5516,N_5648);
nor U6163 (N_6163,N_5783,N_5587);
nor U6164 (N_6164,N_5565,N_5963);
or U6165 (N_6165,N_5800,N_5554);
and U6166 (N_6166,N_5758,N_5992);
nand U6167 (N_6167,N_5504,N_5911);
or U6168 (N_6168,N_5921,N_5786);
or U6169 (N_6169,N_5889,N_5670);
or U6170 (N_6170,N_5636,N_5891);
or U6171 (N_6171,N_5971,N_5727);
nor U6172 (N_6172,N_5614,N_5702);
and U6173 (N_6173,N_5656,N_5501);
nand U6174 (N_6174,N_5814,N_5694);
xor U6175 (N_6175,N_5527,N_5804);
or U6176 (N_6176,N_5590,N_5640);
and U6177 (N_6177,N_5775,N_5906);
or U6178 (N_6178,N_5863,N_5681);
or U6179 (N_6179,N_5693,N_5667);
nor U6180 (N_6180,N_5799,N_5708);
xnor U6181 (N_6181,N_5820,N_5886);
nor U6182 (N_6182,N_5937,N_5794);
or U6183 (N_6183,N_5669,N_5506);
xor U6184 (N_6184,N_5589,N_5509);
nand U6185 (N_6185,N_5755,N_5539);
nand U6186 (N_6186,N_5862,N_5519);
nand U6187 (N_6187,N_5581,N_5981);
xor U6188 (N_6188,N_5592,N_5528);
or U6189 (N_6189,N_5955,N_5721);
and U6190 (N_6190,N_5807,N_5833);
and U6191 (N_6191,N_5832,N_5880);
nor U6192 (N_6192,N_5646,N_5601);
xnor U6193 (N_6193,N_5892,N_5505);
xnor U6194 (N_6194,N_5673,N_5649);
or U6195 (N_6195,N_5726,N_5660);
and U6196 (N_6196,N_5966,N_5724);
nor U6197 (N_6197,N_5690,N_5792);
nor U6198 (N_6198,N_5744,N_5700);
or U6199 (N_6199,N_5532,N_5713);
and U6200 (N_6200,N_5620,N_5843);
or U6201 (N_6201,N_5585,N_5701);
or U6202 (N_6202,N_5747,N_5544);
xor U6203 (N_6203,N_5552,N_5736);
or U6204 (N_6204,N_5728,N_5905);
nor U6205 (N_6205,N_5644,N_5699);
nand U6206 (N_6206,N_5668,N_5836);
and U6207 (N_6207,N_5944,N_5632);
nor U6208 (N_6208,N_5935,N_5848);
and U6209 (N_6209,N_5970,N_5770);
xnor U6210 (N_6210,N_5593,N_5558);
nand U6211 (N_6211,N_5518,N_5530);
and U6212 (N_6212,N_5856,N_5666);
nand U6213 (N_6213,N_5512,N_5931);
xnor U6214 (N_6214,N_5522,N_5912);
nor U6215 (N_6215,N_5990,N_5622);
nor U6216 (N_6216,N_5631,N_5778);
xnor U6217 (N_6217,N_5684,N_5918);
and U6218 (N_6218,N_5550,N_5576);
and U6219 (N_6219,N_5847,N_5928);
or U6220 (N_6220,N_5896,N_5782);
or U6221 (N_6221,N_5580,N_5627);
and U6222 (N_6222,N_5611,N_5541);
and U6223 (N_6223,N_5624,N_5887);
nor U6224 (N_6224,N_5730,N_5650);
xnor U6225 (N_6225,N_5825,N_5733);
or U6226 (N_6226,N_5748,N_5776);
nand U6227 (N_6227,N_5857,N_5787);
and U6228 (N_6228,N_5615,N_5872);
nor U6229 (N_6229,N_5989,N_5982);
xor U6230 (N_6230,N_5564,N_5774);
and U6231 (N_6231,N_5577,N_5607);
xnor U6232 (N_6232,N_5616,N_5662);
and U6233 (N_6233,N_5881,N_5703);
and U6234 (N_6234,N_5824,N_5566);
nand U6235 (N_6235,N_5973,N_5737);
and U6236 (N_6236,N_5993,N_5910);
nand U6237 (N_6237,N_5785,N_5619);
and U6238 (N_6238,N_5625,N_5757);
nand U6239 (N_6239,N_5704,N_5657);
xor U6240 (N_6240,N_5573,N_5535);
nor U6241 (N_6241,N_5894,N_5806);
nor U6242 (N_6242,N_5602,N_5925);
nor U6243 (N_6243,N_5821,N_5817);
nand U6244 (N_6244,N_5659,N_5827);
and U6245 (N_6245,N_5525,N_5920);
nand U6246 (N_6246,N_5596,N_5756);
nand U6247 (N_6247,N_5633,N_5706);
xnor U6248 (N_6248,N_5718,N_5597);
or U6249 (N_6249,N_5500,N_5720);
xor U6250 (N_6250,N_5593,N_5682);
and U6251 (N_6251,N_5722,N_5851);
nor U6252 (N_6252,N_5776,N_5815);
xor U6253 (N_6253,N_5743,N_5692);
or U6254 (N_6254,N_5528,N_5506);
and U6255 (N_6255,N_5949,N_5538);
nand U6256 (N_6256,N_5755,N_5530);
nor U6257 (N_6257,N_5572,N_5883);
xor U6258 (N_6258,N_5548,N_5805);
nand U6259 (N_6259,N_5743,N_5970);
nor U6260 (N_6260,N_5780,N_5753);
nor U6261 (N_6261,N_5882,N_5808);
nand U6262 (N_6262,N_5818,N_5995);
or U6263 (N_6263,N_5623,N_5957);
xor U6264 (N_6264,N_5817,N_5546);
nand U6265 (N_6265,N_5702,N_5678);
and U6266 (N_6266,N_5891,N_5601);
xor U6267 (N_6267,N_5781,N_5676);
nand U6268 (N_6268,N_5619,N_5924);
nand U6269 (N_6269,N_5673,N_5913);
and U6270 (N_6270,N_5502,N_5846);
nand U6271 (N_6271,N_5524,N_5820);
and U6272 (N_6272,N_5935,N_5594);
nand U6273 (N_6273,N_5967,N_5831);
nor U6274 (N_6274,N_5941,N_5704);
nand U6275 (N_6275,N_5640,N_5574);
xor U6276 (N_6276,N_5924,N_5600);
or U6277 (N_6277,N_5802,N_5925);
nand U6278 (N_6278,N_5535,N_5942);
nand U6279 (N_6279,N_5919,N_5832);
and U6280 (N_6280,N_5653,N_5558);
nand U6281 (N_6281,N_5896,N_5552);
nand U6282 (N_6282,N_5503,N_5841);
and U6283 (N_6283,N_5622,N_5570);
and U6284 (N_6284,N_5841,N_5662);
xnor U6285 (N_6285,N_5710,N_5567);
nand U6286 (N_6286,N_5723,N_5733);
xor U6287 (N_6287,N_5593,N_5521);
nor U6288 (N_6288,N_5627,N_5625);
or U6289 (N_6289,N_5809,N_5707);
nand U6290 (N_6290,N_5831,N_5747);
or U6291 (N_6291,N_5634,N_5830);
xor U6292 (N_6292,N_5790,N_5823);
nor U6293 (N_6293,N_5705,N_5622);
or U6294 (N_6294,N_5536,N_5840);
or U6295 (N_6295,N_5882,N_5818);
nor U6296 (N_6296,N_5990,N_5709);
and U6297 (N_6297,N_5613,N_5663);
or U6298 (N_6298,N_5531,N_5613);
xnor U6299 (N_6299,N_5962,N_5746);
nor U6300 (N_6300,N_5884,N_5653);
nand U6301 (N_6301,N_5944,N_5551);
or U6302 (N_6302,N_5812,N_5559);
nor U6303 (N_6303,N_5812,N_5853);
or U6304 (N_6304,N_5931,N_5804);
and U6305 (N_6305,N_5585,N_5984);
xnor U6306 (N_6306,N_5851,N_5660);
nand U6307 (N_6307,N_5666,N_5681);
nor U6308 (N_6308,N_5676,N_5595);
nand U6309 (N_6309,N_5579,N_5510);
or U6310 (N_6310,N_5811,N_5535);
nor U6311 (N_6311,N_5900,N_5677);
or U6312 (N_6312,N_5631,N_5629);
or U6313 (N_6313,N_5837,N_5688);
nand U6314 (N_6314,N_5566,N_5556);
xor U6315 (N_6315,N_5520,N_5518);
and U6316 (N_6316,N_5810,N_5806);
nand U6317 (N_6317,N_5502,N_5713);
and U6318 (N_6318,N_5579,N_5987);
nor U6319 (N_6319,N_5658,N_5685);
nor U6320 (N_6320,N_5909,N_5676);
xnor U6321 (N_6321,N_5900,N_5576);
nor U6322 (N_6322,N_5753,N_5697);
nor U6323 (N_6323,N_5818,N_5616);
and U6324 (N_6324,N_5700,N_5746);
xnor U6325 (N_6325,N_5711,N_5628);
nor U6326 (N_6326,N_5842,N_5984);
xor U6327 (N_6327,N_5768,N_5725);
or U6328 (N_6328,N_5584,N_5575);
xor U6329 (N_6329,N_5688,N_5920);
xor U6330 (N_6330,N_5717,N_5668);
nor U6331 (N_6331,N_5622,N_5774);
xnor U6332 (N_6332,N_5823,N_5556);
nand U6333 (N_6333,N_5789,N_5815);
nor U6334 (N_6334,N_5956,N_5960);
nand U6335 (N_6335,N_5746,N_5744);
nor U6336 (N_6336,N_5933,N_5897);
xor U6337 (N_6337,N_5740,N_5532);
nand U6338 (N_6338,N_5738,N_5658);
xnor U6339 (N_6339,N_5622,N_5745);
xor U6340 (N_6340,N_5774,N_5848);
or U6341 (N_6341,N_5805,N_5970);
and U6342 (N_6342,N_5942,N_5998);
xnor U6343 (N_6343,N_5826,N_5694);
nand U6344 (N_6344,N_5881,N_5663);
and U6345 (N_6345,N_5726,N_5859);
nor U6346 (N_6346,N_5675,N_5611);
or U6347 (N_6347,N_5644,N_5586);
xnor U6348 (N_6348,N_5944,N_5789);
or U6349 (N_6349,N_5761,N_5988);
nor U6350 (N_6350,N_5806,N_5553);
and U6351 (N_6351,N_5750,N_5509);
nor U6352 (N_6352,N_5966,N_5500);
or U6353 (N_6353,N_5641,N_5696);
nand U6354 (N_6354,N_5673,N_5654);
or U6355 (N_6355,N_5578,N_5546);
and U6356 (N_6356,N_5976,N_5936);
xnor U6357 (N_6357,N_5784,N_5533);
and U6358 (N_6358,N_5880,N_5948);
or U6359 (N_6359,N_5730,N_5758);
or U6360 (N_6360,N_5596,N_5552);
and U6361 (N_6361,N_5615,N_5764);
and U6362 (N_6362,N_5964,N_5763);
nand U6363 (N_6363,N_5881,N_5501);
nor U6364 (N_6364,N_5797,N_5809);
and U6365 (N_6365,N_5727,N_5746);
or U6366 (N_6366,N_5892,N_5993);
and U6367 (N_6367,N_5553,N_5577);
nor U6368 (N_6368,N_5963,N_5718);
and U6369 (N_6369,N_5998,N_5568);
or U6370 (N_6370,N_5815,N_5751);
and U6371 (N_6371,N_5701,N_5915);
or U6372 (N_6372,N_5923,N_5972);
and U6373 (N_6373,N_5867,N_5764);
or U6374 (N_6374,N_5770,N_5738);
nor U6375 (N_6375,N_5688,N_5572);
or U6376 (N_6376,N_5631,N_5945);
and U6377 (N_6377,N_5743,N_5672);
xor U6378 (N_6378,N_5660,N_5593);
xnor U6379 (N_6379,N_5725,N_5801);
and U6380 (N_6380,N_5546,N_5551);
xor U6381 (N_6381,N_5744,N_5635);
xor U6382 (N_6382,N_5539,N_5837);
xnor U6383 (N_6383,N_5894,N_5777);
nor U6384 (N_6384,N_5795,N_5610);
nand U6385 (N_6385,N_5730,N_5548);
xnor U6386 (N_6386,N_5760,N_5687);
or U6387 (N_6387,N_5772,N_5845);
nand U6388 (N_6388,N_5744,N_5511);
nor U6389 (N_6389,N_5918,N_5588);
nor U6390 (N_6390,N_5603,N_5966);
xnor U6391 (N_6391,N_5776,N_5680);
nand U6392 (N_6392,N_5839,N_5845);
nand U6393 (N_6393,N_5659,N_5625);
nand U6394 (N_6394,N_5640,N_5668);
xnor U6395 (N_6395,N_5745,N_5720);
nand U6396 (N_6396,N_5647,N_5502);
or U6397 (N_6397,N_5912,N_5631);
nor U6398 (N_6398,N_5779,N_5816);
nand U6399 (N_6399,N_5653,N_5665);
or U6400 (N_6400,N_5633,N_5789);
nor U6401 (N_6401,N_5997,N_5567);
xor U6402 (N_6402,N_5632,N_5559);
or U6403 (N_6403,N_5986,N_5932);
and U6404 (N_6404,N_5582,N_5664);
or U6405 (N_6405,N_5730,N_5995);
nor U6406 (N_6406,N_5921,N_5749);
nor U6407 (N_6407,N_5699,N_5583);
nor U6408 (N_6408,N_5771,N_5742);
and U6409 (N_6409,N_5882,N_5530);
and U6410 (N_6410,N_5845,N_5967);
nor U6411 (N_6411,N_5998,N_5926);
and U6412 (N_6412,N_5893,N_5913);
xor U6413 (N_6413,N_5674,N_5571);
and U6414 (N_6414,N_5874,N_5966);
or U6415 (N_6415,N_5706,N_5690);
or U6416 (N_6416,N_5625,N_5940);
xnor U6417 (N_6417,N_5599,N_5619);
xnor U6418 (N_6418,N_5512,N_5718);
and U6419 (N_6419,N_5520,N_5607);
nand U6420 (N_6420,N_5696,N_5655);
nand U6421 (N_6421,N_5638,N_5849);
or U6422 (N_6422,N_5785,N_5732);
nor U6423 (N_6423,N_5743,N_5727);
or U6424 (N_6424,N_5881,N_5653);
or U6425 (N_6425,N_5842,N_5832);
and U6426 (N_6426,N_5928,N_5977);
nand U6427 (N_6427,N_5825,N_5628);
nand U6428 (N_6428,N_5512,N_5891);
xor U6429 (N_6429,N_5860,N_5916);
and U6430 (N_6430,N_5756,N_5876);
or U6431 (N_6431,N_5978,N_5930);
nor U6432 (N_6432,N_5755,N_5596);
xor U6433 (N_6433,N_5907,N_5698);
nand U6434 (N_6434,N_5917,N_5770);
or U6435 (N_6435,N_5799,N_5594);
nor U6436 (N_6436,N_5544,N_5695);
nand U6437 (N_6437,N_5603,N_5948);
nand U6438 (N_6438,N_5981,N_5893);
xnor U6439 (N_6439,N_5769,N_5826);
xnor U6440 (N_6440,N_5934,N_5985);
and U6441 (N_6441,N_5544,N_5550);
or U6442 (N_6442,N_5882,N_5665);
and U6443 (N_6443,N_5526,N_5962);
and U6444 (N_6444,N_5724,N_5554);
nand U6445 (N_6445,N_5786,N_5577);
or U6446 (N_6446,N_5884,N_5690);
nor U6447 (N_6447,N_5543,N_5866);
xnor U6448 (N_6448,N_5955,N_5776);
nand U6449 (N_6449,N_5622,N_5850);
and U6450 (N_6450,N_5514,N_5551);
nor U6451 (N_6451,N_5672,N_5826);
and U6452 (N_6452,N_5638,N_5726);
xor U6453 (N_6453,N_5652,N_5525);
and U6454 (N_6454,N_5773,N_5907);
and U6455 (N_6455,N_5687,N_5509);
or U6456 (N_6456,N_5539,N_5898);
nor U6457 (N_6457,N_5938,N_5580);
nor U6458 (N_6458,N_5940,N_5583);
and U6459 (N_6459,N_5986,N_5809);
and U6460 (N_6460,N_5791,N_5847);
and U6461 (N_6461,N_5806,N_5996);
xor U6462 (N_6462,N_5740,N_5560);
xnor U6463 (N_6463,N_5647,N_5821);
xnor U6464 (N_6464,N_5606,N_5732);
and U6465 (N_6465,N_5941,N_5631);
and U6466 (N_6466,N_5741,N_5978);
nand U6467 (N_6467,N_5837,N_5609);
xor U6468 (N_6468,N_5516,N_5933);
nand U6469 (N_6469,N_5552,N_5971);
or U6470 (N_6470,N_5638,N_5733);
or U6471 (N_6471,N_5811,N_5860);
nor U6472 (N_6472,N_5673,N_5667);
xor U6473 (N_6473,N_5517,N_5726);
or U6474 (N_6474,N_5762,N_5872);
xor U6475 (N_6475,N_5899,N_5832);
xnor U6476 (N_6476,N_5526,N_5542);
nor U6477 (N_6477,N_5931,N_5702);
and U6478 (N_6478,N_5765,N_5953);
xor U6479 (N_6479,N_5870,N_5751);
xor U6480 (N_6480,N_5997,N_5536);
nand U6481 (N_6481,N_5672,N_5781);
xnor U6482 (N_6482,N_5582,N_5834);
and U6483 (N_6483,N_5531,N_5943);
and U6484 (N_6484,N_5902,N_5547);
nand U6485 (N_6485,N_5501,N_5602);
or U6486 (N_6486,N_5596,N_5570);
or U6487 (N_6487,N_5544,N_5913);
xor U6488 (N_6488,N_5924,N_5865);
and U6489 (N_6489,N_5916,N_5945);
and U6490 (N_6490,N_5721,N_5861);
xnor U6491 (N_6491,N_5701,N_5952);
nand U6492 (N_6492,N_5916,N_5522);
nand U6493 (N_6493,N_5690,N_5501);
nand U6494 (N_6494,N_5910,N_5564);
xnor U6495 (N_6495,N_5755,N_5809);
nor U6496 (N_6496,N_5910,N_5521);
xor U6497 (N_6497,N_5891,N_5898);
nand U6498 (N_6498,N_5920,N_5511);
xor U6499 (N_6499,N_5684,N_5937);
and U6500 (N_6500,N_6123,N_6434);
nand U6501 (N_6501,N_6212,N_6244);
xnor U6502 (N_6502,N_6311,N_6352);
or U6503 (N_6503,N_6115,N_6442);
nor U6504 (N_6504,N_6356,N_6259);
xor U6505 (N_6505,N_6204,N_6369);
or U6506 (N_6506,N_6074,N_6421);
nor U6507 (N_6507,N_6000,N_6349);
nor U6508 (N_6508,N_6368,N_6217);
nand U6509 (N_6509,N_6483,N_6094);
or U6510 (N_6510,N_6206,N_6319);
nor U6511 (N_6511,N_6315,N_6072);
nand U6512 (N_6512,N_6213,N_6291);
and U6513 (N_6513,N_6031,N_6242);
xnor U6514 (N_6514,N_6454,N_6284);
nand U6515 (N_6515,N_6260,N_6230);
and U6516 (N_6516,N_6026,N_6139);
nand U6517 (N_6517,N_6295,N_6264);
nor U6518 (N_6518,N_6058,N_6188);
nor U6519 (N_6519,N_6306,N_6451);
xnor U6520 (N_6520,N_6262,N_6080);
nand U6521 (N_6521,N_6109,N_6279);
nand U6522 (N_6522,N_6373,N_6446);
nand U6523 (N_6523,N_6441,N_6430);
and U6524 (N_6524,N_6268,N_6256);
and U6525 (N_6525,N_6463,N_6481);
xnor U6526 (N_6526,N_6363,N_6357);
xor U6527 (N_6527,N_6327,N_6414);
nand U6528 (N_6528,N_6347,N_6056);
and U6529 (N_6529,N_6012,N_6416);
nor U6530 (N_6530,N_6226,N_6101);
and U6531 (N_6531,N_6489,N_6289);
xnor U6532 (N_6532,N_6033,N_6257);
nand U6533 (N_6533,N_6147,N_6035);
and U6534 (N_6534,N_6486,N_6392);
nand U6535 (N_6535,N_6041,N_6344);
nor U6536 (N_6536,N_6415,N_6010);
xnor U6537 (N_6537,N_6020,N_6419);
nand U6538 (N_6538,N_6223,N_6241);
xnor U6539 (N_6539,N_6346,N_6365);
or U6540 (N_6540,N_6117,N_6053);
xnor U6541 (N_6541,N_6364,N_6271);
or U6542 (N_6542,N_6336,N_6297);
nor U6543 (N_6543,N_6119,N_6091);
nor U6544 (N_6544,N_6361,N_6413);
xor U6545 (N_6545,N_6073,N_6371);
xnor U6546 (N_6546,N_6084,N_6394);
or U6547 (N_6547,N_6350,N_6285);
and U6548 (N_6548,N_6039,N_6251);
or U6549 (N_6549,N_6301,N_6405);
xnor U6550 (N_6550,N_6077,N_6219);
or U6551 (N_6551,N_6396,N_6062);
and U6552 (N_6552,N_6351,N_6034);
nand U6553 (N_6553,N_6193,N_6155);
xor U6554 (N_6554,N_6330,N_6304);
and U6555 (N_6555,N_6466,N_6167);
nor U6556 (N_6556,N_6423,N_6049);
or U6557 (N_6557,N_6132,N_6177);
xor U6558 (N_6558,N_6360,N_6013);
and U6559 (N_6559,N_6417,N_6032);
nand U6560 (N_6560,N_6469,N_6222);
nor U6561 (N_6561,N_6467,N_6435);
nand U6562 (N_6562,N_6255,N_6144);
and U6563 (N_6563,N_6444,N_6465);
nor U6564 (N_6564,N_6438,N_6207);
or U6565 (N_6565,N_6341,N_6280);
nand U6566 (N_6566,N_6487,N_6014);
nand U6567 (N_6567,N_6339,N_6168);
and U6568 (N_6568,N_6092,N_6048);
nand U6569 (N_6569,N_6275,N_6431);
nor U6570 (N_6570,N_6105,N_6385);
nor U6571 (N_6571,N_6043,N_6282);
nor U6572 (N_6572,N_6015,N_6247);
nor U6573 (N_6573,N_6436,N_6156);
nand U6574 (N_6574,N_6426,N_6252);
nor U6575 (N_6575,N_6003,N_6358);
or U6576 (N_6576,N_6201,N_6078);
or U6577 (N_6577,N_6118,N_6180);
and U6578 (N_6578,N_6069,N_6008);
nor U6579 (N_6579,N_6300,N_6461);
and U6580 (N_6580,N_6353,N_6239);
nor U6581 (N_6581,N_6173,N_6044);
xor U6582 (N_6582,N_6063,N_6302);
nand U6583 (N_6583,N_6445,N_6471);
nor U6584 (N_6584,N_6211,N_6238);
and U6585 (N_6585,N_6340,N_6307);
nand U6586 (N_6586,N_6397,N_6272);
or U6587 (N_6587,N_6197,N_6348);
and U6588 (N_6588,N_6157,N_6440);
nor U6589 (N_6589,N_6175,N_6002);
nor U6590 (N_6590,N_6288,N_6199);
xnor U6591 (N_6591,N_6064,N_6022);
nor U6592 (N_6592,N_6087,N_6472);
nor U6593 (N_6593,N_6061,N_6292);
nor U6594 (N_6594,N_6057,N_6135);
and U6595 (N_6595,N_6408,N_6420);
xnor U6596 (N_6596,N_6402,N_6484);
nor U6597 (N_6597,N_6198,N_6021);
nand U6598 (N_6598,N_6428,N_6146);
and U6599 (N_6599,N_6138,N_6164);
nand U6600 (N_6600,N_6376,N_6065);
nor U6601 (N_6601,N_6407,N_6089);
and U6602 (N_6602,N_6232,N_6097);
nor U6603 (N_6603,N_6354,N_6382);
xnor U6604 (N_6604,N_6298,N_6178);
and U6605 (N_6605,N_6121,N_6322);
and U6606 (N_6606,N_6149,N_6161);
and U6607 (N_6607,N_6190,N_6389);
nor U6608 (N_6608,N_6130,N_6220);
and U6609 (N_6609,N_6203,N_6393);
nor U6610 (N_6610,N_6458,N_6253);
or U6611 (N_6611,N_6399,N_6030);
nor U6612 (N_6612,N_6208,N_6059);
nand U6613 (N_6613,N_6494,N_6313);
nor U6614 (N_6614,N_6099,N_6482);
nor U6615 (N_6615,N_6098,N_6224);
and U6616 (N_6616,N_6437,N_6497);
or U6617 (N_6617,N_6055,N_6200);
or U6618 (N_6618,N_6390,N_6216);
or U6619 (N_6619,N_6294,N_6479);
or U6620 (N_6620,N_6470,N_6498);
or U6621 (N_6621,N_6066,N_6227);
nand U6622 (N_6622,N_6007,N_6102);
nor U6623 (N_6623,N_6269,N_6004);
and U6624 (N_6624,N_6129,N_6281);
xor U6625 (N_6625,N_6001,N_6141);
nand U6626 (N_6626,N_6192,N_6355);
or U6627 (N_6627,N_6383,N_6303);
nand U6628 (N_6628,N_6116,N_6127);
and U6629 (N_6629,N_6455,N_6112);
or U6630 (N_6630,N_6174,N_6179);
or U6631 (N_6631,N_6338,N_6187);
nand U6632 (N_6632,N_6370,N_6495);
nor U6633 (N_6633,N_6140,N_6305);
nor U6634 (N_6634,N_6337,N_6406);
nand U6635 (N_6635,N_6037,N_6328);
nor U6636 (N_6636,N_6148,N_6321);
and U6637 (N_6637,N_6071,N_6362);
and U6638 (N_6638,N_6153,N_6462);
and U6639 (N_6639,N_6237,N_6134);
or U6640 (N_6640,N_6186,N_6299);
xnor U6641 (N_6641,N_6027,N_6453);
or U6642 (N_6642,N_6496,N_6409);
xnor U6643 (N_6643,N_6016,N_6182);
xnor U6644 (N_6644,N_6286,N_6050);
xor U6645 (N_6645,N_6137,N_6277);
and U6646 (N_6646,N_6070,N_6051);
or U6647 (N_6647,N_6296,N_6185);
xor U6648 (N_6648,N_6183,N_6045);
and U6649 (N_6649,N_6249,N_6060);
xor U6650 (N_6650,N_6374,N_6125);
nor U6651 (N_6651,N_6085,N_6452);
nor U6652 (N_6652,N_6499,N_6011);
or U6653 (N_6653,N_6290,N_6492);
or U6654 (N_6654,N_6473,N_6169);
nand U6655 (N_6655,N_6403,N_6378);
and U6656 (N_6656,N_6410,N_6194);
nand U6657 (N_6657,N_6250,N_6439);
and U6658 (N_6658,N_6145,N_6491);
nor U6659 (N_6659,N_6323,N_6468);
and U6660 (N_6660,N_6176,N_6126);
and U6661 (N_6661,N_6418,N_6448);
or U6662 (N_6662,N_6433,N_6443);
or U6663 (N_6663,N_6228,N_6096);
or U6664 (N_6664,N_6159,N_6375);
or U6665 (N_6665,N_6189,N_6345);
or U6666 (N_6666,N_6236,N_6457);
nand U6667 (N_6667,N_6398,N_6326);
nand U6668 (N_6668,N_6229,N_6088);
or U6669 (N_6669,N_6172,N_6122);
nor U6670 (N_6670,N_6450,N_6047);
xnor U6671 (N_6671,N_6265,N_6171);
or U6672 (N_6672,N_6195,N_6107);
or U6673 (N_6673,N_6331,N_6150);
or U6674 (N_6674,N_6267,N_6422);
nor U6675 (N_6675,N_6191,N_6120);
or U6676 (N_6676,N_6093,N_6395);
xor U6677 (N_6677,N_6005,N_6372);
and U6678 (N_6678,N_6432,N_6215);
or U6679 (N_6679,N_6209,N_6196);
nor U6680 (N_6680,N_6309,N_6076);
xor U6681 (N_6681,N_6427,N_6052);
or U6682 (N_6682,N_6310,N_6480);
xnor U6683 (N_6683,N_6424,N_6036);
xnor U6684 (N_6684,N_6391,N_6377);
nor U6685 (N_6685,N_6166,N_6386);
and U6686 (N_6686,N_6324,N_6090);
xnor U6687 (N_6687,N_6388,N_6283);
and U6688 (N_6688,N_6384,N_6475);
and U6689 (N_6689,N_6308,N_6261);
or U6690 (N_6690,N_6317,N_6009);
and U6691 (N_6691,N_6075,N_6083);
or U6692 (N_6692,N_6273,N_6234);
nand U6693 (N_6693,N_6131,N_6320);
nand U6694 (N_6694,N_6154,N_6142);
nor U6695 (N_6695,N_6263,N_6181);
or U6696 (N_6696,N_6367,N_6029);
nand U6697 (N_6697,N_6160,N_6067);
xnor U6698 (N_6698,N_6425,N_6042);
nand U6699 (N_6699,N_6456,N_6411);
xor U6700 (N_6700,N_6028,N_6184);
and U6701 (N_6701,N_6329,N_6113);
xor U6702 (N_6702,N_6017,N_6225);
xor U6703 (N_6703,N_6151,N_6287);
xnor U6704 (N_6704,N_6046,N_6210);
or U6705 (N_6705,N_6248,N_6401);
or U6706 (N_6706,N_6025,N_6006);
nand U6707 (N_6707,N_6240,N_6143);
or U6708 (N_6708,N_6111,N_6478);
or U6709 (N_6709,N_6202,N_6449);
and U6710 (N_6710,N_6079,N_6040);
xnor U6711 (N_6711,N_6379,N_6100);
or U6712 (N_6712,N_6221,N_6086);
or U6713 (N_6713,N_6266,N_6205);
and U6714 (N_6714,N_6231,N_6332);
xnor U6715 (N_6715,N_6019,N_6276);
nor U6716 (N_6716,N_6124,N_6474);
or U6717 (N_6717,N_6108,N_6464);
nand U6718 (N_6718,N_6429,N_6018);
nand U6719 (N_6719,N_6312,N_6162);
and U6720 (N_6720,N_6245,N_6366);
nor U6721 (N_6721,N_6488,N_6325);
nor U6722 (N_6722,N_6485,N_6243);
nand U6723 (N_6723,N_6106,N_6380);
and U6724 (N_6724,N_6476,N_6165);
nand U6725 (N_6725,N_6278,N_6254);
or U6726 (N_6726,N_6214,N_6128);
and U6727 (N_6727,N_6381,N_6246);
or U6728 (N_6728,N_6333,N_6493);
and U6729 (N_6729,N_6318,N_6316);
or U6730 (N_6730,N_6023,N_6460);
nand U6731 (N_6731,N_6095,N_6334);
or U6732 (N_6732,N_6404,N_6274);
xnor U6733 (N_6733,N_6054,N_6387);
xor U6734 (N_6734,N_6082,N_6342);
and U6735 (N_6735,N_6447,N_6314);
and U6736 (N_6736,N_6110,N_6490);
xor U6737 (N_6737,N_6412,N_6293);
or U6738 (N_6738,N_6038,N_6104);
and U6739 (N_6739,N_6170,N_6459);
xnor U6740 (N_6740,N_6068,N_6233);
xnor U6741 (N_6741,N_6343,N_6270);
xnor U6742 (N_6742,N_6136,N_6103);
nor U6743 (N_6743,N_6163,N_6400);
nand U6744 (N_6744,N_6218,N_6158);
nand U6745 (N_6745,N_6258,N_6024);
and U6746 (N_6746,N_6477,N_6235);
nand U6747 (N_6747,N_6335,N_6359);
or U6748 (N_6748,N_6114,N_6152);
and U6749 (N_6749,N_6081,N_6133);
nand U6750 (N_6750,N_6104,N_6471);
nor U6751 (N_6751,N_6067,N_6386);
nand U6752 (N_6752,N_6064,N_6070);
nand U6753 (N_6753,N_6101,N_6307);
nand U6754 (N_6754,N_6254,N_6209);
and U6755 (N_6755,N_6009,N_6438);
nor U6756 (N_6756,N_6251,N_6370);
xor U6757 (N_6757,N_6353,N_6471);
and U6758 (N_6758,N_6186,N_6287);
nor U6759 (N_6759,N_6190,N_6475);
nor U6760 (N_6760,N_6113,N_6145);
and U6761 (N_6761,N_6159,N_6416);
xor U6762 (N_6762,N_6299,N_6425);
and U6763 (N_6763,N_6339,N_6092);
xor U6764 (N_6764,N_6098,N_6100);
or U6765 (N_6765,N_6433,N_6216);
xnor U6766 (N_6766,N_6030,N_6002);
or U6767 (N_6767,N_6295,N_6056);
and U6768 (N_6768,N_6472,N_6440);
nor U6769 (N_6769,N_6161,N_6321);
nor U6770 (N_6770,N_6218,N_6009);
nand U6771 (N_6771,N_6069,N_6402);
and U6772 (N_6772,N_6109,N_6225);
nor U6773 (N_6773,N_6437,N_6084);
xor U6774 (N_6774,N_6402,N_6290);
nor U6775 (N_6775,N_6057,N_6120);
and U6776 (N_6776,N_6333,N_6386);
nand U6777 (N_6777,N_6306,N_6001);
xor U6778 (N_6778,N_6228,N_6145);
nand U6779 (N_6779,N_6061,N_6400);
and U6780 (N_6780,N_6308,N_6325);
or U6781 (N_6781,N_6415,N_6169);
or U6782 (N_6782,N_6198,N_6333);
nand U6783 (N_6783,N_6066,N_6040);
nand U6784 (N_6784,N_6372,N_6291);
xnor U6785 (N_6785,N_6139,N_6366);
or U6786 (N_6786,N_6066,N_6119);
and U6787 (N_6787,N_6140,N_6010);
xor U6788 (N_6788,N_6273,N_6177);
nor U6789 (N_6789,N_6391,N_6337);
or U6790 (N_6790,N_6284,N_6469);
nor U6791 (N_6791,N_6032,N_6433);
nand U6792 (N_6792,N_6473,N_6422);
nand U6793 (N_6793,N_6447,N_6303);
nor U6794 (N_6794,N_6299,N_6184);
nor U6795 (N_6795,N_6470,N_6422);
or U6796 (N_6796,N_6170,N_6130);
nor U6797 (N_6797,N_6358,N_6129);
xnor U6798 (N_6798,N_6283,N_6275);
nor U6799 (N_6799,N_6460,N_6016);
nand U6800 (N_6800,N_6474,N_6016);
or U6801 (N_6801,N_6024,N_6321);
and U6802 (N_6802,N_6290,N_6203);
nor U6803 (N_6803,N_6045,N_6035);
and U6804 (N_6804,N_6473,N_6120);
and U6805 (N_6805,N_6094,N_6157);
or U6806 (N_6806,N_6474,N_6217);
and U6807 (N_6807,N_6260,N_6308);
and U6808 (N_6808,N_6364,N_6335);
or U6809 (N_6809,N_6291,N_6481);
nor U6810 (N_6810,N_6253,N_6191);
or U6811 (N_6811,N_6344,N_6051);
or U6812 (N_6812,N_6453,N_6145);
nand U6813 (N_6813,N_6084,N_6225);
or U6814 (N_6814,N_6360,N_6305);
nor U6815 (N_6815,N_6411,N_6294);
nand U6816 (N_6816,N_6347,N_6260);
nand U6817 (N_6817,N_6106,N_6470);
xor U6818 (N_6818,N_6288,N_6346);
nor U6819 (N_6819,N_6100,N_6269);
nor U6820 (N_6820,N_6121,N_6204);
nand U6821 (N_6821,N_6132,N_6149);
nor U6822 (N_6822,N_6031,N_6119);
and U6823 (N_6823,N_6496,N_6381);
xnor U6824 (N_6824,N_6355,N_6096);
or U6825 (N_6825,N_6139,N_6473);
and U6826 (N_6826,N_6297,N_6161);
or U6827 (N_6827,N_6484,N_6032);
and U6828 (N_6828,N_6080,N_6187);
xnor U6829 (N_6829,N_6181,N_6034);
and U6830 (N_6830,N_6016,N_6293);
xor U6831 (N_6831,N_6445,N_6233);
nor U6832 (N_6832,N_6201,N_6366);
xor U6833 (N_6833,N_6435,N_6167);
nand U6834 (N_6834,N_6002,N_6197);
nor U6835 (N_6835,N_6265,N_6101);
or U6836 (N_6836,N_6344,N_6492);
or U6837 (N_6837,N_6278,N_6332);
and U6838 (N_6838,N_6084,N_6444);
xnor U6839 (N_6839,N_6080,N_6068);
and U6840 (N_6840,N_6386,N_6210);
and U6841 (N_6841,N_6208,N_6183);
or U6842 (N_6842,N_6128,N_6440);
or U6843 (N_6843,N_6252,N_6408);
or U6844 (N_6844,N_6485,N_6174);
nor U6845 (N_6845,N_6014,N_6494);
and U6846 (N_6846,N_6494,N_6383);
or U6847 (N_6847,N_6113,N_6389);
nand U6848 (N_6848,N_6126,N_6222);
nor U6849 (N_6849,N_6349,N_6319);
nor U6850 (N_6850,N_6327,N_6138);
nor U6851 (N_6851,N_6177,N_6465);
and U6852 (N_6852,N_6185,N_6085);
or U6853 (N_6853,N_6022,N_6109);
nor U6854 (N_6854,N_6128,N_6392);
xor U6855 (N_6855,N_6299,N_6043);
and U6856 (N_6856,N_6470,N_6195);
and U6857 (N_6857,N_6214,N_6493);
nor U6858 (N_6858,N_6036,N_6392);
or U6859 (N_6859,N_6063,N_6357);
nand U6860 (N_6860,N_6469,N_6380);
xnor U6861 (N_6861,N_6202,N_6491);
or U6862 (N_6862,N_6032,N_6283);
and U6863 (N_6863,N_6394,N_6169);
and U6864 (N_6864,N_6499,N_6009);
nor U6865 (N_6865,N_6289,N_6221);
or U6866 (N_6866,N_6333,N_6339);
and U6867 (N_6867,N_6496,N_6167);
or U6868 (N_6868,N_6069,N_6427);
nand U6869 (N_6869,N_6029,N_6378);
xor U6870 (N_6870,N_6435,N_6380);
nand U6871 (N_6871,N_6370,N_6331);
nor U6872 (N_6872,N_6387,N_6029);
nor U6873 (N_6873,N_6028,N_6253);
xnor U6874 (N_6874,N_6108,N_6419);
and U6875 (N_6875,N_6183,N_6417);
nand U6876 (N_6876,N_6199,N_6339);
nand U6877 (N_6877,N_6064,N_6265);
nand U6878 (N_6878,N_6173,N_6118);
nand U6879 (N_6879,N_6124,N_6027);
nor U6880 (N_6880,N_6034,N_6472);
nor U6881 (N_6881,N_6462,N_6101);
and U6882 (N_6882,N_6468,N_6381);
xor U6883 (N_6883,N_6007,N_6256);
or U6884 (N_6884,N_6386,N_6379);
and U6885 (N_6885,N_6419,N_6179);
nor U6886 (N_6886,N_6181,N_6375);
nand U6887 (N_6887,N_6260,N_6222);
or U6888 (N_6888,N_6209,N_6477);
and U6889 (N_6889,N_6147,N_6052);
nor U6890 (N_6890,N_6002,N_6137);
or U6891 (N_6891,N_6093,N_6363);
xor U6892 (N_6892,N_6391,N_6242);
or U6893 (N_6893,N_6418,N_6272);
and U6894 (N_6894,N_6022,N_6229);
xnor U6895 (N_6895,N_6430,N_6174);
or U6896 (N_6896,N_6095,N_6176);
or U6897 (N_6897,N_6081,N_6144);
xnor U6898 (N_6898,N_6364,N_6043);
and U6899 (N_6899,N_6409,N_6434);
and U6900 (N_6900,N_6166,N_6382);
or U6901 (N_6901,N_6408,N_6134);
xnor U6902 (N_6902,N_6211,N_6096);
xor U6903 (N_6903,N_6369,N_6081);
xor U6904 (N_6904,N_6474,N_6401);
xnor U6905 (N_6905,N_6097,N_6372);
xnor U6906 (N_6906,N_6464,N_6398);
nand U6907 (N_6907,N_6030,N_6310);
nand U6908 (N_6908,N_6026,N_6104);
or U6909 (N_6909,N_6290,N_6201);
xor U6910 (N_6910,N_6392,N_6148);
and U6911 (N_6911,N_6213,N_6378);
nand U6912 (N_6912,N_6401,N_6089);
nand U6913 (N_6913,N_6438,N_6145);
and U6914 (N_6914,N_6147,N_6038);
or U6915 (N_6915,N_6482,N_6046);
and U6916 (N_6916,N_6436,N_6269);
and U6917 (N_6917,N_6322,N_6249);
or U6918 (N_6918,N_6039,N_6345);
and U6919 (N_6919,N_6052,N_6494);
or U6920 (N_6920,N_6178,N_6352);
xor U6921 (N_6921,N_6413,N_6385);
xor U6922 (N_6922,N_6382,N_6463);
nor U6923 (N_6923,N_6347,N_6213);
xnor U6924 (N_6924,N_6241,N_6054);
xnor U6925 (N_6925,N_6071,N_6162);
xor U6926 (N_6926,N_6162,N_6434);
and U6927 (N_6927,N_6379,N_6027);
nand U6928 (N_6928,N_6353,N_6307);
or U6929 (N_6929,N_6456,N_6085);
nor U6930 (N_6930,N_6085,N_6006);
xnor U6931 (N_6931,N_6133,N_6155);
or U6932 (N_6932,N_6093,N_6140);
and U6933 (N_6933,N_6237,N_6175);
xnor U6934 (N_6934,N_6264,N_6235);
nor U6935 (N_6935,N_6207,N_6209);
and U6936 (N_6936,N_6125,N_6431);
xnor U6937 (N_6937,N_6469,N_6462);
or U6938 (N_6938,N_6443,N_6025);
and U6939 (N_6939,N_6019,N_6309);
nor U6940 (N_6940,N_6060,N_6155);
nand U6941 (N_6941,N_6179,N_6381);
or U6942 (N_6942,N_6278,N_6231);
and U6943 (N_6943,N_6038,N_6351);
and U6944 (N_6944,N_6059,N_6485);
xor U6945 (N_6945,N_6016,N_6019);
xnor U6946 (N_6946,N_6051,N_6079);
and U6947 (N_6947,N_6138,N_6391);
or U6948 (N_6948,N_6290,N_6078);
or U6949 (N_6949,N_6478,N_6324);
and U6950 (N_6950,N_6374,N_6254);
nor U6951 (N_6951,N_6399,N_6173);
or U6952 (N_6952,N_6183,N_6021);
nand U6953 (N_6953,N_6043,N_6144);
nor U6954 (N_6954,N_6453,N_6143);
nor U6955 (N_6955,N_6077,N_6332);
nand U6956 (N_6956,N_6082,N_6333);
nor U6957 (N_6957,N_6426,N_6254);
nand U6958 (N_6958,N_6086,N_6290);
nor U6959 (N_6959,N_6321,N_6037);
xor U6960 (N_6960,N_6097,N_6063);
xnor U6961 (N_6961,N_6167,N_6038);
xor U6962 (N_6962,N_6325,N_6356);
xor U6963 (N_6963,N_6112,N_6285);
and U6964 (N_6964,N_6226,N_6135);
and U6965 (N_6965,N_6150,N_6038);
nand U6966 (N_6966,N_6237,N_6008);
nand U6967 (N_6967,N_6460,N_6243);
nor U6968 (N_6968,N_6396,N_6458);
nand U6969 (N_6969,N_6277,N_6312);
or U6970 (N_6970,N_6010,N_6383);
or U6971 (N_6971,N_6146,N_6071);
and U6972 (N_6972,N_6222,N_6155);
xor U6973 (N_6973,N_6450,N_6486);
nand U6974 (N_6974,N_6376,N_6400);
and U6975 (N_6975,N_6084,N_6451);
xor U6976 (N_6976,N_6230,N_6444);
nand U6977 (N_6977,N_6382,N_6492);
xor U6978 (N_6978,N_6050,N_6382);
nor U6979 (N_6979,N_6031,N_6045);
or U6980 (N_6980,N_6072,N_6006);
or U6981 (N_6981,N_6444,N_6094);
nor U6982 (N_6982,N_6032,N_6399);
xor U6983 (N_6983,N_6339,N_6159);
xor U6984 (N_6984,N_6343,N_6161);
and U6985 (N_6985,N_6260,N_6259);
nor U6986 (N_6986,N_6264,N_6116);
and U6987 (N_6987,N_6306,N_6031);
nand U6988 (N_6988,N_6119,N_6253);
nand U6989 (N_6989,N_6480,N_6072);
or U6990 (N_6990,N_6267,N_6414);
or U6991 (N_6991,N_6309,N_6100);
and U6992 (N_6992,N_6459,N_6430);
or U6993 (N_6993,N_6003,N_6222);
or U6994 (N_6994,N_6156,N_6145);
or U6995 (N_6995,N_6341,N_6340);
nor U6996 (N_6996,N_6261,N_6442);
xor U6997 (N_6997,N_6092,N_6368);
and U6998 (N_6998,N_6392,N_6343);
nor U6999 (N_6999,N_6119,N_6299);
nand U7000 (N_7000,N_6952,N_6930);
nand U7001 (N_7001,N_6631,N_6560);
or U7002 (N_7002,N_6998,N_6554);
nand U7003 (N_7003,N_6935,N_6629);
nor U7004 (N_7004,N_6904,N_6773);
nor U7005 (N_7005,N_6752,N_6525);
xor U7006 (N_7006,N_6580,N_6852);
xnor U7007 (N_7007,N_6527,N_6769);
nand U7008 (N_7008,N_6612,N_6790);
nand U7009 (N_7009,N_6599,N_6634);
xnor U7010 (N_7010,N_6981,N_6531);
xor U7011 (N_7011,N_6977,N_6655);
and U7012 (N_7012,N_6677,N_6537);
nand U7013 (N_7013,N_6965,N_6901);
or U7014 (N_7014,N_6964,N_6893);
nor U7015 (N_7015,N_6805,N_6586);
or U7016 (N_7016,N_6703,N_6548);
nor U7017 (N_7017,N_6807,N_6989);
nand U7018 (N_7018,N_6855,N_6712);
and U7019 (N_7019,N_6513,N_6653);
nand U7020 (N_7020,N_6948,N_6624);
and U7021 (N_7021,N_6719,N_6927);
nor U7022 (N_7022,N_6605,N_6582);
xnor U7023 (N_7023,N_6867,N_6519);
nand U7024 (N_7024,N_6673,N_6972);
xnor U7025 (N_7025,N_6929,N_6583);
xnor U7026 (N_7026,N_6562,N_6918);
nand U7027 (N_7027,N_6664,N_6798);
and U7028 (N_7028,N_6896,N_6541);
and U7029 (N_7029,N_6863,N_6615);
nor U7030 (N_7030,N_6757,N_6718);
or U7031 (N_7031,N_6759,N_6962);
xor U7032 (N_7032,N_6802,N_6746);
or U7033 (N_7033,N_6956,N_6729);
and U7034 (N_7034,N_6838,N_6941);
or U7035 (N_7035,N_6824,N_6632);
nor U7036 (N_7036,N_6990,N_6728);
or U7037 (N_7037,N_6590,N_6611);
nor U7038 (N_7038,N_6791,N_6925);
nor U7039 (N_7039,N_6564,N_6506);
nor U7040 (N_7040,N_6890,N_6887);
xor U7041 (N_7041,N_6570,N_6799);
nand U7042 (N_7042,N_6765,N_6979);
nand U7043 (N_7043,N_6761,N_6899);
nor U7044 (N_7044,N_6808,N_6920);
nor U7045 (N_7045,N_6986,N_6942);
nand U7046 (N_7046,N_6676,N_6767);
nor U7047 (N_7047,N_6571,N_6687);
or U7048 (N_7048,N_6958,N_6575);
xor U7049 (N_7049,N_6841,N_6716);
and U7050 (N_7050,N_6870,N_6818);
nor U7051 (N_7051,N_6847,N_6715);
xor U7052 (N_7052,N_6937,N_6819);
xor U7053 (N_7053,N_6754,N_6500);
xnor U7054 (N_7054,N_6504,N_6600);
nor U7055 (N_7055,N_6789,N_6666);
and U7056 (N_7056,N_6526,N_6874);
and U7057 (N_7057,N_6686,N_6860);
nor U7058 (N_7058,N_6820,N_6917);
nor U7059 (N_7059,N_6878,N_6762);
xnor U7060 (N_7060,N_6505,N_6821);
or U7061 (N_7061,N_6591,N_6569);
or U7062 (N_7062,N_6559,N_6542);
nand U7063 (N_7063,N_6503,N_6518);
xnor U7064 (N_7064,N_6511,N_6785);
nand U7065 (N_7065,N_6540,N_6833);
nand U7066 (N_7066,N_6816,N_6700);
nand U7067 (N_7067,N_6630,N_6800);
and U7068 (N_7068,N_6581,N_6510);
or U7069 (N_7069,N_6671,N_6501);
or U7070 (N_7070,N_6961,N_6781);
or U7071 (N_7071,N_6638,N_6806);
xor U7072 (N_7072,N_6657,N_6649);
and U7073 (N_7073,N_6845,N_6916);
or U7074 (N_7074,N_6936,N_6668);
nor U7075 (N_7075,N_6868,N_6699);
xor U7076 (N_7076,N_6978,N_6683);
nand U7077 (N_7077,N_6794,N_6603);
nor U7078 (N_7078,N_6714,N_6726);
nor U7079 (N_7079,N_6755,N_6980);
or U7080 (N_7080,N_6859,N_6596);
or U7081 (N_7081,N_6745,N_6897);
or U7082 (N_7082,N_6589,N_6646);
nor U7083 (N_7083,N_6932,N_6803);
xor U7084 (N_7084,N_6843,N_6853);
and U7085 (N_7085,N_6610,N_6934);
and U7086 (N_7086,N_6604,N_6751);
and U7087 (N_7087,N_6840,N_6680);
and U7088 (N_7088,N_6926,N_6656);
nand U7089 (N_7089,N_6543,N_6740);
nor U7090 (N_7090,N_6988,N_6865);
xnor U7091 (N_7091,N_6984,N_6871);
or U7092 (N_7092,N_6593,N_6606);
xor U7093 (N_7093,N_6577,N_6619);
xnor U7094 (N_7094,N_6822,N_6607);
nor U7095 (N_7095,N_6970,N_6732);
nor U7096 (N_7096,N_6563,N_6635);
nand U7097 (N_7097,N_6758,N_6633);
xnor U7098 (N_7098,N_6578,N_6681);
nand U7099 (N_7099,N_6766,N_6849);
and U7100 (N_7100,N_6922,N_6848);
xor U7101 (N_7101,N_6975,N_6689);
nor U7102 (N_7102,N_6795,N_6949);
nor U7103 (N_7103,N_6967,N_6709);
or U7104 (N_7104,N_6879,N_6538);
xor U7105 (N_7105,N_6969,N_6720);
xor U7106 (N_7106,N_6731,N_6695);
nand U7107 (N_7107,N_6875,N_6627);
or U7108 (N_7108,N_6924,N_6973);
nor U7109 (N_7109,N_6517,N_6647);
or U7110 (N_7110,N_6869,N_6594);
xnor U7111 (N_7111,N_6959,N_6639);
nand U7112 (N_7112,N_6992,N_6793);
or U7113 (N_7113,N_6888,N_6707);
nand U7114 (N_7114,N_6530,N_6669);
or U7115 (N_7115,N_6684,N_6748);
or U7116 (N_7116,N_6960,N_6620);
and U7117 (N_7117,N_6921,N_6609);
xnor U7118 (N_7118,N_6643,N_6774);
xor U7119 (N_7119,N_6545,N_6994);
or U7120 (N_7120,N_6648,N_6784);
or U7121 (N_7121,N_6588,N_6705);
and U7122 (N_7122,N_6938,N_6725);
or U7123 (N_7123,N_6617,N_6546);
nor U7124 (N_7124,N_6654,N_6674);
nor U7125 (N_7125,N_6626,N_6650);
and U7126 (N_7126,N_6739,N_6997);
nand U7127 (N_7127,N_6864,N_6601);
or U7128 (N_7128,N_6995,N_6642);
or U7129 (N_7129,N_6966,N_6736);
xnor U7130 (N_7130,N_6968,N_6551);
and U7131 (N_7131,N_6895,N_6856);
and U7132 (N_7132,N_6738,N_6829);
nand U7133 (N_7133,N_6682,N_6618);
nand U7134 (N_7134,N_6651,N_6987);
xnor U7135 (N_7135,N_6713,N_6509);
or U7136 (N_7136,N_6903,N_6636);
xnor U7137 (N_7137,N_6830,N_6982);
or U7138 (N_7138,N_6993,N_6614);
nor U7139 (N_7139,N_6827,N_6733);
nand U7140 (N_7140,N_6837,N_6985);
nand U7141 (N_7141,N_6876,N_6944);
xnor U7142 (N_7142,N_6999,N_6771);
nor U7143 (N_7143,N_6913,N_6850);
nand U7144 (N_7144,N_6931,N_6557);
xor U7145 (N_7145,N_6940,N_6826);
xnor U7146 (N_7146,N_6780,N_6892);
or U7147 (N_7147,N_6957,N_6953);
and U7148 (N_7148,N_6585,N_6690);
nand U7149 (N_7149,N_6549,N_6533);
nor U7150 (N_7150,N_6991,N_6539);
and U7151 (N_7151,N_6882,N_6708);
nor U7152 (N_7152,N_6516,N_6685);
and U7153 (N_7153,N_6675,N_6839);
or U7154 (N_7154,N_6658,N_6584);
nand U7155 (N_7155,N_6529,N_6881);
xor U7156 (N_7156,N_6645,N_6954);
nor U7157 (N_7157,N_6670,N_6678);
xnor U7158 (N_7158,N_6796,N_6747);
and U7159 (N_7159,N_6943,N_6717);
nor U7160 (N_7160,N_6662,N_6950);
xnor U7161 (N_7161,N_6813,N_6788);
xnor U7162 (N_7162,N_6534,N_6622);
xnor U7163 (N_7163,N_6891,N_6861);
or U7164 (N_7164,N_6694,N_6907);
nand U7165 (N_7165,N_6923,N_6933);
nand U7166 (N_7166,N_6663,N_6565);
nand U7167 (N_7167,N_6749,N_6592);
or U7168 (N_7168,N_6919,N_6721);
xor U7169 (N_7169,N_6688,N_6814);
xnor U7170 (N_7170,N_6854,N_6776);
xnor U7171 (N_7171,N_6660,N_6884);
nor U7172 (N_7172,N_6621,N_6797);
or U7173 (N_7173,N_6723,N_6889);
nand U7174 (N_7174,N_6886,N_6768);
xnor U7175 (N_7175,N_6782,N_6727);
nand U7176 (N_7176,N_6520,N_6801);
nor U7177 (N_7177,N_6652,N_6885);
xor U7178 (N_7178,N_6811,N_6900);
nand U7179 (N_7179,N_6698,N_6628);
nand U7180 (N_7180,N_6883,N_6706);
xnor U7181 (N_7181,N_6587,N_6905);
nor U7182 (N_7182,N_6844,N_6775);
nand U7183 (N_7183,N_6521,N_6702);
xnor U7184 (N_7184,N_6877,N_6579);
nor U7185 (N_7185,N_6659,N_6831);
xnor U7186 (N_7186,N_6786,N_6544);
or U7187 (N_7187,N_6693,N_6558);
and U7188 (N_7188,N_6711,N_6710);
xor U7189 (N_7189,N_6597,N_6976);
nor U7190 (N_7190,N_6704,N_6692);
and U7191 (N_7191,N_6846,N_6679);
and U7192 (N_7192,N_6835,N_6939);
and U7193 (N_7193,N_6770,N_6898);
and U7194 (N_7194,N_6779,N_6906);
and U7195 (N_7195,N_6522,N_6825);
and U7196 (N_7196,N_6914,N_6823);
and U7197 (N_7197,N_6756,N_6532);
nand U7198 (N_7198,N_6697,N_6777);
nor U7199 (N_7199,N_6894,N_6857);
and U7200 (N_7200,N_6595,N_6743);
xnor U7201 (N_7201,N_6911,N_6613);
xnor U7202 (N_7202,N_6963,N_6828);
and U7203 (N_7203,N_6744,N_6556);
nor U7204 (N_7204,N_6667,N_6946);
xnor U7205 (N_7205,N_6763,N_6815);
nand U7206 (N_7206,N_6760,N_6514);
or U7207 (N_7207,N_6836,N_6661);
nand U7208 (N_7208,N_6608,N_6536);
and U7209 (N_7209,N_6572,N_6974);
nor U7210 (N_7210,N_6507,N_6996);
xnor U7211 (N_7211,N_6555,N_6741);
xnor U7212 (N_7212,N_6858,N_6512);
or U7213 (N_7213,N_6672,N_6722);
nor U7214 (N_7214,N_6644,N_6523);
and U7215 (N_7215,N_6598,N_6730);
xor U7216 (N_7216,N_6909,N_6502);
and U7217 (N_7217,N_6724,N_6851);
nand U7218 (N_7218,N_6568,N_6912);
and U7219 (N_7219,N_6576,N_6842);
or U7220 (N_7220,N_6625,N_6778);
and U7221 (N_7221,N_6641,N_6866);
xor U7222 (N_7222,N_6508,N_6772);
nor U7223 (N_7223,N_6908,N_6880);
nor U7224 (N_7224,N_6553,N_6561);
xnor U7225 (N_7225,N_6832,N_6812);
xnor U7226 (N_7226,N_6550,N_6947);
nand U7227 (N_7227,N_6623,N_6810);
and U7228 (N_7228,N_6691,N_6616);
xor U7229 (N_7229,N_6817,N_6524);
or U7230 (N_7230,N_6750,N_6872);
or U7231 (N_7231,N_6734,N_6804);
xnor U7232 (N_7232,N_6696,N_6971);
nand U7233 (N_7233,N_6701,N_6910);
and U7234 (N_7234,N_6515,N_6951);
nand U7235 (N_7235,N_6945,N_6637);
xor U7236 (N_7236,N_6566,N_6535);
or U7237 (N_7237,N_6567,N_6640);
xor U7238 (N_7238,N_6862,N_6955);
and U7239 (N_7239,N_6928,N_6787);
or U7240 (N_7240,N_6742,N_6764);
xnor U7241 (N_7241,N_6902,N_6573);
nor U7242 (N_7242,N_6737,N_6574);
or U7243 (N_7243,N_6547,N_6834);
or U7244 (N_7244,N_6915,N_6792);
nand U7245 (N_7245,N_6873,N_6602);
or U7246 (N_7246,N_6735,N_6753);
and U7247 (N_7247,N_6528,N_6783);
xor U7248 (N_7248,N_6665,N_6809);
or U7249 (N_7249,N_6983,N_6552);
nor U7250 (N_7250,N_6749,N_6882);
nor U7251 (N_7251,N_6695,N_6953);
and U7252 (N_7252,N_6651,N_6851);
nor U7253 (N_7253,N_6883,N_6764);
or U7254 (N_7254,N_6735,N_6905);
nor U7255 (N_7255,N_6724,N_6715);
nand U7256 (N_7256,N_6763,N_6539);
nand U7257 (N_7257,N_6580,N_6700);
and U7258 (N_7258,N_6798,N_6606);
or U7259 (N_7259,N_6792,N_6903);
nand U7260 (N_7260,N_6594,N_6732);
nand U7261 (N_7261,N_6909,N_6545);
nor U7262 (N_7262,N_6900,N_6946);
and U7263 (N_7263,N_6807,N_6818);
or U7264 (N_7264,N_6846,N_6749);
and U7265 (N_7265,N_6551,N_6965);
xnor U7266 (N_7266,N_6511,N_6741);
xnor U7267 (N_7267,N_6917,N_6606);
and U7268 (N_7268,N_6683,N_6773);
nand U7269 (N_7269,N_6802,N_6782);
and U7270 (N_7270,N_6897,N_6860);
nand U7271 (N_7271,N_6925,N_6553);
xnor U7272 (N_7272,N_6672,N_6800);
xnor U7273 (N_7273,N_6795,N_6956);
or U7274 (N_7274,N_6777,N_6585);
and U7275 (N_7275,N_6823,N_6526);
and U7276 (N_7276,N_6893,N_6799);
nor U7277 (N_7277,N_6689,N_6788);
nor U7278 (N_7278,N_6845,N_6958);
and U7279 (N_7279,N_6643,N_6509);
xnor U7280 (N_7280,N_6645,N_6893);
nand U7281 (N_7281,N_6504,N_6596);
xnor U7282 (N_7282,N_6537,N_6849);
nand U7283 (N_7283,N_6511,N_6915);
xor U7284 (N_7284,N_6508,N_6696);
or U7285 (N_7285,N_6931,N_6789);
nor U7286 (N_7286,N_6521,N_6637);
nor U7287 (N_7287,N_6768,N_6625);
xor U7288 (N_7288,N_6816,N_6883);
nor U7289 (N_7289,N_6679,N_6905);
nor U7290 (N_7290,N_6996,N_6898);
nand U7291 (N_7291,N_6659,N_6632);
and U7292 (N_7292,N_6971,N_6616);
nand U7293 (N_7293,N_6853,N_6580);
and U7294 (N_7294,N_6945,N_6792);
or U7295 (N_7295,N_6919,N_6928);
and U7296 (N_7296,N_6903,N_6523);
and U7297 (N_7297,N_6993,N_6508);
or U7298 (N_7298,N_6860,N_6523);
nor U7299 (N_7299,N_6524,N_6672);
nor U7300 (N_7300,N_6520,N_6738);
xor U7301 (N_7301,N_6707,N_6857);
xnor U7302 (N_7302,N_6669,N_6646);
nand U7303 (N_7303,N_6647,N_6573);
xnor U7304 (N_7304,N_6616,N_6524);
and U7305 (N_7305,N_6777,N_6832);
or U7306 (N_7306,N_6593,N_6650);
xor U7307 (N_7307,N_6557,N_6575);
xor U7308 (N_7308,N_6585,N_6947);
nor U7309 (N_7309,N_6717,N_6606);
nor U7310 (N_7310,N_6516,N_6607);
nor U7311 (N_7311,N_6895,N_6530);
or U7312 (N_7312,N_6969,N_6608);
nand U7313 (N_7313,N_6636,N_6500);
and U7314 (N_7314,N_6926,N_6947);
nand U7315 (N_7315,N_6602,N_6515);
and U7316 (N_7316,N_6613,N_6942);
nor U7317 (N_7317,N_6524,N_6731);
nor U7318 (N_7318,N_6522,N_6544);
or U7319 (N_7319,N_6887,N_6605);
nor U7320 (N_7320,N_6581,N_6727);
or U7321 (N_7321,N_6819,N_6787);
and U7322 (N_7322,N_6609,N_6689);
nor U7323 (N_7323,N_6733,N_6989);
and U7324 (N_7324,N_6890,N_6681);
or U7325 (N_7325,N_6920,N_6568);
and U7326 (N_7326,N_6528,N_6948);
nor U7327 (N_7327,N_6852,N_6715);
or U7328 (N_7328,N_6634,N_6515);
nand U7329 (N_7329,N_6658,N_6963);
nand U7330 (N_7330,N_6831,N_6844);
or U7331 (N_7331,N_6904,N_6656);
nor U7332 (N_7332,N_6677,N_6526);
nor U7333 (N_7333,N_6862,N_6888);
and U7334 (N_7334,N_6986,N_6811);
xnor U7335 (N_7335,N_6977,N_6551);
xor U7336 (N_7336,N_6904,N_6613);
or U7337 (N_7337,N_6771,N_6714);
or U7338 (N_7338,N_6780,N_6636);
or U7339 (N_7339,N_6850,N_6997);
and U7340 (N_7340,N_6712,N_6678);
or U7341 (N_7341,N_6771,N_6602);
nor U7342 (N_7342,N_6687,N_6976);
xnor U7343 (N_7343,N_6687,N_6589);
or U7344 (N_7344,N_6665,N_6517);
or U7345 (N_7345,N_6729,N_6864);
nor U7346 (N_7346,N_6940,N_6943);
nand U7347 (N_7347,N_6902,N_6838);
xor U7348 (N_7348,N_6515,N_6566);
nand U7349 (N_7349,N_6694,N_6695);
nand U7350 (N_7350,N_6942,N_6946);
xor U7351 (N_7351,N_6716,N_6746);
and U7352 (N_7352,N_6634,N_6729);
or U7353 (N_7353,N_6758,N_6771);
nor U7354 (N_7354,N_6752,N_6722);
or U7355 (N_7355,N_6749,N_6655);
xnor U7356 (N_7356,N_6827,N_6815);
xnor U7357 (N_7357,N_6988,N_6673);
or U7358 (N_7358,N_6874,N_6994);
or U7359 (N_7359,N_6767,N_6750);
or U7360 (N_7360,N_6983,N_6949);
xnor U7361 (N_7361,N_6679,N_6945);
nor U7362 (N_7362,N_6753,N_6923);
and U7363 (N_7363,N_6562,N_6884);
nor U7364 (N_7364,N_6580,N_6574);
or U7365 (N_7365,N_6901,N_6973);
nand U7366 (N_7366,N_6882,N_6542);
and U7367 (N_7367,N_6537,N_6720);
nor U7368 (N_7368,N_6759,N_6787);
xor U7369 (N_7369,N_6564,N_6847);
and U7370 (N_7370,N_6738,N_6753);
or U7371 (N_7371,N_6694,N_6790);
and U7372 (N_7372,N_6557,N_6709);
nor U7373 (N_7373,N_6941,N_6674);
xor U7374 (N_7374,N_6847,N_6798);
or U7375 (N_7375,N_6593,N_6550);
nor U7376 (N_7376,N_6683,N_6765);
xnor U7377 (N_7377,N_6980,N_6600);
nand U7378 (N_7378,N_6830,N_6651);
nor U7379 (N_7379,N_6617,N_6938);
or U7380 (N_7380,N_6847,N_6874);
and U7381 (N_7381,N_6757,N_6652);
and U7382 (N_7382,N_6915,N_6686);
and U7383 (N_7383,N_6751,N_6657);
nor U7384 (N_7384,N_6626,N_6911);
nand U7385 (N_7385,N_6535,N_6639);
and U7386 (N_7386,N_6611,N_6885);
or U7387 (N_7387,N_6999,N_6658);
xnor U7388 (N_7388,N_6511,N_6708);
xor U7389 (N_7389,N_6954,N_6939);
and U7390 (N_7390,N_6969,N_6956);
and U7391 (N_7391,N_6555,N_6561);
and U7392 (N_7392,N_6846,N_6742);
nand U7393 (N_7393,N_6914,N_6614);
and U7394 (N_7394,N_6556,N_6929);
nand U7395 (N_7395,N_6981,N_6856);
nor U7396 (N_7396,N_6736,N_6679);
and U7397 (N_7397,N_6635,N_6790);
nand U7398 (N_7398,N_6508,N_6932);
xor U7399 (N_7399,N_6849,N_6818);
xnor U7400 (N_7400,N_6666,N_6596);
nand U7401 (N_7401,N_6943,N_6953);
xnor U7402 (N_7402,N_6656,N_6898);
nor U7403 (N_7403,N_6623,N_6905);
or U7404 (N_7404,N_6578,N_6660);
nand U7405 (N_7405,N_6693,N_6501);
and U7406 (N_7406,N_6616,N_6966);
xor U7407 (N_7407,N_6737,N_6578);
nor U7408 (N_7408,N_6937,N_6700);
or U7409 (N_7409,N_6562,N_6635);
xor U7410 (N_7410,N_6858,N_6564);
or U7411 (N_7411,N_6910,N_6882);
nor U7412 (N_7412,N_6897,N_6702);
or U7413 (N_7413,N_6712,N_6594);
nand U7414 (N_7414,N_6662,N_6835);
nand U7415 (N_7415,N_6940,N_6762);
nor U7416 (N_7416,N_6842,N_6690);
nand U7417 (N_7417,N_6849,N_6905);
or U7418 (N_7418,N_6533,N_6882);
nand U7419 (N_7419,N_6984,N_6867);
nor U7420 (N_7420,N_6597,N_6640);
nor U7421 (N_7421,N_6667,N_6874);
or U7422 (N_7422,N_6797,N_6722);
nor U7423 (N_7423,N_6905,N_6509);
nand U7424 (N_7424,N_6738,N_6640);
or U7425 (N_7425,N_6828,N_6534);
or U7426 (N_7426,N_6762,N_6648);
or U7427 (N_7427,N_6511,N_6789);
and U7428 (N_7428,N_6688,N_6697);
or U7429 (N_7429,N_6565,N_6584);
nand U7430 (N_7430,N_6930,N_6743);
and U7431 (N_7431,N_6534,N_6506);
nor U7432 (N_7432,N_6898,N_6686);
or U7433 (N_7433,N_6722,N_6603);
nand U7434 (N_7434,N_6835,N_6981);
xnor U7435 (N_7435,N_6656,N_6726);
or U7436 (N_7436,N_6702,N_6719);
and U7437 (N_7437,N_6624,N_6620);
or U7438 (N_7438,N_6594,N_6867);
xnor U7439 (N_7439,N_6578,N_6663);
nand U7440 (N_7440,N_6516,N_6927);
and U7441 (N_7441,N_6534,N_6926);
nand U7442 (N_7442,N_6919,N_6952);
xnor U7443 (N_7443,N_6562,N_6529);
xor U7444 (N_7444,N_6887,N_6875);
or U7445 (N_7445,N_6796,N_6963);
and U7446 (N_7446,N_6562,N_6509);
xor U7447 (N_7447,N_6558,N_6585);
nand U7448 (N_7448,N_6535,N_6669);
nand U7449 (N_7449,N_6553,N_6784);
xor U7450 (N_7450,N_6946,N_6860);
nor U7451 (N_7451,N_6989,N_6683);
or U7452 (N_7452,N_6698,N_6635);
and U7453 (N_7453,N_6865,N_6744);
and U7454 (N_7454,N_6834,N_6993);
nand U7455 (N_7455,N_6685,N_6805);
and U7456 (N_7456,N_6506,N_6772);
nand U7457 (N_7457,N_6634,N_6872);
and U7458 (N_7458,N_6715,N_6865);
and U7459 (N_7459,N_6532,N_6815);
nand U7460 (N_7460,N_6578,N_6983);
or U7461 (N_7461,N_6759,N_6529);
nand U7462 (N_7462,N_6893,N_6566);
and U7463 (N_7463,N_6993,N_6820);
nor U7464 (N_7464,N_6844,N_6922);
and U7465 (N_7465,N_6821,N_6834);
xnor U7466 (N_7466,N_6515,N_6871);
and U7467 (N_7467,N_6671,N_6814);
nand U7468 (N_7468,N_6593,N_6978);
nor U7469 (N_7469,N_6630,N_6705);
xnor U7470 (N_7470,N_6920,N_6744);
xnor U7471 (N_7471,N_6836,N_6952);
or U7472 (N_7472,N_6728,N_6863);
nand U7473 (N_7473,N_6784,N_6595);
nor U7474 (N_7474,N_6735,N_6573);
and U7475 (N_7475,N_6817,N_6858);
nor U7476 (N_7476,N_6694,N_6889);
nor U7477 (N_7477,N_6662,N_6582);
nor U7478 (N_7478,N_6703,N_6634);
nand U7479 (N_7479,N_6812,N_6905);
nor U7480 (N_7480,N_6966,N_6516);
and U7481 (N_7481,N_6890,N_6990);
nor U7482 (N_7482,N_6669,N_6946);
xnor U7483 (N_7483,N_6966,N_6916);
xnor U7484 (N_7484,N_6572,N_6910);
or U7485 (N_7485,N_6977,N_6917);
xnor U7486 (N_7486,N_6978,N_6993);
or U7487 (N_7487,N_6958,N_6788);
or U7488 (N_7488,N_6775,N_6630);
nand U7489 (N_7489,N_6906,N_6514);
nand U7490 (N_7490,N_6614,N_6586);
and U7491 (N_7491,N_6820,N_6789);
or U7492 (N_7492,N_6900,N_6653);
or U7493 (N_7493,N_6608,N_6941);
nand U7494 (N_7494,N_6657,N_6709);
nand U7495 (N_7495,N_6787,N_6551);
and U7496 (N_7496,N_6674,N_6887);
nand U7497 (N_7497,N_6854,N_6674);
xor U7498 (N_7498,N_6703,N_6771);
and U7499 (N_7499,N_6528,N_6902);
or U7500 (N_7500,N_7477,N_7353);
xor U7501 (N_7501,N_7159,N_7111);
nor U7502 (N_7502,N_7137,N_7330);
nor U7503 (N_7503,N_7141,N_7332);
xor U7504 (N_7504,N_7215,N_7211);
nand U7505 (N_7505,N_7284,N_7108);
nor U7506 (N_7506,N_7144,N_7149);
and U7507 (N_7507,N_7299,N_7323);
or U7508 (N_7508,N_7120,N_7013);
nor U7509 (N_7509,N_7088,N_7448);
xor U7510 (N_7510,N_7118,N_7272);
nand U7511 (N_7511,N_7488,N_7124);
and U7512 (N_7512,N_7132,N_7229);
or U7513 (N_7513,N_7079,N_7402);
nor U7514 (N_7514,N_7234,N_7278);
and U7515 (N_7515,N_7087,N_7240);
or U7516 (N_7516,N_7445,N_7051);
nand U7517 (N_7517,N_7400,N_7040);
nand U7518 (N_7518,N_7375,N_7189);
and U7519 (N_7519,N_7414,N_7220);
nand U7520 (N_7520,N_7316,N_7381);
and U7521 (N_7521,N_7483,N_7382);
nor U7522 (N_7522,N_7063,N_7039);
xnor U7523 (N_7523,N_7249,N_7233);
nand U7524 (N_7524,N_7188,N_7122);
and U7525 (N_7525,N_7037,N_7309);
or U7526 (N_7526,N_7101,N_7453);
or U7527 (N_7527,N_7360,N_7153);
nand U7528 (N_7528,N_7374,N_7499);
xnor U7529 (N_7529,N_7175,N_7308);
or U7530 (N_7530,N_7121,N_7471);
nor U7531 (N_7531,N_7091,N_7401);
nand U7532 (N_7532,N_7298,N_7230);
nand U7533 (N_7533,N_7378,N_7135);
xor U7534 (N_7534,N_7254,N_7105);
nand U7535 (N_7535,N_7315,N_7379);
nand U7536 (N_7536,N_7245,N_7327);
and U7537 (N_7537,N_7248,N_7075);
nand U7538 (N_7538,N_7198,N_7313);
nor U7539 (N_7539,N_7421,N_7226);
nor U7540 (N_7540,N_7092,N_7044);
nand U7541 (N_7541,N_7019,N_7251);
xor U7542 (N_7542,N_7406,N_7239);
nor U7543 (N_7543,N_7334,N_7281);
xor U7544 (N_7544,N_7097,N_7388);
xnor U7545 (N_7545,N_7033,N_7270);
and U7546 (N_7546,N_7289,N_7072);
and U7547 (N_7547,N_7224,N_7131);
xor U7548 (N_7548,N_7394,N_7209);
nand U7549 (N_7549,N_7321,N_7459);
nand U7550 (N_7550,N_7020,N_7255);
and U7551 (N_7551,N_7073,N_7271);
xnor U7552 (N_7552,N_7481,N_7086);
or U7553 (N_7553,N_7128,N_7099);
xnor U7554 (N_7554,N_7376,N_7437);
nor U7555 (N_7555,N_7026,N_7286);
nand U7556 (N_7556,N_7493,N_7403);
nand U7557 (N_7557,N_7243,N_7405);
nand U7558 (N_7558,N_7204,N_7432);
and U7559 (N_7559,N_7268,N_7373);
xnor U7560 (N_7560,N_7203,N_7438);
and U7561 (N_7561,N_7168,N_7317);
and U7562 (N_7562,N_7267,N_7146);
or U7563 (N_7563,N_7050,N_7338);
nand U7564 (N_7564,N_7335,N_7192);
or U7565 (N_7565,N_7435,N_7151);
nor U7566 (N_7566,N_7454,N_7365);
nand U7567 (N_7567,N_7498,N_7482);
nand U7568 (N_7568,N_7322,N_7126);
and U7569 (N_7569,N_7028,N_7222);
nor U7570 (N_7570,N_7328,N_7125);
nand U7571 (N_7571,N_7030,N_7319);
nand U7572 (N_7572,N_7417,N_7450);
or U7573 (N_7573,N_7350,N_7458);
nand U7574 (N_7574,N_7468,N_7015);
nor U7575 (N_7575,N_7430,N_7287);
nor U7576 (N_7576,N_7163,N_7367);
or U7577 (N_7577,N_7098,N_7006);
nor U7578 (N_7578,N_7080,N_7195);
nor U7579 (N_7579,N_7444,N_7257);
and U7580 (N_7580,N_7467,N_7193);
nor U7581 (N_7581,N_7480,N_7032);
or U7582 (N_7582,N_7491,N_7462);
or U7583 (N_7583,N_7303,N_7244);
and U7584 (N_7584,N_7312,N_7060);
or U7585 (N_7585,N_7497,N_7442);
and U7586 (N_7586,N_7059,N_7324);
and U7587 (N_7587,N_7306,N_7424);
or U7588 (N_7588,N_7179,N_7280);
or U7589 (N_7589,N_7023,N_7236);
and U7590 (N_7590,N_7354,N_7426);
xor U7591 (N_7591,N_7398,N_7484);
and U7592 (N_7592,N_7336,N_7018);
xor U7593 (N_7593,N_7235,N_7054);
and U7594 (N_7594,N_7219,N_7190);
nand U7595 (N_7595,N_7127,N_7391);
or U7596 (N_7596,N_7486,N_7082);
xor U7597 (N_7597,N_7228,N_7046);
nand U7598 (N_7598,N_7446,N_7207);
xnor U7599 (N_7599,N_7472,N_7463);
or U7600 (N_7600,N_7150,N_7218);
nor U7601 (N_7601,N_7370,N_7156);
nor U7602 (N_7602,N_7174,N_7476);
or U7603 (N_7603,N_7066,N_7343);
xnor U7604 (N_7604,N_7202,N_7451);
and U7605 (N_7605,N_7326,N_7170);
or U7606 (N_7606,N_7371,N_7333);
xnor U7607 (N_7607,N_7293,N_7404);
nand U7608 (N_7608,N_7366,N_7035);
xnor U7609 (N_7609,N_7295,N_7441);
or U7610 (N_7610,N_7173,N_7478);
or U7611 (N_7611,N_7357,N_7112);
nand U7612 (N_7612,N_7157,N_7369);
and U7613 (N_7613,N_7129,N_7297);
nand U7614 (N_7614,N_7021,N_7265);
nor U7615 (N_7615,N_7100,N_7227);
or U7616 (N_7616,N_7455,N_7247);
or U7617 (N_7617,N_7351,N_7264);
or U7618 (N_7618,N_7007,N_7138);
nand U7619 (N_7619,N_7258,N_7183);
or U7620 (N_7620,N_7489,N_7027);
and U7621 (N_7621,N_7384,N_7205);
nor U7622 (N_7622,N_7213,N_7434);
and U7623 (N_7623,N_7031,N_7169);
xor U7624 (N_7624,N_7178,N_7253);
xor U7625 (N_7625,N_7095,N_7428);
nand U7626 (N_7626,N_7440,N_7143);
xor U7627 (N_7627,N_7184,N_7003);
nor U7628 (N_7628,N_7279,N_7275);
nand U7629 (N_7629,N_7277,N_7331);
or U7630 (N_7630,N_7133,N_7110);
and U7631 (N_7631,N_7355,N_7292);
or U7632 (N_7632,N_7083,N_7492);
xor U7633 (N_7633,N_7142,N_7191);
and U7634 (N_7634,N_7147,N_7042);
or U7635 (N_7635,N_7152,N_7294);
and U7636 (N_7636,N_7436,N_7116);
nand U7637 (N_7637,N_7058,N_7305);
and U7638 (N_7638,N_7256,N_7490);
or U7639 (N_7639,N_7301,N_7396);
or U7640 (N_7640,N_7380,N_7025);
nand U7641 (N_7641,N_7109,N_7390);
or U7642 (N_7642,N_7290,N_7415);
or U7643 (N_7643,N_7136,N_7318);
nor U7644 (N_7644,N_7145,N_7241);
or U7645 (N_7645,N_7038,N_7314);
xor U7646 (N_7646,N_7464,N_7345);
xnor U7647 (N_7647,N_7155,N_7212);
and U7648 (N_7648,N_7282,N_7090);
nand U7649 (N_7649,N_7232,N_7160);
nor U7650 (N_7650,N_7016,N_7461);
nand U7651 (N_7651,N_7194,N_7022);
and U7652 (N_7652,N_7012,N_7361);
nand U7653 (N_7653,N_7176,N_7410);
xor U7654 (N_7654,N_7048,N_7061);
nor U7655 (N_7655,N_7199,N_7408);
nand U7656 (N_7656,N_7276,N_7397);
xor U7657 (N_7657,N_7036,N_7250);
nand U7658 (N_7658,N_7217,N_7096);
nor U7659 (N_7659,N_7449,N_7068);
and U7660 (N_7660,N_7005,N_7140);
xor U7661 (N_7661,N_7273,N_7231);
nand U7662 (N_7662,N_7011,N_7416);
or U7663 (N_7663,N_7342,N_7423);
nor U7664 (N_7664,N_7177,N_7344);
nand U7665 (N_7665,N_7165,N_7283);
xnor U7666 (N_7666,N_7307,N_7358);
xor U7667 (N_7667,N_7496,N_7359);
nand U7668 (N_7668,N_7115,N_7412);
and U7669 (N_7669,N_7034,N_7460);
nand U7670 (N_7670,N_7433,N_7352);
xnor U7671 (N_7671,N_7487,N_7377);
nand U7672 (N_7672,N_7356,N_7325);
and U7673 (N_7673,N_7252,N_7055);
nand U7674 (N_7674,N_7425,N_7200);
nand U7675 (N_7675,N_7368,N_7070);
or U7676 (N_7676,N_7167,N_7008);
xnor U7677 (N_7677,N_7420,N_7196);
and U7678 (N_7678,N_7427,N_7071);
xnor U7679 (N_7679,N_7182,N_7078);
xor U7680 (N_7680,N_7164,N_7310);
or U7681 (N_7681,N_7337,N_7262);
nand U7682 (N_7682,N_7085,N_7057);
or U7683 (N_7683,N_7172,N_7069);
nor U7684 (N_7684,N_7413,N_7161);
nand U7685 (N_7685,N_7246,N_7208);
and U7686 (N_7686,N_7004,N_7372);
and U7687 (N_7687,N_7171,N_7049);
nor U7688 (N_7688,N_7002,N_7296);
or U7689 (N_7689,N_7139,N_7320);
nor U7690 (N_7690,N_7485,N_7065);
nor U7691 (N_7691,N_7043,N_7102);
and U7692 (N_7692,N_7429,N_7452);
nor U7693 (N_7693,N_7134,N_7181);
xnor U7694 (N_7694,N_7389,N_7074);
or U7695 (N_7695,N_7117,N_7494);
nand U7696 (N_7696,N_7114,N_7422);
or U7697 (N_7697,N_7288,N_7154);
xor U7698 (N_7698,N_7130,N_7362);
and U7699 (N_7699,N_7443,N_7392);
or U7700 (N_7700,N_7103,N_7045);
nor U7701 (N_7701,N_7495,N_7056);
nand U7702 (N_7702,N_7214,N_7089);
nor U7703 (N_7703,N_7291,N_7067);
xor U7704 (N_7704,N_7340,N_7395);
nand U7705 (N_7705,N_7383,N_7052);
or U7706 (N_7706,N_7162,N_7465);
xnor U7707 (N_7707,N_7064,N_7041);
xor U7708 (N_7708,N_7364,N_7473);
xor U7709 (N_7709,N_7259,N_7341);
nand U7710 (N_7710,N_7479,N_7104);
or U7711 (N_7711,N_7347,N_7393);
xor U7712 (N_7712,N_7223,N_7009);
and U7713 (N_7713,N_7348,N_7387);
or U7714 (N_7714,N_7053,N_7077);
nand U7715 (N_7715,N_7339,N_7260);
nor U7716 (N_7716,N_7457,N_7386);
or U7717 (N_7717,N_7158,N_7062);
nor U7718 (N_7718,N_7411,N_7206);
xnor U7719 (N_7719,N_7261,N_7304);
nor U7720 (N_7720,N_7431,N_7419);
xor U7721 (N_7721,N_7221,N_7076);
nand U7722 (N_7722,N_7385,N_7238);
or U7723 (N_7723,N_7186,N_7000);
xor U7724 (N_7724,N_7123,N_7469);
xor U7725 (N_7725,N_7329,N_7187);
and U7726 (N_7726,N_7407,N_7024);
xor U7727 (N_7727,N_7274,N_7475);
nor U7728 (N_7728,N_7447,N_7201);
xor U7729 (N_7729,N_7399,N_7285);
or U7730 (N_7730,N_7017,N_7197);
and U7731 (N_7731,N_7456,N_7242);
or U7732 (N_7732,N_7107,N_7409);
nand U7733 (N_7733,N_7266,N_7216);
nor U7734 (N_7734,N_7225,N_7029);
nor U7735 (N_7735,N_7113,N_7119);
nor U7736 (N_7736,N_7084,N_7166);
and U7737 (N_7737,N_7148,N_7311);
or U7738 (N_7738,N_7466,N_7363);
nor U7739 (N_7739,N_7014,N_7094);
or U7740 (N_7740,N_7047,N_7474);
xnor U7741 (N_7741,N_7237,N_7210);
or U7742 (N_7742,N_7349,N_7470);
or U7743 (N_7743,N_7302,N_7185);
nor U7744 (N_7744,N_7001,N_7269);
and U7745 (N_7745,N_7010,N_7106);
or U7746 (N_7746,N_7263,N_7081);
and U7747 (N_7747,N_7180,N_7439);
and U7748 (N_7748,N_7300,N_7093);
nand U7749 (N_7749,N_7346,N_7418);
nor U7750 (N_7750,N_7055,N_7290);
nor U7751 (N_7751,N_7245,N_7165);
or U7752 (N_7752,N_7086,N_7314);
xnor U7753 (N_7753,N_7147,N_7088);
or U7754 (N_7754,N_7318,N_7193);
or U7755 (N_7755,N_7282,N_7112);
or U7756 (N_7756,N_7107,N_7292);
nand U7757 (N_7757,N_7238,N_7072);
nand U7758 (N_7758,N_7046,N_7414);
nor U7759 (N_7759,N_7172,N_7145);
nand U7760 (N_7760,N_7327,N_7187);
nor U7761 (N_7761,N_7067,N_7237);
xnor U7762 (N_7762,N_7438,N_7362);
xnor U7763 (N_7763,N_7433,N_7160);
nor U7764 (N_7764,N_7249,N_7328);
or U7765 (N_7765,N_7409,N_7213);
xor U7766 (N_7766,N_7227,N_7194);
or U7767 (N_7767,N_7303,N_7455);
xnor U7768 (N_7768,N_7156,N_7228);
or U7769 (N_7769,N_7041,N_7221);
or U7770 (N_7770,N_7164,N_7473);
nand U7771 (N_7771,N_7388,N_7434);
nand U7772 (N_7772,N_7065,N_7119);
or U7773 (N_7773,N_7461,N_7449);
nand U7774 (N_7774,N_7358,N_7468);
xor U7775 (N_7775,N_7291,N_7441);
nand U7776 (N_7776,N_7084,N_7061);
or U7777 (N_7777,N_7199,N_7353);
xor U7778 (N_7778,N_7055,N_7374);
and U7779 (N_7779,N_7250,N_7143);
nor U7780 (N_7780,N_7140,N_7300);
nand U7781 (N_7781,N_7251,N_7256);
xor U7782 (N_7782,N_7315,N_7058);
nor U7783 (N_7783,N_7151,N_7144);
and U7784 (N_7784,N_7109,N_7114);
nor U7785 (N_7785,N_7049,N_7005);
nand U7786 (N_7786,N_7000,N_7455);
xor U7787 (N_7787,N_7398,N_7107);
nor U7788 (N_7788,N_7328,N_7414);
nand U7789 (N_7789,N_7131,N_7258);
xor U7790 (N_7790,N_7312,N_7417);
or U7791 (N_7791,N_7404,N_7313);
xnor U7792 (N_7792,N_7494,N_7038);
and U7793 (N_7793,N_7383,N_7027);
and U7794 (N_7794,N_7081,N_7297);
and U7795 (N_7795,N_7301,N_7380);
or U7796 (N_7796,N_7063,N_7160);
or U7797 (N_7797,N_7272,N_7356);
or U7798 (N_7798,N_7268,N_7220);
xnor U7799 (N_7799,N_7357,N_7092);
nor U7800 (N_7800,N_7200,N_7169);
and U7801 (N_7801,N_7464,N_7463);
or U7802 (N_7802,N_7020,N_7053);
xnor U7803 (N_7803,N_7198,N_7118);
nor U7804 (N_7804,N_7054,N_7434);
nand U7805 (N_7805,N_7221,N_7153);
nor U7806 (N_7806,N_7055,N_7292);
or U7807 (N_7807,N_7040,N_7295);
xnor U7808 (N_7808,N_7173,N_7417);
and U7809 (N_7809,N_7436,N_7178);
xnor U7810 (N_7810,N_7131,N_7147);
and U7811 (N_7811,N_7004,N_7092);
xnor U7812 (N_7812,N_7200,N_7272);
and U7813 (N_7813,N_7197,N_7332);
xor U7814 (N_7814,N_7418,N_7413);
and U7815 (N_7815,N_7248,N_7240);
xnor U7816 (N_7816,N_7173,N_7493);
xnor U7817 (N_7817,N_7030,N_7476);
and U7818 (N_7818,N_7038,N_7265);
nor U7819 (N_7819,N_7028,N_7269);
nor U7820 (N_7820,N_7168,N_7461);
or U7821 (N_7821,N_7004,N_7082);
xor U7822 (N_7822,N_7255,N_7440);
nand U7823 (N_7823,N_7395,N_7058);
and U7824 (N_7824,N_7292,N_7051);
nor U7825 (N_7825,N_7421,N_7245);
nor U7826 (N_7826,N_7428,N_7219);
or U7827 (N_7827,N_7414,N_7374);
nand U7828 (N_7828,N_7013,N_7276);
or U7829 (N_7829,N_7075,N_7403);
or U7830 (N_7830,N_7178,N_7340);
or U7831 (N_7831,N_7032,N_7338);
or U7832 (N_7832,N_7109,N_7436);
nand U7833 (N_7833,N_7028,N_7387);
or U7834 (N_7834,N_7468,N_7050);
nor U7835 (N_7835,N_7472,N_7355);
or U7836 (N_7836,N_7039,N_7275);
and U7837 (N_7837,N_7206,N_7170);
nand U7838 (N_7838,N_7196,N_7312);
and U7839 (N_7839,N_7212,N_7309);
nand U7840 (N_7840,N_7006,N_7385);
nor U7841 (N_7841,N_7054,N_7426);
nor U7842 (N_7842,N_7291,N_7112);
or U7843 (N_7843,N_7476,N_7403);
nand U7844 (N_7844,N_7296,N_7065);
nand U7845 (N_7845,N_7027,N_7219);
nand U7846 (N_7846,N_7463,N_7462);
nor U7847 (N_7847,N_7496,N_7362);
or U7848 (N_7848,N_7183,N_7226);
and U7849 (N_7849,N_7410,N_7459);
or U7850 (N_7850,N_7132,N_7048);
nand U7851 (N_7851,N_7037,N_7110);
nor U7852 (N_7852,N_7407,N_7410);
and U7853 (N_7853,N_7281,N_7099);
xnor U7854 (N_7854,N_7068,N_7488);
and U7855 (N_7855,N_7374,N_7362);
or U7856 (N_7856,N_7071,N_7101);
and U7857 (N_7857,N_7212,N_7108);
nand U7858 (N_7858,N_7171,N_7069);
nor U7859 (N_7859,N_7425,N_7456);
and U7860 (N_7860,N_7268,N_7162);
or U7861 (N_7861,N_7256,N_7226);
or U7862 (N_7862,N_7018,N_7002);
xnor U7863 (N_7863,N_7015,N_7116);
nand U7864 (N_7864,N_7240,N_7046);
nand U7865 (N_7865,N_7189,N_7114);
nand U7866 (N_7866,N_7413,N_7018);
nor U7867 (N_7867,N_7494,N_7158);
xor U7868 (N_7868,N_7316,N_7161);
and U7869 (N_7869,N_7020,N_7163);
nand U7870 (N_7870,N_7376,N_7083);
xnor U7871 (N_7871,N_7351,N_7194);
nand U7872 (N_7872,N_7327,N_7057);
nor U7873 (N_7873,N_7455,N_7317);
and U7874 (N_7874,N_7381,N_7018);
nor U7875 (N_7875,N_7452,N_7391);
and U7876 (N_7876,N_7069,N_7232);
xor U7877 (N_7877,N_7318,N_7152);
nor U7878 (N_7878,N_7384,N_7403);
and U7879 (N_7879,N_7215,N_7355);
nand U7880 (N_7880,N_7355,N_7441);
nand U7881 (N_7881,N_7197,N_7274);
and U7882 (N_7882,N_7196,N_7493);
and U7883 (N_7883,N_7383,N_7070);
xnor U7884 (N_7884,N_7220,N_7237);
xnor U7885 (N_7885,N_7181,N_7294);
and U7886 (N_7886,N_7426,N_7061);
nor U7887 (N_7887,N_7041,N_7181);
nor U7888 (N_7888,N_7123,N_7016);
nand U7889 (N_7889,N_7354,N_7057);
nand U7890 (N_7890,N_7260,N_7012);
or U7891 (N_7891,N_7352,N_7241);
and U7892 (N_7892,N_7470,N_7056);
nor U7893 (N_7893,N_7344,N_7448);
or U7894 (N_7894,N_7428,N_7215);
and U7895 (N_7895,N_7091,N_7274);
nor U7896 (N_7896,N_7412,N_7108);
or U7897 (N_7897,N_7389,N_7010);
xor U7898 (N_7898,N_7083,N_7007);
or U7899 (N_7899,N_7456,N_7336);
xor U7900 (N_7900,N_7409,N_7315);
nor U7901 (N_7901,N_7497,N_7224);
or U7902 (N_7902,N_7472,N_7129);
nand U7903 (N_7903,N_7403,N_7371);
and U7904 (N_7904,N_7131,N_7151);
nor U7905 (N_7905,N_7412,N_7455);
xnor U7906 (N_7906,N_7484,N_7057);
nand U7907 (N_7907,N_7239,N_7277);
and U7908 (N_7908,N_7115,N_7154);
and U7909 (N_7909,N_7411,N_7052);
or U7910 (N_7910,N_7113,N_7007);
nor U7911 (N_7911,N_7440,N_7326);
or U7912 (N_7912,N_7175,N_7148);
nor U7913 (N_7913,N_7424,N_7097);
or U7914 (N_7914,N_7245,N_7172);
nor U7915 (N_7915,N_7090,N_7383);
and U7916 (N_7916,N_7295,N_7447);
or U7917 (N_7917,N_7104,N_7370);
nor U7918 (N_7918,N_7205,N_7282);
and U7919 (N_7919,N_7273,N_7479);
xor U7920 (N_7920,N_7389,N_7258);
or U7921 (N_7921,N_7292,N_7348);
xor U7922 (N_7922,N_7247,N_7348);
and U7923 (N_7923,N_7172,N_7371);
nand U7924 (N_7924,N_7226,N_7019);
nor U7925 (N_7925,N_7221,N_7298);
nand U7926 (N_7926,N_7352,N_7325);
nor U7927 (N_7927,N_7047,N_7461);
or U7928 (N_7928,N_7221,N_7168);
xnor U7929 (N_7929,N_7325,N_7007);
and U7930 (N_7930,N_7311,N_7270);
and U7931 (N_7931,N_7386,N_7356);
nand U7932 (N_7932,N_7403,N_7223);
nor U7933 (N_7933,N_7447,N_7229);
nand U7934 (N_7934,N_7364,N_7218);
and U7935 (N_7935,N_7220,N_7113);
and U7936 (N_7936,N_7097,N_7267);
xor U7937 (N_7937,N_7473,N_7257);
and U7938 (N_7938,N_7186,N_7311);
nand U7939 (N_7939,N_7425,N_7126);
xnor U7940 (N_7940,N_7088,N_7238);
nor U7941 (N_7941,N_7414,N_7122);
nand U7942 (N_7942,N_7004,N_7079);
nor U7943 (N_7943,N_7302,N_7042);
nand U7944 (N_7944,N_7472,N_7165);
xor U7945 (N_7945,N_7279,N_7342);
nor U7946 (N_7946,N_7101,N_7385);
nor U7947 (N_7947,N_7220,N_7047);
and U7948 (N_7948,N_7182,N_7162);
nand U7949 (N_7949,N_7120,N_7425);
or U7950 (N_7950,N_7437,N_7367);
and U7951 (N_7951,N_7423,N_7353);
nand U7952 (N_7952,N_7424,N_7269);
or U7953 (N_7953,N_7078,N_7406);
nor U7954 (N_7954,N_7470,N_7498);
xor U7955 (N_7955,N_7427,N_7080);
nand U7956 (N_7956,N_7397,N_7148);
nand U7957 (N_7957,N_7314,N_7050);
and U7958 (N_7958,N_7007,N_7130);
nor U7959 (N_7959,N_7043,N_7079);
nand U7960 (N_7960,N_7313,N_7160);
nor U7961 (N_7961,N_7213,N_7441);
nand U7962 (N_7962,N_7204,N_7065);
nand U7963 (N_7963,N_7199,N_7311);
xnor U7964 (N_7964,N_7295,N_7102);
xnor U7965 (N_7965,N_7055,N_7466);
nor U7966 (N_7966,N_7228,N_7034);
nor U7967 (N_7967,N_7318,N_7141);
nor U7968 (N_7968,N_7243,N_7370);
xor U7969 (N_7969,N_7290,N_7444);
xnor U7970 (N_7970,N_7216,N_7018);
xnor U7971 (N_7971,N_7128,N_7111);
or U7972 (N_7972,N_7295,N_7315);
xnor U7973 (N_7973,N_7123,N_7142);
nor U7974 (N_7974,N_7264,N_7496);
or U7975 (N_7975,N_7029,N_7348);
nor U7976 (N_7976,N_7087,N_7130);
xor U7977 (N_7977,N_7490,N_7396);
xor U7978 (N_7978,N_7262,N_7493);
nor U7979 (N_7979,N_7088,N_7062);
xor U7980 (N_7980,N_7273,N_7072);
nand U7981 (N_7981,N_7448,N_7407);
or U7982 (N_7982,N_7042,N_7072);
xnor U7983 (N_7983,N_7106,N_7349);
or U7984 (N_7984,N_7155,N_7048);
nand U7985 (N_7985,N_7131,N_7149);
and U7986 (N_7986,N_7395,N_7337);
nand U7987 (N_7987,N_7422,N_7132);
xnor U7988 (N_7988,N_7089,N_7023);
nor U7989 (N_7989,N_7401,N_7145);
and U7990 (N_7990,N_7063,N_7199);
or U7991 (N_7991,N_7104,N_7057);
nand U7992 (N_7992,N_7018,N_7346);
and U7993 (N_7993,N_7401,N_7323);
and U7994 (N_7994,N_7416,N_7342);
and U7995 (N_7995,N_7224,N_7445);
and U7996 (N_7996,N_7259,N_7421);
nor U7997 (N_7997,N_7061,N_7215);
xnor U7998 (N_7998,N_7251,N_7426);
xor U7999 (N_7999,N_7499,N_7167);
or U8000 (N_8000,N_7579,N_7617);
nand U8001 (N_8001,N_7709,N_7689);
nand U8002 (N_8002,N_7647,N_7973);
and U8003 (N_8003,N_7874,N_7911);
and U8004 (N_8004,N_7964,N_7908);
nand U8005 (N_8005,N_7565,N_7905);
and U8006 (N_8006,N_7615,N_7725);
nor U8007 (N_8007,N_7876,N_7504);
and U8008 (N_8008,N_7902,N_7963);
nor U8009 (N_8009,N_7954,N_7640);
nor U8010 (N_8010,N_7551,N_7711);
nor U8011 (N_8011,N_7912,N_7832);
nor U8012 (N_8012,N_7794,N_7655);
nand U8013 (N_8013,N_7920,N_7611);
xor U8014 (N_8014,N_7723,N_7641);
xor U8015 (N_8015,N_7643,N_7774);
or U8016 (N_8016,N_7522,N_7736);
nor U8017 (N_8017,N_7949,N_7695);
nand U8018 (N_8018,N_7502,N_7969);
or U8019 (N_8019,N_7914,N_7581);
and U8020 (N_8020,N_7569,N_7526);
nor U8021 (N_8021,N_7574,N_7557);
xnor U8022 (N_8022,N_7833,N_7770);
or U8023 (N_8023,N_7629,N_7596);
and U8024 (N_8024,N_7663,N_7543);
or U8025 (N_8025,N_7752,N_7505);
nor U8026 (N_8026,N_7534,N_7835);
or U8027 (N_8027,N_7999,N_7877);
nand U8028 (N_8028,N_7607,N_7939);
or U8029 (N_8029,N_7602,N_7523);
nor U8030 (N_8030,N_7866,N_7831);
xor U8031 (N_8031,N_7805,N_7981);
xnor U8032 (N_8032,N_7966,N_7823);
nand U8033 (N_8033,N_7639,N_7600);
nand U8034 (N_8034,N_7788,N_7533);
xnor U8035 (N_8035,N_7809,N_7952);
and U8036 (N_8036,N_7855,N_7759);
xor U8037 (N_8037,N_7651,N_7791);
nor U8038 (N_8038,N_7883,N_7510);
xor U8039 (N_8039,N_7932,N_7553);
xor U8040 (N_8040,N_7782,N_7775);
xor U8041 (N_8041,N_7684,N_7925);
xnor U8042 (N_8042,N_7538,N_7886);
nand U8043 (N_8043,N_7717,N_7573);
nor U8044 (N_8044,N_7900,N_7720);
nand U8045 (N_8045,N_7652,N_7636);
nand U8046 (N_8046,N_7938,N_7645);
xor U8047 (N_8047,N_7556,N_7972);
or U8048 (N_8048,N_7532,N_7758);
nand U8049 (N_8049,N_7901,N_7934);
or U8050 (N_8050,N_7895,N_7859);
or U8051 (N_8051,N_7623,N_7784);
nand U8052 (N_8052,N_7671,N_7847);
or U8053 (N_8053,N_7525,N_7864);
or U8054 (N_8054,N_7757,N_7728);
nor U8055 (N_8055,N_7624,N_7811);
and U8056 (N_8056,N_7941,N_7700);
xnor U8057 (N_8057,N_7904,N_7740);
xnor U8058 (N_8058,N_7810,N_7790);
nand U8059 (N_8059,N_7868,N_7918);
xor U8060 (N_8060,N_7890,N_7732);
nor U8061 (N_8061,N_7715,N_7635);
or U8062 (N_8062,N_7769,N_7796);
nor U8063 (N_8063,N_7985,N_7508);
and U8064 (N_8064,N_7708,N_7781);
nand U8065 (N_8065,N_7706,N_7692);
and U8066 (N_8066,N_7862,N_7967);
nor U8067 (N_8067,N_7899,N_7827);
or U8068 (N_8068,N_7540,N_7677);
and U8069 (N_8069,N_7649,N_7806);
and U8070 (N_8070,N_7539,N_7776);
nand U8071 (N_8071,N_7873,N_7850);
nor U8072 (N_8072,N_7944,N_7586);
nand U8073 (N_8073,N_7755,N_7633);
xnor U8074 (N_8074,N_7846,N_7664);
nand U8075 (N_8075,N_7749,N_7675);
xnor U8076 (N_8076,N_7898,N_7892);
or U8077 (N_8077,N_7962,N_7906);
xnor U8078 (N_8078,N_7991,N_7785);
or U8079 (N_8079,N_7527,N_7764);
nor U8080 (N_8080,N_7848,N_7976);
nor U8081 (N_8081,N_7975,N_7824);
or U8082 (N_8082,N_7628,N_7506);
nand U8083 (N_8083,N_7885,N_7638);
nand U8084 (N_8084,N_7658,N_7562);
nor U8085 (N_8085,N_7860,N_7995);
xor U8086 (N_8086,N_7753,N_7974);
nand U8087 (N_8087,N_7798,N_7993);
nor U8088 (N_8088,N_7683,N_7550);
xor U8089 (N_8089,N_7982,N_7997);
nor U8090 (N_8090,N_7767,N_7878);
nor U8091 (N_8091,N_7891,N_7722);
nor U8092 (N_8092,N_7828,N_7585);
nor U8093 (N_8093,N_7818,N_7697);
or U8094 (N_8094,N_7604,N_7567);
nor U8095 (N_8095,N_7894,N_7968);
and U8096 (N_8096,N_7509,N_7821);
nand U8097 (N_8097,N_7515,N_7744);
nor U8098 (N_8098,N_7836,N_7730);
nand U8099 (N_8099,N_7512,N_7544);
and U8100 (N_8100,N_7632,N_7531);
nor U8101 (N_8101,N_7681,N_7867);
or U8102 (N_8102,N_7698,N_7875);
or U8103 (N_8103,N_7936,N_7977);
or U8104 (N_8104,N_7598,N_7983);
xor U8105 (N_8105,N_7731,N_7880);
and U8106 (N_8106,N_7559,N_7609);
or U8107 (N_8107,N_7958,N_7516);
and U8108 (N_8108,N_7853,N_7924);
and U8109 (N_8109,N_7852,N_7595);
nor U8110 (N_8110,N_7668,N_7584);
nor U8111 (N_8111,N_7676,N_7889);
xor U8112 (N_8112,N_7535,N_7814);
or U8113 (N_8113,N_7729,N_7577);
xnor U8114 (N_8114,N_7678,N_7702);
xnor U8115 (N_8115,N_7923,N_7916);
or U8116 (N_8116,N_7858,N_7674);
xnor U8117 (N_8117,N_7915,N_7503);
and U8118 (N_8118,N_7738,N_7558);
nand U8119 (N_8119,N_7897,N_7800);
and U8120 (N_8120,N_7673,N_7945);
or U8121 (N_8121,N_7951,N_7619);
nand U8122 (N_8122,N_7568,N_7820);
and U8123 (N_8123,N_7998,N_7741);
nand U8124 (N_8124,N_7903,N_7605);
or U8125 (N_8125,N_7802,N_7869);
nand U8126 (N_8126,N_7682,N_7688);
or U8127 (N_8127,N_7771,N_7537);
xor U8128 (N_8128,N_7960,N_7735);
or U8129 (N_8129,N_7825,N_7590);
nor U8130 (N_8130,N_7739,N_7947);
xor U8131 (N_8131,N_7583,N_7829);
nand U8132 (N_8132,N_7884,N_7524);
and U8133 (N_8133,N_7988,N_7815);
xor U8134 (N_8134,N_7801,N_7804);
nand U8135 (N_8135,N_7563,N_7946);
nand U8136 (N_8136,N_7760,N_7787);
nor U8137 (N_8137,N_7888,N_7879);
nor U8138 (N_8138,N_7777,N_7959);
xor U8139 (N_8139,N_7511,N_7546);
nor U8140 (N_8140,N_7909,N_7789);
nor U8141 (N_8141,N_7786,N_7746);
nor U8142 (N_8142,N_7718,N_7965);
xor U8143 (N_8143,N_7703,N_7705);
xnor U8144 (N_8144,N_7528,N_7710);
nor U8145 (N_8145,N_7521,N_7630);
and U8146 (N_8146,N_7845,N_7606);
nor U8147 (N_8147,N_7616,N_7513);
nand U8148 (N_8148,N_7554,N_7566);
or U8149 (N_8149,N_7768,N_7953);
nor U8150 (N_8150,N_7541,N_7816);
or U8151 (N_8151,N_7907,N_7627);
or U8152 (N_8152,N_7561,N_7844);
xor U8153 (N_8153,N_7817,N_7970);
or U8154 (N_8154,N_7765,N_7589);
xor U8155 (N_8155,N_7612,N_7727);
nand U8156 (N_8156,N_7704,N_7956);
nand U8157 (N_8157,N_7662,N_7733);
and U8158 (N_8158,N_7530,N_7854);
nand U8159 (N_8159,N_7992,N_7871);
nand U8160 (N_8160,N_7694,N_7919);
nand U8161 (N_8161,N_7762,N_7849);
nor U8162 (N_8162,N_7693,N_7672);
nand U8163 (N_8163,N_7575,N_7792);
nor U8164 (N_8164,N_7564,N_7646);
xnor U8165 (N_8165,N_7699,N_7716);
xor U8166 (N_8166,N_7592,N_7742);
or U8167 (N_8167,N_7631,N_7656);
and U8168 (N_8168,N_7926,N_7780);
nand U8169 (N_8169,N_7893,N_7648);
or U8170 (N_8170,N_7552,N_7665);
or U8171 (N_8171,N_7734,N_7594);
nor U8172 (N_8172,N_7763,N_7591);
nand U8173 (N_8173,N_7950,N_7813);
xnor U8174 (N_8174,N_7549,N_7870);
and U8175 (N_8175,N_7943,N_7626);
and U8176 (N_8176,N_7984,N_7979);
or U8177 (N_8177,N_7667,N_7857);
xor U8178 (N_8178,N_7642,N_7536);
or U8179 (N_8179,N_7547,N_7657);
nor U8180 (N_8180,N_7929,N_7834);
xnor U8181 (N_8181,N_7987,N_7696);
nand U8182 (N_8182,N_7935,N_7601);
nor U8183 (N_8183,N_7588,N_7756);
or U8184 (N_8184,N_7913,N_7778);
or U8185 (N_8185,N_7518,N_7882);
and U8186 (N_8186,N_7955,N_7865);
nand U8187 (N_8187,N_7707,N_7807);
xnor U8188 (N_8188,N_7654,N_7793);
and U8189 (N_8189,N_7921,N_7578);
xnor U8190 (N_8190,N_7761,N_7957);
nand U8191 (N_8191,N_7773,N_7940);
xnor U8192 (N_8192,N_7856,N_7724);
nand U8193 (N_8193,N_7830,N_7726);
nand U8194 (N_8194,N_7634,N_7837);
nor U8195 (N_8195,N_7661,N_7961);
nor U8196 (N_8196,N_7520,N_7529);
nor U8197 (N_8197,N_7670,N_7599);
nand U8198 (N_8198,N_7686,N_7861);
or U8199 (N_8199,N_7989,N_7701);
nand U8200 (N_8200,N_7603,N_7560);
xor U8201 (N_8201,N_7712,N_7679);
and U8202 (N_8202,N_7795,N_7803);
or U8203 (N_8203,N_7622,N_7571);
or U8204 (N_8204,N_7841,N_7650);
and U8205 (N_8205,N_7822,N_7620);
xnor U8206 (N_8206,N_7501,N_7517);
nor U8207 (N_8207,N_7881,N_7500);
nand U8208 (N_8208,N_7930,N_7576);
nand U8209 (N_8209,N_7779,N_7719);
nand U8210 (N_8210,N_7843,N_7548);
xor U8211 (N_8211,N_7910,N_7863);
or U8212 (N_8212,N_7986,N_7713);
nor U8213 (N_8213,N_7937,N_7754);
nand U8214 (N_8214,N_7747,N_7545);
or U8215 (N_8215,N_7570,N_7519);
nand U8216 (N_8216,N_7572,N_7721);
nor U8217 (N_8217,N_7597,N_7582);
xor U8218 (N_8218,N_7990,N_7842);
and U8219 (N_8219,N_7772,N_7980);
nor U8220 (N_8220,N_7614,N_7743);
xor U8221 (N_8221,N_7687,N_7610);
and U8222 (N_8222,N_7542,N_7839);
xor U8223 (N_8223,N_7872,N_7851);
nand U8224 (N_8224,N_7887,N_7751);
nor U8225 (N_8225,N_7927,N_7690);
nand U8226 (N_8226,N_7808,N_7797);
xnor U8227 (N_8227,N_7948,N_7660);
nor U8228 (N_8228,N_7838,N_7587);
and U8229 (N_8229,N_7766,N_7621);
nand U8230 (N_8230,N_7737,N_7637);
or U8231 (N_8231,N_7799,N_7593);
or U8232 (N_8232,N_7896,N_7931);
nor U8233 (N_8233,N_7691,N_7608);
xor U8234 (N_8234,N_7783,N_7928);
xor U8235 (N_8235,N_7971,N_7922);
or U8236 (N_8236,N_7653,N_7996);
nand U8237 (N_8237,N_7507,N_7826);
nor U8238 (N_8238,N_7840,N_7514);
and U8239 (N_8239,N_7812,N_7745);
nand U8240 (N_8240,N_7680,N_7625);
xnor U8241 (N_8241,N_7659,N_7748);
or U8242 (N_8242,N_7917,N_7669);
or U8243 (N_8243,N_7819,N_7618);
nor U8244 (N_8244,N_7685,N_7978);
or U8245 (N_8245,N_7555,N_7994);
nor U8246 (N_8246,N_7750,N_7942);
and U8247 (N_8247,N_7644,N_7933);
nand U8248 (N_8248,N_7580,N_7666);
nor U8249 (N_8249,N_7714,N_7613);
nand U8250 (N_8250,N_7964,N_7551);
xor U8251 (N_8251,N_7911,N_7506);
nor U8252 (N_8252,N_7561,N_7635);
or U8253 (N_8253,N_7864,N_7682);
xnor U8254 (N_8254,N_7908,N_7788);
nor U8255 (N_8255,N_7881,N_7666);
nand U8256 (N_8256,N_7570,N_7569);
nand U8257 (N_8257,N_7514,N_7587);
nor U8258 (N_8258,N_7739,N_7610);
xor U8259 (N_8259,N_7649,N_7610);
nor U8260 (N_8260,N_7621,N_7849);
nand U8261 (N_8261,N_7642,N_7573);
xor U8262 (N_8262,N_7700,N_7574);
nor U8263 (N_8263,N_7638,N_7966);
xnor U8264 (N_8264,N_7671,N_7938);
nor U8265 (N_8265,N_7803,N_7818);
or U8266 (N_8266,N_7635,N_7508);
and U8267 (N_8267,N_7691,N_7964);
xor U8268 (N_8268,N_7856,N_7912);
nor U8269 (N_8269,N_7983,N_7866);
xor U8270 (N_8270,N_7810,N_7504);
and U8271 (N_8271,N_7896,N_7968);
or U8272 (N_8272,N_7566,N_7777);
nand U8273 (N_8273,N_7776,N_7830);
or U8274 (N_8274,N_7671,N_7903);
xnor U8275 (N_8275,N_7536,N_7891);
xor U8276 (N_8276,N_7976,N_7591);
and U8277 (N_8277,N_7650,N_7911);
nand U8278 (N_8278,N_7610,N_7792);
or U8279 (N_8279,N_7884,N_7950);
nand U8280 (N_8280,N_7670,N_7598);
or U8281 (N_8281,N_7889,N_7911);
xor U8282 (N_8282,N_7969,N_7735);
xnor U8283 (N_8283,N_7508,N_7835);
nand U8284 (N_8284,N_7991,N_7909);
xor U8285 (N_8285,N_7757,N_7664);
nor U8286 (N_8286,N_7536,N_7727);
and U8287 (N_8287,N_7820,N_7923);
nor U8288 (N_8288,N_7987,N_7709);
nor U8289 (N_8289,N_7504,N_7952);
nor U8290 (N_8290,N_7700,N_7835);
nor U8291 (N_8291,N_7971,N_7820);
and U8292 (N_8292,N_7879,N_7549);
xor U8293 (N_8293,N_7504,N_7708);
xor U8294 (N_8294,N_7802,N_7841);
and U8295 (N_8295,N_7627,N_7585);
and U8296 (N_8296,N_7732,N_7788);
xnor U8297 (N_8297,N_7651,N_7891);
xor U8298 (N_8298,N_7765,N_7581);
nor U8299 (N_8299,N_7809,N_7886);
xor U8300 (N_8300,N_7669,N_7523);
or U8301 (N_8301,N_7705,N_7650);
nor U8302 (N_8302,N_7853,N_7567);
nor U8303 (N_8303,N_7781,N_7794);
nor U8304 (N_8304,N_7679,N_7763);
and U8305 (N_8305,N_7500,N_7983);
and U8306 (N_8306,N_7886,N_7864);
and U8307 (N_8307,N_7799,N_7608);
and U8308 (N_8308,N_7573,N_7809);
or U8309 (N_8309,N_7600,N_7560);
xnor U8310 (N_8310,N_7528,N_7890);
or U8311 (N_8311,N_7574,N_7664);
xor U8312 (N_8312,N_7910,N_7959);
nand U8313 (N_8313,N_7659,N_7963);
or U8314 (N_8314,N_7657,N_7999);
nand U8315 (N_8315,N_7607,N_7685);
nor U8316 (N_8316,N_7888,N_7760);
and U8317 (N_8317,N_7700,N_7928);
xor U8318 (N_8318,N_7727,N_7558);
and U8319 (N_8319,N_7674,N_7849);
nand U8320 (N_8320,N_7920,N_7816);
nand U8321 (N_8321,N_7898,N_7896);
xnor U8322 (N_8322,N_7681,N_7554);
xor U8323 (N_8323,N_7620,N_7568);
nand U8324 (N_8324,N_7902,N_7523);
or U8325 (N_8325,N_7637,N_7694);
xor U8326 (N_8326,N_7535,N_7883);
or U8327 (N_8327,N_7580,N_7551);
nor U8328 (N_8328,N_7619,N_7959);
xnor U8329 (N_8329,N_7998,N_7795);
or U8330 (N_8330,N_7582,N_7561);
xor U8331 (N_8331,N_7615,N_7900);
nand U8332 (N_8332,N_7908,N_7837);
nand U8333 (N_8333,N_7766,N_7979);
and U8334 (N_8334,N_7697,N_7523);
and U8335 (N_8335,N_7601,N_7864);
or U8336 (N_8336,N_7846,N_7967);
nor U8337 (N_8337,N_7607,N_7551);
and U8338 (N_8338,N_7881,N_7624);
xor U8339 (N_8339,N_7569,N_7724);
nor U8340 (N_8340,N_7751,N_7932);
or U8341 (N_8341,N_7648,N_7917);
and U8342 (N_8342,N_7935,N_7564);
xnor U8343 (N_8343,N_7507,N_7522);
and U8344 (N_8344,N_7771,N_7746);
or U8345 (N_8345,N_7810,N_7519);
and U8346 (N_8346,N_7558,N_7625);
nor U8347 (N_8347,N_7519,N_7854);
and U8348 (N_8348,N_7637,N_7739);
and U8349 (N_8349,N_7874,N_7820);
nor U8350 (N_8350,N_7672,N_7817);
and U8351 (N_8351,N_7763,N_7529);
and U8352 (N_8352,N_7829,N_7882);
nand U8353 (N_8353,N_7831,N_7828);
nor U8354 (N_8354,N_7898,N_7914);
nor U8355 (N_8355,N_7924,N_7586);
xor U8356 (N_8356,N_7677,N_7583);
xnor U8357 (N_8357,N_7695,N_7611);
xnor U8358 (N_8358,N_7965,N_7734);
nand U8359 (N_8359,N_7586,N_7997);
or U8360 (N_8360,N_7647,N_7991);
nor U8361 (N_8361,N_7925,N_7715);
or U8362 (N_8362,N_7747,N_7561);
and U8363 (N_8363,N_7504,N_7950);
and U8364 (N_8364,N_7585,N_7882);
and U8365 (N_8365,N_7711,N_7954);
xnor U8366 (N_8366,N_7613,N_7852);
xor U8367 (N_8367,N_7551,N_7556);
xor U8368 (N_8368,N_7604,N_7642);
nor U8369 (N_8369,N_7859,N_7539);
or U8370 (N_8370,N_7971,N_7953);
or U8371 (N_8371,N_7639,N_7586);
and U8372 (N_8372,N_7518,N_7730);
nor U8373 (N_8373,N_7775,N_7923);
and U8374 (N_8374,N_7657,N_7971);
or U8375 (N_8375,N_7944,N_7697);
nand U8376 (N_8376,N_7730,N_7674);
nand U8377 (N_8377,N_7898,N_7931);
or U8378 (N_8378,N_7655,N_7826);
and U8379 (N_8379,N_7857,N_7709);
or U8380 (N_8380,N_7653,N_7781);
nand U8381 (N_8381,N_7792,N_7767);
or U8382 (N_8382,N_7832,N_7928);
nor U8383 (N_8383,N_7929,N_7842);
xnor U8384 (N_8384,N_7745,N_7919);
xnor U8385 (N_8385,N_7854,N_7735);
and U8386 (N_8386,N_7649,N_7585);
or U8387 (N_8387,N_7992,N_7759);
or U8388 (N_8388,N_7802,N_7839);
nor U8389 (N_8389,N_7848,N_7527);
and U8390 (N_8390,N_7559,N_7723);
and U8391 (N_8391,N_7840,N_7527);
or U8392 (N_8392,N_7910,N_7964);
xor U8393 (N_8393,N_7729,N_7813);
nor U8394 (N_8394,N_7563,N_7640);
nor U8395 (N_8395,N_7719,N_7780);
xnor U8396 (N_8396,N_7684,N_7715);
xnor U8397 (N_8397,N_7996,N_7546);
nor U8398 (N_8398,N_7622,N_7829);
and U8399 (N_8399,N_7754,N_7896);
xor U8400 (N_8400,N_7519,N_7968);
or U8401 (N_8401,N_7520,N_7658);
or U8402 (N_8402,N_7753,N_7890);
and U8403 (N_8403,N_7801,N_7949);
nor U8404 (N_8404,N_7664,N_7560);
nand U8405 (N_8405,N_7676,N_7761);
nor U8406 (N_8406,N_7730,N_7963);
nor U8407 (N_8407,N_7628,N_7526);
and U8408 (N_8408,N_7708,N_7638);
nor U8409 (N_8409,N_7582,N_7750);
or U8410 (N_8410,N_7781,N_7755);
or U8411 (N_8411,N_7653,N_7526);
or U8412 (N_8412,N_7881,N_7529);
or U8413 (N_8413,N_7892,N_7640);
xor U8414 (N_8414,N_7803,N_7879);
and U8415 (N_8415,N_7940,N_7913);
or U8416 (N_8416,N_7613,N_7814);
nand U8417 (N_8417,N_7873,N_7674);
xnor U8418 (N_8418,N_7555,N_7802);
or U8419 (N_8419,N_7632,N_7570);
or U8420 (N_8420,N_7510,N_7735);
xnor U8421 (N_8421,N_7583,N_7918);
or U8422 (N_8422,N_7834,N_7634);
nand U8423 (N_8423,N_7898,N_7717);
and U8424 (N_8424,N_7845,N_7514);
nand U8425 (N_8425,N_7730,N_7687);
nor U8426 (N_8426,N_7562,N_7754);
nand U8427 (N_8427,N_7994,N_7661);
nor U8428 (N_8428,N_7550,N_7912);
nand U8429 (N_8429,N_7538,N_7643);
nand U8430 (N_8430,N_7733,N_7596);
nor U8431 (N_8431,N_7545,N_7844);
xor U8432 (N_8432,N_7801,N_7605);
nor U8433 (N_8433,N_7737,N_7630);
or U8434 (N_8434,N_7516,N_7706);
nor U8435 (N_8435,N_7981,N_7873);
xnor U8436 (N_8436,N_7777,N_7912);
nor U8437 (N_8437,N_7796,N_7965);
nand U8438 (N_8438,N_7989,N_7699);
xnor U8439 (N_8439,N_7852,N_7688);
xor U8440 (N_8440,N_7874,N_7989);
xnor U8441 (N_8441,N_7981,N_7524);
or U8442 (N_8442,N_7783,N_7574);
or U8443 (N_8443,N_7984,N_7921);
xnor U8444 (N_8444,N_7743,N_7819);
nand U8445 (N_8445,N_7717,N_7977);
xnor U8446 (N_8446,N_7755,N_7805);
and U8447 (N_8447,N_7738,N_7897);
or U8448 (N_8448,N_7904,N_7891);
xor U8449 (N_8449,N_7628,N_7522);
nor U8450 (N_8450,N_7634,N_7888);
nor U8451 (N_8451,N_7987,N_7636);
nor U8452 (N_8452,N_7705,N_7558);
nor U8453 (N_8453,N_7572,N_7916);
nand U8454 (N_8454,N_7994,N_7581);
nor U8455 (N_8455,N_7670,N_7883);
xnor U8456 (N_8456,N_7804,N_7709);
nand U8457 (N_8457,N_7672,N_7984);
and U8458 (N_8458,N_7675,N_7806);
or U8459 (N_8459,N_7914,N_7851);
xnor U8460 (N_8460,N_7837,N_7757);
nor U8461 (N_8461,N_7778,N_7611);
nand U8462 (N_8462,N_7645,N_7557);
or U8463 (N_8463,N_7712,N_7771);
xnor U8464 (N_8464,N_7854,N_7670);
nand U8465 (N_8465,N_7851,N_7994);
or U8466 (N_8466,N_7784,N_7617);
and U8467 (N_8467,N_7716,N_7616);
and U8468 (N_8468,N_7578,N_7575);
xnor U8469 (N_8469,N_7662,N_7539);
and U8470 (N_8470,N_7974,N_7648);
xor U8471 (N_8471,N_7661,N_7830);
xor U8472 (N_8472,N_7651,N_7544);
or U8473 (N_8473,N_7503,N_7895);
nor U8474 (N_8474,N_7833,N_7832);
and U8475 (N_8475,N_7595,N_7716);
or U8476 (N_8476,N_7963,N_7597);
nor U8477 (N_8477,N_7902,N_7718);
or U8478 (N_8478,N_7991,N_7678);
nor U8479 (N_8479,N_7531,N_7774);
xor U8480 (N_8480,N_7918,N_7677);
nand U8481 (N_8481,N_7874,N_7981);
xor U8482 (N_8482,N_7650,N_7932);
xor U8483 (N_8483,N_7923,N_7798);
and U8484 (N_8484,N_7826,N_7893);
nor U8485 (N_8485,N_7634,N_7991);
and U8486 (N_8486,N_7939,N_7683);
nor U8487 (N_8487,N_7787,N_7877);
and U8488 (N_8488,N_7652,N_7833);
or U8489 (N_8489,N_7825,N_7791);
nor U8490 (N_8490,N_7722,N_7704);
xor U8491 (N_8491,N_7551,N_7636);
nand U8492 (N_8492,N_7589,N_7786);
nor U8493 (N_8493,N_7935,N_7532);
xor U8494 (N_8494,N_7529,N_7698);
and U8495 (N_8495,N_7990,N_7756);
and U8496 (N_8496,N_7660,N_7526);
nand U8497 (N_8497,N_7519,N_7872);
xor U8498 (N_8498,N_7906,N_7550);
xnor U8499 (N_8499,N_7535,N_7889);
xnor U8500 (N_8500,N_8445,N_8102);
nand U8501 (N_8501,N_8186,N_8428);
nand U8502 (N_8502,N_8296,N_8224);
and U8503 (N_8503,N_8434,N_8150);
or U8504 (N_8504,N_8392,N_8446);
nor U8505 (N_8505,N_8462,N_8163);
nor U8506 (N_8506,N_8087,N_8376);
nand U8507 (N_8507,N_8255,N_8030);
or U8508 (N_8508,N_8318,N_8013);
xnor U8509 (N_8509,N_8362,N_8471);
or U8510 (N_8510,N_8088,N_8472);
nor U8511 (N_8511,N_8114,N_8327);
nor U8512 (N_8512,N_8099,N_8192);
or U8513 (N_8513,N_8419,N_8009);
or U8514 (N_8514,N_8203,N_8231);
nand U8515 (N_8515,N_8389,N_8242);
nor U8516 (N_8516,N_8152,N_8371);
nor U8517 (N_8517,N_8041,N_8122);
nor U8518 (N_8518,N_8218,N_8006);
and U8519 (N_8519,N_8024,N_8490);
and U8520 (N_8520,N_8207,N_8067);
nand U8521 (N_8521,N_8279,N_8495);
nor U8522 (N_8522,N_8104,N_8251);
xnor U8523 (N_8523,N_8200,N_8314);
or U8524 (N_8524,N_8188,N_8345);
or U8525 (N_8525,N_8388,N_8351);
or U8526 (N_8526,N_8005,N_8299);
xnor U8527 (N_8527,N_8414,N_8265);
and U8528 (N_8528,N_8425,N_8205);
and U8529 (N_8529,N_8080,N_8078);
or U8530 (N_8530,N_8451,N_8011);
nand U8531 (N_8531,N_8461,N_8032);
xor U8532 (N_8532,N_8131,N_8214);
nor U8533 (N_8533,N_8086,N_8381);
nor U8534 (N_8534,N_8353,N_8499);
and U8535 (N_8535,N_8328,N_8177);
nor U8536 (N_8536,N_8473,N_8089);
or U8537 (N_8537,N_8485,N_8158);
nor U8538 (N_8538,N_8190,N_8393);
or U8539 (N_8539,N_8326,N_8491);
and U8540 (N_8540,N_8139,N_8031);
xnor U8541 (N_8541,N_8054,N_8494);
and U8542 (N_8542,N_8208,N_8240);
nand U8543 (N_8543,N_8154,N_8386);
or U8544 (N_8544,N_8250,N_8145);
and U8545 (N_8545,N_8452,N_8341);
xor U8546 (N_8546,N_8406,N_8090);
nand U8547 (N_8547,N_8226,N_8420);
or U8548 (N_8548,N_8132,N_8256);
nor U8549 (N_8549,N_8404,N_8047);
nor U8550 (N_8550,N_8426,N_8480);
and U8551 (N_8551,N_8064,N_8412);
xor U8552 (N_8552,N_8295,N_8026);
or U8553 (N_8553,N_8292,N_8140);
nor U8554 (N_8554,N_8243,N_8021);
and U8555 (N_8555,N_8234,N_8098);
or U8556 (N_8556,N_8123,N_8229);
nand U8557 (N_8557,N_8146,N_8320);
or U8558 (N_8558,N_8394,N_8276);
nand U8559 (N_8559,N_8117,N_8331);
or U8560 (N_8560,N_8179,N_8033);
nor U8561 (N_8561,N_8058,N_8196);
or U8562 (N_8562,N_8217,N_8144);
nand U8563 (N_8563,N_8194,N_8361);
or U8564 (N_8564,N_8227,N_8138);
xor U8565 (N_8565,N_8010,N_8166);
or U8566 (N_8566,N_8252,N_8288);
nor U8567 (N_8567,N_8346,N_8258);
nand U8568 (N_8568,N_8468,N_8036);
nand U8569 (N_8569,N_8083,N_8421);
and U8570 (N_8570,N_8336,N_8043);
nand U8571 (N_8571,N_8093,N_8284);
nor U8572 (N_8572,N_8180,N_8055);
nor U8573 (N_8573,N_8219,N_8246);
or U8574 (N_8574,N_8034,N_8312);
xnor U8575 (N_8575,N_8113,N_8498);
nor U8576 (N_8576,N_8316,N_8198);
xnor U8577 (N_8577,N_8079,N_8437);
xnor U8578 (N_8578,N_8359,N_8189);
xnor U8579 (N_8579,N_8081,N_8489);
xnor U8580 (N_8580,N_8294,N_8211);
nand U8581 (N_8581,N_8176,N_8474);
or U8582 (N_8582,N_8103,N_8470);
nand U8583 (N_8583,N_8124,N_8348);
nor U8584 (N_8584,N_8457,N_8249);
and U8585 (N_8585,N_8382,N_8477);
or U8586 (N_8586,N_8197,N_8168);
nor U8587 (N_8587,N_8486,N_8069);
nor U8588 (N_8588,N_8370,N_8304);
nand U8589 (N_8589,N_8161,N_8478);
and U8590 (N_8590,N_8051,N_8379);
xor U8591 (N_8591,N_8440,N_8096);
xor U8592 (N_8592,N_8280,N_8398);
or U8593 (N_8593,N_8149,N_8071);
or U8594 (N_8594,N_8357,N_8308);
or U8595 (N_8595,N_8247,N_8016);
nor U8596 (N_8596,N_8142,N_8063);
nand U8597 (N_8597,N_8003,N_8097);
nand U8598 (N_8598,N_8027,N_8044);
nor U8599 (N_8599,N_8125,N_8390);
and U8600 (N_8600,N_8395,N_8143);
and U8601 (N_8601,N_8048,N_8397);
xnor U8602 (N_8602,N_8482,N_8402);
or U8603 (N_8603,N_8156,N_8065);
and U8604 (N_8604,N_8342,N_8344);
xor U8605 (N_8605,N_8193,N_8422);
nand U8606 (N_8606,N_8171,N_8223);
or U8607 (N_8607,N_8002,N_8059);
or U8608 (N_8608,N_8343,N_8245);
nand U8609 (N_8609,N_8233,N_8259);
xnor U8610 (N_8610,N_8238,N_8228);
nor U8611 (N_8611,N_8385,N_8378);
or U8612 (N_8612,N_8297,N_8022);
xnor U8613 (N_8613,N_8306,N_8372);
and U8614 (N_8614,N_8195,N_8281);
nor U8615 (N_8615,N_8173,N_8355);
and U8616 (N_8616,N_8282,N_8191);
or U8617 (N_8617,N_8453,N_8384);
nor U8618 (N_8618,N_8286,N_8014);
nor U8619 (N_8619,N_8025,N_8263);
nor U8620 (N_8620,N_8182,N_8164);
and U8621 (N_8621,N_8201,N_8109);
and U8622 (N_8622,N_8447,N_8137);
and U8623 (N_8623,N_8315,N_8349);
and U8624 (N_8624,N_8220,N_8264);
nand U8625 (N_8625,N_8313,N_8070);
or U8626 (N_8626,N_8038,N_8007);
or U8627 (N_8627,N_8028,N_8112);
and U8628 (N_8628,N_8206,N_8374);
or U8629 (N_8629,N_8363,N_8438);
xnor U8630 (N_8630,N_8293,N_8039);
nand U8631 (N_8631,N_8111,N_8460);
nand U8632 (N_8632,N_8052,N_8317);
xor U8633 (N_8633,N_8001,N_8432);
nor U8634 (N_8634,N_8339,N_8147);
nand U8635 (N_8635,N_8085,N_8366);
xor U8636 (N_8636,N_8105,N_8153);
xnor U8637 (N_8637,N_8274,N_8133);
nand U8638 (N_8638,N_8107,N_8298);
nor U8639 (N_8639,N_8458,N_8488);
xnor U8640 (N_8640,N_8347,N_8209);
nand U8641 (N_8641,N_8060,N_8450);
xor U8642 (N_8642,N_8354,N_8202);
nand U8643 (N_8643,N_8178,N_8364);
xnor U8644 (N_8644,N_8023,N_8165);
nor U8645 (N_8645,N_8268,N_8415);
xnor U8646 (N_8646,N_8467,N_8322);
and U8647 (N_8647,N_8020,N_8260);
or U8648 (N_8648,N_8046,N_8424);
xnor U8649 (N_8649,N_8285,N_8019);
nand U8650 (N_8650,N_8056,N_8305);
or U8651 (N_8651,N_8082,N_8230);
xor U8652 (N_8652,N_8101,N_8466);
nor U8653 (N_8653,N_8204,N_8443);
and U8654 (N_8654,N_8187,N_8335);
and U8655 (N_8655,N_8235,N_8045);
or U8656 (N_8656,N_8456,N_8319);
xnor U8657 (N_8657,N_8405,N_8075);
xor U8658 (N_8658,N_8053,N_8411);
xor U8659 (N_8659,N_8118,N_8135);
nand U8660 (N_8660,N_8169,N_8329);
xnor U8661 (N_8661,N_8377,N_8273);
nand U8662 (N_8662,N_8232,N_8254);
and U8663 (N_8663,N_8418,N_8479);
nor U8664 (N_8664,N_8492,N_8072);
nor U8665 (N_8665,N_8387,N_8066);
or U8666 (N_8666,N_8403,N_8134);
nand U8667 (N_8667,N_8035,N_8391);
xor U8668 (N_8668,N_8004,N_8215);
nand U8669 (N_8669,N_8162,N_8433);
xnor U8670 (N_8670,N_8119,N_8184);
nand U8671 (N_8671,N_8100,N_8185);
or U8672 (N_8672,N_8091,N_8222);
nand U8673 (N_8673,N_8108,N_8040);
nand U8674 (N_8674,N_8413,N_8455);
xor U8675 (N_8675,N_8018,N_8309);
and U8676 (N_8676,N_8278,N_8431);
or U8677 (N_8677,N_8487,N_8483);
or U8678 (N_8678,N_8074,N_8175);
and U8679 (N_8679,N_8429,N_8465);
nor U8680 (N_8680,N_8350,N_8283);
and U8681 (N_8681,N_8365,N_8307);
or U8682 (N_8682,N_8449,N_8241);
or U8683 (N_8683,N_8049,N_8401);
nand U8684 (N_8684,N_8257,N_8213);
nor U8685 (N_8685,N_8266,N_8287);
nor U8686 (N_8686,N_8454,N_8076);
xor U8687 (N_8687,N_8225,N_8464);
and U8688 (N_8688,N_8126,N_8267);
nor U8689 (N_8689,N_8157,N_8476);
nand U8690 (N_8690,N_8311,N_8248);
or U8691 (N_8691,N_8210,N_8172);
xor U8692 (N_8692,N_8399,N_8121);
nor U8693 (N_8693,N_8442,N_8077);
xnor U8694 (N_8694,N_8110,N_8360);
nand U8695 (N_8695,N_8130,N_8237);
nor U8696 (N_8696,N_8330,N_8496);
xnor U8697 (N_8697,N_8050,N_8160);
nor U8698 (N_8698,N_8106,N_8324);
and U8699 (N_8699,N_8310,N_8373);
nand U8700 (N_8700,N_8136,N_8272);
nor U8701 (N_8701,N_8095,N_8352);
or U8702 (N_8702,N_8061,N_8369);
nor U8703 (N_8703,N_8000,N_8430);
or U8704 (N_8704,N_8261,N_8356);
nand U8705 (N_8705,N_8417,N_8170);
or U8706 (N_8706,N_8441,N_8380);
and U8707 (N_8707,N_8435,N_8244);
or U8708 (N_8708,N_8289,N_8116);
and U8709 (N_8709,N_8155,N_8332);
or U8710 (N_8710,N_8409,N_8338);
xnor U8711 (N_8711,N_8015,N_8129);
nand U8712 (N_8712,N_8375,N_8383);
and U8713 (N_8713,N_8448,N_8325);
or U8714 (N_8714,N_8277,N_8368);
nand U8715 (N_8715,N_8358,N_8408);
or U8716 (N_8716,N_8239,N_8475);
nor U8717 (N_8717,N_8151,N_8340);
and U8718 (N_8718,N_8084,N_8291);
and U8719 (N_8719,N_8174,N_8396);
or U8720 (N_8720,N_8062,N_8423);
or U8721 (N_8721,N_8416,N_8262);
and U8722 (N_8722,N_8493,N_8290);
xnor U8723 (N_8723,N_8008,N_8302);
and U8724 (N_8724,N_8181,N_8199);
and U8725 (N_8725,N_8057,N_8400);
or U8726 (N_8726,N_8436,N_8444);
xnor U8727 (N_8727,N_8212,N_8275);
nor U8728 (N_8728,N_8127,N_8183);
xnor U8729 (N_8729,N_8141,N_8037);
nand U8730 (N_8730,N_8410,N_8469);
nor U8731 (N_8731,N_8333,N_8323);
nor U8732 (N_8732,N_8270,N_8068);
xor U8733 (N_8733,N_8271,N_8484);
xor U8734 (N_8734,N_8321,N_8042);
nand U8735 (N_8735,N_8159,N_8017);
nand U8736 (N_8736,N_8367,N_8481);
xnor U8737 (N_8737,N_8463,N_8120);
nand U8738 (N_8738,N_8253,N_8337);
nor U8739 (N_8739,N_8427,N_8092);
or U8740 (N_8740,N_8029,N_8115);
nand U8741 (N_8741,N_8221,N_8303);
nor U8742 (N_8742,N_8269,N_8148);
or U8743 (N_8743,N_8407,N_8300);
nor U8744 (N_8744,N_8439,N_8216);
nand U8745 (N_8745,N_8497,N_8073);
nor U8746 (N_8746,N_8301,N_8167);
and U8747 (N_8747,N_8334,N_8128);
and U8748 (N_8748,N_8012,N_8236);
xor U8749 (N_8749,N_8459,N_8094);
xnor U8750 (N_8750,N_8422,N_8499);
or U8751 (N_8751,N_8294,N_8056);
nand U8752 (N_8752,N_8275,N_8043);
xor U8753 (N_8753,N_8149,N_8162);
or U8754 (N_8754,N_8291,N_8413);
or U8755 (N_8755,N_8450,N_8299);
nor U8756 (N_8756,N_8202,N_8188);
nand U8757 (N_8757,N_8464,N_8399);
nor U8758 (N_8758,N_8199,N_8464);
nand U8759 (N_8759,N_8046,N_8015);
xnor U8760 (N_8760,N_8257,N_8392);
nand U8761 (N_8761,N_8215,N_8447);
nand U8762 (N_8762,N_8211,N_8180);
xnor U8763 (N_8763,N_8480,N_8029);
nand U8764 (N_8764,N_8001,N_8284);
xnor U8765 (N_8765,N_8380,N_8178);
xnor U8766 (N_8766,N_8103,N_8270);
or U8767 (N_8767,N_8001,N_8202);
nand U8768 (N_8768,N_8151,N_8026);
nand U8769 (N_8769,N_8091,N_8157);
xnor U8770 (N_8770,N_8388,N_8242);
and U8771 (N_8771,N_8408,N_8050);
nand U8772 (N_8772,N_8122,N_8307);
nor U8773 (N_8773,N_8140,N_8451);
and U8774 (N_8774,N_8240,N_8198);
xor U8775 (N_8775,N_8424,N_8135);
xnor U8776 (N_8776,N_8137,N_8440);
or U8777 (N_8777,N_8388,N_8114);
nor U8778 (N_8778,N_8207,N_8357);
or U8779 (N_8779,N_8143,N_8237);
nor U8780 (N_8780,N_8239,N_8169);
nand U8781 (N_8781,N_8447,N_8465);
nand U8782 (N_8782,N_8497,N_8105);
xnor U8783 (N_8783,N_8007,N_8424);
or U8784 (N_8784,N_8416,N_8351);
and U8785 (N_8785,N_8459,N_8052);
and U8786 (N_8786,N_8011,N_8387);
or U8787 (N_8787,N_8190,N_8442);
or U8788 (N_8788,N_8090,N_8363);
nand U8789 (N_8789,N_8330,N_8216);
nor U8790 (N_8790,N_8352,N_8217);
xnor U8791 (N_8791,N_8030,N_8398);
or U8792 (N_8792,N_8301,N_8020);
nor U8793 (N_8793,N_8073,N_8243);
xnor U8794 (N_8794,N_8416,N_8428);
xor U8795 (N_8795,N_8007,N_8289);
or U8796 (N_8796,N_8363,N_8165);
xor U8797 (N_8797,N_8457,N_8192);
nand U8798 (N_8798,N_8023,N_8463);
and U8799 (N_8799,N_8098,N_8312);
and U8800 (N_8800,N_8050,N_8479);
or U8801 (N_8801,N_8439,N_8056);
nor U8802 (N_8802,N_8210,N_8021);
or U8803 (N_8803,N_8086,N_8247);
xnor U8804 (N_8804,N_8227,N_8326);
and U8805 (N_8805,N_8312,N_8067);
and U8806 (N_8806,N_8224,N_8200);
nand U8807 (N_8807,N_8164,N_8173);
xnor U8808 (N_8808,N_8474,N_8254);
or U8809 (N_8809,N_8146,N_8014);
or U8810 (N_8810,N_8098,N_8413);
or U8811 (N_8811,N_8014,N_8482);
nor U8812 (N_8812,N_8229,N_8351);
nor U8813 (N_8813,N_8244,N_8143);
nor U8814 (N_8814,N_8270,N_8416);
and U8815 (N_8815,N_8401,N_8264);
xor U8816 (N_8816,N_8434,N_8345);
xnor U8817 (N_8817,N_8370,N_8124);
and U8818 (N_8818,N_8127,N_8334);
nor U8819 (N_8819,N_8104,N_8318);
xor U8820 (N_8820,N_8370,N_8420);
or U8821 (N_8821,N_8251,N_8482);
or U8822 (N_8822,N_8284,N_8088);
xnor U8823 (N_8823,N_8058,N_8237);
nor U8824 (N_8824,N_8010,N_8193);
nand U8825 (N_8825,N_8475,N_8099);
or U8826 (N_8826,N_8092,N_8079);
xnor U8827 (N_8827,N_8118,N_8489);
xor U8828 (N_8828,N_8407,N_8030);
nand U8829 (N_8829,N_8121,N_8381);
or U8830 (N_8830,N_8423,N_8034);
nand U8831 (N_8831,N_8404,N_8313);
nand U8832 (N_8832,N_8460,N_8385);
xnor U8833 (N_8833,N_8498,N_8087);
nor U8834 (N_8834,N_8195,N_8394);
xnor U8835 (N_8835,N_8173,N_8422);
nand U8836 (N_8836,N_8392,N_8414);
nand U8837 (N_8837,N_8188,N_8019);
xor U8838 (N_8838,N_8007,N_8461);
nand U8839 (N_8839,N_8078,N_8380);
or U8840 (N_8840,N_8218,N_8454);
nand U8841 (N_8841,N_8491,N_8465);
or U8842 (N_8842,N_8314,N_8333);
nor U8843 (N_8843,N_8014,N_8273);
nand U8844 (N_8844,N_8086,N_8495);
nand U8845 (N_8845,N_8072,N_8226);
nor U8846 (N_8846,N_8408,N_8381);
nand U8847 (N_8847,N_8036,N_8087);
nor U8848 (N_8848,N_8180,N_8016);
and U8849 (N_8849,N_8095,N_8224);
nand U8850 (N_8850,N_8478,N_8112);
and U8851 (N_8851,N_8386,N_8398);
or U8852 (N_8852,N_8329,N_8031);
xnor U8853 (N_8853,N_8181,N_8285);
nand U8854 (N_8854,N_8346,N_8452);
xor U8855 (N_8855,N_8051,N_8392);
nand U8856 (N_8856,N_8496,N_8177);
xor U8857 (N_8857,N_8150,N_8232);
or U8858 (N_8858,N_8174,N_8401);
or U8859 (N_8859,N_8141,N_8333);
nor U8860 (N_8860,N_8005,N_8243);
nor U8861 (N_8861,N_8036,N_8335);
xnor U8862 (N_8862,N_8312,N_8418);
or U8863 (N_8863,N_8148,N_8233);
nand U8864 (N_8864,N_8008,N_8257);
or U8865 (N_8865,N_8151,N_8353);
xnor U8866 (N_8866,N_8120,N_8390);
xor U8867 (N_8867,N_8470,N_8412);
and U8868 (N_8868,N_8395,N_8180);
or U8869 (N_8869,N_8125,N_8414);
and U8870 (N_8870,N_8219,N_8449);
nand U8871 (N_8871,N_8033,N_8150);
xor U8872 (N_8872,N_8264,N_8343);
xor U8873 (N_8873,N_8432,N_8240);
nor U8874 (N_8874,N_8282,N_8027);
xor U8875 (N_8875,N_8041,N_8260);
and U8876 (N_8876,N_8151,N_8265);
nand U8877 (N_8877,N_8413,N_8492);
or U8878 (N_8878,N_8004,N_8126);
xor U8879 (N_8879,N_8054,N_8143);
or U8880 (N_8880,N_8420,N_8023);
xor U8881 (N_8881,N_8347,N_8291);
nor U8882 (N_8882,N_8357,N_8090);
xor U8883 (N_8883,N_8198,N_8245);
nor U8884 (N_8884,N_8170,N_8461);
or U8885 (N_8885,N_8042,N_8225);
xor U8886 (N_8886,N_8197,N_8471);
or U8887 (N_8887,N_8137,N_8206);
nand U8888 (N_8888,N_8433,N_8049);
nand U8889 (N_8889,N_8413,N_8197);
nand U8890 (N_8890,N_8290,N_8096);
and U8891 (N_8891,N_8018,N_8405);
nor U8892 (N_8892,N_8263,N_8318);
nand U8893 (N_8893,N_8449,N_8019);
or U8894 (N_8894,N_8148,N_8150);
nand U8895 (N_8895,N_8219,N_8462);
xnor U8896 (N_8896,N_8268,N_8219);
nor U8897 (N_8897,N_8021,N_8064);
nor U8898 (N_8898,N_8179,N_8321);
nand U8899 (N_8899,N_8073,N_8317);
nor U8900 (N_8900,N_8423,N_8015);
or U8901 (N_8901,N_8227,N_8283);
and U8902 (N_8902,N_8065,N_8090);
xor U8903 (N_8903,N_8471,N_8025);
and U8904 (N_8904,N_8017,N_8037);
nand U8905 (N_8905,N_8225,N_8469);
xor U8906 (N_8906,N_8106,N_8312);
or U8907 (N_8907,N_8301,N_8329);
or U8908 (N_8908,N_8157,N_8385);
and U8909 (N_8909,N_8329,N_8078);
xor U8910 (N_8910,N_8095,N_8248);
xor U8911 (N_8911,N_8297,N_8435);
nand U8912 (N_8912,N_8201,N_8366);
nor U8913 (N_8913,N_8092,N_8011);
or U8914 (N_8914,N_8479,N_8303);
xor U8915 (N_8915,N_8082,N_8166);
or U8916 (N_8916,N_8118,N_8355);
nor U8917 (N_8917,N_8490,N_8099);
nand U8918 (N_8918,N_8295,N_8435);
or U8919 (N_8919,N_8393,N_8191);
nand U8920 (N_8920,N_8496,N_8110);
nor U8921 (N_8921,N_8045,N_8275);
nor U8922 (N_8922,N_8411,N_8083);
nor U8923 (N_8923,N_8293,N_8230);
and U8924 (N_8924,N_8166,N_8449);
xnor U8925 (N_8925,N_8458,N_8462);
and U8926 (N_8926,N_8385,N_8474);
nor U8927 (N_8927,N_8446,N_8399);
nand U8928 (N_8928,N_8025,N_8237);
and U8929 (N_8929,N_8337,N_8308);
or U8930 (N_8930,N_8150,N_8402);
nand U8931 (N_8931,N_8203,N_8369);
or U8932 (N_8932,N_8096,N_8185);
or U8933 (N_8933,N_8190,N_8103);
or U8934 (N_8934,N_8147,N_8230);
and U8935 (N_8935,N_8434,N_8083);
nand U8936 (N_8936,N_8357,N_8398);
nand U8937 (N_8937,N_8233,N_8005);
xnor U8938 (N_8938,N_8412,N_8024);
nor U8939 (N_8939,N_8067,N_8402);
or U8940 (N_8940,N_8393,N_8025);
and U8941 (N_8941,N_8249,N_8136);
and U8942 (N_8942,N_8353,N_8264);
xor U8943 (N_8943,N_8466,N_8136);
and U8944 (N_8944,N_8045,N_8120);
or U8945 (N_8945,N_8065,N_8469);
xnor U8946 (N_8946,N_8095,N_8478);
xor U8947 (N_8947,N_8000,N_8279);
xor U8948 (N_8948,N_8069,N_8250);
and U8949 (N_8949,N_8166,N_8253);
nor U8950 (N_8950,N_8302,N_8409);
nand U8951 (N_8951,N_8157,N_8013);
nor U8952 (N_8952,N_8347,N_8010);
and U8953 (N_8953,N_8186,N_8250);
nor U8954 (N_8954,N_8265,N_8277);
xor U8955 (N_8955,N_8182,N_8220);
and U8956 (N_8956,N_8292,N_8427);
or U8957 (N_8957,N_8193,N_8173);
xnor U8958 (N_8958,N_8306,N_8315);
nand U8959 (N_8959,N_8295,N_8242);
xor U8960 (N_8960,N_8378,N_8226);
xnor U8961 (N_8961,N_8309,N_8154);
or U8962 (N_8962,N_8103,N_8433);
or U8963 (N_8963,N_8211,N_8214);
or U8964 (N_8964,N_8363,N_8171);
or U8965 (N_8965,N_8311,N_8084);
nor U8966 (N_8966,N_8225,N_8115);
nor U8967 (N_8967,N_8022,N_8085);
nor U8968 (N_8968,N_8161,N_8387);
xnor U8969 (N_8969,N_8186,N_8413);
nor U8970 (N_8970,N_8499,N_8347);
or U8971 (N_8971,N_8444,N_8443);
nand U8972 (N_8972,N_8189,N_8022);
xnor U8973 (N_8973,N_8356,N_8199);
xor U8974 (N_8974,N_8439,N_8493);
and U8975 (N_8975,N_8020,N_8003);
and U8976 (N_8976,N_8339,N_8267);
nor U8977 (N_8977,N_8335,N_8278);
and U8978 (N_8978,N_8072,N_8076);
xnor U8979 (N_8979,N_8086,N_8164);
xnor U8980 (N_8980,N_8161,N_8470);
or U8981 (N_8981,N_8403,N_8320);
or U8982 (N_8982,N_8143,N_8279);
nand U8983 (N_8983,N_8088,N_8413);
or U8984 (N_8984,N_8181,N_8064);
and U8985 (N_8985,N_8273,N_8452);
xor U8986 (N_8986,N_8196,N_8404);
nand U8987 (N_8987,N_8087,N_8434);
or U8988 (N_8988,N_8426,N_8345);
or U8989 (N_8989,N_8478,N_8326);
xnor U8990 (N_8990,N_8160,N_8188);
and U8991 (N_8991,N_8191,N_8481);
nor U8992 (N_8992,N_8055,N_8316);
and U8993 (N_8993,N_8422,N_8431);
nand U8994 (N_8994,N_8284,N_8378);
nor U8995 (N_8995,N_8074,N_8290);
nor U8996 (N_8996,N_8105,N_8422);
nor U8997 (N_8997,N_8071,N_8382);
and U8998 (N_8998,N_8075,N_8247);
xnor U8999 (N_8999,N_8419,N_8306);
xnor U9000 (N_9000,N_8632,N_8732);
and U9001 (N_9001,N_8568,N_8612);
or U9002 (N_9002,N_8955,N_8771);
xnor U9003 (N_9003,N_8969,N_8639);
nor U9004 (N_9004,N_8640,N_8703);
nand U9005 (N_9005,N_8839,N_8963);
nand U9006 (N_9006,N_8546,N_8702);
and U9007 (N_9007,N_8528,N_8823);
xnor U9008 (N_9008,N_8717,N_8502);
xor U9009 (N_9009,N_8781,N_8956);
nor U9010 (N_9010,N_8851,N_8872);
nand U9011 (N_9011,N_8886,N_8641);
xnor U9012 (N_9012,N_8626,N_8980);
or U9013 (N_9013,N_8767,N_8898);
nor U9014 (N_9014,N_8929,N_8930);
or U9015 (N_9015,N_8696,N_8993);
nand U9016 (N_9016,N_8710,N_8936);
nor U9017 (N_9017,N_8619,N_8654);
or U9018 (N_9018,N_8725,N_8551);
nor U9019 (N_9019,N_8585,N_8916);
nand U9020 (N_9020,N_8997,N_8665);
and U9021 (N_9021,N_8713,N_8706);
nor U9022 (N_9022,N_8743,N_8874);
nand U9023 (N_9023,N_8704,N_8514);
and U9024 (N_9024,N_8797,N_8727);
xor U9025 (N_9025,N_8854,N_8842);
or U9026 (N_9026,N_8584,N_8790);
and U9027 (N_9027,N_8804,N_8628);
xor U9028 (N_9028,N_8720,N_8596);
and U9029 (N_9029,N_8660,N_8622);
xor U9030 (N_9030,N_8992,N_8763);
nand U9031 (N_9031,N_8788,N_8933);
and U9032 (N_9032,N_8850,N_8981);
nor U9033 (N_9033,N_8540,N_8574);
xor U9034 (N_9034,N_8545,N_8547);
xnor U9035 (N_9035,N_8554,N_8719);
nand U9036 (N_9036,N_8723,N_8533);
xor U9037 (N_9037,N_8739,N_8906);
nand U9038 (N_9038,N_8867,N_8532);
nand U9039 (N_9039,N_8796,N_8896);
nor U9040 (N_9040,N_8889,N_8650);
nor U9041 (N_9041,N_8515,N_8937);
and U9042 (N_9042,N_8964,N_8844);
nor U9043 (N_9043,N_8620,N_8864);
and U9044 (N_9044,N_8976,N_8926);
or U9045 (N_9045,N_8892,N_8536);
xor U9046 (N_9046,N_8543,N_8559);
nor U9047 (N_9047,N_8931,N_8870);
nor U9048 (N_9048,N_8830,N_8700);
and U9049 (N_9049,N_8847,N_8592);
xnor U9050 (N_9050,N_8738,N_8808);
or U9051 (N_9051,N_8576,N_8670);
nor U9052 (N_9052,N_8748,N_8950);
nand U9053 (N_9053,N_8637,N_8920);
xnor U9054 (N_9054,N_8942,N_8667);
and U9055 (N_9055,N_8778,N_8745);
nor U9056 (N_9056,N_8875,N_8954);
nand U9057 (N_9057,N_8671,N_8908);
nor U9058 (N_9058,N_8734,N_8986);
xor U9059 (N_9059,N_8856,N_8770);
or U9060 (N_9060,N_8960,N_8567);
nor U9061 (N_9061,N_8646,N_8834);
nor U9062 (N_9062,N_8691,N_8918);
nor U9063 (N_9063,N_8518,N_8746);
and U9064 (N_9064,N_8812,N_8761);
nand U9065 (N_9065,N_8973,N_8894);
nand U9066 (N_9066,N_8901,N_8837);
and U9067 (N_9067,N_8541,N_8990);
nand U9068 (N_9068,N_8962,N_8582);
or U9069 (N_9069,N_8765,N_8983);
nand U9070 (N_9070,N_8625,N_8694);
and U9071 (N_9071,N_8932,N_8643);
nand U9072 (N_9072,N_8644,N_8633);
nand U9073 (N_9073,N_8750,N_8838);
nand U9074 (N_9074,N_8747,N_8594);
and U9075 (N_9075,N_8740,N_8511);
xnor U9076 (N_9076,N_8614,N_8831);
nor U9077 (N_9077,N_8523,N_8708);
nand U9078 (N_9078,N_8814,N_8751);
and U9079 (N_9079,N_8940,N_8501);
xor U9080 (N_9080,N_8583,N_8537);
nand U9081 (N_9081,N_8853,N_8510);
nor U9082 (N_9082,N_8590,N_8873);
and U9083 (N_9083,N_8773,N_8601);
and U9084 (N_9084,N_8946,N_8705);
and U9085 (N_9085,N_8552,N_8564);
nand U9086 (N_9086,N_8688,N_8542);
nand U9087 (N_9087,N_8709,N_8909);
and U9088 (N_9088,N_8604,N_8925);
nand U9089 (N_9089,N_8645,N_8549);
nand U9090 (N_9090,N_8818,N_8826);
xnor U9091 (N_9091,N_8887,N_8504);
or U9092 (N_9092,N_8791,N_8520);
xnor U9093 (N_9093,N_8698,N_8726);
nor U9094 (N_9094,N_8967,N_8524);
nand U9095 (N_9095,N_8935,N_8664);
and U9096 (N_9096,N_8681,N_8807);
nand U9097 (N_9097,N_8675,N_8952);
xor U9098 (N_9098,N_8764,N_8957);
and U9099 (N_9099,N_8958,N_8975);
nor U9100 (N_9100,N_8548,N_8599);
or U9101 (N_9101,N_8924,N_8938);
and U9102 (N_9102,N_8652,N_8903);
nor U9103 (N_9103,N_8662,N_8939);
xnor U9104 (N_9104,N_8752,N_8813);
or U9105 (N_9105,N_8859,N_8657);
or U9106 (N_9106,N_8538,N_8849);
nor U9107 (N_9107,N_8597,N_8701);
xnor U9108 (N_9108,N_8985,N_8737);
or U9109 (N_9109,N_8655,N_8827);
xnor U9110 (N_9110,N_8911,N_8840);
and U9111 (N_9111,N_8769,N_8885);
nand U9112 (N_9112,N_8776,N_8522);
nor U9113 (N_9113,N_8890,N_8786);
and U9114 (N_9114,N_8679,N_8825);
or U9115 (N_9115,N_8998,N_8507);
and U9116 (N_9116,N_8759,N_8697);
and U9117 (N_9117,N_8577,N_8971);
xnor U9118 (N_9118,N_8782,N_8621);
and U9119 (N_9119,N_8672,N_8736);
nor U9120 (N_9120,N_8863,N_8616);
nor U9121 (N_9121,N_8907,N_8815);
or U9122 (N_9122,N_8729,N_8692);
nand U9123 (N_9123,N_8772,N_8517);
nand U9124 (N_9124,N_8603,N_8566);
and U9125 (N_9125,N_8579,N_8755);
nor U9126 (N_9126,N_8774,N_8902);
nand U9127 (N_9127,N_8521,N_8999);
nand U9128 (N_9128,N_8730,N_8915);
or U9129 (N_9129,N_8984,N_8819);
or U9130 (N_9130,N_8500,N_8780);
nor U9131 (N_9131,N_8891,N_8754);
nor U9132 (N_9132,N_8580,N_8927);
and U9133 (N_9133,N_8731,N_8715);
nand U9134 (N_9134,N_8631,N_8760);
or U9135 (N_9135,N_8888,N_8712);
nand U9136 (N_9136,N_8558,N_8525);
xor U9137 (N_9137,N_8508,N_8968);
xnor U9138 (N_9138,N_8795,N_8811);
nor U9139 (N_9139,N_8647,N_8615);
xnor U9140 (N_9140,N_8724,N_8635);
nand U9141 (N_9141,N_8591,N_8919);
xnor U9142 (N_9142,N_8868,N_8741);
nand U9143 (N_9143,N_8570,N_8677);
nand U9144 (N_9144,N_8959,N_8663);
or U9145 (N_9145,N_8505,N_8733);
and U9146 (N_9146,N_8996,N_8693);
xor U9147 (N_9147,N_8882,N_8821);
or U9148 (N_9148,N_8792,N_8953);
and U9149 (N_9149,N_8910,N_8995);
and U9150 (N_9150,N_8608,N_8846);
nor U9151 (N_9151,N_8714,N_8602);
and U9152 (N_9152,N_8707,N_8895);
xnor U9153 (N_9153,N_8649,N_8877);
or U9154 (N_9154,N_8744,N_8600);
xnor U9155 (N_9155,N_8575,N_8832);
nor U9156 (N_9156,N_8685,N_8735);
nand U9157 (N_9157,N_8913,N_8562);
and U9158 (N_9158,N_8800,N_8648);
nor U9159 (N_9159,N_8988,N_8711);
nand U9160 (N_9160,N_8923,N_8561);
xor U9161 (N_9161,N_8878,N_8991);
or U9162 (N_9162,N_8573,N_8829);
nand U9163 (N_9163,N_8972,N_8607);
nor U9164 (N_9164,N_8512,N_8673);
or U9165 (N_9165,N_8506,N_8810);
nand U9166 (N_9166,N_8539,N_8948);
nand U9167 (N_9167,N_8636,N_8678);
xor U9168 (N_9168,N_8684,N_8861);
or U9169 (N_9169,N_8572,N_8722);
nor U9170 (N_9170,N_8793,N_8535);
or U9171 (N_9171,N_8529,N_8917);
and U9172 (N_9172,N_8852,N_8605);
nand U9173 (N_9173,N_8634,N_8556);
nand U9174 (N_9174,N_8593,N_8966);
xor U9175 (N_9175,N_8928,N_8978);
nand U9176 (N_9176,N_8860,N_8669);
or U9177 (N_9177,N_8799,N_8588);
xor U9178 (N_9178,N_8947,N_8526);
and U9179 (N_9179,N_8893,N_8982);
or U9180 (N_9180,N_8941,N_8961);
nand U9181 (N_9181,N_8563,N_8519);
and U9182 (N_9182,N_8695,N_8809);
xor U9183 (N_9183,N_8527,N_8845);
or U9184 (N_9184,N_8784,N_8656);
xnor U9185 (N_9185,N_8611,N_8618);
and U9186 (N_9186,N_8912,N_8905);
nor U9187 (N_9187,N_8989,N_8638);
xnor U9188 (N_9188,N_8749,N_8965);
nor U9189 (N_9189,N_8945,N_8803);
nand U9190 (N_9190,N_8560,N_8550);
or U9191 (N_9191,N_8798,N_8659);
xnor U9192 (N_9192,N_8943,N_8897);
xnor U9193 (N_9193,N_8627,N_8865);
or U9194 (N_9194,N_8802,N_8879);
nor U9195 (N_9195,N_8630,N_8820);
nand U9196 (N_9196,N_8589,N_8974);
or U9197 (N_9197,N_8758,N_8753);
and U9198 (N_9198,N_8794,N_8822);
xnor U9199 (N_9199,N_8987,N_8686);
and U9200 (N_9200,N_8555,N_8553);
or U9201 (N_9201,N_8816,N_8949);
or U9202 (N_9202,N_8516,N_8848);
xor U9203 (N_9203,N_8742,N_8801);
xnor U9204 (N_9204,N_8690,N_8951);
or U9205 (N_9205,N_8833,N_8858);
or U9206 (N_9206,N_8674,N_8544);
and U9207 (N_9207,N_8862,N_8586);
xnor U9208 (N_9208,N_8721,N_8728);
or U9209 (N_9209,N_8768,N_8689);
nand U9210 (N_9210,N_8922,N_8606);
or U9211 (N_9211,N_8977,N_8530);
and U9212 (N_9212,N_8871,N_8789);
or U9213 (N_9213,N_8653,N_8914);
nand U9214 (N_9214,N_8970,N_8531);
and U9215 (N_9215,N_8699,N_8757);
or U9216 (N_9216,N_8824,N_8718);
or U9217 (N_9217,N_8869,N_8835);
xnor U9218 (N_9218,N_8880,N_8766);
or U9219 (N_9219,N_8876,N_8651);
nor U9220 (N_9220,N_8623,N_8534);
and U9221 (N_9221,N_8944,N_8569);
xor U9222 (N_9222,N_8883,N_8884);
or U9223 (N_9223,N_8785,N_8881);
nand U9224 (N_9224,N_8843,N_8610);
xor U9225 (N_9225,N_8609,N_8775);
or U9226 (N_9226,N_8777,N_8666);
or U9227 (N_9227,N_8817,N_8994);
or U9228 (N_9228,N_8828,N_8503);
nand U9229 (N_9229,N_8598,N_8783);
xor U9230 (N_9230,N_8578,N_8934);
and U9231 (N_9231,N_8565,N_8904);
or U9232 (N_9232,N_8787,N_8899);
nand U9233 (N_9233,N_8624,N_8682);
and U9234 (N_9234,N_8629,N_8658);
and U9235 (N_9235,N_8642,N_8841);
nand U9236 (N_9236,N_8668,N_8687);
nor U9237 (N_9237,N_8836,N_8680);
or U9238 (N_9238,N_8571,N_8587);
xnor U9239 (N_9239,N_8762,N_8806);
nand U9240 (N_9240,N_8716,N_8513);
nand U9241 (N_9241,N_8676,N_8613);
nor U9242 (N_9242,N_8509,N_8557);
nand U9243 (N_9243,N_8866,N_8805);
nand U9244 (N_9244,N_8979,N_8617);
nand U9245 (N_9245,N_8921,N_8595);
and U9246 (N_9246,N_8683,N_8756);
nand U9247 (N_9247,N_8779,N_8855);
nand U9248 (N_9248,N_8661,N_8900);
and U9249 (N_9249,N_8581,N_8857);
and U9250 (N_9250,N_8971,N_8780);
or U9251 (N_9251,N_8534,N_8951);
or U9252 (N_9252,N_8712,N_8819);
xor U9253 (N_9253,N_8619,N_8873);
nand U9254 (N_9254,N_8730,N_8529);
xnor U9255 (N_9255,N_8755,N_8853);
nor U9256 (N_9256,N_8524,N_8759);
or U9257 (N_9257,N_8583,N_8835);
nand U9258 (N_9258,N_8650,N_8934);
xnor U9259 (N_9259,N_8633,N_8528);
xnor U9260 (N_9260,N_8917,N_8701);
nor U9261 (N_9261,N_8908,N_8955);
or U9262 (N_9262,N_8995,N_8875);
and U9263 (N_9263,N_8781,N_8919);
nor U9264 (N_9264,N_8688,N_8640);
xor U9265 (N_9265,N_8700,N_8969);
nor U9266 (N_9266,N_8802,N_8743);
nor U9267 (N_9267,N_8588,N_8642);
or U9268 (N_9268,N_8966,N_8983);
and U9269 (N_9269,N_8635,N_8581);
xor U9270 (N_9270,N_8596,N_8978);
xnor U9271 (N_9271,N_8876,N_8506);
nor U9272 (N_9272,N_8517,N_8815);
xnor U9273 (N_9273,N_8673,N_8664);
and U9274 (N_9274,N_8590,N_8958);
xnor U9275 (N_9275,N_8611,N_8870);
xor U9276 (N_9276,N_8962,N_8623);
nor U9277 (N_9277,N_8790,N_8736);
nand U9278 (N_9278,N_8764,N_8634);
or U9279 (N_9279,N_8864,N_8853);
or U9280 (N_9280,N_8776,N_8819);
nand U9281 (N_9281,N_8539,N_8992);
nand U9282 (N_9282,N_8960,N_8644);
nand U9283 (N_9283,N_8669,N_8869);
nand U9284 (N_9284,N_8658,N_8548);
or U9285 (N_9285,N_8867,N_8921);
or U9286 (N_9286,N_8782,N_8870);
nand U9287 (N_9287,N_8613,N_8822);
and U9288 (N_9288,N_8987,N_8604);
nand U9289 (N_9289,N_8584,N_8590);
or U9290 (N_9290,N_8684,N_8555);
nor U9291 (N_9291,N_8781,N_8501);
xnor U9292 (N_9292,N_8906,N_8763);
and U9293 (N_9293,N_8911,N_8950);
xor U9294 (N_9294,N_8966,N_8714);
and U9295 (N_9295,N_8733,N_8936);
xnor U9296 (N_9296,N_8892,N_8563);
or U9297 (N_9297,N_8789,N_8907);
or U9298 (N_9298,N_8967,N_8755);
nor U9299 (N_9299,N_8783,N_8796);
and U9300 (N_9300,N_8513,N_8673);
and U9301 (N_9301,N_8864,N_8881);
nand U9302 (N_9302,N_8788,N_8766);
or U9303 (N_9303,N_8705,N_8978);
and U9304 (N_9304,N_8740,N_8897);
nor U9305 (N_9305,N_8500,N_8504);
nor U9306 (N_9306,N_8940,N_8527);
xnor U9307 (N_9307,N_8512,N_8892);
xnor U9308 (N_9308,N_8772,N_8803);
xnor U9309 (N_9309,N_8848,N_8947);
and U9310 (N_9310,N_8977,N_8763);
and U9311 (N_9311,N_8545,N_8879);
xor U9312 (N_9312,N_8872,N_8758);
xor U9313 (N_9313,N_8518,N_8684);
nand U9314 (N_9314,N_8715,N_8868);
nor U9315 (N_9315,N_8914,N_8956);
nand U9316 (N_9316,N_8525,N_8533);
nand U9317 (N_9317,N_8905,N_8920);
nand U9318 (N_9318,N_8772,N_8773);
and U9319 (N_9319,N_8906,N_8857);
or U9320 (N_9320,N_8727,N_8722);
xnor U9321 (N_9321,N_8750,N_8854);
and U9322 (N_9322,N_8505,N_8749);
xor U9323 (N_9323,N_8546,N_8864);
or U9324 (N_9324,N_8926,N_8647);
nor U9325 (N_9325,N_8507,N_8844);
xnor U9326 (N_9326,N_8876,N_8546);
and U9327 (N_9327,N_8620,N_8947);
nor U9328 (N_9328,N_8627,N_8874);
or U9329 (N_9329,N_8965,N_8708);
nor U9330 (N_9330,N_8978,N_8846);
or U9331 (N_9331,N_8635,N_8691);
nor U9332 (N_9332,N_8668,N_8561);
and U9333 (N_9333,N_8976,N_8663);
or U9334 (N_9334,N_8701,N_8918);
or U9335 (N_9335,N_8598,N_8677);
xnor U9336 (N_9336,N_8853,N_8845);
and U9337 (N_9337,N_8650,N_8611);
xor U9338 (N_9338,N_8988,N_8535);
nor U9339 (N_9339,N_8879,N_8976);
or U9340 (N_9340,N_8735,N_8918);
nor U9341 (N_9341,N_8790,N_8925);
xnor U9342 (N_9342,N_8968,N_8557);
nor U9343 (N_9343,N_8658,N_8690);
xor U9344 (N_9344,N_8793,N_8986);
or U9345 (N_9345,N_8687,N_8887);
xnor U9346 (N_9346,N_8561,N_8767);
and U9347 (N_9347,N_8742,N_8510);
or U9348 (N_9348,N_8847,N_8797);
nor U9349 (N_9349,N_8666,N_8957);
xnor U9350 (N_9350,N_8913,N_8632);
or U9351 (N_9351,N_8608,N_8636);
or U9352 (N_9352,N_8781,N_8511);
xnor U9353 (N_9353,N_8517,N_8676);
and U9354 (N_9354,N_8826,N_8693);
nor U9355 (N_9355,N_8560,N_8670);
and U9356 (N_9356,N_8844,N_8990);
nand U9357 (N_9357,N_8501,N_8848);
nand U9358 (N_9358,N_8724,N_8544);
nand U9359 (N_9359,N_8661,N_8824);
nand U9360 (N_9360,N_8659,N_8676);
nor U9361 (N_9361,N_8705,N_8654);
xnor U9362 (N_9362,N_8924,N_8558);
or U9363 (N_9363,N_8639,N_8959);
xnor U9364 (N_9364,N_8915,N_8841);
or U9365 (N_9365,N_8798,N_8906);
or U9366 (N_9366,N_8536,N_8711);
and U9367 (N_9367,N_8826,N_8712);
xor U9368 (N_9368,N_8963,N_8795);
nor U9369 (N_9369,N_8586,N_8893);
nand U9370 (N_9370,N_8676,N_8988);
or U9371 (N_9371,N_8513,N_8500);
or U9372 (N_9372,N_8790,N_8640);
nand U9373 (N_9373,N_8824,N_8802);
nand U9374 (N_9374,N_8686,N_8717);
or U9375 (N_9375,N_8652,N_8714);
nor U9376 (N_9376,N_8840,N_8756);
xor U9377 (N_9377,N_8813,N_8896);
xnor U9378 (N_9378,N_8982,N_8547);
nand U9379 (N_9379,N_8781,N_8735);
and U9380 (N_9380,N_8950,N_8973);
xor U9381 (N_9381,N_8866,N_8841);
or U9382 (N_9382,N_8844,N_8982);
or U9383 (N_9383,N_8972,N_8709);
xnor U9384 (N_9384,N_8970,N_8870);
nand U9385 (N_9385,N_8893,N_8761);
or U9386 (N_9386,N_8834,N_8856);
nor U9387 (N_9387,N_8977,N_8903);
nor U9388 (N_9388,N_8859,N_8989);
nand U9389 (N_9389,N_8818,N_8687);
nand U9390 (N_9390,N_8693,N_8677);
nor U9391 (N_9391,N_8575,N_8850);
nor U9392 (N_9392,N_8777,N_8552);
and U9393 (N_9393,N_8676,N_8857);
and U9394 (N_9394,N_8962,N_8678);
and U9395 (N_9395,N_8620,N_8990);
xnor U9396 (N_9396,N_8884,N_8762);
and U9397 (N_9397,N_8671,N_8941);
nand U9398 (N_9398,N_8828,N_8836);
nand U9399 (N_9399,N_8982,N_8631);
nor U9400 (N_9400,N_8874,N_8906);
or U9401 (N_9401,N_8762,N_8721);
and U9402 (N_9402,N_8658,N_8895);
and U9403 (N_9403,N_8736,N_8945);
xor U9404 (N_9404,N_8575,N_8750);
and U9405 (N_9405,N_8844,N_8856);
xor U9406 (N_9406,N_8573,N_8877);
xnor U9407 (N_9407,N_8736,N_8993);
nor U9408 (N_9408,N_8688,N_8575);
or U9409 (N_9409,N_8721,N_8794);
or U9410 (N_9410,N_8595,N_8610);
nor U9411 (N_9411,N_8752,N_8833);
nand U9412 (N_9412,N_8832,N_8680);
nand U9413 (N_9413,N_8590,N_8683);
xnor U9414 (N_9414,N_8717,N_8575);
and U9415 (N_9415,N_8684,N_8689);
and U9416 (N_9416,N_8570,N_8624);
nor U9417 (N_9417,N_8892,N_8997);
and U9418 (N_9418,N_8750,N_8585);
and U9419 (N_9419,N_8596,N_8689);
xor U9420 (N_9420,N_8742,N_8771);
and U9421 (N_9421,N_8508,N_8502);
xnor U9422 (N_9422,N_8648,N_8635);
and U9423 (N_9423,N_8897,N_8813);
nor U9424 (N_9424,N_8682,N_8609);
nor U9425 (N_9425,N_8854,N_8702);
or U9426 (N_9426,N_8948,N_8548);
and U9427 (N_9427,N_8607,N_8708);
and U9428 (N_9428,N_8767,N_8503);
xnor U9429 (N_9429,N_8689,N_8950);
xor U9430 (N_9430,N_8925,N_8887);
and U9431 (N_9431,N_8940,N_8878);
nand U9432 (N_9432,N_8607,N_8587);
xnor U9433 (N_9433,N_8599,N_8684);
nor U9434 (N_9434,N_8762,N_8619);
and U9435 (N_9435,N_8747,N_8842);
nor U9436 (N_9436,N_8892,N_8616);
and U9437 (N_9437,N_8842,N_8906);
nand U9438 (N_9438,N_8958,N_8955);
and U9439 (N_9439,N_8540,N_8558);
nor U9440 (N_9440,N_8500,N_8763);
or U9441 (N_9441,N_8982,N_8976);
nand U9442 (N_9442,N_8854,N_8853);
xnor U9443 (N_9443,N_8712,N_8539);
nor U9444 (N_9444,N_8890,N_8612);
xnor U9445 (N_9445,N_8513,N_8810);
and U9446 (N_9446,N_8735,N_8864);
nor U9447 (N_9447,N_8698,N_8562);
nand U9448 (N_9448,N_8826,N_8822);
and U9449 (N_9449,N_8662,N_8778);
nor U9450 (N_9450,N_8835,N_8748);
and U9451 (N_9451,N_8503,N_8931);
nor U9452 (N_9452,N_8895,N_8553);
xnor U9453 (N_9453,N_8988,N_8968);
nand U9454 (N_9454,N_8859,N_8561);
xor U9455 (N_9455,N_8898,N_8685);
or U9456 (N_9456,N_8674,N_8965);
nor U9457 (N_9457,N_8843,N_8654);
and U9458 (N_9458,N_8995,N_8937);
or U9459 (N_9459,N_8529,N_8994);
and U9460 (N_9460,N_8602,N_8890);
and U9461 (N_9461,N_8939,N_8519);
nand U9462 (N_9462,N_8754,N_8750);
and U9463 (N_9463,N_8953,N_8860);
or U9464 (N_9464,N_8899,N_8573);
nor U9465 (N_9465,N_8656,N_8762);
or U9466 (N_9466,N_8764,N_8967);
nand U9467 (N_9467,N_8631,N_8693);
or U9468 (N_9468,N_8712,N_8752);
or U9469 (N_9469,N_8802,N_8783);
or U9470 (N_9470,N_8686,N_8644);
nand U9471 (N_9471,N_8526,N_8807);
nand U9472 (N_9472,N_8919,N_8883);
and U9473 (N_9473,N_8725,N_8956);
nand U9474 (N_9474,N_8502,N_8709);
nand U9475 (N_9475,N_8912,N_8600);
nor U9476 (N_9476,N_8761,N_8977);
or U9477 (N_9477,N_8654,N_8584);
xor U9478 (N_9478,N_8887,N_8873);
or U9479 (N_9479,N_8711,N_8527);
xnor U9480 (N_9480,N_8857,N_8879);
and U9481 (N_9481,N_8551,N_8623);
nand U9482 (N_9482,N_8883,N_8702);
nor U9483 (N_9483,N_8783,N_8826);
or U9484 (N_9484,N_8886,N_8574);
nand U9485 (N_9485,N_8971,N_8773);
nor U9486 (N_9486,N_8918,N_8720);
xnor U9487 (N_9487,N_8834,N_8517);
or U9488 (N_9488,N_8772,N_8839);
nand U9489 (N_9489,N_8891,N_8834);
and U9490 (N_9490,N_8776,N_8558);
and U9491 (N_9491,N_8836,N_8817);
or U9492 (N_9492,N_8707,N_8607);
or U9493 (N_9493,N_8674,N_8633);
nand U9494 (N_9494,N_8724,N_8888);
nor U9495 (N_9495,N_8603,N_8870);
nor U9496 (N_9496,N_8929,N_8520);
and U9497 (N_9497,N_8874,N_8980);
and U9498 (N_9498,N_8716,N_8956);
and U9499 (N_9499,N_8904,N_8602);
nand U9500 (N_9500,N_9196,N_9138);
nor U9501 (N_9501,N_9272,N_9376);
xnor U9502 (N_9502,N_9336,N_9268);
and U9503 (N_9503,N_9467,N_9393);
nand U9504 (N_9504,N_9029,N_9315);
and U9505 (N_9505,N_9219,N_9195);
and U9506 (N_9506,N_9211,N_9077);
and U9507 (N_9507,N_9079,N_9139);
and U9508 (N_9508,N_9399,N_9004);
and U9509 (N_9509,N_9396,N_9224);
nand U9510 (N_9510,N_9416,N_9206);
or U9511 (N_9511,N_9190,N_9075);
and U9512 (N_9512,N_9185,N_9241);
xnor U9513 (N_9513,N_9250,N_9403);
xnor U9514 (N_9514,N_9228,N_9094);
nand U9515 (N_9515,N_9059,N_9063);
nand U9516 (N_9516,N_9323,N_9445);
and U9517 (N_9517,N_9245,N_9027);
nand U9518 (N_9518,N_9036,N_9242);
xor U9519 (N_9519,N_9477,N_9351);
or U9520 (N_9520,N_9115,N_9026);
and U9521 (N_9521,N_9292,N_9400);
or U9522 (N_9522,N_9287,N_9042);
or U9523 (N_9523,N_9488,N_9342);
or U9524 (N_9524,N_9299,N_9105);
nor U9525 (N_9525,N_9343,N_9111);
xnor U9526 (N_9526,N_9289,N_9015);
and U9527 (N_9527,N_9433,N_9064);
or U9528 (N_9528,N_9310,N_9135);
xnor U9529 (N_9529,N_9402,N_9177);
or U9530 (N_9530,N_9198,N_9340);
nand U9531 (N_9531,N_9216,N_9176);
nand U9532 (N_9532,N_9392,N_9204);
or U9533 (N_9533,N_9009,N_9114);
and U9534 (N_9534,N_9005,N_9280);
xnor U9535 (N_9535,N_9309,N_9412);
nand U9536 (N_9536,N_9408,N_9207);
and U9537 (N_9537,N_9189,N_9048);
nand U9538 (N_9538,N_9043,N_9334);
nor U9539 (N_9539,N_9200,N_9083);
and U9540 (N_9540,N_9047,N_9012);
or U9541 (N_9541,N_9007,N_9188);
or U9542 (N_9542,N_9371,N_9273);
xnor U9543 (N_9543,N_9421,N_9499);
nand U9544 (N_9544,N_9161,N_9428);
or U9545 (N_9545,N_9031,N_9441);
xor U9546 (N_9546,N_9203,N_9303);
nor U9547 (N_9547,N_9129,N_9410);
xor U9548 (N_9548,N_9008,N_9264);
or U9549 (N_9549,N_9308,N_9293);
nor U9550 (N_9550,N_9236,N_9167);
nand U9551 (N_9551,N_9178,N_9247);
or U9552 (N_9552,N_9430,N_9277);
nand U9553 (N_9553,N_9013,N_9267);
and U9554 (N_9554,N_9345,N_9102);
nor U9555 (N_9555,N_9084,N_9088);
nand U9556 (N_9556,N_9360,N_9082);
nor U9557 (N_9557,N_9095,N_9490);
nor U9558 (N_9558,N_9150,N_9210);
xnor U9559 (N_9559,N_9076,N_9483);
or U9560 (N_9560,N_9018,N_9482);
nand U9561 (N_9561,N_9122,N_9067);
nand U9562 (N_9562,N_9413,N_9035);
nand U9563 (N_9563,N_9370,N_9327);
nor U9564 (N_9564,N_9163,N_9024);
and U9565 (N_9565,N_9324,N_9225);
nor U9566 (N_9566,N_9325,N_9132);
and U9567 (N_9567,N_9263,N_9186);
nand U9568 (N_9568,N_9212,N_9034);
xor U9569 (N_9569,N_9479,N_9126);
nor U9570 (N_9570,N_9125,N_9385);
nor U9571 (N_9571,N_9422,N_9427);
xor U9572 (N_9572,N_9143,N_9418);
and U9573 (N_9573,N_9113,N_9232);
and U9574 (N_9574,N_9107,N_9357);
xnor U9575 (N_9575,N_9191,N_9246);
xnor U9576 (N_9576,N_9087,N_9470);
and U9577 (N_9577,N_9316,N_9326);
xor U9578 (N_9578,N_9466,N_9174);
nor U9579 (N_9579,N_9202,N_9002);
and U9580 (N_9580,N_9085,N_9497);
nand U9581 (N_9581,N_9223,N_9380);
nand U9582 (N_9582,N_9081,N_9361);
xnor U9583 (N_9583,N_9106,N_9367);
or U9584 (N_9584,N_9305,N_9050);
xnor U9585 (N_9585,N_9220,N_9151);
xnor U9586 (N_9586,N_9213,N_9350);
xnor U9587 (N_9587,N_9030,N_9382);
nand U9588 (N_9588,N_9281,N_9072);
and U9589 (N_9589,N_9182,N_9054);
or U9590 (N_9590,N_9230,N_9259);
xnor U9591 (N_9591,N_9068,N_9239);
or U9592 (N_9592,N_9271,N_9362);
or U9593 (N_9593,N_9374,N_9387);
nand U9594 (N_9594,N_9258,N_9417);
and U9595 (N_9595,N_9158,N_9244);
nand U9596 (N_9596,N_9153,N_9330);
or U9597 (N_9597,N_9217,N_9291);
nand U9598 (N_9598,N_9473,N_9146);
nand U9599 (N_9599,N_9116,N_9295);
nand U9600 (N_9600,N_9450,N_9061);
nor U9601 (N_9601,N_9347,N_9491);
and U9602 (N_9602,N_9180,N_9051);
or U9603 (N_9603,N_9437,N_9498);
or U9604 (N_9604,N_9155,N_9199);
nand U9605 (N_9605,N_9165,N_9468);
nand U9606 (N_9606,N_9233,N_9356);
nand U9607 (N_9607,N_9306,N_9120);
xor U9608 (N_9608,N_9436,N_9016);
nor U9609 (N_9609,N_9251,N_9025);
nor U9610 (N_9610,N_9020,N_9152);
nor U9611 (N_9611,N_9331,N_9112);
xor U9612 (N_9612,N_9156,N_9157);
nand U9613 (N_9613,N_9221,N_9208);
and U9614 (N_9614,N_9071,N_9487);
and U9615 (N_9615,N_9270,N_9010);
and U9616 (N_9616,N_9038,N_9046);
nor U9617 (N_9617,N_9352,N_9425);
or U9618 (N_9618,N_9288,N_9274);
nor U9619 (N_9619,N_9069,N_9240);
xnor U9620 (N_9620,N_9184,N_9290);
xnor U9621 (N_9621,N_9472,N_9283);
nor U9622 (N_9622,N_9160,N_9443);
or U9623 (N_9623,N_9354,N_9006);
nand U9624 (N_9624,N_9108,N_9057);
or U9625 (N_9625,N_9183,N_9368);
nand U9626 (N_9626,N_9379,N_9481);
xnor U9627 (N_9627,N_9044,N_9099);
and U9628 (N_9628,N_9179,N_9296);
nor U9629 (N_9629,N_9276,N_9346);
xor U9630 (N_9630,N_9110,N_9214);
nor U9631 (N_9631,N_9381,N_9091);
nand U9632 (N_9632,N_9017,N_9149);
nand U9633 (N_9633,N_9318,N_9429);
xnor U9634 (N_9634,N_9444,N_9415);
nor U9635 (N_9635,N_9397,N_9121);
and U9636 (N_9636,N_9137,N_9353);
nand U9637 (N_9637,N_9119,N_9260);
nor U9638 (N_9638,N_9307,N_9476);
or U9639 (N_9639,N_9066,N_9058);
nor U9640 (N_9640,N_9278,N_9133);
nor U9641 (N_9641,N_9118,N_9117);
or U9642 (N_9642,N_9448,N_9359);
nand U9643 (N_9643,N_9169,N_9344);
nor U9644 (N_9644,N_9011,N_9222);
and U9645 (N_9645,N_9098,N_9431);
or U9646 (N_9646,N_9124,N_9435);
xnor U9647 (N_9647,N_9432,N_9145);
or U9648 (N_9648,N_9337,N_9140);
and U9649 (N_9649,N_9170,N_9341);
xnor U9650 (N_9650,N_9201,N_9489);
or U9651 (N_9651,N_9453,N_9451);
xnor U9652 (N_9652,N_9405,N_9073);
nor U9653 (N_9653,N_9449,N_9434);
nor U9654 (N_9654,N_9023,N_9363);
nand U9655 (N_9655,N_9197,N_9457);
nor U9656 (N_9656,N_9314,N_9218);
nor U9657 (N_9657,N_9492,N_9089);
and U9658 (N_9658,N_9384,N_9404);
and U9659 (N_9659,N_9227,N_9231);
and U9660 (N_9660,N_9313,N_9053);
nor U9661 (N_9661,N_9109,N_9101);
and U9662 (N_9662,N_9304,N_9423);
nand U9663 (N_9663,N_9456,N_9056);
and U9664 (N_9664,N_9414,N_9266);
nor U9665 (N_9665,N_9333,N_9471);
nand U9666 (N_9666,N_9033,N_9398);
and U9667 (N_9667,N_9144,N_9253);
xnor U9668 (N_9668,N_9328,N_9461);
or U9669 (N_9669,N_9000,N_9100);
xnor U9670 (N_9670,N_9459,N_9238);
xnor U9671 (N_9671,N_9474,N_9485);
nand U9672 (N_9672,N_9041,N_9080);
or U9673 (N_9673,N_9162,N_9424);
and U9674 (N_9674,N_9355,N_9406);
nor U9675 (N_9675,N_9319,N_9104);
and U9676 (N_9676,N_9465,N_9426);
xor U9677 (N_9677,N_9062,N_9142);
or U9678 (N_9678,N_9302,N_9300);
nand U9679 (N_9679,N_9411,N_9123);
nor U9680 (N_9680,N_9021,N_9348);
and U9681 (N_9681,N_9147,N_9248);
nand U9682 (N_9682,N_9173,N_9286);
xnor U9683 (N_9683,N_9494,N_9037);
and U9684 (N_9684,N_9269,N_9065);
and U9685 (N_9685,N_9265,N_9389);
nand U9686 (N_9686,N_9395,N_9373);
nand U9687 (N_9687,N_9294,N_9317);
or U9688 (N_9688,N_9226,N_9475);
or U9689 (N_9689,N_9285,N_9255);
nor U9690 (N_9690,N_9312,N_9455);
or U9691 (N_9691,N_9469,N_9480);
or U9692 (N_9692,N_9349,N_9193);
nand U9693 (N_9693,N_9166,N_9297);
xor U9694 (N_9694,N_9243,N_9298);
nand U9695 (N_9695,N_9366,N_9194);
xnor U9696 (N_9696,N_9172,N_9168);
xnor U9697 (N_9697,N_9128,N_9320);
or U9698 (N_9698,N_9256,N_9181);
nand U9699 (N_9699,N_9358,N_9329);
nand U9700 (N_9700,N_9311,N_9390);
nand U9701 (N_9701,N_9388,N_9339);
or U9702 (N_9702,N_9279,N_9154);
and U9703 (N_9703,N_9159,N_9442);
and U9704 (N_9704,N_9164,N_9321);
nor U9705 (N_9705,N_9103,N_9014);
or U9706 (N_9706,N_9301,N_9493);
nor U9707 (N_9707,N_9086,N_9275);
or U9708 (N_9708,N_9458,N_9141);
or U9709 (N_9709,N_9391,N_9254);
nand U9710 (N_9710,N_9070,N_9028);
or U9711 (N_9711,N_9439,N_9486);
nor U9712 (N_9712,N_9127,N_9192);
or U9713 (N_9713,N_9369,N_9052);
nand U9714 (N_9714,N_9209,N_9401);
or U9715 (N_9715,N_9136,N_9261);
xnor U9716 (N_9716,N_9394,N_9229);
or U9717 (N_9717,N_9175,N_9215);
or U9718 (N_9718,N_9187,N_9032);
nand U9719 (N_9719,N_9205,N_9090);
xnor U9720 (N_9720,N_9484,N_9332);
and U9721 (N_9721,N_9420,N_9235);
xor U9722 (N_9722,N_9252,N_9171);
nor U9723 (N_9723,N_9019,N_9454);
or U9724 (N_9724,N_9234,N_9003);
nor U9725 (N_9725,N_9365,N_9460);
nand U9726 (N_9726,N_9364,N_9134);
xnor U9727 (N_9727,N_9096,N_9040);
or U9728 (N_9728,N_9262,N_9372);
or U9729 (N_9729,N_9447,N_9049);
or U9730 (N_9730,N_9496,N_9375);
xnor U9731 (N_9731,N_9438,N_9092);
and U9732 (N_9732,N_9074,N_9495);
and U9733 (N_9733,N_9464,N_9383);
nor U9734 (N_9734,N_9237,N_9322);
nor U9735 (N_9735,N_9377,N_9335);
xor U9736 (N_9736,N_9478,N_9386);
or U9737 (N_9737,N_9097,N_9452);
xnor U9738 (N_9738,N_9257,N_9078);
nand U9739 (N_9739,N_9440,N_9462);
xnor U9740 (N_9740,N_9148,N_9060);
nor U9741 (N_9741,N_9001,N_9093);
nor U9742 (N_9742,N_9249,N_9409);
xnor U9743 (N_9743,N_9378,N_9130);
nor U9744 (N_9744,N_9055,N_9419);
or U9745 (N_9745,N_9338,N_9407);
and U9746 (N_9746,N_9463,N_9045);
or U9747 (N_9747,N_9284,N_9446);
xor U9748 (N_9748,N_9282,N_9022);
xnor U9749 (N_9749,N_9131,N_9039);
or U9750 (N_9750,N_9364,N_9042);
xor U9751 (N_9751,N_9377,N_9153);
or U9752 (N_9752,N_9359,N_9146);
or U9753 (N_9753,N_9012,N_9095);
xor U9754 (N_9754,N_9238,N_9022);
nand U9755 (N_9755,N_9207,N_9496);
or U9756 (N_9756,N_9116,N_9144);
xnor U9757 (N_9757,N_9174,N_9444);
or U9758 (N_9758,N_9401,N_9340);
and U9759 (N_9759,N_9244,N_9292);
xnor U9760 (N_9760,N_9109,N_9280);
nor U9761 (N_9761,N_9366,N_9212);
nand U9762 (N_9762,N_9390,N_9037);
nor U9763 (N_9763,N_9118,N_9457);
nor U9764 (N_9764,N_9252,N_9424);
and U9765 (N_9765,N_9401,N_9118);
nand U9766 (N_9766,N_9089,N_9391);
nand U9767 (N_9767,N_9164,N_9198);
and U9768 (N_9768,N_9255,N_9228);
and U9769 (N_9769,N_9125,N_9132);
or U9770 (N_9770,N_9274,N_9086);
xnor U9771 (N_9771,N_9335,N_9046);
xnor U9772 (N_9772,N_9214,N_9450);
nand U9773 (N_9773,N_9436,N_9306);
nand U9774 (N_9774,N_9105,N_9168);
or U9775 (N_9775,N_9049,N_9235);
or U9776 (N_9776,N_9336,N_9275);
and U9777 (N_9777,N_9259,N_9422);
and U9778 (N_9778,N_9241,N_9345);
or U9779 (N_9779,N_9161,N_9363);
or U9780 (N_9780,N_9242,N_9048);
and U9781 (N_9781,N_9059,N_9019);
nand U9782 (N_9782,N_9021,N_9462);
and U9783 (N_9783,N_9357,N_9120);
nand U9784 (N_9784,N_9371,N_9296);
or U9785 (N_9785,N_9108,N_9407);
and U9786 (N_9786,N_9481,N_9418);
nand U9787 (N_9787,N_9115,N_9396);
or U9788 (N_9788,N_9309,N_9377);
or U9789 (N_9789,N_9031,N_9483);
and U9790 (N_9790,N_9202,N_9474);
nand U9791 (N_9791,N_9165,N_9441);
nand U9792 (N_9792,N_9148,N_9255);
or U9793 (N_9793,N_9057,N_9065);
nand U9794 (N_9794,N_9137,N_9468);
xnor U9795 (N_9795,N_9428,N_9028);
or U9796 (N_9796,N_9141,N_9029);
xnor U9797 (N_9797,N_9234,N_9166);
nand U9798 (N_9798,N_9152,N_9266);
and U9799 (N_9799,N_9138,N_9224);
xor U9800 (N_9800,N_9002,N_9176);
nand U9801 (N_9801,N_9070,N_9188);
nand U9802 (N_9802,N_9408,N_9388);
and U9803 (N_9803,N_9059,N_9456);
nand U9804 (N_9804,N_9116,N_9049);
nand U9805 (N_9805,N_9334,N_9396);
nand U9806 (N_9806,N_9161,N_9258);
nor U9807 (N_9807,N_9035,N_9161);
nor U9808 (N_9808,N_9350,N_9417);
or U9809 (N_9809,N_9168,N_9466);
xor U9810 (N_9810,N_9450,N_9299);
or U9811 (N_9811,N_9044,N_9346);
nor U9812 (N_9812,N_9252,N_9250);
or U9813 (N_9813,N_9379,N_9436);
and U9814 (N_9814,N_9480,N_9258);
nand U9815 (N_9815,N_9395,N_9306);
xnor U9816 (N_9816,N_9092,N_9301);
and U9817 (N_9817,N_9177,N_9424);
xor U9818 (N_9818,N_9285,N_9478);
xor U9819 (N_9819,N_9441,N_9342);
or U9820 (N_9820,N_9116,N_9124);
or U9821 (N_9821,N_9328,N_9453);
nand U9822 (N_9822,N_9393,N_9080);
nand U9823 (N_9823,N_9289,N_9104);
nor U9824 (N_9824,N_9022,N_9088);
or U9825 (N_9825,N_9189,N_9343);
or U9826 (N_9826,N_9224,N_9191);
nand U9827 (N_9827,N_9279,N_9142);
or U9828 (N_9828,N_9224,N_9373);
nand U9829 (N_9829,N_9339,N_9026);
or U9830 (N_9830,N_9317,N_9492);
xnor U9831 (N_9831,N_9491,N_9160);
and U9832 (N_9832,N_9453,N_9478);
nand U9833 (N_9833,N_9363,N_9198);
nand U9834 (N_9834,N_9125,N_9128);
or U9835 (N_9835,N_9400,N_9359);
nor U9836 (N_9836,N_9313,N_9199);
and U9837 (N_9837,N_9477,N_9236);
and U9838 (N_9838,N_9458,N_9467);
xnor U9839 (N_9839,N_9452,N_9310);
or U9840 (N_9840,N_9379,N_9414);
xnor U9841 (N_9841,N_9222,N_9474);
and U9842 (N_9842,N_9448,N_9343);
nor U9843 (N_9843,N_9141,N_9350);
and U9844 (N_9844,N_9198,N_9234);
xor U9845 (N_9845,N_9132,N_9006);
and U9846 (N_9846,N_9029,N_9443);
or U9847 (N_9847,N_9182,N_9409);
and U9848 (N_9848,N_9140,N_9304);
and U9849 (N_9849,N_9258,N_9026);
nand U9850 (N_9850,N_9184,N_9124);
xor U9851 (N_9851,N_9045,N_9308);
xor U9852 (N_9852,N_9034,N_9340);
nor U9853 (N_9853,N_9449,N_9318);
and U9854 (N_9854,N_9494,N_9493);
or U9855 (N_9855,N_9018,N_9422);
nand U9856 (N_9856,N_9441,N_9015);
and U9857 (N_9857,N_9260,N_9281);
and U9858 (N_9858,N_9292,N_9060);
and U9859 (N_9859,N_9131,N_9092);
nor U9860 (N_9860,N_9429,N_9309);
nor U9861 (N_9861,N_9036,N_9128);
nand U9862 (N_9862,N_9156,N_9235);
nor U9863 (N_9863,N_9404,N_9067);
xnor U9864 (N_9864,N_9380,N_9325);
and U9865 (N_9865,N_9318,N_9372);
or U9866 (N_9866,N_9440,N_9432);
nand U9867 (N_9867,N_9329,N_9005);
and U9868 (N_9868,N_9374,N_9022);
nand U9869 (N_9869,N_9224,N_9253);
or U9870 (N_9870,N_9318,N_9306);
and U9871 (N_9871,N_9409,N_9315);
and U9872 (N_9872,N_9219,N_9015);
nand U9873 (N_9873,N_9329,N_9454);
or U9874 (N_9874,N_9335,N_9379);
and U9875 (N_9875,N_9003,N_9411);
xor U9876 (N_9876,N_9001,N_9320);
xor U9877 (N_9877,N_9008,N_9009);
xor U9878 (N_9878,N_9463,N_9425);
nand U9879 (N_9879,N_9151,N_9233);
nor U9880 (N_9880,N_9063,N_9115);
nor U9881 (N_9881,N_9067,N_9431);
nor U9882 (N_9882,N_9358,N_9149);
nor U9883 (N_9883,N_9177,N_9277);
nor U9884 (N_9884,N_9242,N_9229);
or U9885 (N_9885,N_9288,N_9157);
nor U9886 (N_9886,N_9391,N_9436);
nand U9887 (N_9887,N_9052,N_9286);
or U9888 (N_9888,N_9345,N_9435);
and U9889 (N_9889,N_9173,N_9081);
or U9890 (N_9890,N_9374,N_9161);
or U9891 (N_9891,N_9440,N_9275);
and U9892 (N_9892,N_9006,N_9465);
nand U9893 (N_9893,N_9355,N_9216);
and U9894 (N_9894,N_9126,N_9061);
nand U9895 (N_9895,N_9209,N_9050);
and U9896 (N_9896,N_9000,N_9379);
and U9897 (N_9897,N_9041,N_9306);
and U9898 (N_9898,N_9378,N_9491);
nor U9899 (N_9899,N_9132,N_9229);
xor U9900 (N_9900,N_9212,N_9285);
and U9901 (N_9901,N_9015,N_9029);
or U9902 (N_9902,N_9316,N_9237);
xnor U9903 (N_9903,N_9330,N_9429);
and U9904 (N_9904,N_9208,N_9364);
or U9905 (N_9905,N_9152,N_9008);
and U9906 (N_9906,N_9366,N_9029);
nor U9907 (N_9907,N_9381,N_9158);
xnor U9908 (N_9908,N_9369,N_9445);
nor U9909 (N_9909,N_9292,N_9474);
or U9910 (N_9910,N_9398,N_9348);
or U9911 (N_9911,N_9008,N_9299);
or U9912 (N_9912,N_9063,N_9001);
xnor U9913 (N_9913,N_9251,N_9023);
nand U9914 (N_9914,N_9143,N_9479);
nand U9915 (N_9915,N_9025,N_9159);
and U9916 (N_9916,N_9055,N_9086);
xor U9917 (N_9917,N_9153,N_9020);
nor U9918 (N_9918,N_9406,N_9156);
nor U9919 (N_9919,N_9403,N_9005);
and U9920 (N_9920,N_9130,N_9326);
or U9921 (N_9921,N_9491,N_9369);
xor U9922 (N_9922,N_9314,N_9311);
nand U9923 (N_9923,N_9351,N_9166);
or U9924 (N_9924,N_9267,N_9394);
nand U9925 (N_9925,N_9124,N_9469);
or U9926 (N_9926,N_9395,N_9180);
and U9927 (N_9927,N_9137,N_9398);
nand U9928 (N_9928,N_9336,N_9405);
and U9929 (N_9929,N_9027,N_9211);
xor U9930 (N_9930,N_9364,N_9007);
xor U9931 (N_9931,N_9393,N_9464);
and U9932 (N_9932,N_9349,N_9499);
nand U9933 (N_9933,N_9444,N_9202);
nor U9934 (N_9934,N_9360,N_9002);
nand U9935 (N_9935,N_9201,N_9408);
nor U9936 (N_9936,N_9314,N_9151);
or U9937 (N_9937,N_9240,N_9166);
or U9938 (N_9938,N_9452,N_9213);
nand U9939 (N_9939,N_9106,N_9370);
xor U9940 (N_9940,N_9331,N_9330);
and U9941 (N_9941,N_9182,N_9386);
and U9942 (N_9942,N_9243,N_9350);
xor U9943 (N_9943,N_9462,N_9077);
or U9944 (N_9944,N_9283,N_9435);
and U9945 (N_9945,N_9455,N_9100);
xnor U9946 (N_9946,N_9154,N_9292);
or U9947 (N_9947,N_9352,N_9196);
and U9948 (N_9948,N_9189,N_9383);
or U9949 (N_9949,N_9399,N_9431);
xor U9950 (N_9950,N_9149,N_9415);
and U9951 (N_9951,N_9434,N_9137);
nand U9952 (N_9952,N_9207,N_9228);
and U9953 (N_9953,N_9317,N_9311);
nand U9954 (N_9954,N_9311,N_9002);
and U9955 (N_9955,N_9233,N_9317);
and U9956 (N_9956,N_9130,N_9364);
and U9957 (N_9957,N_9068,N_9243);
nand U9958 (N_9958,N_9423,N_9172);
and U9959 (N_9959,N_9331,N_9012);
and U9960 (N_9960,N_9367,N_9480);
nand U9961 (N_9961,N_9120,N_9431);
xnor U9962 (N_9962,N_9034,N_9248);
and U9963 (N_9963,N_9488,N_9313);
xnor U9964 (N_9964,N_9264,N_9238);
nor U9965 (N_9965,N_9493,N_9390);
or U9966 (N_9966,N_9410,N_9130);
and U9967 (N_9967,N_9079,N_9111);
nand U9968 (N_9968,N_9366,N_9378);
nor U9969 (N_9969,N_9301,N_9294);
nand U9970 (N_9970,N_9304,N_9027);
xor U9971 (N_9971,N_9313,N_9311);
or U9972 (N_9972,N_9123,N_9484);
or U9973 (N_9973,N_9395,N_9356);
or U9974 (N_9974,N_9474,N_9353);
or U9975 (N_9975,N_9214,N_9465);
and U9976 (N_9976,N_9320,N_9125);
and U9977 (N_9977,N_9468,N_9444);
or U9978 (N_9978,N_9035,N_9041);
nor U9979 (N_9979,N_9367,N_9025);
nor U9980 (N_9980,N_9179,N_9453);
or U9981 (N_9981,N_9073,N_9199);
xor U9982 (N_9982,N_9169,N_9311);
xor U9983 (N_9983,N_9346,N_9199);
xnor U9984 (N_9984,N_9017,N_9431);
nor U9985 (N_9985,N_9101,N_9436);
xnor U9986 (N_9986,N_9152,N_9127);
or U9987 (N_9987,N_9388,N_9181);
or U9988 (N_9988,N_9264,N_9147);
nand U9989 (N_9989,N_9009,N_9078);
or U9990 (N_9990,N_9264,N_9036);
nand U9991 (N_9991,N_9394,N_9266);
or U9992 (N_9992,N_9428,N_9401);
xor U9993 (N_9993,N_9003,N_9115);
or U9994 (N_9994,N_9085,N_9103);
nand U9995 (N_9995,N_9173,N_9051);
and U9996 (N_9996,N_9149,N_9225);
and U9997 (N_9997,N_9282,N_9014);
nand U9998 (N_9998,N_9194,N_9100);
nand U9999 (N_9999,N_9064,N_9266);
nand UO_0 (O_0,N_9686,N_9664);
nand UO_1 (O_1,N_9536,N_9769);
xnor UO_2 (O_2,N_9533,N_9682);
nand UO_3 (O_3,N_9599,N_9576);
or UO_4 (O_4,N_9581,N_9616);
nor UO_5 (O_5,N_9993,N_9757);
xor UO_6 (O_6,N_9890,N_9504);
nand UO_7 (O_7,N_9821,N_9540);
xor UO_8 (O_8,N_9649,N_9822);
and UO_9 (O_9,N_9713,N_9749);
xnor UO_10 (O_10,N_9564,N_9516);
nand UO_11 (O_11,N_9752,N_9955);
xnor UO_12 (O_12,N_9781,N_9835);
xor UO_13 (O_13,N_9964,N_9983);
xor UO_14 (O_14,N_9638,N_9613);
or UO_15 (O_15,N_9839,N_9689);
nand UO_16 (O_16,N_9943,N_9895);
and UO_17 (O_17,N_9913,N_9871);
and UO_18 (O_18,N_9830,N_9806);
xnor UO_19 (O_19,N_9941,N_9783);
and UO_20 (O_20,N_9706,N_9553);
nand UO_21 (O_21,N_9519,N_9787);
or UO_22 (O_22,N_9918,N_9676);
xnor UO_23 (O_23,N_9730,N_9663);
nand UO_24 (O_24,N_9693,N_9865);
or UO_25 (O_25,N_9674,N_9524);
xnor UO_26 (O_26,N_9583,N_9776);
and UO_27 (O_27,N_9579,N_9514);
xor UO_28 (O_28,N_9506,N_9747);
xor UO_29 (O_29,N_9812,N_9860);
or UO_30 (O_30,N_9782,N_9546);
and UO_31 (O_31,N_9665,N_9946);
or UO_32 (O_32,N_9659,N_9673);
nand UO_33 (O_33,N_9523,N_9679);
and UO_34 (O_34,N_9697,N_9695);
nand UO_35 (O_35,N_9605,N_9735);
or UO_36 (O_36,N_9500,N_9932);
or UO_37 (O_37,N_9739,N_9696);
nand UO_38 (O_38,N_9887,N_9882);
nor UO_39 (O_39,N_9520,N_9685);
nor UO_40 (O_40,N_9753,N_9791);
xor UO_41 (O_41,N_9615,N_9784);
and UO_42 (O_42,N_9870,N_9926);
nand UO_43 (O_43,N_9744,N_9774);
xnor UO_44 (O_44,N_9991,N_9601);
and UO_45 (O_45,N_9759,N_9568);
and UO_46 (O_46,N_9900,N_9919);
nand UO_47 (O_47,N_9763,N_9603);
xnor UO_48 (O_48,N_9598,N_9852);
and UO_49 (O_49,N_9803,N_9915);
and UO_50 (O_50,N_9916,N_9814);
nor UO_51 (O_51,N_9580,N_9582);
xnor UO_52 (O_52,N_9847,N_9513);
nor UO_53 (O_53,N_9981,N_9980);
or UO_54 (O_54,N_9878,N_9577);
xnor UO_55 (O_55,N_9646,N_9848);
or UO_56 (O_56,N_9728,N_9829);
xnor UO_57 (O_57,N_9873,N_9670);
xnor UO_58 (O_58,N_9813,N_9794);
xor UO_59 (O_59,N_9905,N_9864);
or UO_60 (O_60,N_9563,N_9885);
or UO_61 (O_61,N_9573,N_9570);
and UO_62 (O_62,N_9779,N_9544);
xor UO_63 (O_63,N_9700,N_9949);
nand UO_64 (O_64,N_9633,N_9771);
nor UO_65 (O_65,N_9656,N_9762);
nand UO_66 (O_66,N_9718,N_9736);
or UO_67 (O_67,N_9600,N_9721);
nor UO_68 (O_68,N_9876,N_9966);
xor UO_69 (O_69,N_9987,N_9979);
nand UO_70 (O_70,N_9856,N_9967);
nor UO_71 (O_71,N_9588,N_9775);
or UO_72 (O_72,N_9716,N_9960);
or UO_73 (O_73,N_9508,N_9522);
and UO_74 (O_74,N_9515,N_9602);
and UO_75 (O_75,N_9559,N_9858);
nor UO_76 (O_76,N_9881,N_9707);
nor UO_77 (O_77,N_9512,N_9518);
xnor UO_78 (O_78,N_9709,N_9554);
nor UO_79 (O_79,N_9810,N_9597);
nand UO_80 (O_80,N_9802,N_9891);
nand UO_81 (O_81,N_9502,N_9666);
xnor UO_82 (O_82,N_9773,N_9703);
or UO_83 (O_83,N_9903,N_9874);
nand UO_84 (O_84,N_9765,N_9928);
or UO_85 (O_85,N_9862,N_9975);
xnor UO_86 (O_86,N_9832,N_9608);
and UO_87 (O_87,N_9974,N_9907);
nor UO_88 (O_88,N_9959,N_9884);
nand UO_89 (O_89,N_9619,N_9680);
or UO_90 (O_90,N_9797,N_9574);
nor UO_91 (O_91,N_9965,N_9953);
and UO_92 (O_92,N_9808,N_9995);
xor UO_93 (O_93,N_9737,N_9732);
and UO_94 (O_94,N_9910,N_9526);
nand UO_95 (O_95,N_9948,N_9755);
and UO_96 (O_96,N_9795,N_9777);
nor UO_97 (O_97,N_9655,N_9584);
and UO_98 (O_98,N_9618,N_9897);
and UO_99 (O_99,N_9911,N_9801);
or UO_100 (O_100,N_9694,N_9868);
or UO_101 (O_101,N_9717,N_9637);
and UO_102 (O_102,N_9780,N_9660);
or UO_103 (O_103,N_9569,N_9990);
nor UO_104 (O_104,N_9701,N_9836);
and UO_105 (O_105,N_9669,N_9840);
or UO_106 (O_106,N_9846,N_9982);
or UO_107 (O_107,N_9617,N_9898);
nor UO_108 (O_108,N_9796,N_9741);
nor UO_109 (O_109,N_9989,N_9889);
and UO_110 (O_110,N_9947,N_9509);
nand UO_111 (O_111,N_9527,N_9719);
nor UO_112 (O_112,N_9970,N_9997);
nor UO_113 (O_113,N_9790,N_9789);
nand UO_114 (O_114,N_9978,N_9675);
nand UO_115 (O_115,N_9611,N_9688);
and UO_116 (O_116,N_9699,N_9861);
and UO_117 (O_117,N_9909,N_9844);
nand UO_118 (O_118,N_9623,N_9825);
nor UO_119 (O_119,N_9788,N_9604);
and UO_120 (O_120,N_9552,N_9992);
xnor UO_121 (O_121,N_9543,N_9743);
nor UO_122 (O_122,N_9920,N_9940);
xnor UO_123 (O_123,N_9756,N_9772);
or UO_124 (O_124,N_9935,N_9770);
and UO_125 (O_125,N_9977,N_9555);
or UO_126 (O_126,N_9845,N_9572);
xor UO_127 (O_127,N_9671,N_9562);
or UO_128 (O_128,N_9786,N_9733);
and UO_129 (O_129,N_9807,N_9609);
xor UO_130 (O_130,N_9621,N_9968);
and UO_131 (O_131,N_9565,N_9505);
and UO_132 (O_132,N_9537,N_9971);
or UO_133 (O_133,N_9921,N_9793);
and UO_134 (O_134,N_9691,N_9930);
and UO_135 (O_135,N_9624,N_9651);
nand UO_136 (O_136,N_9556,N_9531);
xor UO_137 (O_137,N_9571,N_9853);
xnor UO_138 (O_138,N_9710,N_9585);
nand UO_139 (O_139,N_9662,N_9800);
xor UO_140 (O_140,N_9880,N_9541);
or UO_141 (O_141,N_9678,N_9539);
xnor UO_142 (O_142,N_9833,N_9841);
or UO_143 (O_143,N_9622,N_9607);
or UO_144 (O_144,N_9933,N_9723);
xnor UO_145 (O_145,N_9838,N_9594);
xor UO_146 (O_146,N_9866,N_9837);
nor UO_147 (O_147,N_9925,N_9742);
or UO_148 (O_148,N_9785,N_9904);
xor UO_149 (O_149,N_9896,N_9628);
or UO_150 (O_150,N_9994,N_9908);
or UO_151 (O_151,N_9892,N_9627);
nor UO_152 (O_152,N_9625,N_9647);
and UO_153 (O_153,N_9528,N_9818);
nand UO_154 (O_154,N_9681,N_9958);
and UO_155 (O_155,N_9768,N_9614);
nor UO_156 (O_156,N_9766,N_9740);
nor UO_157 (O_157,N_9767,N_9550);
nor UO_158 (O_158,N_9629,N_9653);
xor UO_159 (O_159,N_9729,N_9626);
or UO_160 (O_160,N_9636,N_9996);
or UO_161 (O_161,N_9722,N_9640);
xor UO_162 (O_162,N_9944,N_9809);
or UO_163 (O_163,N_9683,N_9901);
or UO_164 (O_164,N_9883,N_9923);
xor UO_165 (O_165,N_9872,N_9587);
xor UO_166 (O_166,N_9855,N_9798);
xor UO_167 (O_167,N_9917,N_9750);
nand UO_168 (O_168,N_9596,N_9819);
nand UO_169 (O_169,N_9507,N_9510);
or UO_170 (O_170,N_9912,N_9654);
or UO_171 (O_171,N_9863,N_9942);
and UO_172 (O_172,N_9645,N_9644);
and UO_173 (O_173,N_9778,N_9692);
and UO_174 (O_174,N_9529,N_9893);
and UO_175 (O_175,N_9593,N_9672);
nand UO_176 (O_176,N_9999,N_9936);
or UO_177 (O_177,N_9760,N_9525);
xor UO_178 (O_178,N_9561,N_9850);
nor UO_179 (O_179,N_9612,N_9632);
xnor UO_180 (O_180,N_9922,N_9648);
nor UO_181 (O_181,N_9986,N_9545);
nor UO_182 (O_182,N_9690,N_9642);
nand UO_183 (O_183,N_9557,N_9859);
nor UO_184 (O_184,N_9963,N_9879);
nor UO_185 (O_185,N_9724,N_9914);
xnor UO_186 (O_186,N_9877,N_9501);
and UO_187 (O_187,N_9824,N_9590);
nor UO_188 (O_188,N_9754,N_9641);
nand UO_189 (O_189,N_9726,N_9708);
and UO_190 (O_190,N_9575,N_9532);
nand UO_191 (O_191,N_9761,N_9823);
xor UO_192 (O_192,N_9684,N_9843);
or UO_193 (O_193,N_9738,N_9551);
nand UO_194 (O_194,N_9639,N_9988);
and UO_195 (O_195,N_9972,N_9712);
nor UO_196 (O_196,N_9702,N_9857);
nand UO_197 (O_197,N_9951,N_9745);
nor UO_198 (O_198,N_9704,N_9976);
and UO_199 (O_199,N_9530,N_9589);
xnor UO_200 (O_200,N_9620,N_9998);
or UO_201 (O_201,N_9630,N_9985);
and UO_202 (O_202,N_9535,N_9867);
or UO_203 (O_203,N_9503,N_9937);
or UO_204 (O_204,N_9711,N_9714);
xor UO_205 (O_205,N_9652,N_9854);
nand UO_206 (O_206,N_9635,N_9817);
xnor UO_207 (O_207,N_9658,N_9816);
and UO_208 (O_208,N_9547,N_9952);
nor UO_209 (O_209,N_9827,N_9746);
and UO_210 (O_210,N_9668,N_9610);
nand UO_211 (O_211,N_9657,N_9548);
or UO_212 (O_212,N_9924,N_9899);
and UO_213 (O_213,N_9815,N_9849);
nand UO_214 (O_214,N_9725,N_9631);
nor UO_215 (O_215,N_9834,N_9939);
nor UO_216 (O_216,N_9586,N_9606);
and UO_217 (O_217,N_9560,N_9826);
or UO_218 (O_218,N_9591,N_9938);
xnor UO_219 (O_219,N_9805,N_9727);
nand UO_220 (O_220,N_9961,N_9894);
nand UO_221 (O_221,N_9534,N_9984);
nor UO_222 (O_222,N_9764,N_9578);
xnor UO_223 (O_223,N_9969,N_9831);
or UO_224 (O_224,N_9698,N_9875);
and UO_225 (O_225,N_9643,N_9566);
nand UO_226 (O_226,N_9799,N_9811);
nor UO_227 (O_227,N_9731,N_9634);
nor UO_228 (O_228,N_9558,N_9842);
xnor UO_229 (O_229,N_9820,N_9705);
and UO_230 (O_230,N_9929,N_9954);
or UO_231 (O_231,N_9720,N_9661);
nor UO_232 (O_232,N_9521,N_9748);
and UO_233 (O_233,N_9567,N_9595);
nand UO_234 (O_234,N_9906,N_9828);
or UO_235 (O_235,N_9804,N_9538);
xnor UO_236 (O_236,N_9956,N_9886);
nand UO_237 (O_237,N_9751,N_9931);
and UO_238 (O_238,N_9973,N_9945);
nand UO_239 (O_239,N_9715,N_9687);
nand UO_240 (O_240,N_9851,N_9888);
or UO_241 (O_241,N_9592,N_9650);
and UO_242 (O_242,N_9667,N_9957);
nand UO_243 (O_243,N_9758,N_9934);
nand UO_244 (O_244,N_9511,N_9734);
and UO_245 (O_245,N_9950,N_9677);
xnor UO_246 (O_246,N_9517,N_9542);
nor UO_247 (O_247,N_9902,N_9962);
nor UO_248 (O_248,N_9549,N_9792);
or UO_249 (O_249,N_9869,N_9927);
or UO_250 (O_250,N_9998,N_9553);
or UO_251 (O_251,N_9715,N_9865);
nor UO_252 (O_252,N_9691,N_9509);
or UO_253 (O_253,N_9950,N_9936);
nor UO_254 (O_254,N_9578,N_9974);
xor UO_255 (O_255,N_9898,N_9786);
nor UO_256 (O_256,N_9916,N_9717);
nor UO_257 (O_257,N_9597,N_9598);
and UO_258 (O_258,N_9579,N_9701);
xor UO_259 (O_259,N_9865,N_9797);
and UO_260 (O_260,N_9709,N_9635);
xnor UO_261 (O_261,N_9762,N_9529);
or UO_262 (O_262,N_9992,N_9590);
xnor UO_263 (O_263,N_9696,N_9719);
or UO_264 (O_264,N_9755,N_9829);
nand UO_265 (O_265,N_9833,N_9929);
nand UO_266 (O_266,N_9676,N_9855);
nor UO_267 (O_267,N_9956,N_9554);
and UO_268 (O_268,N_9824,N_9568);
nand UO_269 (O_269,N_9734,N_9673);
or UO_270 (O_270,N_9553,N_9845);
xor UO_271 (O_271,N_9957,N_9902);
or UO_272 (O_272,N_9522,N_9776);
or UO_273 (O_273,N_9694,N_9898);
and UO_274 (O_274,N_9792,N_9898);
nand UO_275 (O_275,N_9766,N_9737);
nor UO_276 (O_276,N_9684,N_9547);
xnor UO_277 (O_277,N_9964,N_9948);
xnor UO_278 (O_278,N_9816,N_9662);
xnor UO_279 (O_279,N_9548,N_9703);
xnor UO_280 (O_280,N_9872,N_9903);
xor UO_281 (O_281,N_9969,N_9586);
xor UO_282 (O_282,N_9955,N_9739);
xor UO_283 (O_283,N_9794,N_9947);
nand UO_284 (O_284,N_9871,N_9559);
xor UO_285 (O_285,N_9945,N_9872);
xor UO_286 (O_286,N_9580,N_9915);
or UO_287 (O_287,N_9814,N_9837);
or UO_288 (O_288,N_9653,N_9556);
and UO_289 (O_289,N_9931,N_9749);
nor UO_290 (O_290,N_9681,N_9766);
nor UO_291 (O_291,N_9713,N_9895);
and UO_292 (O_292,N_9596,N_9738);
and UO_293 (O_293,N_9785,N_9689);
or UO_294 (O_294,N_9700,N_9864);
and UO_295 (O_295,N_9965,N_9904);
or UO_296 (O_296,N_9566,N_9721);
xnor UO_297 (O_297,N_9828,N_9865);
or UO_298 (O_298,N_9715,N_9859);
nand UO_299 (O_299,N_9746,N_9924);
and UO_300 (O_300,N_9758,N_9745);
and UO_301 (O_301,N_9836,N_9667);
xnor UO_302 (O_302,N_9709,N_9872);
nand UO_303 (O_303,N_9780,N_9626);
and UO_304 (O_304,N_9898,N_9851);
nor UO_305 (O_305,N_9804,N_9828);
xor UO_306 (O_306,N_9589,N_9523);
and UO_307 (O_307,N_9736,N_9996);
nor UO_308 (O_308,N_9581,N_9953);
nor UO_309 (O_309,N_9908,N_9571);
nor UO_310 (O_310,N_9693,N_9806);
nor UO_311 (O_311,N_9783,N_9805);
xor UO_312 (O_312,N_9628,N_9771);
nor UO_313 (O_313,N_9795,N_9896);
and UO_314 (O_314,N_9747,N_9552);
or UO_315 (O_315,N_9877,N_9943);
nand UO_316 (O_316,N_9613,N_9917);
or UO_317 (O_317,N_9510,N_9952);
xnor UO_318 (O_318,N_9663,N_9655);
xor UO_319 (O_319,N_9635,N_9864);
nor UO_320 (O_320,N_9945,N_9905);
nand UO_321 (O_321,N_9831,N_9645);
xor UO_322 (O_322,N_9639,N_9504);
or UO_323 (O_323,N_9858,N_9915);
xnor UO_324 (O_324,N_9776,N_9592);
and UO_325 (O_325,N_9854,N_9723);
nand UO_326 (O_326,N_9563,N_9601);
xnor UO_327 (O_327,N_9762,N_9551);
nand UO_328 (O_328,N_9785,N_9544);
nand UO_329 (O_329,N_9676,N_9981);
xnor UO_330 (O_330,N_9874,N_9592);
nor UO_331 (O_331,N_9870,N_9760);
nand UO_332 (O_332,N_9870,N_9660);
xnor UO_333 (O_333,N_9580,N_9873);
and UO_334 (O_334,N_9643,N_9585);
xnor UO_335 (O_335,N_9893,N_9919);
or UO_336 (O_336,N_9764,N_9572);
nand UO_337 (O_337,N_9838,N_9698);
nand UO_338 (O_338,N_9896,N_9988);
and UO_339 (O_339,N_9920,N_9939);
nor UO_340 (O_340,N_9983,N_9888);
and UO_341 (O_341,N_9859,N_9974);
and UO_342 (O_342,N_9880,N_9669);
xor UO_343 (O_343,N_9921,N_9813);
or UO_344 (O_344,N_9515,N_9851);
xor UO_345 (O_345,N_9581,N_9874);
or UO_346 (O_346,N_9979,N_9650);
nand UO_347 (O_347,N_9613,N_9965);
xnor UO_348 (O_348,N_9740,N_9794);
and UO_349 (O_349,N_9557,N_9800);
xnor UO_350 (O_350,N_9980,N_9883);
nand UO_351 (O_351,N_9656,N_9941);
nand UO_352 (O_352,N_9610,N_9833);
nand UO_353 (O_353,N_9731,N_9546);
or UO_354 (O_354,N_9936,N_9593);
nand UO_355 (O_355,N_9832,N_9771);
or UO_356 (O_356,N_9947,N_9633);
and UO_357 (O_357,N_9976,N_9666);
nor UO_358 (O_358,N_9623,N_9839);
nand UO_359 (O_359,N_9599,N_9902);
nand UO_360 (O_360,N_9775,N_9817);
and UO_361 (O_361,N_9540,N_9829);
nor UO_362 (O_362,N_9912,N_9934);
nand UO_363 (O_363,N_9746,N_9981);
nand UO_364 (O_364,N_9649,N_9727);
or UO_365 (O_365,N_9705,N_9614);
and UO_366 (O_366,N_9583,N_9507);
nand UO_367 (O_367,N_9668,N_9768);
xor UO_368 (O_368,N_9860,N_9843);
xnor UO_369 (O_369,N_9998,N_9600);
nand UO_370 (O_370,N_9948,N_9841);
nand UO_371 (O_371,N_9770,N_9619);
nand UO_372 (O_372,N_9537,N_9824);
nand UO_373 (O_373,N_9937,N_9898);
and UO_374 (O_374,N_9812,N_9666);
or UO_375 (O_375,N_9643,N_9982);
or UO_376 (O_376,N_9934,N_9829);
xnor UO_377 (O_377,N_9653,N_9508);
xor UO_378 (O_378,N_9830,N_9656);
nand UO_379 (O_379,N_9735,N_9627);
nand UO_380 (O_380,N_9575,N_9849);
nor UO_381 (O_381,N_9645,N_9733);
and UO_382 (O_382,N_9749,N_9714);
xor UO_383 (O_383,N_9569,N_9618);
nor UO_384 (O_384,N_9617,N_9596);
and UO_385 (O_385,N_9538,N_9945);
and UO_386 (O_386,N_9644,N_9673);
xnor UO_387 (O_387,N_9772,N_9966);
nor UO_388 (O_388,N_9637,N_9982);
or UO_389 (O_389,N_9683,N_9867);
or UO_390 (O_390,N_9803,N_9902);
xnor UO_391 (O_391,N_9865,N_9959);
xnor UO_392 (O_392,N_9872,N_9609);
or UO_393 (O_393,N_9711,N_9797);
nand UO_394 (O_394,N_9565,N_9669);
xor UO_395 (O_395,N_9892,N_9949);
xor UO_396 (O_396,N_9832,N_9840);
nand UO_397 (O_397,N_9851,N_9516);
xnor UO_398 (O_398,N_9989,N_9688);
or UO_399 (O_399,N_9826,N_9655);
nor UO_400 (O_400,N_9968,N_9744);
xor UO_401 (O_401,N_9594,N_9908);
nand UO_402 (O_402,N_9583,N_9719);
and UO_403 (O_403,N_9523,N_9558);
nor UO_404 (O_404,N_9823,N_9500);
xor UO_405 (O_405,N_9560,N_9768);
or UO_406 (O_406,N_9693,N_9566);
nor UO_407 (O_407,N_9519,N_9546);
nand UO_408 (O_408,N_9742,N_9692);
and UO_409 (O_409,N_9777,N_9643);
xor UO_410 (O_410,N_9959,N_9975);
and UO_411 (O_411,N_9945,N_9921);
nor UO_412 (O_412,N_9824,N_9942);
nor UO_413 (O_413,N_9975,N_9664);
or UO_414 (O_414,N_9659,N_9657);
and UO_415 (O_415,N_9541,N_9913);
nor UO_416 (O_416,N_9521,N_9856);
and UO_417 (O_417,N_9839,N_9985);
xor UO_418 (O_418,N_9845,N_9936);
and UO_419 (O_419,N_9634,N_9935);
and UO_420 (O_420,N_9532,N_9878);
nor UO_421 (O_421,N_9849,N_9701);
or UO_422 (O_422,N_9935,N_9908);
nor UO_423 (O_423,N_9577,N_9615);
and UO_424 (O_424,N_9515,N_9548);
and UO_425 (O_425,N_9780,N_9969);
xor UO_426 (O_426,N_9678,N_9782);
nand UO_427 (O_427,N_9888,N_9604);
nand UO_428 (O_428,N_9656,N_9814);
nand UO_429 (O_429,N_9949,N_9740);
and UO_430 (O_430,N_9936,N_9919);
nand UO_431 (O_431,N_9635,N_9858);
nand UO_432 (O_432,N_9873,N_9951);
nand UO_433 (O_433,N_9651,N_9717);
nand UO_434 (O_434,N_9879,N_9635);
xnor UO_435 (O_435,N_9999,N_9788);
nor UO_436 (O_436,N_9580,N_9655);
nand UO_437 (O_437,N_9752,N_9703);
or UO_438 (O_438,N_9670,N_9945);
nor UO_439 (O_439,N_9764,N_9942);
nor UO_440 (O_440,N_9903,N_9693);
xnor UO_441 (O_441,N_9815,N_9525);
nand UO_442 (O_442,N_9893,N_9955);
nand UO_443 (O_443,N_9548,N_9732);
or UO_444 (O_444,N_9819,N_9609);
and UO_445 (O_445,N_9627,N_9827);
and UO_446 (O_446,N_9582,N_9799);
or UO_447 (O_447,N_9575,N_9551);
nor UO_448 (O_448,N_9590,N_9916);
nor UO_449 (O_449,N_9572,N_9940);
xor UO_450 (O_450,N_9754,N_9832);
xnor UO_451 (O_451,N_9517,N_9984);
or UO_452 (O_452,N_9531,N_9707);
and UO_453 (O_453,N_9851,N_9967);
nand UO_454 (O_454,N_9926,N_9956);
nor UO_455 (O_455,N_9814,N_9779);
and UO_456 (O_456,N_9899,N_9530);
nand UO_457 (O_457,N_9893,N_9716);
nor UO_458 (O_458,N_9852,N_9714);
nand UO_459 (O_459,N_9526,N_9818);
or UO_460 (O_460,N_9550,N_9593);
xor UO_461 (O_461,N_9623,N_9741);
xor UO_462 (O_462,N_9859,N_9784);
and UO_463 (O_463,N_9942,N_9871);
xnor UO_464 (O_464,N_9895,N_9644);
or UO_465 (O_465,N_9913,N_9786);
nand UO_466 (O_466,N_9676,N_9638);
or UO_467 (O_467,N_9726,N_9674);
and UO_468 (O_468,N_9613,N_9725);
and UO_469 (O_469,N_9534,N_9539);
xor UO_470 (O_470,N_9645,N_9805);
or UO_471 (O_471,N_9878,N_9552);
nor UO_472 (O_472,N_9788,N_9676);
xnor UO_473 (O_473,N_9578,N_9973);
nand UO_474 (O_474,N_9529,N_9707);
nand UO_475 (O_475,N_9854,N_9634);
or UO_476 (O_476,N_9654,N_9632);
nand UO_477 (O_477,N_9772,N_9812);
or UO_478 (O_478,N_9992,N_9672);
and UO_479 (O_479,N_9526,N_9586);
nand UO_480 (O_480,N_9718,N_9820);
or UO_481 (O_481,N_9728,N_9933);
nand UO_482 (O_482,N_9685,N_9703);
or UO_483 (O_483,N_9708,N_9718);
or UO_484 (O_484,N_9531,N_9787);
or UO_485 (O_485,N_9905,N_9833);
or UO_486 (O_486,N_9872,N_9687);
xnor UO_487 (O_487,N_9507,N_9647);
xnor UO_488 (O_488,N_9599,N_9595);
nand UO_489 (O_489,N_9845,N_9903);
xnor UO_490 (O_490,N_9961,N_9838);
nor UO_491 (O_491,N_9625,N_9856);
nor UO_492 (O_492,N_9848,N_9638);
or UO_493 (O_493,N_9995,N_9959);
xor UO_494 (O_494,N_9815,N_9771);
or UO_495 (O_495,N_9570,N_9805);
nor UO_496 (O_496,N_9712,N_9540);
and UO_497 (O_497,N_9763,N_9570);
and UO_498 (O_498,N_9745,N_9800);
and UO_499 (O_499,N_9724,N_9909);
nor UO_500 (O_500,N_9929,N_9910);
or UO_501 (O_501,N_9864,N_9617);
xor UO_502 (O_502,N_9695,N_9960);
nor UO_503 (O_503,N_9902,N_9688);
nand UO_504 (O_504,N_9821,N_9722);
nand UO_505 (O_505,N_9881,N_9524);
nor UO_506 (O_506,N_9504,N_9544);
xor UO_507 (O_507,N_9946,N_9849);
nand UO_508 (O_508,N_9955,N_9518);
nand UO_509 (O_509,N_9626,N_9769);
nand UO_510 (O_510,N_9992,N_9760);
and UO_511 (O_511,N_9619,N_9900);
or UO_512 (O_512,N_9652,N_9722);
xor UO_513 (O_513,N_9732,N_9815);
nand UO_514 (O_514,N_9897,N_9764);
nor UO_515 (O_515,N_9713,N_9913);
or UO_516 (O_516,N_9769,N_9640);
and UO_517 (O_517,N_9804,N_9790);
or UO_518 (O_518,N_9931,N_9643);
nor UO_519 (O_519,N_9795,N_9881);
nand UO_520 (O_520,N_9995,N_9993);
nand UO_521 (O_521,N_9917,N_9876);
nand UO_522 (O_522,N_9572,N_9917);
nand UO_523 (O_523,N_9735,N_9601);
xnor UO_524 (O_524,N_9998,N_9853);
xor UO_525 (O_525,N_9606,N_9591);
and UO_526 (O_526,N_9632,N_9606);
nor UO_527 (O_527,N_9692,N_9919);
nand UO_528 (O_528,N_9557,N_9745);
nand UO_529 (O_529,N_9511,N_9943);
and UO_530 (O_530,N_9916,N_9997);
nand UO_531 (O_531,N_9983,N_9761);
and UO_532 (O_532,N_9672,N_9660);
or UO_533 (O_533,N_9975,N_9738);
nor UO_534 (O_534,N_9565,N_9854);
xor UO_535 (O_535,N_9688,N_9966);
and UO_536 (O_536,N_9715,N_9743);
or UO_537 (O_537,N_9662,N_9777);
nor UO_538 (O_538,N_9909,N_9732);
xor UO_539 (O_539,N_9767,N_9691);
and UO_540 (O_540,N_9556,N_9738);
or UO_541 (O_541,N_9807,N_9612);
xor UO_542 (O_542,N_9911,N_9792);
or UO_543 (O_543,N_9919,N_9950);
nand UO_544 (O_544,N_9560,N_9841);
or UO_545 (O_545,N_9684,N_9860);
and UO_546 (O_546,N_9694,N_9520);
and UO_547 (O_547,N_9509,N_9849);
or UO_548 (O_548,N_9655,N_9519);
nand UO_549 (O_549,N_9818,N_9933);
nor UO_550 (O_550,N_9795,N_9544);
and UO_551 (O_551,N_9857,N_9598);
xor UO_552 (O_552,N_9502,N_9584);
or UO_553 (O_553,N_9541,N_9668);
nand UO_554 (O_554,N_9945,N_9770);
and UO_555 (O_555,N_9624,N_9725);
nand UO_556 (O_556,N_9946,N_9541);
nand UO_557 (O_557,N_9535,N_9950);
xor UO_558 (O_558,N_9635,N_9567);
nor UO_559 (O_559,N_9672,N_9600);
xnor UO_560 (O_560,N_9812,N_9536);
nand UO_561 (O_561,N_9882,N_9739);
xor UO_562 (O_562,N_9777,N_9647);
nand UO_563 (O_563,N_9588,N_9646);
or UO_564 (O_564,N_9511,N_9750);
nand UO_565 (O_565,N_9889,N_9673);
nand UO_566 (O_566,N_9734,N_9652);
or UO_567 (O_567,N_9755,N_9676);
nor UO_568 (O_568,N_9904,N_9672);
and UO_569 (O_569,N_9545,N_9552);
and UO_570 (O_570,N_9966,N_9771);
and UO_571 (O_571,N_9885,N_9735);
or UO_572 (O_572,N_9814,N_9934);
nand UO_573 (O_573,N_9789,N_9845);
xor UO_574 (O_574,N_9741,N_9534);
or UO_575 (O_575,N_9527,N_9854);
xnor UO_576 (O_576,N_9509,N_9781);
nand UO_577 (O_577,N_9945,N_9790);
or UO_578 (O_578,N_9881,N_9639);
nor UO_579 (O_579,N_9674,N_9943);
xnor UO_580 (O_580,N_9840,N_9552);
and UO_581 (O_581,N_9732,N_9995);
nand UO_582 (O_582,N_9956,N_9951);
nand UO_583 (O_583,N_9749,N_9510);
and UO_584 (O_584,N_9899,N_9822);
or UO_585 (O_585,N_9754,N_9549);
nor UO_586 (O_586,N_9877,N_9783);
or UO_587 (O_587,N_9720,N_9676);
and UO_588 (O_588,N_9703,N_9542);
nand UO_589 (O_589,N_9627,N_9521);
or UO_590 (O_590,N_9815,N_9673);
and UO_591 (O_591,N_9928,N_9929);
nand UO_592 (O_592,N_9600,N_9889);
xnor UO_593 (O_593,N_9838,N_9944);
nand UO_594 (O_594,N_9839,N_9743);
xor UO_595 (O_595,N_9981,N_9699);
xor UO_596 (O_596,N_9621,N_9903);
nand UO_597 (O_597,N_9988,N_9694);
nand UO_598 (O_598,N_9875,N_9860);
nand UO_599 (O_599,N_9825,N_9874);
xor UO_600 (O_600,N_9914,N_9959);
xnor UO_601 (O_601,N_9609,N_9843);
xnor UO_602 (O_602,N_9858,N_9770);
nand UO_603 (O_603,N_9730,N_9689);
or UO_604 (O_604,N_9570,N_9612);
nand UO_605 (O_605,N_9822,N_9722);
or UO_606 (O_606,N_9893,N_9606);
nor UO_607 (O_607,N_9669,N_9723);
or UO_608 (O_608,N_9503,N_9994);
nor UO_609 (O_609,N_9901,N_9629);
and UO_610 (O_610,N_9982,N_9543);
xor UO_611 (O_611,N_9571,N_9768);
or UO_612 (O_612,N_9920,N_9758);
and UO_613 (O_613,N_9910,N_9533);
xor UO_614 (O_614,N_9832,N_9761);
and UO_615 (O_615,N_9563,N_9887);
xnor UO_616 (O_616,N_9993,N_9588);
nor UO_617 (O_617,N_9996,N_9984);
nor UO_618 (O_618,N_9530,N_9681);
or UO_619 (O_619,N_9843,N_9744);
or UO_620 (O_620,N_9547,N_9681);
and UO_621 (O_621,N_9764,N_9765);
or UO_622 (O_622,N_9513,N_9617);
nand UO_623 (O_623,N_9919,N_9856);
nor UO_624 (O_624,N_9617,N_9761);
or UO_625 (O_625,N_9989,N_9799);
or UO_626 (O_626,N_9672,N_9621);
nand UO_627 (O_627,N_9958,N_9890);
nor UO_628 (O_628,N_9607,N_9946);
and UO_629 (O_629,N_9581,N_9678);
or UO_630 (O_630,N_9841,N_9521);
nand UO_631 (O_631,N_9526,N_9724);
nor UO_632 (O_632,N_9948,N_9796);
and UO_633 (O_633,N_9792,N_9630);
and UO_634 (O_634,N_9675,N_9879);
nand UO_635 (O_635,N_9638,N_9642);
and UO_636 (O_636,N_9602,N_9524);
xor UO_637 (O_637,N_9647,N_9749);
or UO_638 (O_638,N_9885,N_9566);
nor UO_639 (O_639,N_9842,N_9793);
nand UO_640 (O_640,N_9649,N_9916);
or UO_641 (O_641,N_9913,N_9739);
or UO_642 (O_642,N_9720,N_9796);
nor UO_643 (O_643,N_9879,N_9897);
or UO_644 (O_644,N_9887,N_9853);
nor UO_645 (O_645,N_9705,N_9660);
xor UO_646 (O_646,N_9984,N_9664);
or UO_647 (O_647,N_9559,N_9749);
nor UO_648 (O_648,N_9627,N_9550);
nand UO_649 (O_649,N_9776,N_9902);
nor UO_650 (O_650,N_9864,N_9971);
nand UO_651 (O_651,N_9690,N_9563);
xnor UO_652 (O_652,N_9942,N_9800);
or UO_653 (O_653,N_9931,N_9860);
nand UO_654 (O_654,N_9597,N_9761);
and UO_655 (O_655,N_9642,N_9712);
and UO_656 (O_656,N_9656,N_9881);
nor UO_657 (O_657,N_9919,N_9781);
nor UO_658 (O_658,N_9682,N_9534);
and UO_659 (O_659,N_9638,N_9950);
and UO_660 (O_660,N_9694,N_9826);
or UO_661 (O_661,N_9726,N_9561);
or UO_662 (O_662,N_9750,N_9781);
xnor UO_663 (O_663,N_9692,N_9532);
or UO_664 (O_664,N_9632,N_9583);
or UO_665 (O_665,N_9612,N_9917);
and UO_666 (O_666,N_9979,N_9886);
xnor UO_667 (O_667,N_9679,N_9608);
nand UO_668 (O_668,N_9768,N_9564);
xnor UO_669 (O_669,N_9507,N_9601);
or UO_670 (O_670,N_9722,N_9980);
nor UO_671 (O_671,N_9854,N_9778);
and UO_672 (O_672,N_9884,N_9954);
nor UO_673 (O_673,N_9549,N_9931);
and UO_674 (O_674,N_9810,N_9705);
nor UO_675 (O_675,N_9579,N_9689);
and UO_676 (O_676,N_9945,N_9645);
nand UO_677 (O_677,N_9574,N_9634);
or UO_678 (O_678,N_9771,N_9510);
nor UO_679 (O_679,N_9530,N_9639);
nor UO_680 (O_680,N_9720,N_9906);
nor UO_681 (O_681,N_9954,N_9542);
nand UO_682 (O_682,N_9834,N_9790);
nor UO_683 (O_683,N_9696,N_9504);
or UO_684 (O_684,N_9947,N_9616);
xor UO_685 (O_685,N_9865,N_9606);
xnor UO_686 (O_686,N_9524,N_9874);
nor UO_687 (O_687,N_9919,N_9897);
xnor UO_688 (O_688,N_9627,N_9648);
nor UO_689 (O_689,N_9556,N_9922);
and UO_690 (O_690,N_9564,N_9935);
xor UO_691 (O_691,N_9960,N_9983);
and UO_692 (O_692,N_9547,N_9796);
nor UO_693 (O_693,N_9794,N_9846);
xor UO_694 (O_694,N_9581,N_9656);
nor UO_695 (O_695,N_9649,N_9675);
and UO_696 (O_696,N_9940,N_9904);
xnor UO_697 (O_697,N_9960,N_9893);
nand UO_698 (O_698,N_9845,N_9979);
xnor UO_699 (O_699,N_9539,N_9980);
and UO_700 (O_700,N_9723,N_9813);
nand UO_701 (O_701,N_9590,N_9861);
nand UO_702 (O_702,N_9925,N_9590);
nor UO_703 (O_703,N_9530,N_9578);
xor UO_704 (O_704,N_9919,N_9679);
or UO_705 (O_705,N_9799,N_9898);
or UO_706 (O_706,N_9647,N_9741);
nand UO_707 (O_707,N_9607,N_9829);
xnor UO_708 (O_708,N_9635,N_9995);
xnor UO_709 (O_709,N_9997,N_9830);
xnor UO_710 (O_710,N_9552,N_9514);
nand UO_711 (O_711,N_9891,N_9580);
or UO_712 (O_712,N_9516,N_9865);
and UO_713 (O_713,N_9943,N_9856);
and UO_714 (O_714,N_9690,N_9707);
nor UO_715 (O_715,N_9848,N_9980);
nor UO_716 (O_716,N_9709,N_9687);
nand UO_717 (O_717,N_9574,N_9721);
nor UO_718 (O_718,N_9953,N_9784);
or UO_719 (O_719,N_9833,N_9960);
xor UO_720 (O_720,N_9533,N_9851);
nor UO_721 (O_721,N_9519,N_9789);
or UO_722 (O_722,N_9862,N_9537);
nand UO_723 (O_723,N_9658,N_9823);
and UO_724 (O_724,N_9735,N_9730);
nor UO_725 (O_725,N_9640,N_9733);
nand UO_726 (O_726,N_9628,N_9788);
nor UO_727 (O_727,N_9789,N_9706);
xor UO_728 (O_728,N_9710,N_9985);
and UO_729 (O_729,N_9555,N_9841);
nand UO_730 (O_730,N_9687,N_9799);
xnor UO_731 (O_731,N_9939,N_9995);
or UO_732 (O_732,N_9960,N_9675);
xor UO_733 (O_733,N_9932,N_9664);
nor UO_734 (O_734,N_9506,N_9519);
nor UO_735 (O_735,N_9958,N_9795);
nor UO_736 (O_736,N_9898,N_9580);
or UO_737 (O_737,N_9822,N_9551);
nor UO_738 (O_738,N_9960,N_9669);
and UO_739 (O_739,N_9965,N_9935);
and UO_740 (O_740,N_9645,N_9891);
xnor UO_741 (O_741,N_9873,N_9845);
nor UO_742 (O_742,N_9740,N_9684);
nor UO_743 (O_743,N_9993,N_9619);
nor UO_744 (O_744,N_9919,N_9803);
xnor UO_745 (O_745,N_9945,N_9531);
nand UO_746 (O_746,N_9935,N_9754);
nand UO_747 (O_747,N_9898,N_9791);
nor UO_748 (O_748,N_9539,N_9928);
nand UO_749 (O_749,N_9532,N_9903);
nor UO_750 (O_750,N_9714,N_9525);
or UO_751 (O_751,N_9844,N_9796);
nand UO_752 (O_752,N_9755,N_9701);
or UO_753 (O_753,N_9961,N_9956);
nand UO_754 (O_754,N_9611,N_9771);
and UO_755 (O_755,N_9572,N_9870);
and UO_756 (O_756,N_9595,N_9601);
or UO_757 (O_757,N_9560,N_9971);
xnor UO_758 (O_758,N_9756,N_9856);
or UO_759 (O_759,N_9901,N_9504);
or UO_760 (O_760,N_9924,N_9722);
xnor UO_761 (O_761,N_9728,N_9808);
and UO_762 (O_762,N_9599,N_9742);
nor UO_763 (O_763,N_9944,N_9977);
xnor UO_764 (O_764,N_9814,N_9616);
and UO_765 (O_765,N_9740,N_9869);
or UO_766 (O_766,N_9849,N_9629);
and UO_767 (O_767,N_9801,N_9711);
nor UO_768 (O_768,N_9720,N_9816);
xor UO_769 (O_769,N_9876,N_9870);
nor UO_770 (O_770,N_9780,N_9589);
and UO_771 (O_771,N_9610,N_9674);
nor UO_772 (O_772,N_9984,N_9673);
xor UO_773 (O_773,N_9802,N_9601);
xor UO_774 (O_774,N_9620,N_9673);
and UO_775 (O_775,N_9605,N_9523);
nor UO_776 (O_776,N_9504,N_9973);
nor UO_777 (O_777,N_9552,N_9577);
xor UO_778 (O_778,N_9579,N_9577);
nor UO_779 (O_779,N_9556,N_9968);
nand UO_780 (O_780,N_9541,N_9985);
xnor UO_781 (O_781,N_9872,N_9958);
nor UO_782 (O_782,N_9947,N_9507);
and UO_783 (O_783,N_9583,N_9968);
nand UO_784 (O_784,N_9706,N_9809);
or UO_785 (O_785,N_9755,N_9631);
xor UO_786 (O_786,N_9825,N_9709);
nand UO_787 (O_787,N_9748,N_9901);
and UO_788 (O_788,N_9971,N_9865);
or UO_789 (O_789,N_9549,N_9821);
and UO_790 (O_790,N_9787,N_9841);
or UO_791 (O_791,N_9853,N_9657);
xor UO_792 (O_792,N_9880,N_9516);
nor UO_793 (O_793,N_9846,N_9922);
nand UO_794 (O_794,N_9506,N_9715);
or UO_795 (O_795,N_9519,N_9508);
or UO_796 (O_796,N_9783,N_9672);
nor UO_797 (O_797,N_9925,N_9775);
nor UO_798 (O_798,N_9601,N_9581);
xor UO_799 (O_799,N_9862,N_9951);
and UO_800 (O_800,N_9709,N_9813);
and UO_801 (O_801,N_9750,N_9974);
nand UO_802 (O_802,N_9920,N_9837);
nand UO_803 (O_803,N_9939,N_9521);
xnor UO_804 (O_804,N_9821,N_9841);
nand UO_805 (O_805,N_9619,N_9841);
or UO_806 (O_806,N_9849,N_9772);
or UO_807 (O_807,N_9670,N_9637);
xor UO_808 (O_808,N_9967,N_9831);
nor UO_809 (O_809,N_9953,N_9868);
xor UO_810 (O_810,N_9991,N_9729);
xor UO_811 (O_811,N_9733,N_9787);
nor UO_812 (O_812,N_9611,N_9547);
or UO_813 (O_813,N_9890,N_9864);
nor UO_814 (O_814,N_9604,N_9851);
and UO_815 (O_815,N_9633,N_9595);
xor UO_816 (O_816,N_9951,N_9522);
nor UO_817 (O_817,N_9687,N_9954);
xor UO_818 (O_818,N_9591,N_9785);
nor UO_819 (O_819,N_9633,N_9654);
or UO_820 (O_820,N_9872,N_9699);
or UO_821 (O_821,N_9528,N_9664);
or UO_822 (O_822,N_9990,N_9517);
xor UO_823 (O_823,N_9541,N_9884);
or UO_824 (O_824,N_9934,N_9982);
nand UO_825 (O_825,N_9623,N_9661);
nor UO_826 (O_826,N_9975,N_9836);
nand UO_827 (O_827,N_9821,N_9997);
nand UO_828 (O_828,N_9715,N_9951);
or UO_829 (O_829,N_9836,N_9796);
and UO_830 (O_830,N_9946,N_9905);
and UO_831 (O_831,N_9844,N_9933);
xor UO_832 (O_832,N_9593,N_9633);
and UO_833 (O_833,N_9589,N_9827);
nor UO_834 (O_834,N_9747,N_9761);
or UO_835 (O_835,N_9634,N_9647);
and UO_836 (O_836,N_9681,N_9899);
nand UO_837 (O_837,N_9916,N_9891);
or UO_838 (O_838,N_9923,N_9616);
or UO_839 (O_839,N_9616,N_9759);
or UO_840 (O_840,N_9858,N_9788);
nor UO_841 (O_841,N_9716,N_9997);
nor UO_842 (O_842,N_9929,N_9918);
and UO_843 (O_843,N_9651,N_9617);
or UO_844 (O_844,N_9511,N_9652);
nor UO_845 (O_845,N_9500,N_9709);
nand UO_846 (O_846,N_9790,N_9998);
nor UO_847 (O_847,N_9651,N_9908);
nor UO_848 (O_848,N_9779,N_9993);
nand UO_849 (O_849,N_9609,N_9797);
or UO_850 (O_850,N_9720,N_9728);
nor UO_851 (O_851,N_9579,N_9952);
or UO_852 (O_852,N_9550,N_9556);
nor UO_853 (O_853,N_9731,N_9563);
or UO_854 (O_854,N_9762,N_9711);
nor UO_855 (O_855,N_9816,N_9815);
or UO_856 (O_856,N_9895,N_9997);
xnor UO_857 (O_857,N_9632,N_9911);
or UO_858 (O_858,N_9911,N_9591);
nor UO_859 (O_859,N_9818,N_9727);
xnor UO_860 (O_860,N_9911,N_9712);
nand UO_861 (O_861,N_9557,N_9647);
nand UO_862 (O_862,N_9565,N_9707);
or UO_863 (O_863,N_9945,N_9807);
nand UO_864 (O_864,N_9535,N_9769);
or UO_865 (O_865,N_9882,N_9546);
or UO_866 (O_866,N_9664,N_9986);
nor UO_867 (O_867,N_9572,N_9898);
xor UO_868 (O_868,N_9705,N_9648);
or UO_869 (O_869,N_9606,N_9668);
xor UO_870 (O_870,N_9887,N_9656);
nor UO_871 (O_871,N_9849,N_9547);
and UO_872 (O_872,N_9900,N_9993);
xnor UO_873 (O_873,N_9883,N_9839);
nor UO_874 (O_874,N_9856,N_9726);
xnor UO_875 (O_875,N_9516,N_9929);
nor UO_876 (O_876,N_9770,N_9524);
xnor UO_877 (O_877,N_9860,N_9526);
or UO_878 (O_878,N_9531,N_9752);
xor UO_879 (O_879,N_9685,N_9615);
and UO_880 (O_880,N_9667,N_9970);
and UO_881 (O_881,N_9955,N_9506);
xnor UO_882 (O_882,N_9989,N_9639);
nand UO_883 (O_883,N_9756,N_9604);
and UO_884 (O_884,N_9806,N_9609);
and UO_885 (O_885,N_9815,N_9620);
xor UO_886 (O_886,N_9714,N_9694);
nor UO_887 (O_887,N_9794,N_9912);
or UO_888 (O_888,N_9858,N_9869);
and UO_889 (O_889,N_9605,N_9744);
xnor UO_890 (O_890,N_9868,N_9649);
or UO_891 (O_891,N_9787,N_9696);
nor UO_892 (O_892,N_9673,N_9510);
xnor UO_893 (O_893,N_9729,N_9975);
nand UO_894 (O_894,N_9812,N_9858);
or UO_895 (O_895,N_9557,N_9708);
nor UO_896 (O_896,N_9856,N_9572);
nor UO_897 (O_897,N_9894,N_9620);
and UO_898 (O_898,N_9839,N_9971);
and UO_899 (O_899,N_9537,N_9605);
and UO_900 (O_900,N_9663,N_9782);
nand UO_901 (O_901,N_9613,N_9576);
nor UO_902 (O_902,N_9944,N_9894);
and UO_903 (O_903,N_9949,N_9812);
or UO_904 (O_904,N_9820,N_9872);
and UO_905 (O_905,N_9744,N_9723);
or UO_906 (O_906,N_9599,N_9783);
and UO_907 (O_907,N_9637,N_9951);
nor UO_908 (O_908,N_9672,N_9618);
and UO_909 (O_909,N_9672,N_9673);
nor UO_910 (O_910,N_9909,N_9685);
or UO_911 (O_911,N_9704,N_9914);
nor UO_912 (O_912,N_9953,N_9831);
and UO_913 (O_913,N_9643,N_9824);
or UO_914 (O_914,N_9717,N_9508);
or UO_915 (O_915,N_9589,N_9739);
and UO_916 (O_916,N_9907,N_9964);
xor UO_917 (O_917,N_9750,N_9644);
xnor UO_918 (O_918,N_9741,N_9651);
nor UO_919 (O_919,N_9677,N_9635);
nand UO_920 (O_920,N_9978,N_9652);
or UO_921 (O_921,N_9809,N_9699);
nand UO_922 (O_922,N_9637,N_9649);
nand UO_923 (O_923,N_9505,N_9970);
or UO_924 (O_924,N_9549,N_9947);
nand UO_925 (O_925,N_9777,N_9789);
nor UO_926 (O_926,N_9720,N_9781);
nand UO_927 (O_927,N_9645,N_9835);
or UO_928 (O_928,N_9893,N_9679);
nor UO_929 (O_929,N_9957,N_9975);
nand UO_930 (O_930,N_9594,N_9923);
and UO_931 (O_931,N_9889,N_9644);
nor UO_932 (O_932,N_9785,N_9750);
and UO_933 (O_933,N_9778,N_9745);
or UO_934 (O_934,N_9825,N_9554);
nor UO_935 (O_935,N_9747,N_9676);
and UO_936 (O_936,N_9801,N_9665);
nand UO_937 (O_937,N_9911,N_9519);
and UO_938 (O_938,N_9948,N_9800);
xnor UO_939 (O_939,N_9616,N_9693);
and UO_940 (O_940,N_9796,N_9590);
nand UO_941 (O_941,N_9847,N_9738);
xnor UO_942 (O_942,N_9814,N_9905);
nor UO_943 (O_943,N_9785,N_9936);
xor UO_944 (O_944,N_9870,N_9519);
nand UO_945 (O_945,N_9571,N_9863);
xor UO_946 (O_946,N_9696,N_9887);
and UO_947 (O_947,N_9705,N_9775);
xor UO_948 (O_948,N_9643,N_9750);
xnor UO_949 (O_949,N_9933,N_9619);
nor UO_950 (O_950,N_9825,N_9958);
nand UO_951 (O_951,N_9662,N_9807);
and UO_952 (O_952,N_9609,N_9523);
nand UO_953 (O_953,N_9818,N_9855);
xnor UO_954 (O_954,N_9721,N_9865);
xor UO_955 (O_955,N_9517,N_9760);
xor UO_956 (O_956,N_9993,N_9762);
or UO_957 (O_957,N_9678,N_9939);
nor UO_958 (O_958,N_9989,N_9929);
xor UO_959 (O_959,N_9620,N_9737);
xor UO_960 (O_960,N_9758,N_9590);
or UO_961 (O_961,N_9822,N_9961);
or UO_962 (O_962,N_9984,N_9644);
nand UO_963 (O_963,N_9892,N_9815);
and UO_964 (O_964,N_9805,N_9532);
and UO_965 (O_965,N_9697,N_9787);
and UO_966 (O_966,N_9996,N_9572);
nand UO_967 (O_967,N_9801,N_9923);
nand UO_968 (O_968,N_9762,N_9661);
nor UO_969 (O_969,N_9661,N_9699);
and UO_970 (O_970,N_9952,N_9558);
xnor UO_971 (O_971,N_9545,N_9835);
nand UO_972 (O_972,N_9585,N_9901);
or UO_973 (O_973,N_9507,N_9799);
xor UO_974 (O_974,N_9747,N_9746);
nand UO_975 (O_975,N_9615,N_9583);
xnor UO_976 (O_976,N_9836,N_9532);
and UO_977 (O_977,N_9930,N_9861);
and UO_978 (O_978,N_9535,N_9678);
nand UO_979 (O_979,N_9962,N_9842);
nand UO_980 (O_980,N_9673,N_9598);
xnor UO_981 (O_981,N_9988,N_9594);
and UO_982 (O_982,N_9905,N_9542);
or UO_983 (O_983,N_9540,N_9995);
or UO_984 (O_984,N_9588,N_9750);
and UO_985 (O_985,N_9687,N_9645);
or UO_986 (O_986,N_9949,N_9573);
nand UO_987 (O_987,N_9912,N_9586);
xor UO_988 (O_988,N_9631,N_9601);
nor UO_989 (O_989,N_9615,N_9511);
and UO_990 (O_990,N_9524,N_9783);
nor UO_991 (O_991,N_9883,N_9911);
or UO_992 (O_992,N_9603,N_9844);
xnor UO_993 (O_993,N_9819,N_9706);
and UO_994 (O_994,N_9933,N_9577);
nor UO_995 (O_995,N_9996,N_9635);
or UO_996 (O_996,N_9561,N_9999);
nor UO_997 (O_997,N_9590,N_9501);
and UO_998 (O_998,N_9505,N_9898);
and UO_999 (O_999,N_9914,N_9613);
or UO_1000 (O_1000,N_9719,N_9753);
xnor UO_1001 (O_1001,N_9992,N_9532);
nor UO_1002 (O_1002,N_9688,N_9623);
or UO_1003 (O_1003,N_9960,N_9760);
and UO_1004 (O_1004,N_9676,N_9877);
xor UO_1005 (O_1005,N_9902,N_9519);
or UO_1006 (O_1006,N_9536,N_9991);
and UO_1007 (O_1007,N_9654,N_9879);
and UO_1008 (O_1008,N_9928,N_9932);
and UO_1009 (O_1009,N_9959,N_9726);
and UO_1010 (O_1010,N_9553,N_9665);
or UO_1011 (O_1011,N_9812,N_9595);
nor UO_1012 (O_1012,N_9895,N_9500);
and UO_1013 (O_1013,N_9504,N_9772);
nor UO_1014 (O_1014,N_9707,N_9714);
nand UO_1015 (O_1015,N_9648,N_9548);
xnor UO_1016 (O_1016,N_9722,N_9644);
nand UO_1017 (O_1017,N_9789,N_9873);
nand UO_1018 (O_1018,N_9565,N_9535);
or UO_1019 (O_1019,N_9726,N_9522);
xnor UO_1020 (O_1020,N_9728,N_9632);
or UO_1021 (O_1021,N_9768,N_9775);
or UO_1022 (O_1022,N_9699,N_9999);
nand UO_1023 (O_1023,N_9906,N_9984);
nor UO_1024 (O_1024,N_9977,N_9870);
nand UO_1025 (O_1025,N_9836,N_9582);
nand UO_1026 (O_1026,N_9585,N_9706);
nand UO_1027 (O_1027,N_9510,N_9901);
or UO_1028 (O_1028,N_9504,N_9791);
nand UO_1029 (O_1029,N_9715,N_9725);
xor UO_1030 (O_1030,N_9644,N_9736);
and UO_1031 (O_1031,N_9613,N_9608);
or UO_1032 (O_1032,N_9801,N_9750);
nand UO_1033 (O_1033,N_9599,N_9666);
xor UO_1034 (O_1034,N_9710,N_9653);
xnor UO_1035 (O_1035,N_9855,N_9865);
nand UO_1036 (O_1036,N_9761,N_9536);
nor UO_1037 (O_1037,N_9716,N_9526);
nand UO_1038 (O_1038,N_9773,N_9665);
nor UO_1039 (O_1039,N_9979,N_9760);
nand UO_1040 (O_1040,N_9703,N_9739);
nor UO_1041 (O_1041,N_9942,N_9709);
nand UO_1042 (O_1042,N_9527,N_9979);
and UO_1043 (O_1043,N_9729,N_9551);
nor UO_1044 (O_1044,N_9750,N_9730);
xnor UO_1045 (O_1045,N_9846,N_9750);
and UO_1046 (O_1046,N_9960,N_9702);
nor UO_1047 (O_1047,N_9667,N_9545);
nor UO_1048 (O_1048,N_9599,N_9831);
xor UO_1049 (O_1049,N_9974,N_9712);
xor UO_1050 (O_1050,N_9857,N_9994);
and UO_1051 (O_1051,N_9853,N_9702);
nand UO_1052 (O_1052,N_9756,N_9730);
and UO_1053 (O_1053,N_9975,N_9796);
nor UO_1054 (O_1054,N_9717,N_9856);
nor UO_1055 (O_1055,N_9830,N_9845);
xnor UO_1056 (O_1056,N_9800,N_9649);
and UO_1057 (O_1057,N_9839,N_9531);
or UO_1058 (O_1058,N_9884,N_9841);
nand UO_1059 (O_1059,N_9737,N_9788);
nand UO_1060 (O_1060,N_9982,N_9587);
or UO_1061 (O_1061,N_9731,N_9515);
or UO_1062 (O_1062,N_9513,N_9850);
nor UO_1063 (O_1063,N_9942,N_9904);
nand UO_1064 (O_1064,N_9715,N_9933);
nor UO_1065 (O_1065,N_9753,N_9863);
nand UO_1066 (O_1066,N_9515,N_9623);
nor UO_1067 (O_1067,N_9735,N_9704);
and UO_1068 (O_1068,N_9870,N_9748);
nor UO_1069 (O_1069,N_9662,N_9784);
nor UO_1070 (O_1070,N_9627,N_9653);
and UO_1071 (O_1071,N_9820,N_9878);
xor UO_1072 (O_1072,N_9507,N_9886);
and UO_1073 (O_1073,N_9884,N_9933);
nand UO_1074 (O_1074,N_9767,N_9788);
or UO_1075 (O_1075,N_9542,N_9782);
and UO_1076 (O_1076,N_9515,N_9558);
or UO_1077 (O_1077,N_9651,N_9594);
nand UO_1078 (O_1078,N_9816,N_9814);
nor UO_1079 (O_1079,N_9824,N_9918);
or UO_1080 (O_1080,N_9824,N_9963);
xnor UO_1081 (O_1081,N_9842,N_9874);
nand UO_1082 (O_1082,N_9778,N_9971);
nand UO_1083 (O_1083,N_9841,N_9856);
or UO_1084 (O_1084,N_9921,N_9638);
or UO_1085 (O_1085,N_9842,N_9865);
nor UO_1086 (O_1086,N_9896,N_9691);
nor UO_1087 (O_1087,N_9685,N_9773);
or UO_1088 (O_1088,N_9535,N_9872);
or UO_1089 (O_1089,N_9775,N_9580);
or UO_1090 (O_1090,N_9868,N_9615);
xor UO_1091 (O_1091,N_9742,N_9731);
nand UO_1092 (O_1092,N_9682,N_9588);
xnor UO_1093 (O_1093,N_9745,N_9518);
and UO_1094 (O_1094,N_9891,N_9756);
and UO_1095 (O_1095,N_9845,N_9923);
xnor UO_1096 (O_1096,N_9883,N_9616);
xor UO_1097 (O_1097,N_9541,N_9861);
nand UO_1098 (O_1098,N_9796,N_9919);
or UO_1099 (O_1099,N_9717,N_9641);
nor UO_1100 (O_1100,N_9798,N_9853);
xor UO_1101 (O_1101,N_9519,N_9705);
nand UO_1102 (O_1102,N_9922,N_9776);
nor UO_1103 (O_1103,N_9901,N_9932);
nand UO_1104 (O_1104,N_9707,N_9762);
xnor UO_1105 (O_1105,N_9932,N_9954);
xnor UO_1106 (O_1106,N_9762,N_9602);
or UO_1107 (O_1107,N_9547,N_9558);
xor UO_1108 (O_1108,N_9905,N_9719);
nor UO_1109 (O_1109,N_9709,N_9794);
nand UO_1110 (O_1110,N_9516,N_9875);
or UO_1111 (O_1111,N_9851,N_9704);
or UO_1112 (O_1112,N_9855,N_9510);
nor UO_1113 (O_1113,N_9965,N_9971);
xor UO_1114 (O_1114,N_9611,N_9516);
nor UO_1115 (O_1115,N_9517,N_9717);
or UO_1116 (O_1116,N_9593,N_9794);
xnor UO_1117 (O_1117,N_9669,N_9722);
nor UO_1118 (O_1118,N_9719,N_9709);
or UO_1119 (O_1119,N_9736,N_9609);
or UO_1120 (O_1120,N_9972,N_9767);
xnor UO_1121 (O_1121,N_9775,N_9553);
nor UO_1122 (O_1122,N_9762,N_9567);
nand UO_1123 (O_1123,N_9790,N_9581);
nor UO_1124 (O_1124,N_9804,N_9969);
xnor UO_1125 (O_1125,N_9590,N_9835);
or UO_1126 (O_1126,N_9728,N_9929);
and UO_1127 (O_1127,N_9953,N_9907);
nor UO_1128 (O_1128,N_9877,N_9841);
nor UO_1129 (O_1129,N_9938,N_9783);
nand UO_1130 (O_1130,N_9881,N_9616);
nand UO_1131 (O_1131,N_9794,N_9805);
and UO_1132 (O_1132,N_9790,N_9743);
nor UO_1133 (O_1133,N_9885,N_9688);
and UO_1134 (O_1134,N_9687,N_9502);
or UO_1135 (O_1135,N_9579,N_9921);
nand UO_1136 (O_1136,N_9723,N_9873);
xor UO_1137 (O_1137,N_9573,N_9581);
or UO_1138 (O_1138,N_9741,N_9900);
and UO_1139 (O_1139,N_9894,N_9998);
nand UO_1140 (O_1140,N_9576,N_9892);
or UO_1141 (O_1141,N_9651,N_9642);
and UO_1142 (O_1142,N_9693,N_9926);
xor UO_1143 (O_1143,N_9791,N_9638);
or UO_1144 (O_1144,N_9767,N_9529);
or UO_1145 (O_1145,N_9919,N_9573);
or UO_1146 (O_1146,N_9891,N_9545);
xnor UO_1147 (O_1147,N_9664,N_9623);
nor UO_1148 (O_1148,N_9975,N_9616);
xor UO_1149 (O_1149,N_9850,N_9771);
nand UO_1150 (O_1150,N_9600,N_9944);
or UO_1151 (O_1151,N_9633,N_9901);
or UO_1152 (O_1152,N_9564,N_9740);
nand UO_1153 (O_1153,N_9932,N_9612);
xnor UO_1154 (O_1154,N_9752,N_9589);
nor UO_1155 (O_1155,N_9867,N_9530);
nor UO_1156 (O_1156,N_9629,N_9525);
or UO_1157 (O_1157,N_9922,N_9862);
or UO_1158 (O_1158,N_9841,N_9801);
xor UO_1159 (O_1159,N_9949,N_9822);
or UO_1160 (O_1160,N_9593,N_9952);
xor UO_1161 (O_1161,N_9989,N_9895);
or UO_1162 (O_1162,N_9924,N_9757);
nand UO_1163 (O_1163,N_9805,N_9960);
nand UO_1164 (O_1164,N_9627,N_9664);
xor UO_1165 (O_1165,N_9889,N_9724);
nor UO_1166 (O_1166,N_9768,N_9905);
or UO_1167 (O_1167,N_9920,N_9985);
or UO_1168 (O_1168,N_9635,N_9689);
xnor UO_1169 (O_1169,N_9886,N_9544);
nor UO_1170 (O_1170,N_9892,N_9823);
nand UO_1171 (O_1171,N_9674,N_9934);
nor UO_1172 (O_1172,N_9670,N_9806);
or UO_1173 (O_1173,N_9635,N_9707);
nor UO_1174 (O_1174,N_9536,N_9808);
nor UO_1175 (O_1175,N_9601,N_9799);
nor UO_1176 (O_1176,N_9502,N_9549);
or UO_1177 (O_1177,N_9625,N_9681);
xnor UO_1178 (O_1178,N_9739,N_9697);
xor UO_1179 (O_1179,N_9918,N_9572);
nand UO_1180 (O_1180,N_9510,N_9592);
xor UO_1181 (O_1181,N_9650,N_9960);
nor UO_1182 (O_1182,N_9716,N_9758);
and UO_1183 (O_1183,N_9532,N_9612);
nand UO_1184 (O_1184,N_9712,N_9842);
nand UO_1185 (O_1185,N_9819,N_9758);
and UO_1186 (O_1186,N_9582,N_9714);
and UO_1187 (O_1187,N_9721,N_9994);
xnor UO_1188 (O_1188,N_9696,N_9725);
nand UO_1189 (O_1189,N_9626,N_9968);
nor UO_1190 (O_1190,N_9664,N_9674);
xnor UO_1191 (O_1191,N_9550,N_9543);
or UO_1192 (O_1192,N_9601,N_9537);
and UO_1193 (O_1193,N_9585,N_9671);
nand UO_1194 (O_1194,N_9935,N_9582);
or UO_1195 (O_1195,N_9570,N_9726);
or UO_1196 (O_1196,N_9789,N_9694);
nor UO_1197 (O_1197,N_9701,N_9827);
and UO_1198 (O_1198,N_9893,N_9813);
xor UO_1199 (O_1199,N_9534,N_9677);
nand UO_1200 (O_1200,N_9914,N_9523);
and UO_1201 (O_1201,N_9857,N_9903);
and UO_1202 (O_1202,N_9555,N_9664);
and UO_1203 (O_1203,N_9520,N_9938);
and UO_1204 (O_1204,N_9538,N_9832);
nand UO_1205 (O_1205,N_9569,N_9916);
and UO_1206 (O_1206,N_9769,N_9632);
or UO_1207 (O_1207,N_9569,N_9804);
xnor UO_1208 (O_1208,N_9543,N_9737);
and UO_1209 (O_1209,N_9719,N_9616);
xnor UO_1210 (O_1210,N_9612,N_9583);
or UO_1211 (O_1211,N_9867,N_9552);
and UO_1212 (O_1212,N_9621,N_9805);
and UO_1213 (O_1213,N_9511,N_9808);
xor UO_1214 (O_1214,N_9587,N_9731);
or UO_1215 (O_1215,N_9876,N_9726);
or UO_1216 (O_1216,N_9848,N_9689);
and UO_1217 (O_1217,N_9597,N_9788);
and UO_1218 (O_1218,N_9820,N_9775);
and UO_1219 (O_1219,N_9722,N_9975);
or UO_1220 (O_1220,N_9554,N_9978);
or UO_1221 (O_1221,N_9989,N_9885);
xor UO_1222 (O_1222,N_9733,N_9548);
nand UO_1223 (O_1223,N_9671,N_9884);
nor UO_1224 (O_1224,N_9538,N_9734);
and UO_1225 (O_1225,N_9744,N_9820);
and UO_1226 (O_1226,N_9730,N_9988);
nor UO_1227 (O_1227,N_9792,N_9795);
nor UO_1228 (O_1228,N_9718,N_9985);
xor UO_1229 (O_1229,N_9765,N_9669);
nor UO_1230 (O_1230,N_9691,N_9522);
nor UO_1231 (O_1231,N_9565,N_9530);
nor UO_1232 (O_1232,N_9650,N_9920);
and UO_1233 (O_1233,N_9849,N_9527);
and UO_1234 (O_1234,N_9914,N_9877);
nor UO_1235 (O_1235,N_9683,N_9706);
nand UO_1236 (O_1236,N_9630,N_9940);
xor UO_1237 (O_1237,N_9652,N_9519);
and UO_1238 (O_1238,N_9854,N_9586);
or UO_1239 (O_1239,N_9687,N_9855);
or UO_1240 (O_1240,N_9581,N_9862);
or UO_1241 (O_1241,N_9523,N_9957);
nand UO_1242 (O_1242,N_9827,N_9843);
xnor UO_1243 (O_1243,N_9770,N_9877);
nand UO_1244 (O_1244,N_9936,N_9767);
or UO_1245 (O_1245,N_9994,N_9695);
nand UO_1246 (O_1246,N_9862,N_9827);
xor UO_1247 (O_1247,N_9768,N_9719);
and UO_1248 (O_1248,N_9642,N_9674);
nand UO_1249 (O_1249,N_9667,N_9619);
nor UO_1250 (O_1250,N_9795,N_9561);
or UO_1251 (O_1251,N_9720,N_9863);
or UO_1252 (O_1252,N_9713,N_9875);
nand UO_1253 (O_1253,N_9566,N_9575);
and UO_1254 (O_1254,N_9552,N_9897);
xnor UO_1255 (O_1255,N_9687,N_9674);
xnor UO_1256 (O_1256,N_9641,N_9887);
and UO_1257 (O_1257,N_9753,N_9736);
or UO_1258 (O_1258,N_9840,N_9605);
or UO_1259 (O_1259,N_9637,N_9855);
or UO_1260 (O_1260,N_9560,N_9961);
nor UO_1261 (O_1261,N_9523,N_9783);
nand UO_1262 (O_1262,N_9542,N_9960);
and UO_1263 (O_1263,N_9699,N_9820);
and UO_1264 (O_1264,N_9767,N_9967);
and UO_1265 (O_1265,N_9738,N_9710);
nor UO_1266 (O_1266,N_9737,N_9842);
and UO_1267 (O_1267,N_9779,N_9998);
and UO_1268 (O_1268,N_9626,N_9732);
or UO_1269 (O_1269,N_9972,N_9800);
xor UO_1270 (O_1270,N_9612,N_9520);
and UO_1271 (O_1271,N_9816,N_9566);
and UO_1272 (O_1272,N_9983,N_9589);
xor UO_1273 (O_1273,N_9878,N_9559);
and UO_1274 (O_1274,N_9503,N_9880);
nor UO_1275 (O_1275,N_9528,N_9770);
xor UO_1276 (O_1276,N_9842,N_9955);
nor UO_1277 (O_1277,N_9744,N_9703);
nand UO_1278 (O_1278,N_9618,N_9548);
xnor UO_1279 (O_1279,N_9942,N_9986);
and UO_1280 (O_1280,N_9846,N_9541);
nor UO_1281 (O_1281,N_9830,N_9516);
nand UO_1282 (O_1282,N_9537,N_9561);
nand UO_1283 (O_1283,N_9767,N_9756);
xor UO_1284 (O_1284,N_9630,N_9752);
or UO_1285 (O_1285,N_9586,N_9616);
nor UO_1286 (O_1286,N_9626,N_9548);
and UO_1287 (O_1287,N_9921,N_9814);
or UO_1288 (O_1288,N_9878,N_9923);
nor UO_1289 (O_1289,N_9622,N_9952);
nor UO_1290 (O_1290,N_9911,N_9772);
xnor UO_1291 (O_1291,N_9650,N_9819);
or UO_1292 (O_1292,N_9683,N_9615);
or UO_1293 (O_1293,N_9844,N_9791);
and UO_1294 (O_1294,N_9655,N_9665);
or UO_1295 (O_1295,N_9623,N_9674);
xnor UO_1296 (O_1296,N_9725,N_9698);
nor UO_1297 (O_1297,N_9670,N_9819);
nor UO_1298 (O_1298,N_9989,N_9875);
xnor UO_1299 (O_1299,N_9745,N_9957);
or UO_1300 (O_1300,N_9827,N_9795);
nand UO_1301 (O_1301,N_9623,N_9730);
nand UO_1302 (O_1302,N_9710,N_9939);
nor UO_1303 (O_1303,N_9788,N_9662);
and UO_1304 (O_1304,N_9730,N_9655);
nand UO_1305 (O_1305,N_9660,N_9750);
nand UO_1306 (O_1306,N_9934,N_9572);
nand UO_1307 (O_1307,N_9687,N_9536);
and UO_1308 (O_1308,N_9783,N_9760);
and UO_1309 (O_1309,N_9992,N_9520);
xnor UO_1310 (O_1310,N_9746,N_9667);
nand UO_1311 (O_1311,N_9934,N_9914);
and UO_1312 (O_1312,N_9868,N_9946);
or UO_1313 (O_1313,N_9784,N_9865);
xnor UO_1314 (O_1314,N_9702,N_9931);
nand UO_1315 (O_1315,N_9862,N_9864);
xnor UO_1316 (O_1316,N_9617,N_9837);
xnor UO_1317 (O_1317,N_9988,N_9842);
xnor UO_1318 (O_1318,N_9582,N_9914);
nor UO_1319 (O_1319,N_9824,N_9768);
nor UO_1320 (O_1320,N_9994,N_9733);
xor UO_1321 (O_1321,N_9696,N_9847);
or UO_1322 (O_1322,N_9677,N_9870);
or UO_1323 (O_1323,N_9707,N_9615);
nor UO_1324 (O_1324,N_9581,N_9724);
or UO_1325 (O_1325,N_9981,N_9518);
xor UO_1326 (O_1326,N_9868,N_9530);
nor UO_1327 (O_1327,N_9587,N_9890);
nand UO_1328 (O_1328,N_9567,N_9791);
nor UO_1329 (O_1329,N_9615,N_9846);
nand UO_1330 (O_1330,N_9567,N_9880);
and UO_1331 (O_1331,N_9600,N_9686);
or UO_1332 (O_1332,N_9719,N_9530);
and UO_1333 (O_1333,N_9898,N_9695);
nor UO_1334 (O_1334,N_9759,N_9901);
or UO_1335 (O_1335,N_9892,N_9832);
nor UO_1336 (O_1336,N_9940,N_9847);
nand UO_1337 (O_1337,N_9963,N_9611);
or UO_1338 (O_1338,N_9568,N_9775);
or UO_1339 (O_1339,N_9854,N_9805);
xnor UO_1340 (O_1340,N_9632,N_9791);
nor UO_1341 (O_1341,N_9591,N_9802);
and UO_1342 (O_1342,N_9750,N_9778);
or UO_1343 (O_1343,N_9567,N_9696);
xnor UO_1344 (O_1344,N_9556,N_9695);
xnor UO_1345 (O_1345,N_9879,N_9805);
nor UO_1346 (O_1346,N_9587,N_9513);
or UO_1347 (O_1347,N_9669,N_9504);
nor UO_1348 (O_1348,N_9789,N_9803);
and UO_1349 (O_1349,N_9622,N_9640);
xor UO_1350 (O_1350,N_9581,N_9934);
nor UO_1351 (O_1351,N_9674,N_9545);
or UO_1352 (O_1352,N_9740,N_9991);
nand UO_1353 (O_1353,N_9624,N_9672);
or UO_1354 (O_1354,N_9570,N_9604);
xor UO_1355 (O_1355,N_9745,N_9947);
nand UO_1356 (O_1356,N_9515,N_9594);
nand UO_1357 (O_1357,N_9811,N_9620);
nand UO_1358 (O_1358,N_9760,N_9660);
and UO_1359 (O_1359,N_9727,N_9776);
xnor UO_1360 (O_1360,N_9969,N_9904);
nor UO_1361 (O_1361,N_9619,N_9797);
xnor UO_1362 (O_1362,N_9752,N_9615);
nor UO_1363 (O_1363,N_9955,N_9960);
xnor UO_1364 (O_1364,N_9914,N_9930);
or UO_1365 (O_1365,N_9746,N_9653);
xnor UO_1366 (O_1366,N_9556,N_9666);
nand UO_1367 (O_1367,N_9886,N_9946);
xor UO_1368 (O_1368,N_9907,N_9550);
and UO_1369 (O_1369,N_9541,N_9638);
nand UO_1370 (O_1370,N_9922,N_9850);
xor UO_1371 (O_1371,N_9600,N_9527);
or UO_1372 (O_1372,N_9588,N_9570);
nand UO_1373 (O_1373,N_9693,N_9787);
or UO_1374 (O_1374,N_9573,N_9673);
nor UO_1375 (O_1375,N_9612,N_9581);
or UO_1376 (O_1376,N_9624,N_9644);
nor UO_1377 (O_1377,N_9793,N_9504);
nor UO_1378 (O_1378,N_9888,N_9552);
nor UO_1379 (O_1379,N_9661,N_9753);
nand UO_1380 (O_1380,N_9569,N_9611);
or UO_1381 (O_1381,N_9897,N_9779);
nor UO_1382 (O_1382,N_9546,N_9890);
xor UO_1383 (O_1383,N_9831,N_9948);
xnor UO_1384 (O_1384,N_9933,N_9910);
xor UO_1385 (O_1385,N_9888,N_9909);
and UO_1386 (O_1386,N_9687,N_9575);
or UO_1387 (O_1387,N_9885,N_9819);
xor UO_1388 (O_1388,N_9737,N_9847);
nand UO_1389 (O_1389,N_9591,N_9894);
nand UO_1390 (O_1390,N_9560,N_9954);
nor UO_1391 (O_1391,N_9990,N_9656);
xnor UO_1392 (O_1392,N_9979,N_9592);
xor UO_1393 (O_1393,N_9669,N_9638);
nand UO_1394 (O_1394,N_9954,N_9626);
xor UO_1395 (O_1395,N_9980,N_9813);
nand UO_1396 (O_1396,N_9563,N_9995);
and UO_1397 (O_1397,N_9893,N_9844);
nor UO_1398 (O_1398,N_9932,N_9843);
nand UO_1399 (O_1399,N_9833,N_9734);
and UO_1400 (O_1400,N_9955,N_9969);
nand UO_1401 (O_1401,N_9927,N_9904);
and UO_1402 (O_1402,N_9719,N_9576);
or UO_1403 (O_1403,N_9695,N_9935);
nor UO_1404 (O_1404,N_9659,N_9753);
nand UO_1405 (O_1405,N_9611,N_9521);
xor UO_1406 (O_1406,N_9598,N_9969);
or UO_1407 (O_1407,N_9570,N_9831);
nor UO_1408 (O_1408,N_9588,N_9579);
nor UO_1409 (O_1409,N_9999,N_9766);
or UO_1410 (O_1410,N_9719,N_9912);
and UO_1411 (O_1411,N_9581,N_9732);
xor UO_1412 (O_1412,N_9528,N_9674);
nand UO_1413 (O_1413,N_9532,N_9919);
xnor UO_1414 (O_1414,N_9800,N_9856);
or UO_1415 (O_1415,N_9598,N_9648);
nor UO_1416 (O_1416,N_9945,N_9569);
and UO_1417 (O_1417,N_9755,N_9848);
nand UO_1418 (O_1418,N_9782,N_9757);
or UO_1419 (O_1419,N_9747,N_9729);
nor UO_1420 (O_1420,N_9651,N_9550);
xor UO_1421 (O_1421,N_9856,N_9794);
nand UO_1422 (O_1422,N_9600,N_9570);
xor UO_1423 (O_1423,N_9934,N_9556);
xnor UO_1424 (O_1424,N_9801,N_9649);
and UO_1425 (O_1425,N_9768,N_9969);
nand UO_1426 (O_1426,N_9906,N_9564);
nor UO_1427 (O_1427,N_9750,N_9547);
nand UO_1428 (O_1428,N_9603,N_9837);
xor UO_1429 (O_1429,N_9601,N_9620);
nor UO_1430 (O_1430,N_9984,N_9905);
xnor UO_1431 (O_1431,N_9861,N_9842);
nand UO_1432 (O_1432,N_9962,N_9901);
nand UO_1433 (O_1433,N_9565,N_9603);
xnor UO_1434 (O_1434,N_9845,N_9546);
nand UO_1435 (O_1435,N_9830,N_9731);
nor UO_1436 (O_1436,N_9787,N_9819);
and UO_1437 (O_1437,N_9941,N_9967);
nand UO_1438 (O_1438,N_9595,N_9942);
or UO_1439 (O_1439,N_9916,N_9557);
nand UO_1440 (O_1440,N_9721,N_9898);
nor UO_1441 (O_1441,N_9821,N_9959);
xor UO_1442 (O_1442,N_9642,N_9567);
and UO_1443 (O_1443,N_9745,N_9927);
nor UO_1444 (O_1444,N_9853,N_9630);
xor UO_1445 (O_1445,N_9530,N_9998);
nor UO_1446 (O_1446,N_9998,N_9839);
and UO_1447 (O_1447,N_9960,N_9771);
or UO_1448 (O_1448,N_9990,N_9530);
and UO_1449 (O_1449,N_9664,N_9948);
and UO_1450 (O_1450,N_9850,N_9538);
nor UO_1451 (O_1451,N_9634,N_9540);
nor UO_1452 (O_1452,N_9909,N_9557);
and UO_1453 (O_1453,N_9628,N_9663);
nor UO_1454 (O_1454,N_9776,N_9671);
nand UO_1455 (O_1455,N_9801,N_9703);
and UO_1456 (O_1456,N_9626,N_9643);
and UO_1457 (O_1457,N_9681,N_9685);
and UO_1458 (O_1458,N_9587,N_9690);
nor UO_1459 (O_1459,N_9826,N_9849);
or UO_1460 (O_1460,N_9976,N_9741);
xor UO_1461 (O_1461,N_9842,N_9630);
nand UO_1462 (O_1462,N_9872,N_9645);
and UO_1463 (O_1463,N_9702,N_9723);
and UO_1464 (O_1464,N_9937,N_9982);
and UO_1465 (O_1465,N_9586,N_9683);
nor UO_1466 (O_1466,N_9543,N_9517);
xnor UO_1467 (O_1467,N_9503,N_9846);
and UO_1468 (O_1468,N_9721,N_9822);
or UO_1469 (O_1469,N_9868,N_9981);
nor UO_1470 (O_1470,N_9853,N_9592);
or UO_1471 (O_1471,N_9551,N_9663);
or UO_1472 (O_1472,N_9636,N_9754);
xor UO_1473 (O_1473,N_9509,N_9832);
or UO_1474 (O_1474,N_9765,N_9884);
nand UO_1475 (O_1475,N_9782,N_9621);
or UO_1476 (O_1476,N_9852,N_9757);
nand UO_1477 (O_1477,N_9947,N_9562);
xor UO_1478 (O_1478,N_9530,N_9619);
nand UO_1479 (O_1479,N_9683,N_9541);
nor UO_1480 (O_1480,N_9993,N_9598);
and UO_1481 (O_1481,N_9569,N_9581);
nand UO_1482 (O_1482,N_9801,N_9582);
xor UO_1483 (O_1483,N_9616,N_9524);
xor UO_1484 (O_1484,N_9537,N_9894);
nor UO_1485 (O_1485,N_9503,N_9968);
nand UO_1486 (O_1486,N_9548,N_9950);
and UO_1487 (O_1487,N_9640,N_9637);
nand UO_1488 (O_1488,N_9630,N_9796);
xnor UO_1489 (O_1489,N_9740,N_9752);
and UO_1490 (O_1490,N_9602,N_9513);
nand UO_1491 (O_1491,N_9952,N_9984);
nor UO_1492 (O_1492,N_9619,N_9650);
nor UO_1493 (O_1493,N_9903,N_9987);
and UO_1494 (O_1494,N_9903,N_9655);
xor UO_1495 (O_1495,N_9682,N_9655);
or UO_1496 (O_1496,N_9943,N_9979);
nor UO_1497 (O_1497,N_9964,N_9782);
nand UO_1498 (O_1498,N_9702,N_9982);
nand UO_1499 (O_1499,N_9833,N_9812);
endmodule