module basic_500_3000_500_3_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_255,In_335);
nand U1 (N_1,In_221,In_434);
or U2 (N_2,In_382,In_58);
nand U3 (N_3,In_177,In_325);
nor U4 (N_4,In_152,In_431);
or U5 (N_5,In_244,In_373);
nor U6 (N_6,In_27,In_31);
and U7 (N_7,In_486,In_481);
nand U8 (N_8,In_298,In_74);
nand U9 (N_9,In_277,In_406);
or U10 (N_10,In_347,In_357);
or U11 (N_11,In_490,In_168);
nor U12 (N_12,In_243,In_198);
nor U13 (N_13,In_127,In_404);
and U14 (N_14,In_136,In_82);
or U15 (N_15,In_268,In_392);
nand U16 (N_16,In_116,In_11);
and U17 (N_17,In_185,In_409);
and U18 (N_18,In_395,In_300);
or U19 (N_19,In_324,In_179);
or U20 (N_20,In_160,In_366);
or U21 (N_21,In_149,In_446);
nor U22 (N_22,In_259,In_454);
or U23 (N_23,In_414,In_142);
nand U24 (N_24,In_197,In_202);
nand U25 (N_25,In_350,In_119);
and U26 (N_26,In_310,In_263);
nor U27 (N_27,In_181,In_48);
or U28 (N_28,In_172,In_30);
nor U29 (N_29,In_320,In_89);
nand U30 (N_30,In_76,In_187);
and U31 (N_31,In_458,In_412);
xnor U32 (N_32,In_326,In_276);
nand U33 (N_33,In_493,In_1);
nor U34 (N_34,In_459,In_191);
nor U35 (N_35,In_45,In_162);
nand U36 (N_36,In_466,In_489);
or U37 (N_37,In_212,In_75);
nor U38 (N_38,In_90,In_6);
and U39 (N_39,In_380,In_62);
and U40 (N_40,In_261,In_230);
and U41 (N_41,In_102,In_470);
nand U42 (N_42,In_43,In_78);
or U43 (N_43,In_308,In_445);
nand U44 (N_44,In_460,In_497);
nand U45 (N_45,In_296,In_448);
nand U46 (N_46,In_384,In_487);
nand U47 (N_47,In_118,In_484);
and U48 (N_48,In_239,In_87);
nor U49 (N_49,In_428,In_148);
nand U50 (N_50,In_229,In_456);
and U51 (N_51,In_217,In_291);
nor U52 (N_52,In_478,In_423);
or U53 (N_53,In_360,In_196);
and U54 (N_54,In_389,In_402);
nor U55 (N_55,In_67,In_264);
nor U56 (N_56,In_473,In_376);
and U57 (N_57,In_361,In_238);
or U58 (N_58,In_323,In_139);
nand U59 (N_59,In_124,In_88);
nor U60 (N_60,In_132,In_429);
nand U61 (N_61,In_169,In_189);
nor U62 (N_62,In_223,In_39);
nor U63 (N_63,In_386,In_306);
nor U64 (N_64,In_122,In_247);
nand U65 (N_65,In_271,In_292);
nor U66 (N_66,In_248,In_467);
nand U67 (N_67,In_301,In_73);
nor U68 (N_68,In_104,In_42);
or U69 (N_69,In_273,In_170);
or U70 (N_70,In_343,In_495);
nor U71 (N_71,In_345,In_387);
or U72 (N_72,In_200,In_237);
nand U73 (N_73,In_284,In_57);
or U74 (N_74,In_205,In_46);
and U75 (N_75,In_64,In_128);
or U76 (N_76,In_141,In_208);
nor U77 (N_77,In_26,In_265);
and U78 (N_78,In_444,In_316);
or U79 (N_79,In_34,In_77);
and U80 (N_80,In_313,In_0);
and U81 (N_81,In_61,In_130);
nor U82 (N_82,In_391,In_307);
nand U83 (N_83,In_84,In_279);
and U84 (N_84,In_354,In_447);
nand U85 (N_85,In_54,In_146);
nand U86 (N_86,In_385,In_93);
and U87 (N_87,In_358,In_156);
nand U88 (N_88,In_476,In_35);
nand U89 (N_89,In_66,In_13);
or U90 (N_90,In_182,In_443);
and U91 (N_91,In_59,In_186);
nor U92 (N_92,In_234,In_91);
or U93 (N_93,In_214,In_426);
and U94 (N_94,In_477,In_192);
nand U95 (N_95,In_419,In_299);
or U96 (N_96,In_125,In_397);
nand U97 (N_97,In_110,In_94);
nor U98 (N_98,In_209,In_219);
nor U99 (N_99,In_143,In_85);
and U100 (N_100,In_480,In_38);
and U101 (N_101,In_372,In_96);
or U102 (N_102,In_338,In_437);
nand U103 (N_103,In_349,In_44);
and U104 (N_104,In_280,In_52);
nor U105 (N_105,In_494,In_126);
nand U106 (N_106,In_245,In_282);
nand U107 (N_107,In_364,In_346);
nor U108 (N_108,In_450,In_413);
and U109 (N_109,In_368,In_289);
and U110 (N_110,In_251,In_336);
or U111 (N_111,In_131,In_331);
nor U112 (N_112,In_329,In_287);
or U113 (N_113,In_457,In_482);
and U114 (N_114,In_113,In_311);
nand U115 (N_115,In_36,In_314);
nor U116 (N_116,In_328,In_194);
and U117 (N_117,In_496,In_23);
nand U118 (N_118,In_150,In_309);
nor U119 (N_119,In_449,In_252);
nor U120 (N_120,In_28,In_138);
or U121 (N_121,In_40,In_33);
and U122 (N_122,In_474,In_112);
or U123 (N_123,In_218,In_63);
or U124 (N_124,In_2,In_163);
nor U125 (N_125,In_105,In_108);
or U126 (N_126,In_86,In_72);
or U127 (N_127,In_180,In_32);
and U128 (N_128,In_363,In_195);
or U129 (N_129,In_233,In_269);
or U130 (N_130,In_499,In_322);
nor U131 (N_131,In_302,In_398);
or U132 (N_132,In_117,In_107);
nor U133 (N_133,In_415,In_220);
and U134 (N_134,In_461,In_81);
nand U135 (N_135,In_272,In_374);
or U136 (N_136,In_332,In_103);
nor U137 (N_137,In_403,In_190);
or U138 (N_138,In_422,In_10);
nand U139 (N_139,In_383,In_256);
nand U140 (N_140,In_79,In_266);
nor U141 (N_141,In_158,In_370);
nand U142 (N_142,In_174,In_240);
or U143 (N_143,In_5,In_381);
nand U144 (N_144,In_418,In_334);
nor U145 (N_145,In_297,In_399);
nor U146 (N_146,In_135,In_153);
nand U147 (N_147,In_16,In_49);
nand U148 (N_148,In_140,In_222);
nand U149 (N_149,In_9,In_216);
and U150 (N_150,In_455,In_465);
nand U151 (N_151,In_441,In_420);
and U152 (N_152,In_207,In_92);
nand U153 (N_153,In_410,In_171);
nor U154 (N_154,In_405,In_155);
or U155 (N_155,In_283,In_421);
and U156 (N_156,In_442,In_359);
nor U157 (N_157,In_111,In_356);
nand U158 (N_158,In_211,In_451);
or U159 (N_159,In_351,In_417);
and U160 (N_160,In_120,In_365);
and U161 (N_161,In_123,In_471);
nor U162 (N_162,In_249,In_427);
xnor U163 (N_163,In_121,In_167);
and U164 (N_164,In_161,In_452);
nor U165 (N_165,In_462,In_388);
nand U166 (N_166,In_101,In_362);
nor U167 (N_167,In_498,In_151);
nor U168 (N_168,In_137,In_83);
and U169 (N_169,In_232,In_109);
or U170 (N_170,In_15,In_281);
nand U171 (N_171,In_488,In_253);
nor U172 (N_172,In_106,In_201);
nand U173 (N_173,In_193,In_400);
nor U174 (N_174,In_340,In_20);
or U175 (N_175,In_318,In_491);
nor U176 (N_176,In_225,In_468);
nor U177 (N_177,In_242,In_71);
nand U178 (N_178,In_18,In_394);
nand U179 (N_179,In_355,In_213);
nand U180 (N_180,In_275,In_188);
nor U181 (N_181,In_348,In_258);
xor U182 (N_182,In_257,In_164);
nand U183 (N_183,In_432,In_293);
and U184 (N_184,In_353,In_25);
nor U185 (N_185,In_260,In_50);
nor U186 (N_186,In_3,In_166);
or U187 (N_187,In_47,In_436);
or U188 (N_188,In_262,In_184);
nand U189 (N_189,In_479,In_80);
nor U190 (N_190,In_285,In_485);
or U191 (N_191,In_440,In_341);
and U192 (N_192,In_492,In_330);
nand U193 (N_193,In_319,In_159);
or U194 (N_194,In_250,In_235);
nor U195 (N_195,In_37,In_100);
or U196 (N_196,In_288,In_210);
nor U197 (N_197,In_472,In_165);
nand U198 (N_198,In_8,In_65);
nor U199 (N_199,In_99,In_4);
or U200 (N_200,In_241,In_371);
or U201 (N_201,In_295,In_367);
and U202 (N_202,In_176,In_215);
and U203 (N_203,In_224,In_317);
and U204 (N_204,In_227,In_41);
nand U205 (N_205,In_157,In_294);
xnor U206 (N_206,In_430,In_199);
nor U207 (N_207,In_401,In_147);
nand U208 (N_208,In_134,In_393);
and U209 (N_209,In_274,In_464);
or U210 (N_210,In_115,In_453);
and U211 (N_211,In_12,In_321);
or U212 (N_212,In_145,In_439);
nor U213 (N_213,In_144,In_270);
or U214 (N_214,In_315,In_483);
nand U215 (N_215,In_175,In_14);
and U216 (N_216,In_203,In_438);
or U217 (N_217,In_407,In_411);
or U218 (N_218,In_154,In_425);
nor U219 (N_219,In_377,In_7);
or U220 (N_220,In_246,In_408);
and U221 (N_221,In_68,In_342);
xnor U222 (N_222,In_95,In_305);
nor U223 (N_223,In_133,In_396);
nand U224 (N_224,In_55,In_344);
or U225 (N_225,In_333,In_369);
and U226 (N_226,In_339,In_183);
or U227 (N_227,In_24,In_228);
and U228 (N_228,In_278,In_51);
and U229 (N_229,In_114,In_204);
and U230 (N_230,In_60,In_375);
nand U231 (N_231,In_390,In_327);
and U232 (N_232,In_475,In_352);
xor U233 (N_233,In_416,In_56);
or U234 (N_234,In_463,In_433);
nor U235 (N_235,In_129,In_231);
or U236 (N_236,In_98,In_337);
and U237 (N_237,In_290,In_424);
and U238 (N_238,In_178,In_19);
nand U239 (N_239,In_267,In_286);
nor U240 (N_240,In_70,In_69);
or U241 (N_241,In_21,In_97);
nor U242 (N_242,In_312,In_206);
or U243 (N_243,In_435,In_304);
and U244 (N_244,In_254,In_53);
nor U245 (N_245,In_22,In_29);
nand U246 (N_246,In_226,In_378);
nand U247 (N_247,In_469,In_17);
nand U248 (N_248,In_303,In_236);
or U249 (N_249,In_379,In_173);
nor U250 (N_250,In_394,In_416);
nor U251 (N_251,In_158,In_419);
nor U252 (N_252,In_112,In_201);
xor U253 (N_253,In_64,In_410);
or U254 (N_254,In_341,In_165);
and U255 (N_255,In_205,In_472);
nor U256 (N_256,In_48,In_246);
nor U257 (N_257,In_442,In_325);
or U258 (N_258,In_255,In_159);
nand U259 (N_259,In_379,In_259);
and U260 (N_260,In_412,In_355);
nor U261 (N_261,In_242,In_359);
nand U262 (N_262,In_271,In_101);
nand U263 (N_263,In_392,In_478);
and U264 (N_264,In_499,In_65);
nor U265 (N_265,In_296,In_469);
and U266 (N_266,In_416,In_134);
or U267 (N_267,In_99,In_286);
and U268 (N_268,In_481,In_70);
or U269 (N_269,In_17,In_157);
and U270 (N_270,In_31,In_148);
nor U271 (N_271,In_154,In_358);
nand U272 (N_272,In_285,In_53);
nor U273 (N_273,In_391,In_358);
or U274 (N_274,In_339,In_357);
nand U275 (N_275,In_320,In_148);
nand U276 (N_276,In_399,In_167);
or U277 (N_277,In_387,In_484);
nand U278 (N_278,In_420,In_293);
nand U279 (N_279,In_461,In_104);
or U280 (N_280,In_345,In_97);
nand U281 (N_281,In_32,In_94);
and U282 (N_282,In_100,In_6);
nand U283 (N_283,In_411,In_458);
nor U284 (N_284,In_0,In_31);
nand U285 (N_285,In_163,In_166);
nand U286 (N_286,In_189,In_2);
nand U287 (N_287,In_446,In_432);
nor U288 (N_288,In_185,In_418);
or U289 (N_289,In_286,In_312);
and U290 (N_290,In_433,In_400);
nand U291 (N_291,In_252,In_8);
nand U292 (N_292,In_462,In_5);
and U293 (N_293,In_58,In_173);
nand U294 (N_294,In_439,In_141);
and U295 (N_295,In_444,In_325);
nand U296 (N_296,In_247,In_354);
nor U297 (N_297,In_37,In_15);
or U298 (N_298,In_342,In_246);
or U299 (N_299,In_201,In_432);
and U300 (N_300,In_125,In_121);
nor U301 (N_301,In_318,In_288);
and U302 (N_302,In_413,In_429);
nor U303 (N_303,In_390,In_172);
and U304 (N_304,In_83,In_32);
and U305 (N_305,In_98,In_129);
nor U306 (N_306,In_208,In_0);
and U307 (N_307,In_132,In_125);
or U308 (N_308,In_267,In_5);
nand U309 (N_309,In_206,In_239);
or U310 (N_310,In_295,In_14);
and U311 (N_311,In_28,In_32);
nand U312 (N_312,In_305,In_289);
nor U313 (N_313,In_179,In_223);
nor U314 (N_314,In_229,In_216);
or U315 (N_315,In_216,In_210);
nor U316 (N_316,In_101,In_84);
and U317 (N_317,In_424,In_358);
and U318 (N_318,In_348,In_134);
nand U319 (N_319,In_283,In_328);
or U320 (N_320,In_313,In_365);
and U321 (N_321,In_115,In_39);
or U322 (N_322,In_175,In_39);
nand U323 (N_323,In_223,In_464);
nand U324 (N_324,In_206,In_297);
and U325 (N_325,In_134,In_38);
nand U326 (N_326,In_448,In_479);
xnor U327 (N_327,In_253,In_402);
and U328 (N_328,In_447,In_438);
nand U329 (N_329,In_419,In_342);
nand U330 (N_330,In_280,In_98);
nor U331 (N_331,In_182,In_352);
and U332 (N_332,In_313,In_355);
nor U333 (N_333,In_31,In_270);
nor U334 (N_334,In_124,In_28);
and U335 (N_335,In_300,In_67);
nand U336 (N_336,In_111,In_351);
and U337 (N_337,In_253,In_351);
or U338 (N_338,In_390,In_370);
nor U339 (N_339,In_210,In_444);
nor U340 (N_340,In_468,In_58);
nand U341 (N_341,In_160,In_131);
nand U342 (N_342,In_36,In_33);
nand U343 (N_343,In_5,In_297);
nor U344 (N_344,In_50,In_291);
nor U345 (N_345,In_98,In_17);
nor U346 (N_346,In_260,In_400);
nand U347 (N_347,In_242,In_121);
nand U348 (N_348,In_213,In_95);
nand U349 (N_349,In_30,In_274);
nor U350 (N_350,In_127,In_469);
nand U351 (N_351,In_444,In_430);
and U352 (N_352,In_123,In_435);
and U353 (N_353,In_335,In_218);
and U354 (N_354,In_441,In_105);
and U355 (N_355,In_293,In_377);
nand U356 (N_356,In_338,In_157);
and U357 (N_357,In_177,In_479);
nor U358 (N_358,In_95,In_373);
nand U359 (N_359,In_495,In_28);
nor U360 (N_360,In_447,In_389);
and U361 (N_361,In_96,In_67);
nand U362 (N_362,In_325,In_132);
nor U363 (N_363,In_199,In_490);
xor U364 (N_364,In_324,In_370);
nand U365 (N_365,In_341,In_187);
and U366 (N_366,In_422,In_345);
nor U367 (N_367,In_47,In_41);
or U368 (N_368,In_453,In_102);
and U369 (N_369,In_66,In_369);
and U370 (N_370,In_382,In_178);
nand U371 (N_371,In_54,In_210);
nand U372 (N_372,In_73,In_280);
or U373 (N_373,In_412,In_280);
nand U374 (N_374,In_89,In_271);
and U375 (N_375,In_416,In_352);
nor U376 (N_376,In_174,In_56);
or U377 (N_377,In_9,In_272);
nand U378 (N_378,In_246,In_450);
and U379 (N_379,In_118,In_219);
nor U380 (N_380,In_429,In_207);
nand U381 (N_381,In_51,In_19);
nand U382 (N_382,In_438,In_112);
and U383 (N_383,In_146,In_496);
or U384 (N_384,In_228,In_388);
nand U385 (N_385,In_181,In_299);
nand U386 (N_386,In_188,In_238);
and U387 (N_387,In_270,In_244);
nor U388 (N_388,In_354,In_19);
nand U389 (N_389,In_405,In_71);
nor U390 (N_390,In_19,In_205);
nand U391 (N_391,In_202,In_480);
and U392 (N_392,In_77,In_46);
and U393 (N_393,In_448,In_22);
or U394 (N_394,In_411,In_410);
nor U395 (N_395,In_366,In_121);
or U396 (N_396,In_319,In_72);
and U397 (N_397,In_71,In_399);
or U398 (N_398,In_493,In_270);
nand U399 (N_399,In_133,In_426);
nand U400 (N_400,In_116,In_102);
and U401 (N_401,In_301,In_87);
and U402 (N_402,In_61,In_364);
nand U403 (N_403,In_80,In_306);
or U404 (N_404,In_155,In_168);
nand U405 (N_405,In_13,In_72);
nor U406 (N_406,In_86,In_283);
nand U407 (N_407,In_180,In_119);
or U408 (N_408,In_143,In_378);
or U409 (N_409,In_190,In_411);
nand U410 (N_410,In_82,In_354);
and U411 (N_411,In_321,In_329);
nor U412 (N_412,In_71,In_407);
and U413 (N_413,In_6,In_89);
and U414 (N_414,In_47,In_245);
or U415 (N_415,In_249,In_257);
nand U416 (N_416,In_202,In_251);
nand U417 (N_417,In_4,In_473);
nor U418 (N_418,In_366,In_454);
and U419 (N_419,In_16,In_103);
nand U420 (N_420,In_34,In_452);
and U421 (N_421,In_396,In_61);
nand U422 (N_422,In_24,In_39);
and U423 (N_423,In_310,In_127);
nand U424 (N_424,In_451,In_370);
nand U425 (N_425,In_233,In_463);
nand U426 (N_426,In_62,In_374);
nand U427 (N_427,In_466,In_182);
nor U428 (N_428,In_328,In_340);
nor U429 (N_429,In_485,In_257);
nor U430 (N_430,In_477,In_321);
nand U431 (N_431,In_105,In_371);
and U432 (N_432,In_474,In_390);
or U433 (N_433,In_54,In_316);
nand U434 (N_434,In_28,In_114);
nor U435 (N_435,In_256,In_442);
and U436 (N_436,In_199,In_188);
nor U437 (N_437,In_497,In_180);
or U438 (N_438,In_411,In_231);
or U439 (N_439,In_178,In_74);
nand U440 (N_440,In_239,In_252);
and U441 (N_441,In_63,In_455);
nor U442 (N_442,In_396,In_268);
and U443 (N_443,In_464,In_283);
or U444 (N_444,In_228,In_326);
nand U445 (N_445,In_123,In_309);
nand U446 (N_446,In_275,In_199);
nor U447 (N_447,In_43,In_374);
and U448 (N_448,In_184,In_484);
nand U449 (N_449,In_469,In_19);
xor U450 (N_450,In_156,In_350);
and U451 (N_451,In_77,In_235);
or U452 (N_452,In_24,In_475);
nand U453 (N_453,In_459,In_474);
nor U454 (N_454,In_211,In_233);
nand U455 (N_455,In_35,In_303);
and U456 (N_456,In_421,In_301);
or U457 (N_457,In_463,In_365);
or U458 (N_458,In_228,In_163);
nand U459 (N_459,In_307,In_469);
or U460 (N_460,In_382,In_140);
or U461 (N_461,In_381,In_163);
or U462 (N_462,In_449,In_288);
or U463 (N_463,In_447,In_237);
nand U464 (N_464,In_60,In_150);
or U465 (N_465,In_331,In_453);
nand U466 (N_466,In_396,In_314);
or U467 (N_467,In_13,In_416);
nand U468 (N_468,In_50,In_310);
nand U469 (N_469,In_447,In_325);
nand U470 (N_470,In_64,In_304);
nand U471 (N_471,In_446,In_68);
and U472 (N_472,In_88,In_365);
or U473 (N_473,In_281,In_166);
and U474 (N_474,In_138,In_33);
or U475 (N_475,In_305,In_266);
nor U476 (N_476,In_56,In_287);
and U477 (N_477,In_282,In_221);
nand U478 (N_478,In_480,In_10);
and U479 (N_479,In_323,In_12);
nor U480 (N_480,In_133,In_178);
nor U481 (N_481,In_56,In_317);
nor U482 (N_482,In_202,In_255);
nor U483 (N_483,In_255,In_401);
nor U484 (N_484,In_134,In_457);
or U485 (N_485,In_196,In_4);
and U486 (N_486,In_264,In_170);
nand U487 (N_487,In_147,In_240);
nor U488 (N_488,In_142,In_482);
nor U489 (N_489,In_239,In_271);
and U490 (N_490,In_72,In_350);
and U491 (N_491,In_471,In_2);
nor U492 (N_492,In_192,In_278);
and U493 (N_493,In_113,In_44);
and U494 (N_494,In_363,In_56);
and U495 (N_495,In_323,In_176);
and U496 (N_496,In_107,In_386);
or U497 (N_497,In_318,In_12);
and U498 (N_498,In_194,In_25);
or U499 (N_499,In_144,In_338);
nor U500 (N_500,In_146,In_131);
nand U501 (N_501,In_213,In_180);
nand U502 (N_502,In_92,In_417);
or U503 (N_503,In_140,In_267);
nand U504 (N_504,In_412,In_289);
and U505 (N_505,In_356,In_269);
nor U506 (N_506,In_98,In_8);
and U507 (N_507,In_201,In_483);
or U508 (N_508,In_427,In_495);
nand U509 (N_509,In_394,In_368);
or U510 (N_510,In_298,In_479);
nand U511 (N_511,In_320,In_38);
or U512 (N_512,In_233,In_460);
xnor U513 (N_513,In_340,In_73);
and U514 (N_514,In_420,In_14);
and U515 (N_515,In_157,In_396);
and U516 (N_516,In_380,In_236);
or U517 (N_517,In_116,In_482);
and U518 (N_518,In_200,In_110);
nand U519 (N_519,In_211,In_249);
and U520 (N_520,In_478,In_25);
or U521 (N_521,In_347,In_467);
nor U522 (N_522,In_248,In_365);
or U523 (N_523,In_351,In_152);
nor U524 (N_524,In_448,In_94);
or U525 (N_525,In_59,In_434);
and U526 (N_526,In_199,In_22);
nand U527 (N_527,In_181,In_486);
nand U528 (N_528,In_172,In_264);
or U529 (N_529,In_39,In_118);
nand U530 (N_530,In_10,In_475);
and U531 (N_531,In_469,In_121);
nor U532 (N_532,In_53,In_338);
nand U533 (N_533,In_293,In_130);
and U534 (N_534,In_135,In_384);
nand U535 (N_535,In_171,In_127);
nand U536 (N_536,In_401,In_2);
nor U537 (N_537,In_257,In_312);
and U538 (N_538,In_345,In_19);
or U539 (N_539,In_140,In_230);
nor U540 (N_540,In_292,In_275);
and U541 (N_541,In_415,In_462);
nand U542 (N_542,In_136,In_481);
or U543 (N_543,In_486,In_43);
and U544 (N_544,In_476,In_491);
and U545 (N_545,In_199,In_140);
or U546 (N_546,In_259,In_432);
and U547 (N_547,In_438,In_45);
nor U548 (N_548,In_361,In_76);
and U549 (N_549,In_411,In_307);
nor U550 (N_550,In_347,In_167);
or U551 (N_551,In_342,In_473);
nand U552 (N_552,In_352,In_259);
nor U553 (N_553,In_21,In_116);
nor U554 (N_554,In_279,In_6);
or U555 (N_555,In_448,In_325);
and U556 (N_556,In_482,In_487);
nand U557 (N_557,In_60,In_455);
nand U558 (N_558,In_478,In_316);
or U559 (N_559,In_35,In_342);
or U560 (N_560,In_396,In_291);
and U561 (N_561,In_348,In_435);
or U562 (N_562,In_227,In_465);
and U563 (N_563,In_297,In_309);
or U564 (N_564,In_172,In_56);
nand U565 (N_565,In_330,In_285);
and U566 (N_566,In_116,In_87);
and U567 (N_567,In_455,In_149);
nand U568 (N_568,In_228,In_53);
and U569 (N_569,In_442,In_476);
or U570 (N_570,In_375,In_325);
nand U571 (N_571,In_297,In_201);
nor U572 (N_572,In_136,In_330);
or U573 (N_573,In_265,In_427);
nand U574 (N_574,In_348,In_317);
nand U575 (N_575,In_55,In_208);
or U576 (N_576,In_193,In_441);
xnor U577 (N_577,In_193,In_380);
nand U578 (N_578,In_200,In_235);
or U579 (N_579,In_449,In_360);
nor U580 (N_580,In_341,In_348);
xor U581 (N_581,In_150,In_190);
nor U582 (N_582,In_167,In_137);
nor U583 (N_583,In_58,In_395);
or U584 (N_584,In_314,In_203);
xnor U585 (N_585,In_256,In_353);
or U586 (N_586,In_169,In_457);
and U587 (N_587,In_434,In_113);
nand U588 (N_588,In_63,In_449);
or U589 (N_589,In_366,In_252);
nand U590 (N_590,In_484,In_365);
or U591 (N_591,In_498,In_434);
nor U592 (N_592,In_231,In_166);
nor U593 (N_593,In_460,In_489);
nor U594 (N_594,In_431,In_458);
nand U595 (N_595,In_94,In_358);
or U596 (N_596,In_255,In_285);
nor U597 (N_597,In_242,In_484);
and U598 (N_598,In_336,In_397);
and U599 (N_599,In_370,In_97);
nor U600 (N_600,In_130,In_1);
or U601 (N_601,In_79,In_400);
nor U602 (N_602,In_495,In_477);
and U603 (N_603,In_430,In_268);
nor U604 (N_604,In_375,In_208);
nor U605 (N_605,In_319,In_138);
or U606 (N_606,In_176,In_377);
nand U607 (N_607,In_451,In_305);
nor U608 (N_608,In_76,In_106);
nand U609 (N_609,In_467,In_85);
and U610 (N_610,In_402,In_476);
nand U611 (N_611,In_297,In_33);
nor U612 (N_612,In_457,In_473);
or U613 (N_613,In_11,In_89);
nand U614 (N_614,In_396,In_79);
and U615 (N_615,In_128,In_335);
nor U616 (N_616,In_492,In_329);
and U617 (N_617,In_490,In_16);
nor U618 (N_618,In_496,In_4);
and U619 (N_619,In_466,In_325);
and U620 (N_620,In_83,In_396);
nor U621 (N_621,In_443,In_469);
nor U622 (N_622,In_463,In_275);
nand U623 (N_623,In_499,In_424);
nand U624 (N_624,In_74,In_425);
nor U625 (N_625,In_386,In_376);
nor U626 (N_626,In_87,In_421);
and U627 (N_627,In_242,In_185);
and U628 (N_628,In_370,In_402);
or U629 (N_629,In_160,In_193);
nand U630 (N_630,In_62,In_246);
and U631 (N_631,In_269,In_397);
nor U632 (N_632,In_435,In_180);
and U633 (N_633,In_408,In_39);
and U634 (N_634,In_312,In_236);
and U635 (N_635,In_98,In_394);
nand U636 (N_636,In_352,In_239);
or U637 (N_637,In_356,In_79);
or U638 (N_638,In_425,In_323);
nand U639 (N_639,In_179,In_350);
or U640 (N_640,In_167,In_238);
or U641 (N_641,In_369,In_265);
and U642 (N_642,In_419,In_482);
or U643 (N_643,In_397,In_238);
and U644 (N_644,In_301,In_252);
or U645 (N_645,In_46,In_154);
or U646 (N_646,In_28,In_378);
or U647 (N_647,In_352,In_398);
and U648 (N_648,In_224,In_142);
and U649 (N_649,In_468,In_277);
or U650 (N_650,In_164,In_158);
nand U651 (N_651,In_328,In_104);
nor U652 (N_652,In_487,In_412);
nor U653 (N_653,In_240,In_23);
nand U654 (N_654,In_78,In_418);
or U655 (N_655,In_170,In_7);
and U656 (N_656,In_61,In_428);
nor U657 (N_657,In_296,In_161);
nor U658 (N_658,In_175,In_474);
or U659 (N_659,In_247,In_209);
and U660 (N_660,In_7,In_350);
or U661 (N_661,In_265,In_228);
nor U662 (N_662,In_184,In_17);
or U663 (N_663,In_474,In_186);
nor U664 (N_664,In_453,In_1);
nand U665 (N_665,In_453,In_104);
and U666 (N_666,In_480,In_375);
nor U667 (N_667,In_156,In_244);
nor U668 (N_668,In_243,In_387);
and U669 (N_669,In_178,In_247);
nand U670 (N_670,In_134,In_142);
or U671 (N_671,In_382,In_129);
or U672 (N_672,In_293,In_409);
or U673 (N_673,In_113,In_103);
and U674 (N_674,In_494,In_433);
or U675 (N_675,In_321,In_222);
or U676 (N_676,In_193,In_345);
and U677 (N_677,In_425,In_295);
nand U678 (N_678,In_115,In_437);
or U679 (N_679,In_184,In_39);
nor U680 (N_680,In_465,In_53);
nor U681 (N_681,In_228,In_354);
and U682 (N_682,In_322,In_315);
or U683 (N_683,In_308,In_97);
nor U684 (N_684,In_104,In_189);
or U685 (N_685,In_272,In_137);
xor U686 (N_686,In_92,In_465);
or U687 (N_687,In_243,In_262);
and U688 (N_688,In_396,In_51);
or U689 (N_689,In_173,In_81);
or U690 (N_690,In_219,In_445);
and U691 (N_691,In_197,In_167);
nor U692 (N_692,In_89,In_323);
and U693 (N_693,In_100,In_206);
and U694 (N_694,In_274,In_22);
or U695 (N_695,In_102,In_288);
or U696 (N_696,In_41,In_131);
or U697 (N_697,In_77,In_438);
and U698 (N_698,In_255,In_443);
or U699 (N_699,In_4,In_89);
nand U700 (N_700,In_167,In_170);
and U701 (N_701,In_323,In_118);
or U702 (N_702,In_394,In_156);
nor U703 (N_703,In_346,In_362);
or U704 (N_704,In_299,In_476);
nor U705 (N_705,In_104,In_474);
or U706 (N_706,In_78,In_392);
nor U707 (N_707,In_30,In_304);
nand U708 (N_708,In_299,In_382);
and U709 (N_709,In_251,In_35);
or U710 (N_710,In_7,In_237);
and U711 (N_711,In_241,In_361);
nand U712 (N_712,In_237,In_55);
nand U713 (N_713,In_446,In_47);
nand U714 (N_714,In_159,In_403);
nor U715 (N_715,In_314,In_457);
nand U716 (N_716,In_353,In_46);
or U717 (N_717,In_311,In_89);
nand U718 (N_718,In_119,In_495);
and U719 (N_719,In_214,In_412);
nor U720 (N_720,In_129,In_418);
nor U721 (N_721,In_483,In_121);
nor U722 (N_722,In_498,In_290);
nand U723 (N_723,In_397,In_313);
nor U724 (N_724,In_210,In_17);
nor U725 (N_725,In_258,In_455);
and U726 (N_726,In_28,In_313);
nand U727 (N_727,In_244,In_42);
nor U728 (N_728,In_420,In_382);
and U729 (N_729,In_287,In_380);
and U730 (N_730,In_209,In_213);
nand U731 (N_731,In_38,In_104);
nor U732 (N_732,In_262,In_17);
xnor U733 (N_733,In_25,In_493);
and U734 (N_734,In_243,In_28);
nand U735 (N_735,In_196,In_354);
nor U736 (N_736,In_95,In_31);
or U737 (N_737,In_406,In_278);
and U738 (N_738,In_129,In_366);
and U739 (N_739,In_36,In_166);
and U740 (N_740,In_309,In_471);
nand U741 (N_741,In_126,In_29);
nor U742 (N_742,In_27,In_121);
nand U743 (N_743,In_278,In_208);
nand U744 (N_744,In_51,In_297);
and U745 (N_745,In_201,In_425);
and U746 (N_746,In_450,In_115);
and U747 (N_747,In_306,In_416);
or U748 (N_748,In_184,In_488);
nor U749 (N_749,In_361,In_131);
nand U750 (N_750,In_136,In_486);
nand U751 (N_751,In_445,In_482);
or U752 (N_752,In_25,In_140);
and U753 (N_753,In_468,In_135);
or U754 (N_754,In_115,In_336);
nor U755 (N_755,In_339,In_287);
nand U756 (N_756,In_90,In_201);
and U757 (N_757,In_372,In_394);
and U758 (N_758,In_480,In_326);
nand U759 (N_759,In_314,In_338);
nand U760 (N_760,In_421,In_107);
nor U761 (N_761,In_423,In_77);
nand U762 (N_762,In_122,In_416);
or U763 (N_763,In_39,In_45);
and U764 (N_764,In_77,In_108);
nand U765 (N_765,In_65,In_110);
and U766 (N_766,In_329,In_204);
and U767 (N_767,In_254,In_23);
or U768 (N_768,In_175,In_482);
nor U769 (N_769,In_125,In_154);
nor U770 (N_770,In_344,In_498);
and U771 (N_771,In_48,In_357);
and U772 (N_772,In_166,In_311);
or U773 (N_773,In_120,In_246);
nand U774 (N_774,In_177,In_284);
and U775 (N_775,In_318,In_465);
nand U776 (N_776,In_224,In_124);
and U777 (N_777,In_364,In_382);
nand U778 (N_778,In_252,In_19);
nor U779 (N_779,In_16,In_398);
or U780 (N_780,In_85,In_449);
and U781 (N_781,In_182,In_289);
or U782 (N_782,In_246,In_96);
and U783 (N_783,In_276,In_138);
nor U784 (N_784,In_268,In_171);
or U785 (N_785,In_185,In_426);
or U786 (N_786,In_109,In_157);
nand U787 (N_787,In_322,In_272);
or U788 (N_788,In_188,In_113);
or U789 (N_789,In_274,In_169);
nor U790 (N_790,In_365,In_43);
nand U791 (N_791,In_94,In_206);
or U792 (N_792,In_313,In_274);
nand U793 (N_793,In_156,In_267);
nor U794 (N_794,In_147,In_475);
and U795 (N_795,In_204,In_185);
nand U796 (N_796,In_281,In_284);
and U797 (N_797,In_83,In_158);
or U798 (N_798,In_218,In_358);
nor U799 (N_799,In_286,In_212);
nand U800 (N_800,In_290,In_343);
nand U801 (N_801,In_101,In_441);
nor U802 (N_802,In_19,In_388);
and U803 (N_803,In_325,In_329);
nor U804 (N_804,In_356,In_236);
or U805 (N_805,In_146,In_453);
and U806 (N_806,In_178,In_435);
and U807 (N_807,In_186,In_183);
nor U808 (N_808,In_263,In_229);
nand U809 (N_809,In_263,In_410);
xor U810 (N_810,In_432,In_192);
nand U811 (N_811,In_4,In_11);
nand U812 (N_812,In_206,In_464);
nand U813 (N_813,In_82,In_19);
nand U814 (N_814,In_26,In_222);
nand U815 (N_815,In_250,In_161);
nor U816 (N_816,In_182,In_185);
or U817 (N_817,In_485,In_253);
nand U818 (N_818,In_423,In_264);
and U819 (N_819,In_174,In_1);
and U820 (N_820,In_248,In_50);
nand U821 (N_821,In_185,In_448);
nand U822 (N_822,In_431,In_356);
and U823 (N_823,In_392,In_190);
or U824 (N_824,In_467,In_184);
nor U825 (N_825,In_139,In_298);
and U826 (N_826,In_477,In_84);
nor U827 (N_827,In_45,In_285);
or U828 (N_828,In_134,In_382);
and U829 (N_829,In_13,In_465);
nand U830 (N_830,In_362,In_140);
and U831 (N_831,In_367,In_255);
nand U832 (N_832,In_419,In_92);
nand U833 (N_833,In_352,In_172);
or U834 (N_834,In_319,In_54);
or U835 (N_835,In_258,In_109);
or U836 (N_836,In_67,In_339);
nand U837 (N_837,In_440,In_22);
nand U838 (N_838,In_191,In_155);
or U839 (N_839,In_24,In_339);
xnor U840 (N_840,In_160,In_152);
and U841 (N_841,In_17,In_391);
and U842 (N_842,In_403,In_147);
and U843 (N_843,In_482,In_403);
nand U844 (N_844,In_71,In_416);
or U845 (N_845,In_410,In_139);
or U846 (N_846,In_48,In_260);
and U847 (N_847,In_430,In_283);
and U848 (N_848,In_117,In_172);
nor U849 (N_849,In_39,In_86);
nand U850 (N_850,In_80,In_473);
nand U851 (N_851,In_59,In_405);
nand U852 (N_852,In_306,In_221);
and U853 (N_853,In_97,In_128);
nand U854 (N_854,In_245,In_475);
nor U855 (N_855,In_152,In_68);
and U856 (N_856,In_3,In_435);
or U857 (N_857,In_235,In_44);
or U858 (N_858,In_290,In_406);
nor U859 (N_859,In_342,In_307);
or U860 (N_860,In_181,In_498);
or U861 (N_861,In_57,In_96);
nand U862 (N_862,In_75,In_468);
nand U863 (N_863,In_228,In_340);
nor U864 (N_864,In_244,In_211);
xnor U865 (N_865,In_202,In_147);
or U866 (N_866,In_301,In_19);
and U867 (N_867,In_483,In_51);
and U868 (N_868,In_21,In_18);
and U869 (N_869,In_124,In_474);
or U870 (N_870,In_462,In_337);
nor U871 (N_871,In_83,In_410);
or U872 (N_872,In_98,In_177);
nor U873 (N_873,In_444,In_362);
nand U874 (N_874,In_482,In_212);
nand U875 (N_875,In_202,In_358);
nor U876 (N_876,In_153,In_460);
or U877 (N_877,In_233,In_350);
and U878 (N_878,In_380,In_35);
nand U879 (N_879,In_55,In_274);
nor U880 (N_880,In_493,In_59);
or U881 (N_881,In_333,In_161);
nand U882 (N_882,In_326,In_55);
nor U883 (N_883,In_306,In_238);
or U884 (N_884,In_125,In_466);
and U885 (N_885,In_467,In_6);
or U886 (N_886,In_269,In_494);
and U887 (N_887,In_54,In_191);
and U888 (N_888,In_67,In_468);
nor U889 (N_889,In_385,In_51);
and U890 (N_890,In_224,In_318);
nor U891 (N_891,In_208,In_301);
nand U892 (N_892,In_325,In_345);
nor U893 (N_893,In_484,In_431);
xor U894 (N_894,In_34,In_228);
xor U895 (N_895,In_201,In_411);
xnor U896 (N_896,In_462,In_82);
and U897 (N_897,In_152,In_378);
nor U898 (N_898,In_326,In_251);
and U899 (N_899,In_459,In_30);
or U900 (N_900,In_41,In_248);
nor U901 (N_901,In_193,In_150);
nor U902 (N_902,In_15,In_266);
or U903 (N_903,In_325,In_257);
or U904 (N_904,In_279,In_237);
nor U905 (N_905,In_89,In_197);
and U906 (N_906,In_75,In_332);
nor U907 (N_907,In_312,In_487);
and U908 (N_908,In_122,In_231);
or U909 (N_909,In_189,In_274);
nor U910 (N_910,In_439,In_318);
or U911 (N_911,In_462,In_133);
nor U912 (N_912,In_115,In_1);
nor U913 (N_913,In_116,In_211);
nor U914 (N_914,In_335,In_23);
or U915 (N_915,In_346,In_153);
or U916 (N_916,In_409,In_371);
or U917 (N_917,In_51,In_335);
nor U918 (N_918,In_264,In_141);
or U919 (N_919,In_453,In_12);
nand U920 (N_920,In_56,In_84);
and U921 (N_921,In_192,In_21);
nor U922 (N_922,In_273,In_479);
nor U923 (N_923,In_292,In_185);
or U924 (N_924,In_127,In_371);
nor U925 (N_925,In_499,In_287);
and U926 (N_926,In_231,In_226);
and U927 (N_927,In_438,In_57);
and U928 (N_928,In_437,In_469);
nor U929 (N_929,In_142,In_298);
nor U930 (N_930,In_48,In_211);
and U931 (N_931,In_156,In_153);
or U932 (N_932,In_1,In_333);
nor U933 (N_933,In_476,In_401);
and U934 (N_934,In_319,In_244);
nor U935 (N_935,In_196,In_75);
or U936 (N_936,In_480,In_1);
nand U937 (N_937,In_350,In_430);
nand U938 (N_938,In_403,In_420);
nand U939 (N_939,In_285,In_252);
and U940 (N_940,In_383,In_131);
or U941 (N_941,In_203,In_338);
nand U942 (N_942,In_148,In_113);
nand U943 (N_943,In_245,In_254);
nand U944 (N_944,In_112,In_111);
nor U945 (N_945,In_280,In_253);
or U946 (N_946,In_53,In_115);
nor U947 (N_947,In_38,In_412);
or U948 (N_948,In_320,In_47);
nand U949 (N_949,In_358,In_45);
nor U950 (N_950,In_12,In_108);
or U951 (N_951,In_297,In_368);
and U952 (N_952,In_368,In_354);
nor U953 (N_953,In_20,In_476);
and U954 (N_954,In_115,In_226);
nand U955 (N_955,In_329,In_450);
or U956 (N_956,In_329,In_244);
nand U957 (N_957,In_481,In_291);
nand U958 (N_958,In_77,In_205);
and U959 (N_959,In_469,In_375);
and U960 (N_960,In_186,In_187);
and U961 (N_961,In_393,In_215);
or U962 (N_962,In_98,In_48);
nand U963 (N_963,In_234,In_81);
or U964 (N_964,In_19,In_482);
and U965 (N_965,In_107,In_294);
or U966 (N_966,In_325,In_424);
nor U967 (N_967,In_191,In_178);
nand U968 (N_968,In_165,In_45);
nand U969 (N_969,In_309,In_140);
nor U970 (N_970,In_489,In_171);
nand U971 (N_971,In_56,In_193);
and U972 (N_972,In_144,In_72);
nor U973 (N_973,In_116,In_444);
and U974 (N_974,In_269,In_216);
nor U975 (N_975,In_73,In_96);
nand U976 (N_976,In_361,In_161);
or U977 (N_977,In_29,In_265);
nor U978 (N_978,In_92,In_119);
nand U979 (N_979,In_285,In_196);
nand U980 (N_980,In_470,In_73);
nor U981 (N_981,In_68,In_434);
and U982 (N_982,In_406,In_252);
or U983 (N_983,In_329,In_19);
nand U984 (N_984,In_374,In_185);
nor U985 (N_985,In_107,In_159);
and U986 (N_986,In_461,In_265);
and U987 (N_987,In_312,In_185);
nor U988 (N_988,In_497,In_219);
nand U989 (N_989,In_347,In_166);
and U990 (N_990,In_59,In_129);
and U991 (N_991,In_161,In_314);
nand U992 (N_992,In_118,In_20);
and U993 (N_993,In_180,In_470);
or U994 (N_994,In_312,In_293);
or U995 (N_995,In_425,In_81);
nor U996 (N_996,In_138,In_407);
nor U997 (N_997,In_408,In_138);
or U998 (N_998,In_476,In_378);
nor U999 (N_999,In_279,In_11);
nor U1000 (N_1000,N_957,N_666);
and U1001 (N_1001,N_974,N_873);
or U1002 (N_1002,N_388,N_252);
nand U1003 (N_1003,N_211,N_828);
nand U1004 (N_1004,N_85,N_169);
nor U1005 (N_1005,N_155,N_164);
nor U1006 (N_1006,N_330,N_447);
and U1007 (N_1007,N_538,N_460);
and U1008 (N_1008,N_893,N_212);
nand U1009 (N_1009,N_25,N_781);
or U1010 (N_1010,N_333,N_355);
nand U1011 (N_1011,N_379,N_561);
and U1012 (N_1012,N_316,N_632);
and U1013 (N_1013,N_188,N_879);
or U1014 (N_1014,N_329,N_56);
nor U1015 (N_1015,N_687,N_838);
nand U1016 (N_1016,N_131,N_527);
or U1017 (N_1017,N_789,N_314);
and U1018 (N_1018,N_681,N_998);
nor U1019 (N_1019,N_778,N_405);
or U1020 (N_1020,N_842,N_593);
or U1021 (N_1021,N_445,N_891);
nor U1022 (N_1022,N_745,N_702);
or U1023 (N_1023,N_441,N_449);
or U1024 (N_1024,N_907,N_346);
nand U1025 (N_1025,N_911,N_830);
and U1026 (N_1026,N_765,N_611);
nand U1027 (N_1027,N_485,N_18);
or U1028 (N_1028,N_654,N_216);
or U1029 (N_1029,N_499,N_776);
or U1030 (N_1030,N_874,N_864);
nand U1031 (N_1031,N_549,N_756);
nor U1032 (N_1032,N_746,N_440);
nor U1033 (N_1033,N_3,N_937);
or U1034 (N_1034,N_847,N_601);
or U1035 (N_1035,N_53,N_835);
nand U1036 (N_1036,N_165,N_84);
or U1037 (N_1037,N_125,N_850);
nand U1038 (N_1038,N_564,N_978);
and U1039 (N_1039,N_392,N_908);
nor U1040 (N_1040,N_111,N_612);
or U1041 (N_1041,N_452,N_836);
and U1042 (N_1042,N_130,N_77);
nor U1043 (N_1043,N_571,N_709);
nand U1044 (N_1044,N_168,N_105);
nor U1045 (N_1045,N_656,N_455);
or U1046 (N_1046,N_71,N_610);
nand U1047 (N_1047,N_132,N_143);
or U1048 (N_1048,N_385,N_432);
nor U1049 (N_1049,N_990,N_283);
nand U1050 (N_1050,N_587,N_117);
nor U1051 (N_1051,N_672,N_40);
or U1052 (N_1052,N_288,N_938);
or U1053 (N_1053,N_903,N_173);
nor U1054 (N_1054,N_241,N_416);
nand U1055 (N_1055,N_180,N_403);
or U1056 (N_1056,N_896,N_674);
or U1057 (N_1057,N_556,N_365);
or U1058 (N_1058,N_997,N_194);
and U1059 (N_1059,N_213,N_785);
or U1060 (N_1060,N_635,N_665);
nor U1061 (N_1061,N_918,N_516);
nand U1062 (N_1062,N_332,N_679);
nor U1063 (N_1063,N_179,N_472);
nor U1064 (N_1064,N_711,N_774);
nand U1065 (N_1065,N_890,N_536);
nor U1066 (N_1066,N_588,N_70);
and U1067 (N_1067,N_250,N_518);
and U1068 (N_1068,N_382,N_510);
nor U1069 (N_1069,N_706,N_210);
or U1070 (N_1070,N_359,N_474);
nor U1071 (N_1071,N_16,N_232);
or U1072 (N_1072,N_264,N_772);
nor U1073 (N_1073,N_470,N_892);
and U1074 (N_1074,N_708,N_968);
nand U1075 (N_1075,N_15,N_428);
or U1076 (N_1076,N_186,N_0);
nand U1077 (N_1077,N_504,N_620);
and U1078 (N_1078,N_336,N_613);
nand U1079 (N_1079,N_668,N_435);
nor U1080 (N_1080,N_47,N_55);
nand U1081 (N_1081,N_716,N_791);
and U1082 (N_1082,N_985,N_374);
nand U1083 (N_1083,N_973,N_685);
nand U1084 (N_1084,N_949,N_418);
nand U1085 (N_1085,N_138,N_952);
nand U1086 (N_1086,N_172,N_68);
nand U1087 (N_1087,N_79,N_39);
or U1088 (N_1088,N_479,N_285);
nor U1089 (N_1089,N_511,N_573);
and U1090 (N_1090,N_565,N_191);
nand U1091 (N_1091,N_703,N_292);
nand U1092 (N_1092,N_944,N_487);
nor U1093 (N_1093,N_348,N_742);
or U1094 (N_1094,N_266,N_956);
and U1095 (N_1095,N_78,N_491);
and U1096 (N_1096,N_370,N_151);
nor U1097 (N_1097,N_701,N_969);
nor U1098 (N_1098,N_103,N_768);
nor U1099 (N_1099,N_489,N_614);
or U1100 (N_1100,N_800,N_921);
nor U1101 (N_1101,N_296,N_256);
nor U1102 (N_1102,N_664,N_135);
or U1103 (N_1103,N_503,N_790);
nand U1104 (N_1104,N_263,N_784);
and U1105 (N_1105,N_675,N_943);
nand U1106 (N_1106,N_696,N_655);
nor U1107 (N_1107,N_667,N_96);
nand U1108 (N_1108,N_539,N_744);
nand U1109 (N_1109,N_76,N_760);
or U1110 (N_1110,N_699,N_228);
nand U1111 (N_1111,N_397,N_112);
nand U1112 (N_1112,N_698,N_290);
and U1113 (N_1113,N_933,N_605);
nand U1114 (N_1114,N_609,N_748);
nor U1115 (N_1115,N_486,N_235);
nor U1116 (N_1116,N_197,N_532);
or U1117 (N_1117,N_851,N_924);
or U1118 (N_1118,N_129,N_458);
nand U1119 (N_1119,N_773,N_726);
nand U1120 (N_1120,N_728,N_108);
and U1121 (N_1121,N_976,N_753);
nor U1122 (N_1122,N_647,N_488);
nor U1123 (N_1123,N_963,N_967);
nor U1124 (N_1124,N_592,N_683);
or U1125 (N_1125,N_451,N_826);
or U1126 (N_1126,N_399,N_528);
nand U1127 (N_1127,N_951,N_350);
or U1128 (N_1128,N_187,N_810);
nand U1129 (N_1129,N_886,N_860);
nand U1130 (N_1130,N_803,N_960);
and U1131 (N_1131,N_580,N_747);
and U1132 (N_1132,N_730,N_214);
or U1133 (N_1133,N_302,N_567);
nor U1134 (N_1134,N_648,N_575);
nand U1135 (N_1135,N_551,N_900);
and U1136 (N_1136,N_846,N_183);
or U1137 (N_1137,N_877,N_775);
and U1138 (N_1138,N_340,N_88);
and U1139 (N_1139,N_940,N_141);
nand U1140 (N_1140,N_331,N_731);
nor U1141 (N_1141,N_64,N_21);
or U1142 (N_1142,N_466,N_268);
or U1143 (N_1143,N_688,N_325);
nor U1144 (N_1144,N_59,N_931);
nand U1145 (N_1145,N_626,N_693);
and U1146 (N_1146,N_616,N_855);
and U1147 (N_1147,N_414,N_691);
nor U1148 (N_1148,N_75,N_157);
nor U1149 (N_1149,N_83,N_30);
nand U1150 (N_1150,N_942,N_427);
or U1151 (N_1151,N_324,N_396);
or U1152 (N_1152,N_408,N_307);
and U1153 (N_1153,N_36,N_249);
nor U1154 (N_1154,N_782,N_865);
nor U1155 (N_1155,N_401,N_184);
and U1156 (N_1156,N_856,N_65);
nor U1157 (N_1157,N_872,N_448);
nor U1158 (N_1158,N_522,N_913);
xor U1159 (N_1159,N_542,N_787);
or U1160 (N_1160,N_357,N_992);
and U1161 (N_1161,N_994,N_34);
or U1162 (N_1162,N_66,N_583);
and U1163 (N_1163,N_69,N_404);
and U1164 (N_1164,N_136,N_193);
and U1165 (N_1165,N_335,N_255);
nor U1166 (N_1166,N_398,N_321);
and U1167 (N_1167,N_337,N_537);
nand U1168 (N_1168,N_148,N_553);
nor U1169 (N_1169,N_869,N_298);
nand U1170 (N_1170,N_391,N_928);
nand U1171 (N_1171,N_300,N_282);
nand U1172 (N_1172,N_160,N_27);
or U1173 (N_1173,N_431,N_502);
nor U1174 (N_1174,N_97,N_955);
nand U1175 (N_1175,N_102,N_645);
and U1176 (N_1176,N_607,N_277);
or U1177 (N_1177,N_552,N_154);
xnor U1178 (N_1178,N_811,N_548);
or U1179 (N_1179,N_736,N_63);
or U1180 (N_1180,N_818,N_189);
nor U1181 (N_1181,N_729,N_858);
or U1182 (N_1182,N_771,N_630);
nand U1183 (N_1183,N_145,N_101);
or U1184 (N_1184,N_281,N_638);
or U1185 (N_1185,N_659,N_11);
or U1186 (N_1186,N_286,N_737);
nand U1187 (N_1187,N_496,N_498);
nand U1188 (N_1188,N_217,N_48);
nor U1189 (N_1189,N_305,N_159);
or U1190 (N_1190,N_10,N_12);
or U1191 (N_1191,N_854,N_462);
nor U1192 (N_1192,N_415,N_207);
and U1193 (N_1193,N_393,N_425);
nand U1194 (N_1194,N_410,N_766);
and U1195 (N_1195,N_58,N_291);
and U1196 (N_1196,N_520,N_663);
and U1197 (N_1197,N_843,N_424);
xor U1198 (N_1198,N_371,N_725);
nor U1199 (N_1199,N_293,N_259);
or U1200 (N_1200,N_807,N_899);
or U1201 (N_1201,N_671,N_310);
nor U1202 (N_1202,N_246,N_334);
nand U1203 (N_1203,N_377,N_999);
or U1204 (N_1204,N_895,N_430);
nor U1205 (N_1205,N_351,N_954);
and U1206 (N_1206,N_114,N_739);
nor U1207 (N_1207,N_868,N_303);
or U1208 (N_1208,N_146,N_912);
or U1209 (N_1209,N_144,N_347);
nor U1210 (N_1210,N_684,N_167);
or U1211 (N_1211,N_544,N_915);
nand U1212 (N_1212,N_966,N_578);
xnor U1213 (N_1213,N_586,N_859);
or U1214 (N_1214,N_342,N_9);
and U1215 (N_1215,N_982,N_318);
nor U1216 (N_1216,N_832,N_761);
and U1217 (N_1217,N_450,N_390);
or U1218 (N_1218,N_625,N_320);
and U1219 (N_1219,N_732,N_794);
nor U1220 (N_1220,N_808,N_429);
nand U1221 (N_1221,N_653,N_934);
nand U1222 (N_1222,N_526,N_220);
nor U1223 (N_1223,N_829,N_524);
nor U1224 (N_1224,N_273,N_417);
or U1225 (N_1225,N_769,N_411);
and U1226 (N_1226,N_670,N_546);
nand U1227 (N_1227,N_602,N_555);
nand U1228 (N_1228,N_735,N_633);
and U1229 (N_1229,N_916,N_792);
nand U1230 (N_1230,N_274,N_161);
or U1231 (N_1231,N_473,N_94);
nor U1232 (N_1232,N_834,N_33);
or U1233 (N_1233,N_227,N_92);
nand U1234 (N_1234,N_170,N_322);
nand U1235 (N_1235,N_755,N_381);
and U1236 (N_1236,N_42,N_917);
and U1237 (N_1237,N_1,N_584);
or U1238 (N_1238,N_880,N_793);
nand U1239 (N_1239,N_799,N_280);
and U1240 (N_1240,N_433,N_641);
nor U1241 (N_1241,N_465,N_513);
and U1242 (N_1242,N_500,N_150);
nand U1243 (N_1243,N_929,N_311);
nand U1244 (N_1244,N_245,N_953);
nor U1245 (N_1245,N_505,N_327);
or U1246 (N_1246,N_878,N_461);
or U1247 (N_1247,N_741,N_295);
nor U1248 (N_1248,N_313,N_243);
nand U1249 (N_1249,N_927,N_981);
or U1250 (N_1250,N_242,N_517);
and U1251 (N_1251,N_849,N_743);
and U1252 (N_1252,N_560,N_82);
nand U1253 (N_1253,N_669,N_876);
or U1254 (N_1254,N_362,N_545);
and U1255 (N_1255,N_80,N_475);
nand U1256 (N_1256,N_889,N_205);
or U1257 (N_1257,N_99,N_363);
nor U1258 (N_1258,N_468,N_986);
or U1259 (N_1259,N_471,N_176);
nand U1260 (N_1260,N_270,N_871);
and U1261 (N_1261,N_219,N_284);
or U1262 (N_1262,N_901,N_673);
nand U1263 (N_1263,N_221,N_533);
or U1264 (N_1264,N_478,N_617);
and U1265 (N_1265,N_23,N_525);
or U1266 (N_1266,N_20,N_910);
nor U1267 (N_1267,N_883,N_113);
nor U1268 (N_1268,N_24,N_361);
nand U1269 (N_1269,N_650,N_175);
and U1270 (N_1270,N_31,N_225);
nor U1271 (N_1271,N_271,N_805);
nor U1272 (N_1272,N_759,N_875);
nor U1273 (N_1273,N_939,N_240);
nor U1274 (N_1274,N_109,N_950);
nor U1275 (N_1275,N_62,N_770);
xor U1276 (N_1276,N_804,N_695);
or U1277 (N_1277,N_712,N_570);
nor U1278 (N_1278,N_733,N_162);
nor U1279 (N_1279,N_577,N_163);
or U1280 (N_1280,N_238,N_233);
nand U1281 (N_1281,N_477,N_493);
nor U1282 (N_1282,N_824,N_356);
nand U1283 (N_1283,N_642,N_833);
and U1284 (N_1284,N_234,N_482);
nor U1285 (N_1285,N_369,N_959);
nor U1286 (N_1286,N_122,N_541);
nor U1287 (N_1287,N_386,N_209);
nor U1288 (N_1288,N_267,N_754);
or U1289 (N_1289,N_190,N_993);
nand U1290 (N_1290,N_905,N_715);
nand U1291 (N_1291,N_975,N_140);
or U1292 (N_1292,N_783,N_367);
nand U1293 (N_1293,N_618,N_652);
nor U1294 (N_1294,N_662,N_74);
or U1295 (N_1295,N_598,N_501);
and U1296 (N_1296,N_139,N_831);
nand U1297 (N_1297,N_198,N_50);
and U1298 (N_1298,N_962,N_349);
nand U1299 (N_1299,N_757,N_530);
nand U1300 (N_1300,N_239,N_989);
nor U1301 (N_1301,N_278,N_629);
or U1302 (N_1302,N_121,N_697);
and U1303 (N_1303,N_802,N_258);
or U1304 (N_1304,N_559,N_983);
nor U1305 (N_1305,N_558,N_623);
nor U1306 (N_1306,N_970,N_294);
nand U1307 (N_1307,N_853,N_437);
and U1308 (N_1308,N_694,N_977);
nand U1309 (N_1309,N_705,N_945);
or U1310 (N_1310,N_758,N_195);
nand U1311 (N_1311,N_467,N_67);
and U1312 (N_1312,N_158,N_738);
nor U1313 (N_1313,N_229,N_506);
and U1314 (N_1314,N_287,N_199);
or U1315 (N_1315,N_224,N_202);
and U1316 (N_1316,N_231,N_627);
nand U1317 (N_1317,N_120,N_579);
and U1318 (N_1318,N_987,N_395);
nand U1319 (N_1319,N_54,N_384);
nand U1320 (N_1320,N_196,N_866);
nor U1321 (N_1321,N_837,N_319);
and U1322 (N_1322,N_740,N_204);
nand U1323 (N_1323,N_707,N_814);
xnor U1324 (N_1324,N_534,N_628);
nand U1325 (N_1325,N_649,N_749);
or U1326 (N_1326,N_515,N_402);
nand U1327 (N_1327,N_123,N_723);
and U1328 (N_1328,N_572,N_606);
nand U1329 (N_1329,N_87,N_603);
nand U1330 (N_1330,N_244,N_301);
nand U1331 (N_1331,N_444,N_91);
and U1332 (N_1332,N_798,N_454);
nor U1333 (N_1333,N_710,N_44);
and U1334 (N_1334,N_387,N_643);
and U1335 (N_1335,N_812,N_594);
nand U1336 (N_1336,N_115,N_909);
nand U1337 (N_1337,N_275,N_845);
and U1338 (N_1338,N_888,N_7);
nor U1339 (N_1339,N_817,N_407);
or U1340 (N_1340,N_152,N_262);
or U1341 (N_1341,N_870,N_988);
or U1342 (N_1342,N_700,N_480);
nand U1343 (N_1343,N_971,N_727);
or U1344 (N_1344,N_306,N_752);
nor U1345 (N_1345,N_299,N_339);
nand U1346 (N_1346,N_438,N_353);
or U1347 (N_1347,N_93,N_439);
and U1348 (N_1348,N_61,N_932);
and U1349 (N_1349,N_677,N_636);
and U1350 (N_1350,N_14,N_106);
nand U1351 (N_1351,N_98,N_236);
or U1352 (N_1352,N_453,N_965);
nor U1353 (N_1353,N_208,N_394);
nand U1354 (N_1354,N_621,N_964);
nor U1355 (N_1355,N_45,N_328);
nor U1356 (N_1356,N_780,N_116);
and U1357 (N_1357,N_156,N_599);
or U1358 (N_1358,N_389,N_750);
nand U1359 (N_1359,N_995,N_574);
nor U1360 (N_1360,N_763,N_421);
nand U1361 (N_1361,N_72,N_481);
or U1362 (N_1362,N_137,N_519);
nand U1363 (N_1363,N_713,N_341);
nor U1364 (N_1364,N_585,N_867);
nor U1365 (N_1365,N_717,N_247);
and U1366 (N_1366,N_107,N_128);
nor U1367 (N_1367,N_682,N_272);
or U1368 (N_1368,N_142,N_852);
or U1369 (N_1369,N_581,N_366);
nor U1370 (N_1370,N_185,N_495);
nor U1371 (N_1371,N_308,N_930);
nor U1372 (N_1372,N_413,N_380);
and U1373 (N_1373,N_261,N_133);
or U1374 (N_1374,N_651,N_215);
or U1375 (N_1375,N_41,N_885);
nor U1376 (N_1376,N_35,N_821);
nor U1377 (N_1377,N_436,N_680);
nand U1378 (N_1378,N_984,N_338);
and U1379 (N_1379,N_237,N_373);
and U1380 (N_1380,N_557,N_86);
and U1381 (N_1381,N_762,N_312);
or U1382 (N_1382,N_947,N_223);
or U1383 (N_1383,N_920,N_149);
nor U1384 (N_1384,N_619,N_344);
nand U1385 (N_1385,N_218,N_529);
or U1386 (N_1386,N_343,N_568);
nand U1387 (N_1387,N_19,N_73);
nor U1388 (N_1388,N_690,N_823);
nand U1389 (N_1389,N_596,N_358);
nand U1390 (N_1390,N_660,N_315);
or U1391 (N_1391,N_898,N_29);
nand U1392 (N_1392,N_276,N_22);
nand U1393 (N_1393,N_914,N_839);
nor U1394 (N_1394,N_523,N_841);
or U1395 (N_1395,N_269,N_622);
nand U1396 (N_1396,N_719,N_861);
xor U1397 (N_1397,N_206,N_352);
or U1398 (N_1398,N_95,N_492);
nor U1399 (N_1399,N_597,N_819);
nor U1400 (N_1400,N_323,N_126);
nand U1401 (N_1401,N_509,N_925);
or U1402 (N_1402,N_81,N_354);
nor U1403 (N_1403,N_192,N_809);
and U1404 (N_1404,N_661,N_721);
and U1405 (N_1405,N_372,N_426);
nor U1406 (N_1406,N_566,N_521);
nand U1407 (N_1407,N_406,N_483);
nor U1408 (N_1408,N_595,N_200);
nand U1409 (N_1409,N_4,N_806);
nand U1410 (N_1410,N_419,N_822);
and U1411 (N_1411,N_718,N_547);
nand U1412 (N_1412,N_562,N_902);
nand U1413 (N_1413,N_17,N_251);
nor U1414 (N_1414,N_904,N_825);
nor U1415 (N_1415,N_923,N_815);
nor U1416 (N_1416,N_177,N_494);
or U1417 (N_1417,N_38,N_52);
nand U1418 (N_1418,N_919,N_827);
nand U1419 (N_1419,N_412,N_801);
nor U1420 (N_1420,N_375,N_46);
and U1421 (N_1421,N_991,N_464);
nor U1422 (N_1422,N_936,N_118);
and U1423 (N_1423,N_786,N_124);
nand U1424 (N_1424,N_174,N_639);
or U1425 (N_1425,N_476,N_222);
nand U1426 (N_1426,N_253,N_980);
or U1427 (N_1427,N_897,N_345);
and U1428 (N_1428,N_882,N_576);
and U1429 (N_1429,N_51,N_604);
or U1430 (N_1430,N_631,N_884);
nand U1431 (N_1431,N_941,N_686);
nand U1432 (N_1432,N_857,N_796);
nand U1433 (N_1433,N_304,N_569);
and U1434 (N_1434,N_996,N_862);
or U1435 (N_1435,N_90,N_724);
nand U1436 (N_1436,N_497,N_531);
and U1437 (N_1437,N_226,N_820);
nand U1438 (N_1438,N_767,N_935);
or U1439 (N_1439,N_420,N_615);
or U1440 (N_1440,N_779,N_844);
or U1441 (N_1441,N_948,N_8);
nand U1442 (N_1442,N_507,N_201);
nand U1443 (N_1443,N_309,N_230);
nand U1444 (N_1444,N_676,N_104);
nor U1445 (N_1445,N_134,N_317);
nand U1446 (N_1446,N_127,N_60);
nor U1447 (N_1447,N_171,N_657);
nor U1448 (N_1448,N_469,N_751);
nor U1449 (N_1449,N_364,N_508);
nand U1450 (N_1450,N_297,N_265);
nor U1451 (N_1451,N_147,N_926);
or U1452 (N_1452,N_906,N_490);
nor U1453 (N_1453,N_590,N_863);
and U1454 (N_1454,N_840,N_714);
nor U1455 (N_1455,N_254,N_5);
and U1456 (N_1456,N_816,N_457);
nand U1457 (N_1457,N_89,N_514);
nor U1458 (N_1458,N_894,N_777);
or U1459 (N_1459,N_32,N_582);
and U1460 (N_1460,N_26,N_376);
nor U1461 (N_1461,N_543,N_442);
and U1462 (N_1462,N_153,N_646);
and U1463 (N_1463,N_634,N_788);
nor U1464 (N_1464,N_689,N_704);
nand U1465 (N_1465,N_257,N_540);
nor U1466 (N_1466,N_881,N_166);
and U1467 (N_1467,N_400,N_378);
nor U1468 (N_1468,N_734,N_456);
nand U1469 (N_1469,N_459,N_887);
nand U1470 (N_1470,N_637,N_624);
or U1471 (N_1471,N_446,N_550);
or U1472 (N_1472,N_13,N_972);
nor U1473 (N_1473,N_368,N_119);
nand U1474 (N_1474,N_260,N_182);
or U1475 (N_1475,N_443,N_946);
nor U1476 (N_1476,N_644,N_563);
and U1477 (N_1477,N_248,N_591);
or U1478 (N_1478,N_203,N_423);
or U1479 (N_1479,N_178,N_764);
nand U1480 (N_1480,N_848,N_28);
nor U1481 (N_1481,N_795,N_722);
and U1482 (N_1482,N_658,N_110);
nand U1483 (N_1483,N_49,N_409);
or U1484 (N_1484,N_43,N_434);
and U1485 (N_1485,N_360,N_589);
or U1486 (N_1486,N_463,N_6);
and U1487 (N_1487,N_922,N_600);
nor U1488 (N_1488,N_554,N_797);
or U1489 (N_1489,N_484,N_181);
and U1490 (N_1490,N_326,N_608);
and U1491 (N_1491,N_2,N_678);
or U1492 (N_1492,N_57,N_279);
nor U1493 (N_1493,N_100,N_512);
nand U1494 (N_1494,N_958,N_289);
or U1495 (N_1495,N_37,N_692);
nor U1496 (N_1496,N_813,N_979);
nand U1497 (N_1497,N_383,N_422);
nor U1498 (N_1498,N_640,N_720);
and U1499 (N_1499,N_535,N_961);
and U1500 (N_1500,N_723,N_365);
and U1501 (N_1501,N_833,N_390);
and U1502 (N_1502,N_362,N_507);
and U1503 (N_1503,N_602,N_447);
nor U1504 (N_1504,N_437,N_686);
nand U1505 (N_1505,N_753,N_515);
nor U1506 (N_1506,N_97,N_406);
nor U1507 (N_1507,N_895,N_32);
nand U1508 (N_1508,N_832,N_666);
nor U1509 (N_1509,N_489,N_79);
nor U1510 (N_1510,N_593,N_188);
nand U1511 (N_1511,N_682,N_223);
or U1512 (N_1512,N_730,N_833);
and U1513 (N_1513,N_764,N_558);
or U1514 (N_1514,N_448,N_915);
nand U1515 (N_1515,N_0,N_695);
nand U1516 (N_1516,N_91,N_716);
and U1517 (N_1517,N_963,N_95);
or U1518 (N_1518,N_709,N_901);
nor U1519 (N_1519,N_125,N_63);
nor U1520 (N_1520,N_815,N_754);
or U1521 (N_1521,N_491,N_511);
nor U1522 (N_1522,N_50,N_797);
and U1523 (N_1523,N_445,N_440);
xnor U1524 (N_1524,N_658,N_916);
nor U1525 (N_1525,N_924,N_613);
xor U1526 (N_1526,N_809,N_478);
and U1527 (N_1527,N_665,N_866);
nor U1528 (N_1528,N_352,N_790);
and U1529 (N_1529,N_53,N_70);
or U1530 (N_1530,N_886,N_413);
or U1531 (N_1531,N_882,N_392);
nor U1532 (N_1532,N_582,N_942);
and U1533 (N_1533,N_461,N_465);
and U1534 (N_1534,N_416,N_838);
or U1535 (N_1535,N_808,N_211);
and U1536 (N_1536,N_334,N_943);
nand U1537 (N_1537,N_55,N_760);
or U1538 (N_1538,N_360,N_9);
nand U1539 (N_1539,N_127,N_366);
and U1540 (N_1540,N_377,N_795);
or U1541 (N_1541,N_405,N_662);
or U1542 (N_1542,N_553,N_510);
nand U1543 (N_1543,N_769,N_917);
or U1544 (N_1544,N_128,N_272);
or U1545 (N_1545,N_423,N_411);
or U1546 (N_1546,N_480,N_360);
or U1547 (N_1547,N_908,N_581);
nor U1548 (N_1548,N_65,N_215);
or U1549 (N_1549,N_39,N_395);
nand U1550 (N_1550,N_101,N_226);
nor U1551 (N_1551,N_567,N_420);
nor U1552 (N_1552,N_147,N_924);
nand U1553 (N_1553,N_848,N_781);
and U1554 (N_1554,N_612,N_980);
or U1555 (N_1555,N_45,N_809);
or U1556 (N_1556,N_489,N_633);
nand U1557 (N_1557,N_912,N_765);
nand U1558 (N_1558,N_713,N_444);
nand U1559 (N_1559,N_537,N_18);
nor U1560 (N_1560,N_310,N_144);
nor U1561 (N_1561,N_714,N_50);
nand U1562 (N_1562,N_153,N_119);
or U1563 (N_1563,N_187,N_486);
and U1564 (N_1564,N_976,N_290);
and U1565 (N_1565,N_934,N_838);
and U1566 (N_1566,N_894,N_83);
and U1567 (N_1567,N_581,N_122);
and U1568 (N_1568,N_209,N_54);
nor U1569 (N_1569,N_448,N_997);
and U1570 (N_1570,N_811,N_539);
and U1571 (N_1571,N_562,N_875);
nor U1572 (N_1572,N_59,N_829);
and U1573 (N_1573,N_260,N_929);
or U1574 (N_1574,N_141,N_699);
nand U1575 (N_1575,N_22,N_590);
nand U1576 (N_1576,N_548,N_770);
and U1577 (N_1577,N_534,N_95);
nor U1578 (N_1578,N_580,N_916);
xor U1579 (N_1579,N_966,N_44);
or U1580 (N_1580,N_652,N_998);
nor U1581 (N_1581,N_552,N_66);
and U1582 (N_1582,N_386,N_862);
nand U1583 (N_1583,N_321,N_652);
nor U1584 (N_1584,N_938,N_807);
nor U1585 (N_1585,N_588,N_895);
and U1586 (N_1586,N_506,N_391);
nand U1587 (N_1587,N_435,N_53);
nor U1588 (N_1588,N_195,N_985);
nand U1589 (N_1589,N_527,N_258);
nor U1590 (N_1590,N_115,N_234);
nor U1591 (N_1591,N_498,N_61);
or U1592 (N_1592,N_472,N_572);
or U1593 (N_1593,N_657,N_214);
nor U1594 (N_1594,N_602,N_200);
or U1595 (N_1595,N_694,N_128);
or U1596 (N_1596,N_621,N_31);
and U1597 (N_1597,N_708,N_772);
nand U1598 (N_1598,N_893,N_430);
nor U1599 (N_1599,N_613,N_973);
nor U1600 (N_1600,N_619,N_295);
and U1601 (N_1601,N_78,N_462);
or U1602 (N_1602,N_794,N_736);
nand U1603 (N_1603,N_604,N_788);
nand U1604 (N_1604,N_700,N_146);
or U1605 (N_1605,N_329,N_323);
or U1606 (N_1606,N_559,N_982);
nor U1607 (N_1607,N_199,N_252);
nand U1608 (N_1608,N_155,N_494);
and U1609 (N_1609,N_621,N_982);
or U1610 (N_1610,N_378,N_494);
nand U1611 (N_1611,N_304,N_36);
nand U1612 (N_1612,N_109,N_52);
and U1613 (N_1613,N_243,N_281);
or U1614 (N_1614,N_85,N_856);
and U1615 (N_1615,N_518,N_708);
nor U1616 (N_1616,N_288,N_924);
or U1617 (N_1617,N_719,N_676);
nor U1618 (N_1618,N_157,N_591);
and U1619 (N_1619,N_942,N_308);
or U1620 (N_1620,N_98,N_458);
or U1621 (N_1621,N_658,N_152);
and U1622 (N_1622,N_6,N_504);
or U1623 (N_1623,N_226,N_367);
and U1624 (N_1624,N_534,N_458);
nor U1625 (N_1625,N_854,N_340);
xor U1626 (N_1626,N_742,N_513);
nand U1627 (N_1627,N_789,N_37);
nand U1628 (N_1628,N_791,N_871);
and U1629 (N_1629,N_443,N_419);
or U1630 (N_1630,N_438,N_831);
or U1631 (N_1631,N_875,N_694);
or U1632 (N_1632,N_253,N_82);
nor U1633 (N_1633,N_411,N_635);
or U1634 (N_1634,N_916,N_359);
nand U1635 (N_1635,N_937,N_685);
nand U1636 (N_1636,N_638,N_811);
and U1637 (N_1637,N_992,N_961);
or U1638 (N_1638,N_51,N_994);
nor U1639 (N_1639,N_825,N_202);
or U1640 (N_1640,N_609,N_258);
nor U1641 (N_1641,N_449,N_200);
nand U1642 (N_1642,N_220,N_368);
nand U1643 (N_1643,N_136,N_699);
nor U1644 (N_1644,N_263,N_609);
and U1645 (N_1645,N_530,N_163);
nand U1646 (N_1646,N_929,N_299);
nor U1647 (N_1647,N_182,N_436);
nor U1648 (N_1648,N_670,N_414);
or U1649 (N_1649,N_44,N_588);
or U1650 (N_1650,N_350,N_636);
or U1651 (N_1651,N_18,N_42);
nor U1652 (N_1652,N_321,N_405);
nand U1653 (N_1653,N_437,N_915);
nor U1654 (N_1654,N_659,N_414);
nor U1655 (N_1655,N_628,N_779);
nor U1656 (N_1656,N_110,N_447);
and U1657 (N_1657,N_846,N_936);
and U1658 (N_1658,N_12,N_470);
and U1659 (N_1659,N_111,N_879);
nor U1660 (N_1660,N_918,N_931);
nand U1661 (N_1661,N_277,N_475);
or U1662 (N_1662,N_15,N_473);
or U1663 (N_1663,N_792,N_605);
nand U1664 (N_1664,N_947,N_539);
and U1665 (N_1665,N_388,N_166);
or U1666 (N_1666,N_508,N_161);
or U1667 (N_1667,N_376,N_1);
nor U1668 (N_1668,N_550,N_202);
and U1669 (N_1669,N_39,N_731);
and U1670 (N_1670,N_146,N_763);
nand U1671 (N_1671,N_142,N_207);
nand U1672 (N_1672,N_307,N_498);
and U1673 (N_1673,N_225,N_279);
nand U1674 (N_1674,N_266,N_616);
nand U1675 (N_1675,N_474,N_114);
or U1676 (N_1676,N_37,N_874);
xor U1677 (N_1677,N_394,N_933);
or U1678 (N_1678,N_527,N_626);
or U1679 (N_1679,N_848,N_811);
and U1680 (N_1680,N_601,N_23);
nand U1681 (N_1681,N_397,N_789);
nor U1682 (N_1682,N_280,N_377);
and U1683 (N_1683,N_370,N_874);
and U1684 (N_1684,N_549,N_793);
nand U1685 (N_1685,N_210,N_286);
or U1686 (N_1686,N_798,N_956);
and U1687 (N_1687,N_364,N_179);
nor U1688 (N_1688,N_825,N_666);
or U1689 (N_1689,N_333,N_118);
or U1690 (N_1690,N_803,N_432);
nor U1691 (N_1691,N_679,N_835);
and U1692 (N_1692,N_470,N_824);
or U1693 (N_1693,N_776,N_131);
nand U1694 (N_1694,N_838,N_625);
and U1695 (N_1695,N_529,N_301);
and U1696 (N_1696,N_25,N_920);
or U1697 (N_1697,N_495,N_137);
or U1698 (N_1698,N_133,N_196);
or U1699 (N_1699,N_91,N_508);
nor U1700 (N_1700,N_485,N_816);
or U1701 (N_1701,N_303,N_922);
nand U1702 (N_1702,N_967,N_246);
nand U1703 (N_1703,N_540,N_747);
nand U1704 (N_1704,N_747,N_368);
or U1705 (N_1705,N_564,N_937);
nand U1706 (N_1706,N_746,N_961);
or U1707 (N_1707,N_413,N_381);
and U1708 (N_1708,N_981,N_468);
and U1709 (N_1709,N_770,N_630);
nand U1710 (N_1710,N_328,N_152);
xor U1711 (N_1711,N_717,N_295);
or U1712 (N_1712,N_603,N_2);
nand U1713 (N_1713,N_657,N_226);
or U1714 (N_1714,N_268,N_233);
nand U1715 (N_1715,N_782,N_642);
nand U1716 (N_1716,N_996,N_558);
and U1717 (N_1717,N_985,N_600);
nor U1718 (N_1718,N_637,N_119);
and U1719 (N_1719,N_573,N_223);
nand U1720 (N_1720,N_418,N_551);
and U1721 (N_1721,N_488,N_846);
nor U1722 (N_1722,N_617,N_122);
or U1723 (N_1723,N_128,N_120);
and U1724 (N_1724,N_665,N_394);
nor U1725 (N_1725,N_587,N_392);
nand U1726 (N_1726,N_207,N_865);
or U1727 (N_1727,N_962,N_603);
nor U1728 (N_1728,N_766,N_519);
or U1729 (N_1729,N_81,N_245);
or U1730 (N_1730,N_91,N_886);
nor U1731 (N_1731,N_556,N_950);
and U1732 (N_1732,N_94,N_870);
or U1733 (N_1733,N_224,N_886);
or U1734 (N_1734,N_264,N_132);
and U1735 (N_1735,N_294,N_873);
or U1736 (N_1736,N_221,N_899);
nand U1737 (N_1737,N_867,N_279);
and U1738 (N_1738,N_663,N_448);
nor U1739 (N_1739,N_619,N_216);
nand U1740 (N_1740,N_296,N_559);
nor U1741 (N_1741,N_624,N_665);
nand U1742 (N_1742,N_259,N_658);
nand U1743 (N_1743,N_215,N_107);
nand U1744 (N_1744,N_974,N_935);
nand U1745 (N_1745,N_440,N_295);
and U1746 (N_1746,N_284,N_339);
nor U1747 (N_1747,N_204,N_582);
nand U1748 (N_1748,N_411,N_248);
and U1749 (N_1749,N_77,N_373);
or U1750 (N_1750,N_414,N_880);
nor U1751 (N_1751,N_302,N_695);
and U1752 (N_1752,N_441,N_419);
and U1753 (N_1753,N_963,N_626);
and U1754 (N_1754,N_523,N_346);
nand U1755 (N_1755,N_150,N_615);
nor U1756 (N_1756,N_279,N_387);
or U1757 (N_1757,N_846,N_262);
nor U1758 (N_1758,N_714,N_940);
nor U1759 (N_1759,N_385,N_291);
or U1760 (N_1760,N_441,N_776);
and U1761 (N_1761,N_697,N_522);
nor U1762 (N_1762,N_626,N_762);
nor U1763 (N_1763,N_643,N_702);
xor U1764 (N_1764,N_760,N_909);
and U1765 (N_1765,N_583,N_519);
xnor U1766 (N_1766,N_678,N_299);
nor U1767 (N_1767,N_549,N_432);
nand U1768 (N_1768,N_575,N_546);
or U1769 (N_1769,N_723,N_370);
and U1770 (N_1770,N_800,N_50);
and U1771 (N_1771,N_882,N_745);
nand U1772 (N_1772,N_294,N_84);
nor U1773 (N_1773,N_11,N_643);
or U1774 (N_1774,N_195,N_553);
and U1775 (N_1775,N_143,N_972);
nand U1776 (N_1776,N_113,N_894);
and U1777 (N_1777,N_137,N_110);
or U1778 (N_1778,N_876,N_342);
and U1779 (N_1779,N_906,N_621);
and U1780 (N_1780,N_407,N_372);
or U1781 (N_1781,N_3,N_679);
nor U1782 (N_1782,N_705,N_723);
nand U1783 (N_1783,N_814,N_781);
nand U1784 (N_1784,N_815,N_555);
or U1785 (N_1785,N_786,N_869);
or U1786 (N_1786,N_819,N_285);
nor U1787 (N_1787,N_813,N_628);
or U1788 (N_1788,N_857,N_480);
and U1789 (N_1789,N_937,N_355);
or U1790 (N_1790,N_547,N_947);
nor U1791 (N_1791,N_286,N_603);
nor U1792 (N_1792,N_339,N_337);
nor U1793 (N_1793,N_315,N_250);
nor U1794 (N_1794,N_988,N_228);
nor U1795 (N_1795,N_142,N_132);
or U1796 (N_1796,N_475,N_44);
nand U1797 (N_1797,N_819,N_537);
nor U1798 (N_1798,N_944,N_385);
nor U1799 (N_1799,N_153,N_958);
or U1800 (N_1800,N_724,N_805);
nor U1801 (N_1801,N_542,N_420);
and U1802 (N_1802,N_985,N_393);
and U1803 (N_1803,N_72,N_177);
nor U1804 (N_1804,N_635,N_829);
nor U1805 (N_1805,N_929,N_956);
nor U1806 (N_1806,N_723,N_105);
nor U1807 (N_1807,N_915,N_774);
nand U1808 (N_1808,N_451,N_238);
or U1809 (N_1809,N_615,N_209);
and U1810 (N_1810,N_507,N_105);
or U1811 (N_1811,N_696,N_190);
nor U1812 (N_1812,N_44,N_575);
or U1813 (N_1813,N_194,N_30);
nand U1814 (N_1814,N_248,N_267);
and U1815 (N_1815,N_211,N_633);
and U1816 (N_1816,N_11,N_993);
or U1817 (N_1817,N_613,N_992);
nor U1818 (N_1818,N_170,N_319);
or U1819 (N_1819,N_852,N_229);
nor U1820 (N_1820,N_333,N_159);
or U1821 (N_1821,N_507,N_559);
or U1822 (N_1822,N_888,N_813);
nand U1823 (N_1823,N_458,N_391);
and U1824 (N_1824,N_12,N_766);
and U1825 (N_1825,N_352,N_216);
nor U1826 (N_1826,N_915,N_277);
nor U1827 (N_1827,N_228,N_982);
and U1828 (N_1828,N_152,N_280);
or U1829 (N_1829,N_891,N_878);
nand U1830 (N_1830,N_706,N_939);
nand U1831 (N_1831,N_979,N_903);
nand U1832 (N_1832,N_434,N_295);
and U1833 (N_1833,N_23,N_360);
and U1834 (N_1834,N_741,N_988);
nor U1835 (N_1835,N_8,N_20);
nor U1836 (N_1836,N_697,N_188);
nand U1837 (N_1837,N_514,N_905);
nand U1838 (N_1838,N_821,N_968);
nor U1839 (N_1839,N_686,N_358);
or U1840 (N_1840,N_855,N_743);
nand U1841 (N_1841,N_89,N_947);
nand U1842 (N_1842,N_770,N_262);
or U1843 (N_1843,N_317,N_683);
nor U1844 (N_1844,N_438,N_830);
and U1845 (N_1845,N_382,N_154);
and U1846 (N_1846,N_167,N_968);
and U1847 (N_1847,N_230,N_577);
and U1848 (N_1848,N_648,N_337);
nor U1849 (N_1849,N_23,N_40);
nand U1850 (N_1850,N_408,N_434);
nor U1851 (N_1851,N_281,N_174);
or U1852 (N_1852,N_888,N_28);
or U1853 (N_1853,N_338,N_513);
nor U1854 (N_1854,N_106,N_881);
nor U1855 (N_1855,N_945,N_992);
nand U1856 (N_1856,N_983,N_760);
xnor U1857 (N_1857,N_136,N_114);
and U1858 (N_1858,N_927,N_859);
nand U1859 (N_1859,N_435,N_649);
and U1860 (N_1860,N_93,N_568);
or U1861 (N_1861,N_645,N_967);
and U1862 (N_1862,N_511,N_620);
or U1863 (N_1863,N_842,N_5);
and U1864 (N_1864,N_781,N_957);
xnor U1865 (N_1865,N_821,N_419);
nor U1866 (N_1866,N_747,N_431);
or U1867 (N_1867,N_206,N_675);
and U1868 (N_1868,N_155,N_179);
xnor U1869 (N_1869,N_165,N_624);
nor U1870 (N_1870,N_205,N_371);
and U1871 (N_1871,N_968,N_698);
and U1872 (N_1872,N_1,N_688);
and U1873 (N_1873,N_327,N_630);
and U1874 (N_1874,N_810,N_607);
or U1875 (N_1875,N_335,N_390);
or U1876 (N_1876,N_832,N_160);
nor U1877 (N_1877,N_574,N_955);
or U1878 (N_1878,N_58,N_718);
nand U1879 (N_1879,N_486,N_843);
nand U1880 (N_1880,N_49,N_29);
and U1881 (N_1881,N_874,N_322);
or U1882 (N_1882,N_94,N_746);
or U1883 (N_1883,N_744,N_749);
nand U1884 (N_1884,N_510,N_284);
or U1885 (N_1885,N_386,N_631);
nand U1886 (N_1886,N_104,N_150);
and U1887 (N_1887,N_20,N_720);
and U1888 (N_1888,N_758,N_840);
or U1889 (N_1889,N_111,N_739);
or U1890 (N_1890,N_240,N_522);
and U1891 (N_1891,N_163,N_311);
nand U1892 (N_1892,N_159,N_58);
nor U1893 (N_1893,N_923,N_792);
and U1894 (N_1894,N_556,N_79);
nand U1895 (N_1895,N_846,N_149);
and U1896 (N_1896,N_605,N_65);
or U1897 (N_1897,N_636,N_295);
or U1898 (N_1898,N_358,N_59);
nand U1899 (N_1899,N_51,N_523);
nand U1900 (N_1900,N_902,N_497);
nand U1901 (N_1901,N_735,N_934);
and U1902 (N_1902,N_895,N_292);
or U1903 (N_1903,N_318,N_630);
nand U1904 (N_1904,N_698,N_309);
nor U1905 (N_1905,N_826,N_116);
or U1906 (N_1906,N_950,N_537);
nand U1907 (N_1907,N_598,N_756);
nor U1908 (N_1908,N_519,N_650);
nand U1909 (N_1909,N_416,N_220);
and U1910 (N_1910,N_178,N_687);
and U1911 (N_1911,N_321,N_675);
nor U1912 (N_1912,N_152,N_829);
and U1913 (N_1913,N_203,N_605);
and U1914 (N_1914,N_66,N_310);
nand U1915 (N_1915,N_113,N_464);
or U1916 (N_1916,N_970,N_934);
or U1917 (N_1917,N_709,N_963);
nor U1918 (N_1918,N_747,N_263);
nand U1919 (N_1919,N_997,N_203);
nor U1920 (N_1920,N_879,N_186);
nor U1921 (N_1921,N_349,N_101);
or U1922 (N_1922,N_41,N_143);
and U1923 (N_1923,N_687,N_867);
and U1924 (N_1924,N_283,N_293);
nor U1925 (N_1925,N_60,N_562);
nor U1926 (N_1926,N_352,N_492);
and U1927 (N_1927,N_929,N_802);
nand U1928 (N_1928,N_948,N_539);
or U1929 (N_1929,N_796,N_540);
nor U1930 (N_1930,N_313,N_859);
and U1931 (N_1931,N_446,N_475);
or U1932 (N_1932,N_19,N_984);
nand U1933 (N_1933,N_702,N_538);
or U1934 (N_1934,N_539,N_863);
or U1935 (N_1935,N_678,N_738);
or U1936 (N_1936,N_975,N_185);
nor U1937 (N_1937,N_183,N_284);
and U1938 (N_1938,N_708,N_528);
and U1939 (N_1939,N_506,N_197);
or U1940 (N_1940,N_602,N_257);
and U1941 (N_1941,N_725,N_978);
and U1942 (N_1942,N_988,N_484);
and U1943 (N_1943,N_138,N_126);
nand U1944 (N_1944,N_897,N_375);
and U1945 (N_1945,N_362,N_808);
and U1946 (N_1946,N_391,N_609);
nand U1947 (N_1947,N_413,N_633);
or U1948 (N_1948,N_589,N_384);
nand U1949 (N_1949,N_191,N_161);
nor U1950 (N_1950,N_30,N_999);
and U1951 (N_1951,N_597,N_990);
nor U1952 (N_1952,N_12,N_977);
xnor U1953 (N_1953,N_439,N_394);
nand U1954 (N_1954,N_837,N_753);
or U1955 (N_1955,N_700,N_514);
nand U1956 (N_1956,N_51,N_960);
nand U1957 (N_1957,N_600,N_230);
or U1958 (N_1958,N_699,N_497);
nand U1959 (N_1959,N_991,N_291);
and U1960 (N_1960,N_895,N_97);
and U1961 (N_1961,N_656,N_345);
and U1962 (N_1962,N_667,N_366);
nand U1963 (N_1963,N_126,N_728);
and U1964 (N_1964,N_897,N_97);
nor U1965 (N_1965,N_275,N_74);
nor U1966 (N_1966,N_425,N_979);
nand U1967 (N_1967,N_857,N_367);
or U1968 (N_1968,N_998,N_874);
nand U1969 (N_1969,N_310,N_977);
nand U1970 (N_1970,N_14,N_815);
or U1971 (N_1971,N_445,N_712);
or U1972 (N_1972,N_284,N_652);
nor U1973 (N_1973,N_354,N_87);
or U1974 (N_1974,N_393,N_477);
nor U1975 (N_1975,N_624,N_562);
and U1976 (N_1976,N_680,N_279);
nand U1977 (N_1977,N_427,N_163);
nand U1978 (N_1978,N_615,N_674);
nand U1979 (N_1979,N_919,N_999);
nor U1980 (N_1980,N_678,N_818);
nand U1981 (N_1981,N_854,N_777);
nor U1982 (N_1982,N_36,N_106);
or U1983 (N_1983,N_462,N_654);
and U1984 (N_1984,N_868,N_221);
nand U1985 (N_1985,N_308,N_708);
or U1986 (N_1986,N_398,N_699);
nor U1987 (N_1987,N_814,N_355);
or U1988 (N_1988,N_683,N_304);
and U1989 (N_1989,N_954,N_830);
or U1990 (N_1990,N_776,N_930);
nand U1991 (N_1991,N_703,N_166);
and U1992 (N_1992,N_834,N_431);
nand U1993 (N_1993,N_991,N_997);
and U1994 (N_1994,N_30,N_23);
or U1995 (N_1995,N_570,N_138);
or U1996 (N_1996,N_56,N_849);
and U1997 (N_1997,N_809,N_996);
or U1998 (N_1998,N_261,N_101);
nand U1999 (N_1999,N_520,N_797);
nor U2000 (N_2000,N_1965,N_1139);
and U2001 (N_2001,N_1629,N_1549);
and U2002 (N_2002,N_1162,N_1964);
nor U2003 (N_2003,N_1967,N_1696);
nand U2004 (N_2004,N_1849,N_1498);
or U2005 (N_2005,N_1485,N_1027);
nor U2006 (N_2006,N_1578,N_1163);
nand U2007 (N_2007,N_1983,N_1368);
or U2008 (N_2008,N_1320,N_1232);
nand U2009 (N_2009,N_1555,N_1581);
nor U2010 (N_2010,N_1376,N_1959);
nand U2011 (N_2011,N_1415,N_1479);
nor U2012 (N_2012,N_1728,N_1272);
and U2013 (N_2013,N_1984,N_1305);
nand U2014 (N_2014,N_1262,N_1781);
nor U2015 (N_2015,N_1921,N_1214);
or U2016 (N_2016,N_1772,N_1987);
or U2017 (N_2017,N_1453,N_1759);
and U2018 (N_2018,N_1803,N_1237);
or U2019 (N_2019,N_1881,N_1534);
nor U2020 (N_2020,N_1186,N_1461);
nor U2021 (N_2021,N_1447,N_1598);
nand U2022 (N_2022,N_1031,N_1934);
nand U2023 (N_2023,N_1033,N_1205);
or U2024 (N_2024,N_1111,N_1559);
nor U2025 (N_2025,N_1301,N_1850);
nor U2026 (N_2026,N_1043,N_1880);
or U2027 (N_2027,N_1502,N_1288);
or U2028 (N_2028,N_1627,N_1411);
and U2029 (N_2029,N_1405,N_1492);
nor U2030 (N_2030,N_1384,N_1594);
nand U2031 (N_2031,N_1805,N_1392);
nor U2032 (N_2032,N_1699,N_1004);
or U2033 (N_2033,N_1532,N_1882);
nor U2034 (N_2034,N_1785,N_1359);
nor U2035 (N_2035,N_1729,N_1653);
and U2036 (N_2036,N_1037,N_1631);
nor U2037 (N_2037,N_1704,N_1654);
or U2038 (N_2038,N_1137,N_1567);
nor U2039 (N_2039,N_1192,N_1593);
nor U2040 (N_2040,N_1830,N_1685);
nand U2041 (N_2041,N_1323,N_1530);
and U2042 (N_2042,N_1480,N_1799);
nand U2043 (N_2043,N_1008,N_1938);
nand U2044 (N_2044,N_1662,N_1933);
and U2045 (N_2045,N_1422,N_1210);
nor U2046 (N_2046,N_1723,N_1292);
and U2047 (N_2047,N_1311,N_1953);
or U2048 (N_2048,N_1143,N_1831);
and U2049 (N_2049,N_1003,N_1331);
or U2050 (N_2050,N_1185,N_1211);
nand U2051 (N_2051,N_1835,N_1448);
or U2052 (N_2052,N_1147,N_1056);
nand U2053 (N_2053,N_1580,N_1219);
nand U2054 (N_2054,N_1416,N_1322);
nand U2055 (N_2055,N_1655,N_1489);
and U2056 (N_2056,N_1700,N_1566);
nand U2057 (N_2057,N_1062,N_1408);
nand U2058 (N_2058,N_1344,N_1092);
and U2059 (N_2059,N_1878,N_1528);
nand U2060 (N_2060,N_1193,N_1628);
or U2061 (N_2061,N_1318,N_1054);
and U2062 (N_2062,N_1079,N_1484);
or U2063 (N_2063,N_1273,N_1619);
nor U2064 (N_2064,N_1464,N_1793);
nand U2065 (N_2065,N_1511,N_1020);
or U2066 (N_2066,N_1533,N_1710);
or U2067 (N_2067,N_1870,N_1516);
and U2068 (N_2068,N_1722,N_1019);
and U2069 (N_2069,N_1382,N_1715);
or U2070 (N_2070,N_1011,N_1081);
nand U2071 (N_2071,N_1109,N_1816);
or U2072 (N_2072,N_1045,N_1885);
nor U2073 (N_2073,N_1267,N_1402);
or U2074 (N_2074,N_1596,N_1616);
nor U2075 (N_2075,N_1960,N_1702);
nor U2076 (N_2076,N_1778,N_1428);
nor U2077 (N_2077,N_1550,N_1689);
nor U2078 (N_2078,N_1971,N_1251);
nand U2079 (N_2079,N_1827,N_1425);
nand U2080 (N_2080,N_1924,N_1949);
or U2081 (N_2081,N_1584,N_1714);
and U2082 (N_2082,N_1014,N_1969);
or U2083 (N_2083,N_1076,N_1023);
nor U2084 (N_2084,N_1086,N_1451);
nand U2085 (N_2085,N_1623,N_1478);
and U2086 (N_2086,N_1200,N_1116);
nand U2087 (N_2087,N_1539,N_1614);
or U2088 (N_2088,N_1907,N_1105);
nand U2089 (N_2089,N_1469,N_1182);
nand U2090 (N_2090,N_1792,N_1026);
nand U2091 (N_2091,N_1632,N_1846);
or U2092 (N_2092,N_1588,N_1776);
and U2093 (N_2093,N_1089,N_1840);
or U2094 (N_2094,N_1687,N_1303);
or U2095 (N_2095,N_1429,N_1753);
nand U2096 (N_2096,N_1366,N_1895);
or U2097 (N_2097,N_1667,N_1352);
nor U2098 (N_2098,N_1042,N_1902);
and U2099 (N_2099,N_1176,N_1737);
nor U2100 (N_2100,N_1823,N_1513);
nand U2101 (N_2101,N_1150,N_1591);
nor U2102 (N_2102,N_1204,N_1286);
or U2103 (N_2103,N_1215,N_1586);
nor U2104 (N_2104,N_1709,N_1634);
or U2105 (N_2105,N_1227,N_1721);
and U2106 (N_2106,N_1196,N_1495);
or U2107 (N_2107,N_1783,N_1678);
nor U2108 (N_2108,N_1865,N_1775);
nand U2109 (N_2109,N_1518,N_1486);
or U2110 (N_2110,N_1526,N_1676);
nand U2111 (N_2111,N_1765,N_1663);
nor U2112 (N_2112,N_1608,N_1963);
or U2113 (N_2113,N_1306,N_1444);
or U2114 (N_2114,N_1679,N_1221);
nand U2115 (N_2115,N_1640,N_1615);
or U2116 (N_2116,N_1674,N_1349);
or U2117 (N_2117,N_1603,N_1957);
or U2118 (N_2118,N_1449,N_1113);
and U2119 (N_2119,N_1929,N_1672);
nor U2120 (N_2120,N_1397,N_1371);
nand U2121 (N_2121,N_1868,N_1355);
nor U2122 (N_2122,N_1597,N_1866);
and U2123 (N_2123,N_1706,N_1841);
nor U2124 (N_2124,N_1183,N_1330);
nand U2125 (N_2125,N_1568,N_1212);
or U2126 (N_2126,N_1304,N_1937);
nand U2127 (N_2127,N_1652,N_1275);
or U2128 (N_2128,N_1930,N_1750);
nand U2129 (N_2129,N_1391,N_1436);
and U2130 (N_2130,N_1546,N_1587);
nor U2131 (N_2131,N_1354,N_1085);
nor U2132 (N_2132,N_1980,N_1263);
nand U2133 (N_2133,N_1158,N_1067);
xor U2134 (N_2134,N_1819,N_1670);
nor U2135 (N_2135,N_1951,N_1133);
nor U2136 (N_2136,N_1357,N_1069);
nand U2137 (N_2137,N_1439,N_1797);
or U2138 (N_2138,N_1916,N_1494);
nor U2139 (N_2139,N_1347,N_1579);
xor U2140 (N_2140,N_1075,N_1038);
and U2141 (N_2141,N_1712,N_1418);
nor U2142 (N_2142,N_1507,N_1256);
nor U2143 (N_2143,N_1350,N_1074);
and U2144 (N_2144,N_1771,N_1159);
nand U2145 (N_2145,N_1861,N_1970);
nor U2146 (N_2146,N_1928,N_1167);
and U2147 (N_2147,N_1954,N_1005);
or U2148 (N_2148,N_1807,N_1543);
and U2149 (N_2149,N_1400,N_1569);
nand U2150 (N_2150,N_1490,N_1034);
nand U2151 (N_2151,N_1442,N_1101);
nor U2152 (N_2152,N_1241,N_1346);
nor U2153 (N_2153,N_1250,N_1601);
nand U2154 (N_2154,N_1246,N_1777);
nand U2155 (N_2155,N_1948,N_1994);
nor U2156 (N_2156,N_1129,N_1072);
and U2157 (N_2157,N_1195,N_1531);
nor U2158 (N_2158,N_1690,N_1590);
nand U2159 (N_2159,N_1972,N_1335);
or U2160 (N_2160,N_1280,N_1319);
nor U2161 (N_2161,N_1225,N_1955);
and U2162 (N_2162,N_1621,N_1973);
nor U2163 (N_2163,N_1500,N_1564);
nor U2164 (N_2164,N_1112,N_1942);
or U2165 (N_2165,N_1844,N_1452);
nor U2166 (N_2166,N_1738,N_1462);
and U2167 (N_2167,N_1595,N_1002);
nand U2168 (N_2168,N_1090,N_1986);
or U2169 (N_2169,N_1474,N_1047);
nor U2170 (N_2170,N_1966,N_1148);
nand U2171 (N_2171,N_1259,N_1604);
or U2172 (N_2172,N_1060,N_1110);
nor U2173 (N_2173,N_1190,N_1958);
nor U2174 (N_2174,N_1134,N_1540);
and U2175 (N_2175,N_1695,N_1433);
nor U2176 (N_2176,N_1410,N_1281);
nand U2177 (N_2177,N_1257,N_1703);
and U2178 (N_2178,N_1454,N_1455);
nor U2179 (N_2179,N_1119,N_1682);
nor U2180 (N_2180,N_1094,N_1693);
nand U2181 (N_2181,N_1735,N_1780);
nor U2182 (N_2182,N_1154,N_1249);
or U2183 (N_2183,N_1097,N_1412);
nand U2184 (N_2184,N_1172,N_1950);
or U2185 (N_2185,N_1363,N_1756);
nand U2186 (N_2186,N_1385,N_1978);
nand U2187 (N_2187,N_1668,N_1909);
or U2188 (N_2188,N_1910,N_1692);
nor U2189 (N_2189,N_1197,N_1658);
or U2190 (N_2190,N_1979,N_1351);
or U2191 (N_2191,N_1188,N_1884);
and U2192 (N_2192,N_1527,N_1510);
or U2193 (N_2193,N_1740,N_1499);
or U2194 (N_2194,N_1763,N_1669);
or U2195 (N_2195,N_1115,N_1893);
and U2196 (N_2196,N_1468,N_1254);
nor U2197 (N_2197,N_1536,N_1173);
nand U2198 (N_2198,N_1261,N_1456);
and U2199 (N_2199,N_1952,N_1913);
nor U2200 (N_2200,N_1218,N_1423);
nand U2201 (N_2201,N_1342,N_1470);
nand U2202 (N_2202,N_1808,N_1570);
or U2203 (N_2203,N_1268,N_1744);
or U2204 (N_2204,N_1684,N_1592);
nor U2205 (N_2205,N_1201,N_1472);
and U2206 (N_2206,N_1477,N_1226);
nor U2207 (N_2207,N_1936,N_1325);
or U2208 (N_2208,N_1923,N_1082);
and U2209 (N_2209,N_1025,N_1968);
and U2210 (N_2210,N_1424,N_1252);
and U2211 (N_2211,N_1997,N_1810);
and U2212 (N_2212,N_1406,N_1369);
nand U2213 (N_2213,N_1758,N_1894);
or U2214 (N_2214,N_1857,N_1639);
nand U2215 (N_2215,N_1488,N_1184);
and U2216 (N_2216,N_1503,N_1548);
nand U2217 (N_2217,N_1786,N_1299);
and U2218 (N_2218,N_1208,N_1605);
and U2219 (N_2219,N_1312,N_1240);
nand U2220 (N_2220,N_1906,N_1838);
nor U2221 (N_2221,N_1073,N_1343);
and U2222 (N_2222,N_1656,N_1381);
nor U2223 (N_2223,N_1845,N_1724);
nor U2224 (N_2224,N_1784,N_1600);
or U2225 (N_2225,N_1044,N_1029);
nand U2226 (N_2226,N_1091,N_1166);
nor U2227 (N_2227,N_1055,N_1675);
and U2228 (N_2228,N_1556,N_1168);
or U2229 (N_2229,N_1234,N_1155);
nand U2230 (N_2230,N_1812,N_1279);
and U2231 (N_2231,N_1927,N_1063);
nor U2232 (N_2232,N_1659,N_1277);
nand U2233 (N_2233,N_1328,N_1388);
nor U2234 (N_2234,N_1160,N_1230);
nor U2235 (N_2235,N_1046,N_1374);
nor U2236 (N_2236,N_1136,N_1242);
nor U2237 (N_2237,N_1883,N_1052);
nand U2238 (N_2238,N_1146,N_1633);
nor U2239 (N_2239,N_1446,N_1859);
nor U2240 (N_2240,N_1367,N_1636);
and U2241 (N_2241,N_1562,N_1879);
or U2242 (N_2242,N_1334,N_1284);
or U2243 (N_2243,N_1806,N_1458);
nand U2244 (N_2244,N_1393,N_1851);
nor U2245 (N_2245,N_1818,N_1657);
nor U2246 (N_2246,N_1773,N_1450);
and U2247 (N_2247,N_1992,N_1058);
nor U2248 (N_2248,N_1701,N_1441);
nor U2249 (N_2249,N_1975,N_1976);
nor U2250 (N_2250,N_1487,N_1749);
or U2251 (N_2251,N_1873,N_1087);
and U2252 (N_2252,N_1544,N_1666);
or U2253 (N_2253,N_1920,N_1216);
or U2254 (N_2254,N_1725,N_1645);
or U2255 (N_2255,N_1040,N_1308);
and U2256 (N_2256,N_1742,N_1716);
or U2257 (N_2257,N_1612,N_1899);
or U2258 (N_2258,N_1169,N_1394);
nand U2259 (N_2259,N_1340,N_1843);
or U2260 (N_2260,N_1779,N_1420);
nor U2261 (N_2261,N_1585,N_1630);
or U2262 (N_2262,N_1705,N_1521);
nand U2263 (N_2263,N_1104,N_1466);
and U2264 (N_2264,N_1985,N_1602);
or U2265 (N_2265,N_1624,N_1083);
nand U2266 (N_2266,N_1289,N_1795);
and U2267 (N_2267,N_1762,N_1419);
or U2268 (N_2268,N_1718,N_1132);
and U2269 (N_2269,N_1329,N_1088);
nand U2270 (N_2270,N_1505,N_1274);
nor U2271 (N_2271,N_1491,N_1788);
or U2272 (N_2272,N_1102,N_1475);
nor U2273 (N_2273,N_1265,N_1457);
nor U2274 (N_2274,N_1825,N_1618);
or U2275 (N_2275,N_1236,N_1348);
nand U2276 (N_2276,N_1814,N_1990);
or U2277 (N_2277,N_1908,N_1686);
nor U2278 (N_2278,N_1125,N_1731);
and U2279 (N_2279,N_1291,N_1199);
nand U2280 (N_2280,N_1260,N_1171);
and U2281 (N_2281,N_1537,N_1151);
nor U2282 (N_2282,N_1837,N_1095);
and U2283 (N_2283,N_1707,N_1413);
nand U2284 (N_2284,N_1012,N_1922);
or U2285 (N_2285,N_1811,N_1370);
and U2286 (N_2286,N_1961,N_1103);
nand U2287 (N_2287,N_1332,N_1789);
and U2288 (N_2288,N_1512,N_1977);
nand U2289 (N_2289,N_1719,N_1571);
or U2290 (N_2290,N_1066,N_1822);
nand U2291 (N_2291,N_1379,N_1123);
and U2292 (N_2292,N_1467,N_1583);
and U2293 (N_2293,N_1180,N_1361);
nor U2294 (N_2294,N_1813,N_1547);
and U2295 (N_2295,N_1313,N_1121);
nor U2296 (N_2296,N_1358,N_1931);
or U2297 (N_2297,N_1515,N_1401);
nand U2298 (N_2298,N_1387,N_1764);
nand U2299 (N_2299,N_1373,N_1755);
nor U2300 (N_2300,N_1287,N_1606);
or U2301 (N_2301,N_1565,N_1770);
or U2302 (N_2302,N_1889,N_1207);
nor U2303 (N_2303,N_1732,N_1691);
nor U2304 (N_2304,N_1124,N_1203);
or U2305 (N_2305,N_1904,N_1622);
nor U2306 (N_2306,N_1736,N_1378);
nand U2307 (N_2307,N_1179,N_1078);
or U2308 (N_2308,N_1222,N_1751);
nand U2309 (N_2309,N_1114,N_1900);
nand U2310 (N_2310,N_1245,N_1673);
or U2311 (N_2311,N_1432,N_1638);
nor U2312 (N_2312,N_1796,N_1403);
nor U2313 (N_2313,N_1981,N_1625);
and U2314 (N_2314,N_1443,N_1372);
or U2315 (N_2315,N_1018,N_1098);
nand U2316 (N_2316,N_1834,N_1582);
nor U2317 (N_2317,N_1238,N_1915);
nand U2318 (N_2318,N_1353,N_1050);
or U2319 (N_2319,N_1962,N_1324);
nor U2320 (N_2320,N_1974,N_1999);
or U2321 (N_2321,N_1080,N_1641);
or U2322 (N_2322,N_1278,N_1496);
or U2323 (N_2323,N_1177,N_1745);
or U2324 (N_2324,N_1535,N_1039);
or U2325 (N_2325,N_1383,N_1142);
nand U2326 (N_2326,N_1314,N_1427);
and U2327 (N_2327,N_1440,N_1741);
or U2328 (N_2328,N_1855,N_1360);
or U2329 (N_2329,N_1522,N_1064);
or U2330 (N_2330,N_1506,N_1465);
or U2331 (N_2331,N_1747,N_1223);
or U2332 (N_2332,N_1084,N_1943);
and U2333 (N_2333,N_1365,N_1228);
or U2334 (N_2334,N_1842,N_1364);
nand U2335 (N_2335,N_1575,N_1181);
and U2336 (N_2336,N_1178,N_1681);
and U2337 (N_2337,N_1926,N_1270);
nand U2338 (N_2338,N_1398,N_1911);
xnor U2339 (N_2339,N_1036,N_1282);
or U2340 (N_2340,N_1804,N_1165);
or U2341 (N_2341,N_1106,N_1501);
nand U2342 (N_2342,N_1000,N_1333);
or U2343 (N_2343,N_1680,N_1414);
or U2344 (N_2344,N_1356,N_1128);
nor U2345 (N_2345,N_1327,N_1220);
or U2346 (N_2346,N_1396,N_1009);
nand U2347 (N_2347,N_1341,N_1892);
nor U2348 (N_2348,N_1613,N_1107);
or U2349 (N_2349,N_1244,N_1239);
and U2350 (N_2350,N_1651,N_1174);
or U2351 (N_2351,N_1130,N_1856);
or U2352 (N_2352,N_1157,N_1828);
nand U2353 (N_2353,N_1646,N_1553);
nor U2354 (N_2354,N_1404,N_1213);
nand U2355 (N_2355,N_1552,N_1170);
and U2356 (N_2356,N_1266,N_1235);
and U2357 (N_2357,N_1126,N_1217);
nand U2358 (N_2358,N_1867,N_1138);
or U2359 (N_2359,N_1068,N_1820);
and U2360 (N_2360,N_1833,N_1677);
or U2361 (N_2361,N_1609,N_1774);
nand U2362 (N_2362,N_1229,N_1497);
and U2363 (N_2363,N_1761,N_1607);
and U2364 (N_2364,N_1149,N_1720);
or U2365 (N_2365,N_1617,N_1471);
and U2366 (N_2366,N_1898,N_1748);
nor U2367 (N_2367,N_1473,N_1946);
nand U2368 (N_2368,N_1848,N_1914);
and U2369 (N_2369,N_1164,N_1529);
and U2370 (N_2370,N_1399,N_1407);
nor U2371 (N_2371,N_1445,N_1483);
or U2372 (N_2372,N_1573,N_1093);
nor U2373 (N_2373,N_1863,N_1649);
nor U2374 (N_2374,N_1853,N_1437);
nor U2375 (N_2375,N_1801,N_1156);
and U2376 (N_2376,N_1599,N_1022);
and U2377 (N_2377,N_1647,N_1919);
or U2378 (N_2378,N_1118,N_1993);
or U2379 (N_2379,N_1610,N_1727);
and U2380 (N_2380,N_1295,N_1708);
and U2381 (N_2381,N_1161,N_1253);
or U2382 (N_2382,N_1336,N_1554);
or U2383 (N_2383,N_1520,N_1191);
nand U2384 (N_2384,N_1611,N_1836);
and U2385 (N_2385,N_1891,N_1460);
nor U2386 (N_2386,N_1665,N_1015);
or U2387 (N_2387,N_1561,N_1525);
nor U2388 (N_2388,N_1264,N_1255);
or U2389 (N_2389,N_1117,N_1194);
nand U2390 (N_2390,N_1875,N_1514);
nor U2391 (N_2391,N_1028,N_1059);
nor U2392 (N_2392,N_1826,N_1872);
nor U2393 (N_2393,N_1989,N_1905);
nor U2394 (N_2394,N_1258,N_1096);
and U2395 (N_2395,N_1637,N_1858);
and U2396 (N_2396,N_1897,N_1996);
and U2397 (N_2397,N_1071,N_1817);
nand U2398 (N_2398,N_1435,N_1852);
or U2399 (N_2399,N_1233,N_1988);
and U2400 (N_2400,N_1459,N_1876);
nand U2401 (N_2401,N_1557,N_1189);
nor U2402 (N_2402,N_1576,N_1053);
nand U2403 (N_2403,N_1635,N_1144);
or U2404 (N_2404,N_1717,N_1560);
nand U2405 (N_2405,N_1296,N_1380);
or U2406 (N_2406,N_1127,N_1896);
nand U2407 (N_2407,N_1202,N_1481);
nor U2408 (N_2408,N_1739,N_1713);
nand U2409 (N_2409,N_1524,N_1829);
nor U2410 (N_2410,N_1757,N_1648);
nand U2411 (N_2411,N_1888,N_1434);
nor U2412 (N_2412,N_1768,N_1297);
nor U2413 (N_2413,N_1935,N_1389);
nand U2414 (N_2414,N_1925,N_1760);
nand U2415 (N_2415,N_1206,N_1944);
or U2416 (N_2416,N_1688,N_1787);
and U2417 (N_2417,N_1298,N_1016);
nor U2418 (N_2418,N_1070,N_1317);
or U2419 (N_2419,N_1509,N_1901);
nor U2420 (N_2420,N_1135,N_1006);
or U2421 (N_2421,N_1890,N_1932);
or U2422 (N_2422,N_1956,N_1290);
or U2423 (N_2423,N_1065,N_1152);
and U2424 (N_2424,N_1991,N_1145);
nor U2425 (N_2425,N_1431,N_1832);
nand U2426 (N_2426,N_1798,N_1493);
nor U2427 (N_2427,N_1545,N_1767);
nand U2428 (N_2428,N_1030,N_1339);
and U2429 (N_2429,N_1698,N_1743);
nor U2430 (N_2430,N_1099,N_1940);
or U2431 (N_2431,N_1057,N_1551);
nor U2432 (N_2432,N_1269,N_1307);
nor U2433 (N_2433,N_1945,N_1995);
or U2434 (N_2434,N_1847,N_1643);
or U2435 (N_2435,N_1815,N_1821);
nand U2436 (N_2436,N_1293,N_1734);
nor U2437 (N_2437,N_1860,N_1276);
nand U2438 (N_2438,N_1886,N_1048);
nand U2439 (N_2439,N_1010,N_1285);
and U2440 (N_2440,N_1800,N_1523);
nor U2441 (N_2441,N_1824,N_1541);
nor U2442 (N_2442,N_1746,N_1912);
nand U2443 (N_2443,N_1542,N_1421);
or U2444 (N_2444,N_1007,N_1001);
or U2445 (N_2445,N_1790,N_1309);
or U2446 (N_2446,N_1917,N_1519);
nor U2447 (N_2447,N_1141,N_1209);
or U2448 (N_2448,N_1642,N_1854);
nand U2449 (N_2449,N_1877,N_1694);
nor U2450 (N_2450,N_1316,N_1733);
or U2451 (N_2451,N_1386,N_1326);
or U2452 (N_2452,N_1041,N_1108);
nand U2453 (N_2453,N_1390,N_1754);
and U2454 (N_2454,N_1315,N_1782);
nand U2455 (N_2455,N_1438,N_1671);
or U2456 (N_2456,N_1021,N_1563);
and U2457 (N_2457,N_1982,N_1409);
nor U2458 (N_2458,N_1310,N_1871);
nor U2459 (N_2459,N_1766,N_1140);
and U2460 (N_2460,N_1187,N_1874);
or U2461 (N_2461,N_1574,N_1794);
and U2462 (N_2462,N_1752,N_1947);
or U2463 (N_2463,N_1711,N_1345);
and U2464 (N_2464,N_1463,N_1869);
nand U2465 (N_2465,N_1664,N_1887);
nor U2466 (N_2466,N_1302,N_1697);
and U2467 (N_2467,N_1175,N_1120);
nand U2468 (N_2468,N_1032,N_1650);
nor U2469 (N_2469,N_1769,N_1482);
nor U2470 (N_2470,N_1049,N_1430);
or U2471 (N_2471,N_1375,N_1283);
and U2472 (N_2472,N_1024,N_1395);
nor U2473 (N_2473,N_1362,N_1300);
nor U2474 (N_2474,N_1271,N_1321);
or U2475 (N_2475,N_1061,N_1504);
nor U2476 (N_2476,N_1538,N_1730);
or U2477 (N_2477,N_1508,N_1100);
or U2478 (N_2478,N_1035,N_1131);
nand U2479 (N_2479,N_1839,N_1294);
or U2480 (N_2480,N_1998,N_1077);
and U2481 (N_2481,N_1247,N_1337);
and U2482 (N_2482,N_1661,N_1683);
and U2483 (N_2483,N_1153,N_1248);
or U2484 (N_2484,N_1426,N_1476);
nand U2485 (N_2485,N_1122,N_1864);
and U2486 (N_2486,N_1791,N_1338);
or U2487 (N_2487,N_1918,N_1013);
and U2488 (N_2488,N_1224,N_1017);
nor U2489 (N_2489,N_1939,N_1941);
nor U2490 (N_2490,N_1644,N_1862);
and U2491 (N_2491,N_1726,N_1243);
nor U2492 (N_2492,N_1377,N_1517);
nor U2493 (N_2493,N_1802,N_1903);
nand U2494 (N_2494,N_1417,N_1660);
nand U2495 (N_2495,N_1572,N_1198);
and U2496 (N_2496,N_1231,N_1809);
xor U2497 (N_2497,N_1589,N_1051);
nand U2498 (N_2498,N_1577,N_1558);
or U2499 (N_2499,N_1626,N_1620);
or U2500 (N_2500,N_1875,N_1116);
or U2501 (N_2501,N_1277,N_1415);
nand U2502 (N_2502,N_1709,N_1508);
and U2503 (N_2503,N_1592,N_1354);
nand U2504 (N_2504,N_1792,N_1431);
and U2505 (N_2505,N_1489,N_1033);
and U2506 (N_2506,N_1505,N_1096);
and U2507 (N_2507,N_1281,N_1264);
nand U2508 (N_2508,N_1950,N_1188);
nor U2509 (N_2509,N_1763,N_1508);
nand U2510 (N_2510,N_1555,N_1499);
nand U2511 (N_2511,N_1970,N_1121);
nor U2512 (N_2512,N_1540,N_1233);
nor U2513 (N_2513,N_1551,N_1677);
and U2514 (N_2514,N_1491,N_1132);
nor U2515 (N_2515,N_1330,N_1231);
or U2516 (N_2516,N_1171,N_1908);
nor U2517 (N_2517,N_1649,N_1021);
nor U2518 (N_2518,N_1805,N_1427);
nor U2519 (N_2519,N_1113,N_1087);
and U2520 (N_2520,N_1972,N_1464);
and U2521 (N_2521,N_1936,N_1391);
or U2522 (N_2522,N_1623,N_1738);
and U2523 (N_2523,N_1439,N_1298);
nor U2524 (N_2524,N_1188,N_1916);
and U2525 (N_2525,N_1954,N_1254);
nor U2526 (N_2526,N_1654,N_1421);
and U2527 (N_2527,N_1725,N_1642);
nand U2528 (N_2528,N_1672,N_1994);
nor U2529 (N_2529,N_1524,N_1013);
and U2530 (N_2530,N_1289,N_1360);
nor U2531 (N_2531,N_1694,N_1227);
or U2532 (N_2532,N_1400,N_1202);
or U2533 (N_2533,N_1973,N_1972);
nand U2534 (N_2534,N_1749,N_1175);
and U2535 (N_2535,N_1346,N_1342);
or U2536 (N_2536,N_1182,N_1300);
nor U2537 (N_2537,N_1389,N_1061);
nor U2538 (N_2538,N_1908,N_1043);
nand U2539 (N_2539,N_1670,N_1050);
nand U2540 (N_2540,N_1113,N_1332);
or U2541 (N_2541,N_1563,N_1337);
or U2542 (N_2542,N_1881,N_1548);
or U2543 (N_2543,N_1701,N_1110);
nor U2544 (N_2544,N_1681,N_1223);
or U2545 (N_2545,N_1087,N_1992);
or U2546 (N_2546,N_1701,N_1934);
nand U2547 (N_2547,N_1979,N_1204);
or U2548 (N_2548,N_1441,N_1660);
or U2549 (N_2549,N_1276,N_1737);
or U2550 (N_2550,N_1993,N_1611);
nand U2551 (N_2551,N_1317,N_1824);
nor U2552 (N_2552,N_1890,N_1843);
nand U2553 (N_2553,N_1915,N_1186);
nand U2554 (N_2554,N_1691,N_1045);
nor U2555 (N_2555,N_1436,N_1295);
and U2556 (N_2556,N_1880,N_1855);
and U2557 (N_2557,N_1536,N_1265);
and U2558 (N_2558,N_1115,N_1887);
nor U2559 (N_2559,N_1390,N_1306);
nor U2560 (N_2560,N_1850,N_1325);
and U2561 (N_2561,N_1803,N_1593);
or U2562 (N_2562,N_1024,N_1460);
nand U2563 (N_2563,N_1192,N_1879);
and U2564 (N_2564,N_1611,N_1687);
or U2565 (N_2565,N_1744,N_1202);
nand U2566 (N_2566,N_1539,N_1872);
and U2567 (N_2567,N_1324,N_1677);
or U2568 (N_2568,N_1259,N_1323);
and U2569 (N_2569,N_1637,N_1841);
and U2570 (N_2570,N_1559,N_1853);
nor U2571 (N_2571,N_1287,N_1547);
or U2572 (N_2572,N_1157,N_1687);
nor U2573 (N_2573,N_1522,N_1849);
nand U2574 (N_2574,N_1277,N_1337);
or U2575 (N_2575,N_1766,N_1084);
nor U2576 (N_2576,N_1787,N_1916);
and U2577 (N_2577,N_1365,N_1896);
and U2578 (N_2578,N_1001,N_1177);
nor U2579 (N_2579,N_1852,N_1693);
nor U2580 (N_2580,N_1117,N_1523);
xnor U2581 (N_2581,N_1015,N_1489);
nand U2582 (N_2582,N_1669,N_1777);
nand U2583 (N_2583,N_1343,N_1898);
nor U2584 (N_2584,N_1848,N_1666);
nor U2585 (N_2585,N_1814,N_1202);
and U2586 (N_2586,N_1578,N_1902);
nand U2587 (N_2587,N_1208,N_1195);
nand U2588 (N_2588,N_1326,N_1808);
or U2589 (N_2589,N_1063,N_1457);
or U2590 (N_2590,N_1792,N_1255);
nand U2591 (N_2591,N_1099,N_1045);
nor U2592 (N_2592,N_1054,N_1981);
and U2593 (N_2593,N_1419,N_1783);
and U2594 (N_2594,N_1657,N_1654);
and U2595 (N_2595,N_1832,N_1449);
nor U2596 (N_2596,N_1802,N_1366);
or U2597 (N_2597,N_1788,N_1607);
and U2598 (N_2598,N_1189,N_1228);
or U2599 (N_2599,N_1854,N_1467);
nor U2600 (N_2600,N_1757,N_1926);
nand U2601 (N_2601,N_1246,N_1638);
and U2602 (N_2602,N_1245,N_1815);
nor U2603 (N_2603,N_1336,N_1167);
and U2604 (N_2604,N_1473,N_1369);
or U2605 (N_2605,N_1976,N_1381);
nand U2606 (N_2606,N_1162,N_1386);
and U2607 (N_2607,N_1918,N_1943);
and U2608 (N_2608,N_1608,N_1381);
nor U2609 (N_2609,N_1310,N_1089);
nor U2610 (N_2610,N_1850,N_1088);
nor U2611 (N_2611,N_1479,N_1892);
nor U2612 (N_2612,N_1585,N_1577);
and U2613 (N_2613,N_1783,N_1273);
and U2614 (N_2614,N_1946,N_1990);
and U2615 (N_2615,N_1706,N_1210);
nor U2616 (N_2616,N_1236,N_1088);
nor U2617 (N_2617,N_1656,N_1606);
nand U2618 (N_2618,N_1366,N_1397);
or U2619 (N_2619,N_1669,N_1611);
xnor U2620 (N_2620,N_1201,N_1165);
nor U2621 (N_2621,N_1901,N_1423);
nor U2622 (N_2622,N_1794,N_1987);
nor U2623 (N_2623,N_1553,N_1288);
nor U2624 (N_2624,N_1869,N_1670);
or U2625 (N_2625,N_1973,N_1397);
or U2626 (N_2626,N_1876,N_1175);
nor U2627 (N_2627,N_1539,N_1914);
nor U2628 (N_2628,N_1702,N_1286);
and U2629 (N_2629,N_1031,N_1529);
and U2630 (N_2630,N_1748,N_1742);
nor U2631 (N_2631,N_1035,N_1068);
and U2632 (N_2632,N_1250,N_1959);
and U2633 (N_2633,N_1292,N_1474);
nor U2634 (N_2634,N_1028,N_1450);
nand U2635 (N_2635,N_1843,N_1794);
and U2636 (N_2636,N_1915,N_1663);
nand U2637 (N_2637,N_1403,N_1172);
nand U2638 (N_2638,N_1975,N_1423);
or U2639 (N_2639,N_1966,N_1670);
or U2640 (N_2640,N_1298,N_1126);
or U2641 (N_2641,N_1379,N_1554);
and U2642 (N_2642,N_1024,N_1193);
nor U2643 (N_2643,N_1424,N_1408);
nor U2644 (N_2644,N_1205,N_1408);
nand U2645 (N_2645,N_1079,N_1927);
nor U2646 (N_2646,N_1417,N_1343);
nor U2647 (N_2647,N_1679,N_1535);
or U2648 (N_2648,N_1299,N_1123);
nand U2649 (N_2649,N_1470,N_1500);
nand U2650 (N_2650,N_1187,N_1540);
or U2651 (N_2651,N_1225,N_1126);
nand U2652 (N_2652,N_1079,N_1662);
nand U2653 (N_2653,N_1053,N_1968);
nor U2654 (N_2654,N_1678,N_1759);
and U2655 (N_2655,N_1018,N_1974);
or U2656 (N_2656,N_1858,N_1261);
and U2657 (N_2657,N_1878,N_1300);
nand U2658 (N_2658,N_1573,N_1635);
and U2659 (N_2659,N_1101,N_1436);
nor U2660 (N_2660,N_1173,N_1252);
nand U2661 (N_2661,N_1436,N_1648);
or U2662 (N_2662,N_1524,N_1319);
nand U2663 (N_2663,N_1949,N_1023);
nand U2664 (N_2664,N_1391,N_1592);
nand U2665 (N_2665,N_1176,N_1278);
or U2666 (N_2666,N_1979,N_1614);
and U2667 (N_2667,N_1724,N_1140);
nand U2668 (N_2668,N_1028,N_1215);
nand U2669 (N_2669,N_1003,N_1213);
nand U2670 (N_2670,N_1424,N_1533);
nor U2671 (N_2671,N_1830,N_1717);
nor U2672 (N_2672,N_1734,N_1618);
or U2673 (N_2673,N_1803,N_1490);
nand U2674 (N_2674,N_1517,N_1557);
and U2675 (N_2675,N_1749,N_1997);
or U2676 (N_2676,N_1299,N_1642);
nand U2677 (N_2677,N_1109,N_1820);
nand U2678 (N_2678,N_1194,N_1205);
nor U2679 (N_2679,N_1137,N_1669);
nor U2680 (N_2680,N_1618,N_1610);
nand U2681 (N_2681,N_1362,N_1282);
and U2682 (N_2682,N_1410,N_1305);
nor U2683 (N_2683,N_1529,N_1854);
or U2684 (N_2684,N_1123,N_1329);
nor U2685 (N_2685,N_1306,N_1557);
nor U2686 (N_2686,N_1202,N_1193);
and U2687 (N_2687,N_1872,N_1392);
or U2688 (N_2688,N_1756,N_1578);
and U2689 (N_2689,N_1373,N_1218);
nand U2690 (N_2690,N_1091,N_1226);
and U2691 (N_2691,N_1784,N_1895);
nand U2692 (N_2692,N_1194,N_1277);
nor U2693 (N_2693,N_1324,N_1633);
and U2694 (N_2694,N_1668,N_1289);
and U2695 (N_2695,N_1266,N_1595);
nand U2696 (N_2696,N_1946,N_1386);
nor U2697 (N_2697,N_1823,N_1339);
or U2698 (N_2698,N_1168,N_1826);
nor U2699 (N_2699,N_1657,N_1660);
or U2700 (N_2700,N_1123,N_1655);
and U2701 (N_2701,N_1450,N_1362);
nand U2702 (N_2702,N_1870,N_1795);
and U2703 (N_2703,N_1167,N_1770);
nand U2704 (N_2704,N_1872,N_1218);
nor U2705 (N_2705,N_1103,N_1442);
and U2706 (N_2706,N_1699,N_1952);
and U2707 (N_2707,N_1727,N_1825);
nor U2708 (N_2708,N_1334,N_1664);
or U2709 (N_2709,N_1232,N_1928);
and U2710 (N_2710,N_1539,N_1522);
and U2711 (N_2711,N_1671,N_1169);
and U2712 (N_2712,N_1944,N_1683);
or U2713 (N_2713,N_1421,N_1758);
nand U2714 (N_2714,N_1934,N_1454);
nand U2715 (N_2715,N_1042,N_1084);
nor U2716 (N_2716,N_1121,N_1759);
nand U2717 (N_2717,N_1528,N_1562);
or U2718 (N_2718,N_1641,N_1100);
nor U2719 (N_2719,N_1538,N_1583);
or U2720 (N_2720,N_1206,N_1383);
or U2721 (N_2721,N_1729,N_1940);
and U2722 (N_2722,N_1906,N_1936);
and U2723 (N_2723,N_1482,N_1574);
and U2724 (N_2724,N_1840,N_1256);
nor U2725 (N_2725,N_1925,N_1630);
and U2726 (N_2726,N_1422,N_1789);
or U2727 (N_2727,N_1488,N_1607);
and U2728 (N_2728,N_1730,N_1194);
xor U2729 (N_2729,N_1541,N_1838);
or U2730 (N_2730,N_1306,N_1961);
nand U2731 (N_2731,N_1380,N_1483);
nor U2732 (N_2732,N_1882,N_1089);
nand U2733 (N_2733,N_1123,N_1369);
and U2734 (N_2734,N_1658,N_1872);
and U2735 (N_2735,N_1319,N_1035);
nand U2736 (N_2736,N_1271,N_1022);
nand U2737 (N_2737,N_1873,N_1434);
nor U2738 (N_2738,N_1672,N_1106);
nand U2739 (N_2739,N_1944,N_1190);
or U2740 (N_2740,N_1128,N_1575);
nor U2741 (N_2741,N_1685,N_1089);
nor U2742 (N_2742,N_1133,N_1643);
and U2743 (N_2743,N_1359,N_1047);
nand U2744 (N_2744,N_1913,N_1848);
or U2745 (N_2745,N_1796,N_1750);
and U2746 (N_2746,N_1692,N_1086);
or U2747 (N_2747,N_1871,N_1820);
and U2748 (N_2748,N_1996,N_1147);
nand U2749 (N_2749,N_1453,N_1431);
nor U2750 (N_2750,N_1674,N_1188);
and U2751 (N_2751,N_1523,N_1846);
nand U2752 (N_2752,N_1615,N_1778);
nand U2753 (N_2753,N_1293,N_1442);
or U2754 (N_2754,N_1642,N_1465);
or U2755 (N_2755,N_1815,N_1044);
or U2756 (N_2756,N_1398,N_1217);
or U2757 (N_2757,N_1769,N_1815);
and U2758 (N_2758,N_1430,N_1956);
nand U2759 (N_2759,N_1537,N_1720);
nand U2760 (N_2760,N_1040,N_1450);
or U2761 (N_2761,N_1573,N_1651);
nand U2762 (N_2762,N_1792,N_1052);
or U2763 (N_2763,N_1892,N_1458);
nand U2764 (N_2764,N_1295,N_1935);
or U2765 (N_2765,N_1468,N_1804);
nand U2766 (N_2766,N_1996,N_1759);
or U2767 (N_2767,N_1587,N_1450);
nor U2768 (N_2768,N_1392,N_1108);
nand U2769 (N_2769,N_1195,N_1693);
and U2770 (N_2770,N_1786,N_1266);
nor U2771 (N_2771,N_1302,N_1466);
or U2772 (N_2772,N_1745,N_1361);
or U2773 (N_2773,N_1779,N_1668);
nand U2774 (N_2774,N_1479,N_1863);
or U2775 (N_2775,N_1627,N_1239);
nand U2776 (N_2776,N_1716,N_1809);
and U2777 (N_2777,N_1665,N_1977);
and U2778 (N_2778,N_1735,N_1702);
nor U2779 (N_2779,N_1274,N_1348);
nand U2780 (N_2780,N_1963,N_1872);
or U2781 (N_2781,N_1776,N_1068);
and U2782 (N_2782,N_1704,N_1313);
nor U2783 (N_2783,N_1442,N_1212);
and U2784 (N_2784,N_1992,N_1066);
nand U2785 (N_2785,N_1712,N_1544);
nor U2786 (N_2786,N_1887,N_1205);
or U2787 (N_2787,N_1676,N_1922);
and U2788 (N_2788,N_1814,N_1761);
nor U2789 (N_2789,N_1157,N_1499);
nand U2790 (N_2790,N_1141,N_1048);
or U2791 (N_2791,N_1648,N_1935);
nand U2792 (N_2792,N_1660,N_1798);
nand U2793 (N_2793,N_1307,N_1207);
nor U2794 (N_2794,N_1751,N_1962);
nand U2795 (N_2795,N_1548,N_1490);
and U2796 (N_2796,N_1291,N_1155);
and U2797 (N_2797,N_1878,N_1181);
or U2798 (N_2798,N_1044,N_1801);
and U2799 (N_2799,N_1808,N_1952);
nand U2800 (N_2800,N_1350,N_1757);
nand U2801 (N_2801,N_1543,N_1823);
or U2802 (N_2802,N_1093,N_1065);
nor U2803 (N_2803,N_1614,N_1821);
nand U2804 (N_2804,N_1784,N_1608);
nor U2805 (N_2805,N_1079,N_1138);
nor U2806 (N_2806,N_1857,N_1684);
nor U2807 (N_2807,N_1125,N_1027);
xor U2808 (N_2808,N_1643,N_1911);
and U2809 (N_2809,N_1011,N_1693);
and U2810 (N_2810,N_1006,N_1627);
or U2811 (N_2811,N_1286,N_1192);
nand U2812 (N_2812,N_1993,N_1102);
and U2813 (N_2813,N_1574,N_1183);
and U2814 (N_2814,N_1488,N_1484);
and U2815 (N_2815,N_1439,N_1559);
nor U2816 (N_2816,N_1938,N_1088);
or U2817 (N_2817,N_1180,N_1372);
or U2818 (N_2818,N_1216,N_1638);
and U2819 (N_2819,N_1941,N_1690);
or U2820 (N_2820,N_1493,N_1570);
or U2821 (N_2821,N_1018,N_1063);
nand U2822 (N_2822,N_1122,N_1635);
or U2823 (N_2823,N_1749,N_1488);
and U2824 (N_2824,N_1061,N_1640);
nor U2825 (N_2825,N_1202,N_1636);
nor U2826 (N_2826,N_1154,N_1692);
xnor U2827 (N_2827,N_1592,N_1904);
and U2828 (N_2828,N_1150,N_1024);
and U2829 (N_2829,N_1507,N_1210);
nand U2830 (N_2830,N_1332,N_1723);
and U2831 (N_2831,N_1539,N_1537);
nand U2832 (N_2832,N_1454,N_1701);
nor U2833 (N_2833,N_1436,N_1833);
and U2834 (N_2834,N_1776,N_1188);
or U2835 (N_2835,N_1270,N_1615);
or U2836 (N_2836,N_1474,N_1418);
nand U2837 (N_2837,N_1411,N_1317);
nor U2838 (N_2838,N_1335,N_1743);
nor U2839 (N_2839,N_1113,N_1211);
nor U2840 (N_2840,N_1180,N_1426);
nor U2841 (N_2841,N_1321,N_1982);
or U2842 (N_2842,N_1045,N_1387);
nand U2843 (N_2843,N_1639,N_1608);
or U2844 (N_2844,N_1759,N_1442);
or U2845 (N_2845,N_1243,N_1077);
or U2846 (N_2846,N_1031,N_1071);
nand U2847 (N_2847,N_1337,N_1477);
nand U2848 (N_2848,N_1611,N_1780);
or U2849 (N_2849,N_1832,N_1865);
or U2850 (N_2850,N_1769,N_1958);
nand U2851 (N_2851,N_1732,N_1605);
and U2852 (N_2852,N_1840,N_1826);
nand U2853 (N_2853,N_1049,N_1082);
and U2854 (N_2854,N_1591,N_1085);
or U2855 (N_2855,N_1018,N_1409);
nor U2856 (N_2856,N_1723,N_1643);
nand U2857 (N_2857,N_1086,N_1625);
or U2858 (N_2858,N_1567,N_1757);
nor U2859 (N_2859,N_1879,N_1889);
nand U2860 (N_2860,N_1697,N_1204);
nor U2861 (N_2861,N_1049,N_1048);
nand U2862 (N_2862,N_1651,N_1992);
or U2863 (N_2863,N_1630,N_1668);
nor U2864 (N_2864,N_1697,N_1719);
or U2865 (N_2865,N_1254,N_1694);
or U2866 (N_2866,N_1080,N_1280);
nand U2867 (N_2867,N_1394,N_1893);
or U2868 (N_2868,N_1512,N_1514);
nand U2869 (N_2869,N_1685,N_1268);
nor U2870 (N_2870,N_1499,N_1896);
nand U2871 (N_2871,N_1981,N_1883);
and U2872 (N_2872,N_1403,N_1662);
or U2873 (N_2873,N_1279,N_1253);
and U2874 (N_2874,N_1144,N_1199);
nand U2875 (N_2875,N_1239,N_1186);
nand U2876 (N_2876,N_1140,N_1356);
nand U2877 (N_2877,N_1247,N_1936);
and U2878 (N_2878,N_1127,N_1386);
and U2879 (N_2879,N_1412,N_1041);
nor U2880 (N_2880,N_1926,N_1861);
or U2881 (N_2881,N_1782,N_1374);
and U2882 (N_2882,N_1401,N_1030);
nand U2883 (N_2883,N_1963,N_1567);
and U2884 (N_2884,N_1746,N_1012);
or U2885 (N_2885,N_1228,N_1939);
nor U2886 (N_2886,N_1043,N_1249);
nand U2887 (N_2887,N_1073,N_1126);
or U2888 (N_2888,N_1722,N_1864);
nor U2889 (N_2889,N_1819,N_1181);
nor U2890 (N_2890,N_1747,N_1165);
nor U2891 (N_2891,N_1198,N_1841);
and U2892 (N_2892,N_1674,N_1735);
nor U2893 (N_2893,N_1147,N_1757);
and U2894 (N_2894,N_1425,N_1132);
xnor U2895 (N_2895,N_1845,N_1066);
nor U2896 (N_2896,N_1145,N_1801);
and U2897 (N_2897,N_1212,N_1936);
or U2898 (N_2898,N_1177,N_1223);
or U2899 (N_2899,N_1710,N_1705);
and U2900 (N_2900,N_1799,N_1549);
and U2901 (N_2901,N_1671,N_1184);
or U2902 (N_2902,N_1140,N_1933);
or U2903 (N_2903,N_1024,N_1884);
nand U2904 (N_2904,N_1860,N_1959);
nand U2905 (N_2905,N_1550,N_1970);
or U2906 (N_2906,N_1034,N_1552);
and U2907 (N_2907,N_1933,N_1976);
and U2908 (N_2908,N_1632,N_1039);
nor U2909 (N_2909,N_1114,N_1001);
and U2910 (N_2910,N_1100,N_1289);
nor U2911 (N_2911,N_1846,N_1722);
and U2912 (N_2912,N_1489,N_1564);
and U2913 (N_2913,N_1968,N_1347);
and U2914 (N_2914,N_1484,N_1793);
or U2915 (N_2915,N_1793,N_1440);
or U2916 (N_2916,N_1810,N_1908);
nor U2917 (N_2917,N_1603,N_1911);
and U2918 (N_2918,N_1402,N_1816);
and U2919 (N_2919,N_1330,N_1964);
or U2920 (N_2920,N_1927,N_1774);
and U2921 (N_2921,N_1108,N_1411);
and U2922 (N_2922,N_1173,N_1315);
or U2923 (N_2923,N_1959,N_1284);
nor U2924 (N_2924,N_1698,N_1012);
and U2925 (N_2925,N_1157,N_1483);
nand U2926 (N_2926,N_1632,N_1545);
nand U2927 (N_2927,N_1223,N_1741);
and U2928 (N_2928,N_1330,N_1439);
and U2929 (N_2929,N_1508,N_1448);
and U2930 (N_2930,N_1894,N_1780);
nor U2931 (N_2931,N_1454,N_1552);
and U2932 (N_2932,N_1434,N_1528);
nor U2933 (N_2933,N_1357,N_1668);
and U2934 (N_2934,N_1966,N_1972);
nand U2935 (N_2935,N_1374,N_1592);
and U2936 (N_2936,N_1724,N_1923);
nor U2937 (N_2937,N_1427,N_1481);
or U2938 (N_2938,N_1450,N_1342);
nand U2939 (N_2939,N_1956,N_1097);
nand U2940 (N_2940,N_1997,N_1611);
nor U2941 (N_2941,N_1672,N_1688);
or U2942 (N_2942,N_1864,N_1364);
nand U2943 (N_2943,N_1511,N_1536);
or U2944 (N_2944,N_1126,N_1241);
or U2945 (N_2945,N_1307,N_1682);
nor U2946 (N_2946,N_1585,N_1523);
and U2947 (N_2947,N_1763,N_1870);
or U2948 (N_2948,N_1289,N_1674);
and U2949 (N_2949,N_1151,N_1466);
and U2950 (N_2950,N_1864,N_1380);
nand U2951 (N_2951,N_1814,N_1383);
and U2952 (N_2952,N_1159,N_1867);
nand U2953 (N_2953,N_1362,N_1755);
nor U2954 (N_2954,N_1941,N_1973);
nor U2955 (N_2955,N_1907,N_1882);
and U2956 (N_2956,N_1086,N_1235);
and U2957 (N_2957,N_1950,N_1415);
nor U2958 (N_2958,N_1312,N_1889);
nor U2959 (N_2959,N_1849,N_1846);
or U2960 (N_2960,N_1866,N_1527);
nand U2961 (N_2961,N_1656,N_1891);
nand U2962 (N_2962,N_1159,N_1717);
and U2963 (N_2963,N_1360,N_1282);
nor U2964 (N_2964,N_1376,N_1676);
nand U2965 (N_2965,N_1805,N_1002);
nor U2966 (N_2966,N_1258,N_1568);
nor U2967 (N_2967,N_1937,N_1529);
nand U2968 (N_2968,N_1466,N_1499);
and U2969 (N_2969,N_1858,N_1435);
nand U2970 (N_2970,N_1624,N_1693);
and U2971 (N_2971,N_1282,N_1640);
nor U2972 (N_2972,N_1177,N_1087);
nand U2973 (N_2973,N_1458,N_1390);
nor U2974 (N_2974,N_1461,N_1051);
xnor U2975 (N_2975,N_1337,N_1442);
nor U2976 (N_2976,N_1151,N_1148);
nand U2977 (N_2977,N_1211,N_1312);
nand U2978 (N_2978,N_1677,N_1210);
or U2979 (N_2979,N_1434,N_1985);
nand U2980 (N_2980,N_1651,N_1252);
and U2981 (N_2981,N_1135,N_1786);
nand U2982 (N_2982,N_1242,N_1908);
or U2983 (N_2983,N_1289,N_1352);
nor U2984 (N_2984,N_1156,N_1033);
and U2985 (N_2985,N_1812,N_1469);
or U2986 (N_2986,N_1969,N_1071);
nor U2987 (N_2987,N_1416,N_1817);
nand U2988 (N_2988,N_1429,N_1300);
nand U2989 (N_2989,N_1720,N_1692);
nor U2990 (N_2990,N_1135,N_1538);
or U2991 (N_2991,N_1826,N_1016);
nor U2992 (N_2992,N_1376,N_1583);
or U2993 (N_2993,N_1083,N_1862);
nand U2994 (N_2994,N_1781,N_1461);
nor U2995 (N_2995,N_1062,N_1253);
nand U2996 (N_2996,N_1517,N_1222);
nand U2997 (N_2997,N_1200,N_1129);
and U2998 (N_2998,N_1299,N_1348);
nor U2999 (N_2999,N_1956,N_1487);
nor UO_0 (O_0,N_2471,N_2310);
and UO_1 (O_1,N_2600,N_2014);
nand UO_2 (O_2,N_2856,N_2671);
nor UO_3 (O_3,N_2392,N_2920);
nand UO_4 (O_4,N_2272,N_2435);
or UO_5 (O_5,N_2874,N_2121);
and UO_6 (O_6,N_2794,N_2726);
nor UO_7 (O_7,N_2728,N_2844);
and UO_8 (O_8,N_2102,N_2253);
and UO_9 (O_9,N_2934,N_2501);
nand UO_10 (O_10,N_2798,N_2936);
or UO_11 (O_11,N_2577,N_2060);
nand UO_12 (O_12,N_2507,N_2927);
nor UO_13 (O_13,N_2169,N_2543);
xor UO_14 (O_14,N_2480,N_2258);
nand UO_15 (O_15,N_2767,N_2656);
and UO_16 (O_16,N_2382,N_2907);
and UO_17 (O_17,N_2911,N_2645);
or UO_18 (O_18,N_2974,N_2181);
or UO_19 (O_19,N_2654,N_2597);
or UO_20 (O_20,N_2700,N_2260);
or UO_21 (O_21,N_2208,N_2815);
and UO_22 (O_22,N_2407,N_2538);
nor UO_23 (O_23,N_2139,N_2192);
nor UO_24 (O_24,N_2360,N_2097);
nor UO_25 (O_25,N_2793,N_2883);
or UO_26 (O_26,N_2216,N_2116);
nand UO_27 (O_27,N_2224,N_2147);
nor UO_28 (O_28,N_2675,N_2799);
or UO_29 (O_29,N_2800,N_2063);
and UO_30 (O_30,N_2344,N_2298);
nor UO_31 (O_31,N_2935,N_2394);
nor UO_32 (O_32,N_2493,N_2648);
or UO_33 (O_33,N_2765,N_2595);
nand UO_34 (O_34,N_2495,N_2980);
or UO_35 (O_35,N_2334,N_2458);
or UO_36 (O_36,N_2960,N_2246);
nor UO_37 (O_37,N_2959,N_2488);
or UO_38 (O_38,N_2894,N_2895);
nor UO_39 (O_39,N_2022,N_2668);
nand UO_40 (O_40,N_2696,N_2770);
nor UO_41 (O_41,N_2066,N_2052);
and UO_42 (O_42,N_2954,N_2876);
nor UO_43 (O_43,N_2418,N_2603);
nor UO_44 (O_44,N_2631,N_2914);
and UO_45 (O_45,N_2313,N_2242);
nand UO_46 (O_46,N_2393,N_2406);
and UO_47 (O_47,N_2463,N_2835);
nor UO_48 (O_48,N_2932,N_2257);
and UO_49 (O_49,N_2346,N_2170);
or UO_50 (O_50,N_2624,N_2602);
or UO_51 (O_51,N_2614,N_2667);
or UO_52 (O_52,N_2905,N_2628);
or UO_53 (O_53,N_2479,N_2664);
or UO_54 (O_54,N_2620,N_2008);
or UO_55 (O_55,N_2723,N_2129);
nor UO_56 (O_56,N_2733,N_2811);
nor UO_57 (O_57,N_2613,N_2150);
or UO_58 (O_58,N_2476,N_2193);
or UO_59 (O_59,N_2683,N_2969);
nor UO_60 (O_60,N_2026,N_2611);
nor UO_61 (O_61,N_2531,N_2437);
and UO_62 (O_62,N_2381,N_2941);
xor UO_63 (O_63,N_2788,N_2474);
nor UO_64 (O_64,N_2366,N_2098);
nor UO_65 (O_65,N_2790,N_2740);
nor UO_66 (O_66,N_2144,N_2870);
and UO_67 (O_67,N_2206,N_2011);
nand UO_68 (O_68,N_2890,N_2515);
nor UO_69 (O_69,N_2957,N_2692);
or UO_70 (O_70,N_2962,N_2842);
xnor UO_71 (O_71,N_2068,N_2402);
nand UO_72 (O_72,N_2689,N_2455);
and UO_73 (O_73,N_2563,N_2293);
or UO_74 (O_74,N_2203,N_2412);
nor UO_75 (O_75,N_2512,N_2235);
and UO_76 (O_76,N_2362,N_2076);
nor UO_77 (O_77,N_2106,N_2358);
nand UO_78 (O_78,N_2442,N_2204);
nand UO_79 (O_79,N_2530,N_2223);
nor UO_80 (O_80,N_2697,N_2998);
or UO_81 (O_81,N_2384,N_2288);
and UO_82 (O_82,N_2274,N_2695);
and UO_83 (O_83,N_2556,N_2137);
nand UO_84 (O_84,N_2179,N_2018);
nor UO_85 (O_85,N_2632,N_2923);
nand UO_86 (O_86,N_2847,N_2649);
and UO_87 (O_87,N_2320,N_2028);
and UO_88 (O_88,N_2329,N_2789);
nor UO_89 (O_89,N_2988,N_2973);
or UO_90 (O_90,N_2503,N_2759);
and UO_91 (O_91,N_2389,N_2713);
nand UO_92 (O_92,N_2627,N_2286);
or UO_93 (O_93,N_2209,N_2825);
nor UO_94 (O_94,N_2449,N_2862);
or UO_95 (O_95,N_2809,N_2783);
or UO_96 (O_96,N_2283,N_2184);
or UO_97 (O_97,N_2079,N_2860);
nand UO_98 (O_98,N_2774,N_2466);
nand UO_99 (O_99,N_2639,N_2231);
nand UO_100 (O_100,N_2889,N_2415);
or UO_101 (O_101,N_2454,N_2157);
nor UO_102 (O_102,N_2254,N_2846);
and UO_103 (O_103,N_2432,N_2222);
nand UO_104 (O_104,N_2071,N_2427);
or UO_105 (O_105,N_2964,N_2250);
and UO_106 (O_106,N_2496,N_2295);
nor UO_107 (O_107,N_2043,N_2307);
or UO_108 (O_108,N_2279,N_2804);
or UO_109 (O_109,N_2325,N_2673);
nand UO_110 (O_110,N_2494,N_2900);
nor UO_111 (O_111,N_2745,N_2153);
nand UO_112 (O_112,N_2898,N_2186);
xnor UO_113 (O_113,N_2044,N_2081);
nand UO_114 (O_114,N_2785,N_2075);
and UO_115 (O_115,N_2984,N_2239);
nand UO_116 (O_116,N_2067,N_2126);
or UO_117 (O_117,N_2269,N_2891);
or UO_118 (O_118,N_2665,N_2688);
or UO_119 (O_119,N_2408,N_2211);
or UO_120 (O_120,N_2359,N_2172);
nand UO_121 (O_121,N_2433,N_2981);
nand UO_122 (O_122,N_2576,N_2951);
and UO_123 (O_123,N_2796,N_2776);
or UO_124 (O_124,N_2875,N_2606);
and UO_125 (O_125,N_2490,N_2566);
and UO_126 (O_126,N_2024,N_2083);
nor UO_127 (O_127,N_2583,N_2963);
nand UO_128 (O_128,N_2766,N_2048);
and UO_129 (O_129,N_2252,N_2428);
or UO_130 (O_130,N_2459,N_2977);
nand UO_131 (O_131,N_2299,N_2489);
and UO_132 (O_132,N_2284,N_2212);
and UO_133 (O_133,N_2735,N_2037);
or UO_134 (O_134,N_2534,N_2089);
nor UO_135 (O_135,N_2722,N_2119);
nand UO_136 (O_136,N_2548,N_2475);
and UO_137 (O_137,N_2705,N_2033);
or UO_138 (O_138,N_2699,N_2646);
and UO_139 (O_139,N_2737,N_2338);
nand UO_140 (O_140,N_2651,N_2240);
or UO_141 (O_141,N_2278,N_2180);
or UO_142 (O_142,N_2040,N_2041);
nand UO_143 (O_143,N_2485,N_2727);
and UO_144 (O_144,N_2472,N_2464);
and UO_145 (O_145,N_2879,N_2130);
nand UO_146 (O_146,N_2808,N_2107);
nor UO_147 (O_147,N_2850,N_2568);
or UO_148 (O_148,N_2542,N_2514);
or UO_149 (O_149,N_2550,N_2837);
or UO_150 (O_150,N_2422,N_2363);
or UO_151 (O_151,N_2443,N_2191);
and UO_152 (O_152,N_2290,N_2520);
or UO_153 (O_153,N_2950,N_2087);
and UO_154 (O_154,N_2902,N_2562);
or UO_155 (O_155,N_2970,N_2677);
and UO_156 (O_156,N_2537,N_2516);
or UO_157 (O_157,N_2376,N_2527);
nor UO_158 (O_158,N_2061,N_2262);
nand UO_159 (O_159,N_2016,N_2831);
and UO_160 (O_160,N_2824,N_2540);
nor UO_161 (O_161,N_2747,N_2084);
nor UO_162 (O_162,N_2975,N_2806);
and UO_163 (O_163,N_2468,N_2917);
nand UO_164 (O_164,N_2072,N_2642);
nor UO_165 (O_165,N_2046,N_2644);
and UO_166 (O_166,N_2884,N_2230);
and UO_167 (O_167,N_2942,N_2364);
nand UO_168 (O_168,N_2482,N_2113);
nor UO_169 (O_169,N_2763,N_2373);
nand UO_170 (O_170,N_2758,N_2456);
nand UO_171 (O_171,N_2779,N_2332);
or UO_172 (O_172,N_2487,N_2967);
or UO_173 (O_173,N_2858,N_2103);
and UO_174 (O_174,N_2465,N_2678);
nand UO_175 (O_175,N_2707,N_2450);
nand UO_176 (O_176,N_2820,N_2391);
nand UO_177 (O_177,N_2196,N_2605);
and UO_178 (O_178,N_2164,N_2730);
nand UO_179 (O_179,N_2712,N_2953);
nand UO_180 (O_180,N_2019,N_2185);
nor UO_181 (O_181,N_2704,N_2167);
and UO_182 (O_182,N_2777,N_2655);
nor UO_183 (O_183,N_2234,N_2275);
or UO_184 (O_184,N_2769,N_2108);
or UO_185 (O_185,N_2241,N_2166);
and UO_186 (O_186,N_2005,N_2227);
and UO_187 (O_187,N_2709,N_2020);
or UO_188 (O_188,N_2719,N_2314);
nor UO_189 (O_189,N_2440,N_2124);
nor UO_190 (O_190,N_2390,N_2931);
nand UO_191 (O_191,N_2899,N_2256);
or UO_192 (O_192,N_2424,N_2528);
and UO_193 (O_193,N_2483,N_2553);
or UO_194 (O_194,N_2729,N_2859);
and UO_195 (O_195,N_2992,N_2682);
and UO_196 (O_196,N_2409,N_2265);
nor UO_197 (O_197,N_2535,N_2361);
or UO_198 (O_198,N_2030,N_2397);
nand UO_199 (O_199,N_2608,N_2764);
and UO_200 (O_200,N_2088,N_2596);
and UO_201 (O_201,N_2989,N_2505);
and UO_202 (O_202,N_2582,N_2817);
or UO_203 (O_203,N_2921,N_2710);
and UO_204 (O_204,N_2457,N_2470);
or UO_205 (O_205,N_2182,N_2047);
and UO_206 (O_206,N_2065,N_2082);
nand UO_207 (O_207,N_2277,N_2195);
or UO_208 (O_208,N_2952,N_2762);
and UO_209 (O_209,N_2610,N_2159);
nor UO_210 (O_210,N_2353,N_2069);
or UO_211 (O_211,N_2784,N_2190);
and UO_212 (O_212,N_2154,N_2786);
nand UO_213 (O_213,N_2405,N_2803);
nand UO_214 (O_214,N_2215,N_2128);
nand UO_215 (O_215,N_2567,N_2885);
and UO_216 (O_216,N_2865,N_2612);
nor UO_217 (O_217,N_2949,N_2342);
or UO_218 (O_218,N_2853,N_2038);
or UO_219 (O_219,N_2285,N_2431);
and UO_220 (O_220,N_2152,N_2916);
nand UO_221 (O_221,N_2377,N_2372);
and UO_222 (O_222,N_2511,N_2795);
and UO_223 (O_223,N_2430,N_2706);
nand UO_224 (O_224,N_2145,N_2607);
or UO_225 (O_225,N_2757,N_2205);
and UO_226 (O_226,N_2845,N_2756);
nand UO_227 (O_227,N_2073,N_2101);
nand UO_228 (O_228,N_2378,N_2635);
nand UO_229 (O_229,N_2855,N_2111);
nor UO_230 (O_230,N_2814,N_2541);
and UO_231 (O_231,N_2301,N_2399);
nor UO_232 (O_232,N_2991,N_2335);
nor UO_233 (O_233,N_2746,N_2059);
nor UO_234 (O_234,N_2708,N_2693);
and UO_235 (O_235,N_2755,N_2267);
and UO_236 (O_236,N_2997,N_2947);
and UO_237 (O_237,N_2536,N_2276);
nand UO_238 (O_238,N_2174,N_2368);
nor UO_239 (O_239,N_2508,N_2074);
nor UO_240 (O_240,N_2615,N_2352);
nand UO_241 (O_241,N_2210,N_2238);
and UO_242 (O_242,N_2581,N_2261);
and UO_243 (O_243,N_2161,N_2266);
and UO_244 (O_244,N_2414,N_2497);
nor UO_245 (O_245,N_2114,N_2888);
and UO_246 (O_246,N_2681,N_2165);
nor UO_247 (O_247,N_2626,N_2395);
and UO_248 (O_248,N_2398,N_2580);
nor UO_249 (O_249,N_2833,N_2134);
and UO_250 (O_250,N_2319,N_2411);
and UO_251 (O_251,N_2138,N_2913);
nor UO_252 (O_252,N_2739,N_2287);
nor UO_253 (O_253,N_2202,N_2573);
nor UO_254 (O_254,N_2662,N_2736);
nand UO_255 (O_255,N_2687,N_2049);
and UO_256 (O_256,N_2303,N_2840);
or UO_257 (O_257,N_2297,N_2976);
nor UO_258 (O_258,N_2080,N_2703);
or UO_259 (O_259,N_2533,N_2569);
or UO_260 (O_260,N_2009,N_2023);
nor UO_261 (O_261,N_2306,N_2259);
nor UO_262 (O_262,N_2908,N_2805);
nand UO_263 (O_263,N_2349,N_2330);
and UO_264 (O_264,N_2343,N_2296);
and UO_265 (O_265,N_2594,N_2961);
or UO_266 (O_266,N_2337,N_2085);
or UO_267 (O_267,N_2634,N_2999);
or UO_268 (O_268,N_2502,N_2738);
nor UO_269 (O_269,N_2958,N_2042);
nor UO_270 (O_270,N_2625,N_2078);
nor UO_271 (O_271,N_2782,N_2219);
nand UO_272 (O_272,N_2136,N_2591);
or UO_273 (O_273,N_2478,N_2618);
or UO_274 (O_274,N_2289,N_2122);
nand UO_275 (O_275,N_2748,N_2519);
nor UO_276 (O_276,N_2807,N_2156);
nand UO_277 (O_277,N_2910,N_2526);
or UO_278 (O_278,N_2968,N_2013);
nor UO_279 (O_279,N_2956,N_2429);
and UO_280 (O_280,N_2369,N_2280);
and UO_281 (O_281,N_2326,N_2674);
or UO_282 (O_282,N_2812,N_2400);
or UO_283 (O_283,N_2302,N_2523);
or UO_284 (O_284,N_2685,N_2421);
nand UO_285 (O_285,N_2987,N_2371);
nand UO_286 (O_286,N_2919,N_2133);
nor UO_287 (O_287,N_2232,N_2281);
or UO_288 (O_288,N_2753,N_2679);
nand UO_289 (O_289,N_2564,N_2050);
nor UO_290 (O_290,N_2140,N_2220);
and UO_291 (O_291,N_2436,N_2903);
nand UO_292 (O_292,N_2641,N_2521);
or UO_293 (O_293,N_2118,N_2652);
nand UO_294 (O_294,N_2441,N_2866);
and UO_295 (O_295,N_2015,N_2544);
or UO_296 (O_296,N_2012,N_2271);
nand UO_297 (O_297,N_2955,N_2893);
and UO_298 (O_298,N_2351,N_2909);
and UO_299 (O_299,N_2173,N_2771);
or UO_300 (O_300,N_2244,N_2110);
nand UO_301 (O_301,N_2663,N_2291);
or UO_302 (O_302,N_2183,N_2341);
or UO_303 (O_303,N_2100,N_2933);
nor UO_304 (O_304,N_2574,N_2832);
nand UO_305 (O_305,N_2754,N_2447);
or UO_306 (O_306,N_2904,N_2247);
nor UO_307 (O_307,N_2946,N_2245);
or UO_308 (O_308,N_2355,N_2228);
or UO_309 (O_309,N_2328,N_2123);
nand UO_310 (O_310,N_2539,N_2057);
and UO_311 (O_311,N_2270,N_2768);
or UO_312 (O_312,N_2029,N_2559);
and UO_313 (O_313,N_2385,N_2781);
and UO_314 (O_314,N_2158,N_2187);
or UO_315 (O_315,N_2621,N_2623);
nor UO_316 (O_316,N_2906,N_2176);
and UO_317 (O_317,N_2401,N_2308);
and UO_318 (O_318,N_2640,N_2882);
nand UO_319 (O_319,N_2481,N_2937);
or UO_320 (O_320,N_2590,N_2823);
nand UO_321 (O_321,N_2318,N_2690);
and UO_322 (O_322,N_2194,N_2661);
and UO_323 (O_323,N_2721,N_2309);
or UO_324 (O_324,N_2096,N_2305);
nor UO_325 (O_325,N_2630,N_2031);
nand UO_326 (O_326,N_2922,N_2571);
nor UO_327 (O_327,N_2001,N_2650);
nand UO_328 (O_328,N_2294,N_2864);
nand UO_329 (O_329,N_2177,N_2869);
nor UO_330 (O_330,N_2064,N_2233);
nand UO_331 (O_331,N_2062,N_2025);
or UO_332 (O_332,N_2370,N_2413);
nand UO_333 (O_333,N_2599,N_2915);
nand UO_334 (O_334,N_2093,N_2506);
nor UO_335 (O_335,N_2213,N_2792);
xnor UO_336 (O_336,N_2939,N_2467);
nor UO_337 (O_337,N_2877,N_2327);
nor UO_338 (O_338,N_2554,N_2822);
and UO_339 (O_339,N_2199,N_2561);
or UO_340 (O_340,N_2629,N_2021);
nor UO_341 (O_341,N_2588,N_2189);
or UO_342 (O_342,N_2090,N_2609);
xnor UO_343 (O_343,N_2996,N_2403);
and UO_344 (O_344,N_2448,N_2943);
or UO_345 (O_345,N_2251,N_2444);
and UO_346 (O_346,N_2249,N_2486);
nor UO_347 (O_347,N_2054,N_2198);
nor UO_348 (O_348,N_2178,N_2818);
nand UO_349 (O_349,N_2148,N_2857);
nand UO_350 (O_350,N_2643,N_2878);
nor UO_351 (O_351,N_2524,N_2861);
or UO_352 (O_352,N_2356,N_2004);
or UO_353 (O_353,N_2834,N_2426);
and UO_354 (O_354,N_2469,N_2810);
or UO_355 (O_355,N_2499,N_2598);
and UO_356 (O_356,N_2484,N_2751);
nand UO_357 (O_357,N_2551,N_2142);
or UO_358 (O_358,N_2146,N_2056);
nor UO_359 (O_359,N_2387,N_2000);
or UO_360 (O_360,N_2852,N_2636);
or UO_361 (O_361,N_2586,N_2993);
and UO_362 (O_362,N_2940,N_2036);
or UO_363 (O_363,N_2659,N_2451);
and UO_364 (O_364,N_2868,N_2694);
and UO_365 (O_365,N_2423,N_2221);
and UO_366 (O_366,N_2357,N_2462);
or UO_367 (O_367,N_2718,N_2510);
nand UO_368 (O_368,N_2006,N_2638);
or UO_369 (O_369,N_2887,N_2155);
nand UO_370 (O_370,N_2839,N_2604);
nor UO_371 (O_371,N_2500,N_2388);
nor UO_372 (O_372,N_2135,N_2039);
or UO_373 (O_373,N_2836,N_2616);
or UO_374 (O_374,N_2622,N_2446);
and UO_375 (O_375,N_2316,N_2034);
and UO_376 (O_376,N_2255,N_2816);
nor UO_377 (O_377,N_2162,N_2077);
nor UO_378 (O_378,N_2901,N_2522);
nor UO_379 (O_379,N_2978,N_2724);
nor UO_380 (O_380,N_2105,N_2143);
or UO_381 (O_381,N_2017,N_2292);
nor UO_382 (O_382,N_2045,N_2593);
or UO_383 (O_383,N_2149,N_2585);
and UO_384 (O_384,N_2002,N_2780);
or UO_385 (O_385,N_2461,N_2880);
or UO_386 (O_386,N_2504,N_2930);
nand UO_387 (O_387,N_2716,N_2498);
or UO_388 (O_388,N_2863,N_2003);
or UO_389 (O_389,N_2396,N_2619);
nor UO_390 (O_390,N_2686,N_2851);
and UO_391 (O_391,N_2035,N_2317);
or UO_392 (O_392,N_2672,N_2971);
and UO_393 (O_393,N_2660,N_2374);
nor UO_394 (O_394,N_2813,N_2701);
or UO_395 (O_395,N_2420,N_2966);
or UO_396 (O_396,N_2350,N_2990);
nor UO_397 (O_397,N_2881,N_2336);
and UO_398 (O_398,N_2867,N_2669);
nand UO_399 (O_399,N_2095,N_2787);
or UO_400 (O_400,N_2315,N_2734);
nor UO_401 (O_401,N_2849,N_2965);
nor UO_402 (O_402,N_2331,N_2218);
nor UO_403 (O_403,N_2547,N_2545);
or UO_404 (O_404,N_2565,N_2743);
and UO_405 (O_405,N_2007,N_2117);
nor UO_406 (O_406,N_2714,N_2175);
nand UO_407 (O_407,N_2439,N_2558);
nor UO_408 (O_408,N_2112,N_2676);
and UO_409 (O_409,N_2827,N_2473);
nor UO_410 (O_410,N_2094,N_2127);
and UO_411 (O_411,N_2365,N_2741);
nand UO_412 (O_412,N_2772,N_2589);
nand UO_413 (O_413,N_2912,N_2452);
and UO_414 (O_414,N_2010,N_2053);
or UO_415 (O_415,N_2282,N_2938);
nand UO_416 (O_416,N_2273,N_2091);
nand UO_417 (O_417,N_2572,N_2725);
or UO_418 (O_418,N_2243,N_2491);
and UO_419 (O_419,N_2854,N_2720);
nor UO_420 (O_420,N_2311,N_2698);
nand UO_421 (O_421,N_2340,N_2555);
nor UO_422 (O_422,N_2732,N_2587);
nand UO_423 (O_423,N_2886,N_2617);
nand UO_424 (O_424,N_2670,N_2477);
nand UO_425 (O_425,N_2099,N_2027);
nand UO_426 (O_426,N_2560,N_2055);
nand UO_427 (O_427,N_2492,N_2323);
nand UO_428 (O_428,N_2226,N_2229);
or UO_429 (O_429,N_2207,N_2120);
nand UO_430 (O_430,N_2918,N_2347);
nand UO_431 (O_431,N_2339,N_2691);
nor UO_432 (O_432,N_2801,N_2092);
nand UO_433 (O_433,N_2945,N_2417);
and UO_434 (O_434,N_2552,N_2263);
and UO_435 (O_435,N_2928,N_2367);
nand UO_436 (O_436,N_2380,N_2197);
nand UO_437 (O_437,N_2983,N_2236);
nand UO_438 (O_438,N_2237,N_2304);
nand UO_439 (O_439,N_2633,N_2826);
nor UO_440 (O_440,N_2819,N_2575);
or UO_441 (O_441,N_2141,N_2985);
or UO_442 (O_442,N_2944,N_2657);
and UO_443 (O_443,N_2929,N_2333);
and UO_444 (O_444,N_2518,N_2248);
nor UO_445 (O_445,N_2354,N_2711);
and UO_446 (O_446,N_2453,N_2445);
nand UO_447 (O_447,N_2517,N_2125);
or UO_448 (O_448,N_2684,N_2438);
or UO_449 (O_449,N_2300,N_2386);
nor UO_450 (O_450,N_2375,N_2637);
nor UO_451 (O_451,N_2972,N_2404);
and UO_452 (O_452,N_2802,N_2897);
and UO_453 (O_453,N_2982,N_2986);
nand UO_454 (O_454,N_2717,N_2460);
or UO_455 (O_455,N_2773,N_2549);
or UO_456 (O_456,N_2873,N_2201);
or UO_457 (O_457,N_2744,N_2171);
nand UO_458 (O_458,N_2115,N_2752);
nand UO_459 (O_459,N_2742,N_2131);
nand UO_460 (O_460,N_2086,N_2715);
nand UO_461 (O_461,N_2322,N_2761);
nor UO_462 (O_462,N_2513,N_2379);
nor UO_463 (O_463,N_2994,N_2838);
nor UO_464 (O_464,N_2821,N_2658);
nand UO_465 (O_465,N_2702,N_2132);
nand UO_466 (O_466,N_2109,N_2828);
nor UO_467 (O_467,N_2532,N_2032);
nor UO_468 (O_468,N_2829,N_2830);
or UO_469 (O_469,N_2995,N_2160);
nor UO_470 (O_470,N_2791,N_2151);
nand UO_471 (O_471,N_2425,N_2509);
nand UO_472 (O_472,N_2653,N_2948);
and UO_473 (O_473,N_2578,N_2546);
nand UO_474 (O_474,N_2321,N_2979);
or UO_475 (O_475,N_2778,N_2217);
nor UO_476 (O_476,N_2841,N_2225);
and UO_477 (O_477,N_2896,N_2525);
or UO_478 (O_478,N_2348,N_2214);
or UO_479 (O_479,N_2680,N_2434);
nand UO_480 (O_480,N_2647,N_2410);
nor UO_481 (O_481,N_2871,N_2345);
nor UO_482 (O_482,N_2570,N_2924);
nand UO_483 (O_483,N_2529,N_2200);
and UO_484 (O_484,N_2168,N_2163);
or UO_485 (O_485,N_2848,N_2872);
nor UO_486 (O_486,N_2584,N_2268);
nand UO_487 (O_487,N_2749,N_2592);
nor UO_488 (O_488,N_2312,N_2925);
nor UO_489 (O_489,N_2557,N_2324);
nor UO_490 (O_490,N_2383,N_2058);
nand UO_491 (O_491,N_2601,N_2188);
nand UO_492 (O_492,N_2666,N_2419);
and UO_493 (O_493,N_2775,N_2070);
or UO_494 (O_494,N_2750,N_2051);
nor UO_495 (O_495,N_2892,N_2797);
or UO_496 (O_496,N_2760,N_2416);
or UO_497 (O_497,N_2104,N_2264);
or UO_498 (O_498,N_2843,N_2731);
nor UO_499 (O_499,N_2579,N_2926);
endmodule