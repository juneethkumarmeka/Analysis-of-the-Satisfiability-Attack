module basic_2000_20000_2500_80_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1055,In_1174);
or U1 (N_1,In_159,In_1863);
nor U2 (N_2,In_19,In_1360);
nand U3 (N_3,In_1592,In_1214);
or U4 (N_4,In_1416,In_1057);
or U5 (N_5,In_162,In_1618);
nand U6 (N_6,In_864,In_634);
or U7 (N_7,In_703,In_8);
nor U8 (N_8,In_1676,In_1304);
and U9 (N_9,In_1436,In_322);
nand U10 (N_10,In_466,In_130);
nand U11 (N_11,In_366,In_356);
nor U12 (N_12,In_488,In_1797);
nand U13 (N_13,In_52,In_494);
xor U14 (N_14,In_370,In_541);
or U15 (N_15,In_1384,In_1501);
nand U16 (N_16,In_1855,In_616);
xnor U17 (N_17,In_1959,In_1255);
nand U18 (N_18,In_502,In_436);
and U19 (N_19,In_486,In_1173);
nand U20 (N_20,In_1429,In_1804);
nand U21 (N_21,In_1956,In_1833);
nand U22 (N_22,In_1886,In_1207);
nand U23 (N_23,In_1748,In_45);
xor U24 (N_24,In_1058,In_1373);
nor U25 (N_25,In_1049,In_630);
and U26 (N_26,In_181,In_1218);
nor U27 (N_27,In_1003,In_1466);
nor U28 (N_28,In_365,In_463);
nor U29 (N_29,In_107,In_372);
nor U30 (N_30,In_913,In_249);
and U31 (N_31,In_982,In_1896);
nor U32 (N_32,In_1019,In_134);
nand U33 (N_33,In_414,In_1341);
and U34 (N_34,In_470,In_718);
and U35 (N_35,In_830,In_32);
nor U36 (N_36,In_1795,In_1302);
xnor U37 (N_37,In_343,In_270);
and U38 (N_38,In_1723,In_195);
nand U39 (N_39,In_554,In_1564);
xnor U40 (N_40,In_1093,In_1550);
nand U41 (N_41,In_581,In_203);
or U42 (N_42,In_1254,In_688);
nor U43 (N_43,In_1771,In_1839);
and U44 (N_44,In_1940,In_1531);
or U45 (N_45,In_699,In_1705);
and U46 (N_46,In_686,In_1699);
nor U47 (N_47,In_1256,In_1890);
and U48 (N_48,In_1397,In_230);
or U49 (N_49,In_14,In_1636);
nand U50 (N_50,In_1925,In_1335);
and U51 (N_51,In_487,In_1900);
nor U52 (N_52,In_1388,In_192);
nand U53 (N_53,In_260,In_919);
or U54 (N_54,In_1758,In_399);
xor U55 (N_55,In_754,In_1004);
nor U56 (N_56,In_313,In_735);
xnor U57 (N_57,In_144,In_835);
and U58 (N_58,In_814,In_1829);
nor U59 (N_59,In_758,In_872);
nand U60 (N_60,In_323,In_1065);
or U61 (N_61,In_821,In_1024);
and U62 (N_62,In_390,In_823);
xor U63 (N_63,In_1337,In_362);
and U64 (N_64,In_388,In_1349);
and U65 (N_65,In_64,In_431);
or U66 (N_66,In_1917,In_1314);
nor U67 (N_67,In_160,In_956);
or U68 (N_68,In_1502,In_1759);
and U69 (N_69,In_600,In_1442);
and U70 (N_70,In_566,In_1725);
nand U71 (N_71,In_248,In_796);
nor U72 (N_72,In_1224,In_100);
nand U73 (N_73,In_1523,In_1062);
xor U74 (N_74,In_1901,In_866);
xnor U75 (N_75,In_1334,In_1104);
xor U76 (N_76,In_1646,In_695);
or U77 (N_77,In_206,In_655);
nor U78 (N_78,In_1897,In_946);
or U79 (N_79,In_559,In_1274);
and U80 (N_80,In_1285,In_257);
xnor U81 (N_81,In_1366,In_951);
nor U82 (N_82,In_1082,In_1033);
nor U83 (N_83,In_674,In_288);
nor U84 (N_84,In_21,In_1496);
or U85 (N_85,In_1432,In_646);
and U86 (N_86,In_826,In_139);
nand U87 (N_87,In_1427,In_1456);
and U88 (N_88,In_250,In_408);
and U89 (N_89,In_20,In_818);
nor U90 (N_90,In_430,In_1541);
or U91 (N_91,In_1162,In_1657);
and U92 (N_92,In_1772,In_1097);
xor U93 (N_93,In_543,In_743);
nand U94 (N_94,In_596,In_1631);
nor U95 (N_95,In_1014,In_305);
nand U96 (N_96,In_276,In_1383);
nand U97 (N_97,In_1094,In_1847);
nor U98 (N_98,In_1719,In_207);
and U99 (N_99,In_193,In_1567);
and U100 (N_100,In_1278,In_560);
nand U101 (N_101,In_1754,In_642);
nand U102 (N_102,In_663,In_1372);
and U103 (N_103,In_772,In_1023);
and U104 (N_104,In_1348,In_1529);
and U105 (N_105,In_1601,In_1327);
or U106 (N_106,In_778,In_673);
xor U107 (N_107,In_259,In_464);
and U108 (N_108,In_698,In_43);
and U109 (N_109,In_369,In_1777);
or U110 (N_110,In_660,In_1559);
or U111 (N_111,In_1110,In_1343);
xor U112 (N_112,In_1967,In_1975);
nor U113 (N_113,In_836,In_434);
nand U114 (N_114,In_1259,In_535);
or U115 (N_115,In_636,In_1151);
nand U116 (N_116,In_593,In_500);
or U117 (N_117,In_832,In_941);
nor U118 (N_118,In_786,In_125);
xnor U119 (N_119,In_1208,In_802);
or U120 (N_120,In_1281,In_1707);
or U121 (N_121,In_1694,In_961);
nor U122 (N_122,In_338,In_256);
nor U123 (N_123,In_167,In_1491);
xor U124 (N_124,In_1415,In_1430);
nor U125 (N_125,In_316,In_1328);
or U126 (N_126,In_1017,In_861);
nor U127 (N_127,In_580,In_839);
xor U128 (N_128,In_635,In_173);
nor U129 (N_129,In_1088,In_1858);
xnor U130 (N_130,In_1930,In_1325);
nand U131 (N_131,In_1691,In_1935);
xor U132 (N_132,In_1828,In_391);
nand U133 (N_133,In_1671,In_321);
or U134 (N_134,In_1981,In_710);
nor U135 (N_135,In_480,In_1878);
nor U136 (N_136,In_817,In_613);
nor U137 (N_137,In_1681,In_185);
nor U138 (N_138,In_1464,In_1363);
nor U139 (N_139,In_1655,In_1459);
xor U140 (N_140,In_1751,In_479);
nand U141 (N_141,In_1879,In_1887);
nor U142 (N_142,In_6,In_459);
nor U143 (N_143,In_1120,In_765);
nor U144 (N_144,In_263,In_751);
and U145 (N_145,In_307,In_849);
or U146 (N_146,In_1376,In_1428);
and U147 (N_147,In_649,In_1472);
or U148 (N_148,In_297,In_1536);
xor U149 (N_149,In_671,In_1245);
xnor U150 (N_150,In_484,In_1808);
nand U151 (N_151,In_1525,In_1244);
and U152 (N_152,In_1022,In_1742);
xnor U153 (N_153,In_1010,In_1047);
nand U154 (N_154,In_429,In_73);
nand U155 (N_155,In_1864,In_86);
and U156 (N_156,In_917,In_217);
nor U157 (N_157,In_172,In_892);
xor U158 (N_158,In_867,In_925);
xor U159 (N_159,In_647,In_211);
or U160 (N_160,In_342,In_1730);
nor U161 (N_161,In_199,In_843);
nor U162 (N_162,In_933,In_1101);
and U163 (N_163,In_1267,In_318);
nand U164 (N_164,In_178,In_1217);
xnor U165 (N_165,In_1139,In_1535);
or U166 (N_166,In_1385,In_1982);
xor U167 (N_167,In_563,In_813);
nand U168 (N_168,In_1508,In_1998);
and U169 (N_169,In_294,In_1654);
nand U170 (N_170,In_1986,In_1412);
nand U171 (N_171,In_883,In_1626);
and U172 (N_172,In_103,In_1928);
xor U173 (N_173,In_1507,In_539);
or U174 (N_174,In_1303,In_1371);
and U175 (N_175,In_672,In_964);
nand U176 (N_176,In_1206,In_1187);
and U177 (N_177,In_1695,In_221);
nor U178 (N_178,In_1499,In_1205);
and U179 (N_179,In_55,In_1013);
nand U180 (N_180,In_869,In_963);
nand U181 (N_181,In_675,In_1046);
or U182 (N_182,In_1961,In_168);
nand U183 (N_183,In_567,In_1942);
nor U184 (N_184,In_1331,In_265);
nor U185 (N_185,In_93,In_22);
or U186 (N_186,In_1934,In_1816);
or U187 (N_187,In_1148,In_1953);
or U188 (N_188,In_1391,In_87);
or U189 (N_189,In_651,In_90);
nand U190 (N_190,In_174,In_656);
or U191 (N_191,In_1015,In_54);
nor U192 (N_192,In_1423,In_451);
nand U193 (N_193,In_555,In_1565);
xor U194 (N_194,In_368,In_677);
nand U195 (N_195,In_186,In_573);
xor U196 (N_196,In_1765,In_1779);
xor U197 (N_197,In_627,In_213);
xor U198 (N_198,In_1786,In_1685);
xor U199 (N_199,In_1638,In_266);
xor U200 (N_200,In_105,In_1913);
and U201 (N_201,In_1538,In_1850);
or U202 (N_202,In_310,In_364);
xnor U203 (N_203,In_960,In_202);
or U204 (N_204,In_1936,In_7);
or U205 (N_205,In_1545,In_1770);
xnor U206 (N_206,In_1239,In_1673);
nand U207 (N_207,In_1875,In_141);
or U208 (N_208,In_709,In_377);
or U209 (N_209,In_472,In_662);
or U210 (N_210,In_1071,In_1556);
nor U211 (N_211,In_165,In_524);
or U212 (N_212,In_1895,In_47);
nor U213 (N_213,In_1111,In_1223);
nand U214 (N_214,In_1659,In_352);
xor U215 (N_215,In_379,In_1486);
nor U216 (N_216,In_1340,In_1095);
nor U217 (N_217,In_1380,In_687);
xnor U218 (N_218,In_16,In_1465);
nor U219 (N_219,In_788,In_943);
nand U220 (N_220,In_1179,In_285);
nor U221 (N_221,In_768,In_1006);
nor U222 (N_222,In_389,In_950);
xnor U223 (N_223,In_58,In_572);
nor U224 (N_224,In_551,In_1774);
nor U225 (N_225,In_278,In_1649);
or U226 (N_226,In_1190,In_1729);
or U227 (N_227,In_66,In_239);
or U228 (N_228,In_387,In_1396);
or U229 (N_229,In_1471,In_80);
nor U230 (N_230,In_465,In_79);
nor U231 (N_231,In_1883,In_1778);
nand U232 (N_232,In_781,In_155);
xnor U233 (N_233,In_309,In_658);
or U234 (N_234,In_719,In_1438);
and U235 (N_235,In_244,In_1718);
xor U236 (N_236,In_77,In_1361);
nand U237 (N_237,In_1399,In_750);
or U238 (N_238,In_1229,In_1509);
xnor U239 (N_239,In_1540,In_1996);
nor U240 (N_240,In_1775,In_1113);
nor U241 (N_241,In_1030,In_1249);
xor U242 (N_242,In_371,In_226);
nand U243 (N_243,In_180,In_808);
nand U244 (N_244,In_1216,In_582);
nand U245 (N_245,In_1378,In_1698);
nor U246 (N_246,In_1419,In_910);
nor U247 (N_247,In_1087,In_979);
and U248 (N_248,In_438,In_863);
and U249 (N_249,In_1112,In_791);
and U250 (N_250,In_908,In_1075);
and U251 (N_251,In_1460,In_540);
xnor U252 (N_252,In_200,In_190);
nor U253 (N_253,In_1530,In_1859);
xor U254 (N_254,In_1791,In_1822);
nand U255 (N_255,N_16,In_95);
xnor U256 (N_256,N_218,In_1821);
nand U257 (N_257,N_196,In_948);
nand U258 (N_258,In_421,In_1226);
or U259 (N_259,In_1286,In_509);
nor U260 (N_260,In_1276,In_746);
nor U261 (N_261,In_763,In_1131);
nand U262 (N_262,In_744,In_1150);
and U263 (N_263,In_1234,In_1992);
nand U264 (N_264,In_238,N_160);
or U265 (N_265,N_221,N_51);
and U266 (N_266,In_1773,In_766);
nand U267 (N_267,In_1827,In_886);
nand U268 (N_268,In_1362,In_1853);
nand U269 (N_269,In_974,In_271);
and U270 (N_270,N_68,N_25);
nor U271 (N_271,In_331,In_998);
xnor U272 (N_272,In_34,In_696);
xnor U273 (N_273,In_548,In_1248);
and U274 (N_274,In_975,In_179);
nand U275 (N_275,N_127,In_1843);
xnor U276 (N_276,N_34,In_59);
xor U277 (N_277,N_120,In_1811);
or U278 (N_278,In_624,In_106);
xnor U279 (N_279,In_603,In_1678);
or U280 (N_280,In_1801,N_248);
nand U281 (N_281,In_1583,In_1924);
or U282 (N_282,In_1102,In_967);
nor U283 (N_283,In_1393,In_1869);
nor U284 (N_284,In_247,In_792);
or U285 (N_285,In_1861,In_684);
nand U286 (N_286,In_231,In_531);
xor U287 (N_287,In_1163,N_147);
or U288 (N_288,In_1236,In_644);
or U289 (N_289,In_939,In_1785);
nand U290 (N_290,N_4,In_1194);
and U291 (N_291,In_1090,In_169);
nand U292 (N_292,In_1974,In_1577);
nor U293 (N_293,In_461,In_1116);
and U294 (N_294,In_1289,In_1143);
or U295 (N_295,In_456,In_855);
nor U296 (N_296,In_771,N_159);
or U297 (N_297,N_152,In_556);
nand U298 (N_298,N_99,N_222);
or U299 (N_299,In_1240,In_1849);
xor U300 (N_300,In_373,In_78);
xor U301 (N_301,In_26,In_1985);
nor U302 (N_302,In_1100,In_1727);
nand U303 (N_303,In_668,N_41);
nand U304 (N_304,In_191,N_190);
nand U305 (N_305,In_282,In_150);
or U306 (N_306,In_659,In_1658);
xor U307 (N_307,N_246,In_787);
nor U308 (N_308,In_110,In_320);
and U309 (N_309,N_140,N_178);
and U310 (N_310,In_1487,In_170);
nand U311 (N_311,In_293,In_76);
nand U312 (N_312,N_189,In_355);
nand U313 (N_313,In_853,In_1783);
or U314 (N_314,In_251,In_1734);
nand U315 (N_315,In_1221,In_1937);
or U316 (N_316,In_208,In_1941);
nor U317 (N_317,N_239,In_592);
nor U318 (N_318,In_586,In_392);
nand U319 (N_319,In_1511,In_631);
xnor U320 (N_320,In_1333,In_605);
nor U321 (N_321,In_1546,In_732);
nand U322 (N_322,In_850,N_36);
nor U323 (N_323,In_1637,In_986);
xnor U324 (N_324,In_1746,N_92);
or U325 (N_325,In_733,In_354);
or U326 (N_326,In_1025,In_1520);
and U327 (N_327,In_1454,In_234);
xor U328 (N_328,In_183,N_94);
nand U329 (N_329,In_1135,In_638);
nand U330 (N_330,In_949,In_728);
and U331 (N_331,In_1933,In_520);
xor U332 (N_332,In_1191,N_45);
xor U333 (N_333,In_1524,In_491);
xor U334 (N_334,In_799,In_1129);
nand U335 (N_335,N_230,In_922);
or U336 (N_336,In_1997,In_1145);
nand U337 (N_337,In_1026,In_1856);
nor U338 (N_338,In_82,N_185);
xnor U339 (N_339,In_1085,In_1845);
xor U340 (N_340,N_176,In_1475);
xor U341 (N_341,In_1892,In_17);
and U342 (N_342,In_1860,In_443);
nand U343 (N_343,In_610,In_1332);
and U344 (N_344,In_1449,In_1506);
xnor U345 (N_345,In_811,In_1377);
xor U346 (N_346,In_755,N_146);
nand U347 (N_347,In_447,In_1769);
nor U348 (N_348,N_137,In_1282);
nor U349 (N_349,In_209,In_1212);
and U350 (N_350,In_166,In_117);
nand U351 (N_351,N_219,In_385);
xor U352 (N_352,In_1086,In_1387);
and U353 (N_353,In_738,N_180);
xor U354 (N_354,In_1405,In_514);
and U355 (N_355,In_403,In_724);
or U356 (N_356,In_928,N_47);
nor U357 (N_357,In_901,In_415);
or U358 (N_358,In_62,In_1735);
xnor U359 (N_359,In_876,In_1979);
nand U360 (N_360,N_149,In_1105);
xor U361 (N_361,N_24,N_102);
or U362 (N_362,In_1789,In_904);
and U363 (N_363,In_1622,In_992);
nand U364 (N_364,In_909,N_174);
or U365 (N_365,In_1932,In_1096);
and U366 (N_366,In_444,N_208);
nand U367 (N_367,N_203,In_1064);
and U368 (N_368,In_595,In_707);
nand U369 (N_369,N_156,In_1570);
nor U370 (N_370,N_214,In_923);
nand U371 (N_371,In_1692,In_882);
and U372 (N_372,In_1166,In_1009);
nand U373 (N_373,In_1539,In_701);
and U374 (N_374,In_784,In_1243);
nor U375 (N_375,In_13,In_324);
nor U376 (N_376,In_261,N_101);
and U377 (N_377,In_116,In_1213);
or U378 (N_378,In_1784,In_433);
nor U379 (N_379,N_145,In_1688);
or U380 (N_380,In_1841,In_332);
xnor U381 (N_381,In_1357,In_1787);
or U382 (N_382,In_553,N_5);
and U383 (N_383,In_1137,In_1666);
nor U384 (N_384,N_193,In_918);
xor U385 (N_385,N_188,In_2);
or U386 (N_386,In_1027,In_905);
or U387 (N_387,N_43,In_1198);
nand U388 (N_388,In_1273,In_1505);
xnor U389 (N_389,In_1620,In_1478);
or U390 (N_390,In_1835,In_907);
or U391 (N_391,In_1242,In_1481);
nor U392 (N_392,In_666,In_1593);
nand U393 (N_393,In_584,In_476);
and U394 (N_394,In_1750,In_1018);
or U395 (N_395,N_199,In_1128);
or U396 (N_396,In_550,In_529);
nor U397 (N_397,N_134,N_56);
or U398 (N_398,In_1687,In_280);
and U399 (N_399,In_669,In_1199);
and U400 (N_400,In_590,In_895);
and U401 (N_401,In_1722,N_210);
nor U402 (N_402,N_155,In_1984);
xor U403 (N_403,In_122,In_968);
nor U404 (N_404,In_827,In_1885);
or U405 (N_405,In_384,In_1756);
nand U406 (N_406,In_145,In_824);
or U407 (N_407,In_1960,In_1837);
or U408 (N_408,In_594,In_657);
nor U409 (N_409,In_304,N_108);
and U410 (N_410,In_518,In_1519);
nor U411 (N_411,In_1921,In_712);
or U412 (N_412,In_1051,N_168);
and U413 (N_413,In_154,In_1706);
or U414 (N_414,In_1528,In_612);
xor U415 (N_415,In_1070,N_226);
or U416 (N_416,In_1445,In_637);
nand U417 (N_417,N_163,In_1211);
xnor U418 (N_418,N_77,N_247);
and U419 (N_419,In_1990,In_361);
and U420 (N_420,N_172,In_452);
or U421 (N_421,In_1156,In_1983);
and U422 (N_422,In_532,In_622);
nor U423 (N_423,In_1020,In_809);
or U424 (N_424,In_1374,In_874);
nor U425 (N_425,In_1728,In_748);
nand U426 (N_426,In_1227,In_398);
nor U427 (N_427,In_1854,In_133);
xor U428 (N_428,In_253,In_120);
and U429 (N_429,In_557,In_1966);
nor U430 (N_430,In_683,In_295);
nand U431 (N_431,In_916,In_1168);
or U432 (N_432,In_1625,In_665);
nor U433 (N_433,In_1521,N_38);
nor U434 (N_434,In_457,In_736);
nor U435 (N_435,In_993,N_202);
nor U436 (N_436,In_1186,In_511);
and U437 (N_437,In_935,In_1246);
nor U438 (N_438,N_13,In_926);
and U439 (N_439,In_608,In_1401);
nor U440 (N_440,In_1381,In_505);
nand U441 (N_441,In_1693,In_136);
or U442 (N_442,In_525,In_471);
and U443 (N_443,N_216,In_1209);
or U444 (N_444,In_109,In_153);
or U445 (N_445,In_989,In_1183);
xor U446 (N_446,In_482,N_33);
nor U447 (N_447,In_1080,In_1595);
xnor U448 (N_448,In_1629,In_1617);
or U449 (N_449,In_1250,In_1158);
or U450 (N_450,In_1846,In_1339);
or U451 (N_451,In_1392,In_123);
or U452 (N_452,In_84,In_860);
and U453 (N_453,In_450,In_1379);
or U454 (N_454,In_845,In_1884);
nand U455 (N_455,In_1737,In_1414);
or U456 (N_456,In_891,In_1597);
or U457 (N_457,In_252,In_819);
nor U458 (N_458,In_279,In_652);
xor U459 (N_459,N_100,In_129);
and U460 (N_460,In_501,In_576);
nor U461 (N_461,In_498,N_138);
nor U462 (N_462,In_1441,In_1196);
or U463 (N_463,In_477,In_1140);
nand U464 (N_464,In_448,In_1317);
or U465 (N_465,In_1572,In_1547);
nand U466 (N_466,In_1098,In_715);
or U467 (N_467,In_1232,N_8);
and U468 (N_468,In_1338,In_1680);
nand U469 (N_469,In_1912,In_602);
and U470 (N_470,In_1117,In_752);
xnor U471 (N_471,In_1910,In_1606);
xor U472 (N_472,In_411,In_737);
or U473 (N_473,In_854,In_1455);
nor U474 (N_474,In_1514,In_625);
nor U475 (N_475,In_797,In_947);
xnor U476 (N_476,In_235,In_633);
or U477 (N_477,N_75,In_921);
and U478 (N_478,In_1566,N_76);
nor U479 (N_479,N_3,In_300);
nand U480 (N_480,In_126,N_238);
xor U481 (N_481,In_46,In_1418);
and U482 (N_482,N_231,N_37);
and U483 (N_483,In_1668,In_749);
and U484 (N_484,In_1813,In_1193);
nand U485 (N_485,In_75,In_629);
or U486 (N_486,In_404,In_700);
and U487 (N_487,In_287,N_175);
and U488 (N_488,In_0,In_831);
nand U489 (N_489,In_920,In_1409);
and U490 (N_490,In_1220,N_93);
xor U491 (N_491,In_938,In_131);
xor U492 (N_492,In_1563,In_1149);
xor U493 (N_493,In_396,In_242);
nor U494 (N_494,N_20,In_577);
nor U495 (N_495,In_135,In_311);
or U496 (N_496,In_1720,In_1359);
xnor U497 (N_497,In_71,In_1130);
xor U498 (N_498,In_1905,In_506);
nand U499 (N_499,N_192,In_1309);
or U500 (N_500,In_1307,N_410);
and U501 (N_501,N_474,N_467);
or U502 (N_502,In_38,In_611);
xnor U503 (N_503,In_680,In_1477);
nor U504 (N_504,In_1633,In_1311);
nor U505 (N_505,N_30,N_370);
or U506 (N_506,In_375,In_1607);
or U507 (N_507,N_267,In_1534);
xor U508 (N_508,In_94,In_1504);
or U509 (N_509,N_142,In_924);
or U510 (N_510,N_454,In_1315);
xnor U511 (N_511,In_1950,In_290);
nor U512 (N_512,N_245,In_690);
or U513 (N_513,In_83,In_522);
xor U514 (N_514,In_382,N_7);
nand U515 (N_515,In_1488,In_1053);
or U516 (N_516,In_1042,In_359);
nor U517 (N_517,In_243,In_1865);
nor U518 (N_518,N_404,In_1346);
nand U519 (N_519,In_1195,In_315);
nor U520 (N_520,In_1189,N_407);
nand U521 (N_521,In_694,N_366);
or U522 (N_522,In_575,In_934);
nor U523 (N_523,In_1741,In_1252);
xnor U524 (N_524,N_337,In_1988);
xor U525 (N_525,N_364,In_156);
and U526 (N_526,In_1484,In_847);
nand U527 (N_527,N_487,N_493);
and U528 (N_528,N_169,In_984);
and U529 (N_529,In_1964,In_1696);
nor U530 (N_530,In_1284,N_330);
and U531 (N_531,In_1980,In_1123);
nor U532 (N_532,N_243,N_396);
and U533 (N_533,In_1115,In_969);
xor U534 (N_534,In_1969,In_91);
nand U535 (N_535,In_25,In_1144);
xor U536 (N_536,In_1512,In_148);
nand U537 (N_537,In_468,In_1736);
nand U538 (N_538,In_360,N_342);
nand U539 (N_539,In_1308,In_1201);
nand U540 (N_540,In_1175,In_41);
and U541 (N_541,In_317,In_1731);
nand U542 (N_542,N_184,In_115);
nand U543 (N_543,In_1968,N_420);
nor U544 (N_544,In_419,N_384);
nor U545 (N_545,N_328,N_340);
nor U546 (N_546,N_472,N_74);
or U547 (N_547,In_1612,N_441);
nor U548 (N_548,In_1448,N_260);
nand U549 (N_549,In_262,In_1877);
and U550 (N_550,In_1747,In_1493);
nand U551 (N_551,N_411,In_1641);
xor U552 (N_552,In_1326,In_264);
and U553 (N_553,In_1323,In_957);
xor U554 (N_554,In_113,In_1739);
xor U555 (N_555,In_704,In_1410);
xor U556 (N_556,N_48,N_57);
or U557 (N_557,N_71,In_132);
xor U558 (N_558,In_897,In_1165);
xor U559 (N_559,In_676,In_48);
nor U560 (N_560,In_473,N_447);
or U561 (N_561,In_1672,N_171);
nor U562 (N_562,In_1836,N_59);
nor U563 (N_563,In_1796,In_760);
or U564 (N_564,In_163,In_1918);
xor U565 (N_565,In_1132,In_1642);
nand U566 (N_566,In_161,In_729);
nor U567 (N_567,In_1630,N_347);
nor U568 (N_568,N_314,In_534);
nand U569 (N_569,In_1495,In_36);
or U570 (N_570,In_1184,In_776);
nor U571 (N_571,In_1876,In_723);
nand U572 (N_572,In_806,In_1761);
and U573 (N_573,In_1639,In_1803);
nor U574 (N_574,In_670,In_536);
nand U575 (N_575,In_401,In_296);
and U576 (N_576,N_424,In_1350);
nand U577 (N_577,In_1032,N_227);
nand U578 (N_578,In_1463,In_1159);
nand U579 (N_579,In_1265,In_713);
nor U580 (N_580,In_1899,In_1825);
or U581 (N_581,In_1920,In_1169);
nand U582 (N_582,N_444,N_109);
nor U583 (N_583,N_97,N_166);
and U584 (N_584,In_1743,In_1697);
xnor U585 (N_585,In_1922,N_50);
and U586 (N_586,In_1907,In_196);
nand U587 (N_587,In_281,In_834);
nand U588 (N_588,In_1702,In_1439);
or U589 (N_589,In_1893,N_325);
nand U590 (N_590,N_321,In_1627);
nand U591 (N_591,N_381,N_73);
and U592 (N_592,In_965,In_1498);
or U593 (N_593,In_1684,In_1081);
xnor U594 (N_594,In_1167,In_1955);
and U595 (N_595,In_777,In_1407);
nand U596 (N_596,In_1682,In_329);
and U597 (N_597,In_708,N_439);
and U598 (N_598,In_337,In_1868);
and U599 (N_599,In_1660,N_430);
nand U600 (N_600,In_994,In_678);
or U601 (N_601,N_177,In_1319);
or U602 (N_602,In_1790,In_903);
xnor U603 (N_603,N_377,In_1903);
and U604 (N_604,In_734,In_842);
nand U605 (N_605,In_664,In_1440);
xor U606 (N_606,N_343,In_1548);
xnor U607 (N_607,In_1798,N_78);
nor U608 (N_608,In_1526,N_287);
nor U609 (N_609,In_731,N_82);
nor U610 (N_610,In_412,In_619);
nor U611 (N_611,In_1870,N_452);
nand U612 (N_612,N_312,In_496);
nand U613 (N_613,In_1532,In_640);
xnor U614 (N_614,N_479,N_197);
nor U615 (N_615,In_1453,N_409);
xnor U616 (N_616,In_23,In_1600);
or U617 (N_617,In_140,In_1831);
nand U618 (N_618,In_1283,In_121);
nand U619 (N_619,N_240,N_170);
xor U620 (N_620,In_607,In_1390);
nor U621 (N_621,In_1479,In_1914);
xnor U622 (N_622,N_496,N_58);
nand U623 (N_623,In_1851,In_1963);
xor U624 (N_624,In_1170,In_380);
and U625 (N_625,In_1527,In_1573);
and U626 (N_626,In_745,In_1776);
and U627 (N_627,N_46,In_1233);
nor U628 (N_628,N_349,In_1814);
nand U629 (N_629,In_711,N_386);
and U630 (N_630,N_72,N_413);
and U631 (N_631,In_966,In_1125);
and U632 (N_632,In_314,N_23);
or U633 (N_633,In_1180,N_300);
or U634 (N_634,In_1063,N_481);
nand U635 (N_635,In_1160,In_717);
nor U636 (N_636,In_1490,In_798);
and U637 (N_637,In_1651,In_1228);
xnor U638 (N_638,In_1818,N_395);
or U639 (N_639,In_621,In_1247);
and U640 (N_640,In_1171,In_114);
nand U641 (N_641,N_465,N_486);
or U642 (N_642,In_407,N_195);
and U643 (N_643,In_291,N_114);
or U644 (N_644,In_803,N_303);
and U645 (N_645,In_1515,N_139);
nor U646 (N_646,N_276,In_801);
and U647 (N_647,In_714,N_209);
or U648 (N_648,N_28,In_1652);
and U649 (N_649,In_1446,In_1643);
or U650 (N_650,In_335,In_1404);
nor U651 (N_651,In_216,In_558);
and U652 (N_652,N_117,In_277);
or U653 (N_653,In_1951,N_275);
nand U654 (N_654,In_944,N_241);
nor U655 (N_655,In_804,In_224);
and U656 (N_656,In_643,In_164);
or U657 (N_657,In_1258,In_825);
nand U658 (N_658,In_69,In_1269);
or U659 (N_659,In_1300,N_442);
xnor U660 (N_660,In_705,In_254);
nor U661 (N_661,In_1154,In_1805);
nand U662 (N_662,In_504,In_393);
and U663 (N_663,In_406,N_440);
nor U664 (N_664,In_571,N_344);
nor U665 (N_665,In_1079,In_653);
nor U666 (N_666,In_70,In_1522);
nor U667 (N_667,N_31,In_976);
and U668 (N_668,N_376,In_833);
nor U669 (N_669,N_453,N_223);
xor U670 (N_670,N_399,In_878);
xor U671 (N_671,N_306,In_1369);
nand U672 (N_672,In_716,In_549);
and U673 (N_673,In_328,N_434);
nand U674 (N_674,In_931,N_144);
xor U675 (N_675,In_1962,N_15);
or U676 (N_676,N_198,N_356);
nand U677 (N_677,In_1400,N_90);
nand U678 (N_678,In_4,In_428);
nand U679 (N_679,N_320,In_222);
nor U680 (N_680,N_284,In_1830);
or U681 (N_681,In_875,N_392);
or U682 (N_682,N_402,In_1717);
nand U683 (N_683,In_1947,N_228);
and U684 (N_684,In_1949,In_348);
xnor U685 (N_685,In_1382,In_1819);
xnor U686 (N_686,In_1842,N_332);
xnor U687 (N_687,In_1800,N_355);
nand U688 (N_688,In_441,In_1425);
xor U689 (N_689,N_485,In_1421);
nor U690 (N_690,In_1683,In_1313);
and U691 (N_691,N_194,In_1007);
nor U692 (N_692,In_585,In_104);
xnor U693 (N_693,In_632,In_1991);
and U694 (N_694,In_1978,N_315);
nor U695 (N_695,In_722,In_1424);
xnor U696 (N_696,In_1291,In_983);
xor U697 (N_697,In_204,In_1726);
or U698 (N_698,In_182,In_769);
nor U699 (N_699,In_1732,In_1271);
nand U700 (N_700,In_1973,N_308);
and U701 (N_701,N_141,In_1443);
nor U702 (N_702,In_1122,N_233);
and U703 (N_703,In_1452,In_1552);
nor U704 (N_704,N_391,In_1408);
and U705 (N_705,In_942,In_474);
xnor U706 (N_706,N_278,N_0);
xor U707 (N_707,In_1911,In_899);
nand U708 (N_708,In_127,In_1894);
and U709 (N_709,N_123,In_108);
nand U710 (N_710,In_726,In_1764);
and U711 (N_711,N_478,In_147);
xnor U712 (N_712,In_39,In_1589);
or U713 (N_713,N_29,In_900);
xor U714 (N_714,In_157,N_310);
or U715 (N_715,In_374,In_810);
nor U716 (N_716,In_858,In_469);
nor U717 (N_717,In_1172,N_187);
nor U718 (N_718,In_783,In_268);
nor U719 (N_719,In_1077,In_1619);
nand U720 (N_720,In_1792,In_545);
xor U721 (N_721,In_807,In_1500);
and U722 (N_722,In_1635,N_322);
and U723 (N_723,In_1866,In_272);
or U724 (N_724,In_1461,N_311);
and U725 (N_725,In_1364,In_1492);
nor U726 (N_726,N_249,N_271);
and U727 (N_727,In_284,N_419);
and U728 (N_728,In_873,In_1287);
nand U729 (N_729,In_962,In_1092);
nor U730 (N_730,In_1124,In_739);
xor U731 (N_731,In_336,In_1050);
nand U732 (N_732,In_1826,In_1489);
and U733 (N_733,N_26,In_530);
or U734 (N_734,In_1675,In_1241);
or U735 (N_735,N_148,In_720);
nor U736 (N_736,In_1005,In_721);
or U737 (N_737,N_212,In_1926);
nand U738 (N_738,N_273,In_340);
nor U739 (N_739,In_815,In_828);
or U740 (N_740,In_1898,In_1663);
nand U741 (N_741,N_61,N_81);
and U742 (N_742,N_242,N_316);
nor U743 (N_743,In_816,In_425);
nand U744 (N_744,N_378,In_753);
or U745 (N_745,N_294,In_1576);
nor U746 (N_746,In_1181,In_615);
xor U747 (N_747,In_955,In_124);
and U748 (N_748,In_1782,In_223);
nor U749 (N_749,In_1971,In_1142);
and U750 (N_750,N_266,N_723);
nor U751 (N_751,In_1001,N_83);
nor U752 (N_752,In_793,N_683);
xor U753 (N_753,N_597,N_572);
and U754 (N_754,In_1031,N_237);
xnor U755 (N_755,In_339,N_253);
and U756 (N_756,In_37,N_466);
or U757 (N_757,In_1185,N_578);
xnor U758 (N_758,N_350,N_293);
nor U759 (N_759,In_1584,In_570);
xor U760 (N_760,N_634,N_653);
nand U761 (N_761,In_111,N_67);
or U762 (N_762,N_79,In_507);
nand U763 (N_763,In_1457,In_526);
nand U764 (N_764,N_104,N_508);
xnor U765 (N_765,In_887,In_427);
or U766 (N_766,In_158,N_42);
or U767 (N_767,In_437,N_555);
nand U768 (N_768,In_682,N_613);
nand U769 (N_769,In_1462,In_1916);
and U770 (N_770,In_1431,In_273);
nand U771 (N_771,N_272,N_415);
nand U772 (N_772,In_1152,N_296);
nand U773 (N_773,In_205,In_1587);
and U774 (N_774,N_397,In_857);
or U775 (N_775,In_275,In_1121);
and U776 (N_776,N_733,In_12);
or U777 (N_777,N_544,N_191);
and U778 (N_778,In_1989,In_852);
and U779 (N_779,In_620,In_1993);
xnor U780 (N_780,In_1146,N_715);
nand U781 (N_781,In_1871,N_514);
and U782 (N_782,N_539,N_27);
nand U783 (N_783,In_229,N_611);
nor U784 (N_784,In_1344,In_1268);
and U785 (N_785,In_1261,In_1483);
or U786 (N_786,In_1296,In_1347);
or U787 (N_787,In_227,N_643);
and U788 (N_788,N_598,N_741);
xor U789 (N_789,In_650,In_28);
nand U790 (N_790,In_1290,In_1215);
nand U791 (N_791,N_552,In_1569);
xnor U792 (N_792,In_1074,In_579);
nand U793 (N_793,In_1141,In_1203);
and U794 (N_794,In_1029,In_197);
xor U795 (N_795,In_568,N_661);
nor U796 (N_796,In_987,In_18);
xnor U797 (N_797,In_1610,In_775);
xor U798 (N_798,N_14,N_18);
or U799 (N_799,In_1356,In_283);
nand U800 (N_800,N_669,In_1752);
and U801 (N_801,N_536,In_1561);
nor U802 (N_802,In_641,N_569);
nor U803 (N_803,In_896,In_542);
xnor U804 (N_804,In_353,N_412);
nand U805 (N_805,N_394,In_1647);
and U806 (N_806,N_666,N_609);
nand U807 (N_807,N_646,In_1945);
nand U808 (N_808,N_457,N_475);
and U809 (N_809,In_405,In_1690);
and U810 (N_810,N_200,In_589);
xor U811 (N_811,N_309,In_1644);
nor U812 (N_812,In_1832,In_645);
and U813 (N_813,In_1557,N_360);
xor U814 (N_814,In_1767,In_689);
xnor U815 (N_815,N_298,In_198);
and U816 (N_816,In_1069,In_119);
and U817 (N_817,N_285,In_201);
xor U818 (N_818,N_55,In_996);
nor U819 (N_819,In_1634,In_599);
or U820 (N_820,In_902,In_508);
or U821 (N_821,N_204,In_267);
xor U822 (N_822,In_1293,In_1012);
nor U823 (N_823,N_205,N_477);
and U824 (N_824,In_569,In_289);
nand U825 (N_825,In_503,In_499);
and U826 (N_826,In_358,In_1406);
xor U827 (N_827,N_701,N_425);
nand U828 (N_828,In_742,In_1091);
nor U829 (N_829,N_580,In_856);
nor U830 (N_830,N_98,In_1650);
and U831 (N_831,N_565,N_125);
or U832 (N_832,In_1740,In_812);
xor U833 (N_833,In_1076,N_220);
nor U834 (N_834,In_1904,N_357);
nand U835 (N_835,N_431,N_749);
or U836 (N_836,In_1398,In_1272);
or U837 (N_837,In_142,In_1755);
nor U838 (N_838,N_464,N_129);
nor U839 (N_839,N_471,In_837);
xor U840 (N_840,In_99,N_250);
nand U841 (N_841,In_626,In_1599);
nand U842 (N_842,In_911,In_1965);
and U843 (N_843,In_1008,In_345);
xor U844 (N_844,N_564,N_96);
and U845 (N_845,In_60,N_705);
and U846 (N_846,In_449,N_283);
or U847 (N_847,In_1824,In_1994);
or U848 (N_848,In_1579,In_1299);
nor U849 (N_849,In_1939,In_977);
nor U850 (N_850,In_65,In_544);
nand U851 (N_851,In_1219,N_585);
and U852 (N_852,In_214,In_1823);
nand U853 (N_853,N_450,N_658);
and U854 (N_854,N_348,In_1045);
and U855 (N_855,N_182,In_1251);
or U856 (N_856,N_383,N_281);
nor U857 (N_857,In_1036,In_697);
nand U858 (N_858,In_870,In_1815);
or U859 (N_859,N_186,In_1689);
and U860 (N_860,N_261,In_521);
xor U861 (N_861,In_458,N_739);
and U862 (N_862,In_1715,In_495);
xor U863 (N_863,In_1450,In_1370);
xnor U864 (N_864,N_252,In_1923);
xnor U865 (N_865,In_1306,In_1237);
and U866 (N_866,N_469,In_194);
nand U867 (N_867,In_492,N_712);
and U868 (N_868,In_1594,In_1809);
xor U869 (N_869,N_638,In_1202);
and U870 (N_870,N_618,N_677);
xor U871 (N_871,In_1210,In_418);
and U872 (N_872,In_898,In_1938);
and U873 (N_873,In_397,In_639);
and U874 (N_874,In_1970,In_493);
or U875 (N_875,In_730,In_1182);
and U876 (N_876,In_588,N_660);
xor U877 (N_877,In_1793,In_1817);
and U878 (N_878,In_1279,N_566);
nor U879 (N_879,N_476,N_740);
or U880 (N_880,N_510,In_1549);
and U881 (N_881,N_255,In_402);
or U882 (N_882,N_387,In_1037);
or U883 (N_883,In_137,N_323);
xnor U884 (N_884,N_263,N_361);
nor U885 (N_885,In_889,In_1176);
and U886 (N_886,N_154,In_286);
nand U887 (N_887,N_495,N_714);
xor U888 (N_888,In_1674,N_560);
nand U889 (N_889,N_706,N_115);
xor U890 (N_890,In_1662,N_563);
nand U891 (N_891,In_741,N_615);
nor U892 (N_892,In_727,N_432);
or U893 (N_893,In_424,In_1780);
nor U894 (N_894,In_1288,In_1799);
nand U895 (N_895,In_1305,N_695);
xor U896 (N_896,In_1048,In_848);
or U897 (N_897,N_502,In_840);
nor U898 (N_898,N_663,In_912);
nand U899 (N_899,In_50,In_871);
nand U900 (N_900,N_329,N_470);
or U901 (N_901,In_357,N_541);
xnor U902 (N_902,In_1603,N_575);
nand U903 (N_903,In_1043,N_610);
or U904 (N_904,In_1016,N_730);
nand U905 (N_905,In_846,In_756);
and U906 (N_906,In_601,In_512);
nand U907 (N_907,In_881,In_138);
nor U908 (N_908,N_234,N_173);
and U909 (N_909,N_726,N_717);
and U910 (N_910,N_151,N_429);
xor U911 (N_911,In_1908,In_1178);
nor U912 (N_912,N_501,N_462);
and U913 (N_913,N_490,N_339);
xor U914 (N_914,In_1109,In_1656);
nand U915 (N_915,In_1312,N_143);
and U916 (N_916,N_206,In_1944);
or U917 (N_917,In_319,In_351);
xor U918 (N_918,N_532,In_1543);
or U919 (N_919,In_269,N_590);
or U920 (N_920,N_473,N_107);
or U921 (N_921,In_400,In_240);
nor U922 (N_922,N_87,In_1473);
nand U923 (N_923,N_594,In_1537);
nand U924 (N_924,In_422,In_298);
xor U925 (N_925,N_416,In_410);
or U926 (N_926,N_433,N_499);
or U927 (N_927,N_236,In_679);
nand U928 (N_928,N_400,In_143);
xor U929 (N_929,In_439,N_333);
nand U930 (N_930,N_605,In_225);
xnor U931 (N_931,In_937,In_1665);
nor U932 (N_932,In_1197,In_1136);
and U933 (N_933,In_893,N_279);
or U934 (N_934,In_1608,N_88);
or U935 (N_935,N_521,In_413);
xor U936 (N_936,N_679,N_737);
nand U937 (N_937,In_1417,N_352);
xnor U938 (N_938,In_945,N_498);
xnor U939 (N_939,N_372,In_255);
nand U940 (N_940,N_671,In_327);
or U941 (N_941,N_491,N_483);
xnor U942 (N_942,In_1753,N_729);
nand U943 (N_943,In_386,N_183);
or U944 (N_944,In_1724,In_1494);
or U945 (N_945,N_535,In_417);
nor U946 (N_946,In_1977,In_1518);
or U947 (N_947,In_1320,N_529);
xor U948 (N_948,N_518,In_1744);
or U949 (N_949,N_65,In_1011);
xor U950 (N_950,N_675,In_1838);
or U951 (N_951,In_952,N_277);
nand U952 (N_952,In_1891,In_1413);
or U953 (N_953,In_561,In_149);
nand U954 (N_954,In_3,N_423);
or U955 (N_955,N_103,In_1872);
and U956 (N_956,In_89,N_53);
nand U957 (N_957,In_81,N_553);
or U958 (N_958,N_244,In_455);
xor U959 (N_959,N_326,N_2);
nand U960 (N_960,In_1106,In_1810);
nor U961 (N_961,N_533,In_475);
xor U962 (N_962,In_1352,In_1434);
nand U963 (N_963,In_859,In_1133);
nand U964 (N_964,In_606,In_767);
xnor U965 (N_965,In_523,In_1035);
or U966 (N_966,N_84,In_1586);
nor U967 (N_967,In_565,N_576);
nor U968 (N_968,In_228,In_890);
nor U969 (N_969,N_617,In_800);
nor U970 (N_970,In_562,N_382);
or U971 (N_971,In_171,In_1588);
or U972 (N_972,In_1367,In_1624);
and U973 (N_973,N_674,In_779);
nor U974 (N_974,N_710,N_119);
or U975 (N_975,In_467,N_673);
nor U976 (N_976,N_334,N_637);
nor U977 (N_977,N_368,N_451);
nand U978 (N_978,In_1517,N_691);
xnor U979 (N_979,In_1999,N_684);
nand U980 (N_980,N_688,In_829);
nor U981 (N_981,N_257,N_649);
or U982 (N_982,In_770,In_152);
nand U983 (N_983,N_438,N_724);
nand U984 (N_984,In_740,N_358);
xnor U985 (N_985,N_274,In_1580);
nand U986 (N_986,N_517,N_619);
nand U987 (N_987,In_1089,N_418);
nand U988 (N_988,N_685,In_1231);
nand U989 (N_989,In_1544,In_667);
nand U990 (N_990,In_454,In_1931);
nand U991 (N_991,N_133,N_550);
xnor U992 (N_992,In_1395,In_972);
nand U993 (N_993,In_764,N_460);
or U994 (N_994,N_426,N_522);
xor U995 (N_995,N_128,N_448);
nor U996 (N_996,In_790,In_1946);
or U997 (N_997,In_1623,In_1068);
xnor U998 (N_998,In_533,In_1604);
nand U999 (N_999,In_1467,N_528);
nor U1000 (N_1000,In_497,In_958);
xor U1001 (N_1001,N_796,In_1470);
and U1002 (N_1002,N_963,N_805);
or U1003 (N_1003,N_779,In_973);
nand U1004 (N_1004,In_971,In_1605);
xnor U1005 (N_1005,In_1403,N_534);
nand U1006 (N_1006,In_1948,N_866);
or U1007 (N_1007,N_595,In_350);
nor U1008 (N_1008,In_1351,In_1295);
nand U1009 (N_1009,In_1107,In_1354);
or U1010 (N_1010,N_346,In_102);
or U1011 (N_1011,N_877,In_1972);
or U1012 (N_1012,In_1664,In_604);
xnor U1013 (N_1013,In_1188,N_633);
xor U1014 (N_1014,N_792,N_996);
xor U1015 (N_1015,N_962,N_390);
nand U1016 (N_1016,In_1648,N_771);
xor U1017 (N_1017,N_854,N_581);
nor U1018 (N_1018,N_887,N_628);
nand U1019 (N_1019,In_478,In_237);
nor U1020 (N_1020,N_629,N_886);
nor U1021 (N_1021,N_853,In_1976);
nor U1022 (N_1022,N_914,In_789);
and U1023 (N_1023,N_213,N_863);
xnor U1024 (N_1024,N_509,In_954);
or U1025 (N_1025,In_1358,N_21);
nor U1026 (N_1026,In_258,N_907);
or U1027 (N_1027,In_341,In_598);
and U1028 (N_1028,N_836,In_184);
and U1029 (N_1029,N_632,N_286);
nand U1030 (N_1030,N_369,In_1760);
and U1031 (N_1031,N_976,N_829);
xnor U1032 (N_1032,N_862,In_1551);
or U1033 (N_1033,In_999,N_991);
xor U1034 (N_1034,N_338,N_767);
and U1035 (N_1035,N_331,In_212);
xor U1036 (N_1036,In_274,In_333);
nor U1037 (N_1037,In_1616,N_876);
nor U1038 (N_1038,In_981,In_1447);
nand U1039 (N_1039,N_871,N_232);
nor U1040 (N_1040,In_1609,In_1640);
or U1041 (N_1041,N_527,N_847);
xor U1042 (N_1042,In_1426,In_1108);
nor U1043 (N_1043,In_1034,N_939);
nor U1044 (N_1044,In_306,N_584);
nand U1045 (N_1045,N_699,In_782);
and U1046 (N_1046,N_708,In_1542);
xor U1047 (N_1047,N_282,In_888);
nor U1048 (N_1048,N_953,N_689);
nand U1049 (N_1049,N_865,N_484);
or U1050 (N_1050,In_1280,In_151);
nor U1051 (N_1051,N_844,N_428);
or U1052 (N_1052,In_617,N_917);
and U1053 (N_1053,N_512,N_157);
nand U1054 (N_1054,N_786,In_96);
xor U1055 (N_1055,N_264,N_612);
xnor U1056 (N_1056,In_1513,In_538);
nor U1057 (N_1057,N_446,In_841);
nand U1058 (N_1058,N_551,In_1482);
and U1059 (N_1059,In_1411,N_816);
nor U1060 (N_1060,N_336,In_761);
nand U1061 (N_1061,In_1857,N_915);
nor U1062 (N_1062,N_875,N_881);
nor U1063 (N_1063,N_289,N_622);
or U1064 (N_1064,In_1632,N_302);
and U1065 (N_1065,N_930,In_1028);
or U1066 (N_1066,N_872,N_943);
nand U1067 (N_1067,N_126,In_303);
xnor U1068 (N_1068,In_219,In_822);
or U1069 (N_1069,In_628,N_577);
or U1070 (N_1070,In_885,In_1873);
and U1071 (N_1071,In_330,N_6);
and U1072 (N_1072,In_1516,In_187);
nor U1073 (N_1073,In_1721,N_954);
or U1074 (N_1074,In_785,N_106);
nor U1075 (N_1075,N_922,N_603);
nand U1076 (N_1076,In_805,N_910);
and U1077 (N_1077,N_422,In_446);
or U1078 (N_1078,N_600,N_838);
and U1079 (N_1079,In_1476,N_870);
nor U1080 (N_1080,N_759,In_1889);
and U1081 (N_1081,In_515,N_9);
and U1082 (N_1082,N_802,N_164);
xnor U1083 (N_1083,N_889,N_22);
and U1084 (N_1084,N_80,N_681);
nor U1085 (N_1085,N_807,N_831);
xor U1086 (N_1086,In_1713,N_401);
nor U1087 (N_1087,N_687,In_1621);
or U1088 (N_1088,N_776,In_1909);
or U1089 (N_1089,N_659,N_647);
nand U1090 (N_1090,In_953,In_445);
and U1091 (N_1091,In_762,N_946);
and U1092 (N_1092,In_1365,In_1437);
and U1093 (N_1093,In_1099,In_1263);
xor U1094 (N_1094,N_630,N_885);
nand U1095 (N_1095,In_1708,In_1661);
nand U1096 (N_1096,N_722,In_236);
xnor U1097 (N_1097,N_111,N_867);
or U1098 (N_1098,N_902,N_955);
and U1099 (N_1099,N_923,In_1781);
nor U1100 (N_1100,N_207,N_967);
or U1101 (N_1101,N_803,N_69);
nor U1102 (N_1102,In_1677,In_1614);
nand U1103 (N_1103,In_1039,N_254);
or U1104 (N_1104,N_225,In_53);
nand U1105 (N_1105,N_427,N_692);
nand U1106 (N_1106,N_849,In_440);
xnor U1107 (N_1107,N_105,In_442);
xor U1108 (N_1108,In_481,In_1126);
xnor U1109 (N_1109,In_1368,N_270);
nor U1110 (N_1110,In_880,N_362);
xnor U1111 (N_1111,N_468,In_1316);
or U1112 (N_1112,N_992,N_855);
xnor U1113 (N_1113,N_903,N_91);
xor U1114 (N_1114,N_817,N_201);
nand U1115 (N_1115,N_795,N_896);
or U1116 (N_1116,N_756,N_327);
nand U1117 (N_1117,N_494,In_1628);
and U1118 (N_1118,N_919,In_112);
and U1119 (N_1119,In_915,N_750);
nand U1120 (N_1120,N_530,N_958);
or U1121 (N_1121,N_813,N_950);
or U1122 (N_1122,N_703,In_56);
or U1123 (N_1123,N_707,In_220);
or U1124 (N_1124,N_70,In_68);
and U1125 (N_1125,N_662,In_1602);
nor U1126 (N_1126,In_302,N_482);
nand U1127 (N_1127,N_821,In_1575);
and U1128 (N_1128,N_547,In_383);
and U1129 (N_1129,In_1222,In_1073);
and U1130 (N_1130,N_654,N_837);
nor U1131 (N_1131,In_1533,In_1679);
nor U1132 (N_1132,N_591,In_176);
and U1133 (N_1133,N_841,In_1270);
or U1134 (N_1134,In_747,In_1275);
nor U1135 (N_1135,N_811,In_51);
xnor U1136 (N_1136,In_1084,N_268);
nand U1137 (N_1137,In_1686,In_527);
and U1138 (N_1138,In_930,N_678);
or U1139 (N_1139,In_1701,N_1);
nor U1140 (N_1140,N_941,N_158);
nand U1141 (N_1141,In_1560,N_754);
nand U1142 (N_1142,N_665,N_280);
nor U1143 (N_1143,In_693,N_635);
nand U1144 (N_1144,In_334,In_215);
or U1145 (N_1145,In_1078,N_616);
nand U1146 (N_1146,In_564,In_1336);
xor U1147 (N_1147,N_713,N_89);
and U1148 (N_1148,N_947,N_113);
or U1149 (N_1149,N_738,In_614);
nand U1150 (N_1150,N_956,In_1235);
xnor U1151 (N_1151,In_349,In_146);
nand U1152 (N_1152,N_301,N_64);
or U1153 (N_1153,In_773,In_9);
nand U1154 (N_1154,N_752,N_744);
nand U1155 (N_1155,N_899,N_960);
and U1156 (N_1156,In_1056,In_1147);
nor U1157 (N_1157,In_1345,N_642);
nor U1158 (N_1158,N_359,N_809);
and U1159 (N_1159,In_5,N_964);
xnor U1160 (N_1160,N_908,In_1958);
nor U1161 (N_1161,N_719,In_623);
or U1162 (N_1162,In_862,N_690);
xnor U1163 (N_1163,N_52,In_1880);
or U1164 (N_1164,N_500,In_1709);
nand U1165 (N_1165,N_589,In_15);
xor U1166 (N_1166,N_952,N_932);
nor U1167 (N_1167,N_570,In_1700);
xor U1168 (N_1168,N_371,N_850);
nand U1169 (N_1169,N_788,N_682);
nand U1170 (N_1170,N_380,In_1716);
or U1171 (N_1171,In_1238,N_116);
or U1172 (N_1172,N_516,N_997);
xnor U1173 (N_1173,In_1200,N_11);
or U1174 (N_1174,N_456,N_725);
and U1175 (N_1175,In_490,N_367);
nor U1176 (N_1176,N_861,N_625);
and U1177 (N_1177,In_1114,N_559);
nor U1178 (N_1178,In_1555,N_913);
nor U1179 (N_1179,N_893,N_969);
or U1180 (N_1180,In_865,In_877);
nand U1181 (N_1181,N_319,N_822);
xor U1182 (N_1182,In_218,In_1510);
nand U1183 (N_1183,N_757,N_858);
and U1184 (N_1184,N_488,N_973);
nand U1185 (N_1185,N_696,In_702);
and U1186 (N_1186,N_124,In_210);
or U1187 (N_1187,In_97,N_489);
and U1188 (N_1188,N_549,In_1888);
and U1189 (N_1189,N_895,In_1788);
nor U1190 (N_1190,N_981,N_455);
nor U1191 (N_1191,N_265,N_927);
xor U1192 (N_1192,In_1294,N_897);
xnor U1193 (N_1193,In_552,In_33);
xor U1194 (N_1194,N_406,N_398);
and U1195 (N_1195,N_975,N_62);
or U1196 (N_1196,N_755,N_672);
nor U1197 (N_1197,N_959,N_17);
xor U1198 (N_1198,N_929,N_736);
and U1199 (N_1199,In_1553,N_839);
nor U1200 (N_1200,N_951,In_67);
nor U1201 (N_1201,N_657,N_883);
or U1202 (N_1202,In_416,In_31);
or U1203 (N_1203,In_591,N_859);
and U1204 (N_1204,In_177,N_365);
nor U1205 (N_1205,N_731,In_936);
or U1206 (N_1206,N_906,N_709);
xnor U1207 (N_1207,N_732,N_970);
nand U1208 (N_1208,N_587,In_681);
xor U1209 (N_1209,In_1264,In_1394);
nand U1210 (N_1210,N_122,In_528);
or U1211 (N_1211,N_989,In_609);
nor U1212 (N_1212,In_312,In_774);
xor U1213 (N_1213,In_578,N_894);
xnor U1214 (N_1214,In_326,In_510);
or U1215 (N_1215,N_291,N_905);
nand U1216 (N_1216,N_670,N_304);
or U1217 (N_1217,N_437,In_1044);
nand U1218 (N_1218,N_39,N_827);
and U1219 (N_1219,In_1852,N_721);
and U1220 (N_1220,N_235,N_351);
nor U1221 (N_1221,In_795,In_1763);
nor U1222 (N_1222,N_363,N_515);
or U1223 (N_1223,In_1164,N_784);
xnor U1224 (N_1224,In_128,In_1613);
xnor U1225 (N_1225,In_1733,In_1954);
or U1226 (N_1226,In_1298,In_1038);
or U1227 (N_1227,In_1021,N_869);
nor U1228 (N_1228,N_648,N_614);
nand U1229 (N_1229,N_986,N_892);
or U1230 (N_1230,N_993,N_414);
nor U1231 (N_1231,N_765,In_409);
and U1232 (N_1232,N_596,N_375);
nand U1233 (N_1233,N_606,N_656);
or U1234 (N_1234,N_345,In_547);
nor U1235 (N_1235,N_66,In_1468);
xor U1236 (N_1236,N_768,N_542);
nor U1237 (N_1237,In_1262,N_987);
nor U1238 (N_1238,In_1806,In_820);
nor U1239 (N_1239,N_44,N_974);
and U1240 (N_1240,N_262,N_639);
nor U1241 (N_1241,N_86,N_808);
nand U1242 (N_1242,N_19,N_258);
nand U1243 (N_1243,In_1257,In_988);
xor U1244 (N_1244,N_621,N_999);
xnor U1245 (N_1245,In_1881,In_27);
nand U1246 (N_1246,In_74,N_888);
and U1247 (N_1247,N_977,N_790);
nor U1248 (N_1248,In_691,In_1310);
xor U1249 (N_1249,In_1995,In_1710);
and U1250 (N_1250,N_568,N_770);
and U1251 (N_1251,N_833,N_1144);
and U1252 (N_1252,N_1096,In_1591);
or U1253 (N_1253,N_698,N_920);
and U1254 (N_1254,In_991,N_599);
nor U1255 (N_1255,In_1670,N_297);
xor U1256 (N_1256,In_1653,N_586);
and U1257 (N_1257,N_608,In_780);
and U1258 (N_1258,N_680,N_781);
nand U1259 (N_1259,N_118,N_1082);
xnor U1260 (N_1260,N_1225,N_980);
and U1261 (N_1261,N_1138,N_644);
nor U1262 (N_1262,In_1389,N_405);
and U1263 (N_1263,N_624,In_1766);
nor U1264 (N_1264,N_1071,N_54);
and U1265 (N_1265,N_938,N_652);
nand U1266 (N_1266,N_763,N_783);
xor U1267 (N_1267,N_513,N_1222);
or U1268 (N_1268,In_868,N_1158);
and U1269 (N_1269,N_935,N_748);
nor U1270 (N_1270,N_890,N_623);
or U1271 (N_1271,N_1053,N_846);
and U1272 (N_1272,N_772,In_1802);
and U1273 (N_1273,N_880,N_526);
and U1274 (N_1274,N_150,In_519);
and U1275 (N_1275,In_1324,In_1667);
or U1276 (N_1276,In_1330,In_1503);
nand U1277 (N_1277,In_24,In_175);
and U1278 (N_1278,N_153,N_546);
xor U1279 (N_1279,N_824,N_702);
xor U1280 (N_1280,N_704,N_1062);
xor U1281 (N_1281,N_1102,In_1927);
or U1282 (N_1282,N_626,N_435);
nor U1283 (N_1283,In_1157,N_1151);
nor U1284 (N_1284,N_1230,N_1049);
or U1285 (N_1285,N_1123,N_1241);
and U1286 (N_1286,In_44,N_957);
or U1287 (N_1287,N_408,N_1001);
nand U1288 (N_1288,In_1474,N_773);
or U1289 (N_1289,In_978,N_313);
or U1290 (N_1290,In_1072,N_251);
and U1291 (N_1291,N_1083,In_423);
or U1292 (N_1292,N_983,N_882);
nor U1293 (N_1293,N_459,In_1738);
xor U1294 (N_1294,N_1040,In_246);
nand U1295 (N_1295,In_42,N_562);
nor U1296 (N_1296,N_1004,In_1000);
xnor U1297 (N_1297,In_1103,N_1186);
nand U1298 (N_1298,N_1226,In_1002);
nand U1299 (N_1299,In_1127,N_543);
and U1300 (N_1300,N_716,N_793);
nand U1301 (N_1301,N_1124,N_1206);
xor U1302 (N_1302,In_927,N_745);
and U1303 (N_1303,N_1129,N_1177);
nand U1304 (N_1304,N_968,N_1009);
xor U1305 (N_1305,N_1201,N_1061);
xnor U1306 (N_1306,N_1200,In_1480);
nor U1307 (N_1307,N_35,N_998);
xor U1308 (N_1308,N_461,N_1136);
nand U1309 (N_1309,N_1204,N_583);
xor U1310 (N_1310,N_1240,In_583);
xor U1311 (N_1311,N_868,N_940);
or U1312 (N_1312,In_1230,In_1469);
xor U1313 (N_1313,In_1353,In_57);
nand U1314 (N_1314,N_1173,N_480);
nand U1315 (N_1315,N_978,N_1088);
nor U1316 (N_1316,N_1018,In_189);
or U1317 (N_1317,N_574,N_1220);
and U1318 (N_1318,In_363,N_1030);
or U1319 (N_1319,In_1253,N_1090);
nand U1320 (N_1320,N_1111,N_814);
and U1321 (N_1321,N_1174,In_346);
nor U1322 (N_1322,N_131,In_1134);
xnor U1323 (N_1323,N_1209,N_1215);
nand U1324 (N_1324,N_1056,In_932);
and U1325 (N_1325,In_1485,In_30);
nor U1326 (N_1326,N_524,In_997);
and U1327 (N_1327,In_1297,N_806);
and U1328 (N_1328,In_1862,N_1003);
or U1329 (N_1329,In_1645,In_1451);
xnor U1330 (N_1330,N_1059,N_1162);
and U1331 (N_1331,N_911,N_664);
nor U1332 (N_1332,N_181,N_307);
nand U1333 (N_1333,N_40,N_1164);
nand U1334 (N_1334,N_1006,N_760);
nand U1335 (N_1335,N_918,N_1227);
nand U1336 (N_1336,N_161,N_1091);
or U1337 (N_1337,N_588,N_1079);
nor U1338 (N_1338,N_1092,N_165);
and U1339 (N_1339,N_761,N_966);
and U1340 (N_1340,In_10,In_1204);
xor U1341 (N_1341,In_376,In_995);
and U1342 (N_1342,N_720,N_1033);
and U1343 (N_1343,N_215,In_1615);
nand U1344 (N_1344,In_460,N_445);
xnor U1345 (N_1345,In_1041,In_1794);
or U1346 (N_1346,In_1322,In_618);
or U1347 (N_1347,In_1422,In_1812);
or U1348 (N_1348,N_511,N_891);
and U1349 (N_1349,N_1085,N_403);
nor U1350 (N_1350,In_308,N_1012);
nor U1351 (N_1351,N_1109,N_1211);
nand U1352 (N_1352,In_1874,N_1043);
and U1353 (N_1353,N_1228,In_1848);
or U1354 (N_1354,N_945,N_1008);
xor U1355 (N_1355,In_1987,In_1266);
nor U1356 (N_1356,N_1234,In_61);
and U1357 (N_1357,N_949,In_1066);
nand U1358 (N_1358,N_1089,N_800);
xor U1359 (N_1359,In_72,N_579);
nor U1360 (N_1360,N_830,N_121);
nor U1361 (N_1361,In_794,N_259);
xor U1362 (N_1362,N_556,N_523);
xnor U1363 (N_1363,In_759,N_295);
or U1364 (N_1364,N_505,N_85);
nor U1365 (N_1365,N_742,N_1191);
nand U1366 (N_1366,N_1233,N_627);
or U1367 (N_1367,N_925,N_1239);
and U1368 (N_1368,N_1148,In_725);
nor U1369 (N_1369,N_995,In_1581);
or U1370 (N_1370,N_1118,N_1041);
and U1371 (N_1371,N_1060,In_597);
xor U1372 (N_1372,N_1167,N_820);
nand U1373 (N_1373,N_1013,N_700);
nand U1374 (N_1374,N_743,In_1757);
and U1375 (N_1375,In_435,In_232);
and U1376 (N_1376,N_1184,In_838);
nand U1377 (N_1377,In_990,N_1027);
xor U1378 (N_1378,In_1957,In_1840);
xnor U1379 (N_1379,N_1183,In_1318);
xor U1380 (N_1380,N_1019,N_1168);
nor U1381 (N_1381,N_1031,N_1028);
xnor U1382 (N_1382,In_1301,N_385);
xnor U1383 (N_1383,N_1141,In_29);
nor U1384 (N_1384,N_540,N_620);
xnor U1385 (N_1385,N_60,N_1107);
xor U1386 (N_1386,N_794,N_531);
nand U1387 (N_1387,N_211,N_1178);
and U1388 (N_1388,N_290,N_751);
xnor U1389 (N_1389,In_654,N_851);
and U1390 (N_1390,In_1119,N_1103);
or U1391 (N_1391,In_1061,N_1156);
and U1392 (N_1392,N_780,N_819);
nand U1393 (N_1393,N_1149,N_718);
and U1394 (N_1394,N_592,N_1142);
or U1395 (N_1395,N_823,N_697);
and U1396 (N_1396,N_1198,N_520);
or U1397 (N_1397,N_1188,N_538);
or U1398 (N_1398,N_965,N_1157);
or U1399 (N_1399,N_1180,N_519);
xnor U1400 (N_1400,In_1153,N_812);
and U1401 (N_1401,N_856,N_668);
or U1402 (N_1402,In_537,N_1122);
and U1403 (N_1403,N_1237,N_972);
nand U1404 (N_1404,N_944,N_764);
nand U1405 (N_1405,N_1104,In_516);
nor U1406 (N_1406,In_517,N_217);
nor U1407 (N_1407,In_1711,N_256);
or U1408 (N_1408,N_694,N_1223);
or U1409 (N_1409,In_1952,N_1025);
or U1410 (N_1410,N_506,In_929);
xnor U1411 (N_1411,N_393,N_909);
or U1412 (N_1412,In_661,N_318);
xnor U1413 (N_1413,N_443,N_834);
nand U1414 (N_1414,N_1016,In_851);
or U1415 (N_1415,N_135,In_1902);
or U1416 (N_1416,In_1052,N_1036);
nand U1417 (N_1417,In_98,N_1093);
nand U1418 (N_1418,N_782,In_1915);
and U1419 (N_1419,N_1171,N_810);
nor U1420 (N_1420,N_828,N_1179);
xor U1421 (N_1421,N_379,In_1161);
or U1422 (N_1422,N_1193,In_1562);
nand U1423 (N_1423,In_92,N_1172);
or U1424 (N_1424,In_1040,N_1146);
xor U1425 (N_1425,In_1060,N_937);
or U1426 (N_1426,In_1292,N_1161);
or U1427 (N_1427,N_785,In_940);
xnor U1428 (N_1428,N_374,In_1598);
nor U1429 (N_1429,In_1,N_288);
or U1430 (N_1430,N_1189,N_601);
and U1431 (N_1431,N_734,N_758);
xor U1432 (N_1432,N_650,N_1087);
and U1433 (N_1433,N_1130,N_354);
nand U1434 (N_1434,N_775,N_985);
xor U1435 (N_1435,N_746,In_985);
or U1436 (N_1436,In_970,In_1882);
nor U1437 (N_1437,N_1219,In_40);
xnor U1438 (N_1438,In_1585,In_292);
and U1439 (N_1439,N_651,N_1246);
nor U1440 (N_1440,N_335,In_1558);
and U1441 (N_1441,N_1022,N_787);
and U1442 (N_1442,N_557,N_1097);
or U1443 (N_1443,N_1098,N_417);
xor U1444 (N_1444,N_818,N_1072);
and U1445 (N_1445,N_545,In_1342);
nor U1446 (N_1446,N_735,N_843);
xnor U1447 (N_1447,N_1106,In_1138);
nor U1448 (N_1448,N_1214,N_835);
and U1449 (N_1449,N_1132,N_1063);
and U1450 (N_1450,N_1113,N_874);
nor U1451 (N_1451,In_1834,In_453);
and U1452 (N_1452,N_979,In_1497);
xnor U1453 (N_1453,N_791,N_842);
or U1454 (N_1454,In_325,In_432);
nor U1455 (N_1455,N_1101,N_1067);
xor U1456 (N_1456,In_1375,N_292);
nand U1457 (N_1457,N_1011,In_1177);
nor U1458 (N_1458,N_825,In_1192);
or U1459 (N_1459,N_1015,N_573);
nand U1460 (N_1460,N_95,N_1133);
or U1461 (N_1461,N_848,N_826);
nand U1462 (N_1462,N_1038,N_63);
nor U1463 (N_1463,N_1137,N_1024);
or U1464 (N_1464,N_988,N_1169);
nor U1465 (N_1465,In_980,In_1321);
nor U1466 (N_1466,N_1086,In_118);
nor U1467 (N_1467,N_1210,N_324);
and U1468 (N_1468,In_1118,In_1669);
and U1469 (N_1469,N_567,In_1329);
nand U1470 (N_1470,N_1166,N_373);
nor U1471 (N_1471,In_1703,N_1170);
or U1472 (N_1472,In_1155,N_1153);
nand U1473 (N_1473,N_353,N_942);
nand U1474 (N_1474,N_341,In_879);
and U1475 (N_1475,N_1010,N_801);
nor U1476 (N_1476,N_1116,In_489);
nand U1477 (N_1477,N_852,In_757);
nand U1478 (N_1478,N_901,N_1020);
and U1479 (N_1479,N_1181,In_1054);
nand U1480 (N_1480,N_1114,N_990);
xnor U1481 (N_1481,N_857,N_525);
nand U1482 (N_1482,N_607,N_1002);
nand U1483 (N_1483,N_1029,N_305);
nand U1484 (N_1484,N_110,In_1590);
and U1485 (N_1485,N_667,In_574);
xnor U1486 (N_1486,N_269,N_1052);
nor U1487 (N_1487,In_1867,N_130);
nand U1488 (N_1488,N_1076,N_504);
xnor U1489 (N_1489,N_1017,N_798);
nand U1490 (N_1490,In_1712,N_898);
or U1491 (N_1491,N_436,N_503);
nor U1492 (N_1492,In_63,In_1596);
and U1493 (N_1493,In_959,In_844);
nand U1494 (N_1494,N_1119,N_1058);
and U1495 (N_1495,N_1217,N_1014);
or U1496 (N_1496,N_1190,N_507);
nand U1497 (N_1497,N_561,In_381);
and U1498 (N_1498,N_924,N_224);
and U1499 (N_1499,In_1943,N_593);
nor U1500 (N_1500,N_1139,N_1331);
xnor U1501 (N_1501,N_1175,N_1465);
nand U1502 (N_1502,N_1325,N_1334);
xor U1503 (N_1503,In_1554,N_1291);
and U1504 (N_1504,N_1486,N_1037);
and U1505 (N_1505,N_1110,N_1380);
and U1506 (N_1506,N_727,N_1248);
nand U1507 (N_1507,N_1476,In_1919);
nand U1508 (N_1508,In_884,N_655);
nand U1509 (N_1509,N_1326,N_1000);
or U1510 (N_1510,N_1152,N_1364);
nand U1511 (N_1511,N_1438,N_1224);
nor U1512 (N_1512,N_928,In_1574);
nand U1513 (N_1513,N_299,N_1268);
xor U1514 (N_1514,N_162,N_497);
nor U1515 (N_1515,N_1403,N_1430);
and U1516 (N_1516,N_1270,N_1046);
nand U1517 (N_1517,N_1277,N_1338);
and U1518 (N_1518,In_1402,N_1254);
xor U1519 (N_1519,N_832,N_1407);
nand U1520 (N_1520,N_537,N_916);
xor U1521 (N_1521,N_1352,N_1398);
or U1522 (N_1522,In_188,N_604);
xnor U1523 (N_1523,N_1069,N_1159);
or U1524 (N_1524,N_711,N_554);
nand U1525 (N_1525,N_1314,N_815);
or U1526 (N_1526,N_1371,N_1044);
nor U1527 (N_1527,N_1284,N_136);
nand U1528 (N_1528,In_894,N_1389);
nor U1529 (N_1529,N_1350,N_1290);
nand U1530 (N_1530,N_112,N_1303);
xnor U1531 (N_1531,N_1187,N_864);
nand U1532 (N_1532,N_1495,N_933);
nand U1533 (N_1533,N_1361,N_1035);
and U1534 (N_1534,N_1442,In_49);
and U1535 (N_1535,In_485,N_1464);
xor U1536 (N_1536,N_777,N_1192);
nor U1537 (N_1537,N_1399,N_492);
or U1538 (N_1538,N_1388,In_395);
or U1539 (N_1539,N_1327,N_1418);
xor U1540 (N_1540,N_1288,N_1381);
or U1541 (N_1541,N_179,N_1365);
xor U1542 (N_1542,N_789,In_1059);
or U1543 (N_1543,N_1112,N_1231);
and U1544 (N_1544,N_1221,N_1499);
xnor U1545 (N_1545,N_878,N_1340);
nand U1546 (N_1546,N_631,N_1251);
nand U1547 (N_1547,In_1568,N_1253);
nor U1548 (N_1548,N_1078,N_388);
and U1549 (N_1549,N_1283,N_1309);
nand U1550 (N_1550,N_1074,N_1354);
and U1551 (N_1551,In_394,N_1462);
nor U1552 (N_1552,N_1306,N_1417);
xnor U1553 (N_1553,N_1321,N_1426);
nand U1554 (N_1554,In_301,In_1714);
or U1555 (N_1555,N_1147,N_1304);
nor U1556 (N_1556,In_685,N_1199);
and U1557 (N_1557,N_1429,N_1134);
nor U1558 (N_1558,N_1126,In_1420);
xnor U1559 (N_1559,In_906,N_1279);
and U1560 (N_1560,N_1094,N_931);
nand U1561 (N_1561,In_1807,In_1929);
xor U1562 (N_1562,N_1026,N_1021);
nor U1563 (N_1563,In_1768,N_1366);
nor U1564 (N_1564,In_241,N_1475);
or U1565 (N_1565,N_1305,N_766);
and U1566 (N_1566,N_1333,N_1160);
xor U1567 (N_1567,N_1405,N_1066);
nand U1568 (N_1568,N_1497,N_1395);
or U1569 (N_1569,N_1266,N_1413);
and U1570 (N_1570,N_1478,N_1117);
xor U1571 (N_1571,N_1121,N_1441);
or U1572 (N_1572,N_1433,N_1460);
or U1573 (N_1573,N_1396,N_1347);
and U1574 (N_1574,N_1477,N_1362);
nor U1575 (N_1575,N_1294,N_1095);
nor U1576 (N_1576,N_762,N_1203);
nor U1577 (N_1577,N_1439,N_1255);
xnor U1578 (N_1578,In_378,In_85);
xnor U1579 (N_1579,N_971,N_1051);
nand U1580 (N_1580,N_1336,N_1348);
and U1581 (N_1581,N_1216,N_1456);
nor U1582 (N_1582,N_982,N_1100);
nand U1583 (N_1583,N_636,In_462);
nor U1584 (N_1584,N_1269,N_1424);
xnor U1585 (N_1585,N_845,N_1498);
or U1586 (N_1586,N_1257,In_344);
and U1587 (N_1587,N_1208,N_1472);
nor U1588 (N_1588,N_1341,N_1264);
and U1589 (N_1589,In_1386,In_35);
nand U1590 (N_1590,N_1384,N_1267);
and U1591 (N_1591,N_1489,N_1406);
xor U1592 (N_1592,N_1259,N_1369);
or U1593 (N_1593,N_1150,In_1582);
nand U1594 (N_1594,N_1034,N_1373);
nand U1595 (N_1595,N_1453,N_1400);
nand U1596 (N_1596,In_1444,N_904);
and U1597 (N_1597,N_1263,N_1084);
or U1598 (N_1598,N_1353,N_1285);
nor U1599 (N_1599,N_1372,N_1411);
or U1600 (N_1600,N_1292,N_1316);
xnor U1601 (N_1601,N_1392,N_1108);
xor U1602 (N_1602,N_778,In_513);
xnor U1603 (N_1603,N_1420,N_1408);
xor U1604 (N_1604,N_1434,N_1415);
nor U1605 (N_1605,N_1448,N_1163);
or U1606 (N_1606,N_1409,N_1330);
and U1607 (N_1607,N_1446,In_426);
nand U1608 (N_1608,N_1185,N_1073);
nand U1609 (N_1609,N_912,N_1443);
or U1610 (N_1610,N_994,N_1458);
or U1611 (N_1611,N_961,N_1493);
xor U1612 (N_1612,N_1232,N_1005);
nand U1613 (N_1613,N_728,In_367);
nor U1614 (N_1614,N_926,N_1466);
or U1615 (N_1615,N_1382,N_1391);
xnor U1616 (N_1616,N_1242,In_233);
and U1617 (N_1617,N_1205,N_1393);
xor U1618 (N_1618,N_1143,N_1485);
nor U1619 (N_1619,N_463,N_1351);
nor U1620 (N_1620,N_1455,N_1329);
xnor U1621 (N_1621,N_1322,N_1480);
or U1622 (N_1622,N_1344,N_1068);
xor U1623 (N_1623,N_1394,N_1436);
nor U1624 (N_1624,N_1310,N_1202);
xnor U1625 (N_1625,N_1401,In_1762);
xnor U1626 (N_1626,N_582,N_1140);
or U1627 (N_1627,N_1299,N_1235);
and U1628 (N_1628,N_1048,N_1377);
and U1629 (N_1629,N_1120,N_1236);
nor U1630 (N_1630,N_12,N_1295);
or U1631 (N_1631,N_1386,N_1479);
xor U1632 (N_1632,N_1282,N_1260);
and U1633 (N_1633,N_167,In_1820);
xnor U1634 (N_1634,In_1458,N_1368);
nor U1635 (N_1635,N_1474,In_1906);
and U1636 (N_1636,N_1057,N_1487);
xnor U1637 (N_1637,N_1482,N_602);
nor U1638 (N_1638,N_1467,N_1425);
or U1639 (N_1639,In_587,In_1260);
and U1640 (N_1640,N_1335,N_1463);
or U1641 (N_1641,In_1611,N_1302);
or U1642 (N_1642,N_1390,N_1451);
or U1643 (N_1643,N_873,N_1452);
nor U1644 (N_1644,N_1182,N_1346);
xor U1645 (N_1645,N_804,N_1432);
nor U1646 (N_1646,In_692,N_1280);
nand U1647 (N_1647,N_1375,N_797);
nor U1648 (N_1648,N_1397,N_317);
and U1649 (N_1649,In_1225,N_1312);
nand U1650 (N_1650,N_1262,N_676);
nor U1651 (N_1651,N_1261,N_1449);
xnor U1652 (N_1652,N_774,In_299);
xor U1653 (N_1653,N_1265,N_1308);
nand U1654 (N_1654,N_1357,N_1339);
xor U1655 (N_1655,N_1212,N_1287);
xnor U1656 (N_1656,N_1278,N_1115);
nand U1657 (N_1657,N_1023,N_1296);
nor U1658 (N_1658,N_1307,N_1176);
or U1659 (N_1659,N_1065,N_1154);
and U1660 (N_1660,N_1337,N_1039);
nand U1661 (N_1661,N_879,N_1249);
xor U1662 (N_1662,N_1358,N_1374);
nor U1663 (N_1663,N_1454,In_914);
or U1664 (N_1664,N_1367,N_1050);
nor U1665 (N_1665,N_1055,N_1483);
xor U1666 (N_1666,N_1328,N_769);
or U1667 (N_1667,N_1473,N_1213);
and U1668 (N_1668,N_1385,N_1297);
nand U1669 (N_1669,N_641,N_1484);
nor U1670 (N_1670,In_1749,N_1468);
or U1671 (N_1671,N_1459,In_1578);
nand U1672 (N_1672,N_1243,In_88);
nor U1673 (N_1673,N_1323,N_1419);
xnor U1674 (N_1674,N_1054,N_421);
nand U1675 (N_1675,N_10,N_1422);
xor U1676 (N_1676,N_1080,N_1298);
xnor U1677 (N_1677,In_1844,N_1319);
nor U1678 (N_1678,N_921,N_1155);
xnor U1679 (N_1679,N_32,In_420);
nand U1680 (N_1680,In_1433,N_1165);
and U1681 (N_1681,In_1067,In_347);
xnor U1682 (N_1682,N_1428,N_1274);
xnor U1683 (N_1683,N_1281,N_1099);
or U1684 (N_1684,N_1194,N_1315);
xnor U1685 (N_1685,N_1356,N_1332);
nor U1686 (N_1686,N_1457,N_1324);
nand U1687 (N_1687,N_1427,N_1450);
xor U1688 (N_1688,N_1077,In_648);
nor U1689 (N_1689,N_389,N_1437);
nand U1690 (N_1690,N_1414,N_1320);
nor U1691 (N_1691,N_936,N_1423);
or U1692 (N_1692,N_1218,N_640);
xor U1693 (N_1693,N_1471,N_1342);
nand U1694 (N_1694,N_1064,N_1127);
or U1695 (N_1695,N_1032,N_1355);
nand U1696 (N_1696,In_245,N_1289);
or U1697 (N_1697,N_1379,N_1440);
nand U1698 (N_1698,N_458,N_1238);
nor U1699 (N_1699,N_1481,N_1445);
or U1700 (N_1700,N_1360,N_49);
xnor U1701 (N_1701,N_1421,N_1469);
and U1702 (N_1702,N_1359,N_132);
nor U1703 (N_1703,N_1229,N_1256);
and U1704 (N_1704,N_1416,In_1277);
xor U1705 (N_1705,N_1250,N_1490);
xnor U1706 (N_1706,N_747,N_1370);
xor U1707 (N_1707,N_686,N_1349);
and U1708 (N_1708,N_840,N_1343);
or U1709 (N_1709,N_1271,In_1355);
or U1710 (N_1710,N_1196,N_1293);
nand U1711 (N_1711,N_1258,N_1488);
or U1712 (N_1712,N_1272,N_1135);
nor U1713 (N_1713,N_1047,N_1276);
or U1714 (N_1714,N_1470,N_1007);
or U1715 (N_1715,N_571,N_1042);
xor U1716 (N_1716,N_753,N_1145);
or U1717 (N_1717,N_1131,N_1492);
xnor U1718 (N_1718,N_1496,N_693);
and U1719 (N_1719,N_900,N_1128);
or U1720 (N_1720,In_1435,N_1378);
or U1721 (N_1721,In_1083,N_1317);
xor U1722 (N_1722,N_1412,N_1081);
nor U1723 (N_1723,N_645,N_1494);
xor U1724 (N_1724,N_1363,N_1444);
or U1725 (N_1725,N_799,N_1410);
nand U1726 (N_1726,N_1461,N_1383);
or U1727 (N_1727,N_1301,N_934);
nor U1728 (N_1728,In_1704,In_546);
and U1729 (N_1729,N_229,N_1125);
xnor U1730 (N_1730,N_1318,N_984);
and U1731 (N_1731,N_1195,N_1387);
xor U1732 (N_1732,N_1075,N_1491);
or U1733 (N_1733,N_1404,N_1435);
nand U1734 (N_1734,N_1431,N_1245);
or U1735 (N_1735,N_1376,N_1447);
xnor U1736 (N_1736,N_1197,N_548);
nor U1737 (N_1737,N_1070,N_1402);
nand U1738 (N_1738,N_1207,N_1252);
or U1739 (N_1739,In_1745,N_860);
nand U1740 (N_1740,N_449,In_101);
nand U1741 (N_1741,N_1345,In_11);
nor U1742 (N_1742,N_1311,N_1247);
nor U1743 (N_1743,N_1273,N_1286);
nor U1744 (N_1744,In_706,N_948);
and U1745 (N_1745,N_1275,N_1300);
nor U1746 (N_1746,N_1045,In_483);
nand U1747 (N_1747,N_1313,N_1105);
xor U1748 (N_1748,N_558,In_1571);
xnor U1749 (N_1749,N_884,N_1244);
xnor U1750 (N_1750,N_1645,N_1635);
nand U1751 (N_1751,N_1585,N_1588);
nor U1752 (N_1752,N_1628,N_1622);
nand U1753 (N_1753,N_1662,N_1601);
xnor U1754 (N_1754,N_1652,N_1669);
and U1755 (N_1755,N_1729,N_1590);
nand U1756 (N_1756,N_1710,N_1515);
and U1757 (N_1757,N_1629,N_1688);
nor U1758 (N_1758,N_1686,N_1538);
and U1759 (N_1759,N_1717,N_1598);
xnor U1760 (N_1760,N_1626,N_1517);
nand U1761 (N_1761,N_1587,N_1728);
or U1762 (N_1762,N_1564,N_1520);
nand U1763 (N_1763,N_1655,N_1519);
and U1764 (N_1764,N_1618,N_1742);
xnor U1765 (N_1765,N_1604,N_1646);
or U1766 (N_1766,N_1595,N_1577);
and U1767 (N_1767,N_1674,N_1625);
or U1768 (N_1768,N_1746,N_1641);
nand U1769 (N_1769,N_1723,N_1580);
xnor U1770 (N_1770,N_1568,N_1738);
and U1771 (N_1771,N_1555,N_1518);
nor U1772 (N_1772,N_1648,N_1593);
nand U1773 (N_1773,N_1698,N_1614);
nor U1774 (N_1774,N_1737,N_1542);
and U1775 (N_1775,N_1512,N_1596);
xnor U1776 (N_1776,N_1511,N_1586);
xnor U1777 (N_1777,N_1687,N_1525);
xnor U1778 (N_1778,N_1666,N_1636);
or U1779 (N_1779,N_1623,N_1536);
xor U1780 (N_1780,N_1701,N_1554);
nor U1781 (N_1781,N_1672,N_1530);
xnor U1782 (N_1782,N_1720,N_1719);
and U1783 (N_1783,N_1600,N_1543);
xor U1784 (N_1784,N_1553,N_1748);
xor U1785 (N_1785,N_1664,N_1749);
or U1786 (N_1786,N_1615,N_1651);
or U1787 (N_1787,N_1691,N_1733);
xor U1788 (N_1788,N_1541,N_1714);
and U1789 (N_1789,N_1579,N_1649);
and U1790 (N_1790,N_1521,N_1613);
xor U1791 (N_1791,N_1703,N_1550);
nor U1792 (N_1792,N_1677,N_1633);
nand U1793 (N_1793,N_1642,N_1726);
and U1794 (N_1794,N_1708,N_1634);
or U1795 (N_1795,N_1574,N_1561);
xor U1796 (N_1796,N_1608,N_1523);
or U1797 (N_1797,N_1583,N_1685);
nand U1798 (N_1798,N_1702,N_1689);
and U1799 (N_1799,N_1697,N_1673);
or U1800 (N_1800,N_1548,N_1684);
and U1801 (N_1801,N_1599,N_1631);
nor U1802 (N_1802,N_1591,N_1531);
xnor U1803 (N_1803,N_1722,N_1718);
and U1804 (N_1804,N_1537,N_1569);
xor U1805 (N_1805,N_1675,N_1572);
and U1806 (N_1806,N_1527,N_1562);
xnor U1807 (N_1807,N_1658,N_1632);
xnor U1808 (N_1808,N_1731,N_1739);
and U1809 (N_1809,N_1667,N_1747);
nor U1810 (N_1810,N_1503,N_1606);
and U1811 (N_1811,N_1567,N_1712);
xnor U1812 (N_1812,N_1612,N_1724);
or U1813 (N_1813,N_1709,N_1610);
nand U1814 (N_1814,N_1681,N_1692);
and U1815 (N_1815,N_1556,N_1700);
nor U1816 (N_1816,N_1559,N_1683);
and U1817 (N_1817,N_1715,N_1547);
xnor U1818 (N_1818,N_1690,N_1603);
xor U1819 (N_1819,N_1506,N_1581);
nor U1820 (N_1820,N_1545,N_1736);
nor U1821 (N_1821,N_1741,N_1540);
nand U1822 (N_1822,N_1505,N_1609);
xnor U1823 (N_1823,N_1637,N_1639);
or U1824 (N_1824,N_1576,N_1529);
xor U1825 (N_1825,N_1693,N_1650);
or U1826 (N_1826,N_1734,N_1696);
nand U1827 (N_1827,N_1528,N_1549);
nand U1828 (N_1828,N_1661,N_1656);
xnor U1829 (N_1829,N_1510,N_1617);
or U1830 (N_1830,N_1566,N_1532);
xnor U1831 (N_1831,N_1565,N_1704);
nand U1832 (N_1832,N_1705,N_1627);
nand U1833 (N_1833,N_1605,N_1716);
xnor U1834 (N_1834,N_1653,N_1557);
xor U1835 (N_1835,N_1743,N_1589);
nor U1836 (N_1836,N_1575,N_1504);
nand U1837 (N_1837,N_1544,N_1644);
xor U1838 (N_1838,N_1670,N_1638);
and U1839 (N_1839,N_1699,N_1727);
xor U1840 (N_1840,N_1578,N_1732);
nor U1841 (N_1841,N_1630,N_1551);
nor U1842 (N_1842,N_1508,N_1501);
xnor U1843 (N_1843,N_1654,N_1745);
nor U1844 (N_1844,N_1721,N_1678);
or U1845 (N_1845,N_1694,N_1707);
nor U1846 (N_1846,N_1558,N_1659);
nand U1847 (N_1847,N_1660,N_1602);
nand U1848 (N_1848,N_1524,N_1647);
nand U1849 (N_1849,N_1725,N_1671);
or U1850 (N_1850,N_1500,N_1507);
nor U1851 (N_1851,N_1616,N_1607);
nand U1852 (N_1852,N_1582,N_1744);
nor U1853 (N_1853,N_1735,N_1679);
nor U1854 (N_1854,N_1665,N_1624);
or U1855 (N_1855,N_1621,N_1570);
nand U1856 (N_1856,N_1573,N_1502);
and U1857 (N_1857,N_1535,N_1516);
and U1858 (N_1858,N_1620,N_1546);
xor U1859 (N_1859,N_1513,N_1713);
nor U1860 (N_1860,N_1552,N_1740);
or U1861 (N_1861,N_1514,N_1730);
nand U1862 (N_1862,N_1584,N_1657);
and U1863 (N_1863,N_1682,N_1680);
and U1864 (N_1864,N_1594,N_1619);
or U1865 (N_1865,N_1509,N_1668);
nor U1866 (N_1866,N_1534,N_1663);
and U1867 (N_1867,N_1711,N_1611);
and U1868 (N_1868,N_1597,N_1676);
and U1869 (N_1869,N_1706,N_1560);
xnor U1870 (N_1870,N_1695,N_1592);
nor U1871 (N_1871,N_1526,N_1522);
nand U1872 (N_1872,N_1643,N_1533);
nor U1873 (N_1873,N_1640,N_1571);
or U1874 (N_1874,N_1563,N_1539);
nor U1875 (N_1875,N_1697,N_1535);
nand U1876 (N_1876,N_1696,N_1591);
or U1877 (N_1877,N_1571,N_1728);
nor U1878 (N_1878,N_1731,N_1662);
xor U1879 (N_1879,N_1612,N_1636);
xnor U1880 (N_1880,N_1555,N_1582);
and U1881 (N_1881,N_1721,N_1707);
or U1882 (N_1882,N_1550,N_1618);
nor U1883 (N_1883,N_1705,N_1564);
nand U1884 (N_1884,N_1735,N_1569);
nand U1885 (N_1885,N_1706,N_1697);
nor U1886 (N_1886,N_1618,N_1511);
nand U1887 (N_1887,N_1544,N_1583);
and U1888 (N_1888,N_1539,N_1561);
and U1889 (N_1889,N_1555,N_1553);
nand U1890 (N_1890,N_1549,N_1552);
xnor U1891 (N_1891,N_1539,N_1703);
nor U1892 (N_1892,N_1696,N_1729);
or U1893 (N_1893,N_1740,N_1526);
or U1894 (N_1894,N_1666,N_1534);
or U1895 (N_1895,N_1700,N_1735);
nand U1896 (N_1896,N_1600,N_1637);
nand U1897 (N_1897,N_1593,N_1579);
and U1898 (N_1898,N_1590,N_1672);
or U1899 (N_1899,N_1685,N_1722);
or U1900 (N_1900,N_1530,N_1646);
nand U1901 (N_1901,N_1500,N_1749);
and U1902 (N_1902,N_1720,N_1685);
xnor U1903 (N_1903,N_1560,N_1625);
or U1904 (N_1904,N_1634,N_1716);
xor U1905 (N_1905,N_1564,N_1627);
nor U1906 (N_1906,N_1733,N_1608);
nand U1907 (N_1907,N_1519,N_1658);
nor U1908 (N_1908,N_1573,N_1629);
and U1909 (N_1909,N_1742,N_1734);
nor U1910 (N_1910,N_1508,N_1742);
nand U1911 (N_1911,N_1555,N_1589);
nor U1912 (N_1912,N_1749,N_1731);
and U1913 (N_1913,N_1694,N_1594);
and U1914 (N_1914,N_1659,N_1550);
and U1915 (N_1915,N_1693,N_1701);
xor U1916 (N_1916,N_1720,N_1623);
and U1917 (N_1917,N_1550,N_1661);
and U1918 (N_1918,N_1690,N_1636);
or U1919 (N_1919,N_1730,N_1650);
nand U1920 (N_1920,N_1691,N_1664);
and U1921 (N_1921,N_1724,N_1655);
nand U1922 (N_1922,N_1563,N_1531);
xnor U1923 (N_1923,N_1585,N_1648);
or U1924 (N_1924,N_1592,N_1663);
xor U1925 (N_1925,N_1680,N_1588);
xnor U1926 (N_1926,N_1614,N_1623);
xor U1927 (N_1927,N_1708,N_1654);
xor U1928 (N_1928,N_1690,N_1609);
nand U1929 (N_1929,N_1636,N_1653);
nor U1930 (N_1930,N_1666,N_1536);
and U1931 (N_1931,N_1650,N_1654);
nor U1932 (N_1932,N_1701,N_1523);
and U1933 (N_1933,N_1666,N_1678);
nand U1934 (N_1934,N_1705,N_1729);
nor U1935 (N_1935,N_1503,N_1595);
nand U1936 (N_1936,N_1551,N_1624);
or U1937 (N_1937,N_1635,N_1513);
nor U1938 (N_1938,N_1559,N_1608);
and U1939 (N_1939,N_1540,N_1618);
nand U1940 (N_1940,N_1561,N_1583);
or U1941 (N_1941,N_1591,N_1511);
nand U1942 (N_1942,N_1659,N_1517);
xnor U1943 (N_1943,N_1712,N_1707);
xor U1944 (N_1944,N_1746,N_1662);
nor U1945 (N_1945,N_1612,N_1592);
xnor U1946 (N_1946,N_1722,N_1515);
and U1947 (N_1947,N_1695,N_1705);
or U1948 (N_1948,N_1634,N_1519);
or U1949 (N_1949,N_1521,N_1595);
or U1950 (N_1950,N_1634,N_1517);
or U1951 (N_1951,N_1612,N_1661);
nand U1952 (N_1952,N_1635,N_1604);
and U1953 (N_1953,N_1607,N_1608);
and U1954 (N_1954,N_1739,N_1511);
or U1955 (N_1955,N_1548,N_1634);
nor U1956 (N_1956,N_1707,N_1717);
or U1957 (N_1957,N_1649,N_1629);
or U1958 (N_1958,N_1501,N_1731);
or U1959 (N_1959,N_1595,N_1733);
and U1960 (N_1960,N_1632,N_1604);
and U1961 (N_1961,N_1729,N_1550);
or U1962 (N_1962,N_1562,N_1560);
or U1963 (N_1963,N_1649,N_1725);
or U1964 (N_1964,N_1550,N_1615);
nand U1965 (N_1965,N_1673,N_1694);
nand U1966 (N_1966,N_1729,N_1637);
nand U1967 (N_1967,N_1579,N_1696);
and U1968 (N_1968,N_1709,N_1653);
and U1969 (N_1969,N_1570,N_1687);
or U1970 (N_1970,N_1611,N_1718);
nand U1971 (N_1971,N_1655,N_1732);
nand U1972 (N_1972,N_1510,N_1589);
nand U1973 (N_1973,N_1592,N_1657);
nor U1974 (N_1974,N_1537,N_1749);
nand U1975 (N_1975,N_1565,N_1743);
or U1976 (N_1976,N_1628,N_1626);
or U1977 (N_1977,N_1716,N_1558);
or U1978 (N_1978,N_1535,N_1648);
and U1979 (N_1979,N_1525,N_1664);
or U1980 (N_1980,N_1734,N_1627);
nand U1981 (N_1981,N_1627,N_1723);
and U1982 (N_1982,N_1741,N_1683);
and U1983 (N_1983,N_1581,N_1540);
xor U1984 (N_1984,N_1614,N_1514);
nand U1985 (N_1985,N_1745,N_1681);
xor U1986 (N_1986,N_1709,N_1671);
and U1987 (N_1987,N_1620,N_1520);
and U1988 (N_1988,N_1528,N_1736);
nor U1989 (N_1989,N_1603,N_1643);
or U1990 (N_1990,N_1576,N_1604);
nor U1991 (N_1991,N_1718,N_1680);
xor U1992 (N_1992,N_1502,N_1688);
and U1993 (N_1993,N_1723,N_1560);
and U1994 (N_1994,N_1641,N_1639);
or U1995 (N_1995,N_1664,N_1730);
nor U1996 (N_1996,N_1663,N_1730);
xnor U1997 (N_1997,N_1589,N_1705);
and U1998 (N_1998,N_1608,N_1526);
nand U1999 (N_1999,N_1663,N_1708);
nor U2000 (N_2000,N_1816,N_1863);
xor U2001 (N_2001,N_1765,N_1870);
and U2002 (N_2002,N_1944,N_1905);
nor U2003 (N_2003,N_1864,N_1878);
or U2004 (N_2004,N_1935,N_1775);
xor U2005 (N_2005,N_1927,N_1914);
xor U2006 (N_2006,N_1912,N_1781);
xnor U2007 (N_2007,N_1777,N_1988);
nand U2008 (N_2008,N_1876,N_1916);
nand U2009 (N_2009,N_1883,N_1847);
or U2010 (N_2010,N_1875,N_1824);
nand U2011 (N_2011,N_1845,N_1807);
and U2012 (N_2012,N_1967,N_1750);
and U2013 (N_2013,N_1762,N_1974);
and U2014 (N_2014,N_1963,N_1831);
xor U2015 (N_2015,N_1932,N_1968);
or U2016 (N_2016,N_1838,N_1756);
and U2017 (N_2017,N_1990,N_1769);
and U2018 (N_2018,N_1774,N_1790);
or U2019 (N_2019,N_1778,N_1837);
nor U2020 (N_2020,N_1871,N_1799);
nor U2021 (N_2021,N_1923,N_1836);
nor U2022 (N_2022,N_1899,N_1810);
xnor U2023 (N_2023,N_1953,N_1853);
and U2024 (N_2024,N_1925,N_1809);
and U2025 (N_2025,N_1798,N_1868);
xnor U2026 (N_2026,N_1893,N_1766);
nand U2027 (N_2027,N_1957,N_1861);
nor U2028 (N_2028,N_1901,N_1813);
nor U2029 (N_2029,N_1977,N_1985);
or U2030 (N_2030,N_1773,N_1970);
nand U2031 (N_2031,N_1779,N_1909);
nor U2032 (N_2032,N_1789,N_1992);
nand U2033 (N_2033,N_1852,N_1751);
or U2034 (N_2034,N_1920,N_1827);
and U2035 (N_2035,N_1811,N_1800);
or U2036 (N_2036,N_1782,N_1894);
and U2037 (N_2037,N_1924,N_1821);
nor U2038 (N_2038,N_1939,N_1946);
xnor U2039 (N_2039,N_1973,N_1805);
and U2040 (N_2040,N_1951,N_1872);
xor U2041 (N_2041,N_1833,N_1846);
nand U2042 (N_2042,N_1928,N_1874);
nor U2043 (N_2043,N_1794,N_1856);
xnor U2044 (N_2044,N_1904,N_1999);
or U2045 (N_2045,N_1767,N_1843);
nor U2046 (N_2046,N_1753,N_1839);
or U2047 (N_2047,N_1884,N_1911);
nor U2048 (N_2048,N_1812,N_1942);
and U2049 (N_2049,N_1897,N_1995);
and U2050 (N_2050,N_1860,N_1896);
xnor U2051 (N_2051,N_1890,N_1961);
and U2052 (N_2052,N_1761,N_1998);
nand U2053 (N_2053,N_1826,N_1855);
nand U2054 (N_2054,N_1832,N_1981);
xnor U2055 (N_2055,N_1908,N_1980);
nand U2056 (N_2056,N_1880,N_1887);
xor U2057 (N_2057,N_1915,N_1776);
nor U2058 (N_2058,N_1784,N_1867);
nor U2059 (N_2059,N_1788,N_1888);
xnor U2060 (N_2060,N_1804,N_1785);
or U2061 (N_2061,N_1922,N_1934);
nor U2062 (N_2062,N_1994,N_1885);
nand U2063 (N_2063,N_1891,N_1969);
nor U2064 (N_2064,N_1921,N_1962);
and U2065 (N_2065,N_1848,N_1823);
xor U2066 (N_2066,N_1964,N_1933);
nor U2067 (N_2067,N_1989,N_1857);
nor U2068 (N_2068,N_1991,N_1941);
and U2069 (N_2069,N_1808,N_1792);
xor U2070 (N_2070,N_1772,N_1892);
nor U2071 (N_2071,N_1907,N_1997);
and U2072 (N_2072,N_1975,N_1768);
or U2073 (N_2073,N_1881,N_1903);
and U2074 (N_2074,N_1926,N_1952);
nand U2075 (N_2075,N_1917,N_1972);
nor U2076 (N_2076,N_1757,N_1954);
nand U2077 (N_2077,N_1976,N_1752);
and U2078 (N_2078,N_1770,N_1787);
and U2079 (N_2079,N_1820,N_1759);
and U2080 (N_2080,N_1818,N_1814);
nor U2081 (N_2081,N_1829,N_1929);
or U2082 (N_2082,N_1877,N_1986);
and U2083 (N_2083,N_1780,N_1950);
nand U2084 (N_2084,N_1858,N_1900);
and U2085 (N_2085,N_1793,N_1949);
nor U2086 (N_2086,N_1865,N_1869);
and U2087 (N_2087,N_1862,N_1987);
and U2088 (N_2088,N_1783,N_1859);
nor U2089 (N_2089,N_1936,N_1898);
nand U2090 (N_2090,N_1947,N_1822);
nor U2091 (N_2091,N_1930,N_1764);
nand U2092 (N_2092,N_1795,N_1802);
or U2093 (N_2093,N_1819,N_1830);
nor U2094 (N_2094,N_1786,N_1983);
and U2095 (N_2095,N_1806,N_1758);
or U2096 (N_2096,N_1797,N_1965);
xnor U2097 (N_2097,N_1948,N_1895);
and U2098 (N_2098,N_1910,N_1979);
and U2099 (N_2099,N_1854,N_1960);
nand U2100 (N_2100,N_1984,N_1791);
nand U2101 (N_2101,N_1817,N_1902);
or U2102 (N_2102,N_1815,N_1993);
nor U2103 (N_2103,N_1754,N_1913);
nor U2104 (N_2104,N_1842,N_1931);
nand U2105 (N_2105,N_1763,N_1834);
xnor U2106 (N_2106,N_1945,N_1849);
nand U2107 (N_2107,N_1840,N_1955);
nor U2108 (N_2108,N_1958,N_1971);
nand U2109 (N_2109,N_1918,N_1886);
nand U2110 (N_2110,N_1873,N_1879);
nor U2111 (N_2111,N_1835,N_1938);
or U2112 (N_2112,N_1959,N_1850);
and U2113 (N_2113,N_1919,N_1940);
xor U2114 (N_2114,N_1796,N_1966);
and U2115 (N_2115,N_1803,N_1828);
or U2116 (N_2116,N_1943,N_1825);
nand U2117 (N_2117,N_1866,N_1978);
or U2118 (N_2118,N_1982,N_1801);
nand U2119 (N_2119,N_1760,N_1841);
nand U2120 (N_2120,N_1755,N_1937);
nand U2121 (N_2121,N_1882,N_1956);
nor U2122 (N_2122,N_1851,N_1844);
and U2123 (N_2123,N_1771,N_1996);
and U2124 (N_2124,N_1889,N_1906);
or U2125 (N_2125,N_1840,N_1857);
nand U2126 (N_2126,N_1951,N_1853);
and U2127 (N_2127,N_1758,N_1777);
nand U2128 (N_2128,N_1836,N_1895);
nor U2129 (N_2129,N_1842,N_1871);
and U2130 (N_2130,N_1993,N_1951);
nor U2131 (N_2131,N_1901,N_1889);
nand U2132 (N_2132,N_1814,N_1989);
xor U2133 (N_2133,N_1910,N_1821);
nor U2134 (N_2134,N_1914,N_1880);
and U2135 (N_2135,N_1890,N_1999);
nand U2136 (N_2136,N_1903,N_1778);
nand U2137 (N_2137,N_1870,N_1993);
and U2138 (N_2138,N_1984,N_1991);
nand U2139 (N_2139,N_1841,N_1816);
or U2140 (N_2140,N_1971,N_1912);
nor U2141 (N_2141,N_1982,N_1805);
nand U2142 (N_2142,N_1974,N_1867);
nor U2143 (N_2143,N_1860,N_1853);
or U2144 (N_2144,N_1922,N_1919);
and U2145 (N_2145,N_1916,N_1752);
and U2146 (N_2146,N_1936,N_1863);
nor U2147 (N_2147,N_1830,N_1905);
nand U2148 (N_2148,N_1917,N_1786);
nand U2149 (N_2149,N_1787,N_1931);
nand U2150 (N_2150,N_1923,N_1929);
nor U2151 (N_2151,N_1961,N_1794);
nor U2152 (N_2152,N_1959,N_1839);
or U2153 (N_2153,N_1862,N_1794);
and U2154 (N_2154,N_1945,N_1761);
xnor U2155 (N_2155,N_1790,N_1914);
or U2156 (N_2156,N_1921,N_1772);
or U2157 (N_2157,N_1968,N_1854);
nand U2158 (N_2158,N_1875,N_1917);
nand U2159 (N_2159,N_1789,N_1918);
and U2160 (N_2160,N_1785,N_1767);
nor U2161 (N_2161,N_1908,N_1993);
nand U2162 (N_2162,N_1757,N_1822);
xor U2163 (N_2163,N_1893,N_1924);
xor U2164 (N_2164,N_1905,N_1921);
and U2165 (N_2165,N_1968,N_1796);
and U2166 (N_2166,N_1921,N_1943);
xor U2167 (N_2167,N_1774,N_1931);
nand U2168 (N_2168,N_1820,N_1817);
nand U2169 (N_2169,N_1922,N_1953);
or U2170 (N_2170,N_1942,N_1934);
xor U2171 (N_2171,N_1898,N_1816);
and U2172 (N_2172,N_1986,N_1941);
and U2173 (N_2173,N_1918,N_1803);
or U2174 (N_2174,N_1754,N_1957);
nor U2175 (N_2175,N_1896,N_1804);
nor U2176 (N_2176,N_1830,N_1848);
nor U2177 (N_2177,N_1813,N_1750);
nor U2178 (N_2178,N_1773,N_1913);
xor U2179 (N_2179,N_1965,N_1963);
and U2180 (N_2180,N_1778,N_1891);
nor U2181 (N_2181,N_1758,N_1750);
and U2182 (N_2182,N_1945,N_1991);
nor U2183 (N_2183,N_1940,N_1865);
or U2184 (N_2184,N_1871,N_1873);
and U2185 (N_2185,N_1994,N_1838);
and U2186 (N_2186,N_1824,N_1770);
nor U2187 (N_2187,N_1755,N_1826);
or U2188 (N_2188,N_1768,N_1817);
nor U2189 (N_2189,N_1868,N_1795);
nand U2190 (N_2190,N_1934,N_1791);
nor U2191 (N_2191,N_1883,N_1843);
or U2192 (N_2192,N_1961,N_1830);
or U2193 (N_2193,N_1869,N_1973);
or U2194 (N_2194,N_1753,N_1913);
and U2195 (N_2195,N_1762,N_1978);
nor U2196 (N_2196,N_1996,N_1815);
and U2197 (N_2197,N_1908,N_1883);
nand U2198 (N_2198,N_1855,N_1858);
or U2199 (N_2199,N_1999,N_1985);
nor U2200 (N_2200,N_1844,N_1969);
nand U2201 (N_2201,N_1964,N_1800);
and U2202 (N_2202,N_1928,N_1905);
nand U2203 (N_2203,N_1859,N_1840);
nor U2204 (N_2204,N_1993,N_1929);
and U2205 (N_2205,N_1874,N_1919);
nand U2206 (N_2206,N_1765,N_1899);
nor U2207 (N_2207,N_1879,N_1837);
nand U2208 (N_2208,N_1850,N_1855);
xnor U2209 (N_2209,N_1880,N_1933);
xnor U2210 (N_2210,N_1763,N_1920);
nand U2211 (N_2211,N_1999,N_1807);
xor U2212 (N_2212,N_1753,N_1883);
nor U2213 (N_2213,N_1836,N_1791);
or U2214 (N_2214,N_1771,N_1944);
and U2215 (N_2215,N_1804,N_1880);
nor U2216 (N_2216,N_1751,N_1903);
and U2217 (N_2217,N_1827,N_1760);
nand U2218 (N_2218,N_1986,N_1858);
and U2219 (N_2219,N_1905,N_1938);
xor U2220 (N_2220,N_1825,N_1840);
xnor U2221 (N_2221,N_1774,N_1995);
xor U2222 (N_2222,N_1765,N_1953);
or U2223 (N_2223,N_1908,N_1913);
or U2224 (N_2224,N_1972,N_1999);
or U2225 (N_2225,N_1829,N_1857);
and U2226 (N_2226,N_1807,N_1836);
or U2227 (N_2227,N_1925,N_1943);
or U2228 (N_2228,N_1771,N_1782);
nand U2229 (N_2229,N_1911,N_1922);
and U2230 (N_2230,N_1953,N_1855);
nor U2231 (N_2231,N_1793,N_1929);
or U2232 (N_2232,N_1879,N_1824);
nand U2233 (N_2233,N_1970,N_1779);
nand U2234 (N_2234,N_1800,N_1784);
or U2235 (N_2235,N_1947,N_1817);
nand U2236 (N_2236,N_1824,N_1757);
nor U2237 (N_2237,N_1807,N_1991);
nor U2238 (N_2238,N_1790,N_1870);
nand U2239 (N_2239,N_1916,N_1856);
or U2240 (N_2240,N_1910,N_1935);
xor U2241 (N_2241,N_1970,N_1881);
or U2242 (N_2242,N_1907,N_1930);
and U2243 (N_2243,N_1819,N_1752);
nor U2244 (N_2244,N_1972,N_1817);
and U2245 (N_2245,N_1759,N_1868);
and U2246 (N_2246,N_1932,N_1768);
xor U2247 (N_2247,N_1751,N_1961);
and U2248 (N_2248,N_1880,N_1926);
xor U2249 (N_2249,N_1945,N_1882);
nor U2250 (N_2250,N_2220,N_2123);
and U2251 (N_2251,N_2075,N_2108);
or U2252 (N_2252,N_2141,N_2156);
or U2253 (N_2253,N_2230,N_2159);
or U2254 (N_2254,N_2055,N_2106);
or U2255 (N_2255,N_2185,N_2048);
xnor U2256 (N_2256,N_2107,N_2078);
xor U2257 (N_2257,N_2236,N_2112);
nand U2258 (N_2258,N_2239,N_2197);
or U2259 (N_2259,N_2100,N_2158);
nor U2260 (N_2260,N_2074,N_2054);
nor U2261 (N_2261,N_2214,N_2136);
nand U2262 (N_2262,N_2202,N_2225);
xor U2263 (N_2263,N_2038,N_2067);
nand U2264 (N_2264,N_2044,N_2232);
or U2265 (N_2265,N_2000,N_2187);
or U2266 (N_2266,N_2026,N_2135);
nand U2267 (N_2267,N_2065,N_2025);
xor U2268 (N_2268,N_2188,N_2186);
xor U2269 (N_2269,N_2234,N_2138);
nand U2270 (N_2270,N_2101,N_2028);
xnor U2271 (N_2271,N_2211,N_2160);
xnor U2272 (N_2272,N_2249,N_2163);
and U2273 (N_2273,N_2098,N_2084);
and U2274 (N_2274,N_2180,N_2068);
or U2275 (N_2275,N_2010,N_2227);
xor U2276 (N_2276,N_2058,N_2210);
nand U2277 (N_2277,N_2140,N_2237);
or U2278 (N_2278,N_2009,N_2029);
nand U2279 (N_2279,N_2036,N_2208);
or U2280 (N_2280,N_2161,N_2045);
nor U2281 (N_2281,N_2189,N_2179);
nor U2282 (N_2282,N_2031,N_2064);
nand U2283 (N_2283,N_2063,N_2097);
xor U2284 (N_2284,N_2165,N_2017);
nand U2285 (N_2285,N_2032,N_2072);
nand U2286 (N_2286,N_2011,N_2228);
and U2287 (N_2287,N_2016,N_2248);
nor U2288 (N_2288,N_2217,N_2083);
or U2289 (N_2289,N_2231,N_2096);
or U2290 (N_2290,N_2233,N_2190);
nor U2291 (N_2291,N_2111,N_2221);
or U2292 (N_2292,N_2222,N_2201);
or U2293 (N_2293,N_2006,N_2018);
or U2294 (N_2294,N_2219,N_2116);
nand U2295 (N_2295,N_2071,N_2204);
or U2296 (N_2296,N_2056,N_2152);
or U2297 (N_2297,N_2093,N_2149);
nand U2298 (N_2298,N_2130,N_2240);
and U2299 (N_2299,N_2019,N_2086);
or U2300 (N_2300,N_2042,N_2057);
xor U2301 (N_2301,N_2076,N_2105);
nand U2302 (N_2302,N_2247,N_2060);
nand U2303 (N_2303,N_2126,N_2050);
xor U2304 (N_2304,N_2139,N_2131);
nor U2305 (N_2305,N_2079,N_2142);
nor U2306 (N_2306,N_2178,N_2242);
nor U2307 (N_2307,N_2162,N_2091);
xor U2308 (N_2308,N_2169,N_2226);
nor U2309 (N_2309,N_2133,N_2132);
or U2310 (N_2310,N_2114,N_2049);
xnor U2311 (N_2311,N_2113,N_2172);
xnor U2312 (N_2312,N_2085,N_2062);
nand U2313 (N_2313,N_2014,N_2200);
nor U2314 (N_2314,N_2215,N_2164);
and U2315 (N_2315,N_2207,N_2046);
xnor U2316 (N_2316,N_2059,N_2246);
nand U2317 (N_2317,N_2243,N_2127);
or U2318 (N_2318,N_2195,N_2024);
and U2319 (N_2319,N_2023,N_2039);
and U2320 (N_2320,N_2129,N_2167);
nor U2321 (N_2321,N_2216,N_2003);
nor U2322 (N_2322,N_2213,N_2244);
and U2323 (N_2323,N_2203,N_2082);
or U2324 (N_2324,N_2033,N_2088);
xnor U2325 (N_2325,N_2122,N_2103);
or U2326 (N_2326,N_2145,N_2128);
and U2327 (N_2327,N_2205,N_2007);
xnor U2328 (N_2328,N_2120,N_2144);
or U2329 (N_2329,N_2021,N_2034);
nand U2330 (N_2330,N_2040,N_2061);
or U2331 (N_2331,N_2070,N_2212);
xor U2332 (N_2332,N_2182,N_2027);
xnor U2333 (N_2333,N_2022,N_2198);
and U2334 (N_2334,N_2125,N_2193);
nor U2335 (N_2335,N_2090,N_2119);
nand U2336 (N_2336,N_2154,N_2087);
xor U2337 (N_2337,N_2109,N_2147);
and U2338 (N_2338,N_2157,N_2043);
xor U2339 (N_2339,N_2168,N_2020);
nand U2340 (N_2340,N_2191,N_2037);
or U2341 (N_2341,N_2175,N_2094);
and U2342 (N_2342,N_2148,N_2104);
nor U2343 (N_2343,N_2013,N_2238);
or U2344 (N_2344,N_2099,N_2176);
and U2345 (N_2345,N_2035,N_2173);
xnor U2346 (N_2346,N_2081,N_2012);
nand U2347 (N_2347,N_2206,N_2121);
nor U2348 (N_2348,N_2137,N_2073);
nor U2349 (N_2349,N_2015,N_2124);
nor U2350 (N_2350,N_2102,N_2218);
xnor U2351 (N_2351,N_2245,N_2199);
nor U2352 (N_2352,N_2052,N_2030);
nand U2353 (N_2353,N_2117,N_2053);
nand U2354 (N_2354,N_2066,N_2005);
xnor U2355 (N_2355,N_2241,N_2184);
nand U2356 (N_2356,N_2224,N_2155);
nand U2357 (N_2357,N_2051,N_2229);
xor U2358 (N_2358,N_2235,N_2004);
nor U2359 (N_2359,N_2181,N_2153);
nand U2360 (N_2360,N_2110,N_2209);
nor U2361 (N_2361,N_2166,N_2192);
nand U2362 (N_2362,N_2080,N_2151);
nor U2363 (N_2363,N_2047,N_2143);
nor U2364 (N_2364,N_2115,N_2170);
and U2365 (N_2365,N_2069,N_2223);
or U2366 (N_2366,N_2194,N_2092);
nand U2367 (N_2367,N_2118,N_2146);
xor U2368 (N_2368,N_2089,N_2196);
nor U2369 (N_2369,N_2177,N_2174);
nand U2370 (N_2370,N_2095,N_2002);
or U2371 (N_2371,N_2134,N_2041);
or U2372 (N_2372,N_2171,N_2183);
nand U2373 (N_2373,N_2008,N_2150);
nand U2374 (N_2374,N_2077,N_2001);
or U2375 (N_2375,N_2240,N_2021);
nor U2376 (N_2376,N_2037,N_2136);
nand U2377 (N_2377,N_2178,N_2132);
nand U2378 (N_2378,N_2182,N_2104);
xor U2379 (N_2379,N_2231,N_2184);
nand U2380 (N_2380,N_2044,N_2071);
nand U2381 (N_2381,N_2217,N_2150);
nand U2382 (N_2382,N_2167,N_2101);
xor U2383 (N_2383,N_2184,N_2238);
nor U2384 (N_2384,N_2109,N_2228);
or U2385 (N_2385,N_2019,N_2058);
nor U2386 (N_2386,N_2070,N_2143);
nand U2387 (N_2387,N_2244,N_2022);
nand U2388 (N_2388,N_2102,N_2208);
or U2389 (N_2389,N_2179,N_2147);
and U2390 (N_2390,N_2116,N_2205);
nor U2391 (N_2391,N_2148,N_2215);
xor U2392 (N_2392,N_2030,N_2018);
or U2393 (N_2393,N_2058,N_2180);
and U2394 (N_2394,N_2178,N_2060);
nor U2395 (N_2395,N_2091,N_2023);
nand U2396 (N_2396,N_2145,N_2134);
or U2397 (N_2397,N_2183,N_2135);
nand U2398 (N_2398,N_2108,N_2236);
xor U2399 (N_2399,N_2127,N_2032);
xnor U2400 (N_2400,N_2235,N_2150);
or U2401 (N_2401,N_2112,N_2053);
nor U2402 (N_2402,N_2054,N_2226);
nand U2403 (N_2403,N_2036,N_2222);
xor U2404 (N_2404,N_2247,N_2111);
and U2405 (N_2405,N_2213,N_2061);
or U2406 (N_2406,N_2218,N_2165);
or U2407 (N_2407,N_2110,N_2220);
xor U2408 (N_2408,N_2079,N_2015);
or U2409 (N_2409,N_2031,N_2099);
nand U2410 (N_2410,N_2080,N_2192);
xor U2411 (N_2411,N_2217,N_2128);
nor U2412 (N_2412,N_2227,N_2045);
nor U2413 (N_2413,N_2247,N_2005);
or U2414 (N_2414,N_2131,N_2156);
nand U2415 (N_2415,N_2237,N_2013);
xor U2416 (N_2416,N_2130,N_2055);
xor U2417 (N_2417,N_2028,N_2072);
xnor U2418 (N_2418,N_2236,N_2075);
nand U2419 (N_2419,N_2193,N_2028);
nand U2420 (N_2420,N_2086,N_2224);
nand U2421 (N_2421,N_2214,N_2026);
xor U2422 (N_2422,N_2236,N_2149);
nor U2423 (N_2423,N_2099,N_2246);
xor U2424 (N_2424,N_2214,N_2031);
nor U2425 (N_2425,N_2115,N_2058);
xnor U2426 (N_2426,N_2247,N_2168);
nand U2427 (N_2427,N_2166,N_2161);
or U2428 (N_2428,N_2048,N_2022);
nor U2429 (N_2429,N_2209,N_2136);
or U2430 (N_2430,N_2039,N_2065);
nand U2431 (N_2431,N_2125,N_2230);
or U2432 (N_2432,N_2020,N_2215);
xor U2433 (N_2433,N_2132,N_2007);
nor U2434 (N_2434,N_2173,N_2165);
xnor U2435 (N_2435,N_2056,N_2236);
xor U2436 (N_2436,N_2064,N_2117);
and U2437 (N_2437,N_2204,N_2058);
and U2438 (N_2438,N_2104,N_2062);
nand U2439 (N_2439,N_2045,N_2175);
nand U2440 (N_2440,N_2095,N_2060);
nand U2441 (N_2441,N_2209,N_2008);
and U2442 (N_2442,N_2175,N_2142);
nor U2443 (N_2443,N_2216,N_2001);
xnor U2444 (N_2444,N_2191,N_2082);
xor U2445 (N_2445,N_2082,N_2249);
and U2446 (N_2446,N_2084,N_2079);
or U2447 (N_2447,N_2077,N_2220);
nor U2448 (N_2448,N_2105,N_2225);
xor U2449 (N_2449,N_2062,N_2034);
nand U2450 (N_2450,N_2136,N_2240);
or U2451 (N_2451,N_2121,N_2069);
or U2452 (N_2452,N_2121,N_2048);
xnor U2453 (N_2453,N_2233,N_2006);
nor U2454 (N_2454,N_2220,N_2240);
nor U2455 (N_2455,N_2089,N_2014);
xnor U2456 (N_2456,N_2235,N_2099);
nand U2457 (N_2457,N_2138,N_2039);
and U2458 (N_2458,N_2027,N_2247);
nand U2459 (N_2459,N_2212,N_2175);
nand U2460 (N_2460,N_2077,N_2002);
nor U2461 (N_2461,N_2205,N_2055);
nor U2462 (N_2462,N_2089,N_2235);
or U2463 (N_2463,N_2062,N_2098);
nand U2464 (N_2464,N_2106,N_2230);
nor U2465 (N_2465,N_2219,N_2174);
or U2466 (N_2466,N_2016,N_2161);
or U2467 (N_2467,N_2248,N_2140);
nor U2468 (N_2468,N_2010,N_2079);
xor U2469 (N_2469,N_2071,N_2112);
nand U2470 (N_2470,N_2105,N_2201);
and U2471 (N_2471,N_2221,N_2134);
xor U2472 (N_2472,N_2167,N_2072);
and U2473 (N_2473,N_2160,N_2176);
xnor U2474 (N_2474,N_2114,N_2246);
or U2475 (N_2475,N_2198,N_2159);
or U2476 (N_2476,N_2021,N_2077);
nand U2477 (N_2477,N_2071,N_2003);
xor U2478 (N_2478,N_2063,N_2067);
nand U2479 (N_2479,N_2108,N_2135);
nor U2480 (N_2480,N_2228,N_2058);
or U2481 (N_2481,N_2056,N_2084);
nor U2482 (N_2482,N_2110,N_2247);
nor U2483 (N_2483,N_2096,N_2050);
or U2484 (N_2484,N_2236,N_2090);
nor U2485 (N_2485,N_2224,N_2126);
and U2486 (N_2486,N_2152,N_2065);
nor U2487 (N_2487,N_2167,N_2012);
nand U2488 (N_2488,N_2095,N_2247);
xor U2489 (N_2489,N_2057,N_2058);
xnor U2490 (N_2490,N_2092,N_2148);
nor U2491 (N_2491,N_2024,N_2065);
or U2492 (N_2492,N_2107,N_2025);
nand U2493 (N_2493,N_2187,N_2115);
and U2494 (N_2494,N_2045,N_2158);
xor U2495 (N_2495,N_2053,N_2094);
and U2496 (N_2496,N_2202,N_2246);
nand U2497 (N_2497,N_2105,N_2164);
xnor U2498 (N_2498,N_2059,N_2013);
and U2499 (N_2499,N_2130,N_2099);
or U2500 (N_2500,N_2499,N_2418);
or U2501 (N_2501,N_2262,N_2291);
and U2502 (N_2502,N_2493,N_2449);
nor U2503 (N_2503,N_2464,N_2277);
and U2504 (N_2504,N_2431,N_2375);
or U2505 (N_2505,N_2426,N_2331);
or U2506 (N_2506,N_2459,N_2402);
or U2507 (N_2507,N_2269,N_2340);
nand U2508 (N_2508,N_2396,N_2364);
nor U2509 (N_2509,N_2400,N_2303);
or U2510 (N_2510,N_2434,N_2383);
xnor U2511 (N_2511,N_2315,N_2466);
nor U2512 (N_2512,N_2322,N_2330);
and U2513 (N_2513,N_2312,N_2429);
xor U2514 (N_2514,N_2279,N_2397);
xor U2515 (N_2515,N_2296,N_2488);
or U2516 (N_2516,N_2411,N_2299);
or U2517 (N_2517,N_2327,N_2250);
and U2518 (N_2518,N_2467,N_2441);
or U2519 (N_2519,N_2274,N_2436);
nor U2520 (N_2520,N_2254,N_2425);
nor U2521 (N_2521,N_2301,N_2391);
xor U2522 (N_2522,N_2353,N_2455);
or U2523 (N_2523,N_2308,N_2275);
nor U2524 (N_2524,N_2395,N_2469);
nand U2525 (N_2525,N_2428,N_2415);
xnor U2526 (N_2526,N_2385,N_2496);
nand U2527 (N_2527,N_2332,N_2316);
and U2528 (N_2528,N_2445,N_2363);
and U2529 (N_2529,N_2284,N_2320);
or U2530 (N_2530,N_2422,N_2382);
xnor U2531 (N_2531,N_2326,N_2255);
and U2532 (N_2532,N_2410,N_2325);
xnor U2533 (N_2533,N_2306,N_2286);
nand U2534 (N_2534,N_2376,N_2440);
xor U2535 (N_2535,N_2430,N_2462);
nand U2536 (N_2536,N_2369,N_2278);
and U2537 (N_2537,N_2358,N_2361);
or U2538 (N_2538,N_2302,N_2367);
and U2539 (N_2539,N_2336,N_2309);
or U2540 (N_2540,N_2494,N_2270);
and U2541 (N_2541,N_2388,N_2341);
nand U2542 (N_2542,N_2354,N_2458);
xor U2543 (N_2543,N_2371,N_2349);
nand U2544 (N_2544,N_2453,N_2352);
nor U2545 (N_2545,N_2448,N_2264);
nand U2546 (N_2546,N_2355,N_2344);
nor U2547 (N_2547,N_2342,N_2404);
xor U2548 (N_2548,N_2319,N_2424);
nand U2549 (N_2549,N_2321,N_2486);
or U2550 (N_2550,N_2399,N_2456);
nand U2551 (N_2551,N_2350,N_2289);
nor U2552 (N_2552,N_2468,N_2446);
nand U2553 (N_2553,N_2317,N_2479);
or U2554 (N_2554,N_2283,N_2265);
and U2555 (N_2555,N_2498,N_2256);
nand U2556 (N_2556,N_2421,N_2427);
nor U2557 (N_2557,N_2282,N_2347);
or U2558 (N_2558,N_2297,N_2345);
or U2559 (N_2559,N_2474,N_2394);
xor U2560 (N_2560,N_2387,N_2314);
nor U2561 (N_2561,N_2378,N_2439);
nor U2562 (N_2562,N_2447,N_2334);
and U2563 (N_2563,N_2271,N_2360);
and U2564 (N_2564,N_2492,N_2380);
or U2565 (N_2565,N_2390,N_2491);
or U2566 (N_2566,N_2293,N_2337);
nand U2567 (N_2567,N_2379,N_2351);
and U2568 (N_2568,N_2401,N_2373);
nor U2569 (N_2569,N_2292,N_2452);
nand U2570 (N_2570,N_2346,N_2497);
or U2571 (N_2571,N_2343,N_2487);
and U2572 (N_2572,N_2423,N_2258);
or U2573 (N_2573,N_2437,N_2295);
nor U2574 (N_2574,N_2368,N_2398);
or U2575 (N_2575,N_2280,N_2267);
nor U2576 (N_2576,N_2417,N_2333);
xnor U2577 (N_2577,N_2414,N_2335);
nor U2578 (N_2578,N_2263,N_2409);
and U2579 (N_2579,N_2370,N_2362);
or U2580 (N_2580,N_2272,N_2465);
or U2581 (N_2581,N_2260,N_2457);
or U2582 (N_2582,N_2359,N_2298);
or U2583 (N_2583,N_2253,N_2485);
and U2584 (N_2584,N_2480,N_2338);
xnor U2585 (N_2585,N_2393,N_2287);
xnor U2586 (N_2586,N_2266,N_2389);
or U2587 (N_2587,N_2419,N_2290);
or U2588 (N_2588,N_2490,N_2416);
nand U2589 (N_2589,N_2386,N_2470);
xor U2590 (N_2590,N_2281,N_2433);
and U2591 (N_2591,N_2377,N_2307);
or U2592 (N_2592,N_2481,N_2285);
nor U2593 (N_2593,N_2460,N_2420);
xor U2594 (N_2594,N_2311,N_2261);
nor U2595 (N_2595,N_2366,N_2450);
xor U2596 (N_2596,N_2339,N_2372);
xor U2597 (N_2597,N_2288,N_2454);
and U2598 (N_2598,N_2305,N_2259);
and U2599 (N_2599,N_2324,N_2471);
xor U2600 (N_2600,N_2356,N_2412);
xor U2601 (N_2601,N_2252,N_2257);
nor U2602 (N_2602,N_2408,N_2473);
nand U2603 (N_2603,N_2329,N_2268);
nand U2604 (N_2604,N_2444,N_2304);
xor U2605 (N_2605,N_2357,N_2328);
and U2606 (N_2606,N_2461,N_2482);
nand U2607 (N_2607,N_2384,N_2276);
nand U2608 (N_2608,N_2413,N_2374);
nand U2609 (N_2609,N_2477,N_2407);
nor U2610 (N_2610,N_2478,N_2310);
or U2611 (N_2611,N_2484,N_2318);
nor U2612 (N_2612,N_2435,N_2463);
nand U2613 (N_2613,N_2300,N_2443);
and U2614 (N_2614,N_2438,N_2251);
nand U2615 (N_2615,N_2403,N_2432);
xnor U2616 (N_2616,N_2442,N_2348);
nand U2617 (N_2617,N_2472,N_2294);
xnor U2618 (N_2618,N_2381,N_2476);
or U2619 (N_2619,N_2392,N_2483);
nand U2620 (N_2620,N_2495,N_2365);
nor U2621 (N_2621,N_2405,N_2273);
and U2622 (N_2622,N_2475,N_2406);
nand U2623 (N_2623,N_2489,N_2451);
xnor U2624 (N_2624,N_2323,N_2313);
xnor U2625 (N_2625,N_2358,N_2274);
or U2626 (N_2626,N_2467,N_2452);
nand U2627 (N_2627,N_2473,N_2447);
nand U2628 (N_2628,N_2419,N_2459);
nand U2629 (N_2629,N_2367,N_2271);
nand U2630 (N_2630,N_2397,N_2291);
xnor U2631 (N_2631,N_2353,N_2421);
and U2632 (N_2632,N_2466,N_2286);
nor U2633 (N_2633,N_2375,N_2412);
or U2634 (N_2634,N_2391,N_2444);
nor U2635 (N_2635,N_2331,N_2316);
or U2636 (N_2636,N_2350,N_2340);
xor U2637 (N_2637,N_2315,N_2327);
and U2638 (N_2638,N_2329,N_2328);
or U2639 (N_2639,N_2456,N_2345);
and U2640 (N_2640,N_2254,N_2278);
nand U2641 (N_2641,N_2347,N_2358);
nor U2642 (N_2642,N_2390,N_2401);
or U2643 (N_2643,N_2464,N_2278);
nor U2644 (N_2644,N_2335,N_2332);
or U2645 (N_2645,N_2346,N_2349);
xor U2646 (N_2646,N_2309,N_2339);
or U2647 (N_2647,N_2420,N_2456);
nand U2648 (N_2648,N_2439,N_2450);
nor U2649 (N_2649,N_2392,N_2251);
nor U2650 (N_2650,N_2289,N_2473);
xnor U2651 (N_2651,N_2359,N_2362);
or U2652 (N_2652,N_2297,N_2253);
xor U2653 (N_2653,N_2393,N_2442);
nor U2654 (N_2654,N_2372,N_2258);
or U2655 (N_2655,N_2275,N_2285);
and U2656 (N_2656,N_2397,N_2461);
nand U2657 (N_2657,N_2413,N_2376);
and U2658 (N_2658,N_2291,N_2311);
xor U2659 (N_2659,N_2473,N_2430);
nand U2660 (N_2660,N_2434,N_2367);
nand U2661 (N_2661,N_2450,N_2477);
nor U2662 (N_2662,N_2267,N_2467);
xor U2663 (N_2663,N_2408,N_2328);
nand U2664 (N_2664,N_2463,N_2452);
and U2665 (N_2665,N_2478,N_2314);
nand U2666 (N_2666,N_2330,N_2258);
nor U2667 (N_2667,N_2384,N_2440);
nand U2668 (N_2668,N_2388,N_2464);
xnor U2669 (N_2669,N_2306,N_2258);
nor U2670 (N_2670,N_2437,N_2405);
xnor U2671 (N_2671,N_2286,N_2427);
or U2672 (N_2672,N_2381,N_2497);
nand U2673 (N_2673,N_2331,N_2485);
xnor U2674 (N_2674,N_2460,N_2407);
and U2675 (N_2675,N_2379,N_2415);
nor U2676 (N_2676,N_2473,N_2424);
nor U2677 (N_2677,N_2373,N_2316);
and U2678 (N_2678,N_2284,N_2488);
xor U2679 (N_2679,N_2428,N_2453);
or U2680 (N_2680,N_2349,N_2334);
or U2681 (N_2681,N_2469,N_2464);
xor U2682 (N_2682,N_2306,N_2458);
nor U2683 (N_2683,N_2447,N_2421);
nand U2684 (N_2684,N_2362,N_2461);
nor U2685 (N_2685,N_2267,N_2380);
and U2686 (N_2686,N_2362,N_2293);
nand U2687 (N_2687,N_2456,N_2395);
and U2688 (N_2688,N_2254,N_2410);
and U2689 (N_2689,N_2348,N_2359);
nand U2690 (N_2690,N_2290,N_2415);
or U2691 (N_2691,N_2343,N_2388);
xor U2692 (N_2692,N_2378,N_2252);
nand U2693 (N_2693,N_2467,N_2361);
xor U2694 (N_2694,N_2415,N_2375);
and U2695 (N_2695,N_2348,N_2376);
nand U2696 (N_2696,N_2485,N_2352);
xor U2697 (N_2697,N_2332,N_2382);
nand U2698 (N_2698,N_2478,N_2437);
xnor U2699 (N_2699,N_2478,N_2459);
and U2700 (N_2700,N_2333,N_2481);
nor U2701 (N_2701,N_2326,N_2353);
xor U2702 (N_2702,N_2270,N_2264);
and U2703 (N_2703,N_2376,N_2459);
nand U2704 (N_2704,N_2448,N_2257);
nor U2705 (N_2705,N_2316,N_2256);
or U2706 (N_2706,N_2263,N_2359);
and U2707 (N_2707,N_2340,N_2341);
xnor U2708 (N_2708,N_2452,N_2277);
or U2709 (N_2709,N_2413,N_2414);
nor U2710 (N_2710,N_2308,N_2470);
nor U2711 (N_2711,N_2291,N_2419);
xor U2712 (N_2712,N_2469,N_2286);
or U2713 (N_2713,N_2455,N_2309);
nor U2714 (N_2714,N_2306,N_2344);
nand U2715 (N_2715,N_2371,N_2391);
nand U2716 (N_2716,N_2292,N_2325);
or U2717 (N_2717,N_2402,N_2315);
nor U2718 (N_2718,N_2304,N_2419);
xor U2719 (N_2719,N_2380,N_2260);
nor U2720 (N_2720,N_2359,N_2424);
or U2721 (N_2721,N_2314,N_2294);
xor U2722 (N_2722,N_2361,N_2436);
xnor U2723 (N_2723,N_2403,N_2399);
xnor U2724 (N_2724,N_2271,N_2426);
or U2725 (N_2725,N_2311,N_2320);
and U2726 (N_2726,N_2291,N_2321);
xnor U2727 (N_2727,N_2376,N_2456);
nand U2728 (N_2728,N_2437,N_2292);
or U2729 (N_2729,N_2437,N_2262);
and U2730 (N_2730,N_2463,N_2257);
nor U2731 (N_2731,N_2397,N_2329);
and U2732 (N_2732,N_2361,N_2414);
or U2733 (N_2733,N_2309,N_2468);
nor U2734 (N_2734,N_2368,N_2288);
nand U2735 (N_2735,N_2470,N_2494);
nand U2736 (N_2736,N_2361,N_2338);
nand U2737 (N_2737,N_2471,N_2451);
and U2738 (N_2738,N_2254,N_2400);
nand U2739 (N_2739,N_2258,N_2400);
or U2740 (N_2740,N_2390,N_2315);
nand U2741 (N_2741,N_2432,N_2404);
xnor U2742 (N_2742,N_2469,N_2428);
xor U2743 (N_2743,N_2404,N_2454);
or U2744 (N_2744,N_2442,N_2434);
or U2745 (N_2745,N_2279,N_2333);
and U2746 (N_2746,N_2488,N_2279);
nor U2747 (N_2747,N_2413,N_2379);
xnor U2748 (N_2748,N_2428,N_2394);
xor U2749 (N_2749,N_2302,N_2499);
and U2750 (N_2750,N_2701,N_2587);
nand U2751 (N_2751,N_2550,N_2574);
nand U2752 (N_2752,N_2710,N_2500);
nand U2753 (N_2753,N_2504,N_2563);
or U2754 (N_2754,N_2729,N_2654);
xnor U2755 (N_2755,N_2501,N_2619);
nor U2756 (N_2756,N_2552,N_2513);
nand U2757 (N_2757,N_2585,N_2560);
and U2758 (N_2758,N_2644,N_2532);
and U2759 (N_2759,N_2695,N_2690);
nor U2760 (N_2760,N_2601,N_2604);
nor U2761 (N_2761,N_2618,N_2684);
xnor U2762 (N_2762,N_2613,N_2638);
or U2763 (N_2763,N_2542,N_2674);
nand U2764 (N_2764,N_2609,N_2508);
or U2765 (N_2765,N_2687,N_2657);
nor U2766 (N_2766,N_2555,N_2553);
xor U2767 (N_2767,N_2645,N_2537);
nand U2768 (N_2768,N_2575,N_2625);
or U2769 (N_2769,N_2681,N_2743);
nand U2770 (N_2770,N_2540,N_2721);
and U2771 (N_2771,N_2534,N_2716);
xnor U2772 (N_2772,N_2636,N_2610);
nor U2773 (N_2773,N_2667,N_2635);
nor U2774 (N_2774,N_2698,N_2649);
nor U2775 (N_2775,N_2682,N_2707);
nor U2776 (N_2776,N_2745,N_2642);
nor U2777 (N_2777,N_2567,N_2617);
xnor U2778 (N_2778,N_2620,N_2577);
xnor U2779 (N_2779,N_2713,N_2648);
or U2780 (N_2780,N_2573,N_2626);
nand U2781 (N_2781,N_2502,N_2584);
and U2782 (N_2782,N_2562,N_2686);
xnor U2783 (N_2783,N_2680,N_2715);
nor U2784 (N_2784,N_2709,N_2679);
or U2785 (N_2785,N_2530,N_2544);
nand U2786 (N_2786,N_2509,N_2748);
or U2787 (N_2787,N_2668,N_2669);
xor U2788 (N_2788,N_2590,N_2592);
and U2789 (N_2789,N_2518,N_2526);
and U2790 (N_2790,N_2511,N_2639);
xor U2791 (N_2791,N_2536,N_2708);
nand U2792 (N_2792,N_2566,N_2616);
or U2793 (N_2793,N_2510,N_2559);
xor U2794 (N_2794,N_2597,N_2699);
nand U2795 (N_2795,N_2614,N_2593);
nand U2796 (N_2796,N_2515,N_2608);
nor U2797 (N_2797,N_2529,N_2576);
nand U2798 (N_2798,N_2637,N_2655);
nor U2799 (N_2799,N_2704,N_2664);
and U2800 (N_2800,N_2611,N_2746);
and U2801 (N_2801,N_2623,N_2653);
xor U2802 (N_2802,N_2683,N_2548);
nand U2803 (N_2803,N_2725,N_2742);
or U2804 (N_2804,N_2523,N_2651);
and U2805 (N_2805,N_2615,N_2561);
or U2806 (N_2806,N_2506,N_2737);
xnor U2807 (N_2807,N_2572,N_2722);
xor U2808 (N_2808,N_2514,N_2528);
and U2809 (N_2809,N_2632,N_2557);
nor U2810 (N_2810,N_2538,N_2724);
nand U2811 (N_2811,N_2723,N_2622);
or U2812 (N_2812,N_2665,N_2578);
or U2813 (N_2813,N_2527,N_2565);
nand U2814 (N_2814,N_2607,N_2582);
and U2815 (N_2815,N_2652,N_2594);
and U2816 (N_2816,N_2519,N_2627);
and U2817 (N_2817,N_2505,N_2630);
xor U2818 (N_2818,N_2606,N_2634);
or U2819 (N_2819,N_2586,N_2705);
nor U2820 (N_2820,N_2629,N_2672);
xor U2821 (N_2821,N_2740,N_2663);
or U2822 (N_2822,N_2579,N_2558);
and U2823 (N_2823,N_2659,N_2605);
nor U2824 (N_2824,N_2547,N_2738);
nand U2825 (N_2825,N_2749,N_2551);
nor U2826 (N_2826,N_2733,N_2744);
nor U2827 (N_2827,N_2660,N_2533);
nand U2828 (N_2828,N_2688,N_2666);
xnor U2829 (N_2829,N_2647,N_2556);
or U2830 (N_2830,N_2641,N_2658);
nand U2831 (N_2831,N_2735,N_2673);
and U2832 (N_2832,N_2522,N_2524);
or U2833 (N_2833,N_2546,N_2697);
nand U2834 (N_2834,N_2650,N_2675);
nor U2835 (N_2835,N_2711,N_2646);
and U2836 (N_2836,N_2696,N_2568);
xor U2837 (N_2837,N_2661,N_2512);
or U2838 (N_2838,N_2599,N_2718);
and U2839 (N_2839,N_2719,N_2685);
nor U2840 (N_2840,N_2693,N_2640);
nor U2841 (N_2841,N_2612,N_2734);
nand U2842 (N_2842,N_2570,N_2535);
and U2843 (N_2843,N_2588,N_2631);
xnor U2844 (N_2844,N_2581,N_2677);
nor U2845 (N_2845,N_2662,N_2521);
or U2846 (N_2846,N_2621,N_2569);
and U2847 (N_2847,N_2595,N_2706);
and U2848 (N_2848,N_2516,N_2525);
and U2849 (N_2849,N_2712,N_2730);
nand U2850 (N_2850,N_2739,N_2580);
and U2851 (N_2851,N_2507,N_2717);
nor U2852 (N_2852,N_2728,N_2602);
xnor U2853 (N_2853,N_2600,N_2549);
nand U2854 (N_2854,N_2656,N_2596);
nor U2855 (N_2855,N_2517,N_2694);
nor U2856 (N_2856,N_2589,N_2624);
nand U2857 (N_2857,N_2678,N_2628);
xnor U2858 (N_2858,N_2503,N_2692);
and U2859 (N_2859,N_2700,N_2539);
xor U2860 (N_2860,N_2736,N_2747);
xnor U2861 (N_2861,N_2531,N_2591);
nand U2862 (N_2862,N_2741,N_2714);
xor U2863 (N_2863,N_2676,N_2726);
nor U2864 (N_2864,N_2720,N_2643);
or U2865 (N_2865,N_2541,N_2520);
and U2866 (N_2866,N_2731,N_2633);
and U2867 (N_2867,N_2554,N_2689);
or U2868 (N_2868,N_2703,N_2727);
nor U2869 (N_2869,N_2583,N_2564);
nand U2870 (N_2870,N_2598,N_2545);
nand U2871 (N_2871,N_2671,N_2702);
xnor U2872 (N_2872,N_2571,N_2543);
and U2873 (N_2873,N_2670,N_2732);
and U2874 (N_2874,N_2691,N_2603);
nand U2875 (N_2875,N_2565,N_2667);
nand U2876 (N_2876,N_2620,N_2648);
xor U2877 (N_2877,N_2591,N_2519);
or U2878 (N_2878,N_2584,N_2731);
or U2879 (N_2879,N_2627,N_2708);
and U2880 (N_2880,N_2728,N_2584);
and U2881 (N_2881,N_2688,N_2709);
or U2882 (N_2882,N_2696,N_2629);
and U2883 (N_2883,N_2608,N_2545);
xnor U2884 (N_2884,N_2601,N_2733);
nand U2885 (N_2885,N_2687,N_2644);
xnor U2886 (N_2886,N_2510,N_2684);
xnor U2887 (N_2887,N_2521,N_2627);
nand U2888 (N_2888,N_2580,N_2558);
nor U2889 (N_2889,N_2738,N_2576);
or U2890 (N_2890,N_2743,N_2646);
nand U2891 (N_2891,N_2641,N_2560);
nand U2892 (N_2892,N_2500,N_2713);
nand U2893 (N_2893,N_2544,N_2716);
nand U2894 (N_2894,N_2607,N_2520);
xnor U2895 (N_2895,N_2610,N_2541);
or U2896 (N_2896,N_2510,N_2708);
nor U2897 (N_2897,N_2561,N_2654);
and U2898 (N_2898,N_2742,N_2612);
and U2899 (N_2899,N_2599,N_2669);
nor U2900 (N_2900,N_2560,N_2568);
nor U2901 (N_2901,N_2632,N_2568);
nand U2902 (N_2902,N_2520,N_2650);
and U2903 (N_2903,N_2508,N_2736);
nand U2904 (N_2904,N_2627,N_2617);
xor U2905 (N_2905,N_2727,N_2581);
xor U2906 (N_2906,N_2706,N_2633);
nor U2907 (N_2907,N_2582,N_2615);
or U2908 (N_2908,N_2553,N_2632);
or U2909 (N_2909,N_2614,N_2527);
nand U2910 (N_2910,N_2691,N_2508);
nor U2911 (N_2911,N_2666,N_2680);
and U2912 (N_2912,N_2599,N_2526);
and U2913 (N_2913,N_2628,N_2505);
and U2914 (N_2914,N_2743,N_2610);
nor U2915 (N_2915,N_2675,N_2720);
and U2916 (N_2916,N_2622,N_2640);
or U2917 (N_2917,N_2681,N_2732);
or U2918 (N_2918,N_2530,N_2694);
nor U2919 (N_2919,N_2689,N_2716);
nand U2920 (N_2920,N_2613,N_2573);
and U2921 (N_2921,N_2718,N_2550);
and U2922 (N_2922,N_2549,N_2656);
xor U2923 (N_2923,N_2663,N_2670);
nand U2924 (N_2924,N_2692,N_2509);
xnor U2925 (N_2925,N_2553,N_2683);
and U2926 (N_2926,N_2626,N_2547);
or U2927 (N_2927,N_2549,N_2513);
nor U2928 (N_2928,N_2710,N_2655);
xnor U2929 (N_2929,N_2634,N_2569);
or U2930 (N_2930,N_2512,N_2505);
nor U2931 (N_2931,N_2576,N_2562);
nand U2932 (N_2932,N_2545,N_2701);
and U2933 (N_2933,N_2669,N_2712);
nand U2934 (N_2934,N_2515,N_2502);
or U2935 (N_2935,N_2699,N_2614);
nor U2936 (N_2936,N_2707,N_2696);
nor U2937 (N_2937,N_2744,N_2572);
and U2938 (N_2938,N_2506,N_2708);
or U2939 (N_2939,N_2611,N_2579);
or U2940 (N_2940,N_2636,N_2665);
xor U2941 (N_2941,N_2556,N_2718);
nor U2942 (N_2942,N_2520,N_2575);
and U2943 (N_2943,N_2601,N_2700);
nor U2944 (N_2944,N_2703,N_2656);
nor U2945 (N_2945,N_2535,N_2522);
nand U2946 (N_2946,N_2531,N_2654);
and U2947 (N_2947,N_2640,N_2558);
and U2948 (N_2948,N_2617,N_2655);
xor U2949 (N_2949,N_2561,N_2517);
nand U2950 (N_2950,N_2664,N_2689);
nand U2951 (N_2951,N_2694,N_2535);
xor U2952 (N_2952,N_2706,N_2695);
nor U2953 (N_2953,N_2663,N_2619);
and U2954 (N_2954,N_2639,N_2603);
nand U2955 (N_2955,N_2652,N_2688);
nor U2956 (N_2956,N_2531,N_2610);
nor U2957 (N_2957,N_2707,N_2727);
and U2958 (N_2958,N_2513,N_2527);
and U2959 (N_2959,N_2682,N_2695);
xnor U2960 (N_2960,N_2731,N_2741);
xor U2961 (N_2961,N_2739,N_2689);
or U2962 (N_2962,N_2529,N_2655);
nand U2963 (N_2963,N_2665,N_2508);
xnor U2964 (N_2964,N_2650,N_2546);
xnor U2965 (N_2965,N_2543,N_2596);
nand U2966 (N_2966,N_2586,N_2588);
nor U2967 (N_2967,N_2724,N_2663);
xnor U2968 (N_2968,N_2650,N_2513);
or U2969 (N_2969,N_2603,N_2514);
xor U2970 (N_2970,N_2678,N_2610);
and U2971 (N_2971,N_2555,N_2676);
nand U2972 (N_2972,N_2722,N_2614);
nor U2973 (N_2973,N_2534,N_2607);
or U2974 (N_2974,N_2589,N_2725);
xor U2975 (N_2975,N_2517,N_2650);
or U2976 (N_2976,N_2616,N_2697);
nand U2977 (N_2977,N_2736,N_2659);
nand U2978 (N_2978,N_2530,N_2571);
nor U2979 (N_2979,N_2634,N_2684);
nand U2980 (N_2980,N_2584,N_2656);
xor U2981 (N_2981,N_2656,N_2557);
or U2982 (N_2982,N_2542,N_2521);
or U2983 (N_2983,N_2717,N_2600);
nor U2984 (N_2984,N_2669,N_2649);
nand U2985 (N_2985,N_2501,N_2551);
xor U2986 (N_2986,N_2677,N_2651);
nand U2987 (N_2987,N_2562,N_2568);
nand U2988 (N_2988,N_2592,N_2584);
nand U2989 (N_2989,N_2523,N_2666);
nor U2990 (N_2990,N_2720,N_2581);
nand U2991 (N_2991,N_2551,N_2694);
and U2992 (N_2992,N_2698,N_2543);
and U2993 (N_2993,N_2701,N_2568);
or U2994 (N_2994,N_2748,N_2584);
xnor U2995 (N_2995,N_2538,N_2522);
nand U2996 (N_2996,N_2650,N_2598);
or U2997 (N_2997,N_2690,N_2646);
and U2998 (N_2998,N_2503,N_2538);
and U2999 (N_2999,N_2721,N_2617);
xor U3000 (N_3000,N_2837,N_2997);
and U3001 (N_3001,N_2941,N_2762);
xnor U3002 (N_3002,N_2964,N_2999);
nand U3003 (N_3003,N_2927,N_2899);
nand U3004 (N_3004,N_2971,N_2800);
or U3005 (N_3005,N_2777,N_2751);
nor U3006 (N_3006,N_2968,N_2926);
and U3007 (N_3007,N_2853,N_2816);
nand U3008 (N_3008,N_2988,N_2907);
or U3009 (N_3009,N_2895,N_2896);
nor U3010 (N_3010,N_2804,N_2921);
and U3011 (N_3011,N_2809,N_2801);
or U3012 (N_3012,N_2924,N_2965);
xnor U3013 (N_3013,N_2756,N_2753);
or U3014 (N_3014,N_2769,N_2948);
nor U3015 (N_3015,N_2981,N_2785);
xor U3016 (N_3016,N_2799,N_2871);
nor U3017 (N_3017,N_2985,N_2780);
or U3018 (N_3018,N_2934,N_2974);
and U3019 (N_3019,N_2930,N_2977);
and U3020 (N_3020,N_2940,N_2812);
and U3021 (N_3021,N_2850,N_2912);
nand U3022 (N_3022,N_2923,N_2944);
or U3023 (N_3023,N_2834,N_2916);
nand U3024 (N_3024,N_2998,N_2768);
and U3025 (N_3025,N_2945,N_2910);
and U3026 (N_3026,N_2958,N_2818);
and U3027 (N_3027,N_2943,N_2770);
nand U3028 (N_3028,N_2849,N_2771);
nand U3029 (N_3029,N_2833,N_2806);
or U3030 (N_3030,N_2906,N_2752);
nor U3031 (N_3031,N_2903,N_2931);
nand U3032 (N_3032,N_2932,N_2784);
nand U3033 (N_3033,N_2877,N_2802);
or U3034 (N_3034,N_2873,N_2959);
xor U3035 (N_3035,N_2897,N_2901);
and U3036 (N_3036,N_2778,N_2767);
or U3037 (N_3037,N_2790,N_2986);
and U3038 (N_3038,N_2920,N_2811);
and U3039 (N_3039,N_2946,N_2835);
and U3040 (N_3040,N_2893,N_2962);
or U3041 (N_3041,N_2840,N_2775);
or U3042 (N_3042,N_2817,N_2982);
and U3043 (N_3043,N_2922,N_2861);
nand U3044 (N_3044,N_2911,N_2908);
and U3045 (N_3045,N_2844,N_2969);
or U3046 (N_3046,N_2819,N_2983);
xnor U3047 (N_3047,N_2894,N_2975);
or U3048 (N_3048,N_2876,N_2832);
xnor U3049 (N_3049,N_2807,N_2867);
and U3050 (N_3050,N_2776,N_2954);
or U3051 (N_3051,N_2956,N_2938);
and U3052 (N_3052,N_2992,N_2848);
nor U3053 (N_3053,N_2760,N_2782);
nand U3054 (N_3054,N_2774,N_2866);
xor U3055 (N_3055,N_2796,N_2973);
xor U3056 (N_3056,N_2781,N_2763);
nand U3057 (N_3057,N_2966,N_2822);
xor U3058 (N_3058,N_2862,N_2885);
nor U3059 (N_3059,N_2839,N_2815);
nand U3060 (N_3060,N_2947,N_2886);
xnor U3061 (N_3061,N_2805,N_2783);
xnor U3062 (N_3062,N_2836,N_2808);
and U3063 (N_3063,N_2798,N_2949);
nor U3064 (N_3064,N_2995,N_2915);
or U3065 (N_3065,N_2792,N_2918);
nand U3066 (N_3066,N_2847,N_2789);
nor U3067 (N_3067,N_2870,N_2810);
or U3068 (N_3068,N_2996,N_2820);
and U3069 (N_3069,N_2972,N_2905);
and U3070 (N_3070,N_2976,N_2856);
nand U3071 (N_3071,N_2786,N_2857);
or U3072 (N_3072,N_2821,N_2991);
nand U3073 (N_3073,N_2765,N_2846);
and U3074 (N_3074,N_2904,N_2967);
or U3075 (N_3075,N_2935,N_2826);
or U3076 (N_3076,N_2990,N_2859);
and U3077 (N_3077,N_2779,N_2900);
and U3078 (N_3078,N_2793,N_2953);
and U3079 (N_3079,N_2872,N_2970);
nand U3080 (N_3080,N_2825,N_2845);
nor U3081 (N_3081,N_2838,N_2961);
and U3082 (N_3082,N_2960,N_2855);
or U3083 (N_3083,N_2913,N_2890);
or U3084 (N_3084,N_2978,N_2902);
nand U3085 (N_3085,N_2863,N_2797);
xnor U3086 (N_3086,N_2984,N_2841);
nand U3087 (N_3087,N_2917,N_2858);
nor U3088 (N_3088,N_2889,N_2980);
nand U3089 (N_3089,N_2898,N_2879);
or U3090 (N_3090,N_2880,N_2942);
nand U3091 (N_3091,N_2757,N_2824);
xnor U3092 (N_3092,N_2925,N_2761);
nand U3093 (N_3093,N_2878,N_2754);
and U3094 (N_3094,N_2952,N_2773);
nand U3095 (N_3095,N_2830,N_2887);
or U3096 (N_3096,N_2955,N_2979);
nand U3097 (N_3097,N_2869,N_2892);
and U3098 (N_3098,N_2759,N_2831);
xor U3099 (N_3099,N_2865,N_2909);
nand U3100 (N_3100,N_2951,N_2884);
and U3101 (N_3101,N_2827,N_2957);
or U3102 (N_3102,N_2928,N_2766);
and U3103 (N_3103,N_2993,N_2852);
nand U3104 (N_3104,N_2888,N_2791);
xor U3105 (N_3105,N_2755,N_2854);
xor U3106 (N_3106,N_2914,N_2764);
nand U3107 (N_3107,N_2963,N_2874);
nor U3108 (N_3108,N_2843,N_2803);
nor U3109 (N_3109,N_2750,N_2794);
or U3110 (N_3110,N_2919,N_2875);
or U3111 (N_3111,N_2772,N_2823);
xor U3112 (N_3112,N_2795,N_2829);
and U3113 (N_3113,N_2989,N_2881);
or U3114 (N_3114,N_2851,N_2987);
nand U3115 (N_3115,N_2828,N_2864);
or U3116 (N_3116,N_2758,N_2842);
nand U3117 (N_3117,N_2787,N_2891);
nor U3118 (N_3118,N_2813,N_2933);
nand U3119 (N_3119,N_2883,N_2936);
nor U3120 (N_3120,N_2788,N_2937);
xor U3121 (N_3121,N_2814,N_2994);
xnor U3122 (N_3122,N_2882,N_2929);
or U3123 (N_3123,N_2868,N_2860);
nand U3124 (N_3124,N_2950,N_2939);
and U3125 (N_3125,N_2753,N_2850);
xnor U3126 (N_3126,N_2797,N_2753);
nand U3127 (N_3127,N_2909,N_2960);
or U3128 (N_3128,N_2926,N_2952);
nand U3129 (N_3129,N_2858,N_2803);
xnor U3130 (N_3130,N_2754,N_2778);
xor U3131 (N_3131,N_2787,N_2800);
and U3132 (N_3132,N_2791,N_2804);
xor U3133 (N_3133,N_2855,N_2785);
nand U3134 (N_3134,N_2823,N_2911);
nand U3135 (N_3135,N_2811,N_2830);
nand U3136 (N_3136,N_2932,N_2869);
nor U3137 (N_3137,N_2831,N_2811);
nand U3138 (N_3138,N_2905,N_2820);
nand U3139 (N_3139,N_2822,N_2974);
xnor U3140 (N_3140,N_2860,N_2904);
nand U3141 (N_3141,N_2931,N_2759);
xnor U3142 (N_3142,N_2940,N_2992);
nand U3143 (N_3143,N_2829,N_2837);
xnor U3144 (N_3144,N_2847,N_2864);
or U3145 (N_3145,N_2905,N_2982);
or U3146 (N_3146,N_2760,N_2830);
and U3147 (N_3147,N_2757,N_2892);
xnor U3148 (N_3148,N_2863,N_2834);
nor U3149 (N_3149,N_2817,N_2810);
nand U3150 (N_3150,N_2757,N_2924);
xnor U3151 (N_3151,N_2917,N_2755);
or U3152 (N_3152,N_2936,N_2955);
and U3153 (N_3153,N_2878,N_2967);
xnor U3154 (N_3154,N_2804,N_2875);
xnor U3155 (N_3155,N_2765,N_2899);
nand U3156 (N_3156,N_2809,N_2844);
or U3157 (N_3157,N_2950,N_2989);
nor U3158 (N_3158,N_2877,N_2820);
or U3159 (N_3159,N_2991,N_2868);
xor U3160 (N_3160,N_2897,N_2958);
nor U3161 (N_3161,N_2856,N_2950);
nand U3162 (N_3162,N_2957,N_2945);
nand U3163 (N_3163,N_2915,N_2992);
xnor U3164 (N_3164,N_2928,N_2935);
or U3165 (N_3165,N_2807,N_2774);
and U3166 (N_3166,N_2839,N_2837);
nor U3167 (N_3167,N_2939,N_2826);
or U3168 (N_3168,N_2827,N_2843);
and U3169 (N_3169,N_2906,N_2768);
nor U3170 (N_3170,N_2940,N_2912);
nand U3171 (N_3171,N_2847,N_2751);
or U3172 (N_3172,N_2976,N_2938);
nor U3173 (N_3173,N_2866,N_2980);
and U3174 (N_3174,N_2993,N_2889);
and U3175 (N_3175,N_2847,N_2809);
nand U3176 (N_3176,N_2938,N_2793);
xnor U3177 (N_3177,N_2950,N_2958);
and U3178 (N_3178,N_2968,N_2841);
and U3179 (N_3179,N_2892,N_2996);
xnor U3180 (N_3180,N_2975,N_2966);
xnor U3181 (N_3181,N_2959,N_2958);
and U3182 (N_3182,N_2974,N_2894);
xor U3183 (N_3183,N_2855,N_2954);
and U3184 (N_3184,N_2814,N_2928);
and U3185 (N_3185,N_2777,N_2954);
and U3186 (N_3186,N_2860,N_2776);
and U3187 (N_3187,N_2756,N_2759);
nand U3188 (N_3188,N_2923,N_2895);
or U3189 (N_3189,N_2982,N_2838);
nand U3190 (N_3190,N_2849,N_2932);
and U3191 (N_3191,N_2948,N_2872);
xnor U3192 (N_3192,N_2937,N_2958);
nor U3193 (N_3193,N_2939,N_2862);
xor U3194 (N_3194,N_2977,N_2761);
xor U3195 (N_3195,N_2995,N_2910);
and U3196 (N_3196,N_2869,N_2789);
and U3197 (N_3197,N_2857,N_2941);
xnor U3198 (N_3198,N_2786,N_2782);
and U3199 (N_3199,N_2842,N_2989);
and U3200 (N_3200,N_2850,N_2757);
or U3201 (N_3201,N_2800,N_2991);
or U3202 (N_3202,N_2917,N_2948);
or U3203 (N_3203,N_2968,N_2850);
or U3204 (N_3204,N_2955,N_2829);
nor U3205 (N_3205,N_2791,N_2851);
nand U3206 (N_3206,N_2933,N_2815);
nor U3207 (N_3207,N_2806,N_2990);
nand U3208 (N_3208,N_2912,N_2771);
xor U3209 (N_3209,N_2853,N_2773);
or U3210 (N_3210,N_2951,N_2797);
and U3211 (N_3211,N_2811,N_2942);
or U3212 (N_3212,N_2871,N_2996);
or U3213 (N_3213,N_2852,N_2907);
xor U3214 (N_3214,N_2809,N_2852);
nor U3215 (N_3215,N_2858,N_2789);
nand U3216 (N_3216,N_2871,N_2767);
xnor U3217 (N_3217,N_2946,N_2766);
or U3218 (N_3218,N_2886,N_2988);
and U3219 (N_3219,N_2858,N_2883);
and U3220 (N_3220,N_2851,N_2844);
nor U3221 (N_3221,N_2759,N_2877);
xor U3222 (N_3222,N_2977,N_2990);
nand U3223 (N_3223,N_2891,N_2962);
nand U3224 (N_3224,N_2851,N_2948);
or U3225 (N_3225,N_2765,N_2818);
nor U3226 (N_3226,N_2965,N_2828);
nand U3227 (N_3227,N_2903,N_2786);
nor U3228 (N_3228,N_2962,N_2902);
or U3229 (N_3229,N_2823,N_2794);
nor U3230 (N_3230,N_2847,N_2994);
xnor U3231 (N_3231,N_2838,N_2753);
xor U3232 (N_3232,N_2860,N_2978);
nor U3233 (N_3233,N_2818,N_2831);
nand U3234 (N_3234,N_2780,N_2860);
nand U3235 (N_3235,N_2973,N_2881);
or U3236 (N_3236,N_2757,N_2805);
nand U3237 (N_3237,N_2847,N_2849);
and U3238 (N_3238,N_2919,N_2844);
nor U3239 (N_3239,N_2910,N_2872);
xnor U3240 (N_3240,N_2905,N_2758);
nand U3241 (N_3241,N_2879,N_2850);
xor U3242 (N_3242,N_2780,N_2889);
or U3243 (N_3243,N_2887,N_2950);
nor U3244 (N_3244,N_2934,N_2972);
xnor U3245 (N_3245,N_2833,N_2936);
and U3246 (N_3246,N_2815,N_2832);
xor U3247 (N_3247,N_2854,N_2800);
xor U3248 (N_3248,N_2811,N_2916);
nand U3249 (N_3249,N_2752,N_2935);
nand U3250 (N_3250,N_3193,N_3163);
and U3251 (N_3251,N_3113,N_3225);
and U3252 (N_3252,N_3122,N_3197);
xnor U3253 (N_3253,N_3043,N_3017);
and U3254 (N_3254,N_3191,N_3192);
nand U3255 (N_3255,N_3246,N_3069);
nand U3256 (N_3256,N_3233,N_3008);
or U3257 (N_3257,N_3140,N_3131);
nor U3258 (N_3258,N_3201,N_3048);
xnor U3259 (N_3259,N_3130,N_3229);
nand U3260 (N_3260,N_3180,N_3175);
nand U3261 (N_3261,N_3143,N_3165);
nor U3262 (N_3262,N_3194,N_3118);
or U3263 (N_3263,N_3188,N_3123);
and U3264 (N_3264,N_3219,N_3042);
nor U3265 (N_3265,N_3059,N_3112);
nor U3266 (N_3266,N_3038,N_3058);
xnor U3267 (N_3267,N_3023,N_3108);
nor U3268 (N_3268,N_3209,N_3154);
xor U3269 (N_3269,N_3011,N_3162);
nor U3270 (N_3270,N_3199,N_3116);
nor U3271 (N_3271,N_3203,N_3189);
nand U3272 (N_3272,N_3215,N_3115);
and U3273 (N_3273,N_3089,N_3249);
or U3274 (N_3274,N_3002,N_3213);
xnor U3275 (N_3275,N_3025,N_3155);
nor U3276 (N_3276,N_3093,N_3073);
or U3277 (N_3277,N_3110,N_3153);
nor U3278 (N_3278,N_3129,N_3171);
xnor U3279 (N_3279,N_3007,N_3047);
nor U3280 (N_3280,N_3032,N_3018);
xor U3281 (N_3281,N_3170,N_3204);
nor U3282 (N_3282,N_3234,N_3138);
nor U3283 (N_3283,N_3237,N_3056);
and U3284 (N_3284,N_3152,N_3211);
or U3285 (N_3285,N_3151,N_3183);
or U3286 (N_3286,N_3166,N_3080);
and U3287 (N_3287,N_3006,N_3092);
nor U3288 (N_3288,N_3095,N_3227);
nand U3289 (N_3289,N_3044,N_3111);
nor U3290 (N_3290,N_3055,N_3016);
nand U3291 (N_3291,N_3223,N_3075);
nand U3292 (N_3292,N_3045,N_3247);
nor U3293 (N_3293,N_3185,N_3212);
nand U3294 (N_3294,N_3026,N_3196);
xor U3295 (N_3295,N_3126,N_3035);
or U3296 (N_3296,N_3179,N_3214);
or U3297 (N_3297,N_3029,N_3109);
nor U3298 (N_3298,N_3049,N_3066);
xor U3299 (N_3299,N_3031,N_3027);
nor U3300 (N_3300,N_3172,N_3051);
xnor U3301 (N_3301,N_3005,N_3024);
and U3302 (N_3302,N_3082,N_3146);
or U3303 (N_3303,N_3070,N_3028);
nor U3304 (N_3304,N_3012,N_3034);
or U3305 (N_3305,N_3217,N_3009);
xor U3306 (N_3306,N_3160,N_3094);
nor U3307 (N_3307,N_3036,N_3063);
and U3308 (N_3308,N_3101,N_3245);
nand U3309 (N_3309,N_3173,N_3064);
nor U3310 (N_3310,N_3068,N_3085);
and U3311 (N_3311,N_3037,N_3079);
nor U3312 (N_3312,N_3087,N_3121);
or U3313 (N_3313,N_3124,N_3176);
and U3314 (N_3314,N_3142,N_3132);
nor U3315 (N_3315,N_3033,N_3205);
xnor U3316 (N_3316,N_3187,N_3039);
or U3317 (N_3317,N_3041,N_3096);
xor U3318 (N_3318,N_3167,N_3241);
nand U3319 (N_3319,N_3052,N_3100);
or U3320 (N_3320,N_3164,N_3057);
nand U3321 (N_3321,N_3014,N_3200);
nor U3322 (N_3322,N_3000,N_3090);
or U3323 (N_3323,N_3065,N_3239);
nand U3324 (N_3324,N_3020,N_3010);
and U3325 (N_3325,N_3147,N_3174);
nand U3326 (N_3326,N_3220,N_3081);
and U3327 (N_3327,N_3190,N_3083);
nand U3328 (N_3328,N_3242,N_3184);
nand U3329 (N_3329,N_3244,N_3019);
xor U3330 (N_3330,N_3248,N_3186);
nand U3331 (N_3331,N_3159,N_3243);
xor U3332 (N_3332,N_3133,N_3210);
nand U3333 (N_3333,N_3022,N_3144);
xnor U3334 (N_3334,N_3145,N_3127);
or U3335 (N_3335,N_3168,N_3054);
and U3336 (N_3336,N_3078,N_3208);
nand U3337 (N_3337,N_3084,N_3003);
and U3338 (N_3338,N_3114,N_3076);
nor U3339 (N_3339,N_3161,N_3169);
nor U3340 (N_3340,N_3021,N_3139);
and U3341 (N_3341,N_3136,N_3178);
and U3342 (N_3342,N_3013,N_3149);
or U3343 (N_3343,N_3232,N_3062);
or U3344 (N_3344,N_3119,N_3088);
or U3345 (N_3345,N_3106,N_3098);
and U3346 (N_3346,N_3207,N_3030);
and U3347 (N_3347,N_3157,N_3102);
or U3348 (N_3348,N_3202,N_3072);
or U3349 (N_3349,N_3060,N_3195);
nor U3350 (N_3350,N_3067,N_3240);
nor U3351 (N_3351,N_3099,N_3107);
nor U3352 (N_3352,N_3218,N_3150);
nor U3353 (N_3353,N_3182,N_3050);
or U3354 (N_3354,N_3226,N_3001);
xnor U3355 (N_3355,N_3074,N_3105);
and U3356 (N_3356,N_3238,N_3177);
nor U3357 (N_3357,N_3071,N_3077);
xor U3358 (N_3358,N_3148,N_3141);
nand U3359 (N_3359,N_3004,N_3120);
and U3360 (N_3360,N_3137,N_3224);
or U3361 (N_3361,N_3015,N_3086);
xnor U3362 (N_3362,N_3221,N_3104);
and U3363 (N_3363,N_3091,N_3231);
nor U3364 (N_3364,N_3230,N_3061);
xnor U3365 (N_3365,N_3128,N_3046);
or U3366 (N_3366,N_3053,N_3040);
and U3367 (N_3367,N_3103,N_3125);
nand U3368 (N_3368,N_3236,N_3156);
xor U3369 (N_3369,N_3134,N_3097);
nand U3370 (N_3370,N_3206,N_3216);
or U3371 (N_3371,N_3181,N_3235);
nand U3372 (N_3372,N_3198,N_3222);
and U3373 (N_3373,N_3158,N_3117);
xor U3374 (N_3374,N_3228,N_3135);
xor U3375 (N_3375,N_3219,N_3193);
nor U3376 (N_3376,N_3223,N_3126);
or U3377 (N_3377,N_3049,N_3246);
or U3378 (N_3378,N_3082,N_3105);
or U3379 (N_3379,N_3044,N_3053);
nand U3380 (N_3380,N_3122,N_3049);
xor U3381 (N_3381,N_3116,N_3214);
or U3382 (N_3382,N_3247,N_3024);
nand U3383 (N_3383,N_3242,N_3003);
nand U3384 (N_3384,N_3012,N_3053);
nor U3385 (N_3385,N_3126,N_3128);
and U3386 (N_3386,N_3158,N_3177);
or U3387 (N_3387,N_3061,N_3118);
nand U3388 (N_3388,N_3244,N_3012);
xor U3389 (N_3389,N_3110,N_3200);
nand U3390 (N_3390,N_3061,N_3185);
and U3391 (N_3391,N_3039,N_3010);
nand U3392 (N_3392,N_3017,N_3035);
or U3393 (N_3393,N_3024,N_3057);
or U3394 (N_3394,N_3120,N_3042);
or U3395 (N_3395,N_3042,N_3197);
and U3396 (N_3396,N_3183,N_3073);
xor U3397 (N_3397,N_3222,N_3118);
nor U3398 (N_3398,N_3100,N_3000);
nor U3399 (N_3399,N_3224,N_3044);
xor U3400 (N_3400,N_3022,N_3184);
xor U3401 (N_3401,N_3237,N_3005);
nand U3402 (N_3402,N_3144,N_3107);
nand U3403 (N_3403,N_3168,N_3141);
and U3404 (N_3404,N_3062,N_3223);
xnor U3405 (N_3405,N_3152,N_3200);
nor U3406 (N_3406,N_3132,N_3171);
nand U3407 (N_3407,N_3131,N_3212);
xor U3408 (N_3408,N_3192,N_3053);
nand U3409 (N_3409,N_3046,N_3047);
nor U3410 (N_3410,N_3158,N_3023);
and U3411 (N_3411,N_3107,N_3119);
nor U3412 (N_3412,N_3156,N_3182);
nor U3413 (N_3413,N_3002,N_3040);
xor U3414 (N_3414,N_3119,N_3098);
xnor U3415 (N_3415,N_3036,N_3120);
xnor U3416 (N_3416,N_3233,N_3121);
and U3417 (N_3417,N_3010,N_3098);
nand U3418 (N_3418,N_3096,N_3145);
nand U3419 (N_3419,N_3208,N_3031);
and U3420 (N_3420,N_3110,N_3213);
nor U3421 (N_3421,N_3215,N_3104);
or U3422 (N_3422,N_3184,N_3219);
nor U3423 (N_3423,N_3119,N_3195);
nor U3424 (N_3424,N_3002,N_3103);
nor U3425 (N_3425,N_3146,N_3032);
nor U3426 (N_3426,N_3142,N_3218);
nand U3427 (N_3427,N_3249,N_3019);
xnor U3428 (N_3428,N_3080,N_3140);
or U3429 (N_3429,N_3024,N_3124);
and U3430 (N_3430,N_3132,N_3120);
xnor U3431 (N_3431,N_3088,N_3019);
nand U3432 (N_3432,N_3151,N_3162);
nand U3433 (N_3433,N_3131,N_3137);
nand U3434 (N_3434,N_3116,N_3129);
nand U3435 (N_3435,N_3055,N_3245);
nand U3436 (N_3436,N_3118,N_3027);
or U3437 (N_3437,N_3201,N_3204);
and U3438 (N_3438,N_3109,N_3013);
or U3439 (N_3439,N_3154,N_3062);
xor U3440 (N_3440,N_3030,N_3218);
nand U3441 (N_3441,N_3035,N_3048);
nand U3442 (N_3442,N_3135,N_3030);
nor U3443 (N_3443,N_3123,N_3004);
and U3444 (N_3444,N_3223,N_3170);
nor U3445 (N_3445,N_3220,N_3067);
xnor U3446 (N_3446,N_3140,N_3132);
nor U3447 (N_3447,N_3158,N_3014);
and U3448 (N_3448,N_3041,N_3160);
or U3449 (N_3449,N_3239,N_3063);
or U3450 (N_3450,N_3116,N_3065);
and U3451 (N_3451,N_3047,N_3066);
nand U3452 (N_3452,N_3165,N_3023);
nand U3453 (N_3453,N_3019,N_3181);
nand U3454 (N_3454,N_3013,N_3144);
and U3455 (N_3455,N_3186,N_3096);
and U3456 (N_3456,N_3094,N_3173);
and U3457 (N_3457,N_3063,N_3070);
and U3458 (N_3458,N_3061,N_3166);
and U3459 (N_3459,N_3050,N_3147);
nand U3460 (N_3460,N_3185,N_3151);
nand U3461 (N_3461,N_3186,N_3204);
xnor U3462 (N_3462,N_3063,N_3228);
nand U3463 (N_3463,N_3068,N_3153);
xor U3464 (N_3464,N_3116,N_3124);
or U3465 (N_3465,N_3189,N_3112);
and U3466 (N_3466,N_3113,N_3192);
nor U3467 (N_3467,N_3218,N_3212);
or U3468 (N_3468,N_3190,N_3160);
nand U3469 (N_3469,N_3021,N_3010);
nand U3470 (N_3470,N_3226,N_3051);
xnor U3471 (N_3471,N_3124,N_3117);
or U3472 (N_3472,N_3086,N_3139);
xnor U3473 (N_3473,N_3142,N_3002);
nand U3474 (N_3474,N_3194,N_3165);
xor U3475 (N_3475,N_3049,N_3207);
nand U3476 (N_3476,N_3037,N_3086);
nand U3477 (N_3477,N_3027,N_3242);
or U3478 (N_3478,N_3010,N_3199);
or U3479 (N_3479,N_3158,N_3207);
nand U3480 (N_3480,N_3032,N_3127);
xnor U3481 (N_3481,N_3030,N_3117);
nor U3482 (N_3482,N_3128,N_3101);
nand U3483 (N_3483,N_3240,N_3096);
xor U3484 (N_3484,N_3047,N_3034);
xnor U3485 (N_3485,N_3056,N_3122);
nor U3486 (N_3486,N_3053,N_3083);
xor U3487 (N_3487,N_3039,N_3151);
or U3488 (N_3488,N_3134,N_3124);
and U3489 (N_3489,N_3140,N_3005);
nor U3490 (N_3490,N_3090,N_3139);
and U3491 (N_3491,N_3125,N_3152);
nor U3492 (N_3492,N_3079,N_3030);
xnor U3493 (N_3493,N_3059,N_3190);
and U3494 (N_3494,N_3000,N_3125);
nand U3495 (N_3495,N_3195,N_3017);
or U3496 (N_3496,N_3151,N_3058);
nor U3497 (N_3497,N_3189,N_3177);
or U3498 (N_3498,N_3076,N_3104);
xor U3499 (N_3499,N_3082,N_3139);
and U3500 (N_3500,N_3488,N_3491);
and U3501 (N_3501,N_3463,N_3264);
xnor U3502 (N_3502,N_3442,N_3428);
nor U3503 (N_3503,N_3464,N_3283);
and U3504 (N_3504,N_3447,N_3468);
or U3505 (N_3505,N_3471,N_3370);
xor U3506 (N_3506,N_3485,N_3494);
xor U3507 (N_3507,N_3361,N_3389);
nand U3508 (N_3508,N_3265,N_3415);
xnor U3509 (N_3509,N_3408,N_3277);
nand U3510 (N_3510,N_3307,N_3337);
and U3511 (N_3511,N_3469,N_3425);
nand U3512 (N_3512,N_3481,N_3490);
or U3513 (N_3513,N_3309,N_3477);
or U3514 (N_3514,N_3317,N_3405);
nand U3515 (N_3515,N_3313,N_3434);
and U3516 (N_3516,N_3263,N_3302);
or U3517 (N_3517,N_3465,N_3461);
xnor U3518 (N_3518,N_3418,N_3303);
or U3519 (N_3519,N_3320,N_3406);
xnor U3520 (N_3520,N_3385,N_3274);
or U3521 (N_3521,N_3430,N_3330);
and U3522 (N_3522,N_3437,N_3279);
or U3523 (N_3523,N_3338,N_3432);
or U3524 (N_3524,N_3484,N_3456);
or U3525 (N_3525,N_3394,N_3280);
nor U3526 (N_3526,N_3399,N_3422);
or U3527 (N_3527,N_3288,N_3278);
and U3528 (N_3528,N_3416,N_3450);
nor U3529 (N_3529,N_3296,N_3275);
and U3530 (N_3530,N_3344,N_3261);
nor U3531 (N_3531,N_3300,N_3446);
xnor U3532 (N_3532,N_3374,N_3487);
or U3533 (N_3533,N_3329,N_3351);
or U3534 (N_3534,N_3332,N_3298);
and U3535 (N_3535,N_3496,N_3276);
nor U3536 (N_3536,N_3397,N_3480);
and U3537 (N_3537,N_3402,N_3258);
nor U3538 (N_3538,N_3323,N_3368);
and U3539 (N_3539,N_3474,N_3305);
nand U3540 (N_3540,N_3380,N_3472);
nand U3541 (N_3541,N_3377,N_3414);
nor U3542 (N_3542,N_3255,N_3401);
or U3543 (N_3543,N_3322,N_3269);
nor U3544 (N_3544,N_3365,N_3343);
or U3545 (N_3545,N_3433,N_3455);
xor U3546 (N_3546,N_3440,N_3346);
or U3547 (N_3547,N_3321,N_3387);
and U3548 (N_3548,N_3376,N_3478);
nor U3549 (N_3549,N_3467,N_3498);
xor U3550 (N_3550,N_3292,N_3452);
nor U3551 (N_3551,N_3395,N_3366);
and U3552 (N_3552,N_3459,N_3407);
nand U3553 (N_3553,N_3358,N_3411);
or U3554 (N_3554,N_3492,N_3423);
and U3555 (N_3555,N_3350,N_3482);
and U3556 (N_3556,N_3340,N_3372);
and U3557 (N_3557,N_3266,N_3383);
or U3558 (N_3558,N_3285,N_3268);
nor U3559 (N_3559,N_3435,N_3308);
nand U3560 (N_3560,N_3250,N_3347);
or U3561 (N_3561,N_3331,N_3354);
nor U3562 (N_3562,N_3345,N_3282);
or U3563 (N_3563,N_3257,N_3431);
nand U3564 (N_3564,N_3339,N_3436);
and U3565 (N_3565,N_3324,N_3475);
or U3566 (N_3566,N_3386,N_3390);
xnor U3567 (N_3567,N_3391,N_3497);
and U3568 (N_3568,N_3449,N_3438);
xnor U3569 (N_3569,N_3448,N_3462);
or U3570 (N_3570,N_3403,N_3404);
nor U3571 (N_3571,N_3342,N_3392);
or U3572 (N_3572,N_3429,N_3336);
nor U3573 (N_3573,N_3284,N_3316);
nand U3574 (N_3574,N_3364,N_3291);
and U3575 (N_3575,N_3454,N_3355);
xor U3576 (N_3576,N_3356,N_3443);
and U3577 (N_3577,N_3259,N_3352);
xnor U3578 (N_3578,N_3427,N_3493);
xor U3579 (N_3579,N_3293,N_3318);
xor U3580 (N_3580,N_3379,N_3333);
or U3581 (N_3581,N_3286,N_3299);
and U3582 (N_3582,N_3260,N_3382);
xor U3583 (N_3583,N_3476,N_3486);
nor U3584 (N_3584,N_3470,N_3326);
and U3585 (N_3585,N_3473,N_3357);
and U3586 (N_3586,N_3360,N_3328);
xor U3587 (N_3587,N_3310,N_3410);
xnor U3588 (N_3588,N_3290,N_3396);
xor U3589 (N_3589,N_3348,N_3419);
nand U3590 (N_3590,N_3256,N_3426);
or U3591 (N_3591,N_3417,N_3499);
or U3592 (N_3592,N_3388,N_3363);
and U3593 (N_3593,N_3319,N_3334);
nand U3594 (N_3594,N_3311,N_3420);
nand U3595 (N_3595,N_3281,N_3267);
nor U3596 (N_3596,N_3445,N_3453);
nor U3597 (N_3597,N_3295,N_3272);
nand U3598 (N_3598,N_3400,N_3335);
nand U3599 (N_3599,N_3362,N_3341);
or U3600 (N_3600,N_3353,N_3271);
nor U3601 (N_3601,N_3252,N_3312);
or U3602 (N_3602,N_3254,N_3439);
nand U3603 (N_3603,N_3375,N_3421);
xor U3604 (N_3604,N_3384,N_3409);
nand U3605 (N_3605,N_3460,N_3458);
nor U3606 (N_3606,N_3251,N_3381);
or U3607 (N_3607,N_3495,N_3479);
nor U3608 (N_3608,N_3413,N_3393);
xor U3609 (N_3609,N_3327,N_3466);
and U3610 (N_3610,N_3304,N_3270);
and U3611 (N_3611,N_3424,N_3441);
nand U3612 (N_3612,N_3349,N_3412);
nor U3613 (N_3613,N_3483,N_3325);
nand U3614 (N_3614,N_3287,N_3301);
and U3615 (N_3615,N_3378,N_3489);
xor U3616 (N_3616,N_3451,N_3253);
or U3617 (N_3617,N_3444,N_3294);
nor U3618 (N_3618,N_3262,N_3273);
xor U3619 (N_3619,N_3457,N_3367);
nor U3620 (N_3620,N_3369,N_3359);
or U3621 (N_3621,N_3297,N_3306);
or U3622 (N_3622,N_3289,N_3315);
nand U3623 (N_3623,N_3373,N_3371);
nand U3624 (N_3624,N_3314,N_3398);
or U3625 (N_3625,N_3258,N_3370);
nand U3626 (N_3626,N_3384,N_3289);
or U3627 (N_3627,N_3402,N_3496);
nand U3628 (N_3628,N_3358,N_3407);
xor U3629 (N_3629,N_3462,N_3312);
or U3630 (N_3630,N_3476,N_3320);
and U3631 (N_3631,N_3258,N_3332);
or U3632 (N_3632,N_3326,N_3336);
and U3633 (N_3633,N_3471,N_3497);
xor U3634 (N_3634,N_3408,N_3251);
nor U3635 (N_3635,N_3404,N_3455);
or U3636 (N_3636,N_3251,N_3429);
xnor U3637 (N_3637,N_3484,N_3449);
nor U3638 (N_3638,N_3458,N_3291);
nor U3639 (N_3639,N_3304,N_3443);
and U3640 (N_3640,N_3408,N_3328);
xor U3641 (N_3641,N_3252,N_3469);
and U3642 (N_3642,N_3434,N_3334);
and U3643 (N_3643,N_3368,N_3406);
xnor U3644 (N_3644,N_3476,N_3309);
or U3645 (N_3645,N_3445,N_3419);
or U3646 (N_3646,N_3486,N_3442);
and U3647 (N_3647,N_3469,N_3417);
xnor U3648 (N_3648,N_3490,N_3370);
nand U3649 (N_3649,N_3261,N_3462);
nor U3650 (N_3650,N_3405,N_3315);
and U3651 (N_3651,N_3264,N_3286);
xor U3652 (N_3652,N_3428,N_3353);
or U3653 (N_3653,N_3361,N_3409);
or U3654 (N_3654,N_3304,N_3451);
nand U3655 (N_3655,N_3454,N_3380);
nor U3656 (N_3656,N_3389,N_3431);
nor U3657 (N_3657,N_3352,N_3274);
or U3658 (N_3658,N_3409,N_3454);
and U3659 (N_3659,N_3286,N_3393);
xor U3660 (N_3660,N_3379,N_3325);
nor U3661 (N_3661,N_3481,N_3495);
xor U3662 (N_3662,N_3353,N_3276);
nand U3663 (N_3663,N_3408,N_3393);
nor U3664 (N_3664,N_3445,N_3300);
and U3665 (N_3665,N_3372,N_3448);
nand U3666 (N_3666,N_3420,N_3339);
nand U3667 (N_3667,N_3369,N_3472);
and U3668 (N_3668,N_3323,N_3307);
nand U3669 (N_3669,N_3346,N_3381);
nand U3670 (N_3670,N_3447,N_3334);
nor U3671 (N_3671,N_3422,N_3293);
nor U3672 (N_3672,N_3485,N_3484);
nor U3673 (N_3673,N_3394,N_3437);
and U3674 (N_3674,N_3270,N_3454);
nor U3675 (N_3675,N_3496,N_3261);
and U3676 (N_3676,N_3292,N_3327);
nor U3677 (N_3677,N_3414,N_3331);
nand U3678 (N_3678,N_3304,N_3403);
nand U3679 (N_3679,N_3333,N_3366);
or U3680 (N_3680,N_3360,N_3473);
nor U3681 (N_3681,N_3449,N_3284);
nand U3682 (N_3682,N_3377,N_3312);
and U3683 (N_3683,N_3453,N_3437);
or U3684 (N_3684,N_3320,N_3385);
nor U3685 (N_3685,N_3282,N_3378);
xnor U3686 (N_3686,N_3471,N_3259);
nand U3687 (N_3687,N_3253,N_3329);
xnor U3688 (N_3688,N_3496,N_3294);
xor U3689 (N_3689,N_3425,N_3338);
nand U3690 (N_3690,N_3367,N_3309);
nand U3691 (N_3691,N_3458,N_3408);
nand U3692 (N_3692,N_3468,N_3451);
or U3693 (N_3693,N_3493,N_3290);
xor U3694 (N_3694,N_3276,N_3459);
or U3695 (N_3695,N_3327,N_3471);
nand U3696 (N_3696,N_3269,N_3252);
xor U3697 (N_3697,N_3351,N_3267);
nor U3698 (N_3698,N_3364,N_3489);
and U3699 (N_3699,N_3276,N_3392);
and U3700 (N_3700,N_3493,N_3436);
or U3701 (N_3701,N_3354,N_3297);
or U3702 (N_3702,N_3383,N_3409);
and U3703 (N_3703,N_3374,N_3342);
xnor U3704 (N_3704,N_3422,N_3473);
xor U3705 (N_3705,N_3296,N_3455);
or U3706 (N_3706,N_3319,N_3261);
xnor U3707 (N_3707,N_3364,N_3443);
and U3708 (N_3708,N_3403,N_3497);
nor U3709 (N_3709,N_3441,N_3273);
or U3710 (N_3710,N_3478,N_3327);
and U3711 (N_3711,N_3441,N_3453);
xnor U3712 (N_3712,N_3382,N_3291);
and U3713 (N_3713,N_3291,N_3490);
and U3714 (N_3714,N_3277,N_3393);
and U3715 (N_3715,N_3370,N_3363);
nand U3716 (N_3716,N_3494,N_3306);
nor U3717 (N_3717,N_3345,N_3474);
xnor U3718 (N_3718,N_3300,N_3291);
xnor U3719 (N_3719,N_3362,N_3438);
and U3720 (N_3720,N_3363,N_3434);
nor U3721 (N_3721,N_3322,N_3458);
xnor U3722 (N_3722,N_3343,N_3408);
nand U3723 (N_3723,N_3496,N_3269);
xnor U3724 (N_3724,N_3263,N_3359);
and U3725 (N_3725,N_3351,N_3326);
nand U3726 (N_3726,N_3398,N_3389);
nand U3727 (N_3727,N_3271,N_3286);
xor U3728 (N_3728,N_3377,N_3293);
nand U3729 (N_3729,N_3316,N_3425);
or U3730 (N_3730,N_3408,N_3318);
and U3731 (N_3731,N_3467,N_3347);
and U3732 (N_3732,N_3320,N_3363);
nand U3733 (N_3733,N_3472,N_3287);
or U3734 (N_3734,N_3406,N_3420);
nand U3735 (N_3735,N_3293,N_3294);
nand U3736 (N_3736,N_3397,N_3393);
nor U3737 (N_3737,N_3372,N_3405);
nor U3738 (N_3738,N_3276,N_3384);
and U3739 (N_3739,N_3264,N_3499);
and U3740 (N_3740,N_3268,N_3408);
xor U3741 (N_3741,N_3348,N_3398);
nor U3742 (N_3742,N_3310,N_3482);
nor U3743 (N_3743,N_3329,N_3392);
and U3744 (N_3744,N_3314,N_3255);
xor U3745 (N_3745,N_3289,N_3349);
xnor U3746 (N_3746,N_3386,N_3372);
xnor U3747 (N_3747,N_3398,N_3444);
and U3748 (N_3748,N_3499,N_3420);
xor U3749 (N_3749,N_3489,N_3483);
nand U3750 (N_3750,N_3599,N_3675);
nand U3751 (N_3751,N_3501,N_3567);
or U3752 (N_3752,N_3720,N_3524);
xnor U3753 (N_3753,N_3657,N_3603);
xnor U3754 (N_3754,N_3612,N_3595);
nand U3755 (N_3755,N_3727,N_3505);
and U3756 (N_3756,N_3562,N_3651);
nor U3757 (N_3757,N_3556,N_3633);
nor U3758 (N_3758,N_3665,N_3632);
and U3759 (N_3759,N_3564,N_3647);
nand U3760 (N_3760,N_3620,N_3604);
nand U3761 (N_3761,N_3581,N_3629);
or U3762 (N_3762,N_3705,N_3573);
nand U3763 (N_3763,N_3710,N_3623);
or U3764 (N_3764,N_3578,N_3683);
and U3765 (N_3765,N_3537,N_3659);
nor U3766 (N_3766,N_3511,N_3534);
nand U3767 (N_3767,N_3697,N_3731);
and U3768 (N_3768,N_3518,N_3570);
and U3769 (N_3769,N_3638,N_3611);
nor U3770 (N_3770,N_3718,N_3698);
xor U3771 (N_3771,N_3666,N_3589);
nor U3772 (N_3772,N_3502,N_3553);
and U3773 (N_3773,N_3580,N_3596);
and U3774 (N_3774,N_3572,N_3601);
nand U3775 (N_3775,N_3500,N_3559);
nand U3776 (N_3776,N_3636,N_3643);
or U3777 (N_3777,N_3723,N_3674);
and U3778 (N_3778,N_3712,N_3520);
xnor U3779 (N_3779,N_3563,N_3726);
nand U3780 (N_3780,N_3746,N_3729);
nor U3781 (N_3781,N_3598,N_3584);
xnor U3782 (N_3782,N_3645,N_3615);
and U3783 (N_3783,N_3652,N_3528);
nor U3784 (N_3784,N_3625,N_3725);
nor U3785 (N_3785,N_3579,N_3531);
or U3786 (N_3786,N_3655,N_3660);
or U3787 (N_3787,N_3715,N_3521);
nor U3788 (N_3788,N_3621,N_3646);
nor U3789 (N_3789,N_3624,N_3716);
nor U3790 (N_3790,N_3680,N_3701);
nand U3791 (N_3791,N_3552,N_3738);
nand U3792 (N_3792,N_3558,N_3508);
nand U3793 (N_3793,N_3530,N_3586);
and U3794 (N_3794,N_3565,N_3679);
or U3795 (N_3795,N_3688,N_3656);
or U3796 (N_3796,N_3614,N_3529);
nor U3797 (N_3797,N_3672,N_3702);
xnor U3798 (N_3798,N_3661,N_3664);
or U3799 (N_3799,N_3618,N_3700);
and U3800 (N_3800,N_3594,N_3554);
nor U3801 (N_3801,N_3551,N_3635);
and U3802 (N_3802,N_3536,N_3736);
nor U3803 (N_3803,N_3662,N_3512);
nor U3804 (N_3804,N_3639,N_3577);
and U3805 (N_3805,N_3732,N_3694);
nor U3806 (N_3806,N_3525,N_3709);
xor U3807 (N_3807,N_3619,N_3569);
or U3808 (N_3808,N_3613,N_3609);
xor U3809 (N_3809,N_3644,N_3587);
nand U3810 (N_3810,N_3591,N_3583);
nor U3811 (N_3811,N_3542,N_3742);
nand U3812 (N_3812,N_3538,N_3676);
nor U3813 (N_3813,N_3574,N_3699);
nor U3814 (N_3814,N_3653,N_3717);
xor U3815 (N_3815,N_3622,N_3745);
nand U3816 (N_3816,N_3548,N_3634);
nand U3817 (N_3817,N_3741,N_3748);
or U3818 (N_3818,N_3515,N_3550);
and U3819 (N_3819,N_3541,N_3503);
xor U3820 (N_3820,N_3734,N_3744);
xnor U3821 (N_3821,N_3728,N_3690);
nand U3822 (N_3822,N_3555,N_3517);
xnor U3823 (N_3823,N_3602,N_3606);
and U3824 (N_3824,N_3608,N_3504);
or U3825 (N_3825,N_3509,N_3730);
xnor U3826 (N_3826,N_3630,N_3575);
or U3827 (N_3827,N_3669,N_3719);
and U3828 (N_3828,N_3631,N_3540);
nor U3829 (N_3829,N_3616,N_3549);
or U3830 (N_3830,N_3686,N_3582);
and U3831 (N_3831,N_3733,N_3641);
nand U3832 (N_3832,N_3506,N_3585);
xor U3833 (N_3833,N_3740,N_3708);
nor U3834 (N_3834,N_3650,N_3628);
nand U3835 (N_3835,N_3626,N_3514);
xnor U3836 (N_3836,N_3667,N_3689);
nor U3837 (N_3837,N_3747,N_3571);
nand U3838 (N_3838,N_3678,N_3670);
and U3839 (N_3839,N_3545,N_3663);
nor U3840 (N_3840,N_3649,N_3658);
and U3841 (N_3841,N_3544,N_3673);
nor U3842 (N_3842,N_3607,N_3714);
nor U3843 (N_3843,N_3510,N_3706);
or U3844 (N_3844,N_3737,N_3576);
or U3845 (N_3845,N_3681,N_3704);
nor U3846 (N_3846,N_3560,N_3677);
nor U3847 (N_3847,N_3668,N_3566);
nor U3848 (N_3848,N_3735,N_3523);
and U3849 (N_3849,N_3724,N_3610);
xor U3850 (N_3850,N_3527,N_3546);
or U3851 (N_3851,N_3627,N_3507);
and U3852 (N_3852,N_3532,N_3597);
nor U3853 (N_3853,N_3695,N_3691);
nor U3854 (N_3854,N_3654,N_3588);
and U3855 (N_3855,N_3547,N_3693);
nor U3856 (N_3856,N_3722,N_3605);
nand U3857 (N_3857,N_3711,N_3671);
xnor U3858 (N_3858,N_3743,N_3590);
xor U3859 (N_3859,N_3749,N_3600);
xnor U3860 (N_3860,N_3557,N_3642);
and U3861 (N_3861,N_3539,N_3516);
or U3862 (N_3862,N_3692,N_3543);
nand U3863 (N_3863,N_3687,N_3721);
xor U3864 (N_3864,N_3640,N_3519);
nand U3865 (N_3865,N_3739,N_3617);
xor U3866 (N_3866,N_3513,N_3682);
and U3867 (N_3867,N_3561,N_3522);
and U3868 (N_3868,N_3568,N_3535);
or U3869 (N_3869,N_3703,N_3637);
nor U3870 (N_3870,N_3592,N_3593);
nand U3871 (N_3871,N_3533,N_3696);
nand U3872 (N_3872,N_3684,N_3526);
xor U3873 (N_3873,N_3648,N_3707);
nand U3874 (N_3874,N_3713,N_3685);
nor U3875 (N_3875,N_3539,N_3575);
nor U3876 (N_3876,N_3599,N_3641);
or U3877 (N_3877,N_3600,N_3568);
and U3878 (N_3878,N_3650,N_3729);
and U3879 (N_3879,N_3581,N_3545);
nand U3880 (N_3880,N_3563,N_3576);
nor U3881 (N_3881,N_3526,N_3558);
or U3882 (N_3882,N_3700,N_3531);
or U3883 (N_3883,N_3510,N_3579);
and U3884 (N_3884,N_3556,N_3640);
nand U3885 (N_3885,N_3531,N_3570);
nand U3886 (N_3886,N_3739,N_3558);
or U3887 (N_3887,N_3731,N_3678);
xnor U3888 (N_3888,N_3572,N_3673);
and U3889 (N_3889,N_3640,N_3713);
nand U3890 (N_3890,N_3648,N_3573);
nand U3891 (N_3891,N_3635,N_3638);
xor U3892 (N_3892,N_3528,N_3635);
nand U3893 (N_3893,N_3673,N_3686);
nand U3894 (N_3894,N_3682,N_3591);
and U3895 (N_3895,N_3504,N_3559);
and U3896 (N_3896,N_3540,N_3539);
xnor U3897 (N_3897,N_3732,N_3624);
nand U3898 (N_3898,N_3617,N_3692);
nand U3899 (N_3899,N_3628,N_3535);
and U3900 (N_3900,N_3544,N_3524);
nand U3901 (N_3901,N_3556,N_3610);
or U3902 (N_3902,N_3631,N_3539);
and U3903 (N_3903,N_3717,N_3735);
or U3904 (N_3904,N_3607,N_3590);
nor U3905 (N_3905,N_3592,N_3701);
or U3906 (N_3906,N_3560,N_3553);
nand U3907 (N_3907,N_3734,N_3557);
or U3908 (N_3908,N_3539,N_3673);
nand U3909 (N_3909,N_3704,N_3651);
or U3910 (N_3910,N_3501,N_3711);
nor U3911 (N_3911,N_3749,N_3735);
xor U3912 (N_3912,N_3639,N_3697);
and U3913 (N_3913,N_3547,N_3721);
or U3914 (N_3914,N_3695,N_3703);
or U3915 (N_3915,N_3582,N_3550);
or U3916 (N_3916,N_3656,N_3554);
and U3917 (N_3917,N_3746,N_3599);
xnor U3918 (N_3918,N_3526,N_3588);
xnor U3919 (N_3919,N_3658,N_3535);
xnor U3920 (N_3920,N_3557,N_3586);
or U3921 (N_3921,N_3718,N_3740);
xnor U3922 (N_3922,N_3697,N_3554);
xor U3923 (N_3923,N_3596,N_3713);
and U3924 (N_3924,N_3611,N_3535);
xor U3925 (N_3925,N_3560,N_3565);
or U3926 (N_3926,N_3550,N_3735);
or U3927 (N_3927,N_3629,N_3697);
nand U3928 (N_3928,N_3535,N_3603);
nand U3929 (N_3929,N_3715,N_3552);
and U3930 (N_3930,N_3721,N_3657);
or U3931 (N_3931,N_3678,N_3655);
xor U3932 (N_3932,N_3677,N_3537);
or U3933 (N_3933,N_3532,N_3523);
or U3934 (N_3934,N_3718,N_3677);
and U3935 (N_3935,N_3747,N_3619);
xnor U3936 (N_3936,N_3748,N_3690);
or U3937 (N_3937,N_3705,N_3718);
nor U3938 (N_3938,N_3635,N_3508);
nor U3939 (N_3939,N_3638,N_3571);
nand U3940 (N_3940,N_3676,N_3510);
xnor U3941 (N_3941,N_3587,N_3635);
nand U3942 (N_3942,N_3557,N_3740);
xnor U3943 (N_3943,N_3652,N_3737);
and U3944 (N_3944,N_3582,N_3748);
or U3945 (N_3945,N_3648,N_3566);
nand U3946 (N_3946,N_3657,N_3736);
or U3947 (N_3947,N_3510,N_3665);
nor U3948 (N_3948,N_3721,N_3561);
and U3949 (N_3949,N_3516,N_3619);
or U3950 (N_3950,N_3681,N_3576);
nand U3951 (N_3951,N_3627,N_3601);
and U3952 (N_3952,N_3601,N_3626);
and U3953 (N_3953,N_3679,N_3541);
nor U3954 (N_3954,N_3599,N_3745);
nand U3955 (N_3955,N_3534,N_3519);
xor U3956 (N_3956,N_3556,N_3703);
or U3957 (N_3957,N_3597,N_3590);
or U3958 (N_3958,N_3666,N_3556);
nand U3959 (N_3959,N_3541,N_3715);
and U3960 (N_3960,N_3644,N_3683);
xnor U3961 (N_3961,N_3526,N_3545);
xor U3962 (N_3962,N_3592,N_3551);
xnor U3963 (N_3963,N_3597,N_3729);
nor U3964 (N_3964,N_3701,N_3682);
nand U3965 (N_3965,N_3517,N_3675);
and U3966 (N_3966,N_3615,N_3596);
or U3967 (N_3967,N_3500,N_3643);
xor U3968 (N_3968,N_3515,N_3629);
or U3969 (N_3969,N_3719,N_3718);
nor U3970 (N_3970,N_3519,N_3555);
or U3971 (N_3971,N_3520,N_3565);
or U3972 (N_3972,N_3749,N_3610);
or U3973 (N_3973,N_3610,N_3671);
or U3974 (N_3974,N_3585,N_3705);
and U3975 (N_3975,N_3717,N_3615);
or U3976 (N_3976,N_3547,N_3646);
and U3977 (N_3977,N_3660,N_3533);
nor U3978 (N_3978,N_3607,N_3721);
nand U3979 (N_3979,N_3540,N_3524);
xnor U3980 (N_3980,N_3639,N_3546);
nand U3981 (N_3981,N_3702,N_3547);
or U3982 (N_3982,N_3668,N_3670);
nor U3983 (N_3983,N_3606,N_3710);
nor U3984 (N_3984,N_3592,N_3743);
and U3985 (N_3985,N_3739,N_3644);
and U3986 (N_3986,N_3572,N_3589);
or U3987 (N_3987,N_3728,N_3672);
xor U3988 (N_3988,N_3643,N_3644);
xnor U3989 (N_3989,N_3675,N_3538);
nand U3990 (N_3990,N_3729,N_3539);
and U3991 (N_3991,N_3559,N_3521);
nor U3992 (N_3992,N_3573,N_3580);
and U3993 (N_3993,N_3588,N_3504);
and U3994 (N_3994,N_3601,N_3611);
and U3995 (N_3995,N_3624,N_3627);
nand U3996 (N_3996,N_3602,N_3663);
xor U3997 (N_3997,N_3522,N_3714);
xor U3998 (N_3998,N_3727,N_3703);
and U3999 (N_3999,N_3731,N_3560);
xnor U4000 (N_4000,N_3837,N_3758);
nor U4001 (N_4001,N_3816,N_3801);
xor U4002 (N_4002,N_3859,N_3875);
xnor U4003 (N_4003,N_3856,N_3921);
and U4004 (N_4004,N_3999,N_3872);
xnor U4005 (N_4005,N_3917,N_3809);
nand U4006 (N_4006,N_3847,N_3838);
or U4007 (N_4007,N_3950,N_3879);
or U4008 (N_4008,N_3840,N_3902);
and U4009 (N_4009,N_3942,N_3858);
nand U4010 (N_4010,N_3947,N_3946);
or U4011 (N_4011,N_3804,N_3795);
or U4012 (N_4012,N_3799,N_3995);
nor U4013 (N_4013,N_3937,N_3752);
nand U4014 (N_4014,N_3963,N_3850);
and U4015 (N_4015,N_3834,N_3911);
or U4016 (N_4016,N_3894,N_3989);
nor U4017 (N_4017,N_3881,N_3796);
and U4018 (N_4018,N_3943,N_3852);
nor U4019 (N_4019,N_3857,N_3813);
nor U4020 (N_4020,N_3843,N_3888);
xnor U4021 (N_4021,N_3776,N_3851);
nor U4022 (N_4022,N_3835,N_3919);
nor U4023 (N_4023,N_3819,N_3922);
and U4024 (N_4024,N_3923,N_3915);
xor U4025 (N_4025,N_3787,N_3833);
and U4026 (N_4026,N_3869,N_3968);
nor U4027 (N_4027,N_3892,N_3970);
and U4028 (N_4028,N_3790,N_3866);
xor U4029 (N_4029,N_3933,N_3750);
and U4030 (N_4030,N_3810,N_3811);
and U4031 (N_4031,N_3757,N_3972);
and U4032 (N_4032,N_3761,N_3964);
xnor U4033 (N_4033,N_3862,N_3770);
or U4034 (N_4034,N_3938,N_3756);
nor U4035 (N_4035,N_3868,N_3836);
xor U4036 (N_4036,N_3829,N_3895);
or U4037 (N_4037,N_3777,N_3969);
nor U4038 (N_4038,N_3769,N_3900);
xor U4039 (N_4039,N_3805,N_3925);
nand U4040 (N_4040,N_3981,N_3903);
and U4041 (N_4041,N_3784,N_3918);
and U4042 (N_4042,N_3967,N_3924);
nand U4043 (N_4043,N_3965,N_3909);
or U4044 (N_4044,N_3846,N_3785);
or U4045 (N_4045,N_3841,N_3788);
and U4046 (N_4046,N_3991,N_3767);
nor U4047 (N_4047,N_3887,N_3808);
nor U4048 (N_4048,N_3765,N_3945);
and U4049 (N_4049,N_3832,N_3860);
or U4050 (N_4050,N_3971,N_3980);
nand U4051 (N_4051,N_3916,N_3984);
and U4052 (N_4052,N_3885,N_3958);
or U4053 (N_4053,N_3996,N_3890);
nor U4054 (N_4054,N_3781,N_3883);
and U4055 (N_4055,N_3842,N_3762);
or U4056 (N_4056,N_3778,N_3782);
or U4057 (N_4057,N_3871,N_3771);
nand U4058 (N_4058,N_3982,N_3951);
nor U4059 (N_4059,N_3953,N_3997);
and U4060 (N_4060,N_3792,N_3960);
nor U4061 (N_4061,N_3974,N_3948);
or U4062 (N_4062,N_3753,N_3914);
nand U4063 (N_4063,N_3814,N_3907);
and U4064 (N_4064,N_3789,N_3825);
nor U4065 (N_4065,N_3961,N_3830);
nor U4066 (N_4066,N_3807,N_3904);
nand U4067 (N_4067,N_3793,N_3978);
nor U4068 (N_4068,N_3998,N_3927);
nor U4069 (N_4069,N_3768,N_3826);
and U4070 (N_4070,N_3763,N_3912);
nor U4071 (N_4071,N_3905,N_3934);
nand U4072 (N_4072,N_3774,N_3820);
xnor U4073 (N_4073,N_3977,N_3880);
nor U4074 (N_4074,N_3992,N_3959);
nor U4075 (N_4075,N_3786,N_3928);
and U4076 (N_4076,N_3944,N_3855);
or U4077 (N_4077,N_3818,N_3764);
xnor U4078 (N_4078,N_3876,N_3821);
or U4079 (N_4079,N_3754,N_3831);
nand U4080 (N_4080,N_3973,N_3863);
nor U4081 (N_4081,N_3898,N_3962);
or U4082 (N_4082,N_3854,N_3983);
xor U4083 (N_4083,N_3791,N_3824);
or U4084 (N_4084,N_3920,N_3844);
and U4085 (N_4085,N_3775,N_3882);
or U4086 (N_4086,N_3957,N_3751);
and U4087 (N_4087,N_3861,N_3952);
nand U4088 (N_4088,N_3899,N_3865);
nor U4089 (N_4089,N_3932,N_3823);
xnor U4090 (N_4090,N_3822,N_3845);
and U4091 (N_4091,N_3812,N_3800);
nor U4092 (N_4092,N_3896,N_3755);
and U4093 (N_4093,N_3955,N_3891);
xor U4094 (N_4094,N_3908,N_3884);
nand U4095 (N_4095,N_3941,N_3798);
nand U4096 (N_4096,N_3929,N_3780);
or U4097 (N_4097,N_3802,N_3940);
nand U4098 (N_4098,N_3779,N_3783);
and U4099 (N_4099,N_3935,N_3772);
and U4100 (N_4100,N_3975,N_3913);
nor U4101 (N_4101,N_3985,N_3873);
and U4102 (N_4102,N_3870,N_3986);
nand U4103 (N_4103,N_3874,N_3901);
or U4104 (N_4104,N_3966,N_3759);
and U4105 (N_4105,N_3848,N_3877);
nand U4106 (N_4106,N_3910,N_3864);
nand U4107 (N_4107,N_3760,N_3797);
xor U4108 (N_4108,N_3878,N_3988);
or U4109 (N_4109,N_3853,N_3990);
xor U4110 (N_4110,N_3794,N_3926);
or U4111 (N_4111,N_3936,N_3766);
nand U4112 (N_4112,N_3897,N_3939);
nand U4113 (N_4113,N_3849,N_3979);
nor U4114 (N_4114,N_3930,N_3949);
and U4115 (N_4115,N_3886,N_3773);
and U4116 (N_4116,N_3976,N_3889);
xor U4117 (N_4117,N_3817,N_3906);
and U4118 (N_4118,N_3956,N_3993);
nand U4119 (N_4119,N_3867,N_3806);
xor U4120 (N_4120,N_3994,N_3815);
nand U4121 (N_4121,N_3954,N_3827);
or U4122 (N_4122,N_3828,N_3803);
nor U4123 (N_4123,N_3839,N_3893);
nand U4124 (N_4124,N_3987,N_3931);
nor U4125 (N_4125,N_3771,N_3874);
xor U4126 (N_4126,N_3962,N_3960);
nand U4127 (N_4127,N_3802,N_3939);
and U4128 (N_4128,N_3851,N_3819);
or U4129 (N_4129,N_3935,N_3765);
xnor U4130 (N_4130,N_3942,N_3965);
nand U4131 (N_4131,N_3916,N_3914);
nor U4132 (N_4132,N_3890,N_3787);
or U4133 (N_4133,N_3991,N_3946);
nor U4134 (N_4134,N_3840,N_3899);
nor U4135 (N_4135,N_3815,N_3803);
nor U4136 (N_4136,N_3830,N_3818);
nor U4137 (N_4137,N_3849,N_3840);
xnor U4138 (N_4138,N_3928,N_3843);
and U4139 (N_4139,N_3923,N_3846);
and U4140 (N_4140,N_3784,N_3754);
xor U4141 (N_4141,N_3835,N_3946);
or U4142 (N_4142,N_3822,N_3981);
nor U4143 (N_4143,N_3767,N_3776);
or U4144 (N_4144,N_3908,N_3790);
nand U4145 (N_4145,N_3772,N_3822);
nor U4146 (N_4146,N_3924,N_3996);
nor U4147 (N_4147,N_3940,N_3824);
nor U4148 (N_4148,N_3949,N_3778);
xnor U4149 (N_4149,N_3860,N_3990);
or U4150 (N_4150,N_3800,N_3983);
nand U4151 (N_4151,N_3954,N_3793);
nand U4152 (N_4152,N_3795,N_3762);
nand U4153 (N_4153,N_3905,N_3912);
nand U4154 (N_4154,N_3795,N_3852);
nand U4155 (N_4155,N_3905,N_3816);
or U4156 (N_4156,N_3852,N_3819);
nor U4157 (N_4157,N_3854,N_3925);
xnor U4158 (N_4158,N_3766,N_3903);
nor U4159 (N_4159,N_3873,N_3893);
xnor U4160 (N_4160,N_3911,N_3902);
and U4161 (N_4161,N_3961,N_3973);
xnor U4162 (N_4162,N_3873,N_3762);
nor U4163 (N_4163,N_3980,N_3931);
or U4164 (N_4164,N_3996,N_3779);
nor U4165 (N_4165,N_3903,N_3873);
nor U4166 (N_4166,N_3940,N_3915);
nor U4167 (N_4167,N_3970,N_3762);
or U4168 (N_4168,N_3964,N_3790);
and U4169 (N_4169,N_3966,N_3985);
nor U4170 (N_4170,N_3771,N_3832);
xor U4171 (N_4171,N_3908,N_3937);
nand U4172 (N_4172,N_3951,N_3856);
nor U4173 (N_4173,N_3925,N_3983);
or U4174 (N_4174,N_3835,N_3762);
nor U4175 (N_4175,N_3750,N_3872);
and U4176 (N_4176,N_3752,N_3932);
nor U4177 (N_4177,N_3929,N_3799);
nand U4178 (N_4178,N_3793,N_3848);
nor U4179 (N_4179,N_3763,N_3818);
nor U4180 (N_4180,N_3917,N_3982);
nor U4181 (N_4181,N_3926,N_3788);
nand U4182 (N_4182,N_3965,N_3847);
nor U4183 (N_4183,N_3824,N_3999);
and U4184 (N_4184,N_3926,N_3973);
nor U4185 (N_4185,N_3935,N_3766);
xnor U4186 (N_4186,N_3890,N_3972);
and U4187 (N_4187,N_3821,N_3783);
nor U4188 (N_4188,N_3804,N_3849);
nand U4189 (N_4189,N_3802,N_3883);
nand U4190 (N_4190,N_3944,N_3912);
nand U4191 (N_4191,N_3772,N_3937);
nor U4192 (N_4192,N_3918,N_3838);
or U4193 (N_4193,N_3804,N_3775);
xor U4194 (N_4194,N_3912,N_3825);
nand U4195 (N_4195,N_3754,N_3964);
nand U4196 (N_4196,N_3841,N_3948);
or U4197 (N_4197,N_3841,N_3925);
nor U4198 (N_4198,N_3974,N_3934);
nor U4199 (N_4199,N_3872,N_3769);
and U4200 (N_4200,N_3950,N_3783);
nor U4201 (N_4201,N_3996,N_3750);
or U4202 (N_4202,N_3937,N_3796);
nor U4203 (N_4203,N_3834,N_3781);
xnor U4204 (N_4204,N_3960,N_3853);
or U4205 (N_4205,N_3810,N_3830);
xor U4206 (N_4206,N_3954,N_3942);
xor U4207 (N_4207,N_3782,N_3787);
nor U4208 (N_4208,N_3922,N_3978);
and U4209 (N_4209,N_3885,N_3966);
xor U4210 (N_4210,N_3950,N_3999);
xor U4211 (N_4211,N_3991,N_3967);
or U4212 (N_4212,N_3866,N_3819);
nand U4213 (N_4213,N_3897,N_3902);
nor U4214 (N_4214,N_3813,N_3799);
and U4215 (N_4215,N_3975,N_3923);
nor U4216 (N_4216,N_3983,N_3894);
and U4217 (N_4217,N_3787,N_3907);
or U4218 (N_4218,N_3994,N_3911);
or U4219 (N_4219,N_3981,N_3904);
nor U4220 (N_4220,N_3961,N_3840);
or U4221 (N_4221,N_3799,N_3977);
nor U4222 (N_4222,N_3821,N_3955);
and U4223 (N_4223,N_3974,N_3773);
nand U4224 (N_4224,N_3998,N_3972);
or U4225 (N_4225,N_3756,N_3834);
and U4226 (N_4226,N_3781,N_3856);
or U4227 (N_4227,N_3876,N_3805);
xnor U4228 (N_4228,N_3950,N_3810);
or U4229 (N_4229,N_3813,N_3771);
xnor U4230 (N_4230,N_3761,N_3984);
nor U4231 (N_4231,N_3967,N_3997);
xnor U4232 (N_4232,N_3930,N_3929);
or U4233 (N_4233,N_3821,N_3875);
and U4234 (N_4234,N_3998,N_3751);
and U4235 (N_4235,N_3932,N_3995);
nor U4236 (N_4236,N_3973,N_3788);
xnor U4237 (N_4237,N_3870,N_3840);
nor U4238 (N_4238,N_3896,N_3853);
or U4239 (N_4239,N_3833,N_3986);
or U4240 (N_4240,N_3778,N_3812);
xor U4241 (N_4241,N_3825,N_3893);
and U4242 (N_4242,N_3944,N_3907);
xnor U4243 (N_4243,N_3794,N_3927);
nor U4244 (N_4244,N_3981,N_3821);
and U4245 (N_4245,N_3795,N_3890);
xor U4246 (N_4246,N_3837,N_3763);
xnor U4247 (N_4247,N_3789,N_3893);
or U4248 (N_4248,N_3885,N_3776);
xor U4249 (N_4249,N_3998,N_3803);
or U4250 (N_4250,N_4189,N_4051);
or U4251 (N_4251,N_4018,N_4159);
and U4252 (N_4252,N_4043,N_4107);
nand U4253 (N_4253,N_4086,N_4032);
xor U4254 (N_4254,N_4034,N_4249);
nand U4255 (N_4255,N_4066,N_4015);
nor U4256 (N_4256,N_4098,N_4230);
or U4257 (N_4257,N_4198,N_4094);
and U4258 (N_4258,N_4220,N_4076);
or U4259 (N_4259,N_4192,N_4138);
xnor U4260 (N_4260,N_4110,N_4025);
xor U4261 (N_4261,N_4170,N_4241);
xor U4262 (N_4262,N_4233,N_4112);
nor U4263 (N_4263,N_4193,N_4119);
and U4264 (N_4264,N_4105,N_4176);
nand U4265 (N_4265,N_4134,N_4153);
nand U4266 (N_4266,N_4007,N_4167);
or U4267 (N_4267,N_4169,N_4190);
nor U4268 (N_4268,N_4040,N_4054);
nor U4269 (N_4269,N_4180,N_4000);
xnor U4270 (N_4270,N_4005,N_4046);
or U4271 (N_4271,N_4215,N_4024);
nor U4272 (N_4272,N_4232,N_4160);
or U4273 (N_4273,N_4069,N_4128);
nand U4274 (N_4274,N_4194,N_4139);
nand U4275 (N_4275,N_4207,N_4129);
or U4276 (N_4276,N_4148,N_4065);
nand U4277 (N_4277,N_4239,N_4223);
and U4278 (N_4278,N_4044,N_4212);
or U4279 (N_4279,N_4081,N_4210);
nand U4280 (N_4280,N_4203,N_4095);
or U4281 (N_4281,N_4012,N_4035);
nand U4282 (N_4282,N_4222,N_4166);
or U4283 (N_4283,N_4003,N_4175);
nand U4284 (N_4284,N_4111,N_4108);
or U4285 (N_4285,N_4201,N_4240);
nor U4286 (N_4286,N_4162,N_4038);
nand U4287 (N_4287,N_4235,N_4191);
nor U4288 (N_4288,N_4161,N_4132);
nor U4289 (N_4289,N_4186,N_4122);
xnor U4290 (N_4290,N_4195,N_4039);
nor U4291 (N_4291,N_4057,N_4197);
nor U4292 (N_4292,N_4187,N_4152);
xnor U4293 (N_4293,N_4089,N_4028);
xnor U4294 (N_4294,N_4023,N_4147);
nand U4295 (N_4295,N_4120,N_4073);
nor U4296 (N_4296,N_4059,N_4080);
and U4297 (N_4297,N_4103,N_4014);
or U4298 (N_4298,N_4131,N_4104);
xor U4299 (N_4299,N_4096,N_4199);
nand U4300 (N_4300,N_4113,N_4145);
and U4301 (N_4301,N_4181,N_4183);
nor U4302 (N_4302,N_4126,N_4174);
xor U4303 (N_4303,N_4085,N_4163);
or U4304 (N_4304,N_4157,N_4135);
and U4305 (N_4305,N_4048,N_4001);
nand U4306 (N_4306,N_4177,N_4061);
nor U4307 (N_4307,N_4021,N_4156);
or U4308 (N_4308,N_4124,N_4151);
nor U4309 (N_4309,N_4226,N_4022);
nand U4310 (N_4310,N_4248,N_4218);
nor U4311 (N_4311,N_4121,N_4228);
or U4312 (N_4312,N_4106,N_4234);
or U4313 (N_4313,N_4062,N_4036);
or U4314 (N_4314,N_4146,N_4208);
or U4315 (N_4315,N_4050,N_4206);
and U4316 (N_4316,N_4141,N_4019);
nor U4317 (N_4317,N_4155,N_4211);
xor U4318 (N_4318,N_4091,N_4002);
xnor U4319 (N_4319,N_4238,N_4053);
nand U4320 (N_4320,N_4116,N_4154);
nor U4321 (N_4321,N_4244,N_4221);
xnor U4322 (N_4322,N_4055,N_4052);
nor U4323 (N_4323,N_4075,N_4205);
nand U4324 (N_4324,N_4168,N_4149);
and U4325 (N_4325,N_4214,N_4045);
nand U4326 (N_4326,N_4172,N_4031);
and U4327 (N_4327,N_4140,N_4229);
nor U4328 (N_4328,N_4144,N_4097);
or U4329 (N_4329,N_4173,N_4142);
nor U4330 (N_4330,N_4063,N_4164);
or U4331 (N_4331,N_4067,N_4017);
xnor U4332 (N_4332,N_4087,N_4109);
nor U4333 (N_4333,N_4064,N_4016);
nand U4334 (N_4334,N_4196,N_4188);
xor U4335 (N_4335,N_4204,N_4184);
or U4336 (N_4336,N_4088,N_4093);
xnor U4337 (N_4337,N_4247,N_4008);
and U4338 (N_4338,N_4243,N_4136);
or U4339 (N_4339,N_4056,N_4101);
xor U4340 (N_4340,N_4165,N_4037);
nor U4341 (N_4341,N_4100,N_4245);
or U4342 (N_4342,N_4125,N_4074);
nand U4343 (N_4343,N_4047,N_4009);
xor U4344 (N_4344,N_4130,N_4225);
nand U4345 (N_4345,N_4082,N_4071);
nor U4346 (N_4346,N_4200,N_4060);
or U4347 (N_4347,N_4114,N_4042);
nand U4348 (N_4348,N_4219,N_4209);
xor U4349 (N_4349,N_4079,N_4185);
or U4350 (N_4350,N_4078,N_4224);
nor U4351 (N_4351,N_4083,N_4236);
and U4352 (N_4352,N_4072,N_4246);
nor U4353 (N_4353,N_4092,N_4137);
or U4354 (N_4354,N_4049,N_4026);
xor U4355 (N_4355,N_4068,N_4171);
nor U4356 (N_4356,N_4020,N_4178);
or U4357 (N_4357,N_4227,N_4127);
xor U4358 (N_4358,N_4099,N_4217);
nor U4359 (N_4359,N_4033,N_4011);
nor U4360 (N_4360,N_4182,N_4090);
nor U4361 (N_4361,N_4027,N_4030);
nand U4362 (N_4362,N_4143,N_4102);
and U4363 (N_4363,N_4213,N_4133);
nor U4364 (N_4364,N_4231,N_4123);
nor U4365 (N_4365,N_4242,N_4029);
and U4366 (N_4366,N_4118,N_4202);
and U4367 (N_4367,N_4070,N_4216);
or U4368 (N_4368,N_4004,N_4179);
xor U4369 (N_4369,N_4058,N_4013);
nor U4370 (N_4370,N_4237,N_4010);
and U4371 (N_4371,N_4117,N_4150);
xor U4372 (N_4372,N_4006,N_4158);
nor U4373 (N_4373,N_4115,N_4041);
and U4374 (N_4374,N_4084,N_4077);
nor U4375 (N_4375,N_4111,N_4028);
nand U4376 (N_4376,N_4061,N_4100);
nor U4377 (N_4377,N_4104,N_4156);
and U4378 (N_4378,N_4109,N_4118);
nand U4379 (N_4379,N_4011,N_4108);
xor U4380 (N_4380,N_4035,N_4208);
and U4381 (N_4381,N_4210,N_4020);
nor U4382 (N_4382,N_4033,N_4015);
or U4383 (N_4383,N_4211,N_4201);
or U4384 (N_4384,N_4005,N_4149);
nand U4385 (N_4385,N_4182,N_4019);
nor U4386 (N_4386,N_4171,N_4168);
nor U4387 (N_4387,N_4058,N_4195);
xnor U4388 (N_4388,N_4025,N_4038);
nand U4389 (N_4389,N_4202,N_4203);
nand U4390 (N_4390,N_4192,N_4081);
or U4391 (N_4391,N_4185,N_4083);
nand U4392 (N_4392,N_4072,N_4204);
nor U4393 (N_4393,N_4155,N_4055);
and U4394 (N_4394,N_4143,N_4241);
nand U4395 (N_4395,N_4210,N_4155);
or U4396 (N_4396,N_4063,N_4143);
or U4397 (N_4397,N_4201,N_4156);
or U4398 (N_4398,N_4120,N_4103);
and U4399 (N_4399,N_4114,N_4071);
or U4400 (N_4400,N_4233,N_4032);
or U4401 (N_4401,N_4180,N_4061);
or U4402 (N_4402,N_4210,N_4069);
or U4403 (N_4403,N_4194,N_4211);
and U4404 (N_4404,N_4010,N_4240);
nor U4405 (N_4405,N_4185,N_4242);
nor U4406 (N_4406,N_4013,N_4060);
and U4407 (N_4407,N_4054,N_4007);
and U4408 (N_4408,N_4125,N_4120);
or U4409 (N_4409,N_4133,N_4029);
and U4410 (N_4410,N_4008,N_4003);
xnor U4411 (N_4411,N_4238,N_4183);
and U4412 (N_4412,N_4164,N_4133);
and U4413 (N_4413,N_4233,N_4101);
nor U4414 (N_4414,N_4089,N_4175);
nand U4415 (N_4415,N_4112,N_4186);
nor U4416 (N_4416,N_4184,N_4182);
and U4417 (N_4417,N_4207,N_4000);
or U4418 (N_4418,N_4038,N_4171);
nand U4419 (N_4419,N_4118,N_4087);
and U4420 (N_4420,N_4049,N_4234);
or U4421 (N_4421,N_4031,N_4137);
xor U4422 (N_4422,N_4013,N_4053);
nor U4423 (N_4423,N_4115,N_4061);
and U4424 (N_4424,N_4137,N_4123);
or U4425 (N_4425,N_4205,N_4148);
xor U4426 (N_4426,N_4047,N_4000);
or U4427 (N_4427,N_4017,N_4089);
or U4428 (N_4428,N_4101,N_4160);
or U4429 (N_4429,N_4083,N_4126);
nor U4430 (N_4430,N_4096,N_4060);
and U4431 (N_4431,N_4150,N_4033);
and U4432 (N_4432,N_4200,N_4044);
or U4433 (N_4433,N_4008,N_4076);
nand U4434 (N_4434,N_4102,N_4022);
xnor U4435 (N_4435,N_4068,N_4063);
xnor U4436 (N_4436,N_4006,N_4037);
or U4437 (N_4437,N_4015,N_4163);
nor U4438 (N_4438,N_4065,N_4083);
and U4439 (N_4439,N_4050,N_4133);
and U4440 (N_4440,N_4208,N_4073);
or U4441 (N_4441,N_4043,N_4173);
or U4442 (N_4442,N_4011,N_4134);
nand U4443 (N_4443,N_4000,N_4018);
or U4444 (N_4444,N_4130,N_4147);
xnor U4445 (N_4445,N_4014,N_4054);
nand U4446 (N_4446,N_4141,N_4170);
xor U4447 (N_4447,N_4050,N_4150);
nand U4448 (N_4448,N_4000,N_4104);
and U4449 (N_4449,N_4114,N_4171);
nand U4450 (N_4450,N_4006,N_4035);
nand U4451 (N_4451,N_4153,N_4067);
xor U4452 (N_4452,N_4180,N_4126);
nor U4453 (N_4453,N_4068,N_4166);
or U4454 (N_4454,N_4065,N_4026);
and U4455 (N_4455,N_4007,N_4211);
or U4456 (N_4456,N_4200,N_4068);
or U4457 (N_4457,N_4105,N_4066);
or U4458 (N_4458,N_4137,N_4024);
nor U4459 (N_4459,N_4047,N_4168);
nand U4460 (N_4460,N_4061,N_4143);
nand U4461 (N_4461,N_4047,N_4128);
or U4462 (N_4462,N_4069,N_4000);
nor U4463 (N_4463,N_4204,N_4161);
or U4464 (N_4464,N_4249,N_4152);
nor U4465 (N_4465,N_4119,N_4098);
xor U4466 (N_4466,N_4062,N_4162);
and U4467 (N_4467,N_4008,N_4089);
and U4468 (N_4468,N_4176,N_4047);
xor U4469 (N_4469,N_4144,N_4189);
xnor U4470 (N_4470,N_4014,N_4219);
xnor U4471 (N_4471,N_4060,N_4105);
xor U4472 (N_4472,N_4068,N_4190);
xnor U4473 (N_4473,N_4142,N_4168);
nor U4474 (N_4474,N_4199,N_4187);
or U4475 (N_4475,N_4087,N_4128);
xor U4476 (N_4476,N_4120,N_4118);
nor U4477 (N_4477,N_4083,N_4084);
nand U4478 (N_4478,N_4142,N_4190);
and U4479 (N_4479,N_4041,N_4201);
nor U4480 (N_4480,N_4025,N_4154);
and U4481 (N_4481,N_4010,N_4146);
and U4482 (N_4482,N_4053,N_4034);
or U4483 (N_4483,N_4139,N_4006);
nand U4484 (N_4484,N_4124,N_4123);
xor U4485 (N_4485,N_4115,N_4160);
and U4486 (N_4486,N_4025,N_4094);
nor U4487 (N_4487,N_4130,N_4066);
nor U4488 (N_4488,N_4097,N_4140);
nand U4489 (N_4489,N_4063,N_4140);
nand U4490 (N_4490,N_4057,N_4132);
nand U4491 (N_4491,N_4130,N_4008);
nand U4492 (N_4492,N_4000,N_4043);
or U4493 (N_4493,N_4168,N_4162);
and U4494 (N_4494,N_4095,N_4213);
nor U4495 (N_4495,N_4047,N_4003);
xor U4496 (N_4496,N_4138,N_4114);
xor U4497 (N_4497,N_4068,N_4246);
nand U4498 (N_4498,N_4028,N_4082);
and U4499 (N_4499,N_4087,N_4148);
and U4500 (N_4500,N_4462,N_4445);
nand U4501 (N_4501,N_4293,N_4383);
nand U4502 (N_4502,N_4255,N_4365);
or U4503 (N_4503,N_4266,N_4295);
or U4504 (N_4504,N_4457,N_4494);
and U4505 (N_4505,N_4416,N_4375);
or U4506 (N_4506,N_4301,N_4449);
and U4507 (N_4507,N_4469,N_4444);
or U4508 (N_4508,N_4490,N_4435);
or U4509 (N_4509,N_4384,N_4361);
nor U4510 (N_4510,N_4348,N_4265);
nor U4511 (N_4511,N_4484,N_4426);
xnor U4512 (N_4512,N_4305,N_4407);
nor U4513 (N_4513,N_4474,N_4308);
or U4514 (N_4514,N_4387,N_4258);
nand U4515 (N_4515,N_4359,N_4313);
xor U4516 (N_4516,N_4456,N_4468);
nor U4517 (N_4517,N_4467,N_4296);
nand U4518 (N_4518,N_4411,N_4423);
nor U4519 (N_4519,N_4309,N_4341);
nand U4520 (N_4520,N_4323,N_4409);
xor U4521 (N_4521,N_4447,N_4488);
xnor U4522 (N_4522,N_4270,N_4406);
xnor U4523 (N_4523,N_4254,N_4472);
nor U4524 (N_4524,N_4355,N_4394);
or U4525 (N_4525,N_4385,N_4331);
and U4526 (N_4526,N_4427,N_4412);
xnor U4527 (N_4527,N_4486,N_4429);
nor U4528 (N_4528,N_4464,N_4369);
nand U4529 (N_4529,N_4317,N_4466);
nand U4530 (N_4530,N_4442,N_4451);
xnor U4531 (N_4531,N_4476,N_4298);
nand U4532 (N_4532,N_4297,N_4352);
xnor U4533 (N_4533,N_4497,N_4342);
nand U4534 (N_4534,N_4414,N_4316);
xor U4535 (N_4535,N_4358,N_4461);
nor U4536 (N_4536,N_4253,N_4366);
and U4537 (N_4537,N_4261,N_4288);
nor U4538 (N_4538,N_4275,N_4346);
nand U4539 (N_4539,N_4344,N_4438);
and U4540 (N_4540,N_4251,N_4374);
or U4541 (N_4541,N_4281,N_4264);
nand U4542 (N_4542,N_4378,N_4436);
nand U4543 (N_4543,N_4470,N_4393);
and U4544 (N_4544,N_4477,N_4340);
xnor U4545 (N_4545,N_4417,N_4455);
or U4546 (N_4546,N_4392,N_4319);
and U4547 (N_4547,N_4441,N_4397);
nand U4548 (N_4548,N_4351,N_4440);
or U4549 (N_4549,N_4424,N_4483);
nand U4550 (N_4550,N_4471,N_4345);
nand U4551 (N_4551,N_4463,N_4380);
xnor U4552 (N_4552,N_4292,N_4300);
and U4553 (N_4553,N_4303,N_4389);
xnor U4554 (N_4554,N_4492,N_4370);
xnor U4555 (N_4555,N_4386,N_4482);
nand U4556 (N_4556,N_4320,N_4291);
and U4557 (N_4557,N_4487,N_4493);
or U4558 (N_4558,N_4395,N_4491);
or U4559 (N_4559,N_4282,N_4428);
or U4560 (N_4560,N_4454,N_4294);
or U4561 (N_4561,N_4439,N_4364);
or U4562 (N_4562,N_4443,N_4408);
and U4563 (N_4563,N_4368,N_4479);
or U4564 (N_4564,N_4353,N_4419);
nor U4565 (N_4565,N_4367,N_4274);
nor U4566 (N_4566,N_4315,N_4250);
or U4567 (N_4567,N_4349,N_4286);
or U4568 (N_4568,N_4334,N_4310);
xor U4569 (N_4569,N_4262,N_4354);
and U4570 (N_4570,N_4458,N_4350);
xor U4571 (N_4571,N_4377,N_4285);
xor U4572 (N_4572,N_4321,N_4306);
and U4573 (N_4573,N_4452,N_4329);
or U4574 (N_4574,N_4421,N_4267);
and U4575 (N_4575,N_4347,N_4327);
nor U4576 (N_4576,N_4263,N_4299);
and U4577 (N_4577,N_4304,N_4257);
and U4578 (N_4578,N_4271,N_4326);
xnor U4579 (N_4579,N_4390,N_4475);
xnor U4580 (N_4580,N_4376,N_4450);
or U4581 (N_4581,N_4430,N_4337);
nor U4582 (N_4582,N_4496,N_4401);
and U4583 (N_4583,N_4318,N_4431);
xor U4584 (N_4584,N_4332,N_4307);
nor U4585 (N_4585,N_4480,N_4391);
nand U4586 (N_4586,N_4379,N_4363);
xor U4587 (N_4587,N_4432,N_4343);
or U4588 (N_4588,N_4495,N_4284);
xnor U4589 (N_4589,N_4272,N_4415);
or U4590 (N_4590,N_4252,N_4398);
and U4591 (N_4591,N_4256,N_4330);
xnor U4592 (N_4592,N_4287,N_4410);
nand U4593 (N_4593,N_4400,N_4357);
or U4594 (N_4594,N_4314,N_4312);
nor U4595 (N_4595,N_4373,N_4459);
xnor U4596 (N_4596,N_4434,N_4372);
and U4597 (N_4597,N_4362,N_4311);
nor U4598 (N_4598,N_4335,N_4290);
xor U4599 (N_4599,N_4403,N_4338);
xor U4600 (N_4600,N_4405,N_4302);
or U4601 (N_4601,N_4268,N_4473);
and U4602 (N_4602,N_4356,N_4324);
or U4603 (N_4603,N_4453,N_4498);
and U4604 (N_4604,N_4280,N_4437);
nor U4605 (N_4605,N_4260,N_4289);
nand U4606 (N_4606,N_4446,N_4399);
or U4607 (N_4607,N_4328,N_4402);
nor U4608 (N_4608,N_4413,N_4322);
and U4609 (N_4609,N_4404,N_4433);
xnor U4610 (N_4610,N_4499,N_4360);
xnor U4611 (N_4611,N_4277,N_4273);
nand U4612 (N_4612,N_4465,N_4478);
and U4613 (N_4613,N_4283,N_4259);
and U4614 (N_4614,N_4460,N_4448);
nand U4615 (N_4615,N_4279,N_4420);
nand U4616 (N_4616,N_4425,N_4396);
nand U4617 (N_4617,N_4485,N_4278);
or U4618 (N_4618,N_4276,N_4336);
nand U4619 (N_4619,N_4481,N_4325);
or U4620 (N_4620,N_4371,N_4382);
nor U4621 (N_4621,N_4388,N_4339);
xnor U4622 (N_4622,N_4422,N_4418);
or U4623 (N_4623,N_4381,N_4333);
nand U4624 (N_4624,N_4489,N_4269);
or U4625 (N_4625,N_4441,N_4257);
nor U4626 (N_4626,N_4343,N_4381);
nand U4627 (N_4627,N_4255,N_4324);
or U4628 (N_4628,N_4303,N_4337);
and U4629 (N_4629,N_4455,N_4336);
nor U4630 (N_4630,N_4301,N_4485);
and U4631 (N_4631,N_4480,N_4408);
nor U4632 (N_4632,N_4387,N_4295);
xnor U4633 (N_4633,N_4452,N_4285);
nand U4634 (N_4634,N_4469,N_4344);
nor U4635 (N_4635,N_4336,N_4473);
or U4636 (N_4636,N_4479,N_4257);
xnor U4637 (N_4637,N_4274,N_4300);
or U4638 (N_4638,N_4467,N_4460);
or U4639 (N_4639,N_4491,N_4357);
xnor U4640 (N_4640,N_4447,N_4388);
nand U4641 (N_4641,N_4362,N_4331);
nor U4642 (N_4642,N_4301,N_4434);
nand U4643 (N_4643,N_4397,N_4348);
nand U4644 (N_4644,N_4340,N_4489);
or U4645 (N_4645,N_4266,N_4448);
nand U4646 (N_4646,N_4339,N_4305);
nand U4647 (N_4647,N_4327,N_4326);
nand U4648 (N_4648,N_4319,N_4305);
and U4649 (N_4649,N_4379,N_4455);
xnor U4650 (N_4650,N_4353,N_4358);
xor U4651 (N_4651,N_4347,N_4251);
nor U4652 (N_4652,N_4371,N_4298);
or U4653 (N_4653,N_4443,N_4438);
nor U4654 (N_4654,N_4307,N_4452);
or U4655 (N_4655,N_4287,N_4487);
or U4656 (N_4656,N_4478,N_4323);
nor U4657 (N_4657,N_4262,N_4308);
and U4658 (N_4658,N_4424,N_4425);
or U4659 (N_4659,N_4301,N_4310);
nor U4660 (N_4660,N_4411,N_4447);
xnor U4661 (N_4661,N_4276,N_4375);
nand U4662 (N_4662,N_4252,N_4325);
xor U4663 (N_4663,N_4337,N_4273);
or U4664 (N_4664,N_4289,N_4378);
nor U4665 (N_4665,N_4331,N_4480);
or U4666 (N_4666,N_4392,N_4305);
or U4667 (N_4667,N_4372,N_4403);
nand U4668 (N_4668,N_4431,N_4438);
nand U4669 (N_4669,N_4374,N_4451);
nand U4670 (N_4670,N_4272,N_4285);
or U4671 (N_4671,N_4495,N_4337);
nor U4672 (N_4672,N_4286,N_4285);
or U4673 (N_4673,N_4476,N_4307);
xnor U4674 (N_4674,N_4460,N_4316);
or U4675 (N_4675,N_4313,N_4495);
nand U4676 (N_4676,N_4396,N_4428);
and U4677 (N_4677,N_4367,N_4478);
and U4678 (N_4678,N_4380,N_4462);
xnor U4679 (N_4679,N_4342,N_4435);
xnor U4680 (N_4680,N_4488,N_4368);
nor U4681 (N_4681,N_4495,N_4317);
nand U4682 (N_4682,N_4366,N_4315);
xnor U4683 (N_4683,N_4316,N_4339);
and U4684 (N_4684,N_4461,N_4302);
nand U4685 (N_4685,N_4331,N_4470);
and U4686 (N_4686,N_4302,N_4458);
and U4687 (N_4687,N_4302,N_4267);
xnor U4688 (N_4688,N_4475,N_4321);
or U4689 (N_4689,N_4293,N_4444);
and U4690 (N_4690,N_4344,N_4310);
or U4691 (N_4691,N_4498,N_4358);
nor U4692 (N_4692,N_4455,N_4442);
nor U4693 (N_4693,N_4378,N_4295);
nand U4694 (N_4694,N_4478,N_4325);
nor U4695 (N_4695,N_4435,N_4302);
or U4696 (N_4696,N_4495,N_4427);
nor U4697 (N_4697,N_4364,N_4344);
and U4698 (N_4698,N_4285,N_4379);
xor U4699 (N_4699,N_4431,N_4417);
nor U4700 (N_4700,N_4475,N_4422);
nor U4701 (N_4701,N_4346,N_4257);
and U4702 (N_4702,N_4463,N_4407);
nor U4703 (N_4703,N_4334,N_4377);
and U4704 (N_4704,N_4320,N_4352);
nor U4705 (N_4705,N_4405,N_4362);
and U4706 (N_4706,N_4350,N_4440);
and U4707 (N_4707,N_4493,N_4438);
or U4708 (N_4708,N_4314,N_4261);
nand U4709 (N_4709,N_4308,N_4298);
xnor U4710 (N_4710,N_4412,N_4430);
nor U4711 (N_4711,N_4357,N_4409);
nand U4712 (N_4712,N_4276,N_4409);
nor U4713 (N_4713,N_4257,N_4335);
nor U4714 (N_4714,N_4397,N_4256);
nand U4715 (N_4715,N_4469,N_4292);
nand U4716 (N_4716,N_4445,N_4441);
or U4717 (N_4717,N_4387,N_4450);
nand U4718 (N_4718,N_4287,N_4444);
nor U4719 (N_4719,N_4273,N_4362);
nand U4720 (N_4720,N_4483,N_4315);
and U4721 (N_4721,N_4457,N_4288);
nor U4722 (N_4722,N_4472,N_4482);
xor U4723 (N_4723,N_4432,N_4497);
nor U4724 (N_4724,N_4315,N_4364);
or U4725 (N_4725,N_4361,N_4445);
nand U4726 (N_4726,N_4429,N_4443);
xnor U4727 (N_4727,N_4416,N_4472);
nand U4728 (N_4728,N_4255,N_4303);
or U4729 (N_4729,N_4494,N_4442);
nand U4730 (N_4730,N_4347,N_4497);
nand U4731 (N_4731,N_4379,N_4402);
or U4732 (N_4732,N_4367,N_4449);
and U4733 (N_4733,N_4410,N_4331);
and U4734 (N_4734,N_4451,N_4295);
nor U4735 (N_4735,N_4256,N_4454);
nand U4736 (N_4736,N_4492,N_4399);
nor U4737 (N_4737,N_4388,N_4305);
and U4738 (N_4738,N_4269,N_4273);
and U4739 (N_4739,N_4299,N_4312);
nand U4740 (N_4740,N_4266,N_4479);
xor U4741 (N_4741,N_4362,N_4421);
nand U4742 (N_4742,N_4399,N_4467);
nor U4743 (N_4743,N_4336,N_4429);
nand U4744 (N_4744,N_4394,N_4309);
nor U4745 (N_4745,N_4266,N_4350);
or U4746 (N_4746,N_4372,N_4279);
or U4747 (N_4747,N_4366,N_4432);
nor U4748 (N_4748,N_4374,N_4279);
and U4749 (N_4749,N_4464,N_4383);
or U4750 (N_4750,N_4562,N_4731);
and U4751 (N_4751,N_4677,N_4663);
and U4752 (N_4752,N_4632,N_4588);
nand U4753 (N_4753,N_4702,N_4564);
and U4754 (N_4754,N_4749,N_4675);
and U4755 (N_4755,N_4746,N_4646);
and U4756 (N_4756,N_4537,N_4549);
and U4757 (N_4757,N_4605,N_4727);
and U4758 (N_4758,N_4643,N_4539);
and U4759 (N_4759,N_4532,N_4649);
and U4760 (N_4760,N_4715,N_4513);
nand U4761 (N_4761,N_4735,N_4680);
and U4762 (N_4762,N_4595,N_4505);
and U4763 (N_4763,N_4614,N_4504);
or U4764 (N_4764,N_4514,N_4618);
nor U4765 (N_4765,N_4623,N_4581);
nand U4766 (N_4766,N_4619,N_4544);
and U4767 (N_4767,N_4707,N_4572);
xnor U4768 (N_4768,N_4589,N_4630);
nor U4769 (N_4769,N_4660,N_4512);
nand U4770 (N_4770,N_4739,N_4701);
nand U4771 (N_4771,N_4672,N_4585);
and U4772 (N_4772,N_4538,N_4547);
nand U4773 (N_4773,N_4716,N_4552);
nand U4774 (N_4774,N_4684,N_4650);
or U4775 (N_4775,N_4615,N_4506);
or U4776 (N_4776,N_4568,N_4669);
nand U4777 (N_4777,N_4719,N_4608);
or U4778 (N_4778,N_4633,N_4690);
nand U4779 (N_4779,N_4732,N_4620);
xor U4780 (N_4780,N_4691,N_4742);
or U4781 (N_4781,N_4673,N_4535);
xnor U4782 (N_4782,N_4587,N_4703);
and U4783 (N_4783,N_4584,N_4726);
nor U4784 (N_4784,N_4668,N_4728);
or U4785 (N_4785,N_4558,N_4555);
and U4786 (N_4786,N_4529,N_4736);
or U4787 (N_4787,N_4502,N_4541);
or U4788 (N_4788,N_4725,N_4644);
nand U4789 (N_4789,N_4627,N_4700);
nor U4790 (N_4790,N_4729,N_4704);
nor U4791 (N_4791,N_4565,N_4523);
nand U4792 (N_4792,N_4510,N_4648);
nor U4793 (N_4793,N_4665,N_4718);
and U4794 (N_4794,N_4607,N_4580);
xor U4795 (N_4795,N_4666,N_4509);
or U4796 (N_4796,N_4517,N_4511);
nor U4797 (N_4797,N_4500,N_4519);
nand U4798 (N_4798,N_4503,N_4696);
xnor U4799 (N_4799,N_4651,N_4508);
nand U4800 (N_4800,N_4686,N_4685);
nor U4801 (N_4801,N_4699,N_4561);
nor U4802 (N_4802,N_4655,N_4566);
nand U4803 (N_4803,N_4583,N_4554);
or U4804 (N_4804,N_4645,N_4638);
nor U4805 (N_4805,N_4559,N_4724);
and U4806 (N_4806,N_4712,N_4659);
nand U4807 (N_4807,N_4639,N_4570);
nand U4808 (N_4808,N_4747,N_4507);
or U4809 (N_4809,N_4654,N_4676);
or U4810 (N_4810,N_4543,N_4657);
nor U4811 (N_4811,N_4625,N_4737);
and U4812 (N_4812,N_4640,N_4634);
and U4813 (N_4813,N_4629,N_4635);
or U4814 (N_4814,N_4730,N_4683);
or U4815 (N_4815,N_4600,N_4743);
nand U4816 (N_4816,N_4551,N_4530);
nor U4817 (N_4817,N_4733,N_4679);
or U4818 (N_4818,N_4597,N_4626);
nand U4819 (N_4819,N_4590,N_4674);
nor U4820 (N_4820,N_4647,N_4560);
and U4821 (N_4821,N_4671,N_4501);
nand U4822 (N_4822,N_4662,N_4661);
or U4823 (N_4823,N_4670,N_4738);
or U4824 (N_4824,N_4522,N_4722);
nor U4825 (N_4825,N_4591,N_4653);
nor U4826 (N_4826,N_4709,N_4579);
xor U4827 (N_4827,N_4598,N_4708);
and U4828 (N_4828,N_4721,N_4692);
or U4829 (N_4829,N_4693,N_4694);
or U4830 (N_4830,N_4741,N_4515);
or U4831 (N_4831,N_4536,N_4621);
or U4832 (N_4832,N_4569,N_4689);
or U4833 (N_4833,N_4631,N_4695);
and U4834 (N_4834,N_4745,N_4710);
or U4835 (N_4835,N_4534,N_4687);
and U4836 (N_4836,N_4622,N_4681);
xnor U4837 (N_4837,N_4593,N_4642);
and U4838 (N_4838,N_4556,N_4575);
and U4839 (N_4839,N_4744,N_4705);
xnor U4840 (N_4840,N_4586,N_4578);
nand U4841 (N_4841,N_4573,N_4557);
and U4842 (N_4842,N_4698,N_4518);
nand U4843 (N_4843,N_4525,N_4697);
nand U4844 (N_4844,N_4542,N_4688);
or U4845 (N_4845,N_4516,N_4599);
nor U4846 (N_4846,N_4740,N_4612);
or U4847 (N_4847,N_4611,N_4540);
nor U4848 (N_4848,N_4571,N_4616);
or U4849 (N_4849,N_4717,N_4610);
nand U4850 (N_4850,N_4577,N_4524);
or U4851 (N_4851,N_4563,N_4678);
nand U4852 (N_4852,N_4628,N_4713);
nor U4853 (N_4853,N_4636,N_4574);
nor U4854 (N_4854,N_4664,N_4613);
xnor U4855 (N_4855,N_4652,N_4720);
xor U4856 (N_4856,N_4682,N_4546);
or U4857 (N_4857,N_4528,N_4533);
nor U4858 (N_4858,N_4527,N_4601);
nand U4859 (N_4859,N_4734,N_4706);
nor U4860 (N_4860,N_4603,N_4748);
xor U4861 (N_4861,N_4596,N_4576);
xor U4862 (N_4862,N_4521,N_4550);
nor U4863 (N_4863,N_4711,N_4531);
or U4864 (N_4864,N_4567,N_4606);
xor U4865 (N_4865,N_4553,N_4617);
nand U4866 (N_4866,N_4545,N_4604);
nand U4867 (N_4867,N_4658,N_4714);
xor U4868 (N_4868,N_4723,N_4667);
and U4869 (N_4869,N_4602,N_4520);
and U4870 (N_4870,N_4582,N_4548);
xor U4871 (N_4871,N_4526,N_4624);
nand U4872 (N_4872,N_4637,N_4594);
nand U4873 (N_4873,N_4592,N_4609);
nor U4874 (N_4874,N_4641,N_4656);
and U4875 (N_4875,N_4677,N_4585);
xor U4876 (N_4876,N_4600,N_4603);
nor U4877 (N_4877,N_4551,N_4635);
nand U4878 (N_4878,N_4582,N_4704);
xor U4879 (N_4879,N_4650,N_4550);
or U4880 (N_4880,N_4699,N_4521);
and U4881 (N_4881,N_4686,N_4634);
xnor U4882 (N_4882,N_4626,N_4631);
nand U4883 (N_4883,N_4590,N_4504);
and U4884 (N_4884,N_4660,N_4616);
nor U4885 (N_4885,N_4735,N_4720);
and U4886 (N_4886,N_4681,N_4729);
nand U4887 (N_4887,N_4614,N_4645);
nand U4888 (N_4888,N_4643,N_4672);
and U4889 (N_4889,N_4509,N_4597);
nor U4890 (N_4890,N_4582,N_4589);
xor U4891 (N_4891,N_4567,N_4585);
nor U4892 (N_4892,N_4726,N_4599);
nand U4893 (N_4893,N_4689,N_4532);
nand U4894 (N_4894,N_4557,N_4615);
and U4895 (N_4895,N_4634,N_4585);
and U4896 (N_4896,N_4702,N_4746);
or U4897 (N_4897,N_4603,N_4648);
and U4898 (N_4898,N_4620,N_4645);
nor U4899 (N_4899,N_4708,N_4631);
nor U4900 (N_4900,N_4525,N_4743);
nand U4901 (N_4901,N_4616,N_4588);
and U4902 (N_4902,N_4533,N_4590);
nand U4903 (N_4903,N_4745,N_4660);
and U4904 (N_4904,N_4748,N_4720);
nor U4905 (N_4905,N_4542,N_4738);
or U4906 (N_4906,N_4568,N_4690);
or U4907 (N_4907,N_4623,N_4559);
and U4908 (N_4908,N_4539,N_4568);
and U4909 (N_4909,N_4587,N_4503);
nor U4910 (N_4910,N_4566,N_4587);
or U4911 (N_4911,N_4512,N_4645);
or U4912 (N_4912,N_4703,N_4510);
nand U4913 (N_4913,N_4584,N_4581);
xor U4914 (N_4914,N_4608,N_4522);
or U4915 (N_4915,N_4537,N_4515);
nor U4916 (N_4916,N_4746,N_4660);
nor U4917 (N_4917,N_4556,N_4704);
and U4918 (N_4918,N_4626,N_4576);
nor U4919 (N_4919,N_4515,N_4665);
nand U4920 (N_4920,N_4666,N_4589);
or U4921 (N_4921,N_4566,N_4673);
and U4922 (N_4922,N_4727,N_4656);
or U4923 (N_4923,N_4512,N_4519);
nor U4924 (N_4924,N_4502,N_4660);
nand U4925 (N_4925,N_4711,N_4726);
nor U4926 (N_4926,N_4727,N_4682);
and U4927 (N_4927,N_4741,N_4626);
and U4928 (N_4928,N_4591,N_4614);
and U4929 (N_4929,N_4651,N_4521);
or U4930 (N_4930,N_4608,N_4517);
nand U4931 (N_4931,N_4669,N_4541);
and U4932 (N_4932,N_4656,N_4702);
nor U4933 (N_4933,N_4533,N_4517);
nand U4934 (N_4934,N_4743,N_4621);
nand U4935 (N_4935,N_4536,N_4606);
and U4936 (N_4936,N_4609,N_4652);
xnor U4937 (N_4937,N_4643,N_4652);
or U4938 (N_4938,N_4659,N_4740);
and U4939 (N_4939,N_4607,N_4638);
nor U4940 (N_4940,N_4571,N_4505);
nand U4941 (N_4941,N_4504,N_4505);
xnor U4942 (N_4942,N_4680,N_4651);
or U4943 (N_4943,N_4523,N_4605);
or U4944 (N_4944,N_4541,N_4634);
and U4945 (N_4945,N_4578,N_4605);
nand U4946 (N_4946,N_4530,N_4686);
nor U4947 (N_4947,N_4533,N_4564);
xnor U4948 (N_4948,N_4528,N_4532);
nor U4949 (N_4949,N_4685,N_4711);
and U4950 (N_4950,N_4556,N_4739);
and U4951 (N_4951,N_4746,N_4569);
xor U4952 (N_4952,N_4662,N_4730);
or U4953 (N_4953,N_4643,N_4700);
nor U4954 (N_4954,N_4548,N_4697);
and U4955 (N_4955,N_4627,N_4584);
and U4956 (N_4956,N_4668,N_4603);
nand U4957 (N_4957,N_4610,N_4674);
xnor U4958 (N_4958,N_4744,N_4737);
and U4959 (N_4959,N_4655,N_4680);
or U4960 (N_4960,N_4621,N_4654);
and U4961 (N_4961,N_4629,N_4599);
or U4962 (N_4962,N_4535,N_4713);
nand U4963 (N_4963,N_4526,N_4514);
nand U4964 (N_4964,N_4500,N_4653);
and U4965 (N_4965,N_4713,N_4707);
and U4966 (N_4966,N_4610,N_4606);
xor U4967 (N_4967,N_4696,N_4635);
xnor U4968 (N_4968,N_4641,N_4588);
nand U4969 (N_4969,N_4583,N_4693);
nand U4970 (N_4970,N_4642,N_4635);
nand U4971 (N_4971,N_4510,N_4724);
and U4972 (N_4972,N_4592,N_4631);
nor U4973 (N_4973,N_4587,N_4520);
xnor U4974 (N_4974,N_4698,N_4607);
nand U4975 (N_4975,N_4669,N_4709);
nor U4976 (N_4976,N_4564,N_4628);
or U4977 (N_4977,N_4538,N_4700);
or U4978 (N_4978,N_4630,N_4676);
and U4979 (N_4979,N_4545,N_4694);
xor U4980 (N_4980,N_4664,N_4691);
nor U4981 (N_4981,N_4736,N_4624);
and U4982 (N_4982,N_4560,N_4735);
or U4983 (N_4983,N_4737,N_4705);
nor U4984 (N_4984,N_4696,N_4597);
and U4985 (N_4985,N_4660,N_4563);
nand U4986 (N_4986,N_4639,N_4626);
xnor U4987 (N_4987,N_4533,N_4550);
and U4988 (N_4988,N_4726,N_4545);
xor U4989 (N_4989,N_4572,N_4700);
nand U4990 (N_4990,N_4535,N_4666);
xnor U4991 (N_4991,N_4583,N_4513);
nor U4992 (N_4992,N_4720,N_4562);
xnor U4993 (N_4993,N_4517,N_4736);
or U4994 (N_4994,N_4730,N_4538);
nand U4995 (N_4995,N_4547,N_4623);
nand U4996 (N_4996,N_4505,N_4652);
or U4997 (N_4997,N_4603,N_4554);
nor U4998 (N_4998,N_4581,N_4556);
xnor U4999 (N_4999,N_4667,N_4742);
nand U5000 (N_5000,N_4900,N_4855);
and U5001 (N_5001,N_4933,N_4818);
nand U5002 (N_5002,N_4792,N_4778);
or U5003 (N_5003,N_4949,N_4891);
and U5004 (N_5004,N_4998,N_4753);
nand U5005 (N_5005,N_4997,N_4847);
nor U5006 (N_5006,N_4972,N_4965);
xnor U5007 (N_5007,N_4815,N_4996);
nand U5008 (N_5008,N_4786,N_4956);
and U5009 (N_5009,N_4806,N_4903);
and U5010 (N_5010,N_4751,N_4887);
nor U5011 (N_5011,N_4927,N_4993);
nor U5012 (N_5012,N_4922,N_4832);
nand U5013 (N_5013,N_4820,N_4861);
or U5014 (N_5014,N_4990,N_4950);
or U5015 (N_5015,N_4981,N_4916);
and U5016 (N_5016,N_4890,N_4945);
and U5017 (N_5017,N_4770,N_4934);
or U5018 (N_5018,N_4964,N_4906);
xnor U5019 (N_5019,N_4931,N_4938);
nor U5020 (N_5020,N_4843,N_4801);
nand U5021 (N_5021,N_4880,N_4853);
xnor U5022 (N_5022,N_4829,N_4794);
nor U5023 (N_5023,N_4932,N_4821);
nand U5024 (N_5024,N_4823,N_4805);
or U5025 (N_5025,N_4907,N_4859);
or U5026 (N_5026,N_4788,N_4873);
nor U5027 (N_5027,N_4935,N_4871);
nor U5028 (N_5028,N_4796,N_4825);
nor U5029 (N_5029,N_4937,N_4799);
and U5030 (N_5030,N_4762,N_4838);
nand U5031 (N_5031,N_4914,N_4874);
or U5032 (N_5032,N_4774,N_4798);
xor U5033 (N_5033,N_4791,N_4962);
and U5034 (N_5034,N_4894,N_4876);
and U5035 (N_5035,N_4883,N_4750);
nor U5036 (N_5036,N_4766,N_4917);
nor U5037 (N_5037,N_4979,N_4973);
xnor U5038 (N_5038,N_4863,N_4999);
nor U5039 (N_5039,N_4957,N_4837);
and U5040 (N_5040,N_4952,N_4854);
xnor U5041 (N_5041,N_4793,N_4913);
and U5042 (N_5042,N_4872,N_4982);
and U5043 (N_5043,N_4976,N_4849);
nand U5044 (N_5044,N_4761,N_4939);
and U5045 (N_5045,N_4944,N_4804);
nand U5046 (N_5046,N_4948,N_4970);
or U5047 (N_5047,N_4882,N_4810);
or U5048 (N_5048,N_4899,N_4985);
or U5049 (N_5049,N_4961,N_4988);
nor U5050 (N_5050,N_4984,N_4827);
nand U5051 (N_5051,N_4878,N_4852);
nor U5052 (N_5052,N_4756,N_4870);
and U5053 (N_5053,N_4908,N_4966);
nor U5054 (N_5054,N_4864,N_4930);
or U5055 (N_5055,N_4812,N_4809);
or U5056 (N_5056,N_4758,N_4803);
nand U5057 (N_5057,N_4919,N_4901);
nor U5058 (N_5058,N_4781,N_4974);
xor U5059 (N_5059,N_4895,N_4875);
and U5060 (N_5060,N_4869,N_4971);
and U5061 (N_5061,N_4777,N_4946);
xnor U5062 (N_5062,N_4771,N_4846);
nor U5063 (N_5063,N_4963,N_4768);
xor U5064 (N_5064,N_4765,N_4851);
xnor U5065 (N_5065,N_4835,N_4828);
xor U5066 (N_5066,N_4755,N_4896);
or U5067 (N_5067,N_4841,N_4831);
and U5068 (N_5068,N_4889,N_4764);
or U5069 (N_5069,N_4968,N_4980);
and U5070 (N_5070,N_4816,N_4780);
xnor U5071 (N_5071,N_4953,N_4858);
or U5072 (N_5072,N_4785,N_4989);
nand U5073 (N_5073,N_4884,N_4995);
or U5074 (N_5074,N_4856,N_4881);
nand U5075 (N_5075,N_4784,N_4954);
nand U5076 (N_5076,N_4915,N_4757);
nor U5077 (N_5077,N_4924,N_4942);
nand U5078 (N_5078,N_4983,N_4842);
or U5079 (N_5079,N_4789,N_4860);
xor U5080 (N_5080,N_4866,N_4886);
nor U5081 (N_5081,N_4902,N_4808);
and U5082 (N_5082,N_4822,N_4754);
and U5083 (N_5083,N_4857,N_4802);
nor U5084 (N_5084,N_4978,N_4797);
xor U5085 (N_5085,N_4830,N_4925);
nor U5086 (N_5086,N_4955,N_4824);
nand U5087 (N_5087,N_4879,N_4994);
xor U5088 (N_5088,N_4897,N_4885);
nand U5089 (N_5089,N_4819,N_4759);
xor U5090 (N_5090,N_4910,N_4840);
nor U5091 (N_5091,N_4975,N_4943);
nor U5092 (N_5092,N_4958,N_4811);
and U5093 (N_5093,N_4839,N_4772);
nand U5094 (N_5094,N_4888,N_4941);
and U5095 (N_5095,N_4905,N_4836);
or U5096 (N_5096,N_4845,N_4767);
nand U5097 (N_5097,N_4800,N_4951);
nand U5098 (N_5098,N_4928,N_4918);
xnor U5099 (N_5099,N_4834,N_4773);
nand U5100 (N_5100,N_4969,N_4790);
and U5101 (N_5101,N_4959,N_4926);
xor U5102 (N_5102,N_4904,N_4862);
nor U5103 (N_5103,N_4817,N_4769);
xor U5104 (N_5104,N_4986,N_4909);
and U5105 (N_5105,N_4987,N_4892);
nor U5106 (N_5106,N_4776,N_4833);
nand U5107 (N_5107,N_4877,N_4848);
xnor U5108 (N_5108,N_4760,N_4921);
and U5109 (N_5109,N_4936,N_4992);
and U5110 (N_5110,N_4763,N_4940);
nor U5111 (N_5111,N_4929,N_4813);
nor U5112 (N_5112,N_4865,N_4911);
nand U5113 (N_5113,N_4920,N_4850);
nand U5114 (N_5114,N_4826,N_4844);
and U5115 (N_5115,N_4947,N_4868);
nor U5116 (N_5116,N_4923,N_4960);
xnor U5117 (N_5117,N_4787,N_4967);
nand U5118 (N_5118,N_4991,N_4898);
or U5119 (N_5119,N_4893,N_4752);
nor U5120 (N_5120,N_4977,N_4807);
or U5121 (N_5121,N_4775,N_4782);
nand U5122 (N_5122,N_4783,N_4814);
xor U5123 (N_5123,N_4795,N_4912);
xor U5124 (N_5124,N_4779,N_4867);
and U5125 (N_5125,N_4823,N_4767);
and U5126 (N_5126,N_4828,N_4928);
nand U5127 (N_5127,N_4884,N_4858);
or U5128 (N_5128,N_4754,N_4951);
nor U5129 (N_5129,N_4963,N_4814);
nor U5130 (N_5130,N_4947,N_4969);
or U5131 (N_5131,N_4775,N_4819);
and U5132 (N_5132,N_4999,N_4986);
and U5133 (N_5133,N_4898,N_4767);
xor U5134 (N_5134,N_4930,N_4764);
xnor U5135 (N_5135,N_4812,N_4785);
nor U5136 (N_5136,N_4774,N_4940);
and U5137 (N_5137,N_4859,N_4994);
nand U5138 (N_5138,N_4969,N_4914);
nor U5139 (N_5139,N_4829,N_4948);
nand U5140 (N_5140,N_4850,N_4823);
nor U5141 (N_5141,N_4855,N_4758);
and U5142 (N_5142,N_4976,N_4843);
nor U5143 (N_5143,N_4905,N_4789);
nand U5144 (N_5144,N_4807,N_4848);
xnor U5145 (N_5145,N_4993,N_4948);
nand U5146 (N_5146,N_4993,N_4918);
and U5147 (N_5147,N_4880,N_4920);
nand U5148 (N_5148,N_4798,N_4871);
nand U5149 (N_5149,N_4822,N_4986);
nor U5150 (N_5150,N_4929,N_4857);
xnor U5151 (N_5151,N_4898,N_4990);
nand U5152 (N_5152,N_4948,N_4836);
xnor U5153 (N_5153,N_4834,N_4968);
and U5154 (N_5154,N_4931,N_4752);
xor U5155 (N_5155,N_4928,N_4820);
nand U5156 (N_5156,N_4838,N_4827);
and U5157 (N_5157,N_4989,N_4864);
nand U5158 (N_5158,N_4990,N_4921);
and U5159 (N_5159,N_4853,N_4958);
nand U5160 (N_5160,N_4759,N_4881);
or U5161 (N_5161,N_4910,N_4861);
nor U5162 (N_5162,N_4804,N_4891);
or U5163 (N_5163,N_4999,N_4953);
or U5164 (N_5164,N_4932,N_4790);
and U5165 (N_5165,N_4865,N_4774);
xnor U5166 (N_5166,N_4842,N_4779);
or U5167 (N_5167,N_4752,N_4769);
or U5168 (N_5168,N_4907,N_4939);
nor U5169 (N_5169,N_4798,N_4851);
and U5170 (N_5170,N_4810,N_4835);
nor U5171 (N_5171,N_4938,N_4823);
or U5172 (N_5172,N_4830,N_4961);
or U5173 (N_5173,N_4761,N_4943);
and U5174 (N_5174,N_4900,N_4807);
and U5175 (N_5175,N_4990,N_4876);
or U5176 (N_5176,N_4943,N_4951);
nor U5177 (N_5177,N_4797,N_4945);
nor U5178 (N_5178,N_4932,N_4852);
xor U5179 (N_5179,N_4996,N_4930);
or U5180 (N_5180,N_4989,N_4845);
nor U5181 (N_5181,N_4922,N_4920);
nand U5182 (N_5182,N_4902,N_4870);
and U5183 (N_5183,N_4754,N_4889);
xor U5184 (N_5184,N_4948,N_4897);
xor U5185 (N_5185,N_4887,N_4984);
and U5186 (N_5186,N_4997,N_4766);
nand U5187 (N_5187,N_4952,N_4763);
and U5188 (N_5188,N_4826,N_4828);
nor U5189 (N_5189,N_4761,N_4977);
xor U5190 (N_5190,N_4938,N_4873);
xnor U5191 (N_5191,N_4755,N_4904);
and U5192 (N_5192,N_4848,N_4964);
nand U5193 (N_5193,N_4792,N_4844);
or U5194 (N_5194,N_4871,N_4895);
or U5195 (N_5195,N_4852,N_4895);
xnor U5196 (N_5196,N_4900,N_4939);
xnor U5197 (N_5197,N_4847,N_4777);
nand U5198 (N_5198,N_4869,N_4963);
nand U5199 (N_5199,N_4867,N_4818);
xnor U5200 (N_5200,N_4785,N_4917);
nor U5201 (N_5201,N_4795,N_4926);
nand U5202 (N_5202,N_4775,N_4997);
xnor U5203 (N_5203,N_4834,N_4850);
and U5204 (N_5204,N_4976,N_4792);
nand U5205 (N_5205,N_4913,N_4863);
nor U5206 (N_5206,N_4877,N_4804);
xnor U5207 (N_5207,N_4861,N_4960);
and U5208 (N_5208,N_4899,N_4800);
nor U5209 (N_5209,N_4840,N_4985);
and U5210 (N_5210,N_4878,N_4881);
xnor U5211 (N_5211,N_4937,N_4949);
nor U5212 (N_5212,N_4774,N_4903);
or U5213 (N_5213,N_4914,N_4884);
or U5214 (N_5214,N_4835,N_4895);
or U5215 (N_5215,N_4859,N_4964);
or U5216 (N_5216,N_4760,N_4979);
or U5217 (N_5217,N_4965,N_4831);
and U5218 (N_5218,N_4963,N_4931);
nand U5219 (N_5219,N_4807,N_4936);
xnor U5220 (N_5220,N_4846,N_4860);
nor U5221 (N_5221,N_4977,N_4750);
nor U5222 (N_5222,N_4953,N_4938);
or U5223 (N_5223,N_4806,N_4935);
nor U5224 (N_5224,N_4960,N_4878);
or U5225 (N_5225,N_4785,N_4853);
and U5226 (N_5226,N_4917,N_4940);
nand U5227 (N_5227,N_4873,N_4988);
and U5228 (N_5228,N_4875,N_4865);
nand U5229 (N_5229,N_4848,N_4869);
or U5230 (N_5230,N_4937,N_4943);
nor U5231 (N_5231,N_4926,N_4998);
nand U5232 (N_5232,N_4977,N_4931);
or U5233 (N_5233,N_4838,N_4932);
nor U5234 (N_5234,N_4996,N_4825);
nand U5235 (N_5235,N_4926,N_4964);
xor U5236 (N_5236,N_4865,N_4766);
nand U5237 (N_5237,N_4805,N_4815);
or U5238 (N_5238,N_4768,N_4880);
nand U5239 (N_5239,N_4785,N_4795);
and U5240 (N_5240,N_4823,N_4997);
nor U5241 (N_5241,N_4786,N_4761);
xnor U5242 (N_5242,N_4793,N_4901);
or U5243 (N_5243,N_4927,N_4881);
nand U5244 (N_5244,N_4933,N_4913);
or U5245 (N_5245,N_4897,N_4813);
or U5246 (N_5246,N_4899,N_4960);
or U5247 (N_5247,N_4780,N_4763);
xor U5248 (N_5248,N_4807,N_4950);
or U5249 (N_5249,N_4908,N_4929);
and U5250 (N_5250,N_5047,N_5128);
nor U5251 (N_5251,N_5075,N_5023);
or U5252 (N_5252,N_5002,N_5152);
nor U5253 (N_5253,N_5151,N_5076);
nor U5254 (N_5254,N_5104,N_5086);
nand U5255 (N_5255,N_5144,N_5026);
or U5256 (N_5256,N_5099,N_5095);
nor U5257 (N_5257,N_5197,N_5078);
or U5258 (N_5258,N_5106,N_5020);
nand U5259 (N_5259,N_5246,N_5040);
nor U5260 (N_5260,N_5221,N_5156);
nor U5261 (N_5261,N_5223,N_5063);
nand U5262 (N_5262,N_5083,N_5001);
and U5263 (N_5263,N_5113,N_5174);
or U5264 (N_5264,N_5013,N_5170);
nand U5265 (N_5265,N_5178,N_5130);
nor U5266 (N_5266,N_5014,N_5089);
nand U5267 (N_5267,N_5044,N_5134);
xnor U5268 (N_5268,N_5045,N_5216);
or U5269 (N_5269,N_5176,N_5060);
nand U5270 (N_5270,N_5005,N_5175);
xnor U5271 (N_5271,N_5192,N_5240);
nor U5272 (N_5272,N_5141,N_5234);
xnor U5273 (N_5273,N_5193,N_5037);
or U5274 (N_5274,N_5015,N_5067);
nand U5275 (N_5275,N_5050,N_5027);
nand U5276 (N_5276,N_5157,N_5158);
and U5277 (N_5277,N_5231,N_5199);
nor U5278 (N_5278,N_5228,N_5055);
and U5279 (N_5279,N_5066,N_5162);
and U5280 (N_5280,N_5011,N_5181);
xor U5281 (N_5281,N_5191,N_5159);
nand U5282 (N_5282,N_5025,N_5200);
nand U5283 (N_5283,N_5125,N_5062);
nand U5284 (N_5284,N_5211,N_5115);
and U5285 (N_5285,N_5167,N_5102);
nor U5286 (N_5286,N_5189,N_5161);
xnor U5287 (N_5287,N_5173,N_5103);
or U5288 (N_5288,N_5204,N_5024);
nand U5289 (N_5289,N_5098,N_5198);
xnor U5290 (N_5290,N_5172,N_5085);
nand U5291 (N_5291,N_5114,N_5006);
and U5292 (N_5292,N_5122,N_5108);
nor U5293 (N_5293,N_5090,N_5029);
nand U5294 (N_5294,N_5057,N_5143);
nand U5295 (N_5295,N_5242,N_5069);
or U5296 (N_5296,N_5244,N_5224);
nand U5297 (N_5297,N_5051,N_5118);
nand U5298 (N_5298,N_5220,N_5196);
nor U5299 (N_5299,N_5245,N_5094);
xor U5300 (N_5300,N_5000,N_5137);
or U5301 (N_5301,N_5180,N_5046);
or U5302 (N_5302,N_5004,N_5022);
or U5303 (N_5303,N_5133,N_5146);
nor U5304 (N_5304,N_5009,N_5209);
or U5305 (N_5305,N_5032,N_5053);
and U5306 (N_5306,N_5121,N_5112);
or U5307 (N_5307,N_5003,N_5168);
xnor U5308 (N_5308,N_5230,N_5194);
or U5309 (N_5309,N_5111,N_5154);
or U5310 (N_5310,N_5235,N_5126);
or U5311 (N_5311,N_5041,N_5215);
nor U5312 (N_5312,N_5109,N_5110);
xnor U5313 (N_5313,N_5177,N_5107);
xnor U5314 (N_5314,N_5249,N_5218);
nor U5315 (N_5315,N_5092,N_5135);
nor U5316 (N_5316,N_5155,N_5219);
nand U5317 (N_5317,N_5236,N_5097);
xnor U5318 (N_5318,N_5101,N_5210);
xor U5319 (N_5319,N_5226,N_5019);
or U5320 (N_5320,N_5016,N_5012);
nand U5321 (N_5321,N_5153,N_5206);
nor U5322 (N_5322,N_5074,N_5187);
nand U5323 (N_5323,N_5018,N_5052);
nor U5324 (N_5324,N_5237,N_5140);
nand U5325 (N_5325,N_5058,N_5150);
and U5326 (N_5326,N_5208,N_5247);
nor U5327 (N_5327,N_5084,N_5127);
xor U5328 (N_5328,N_5243,N_5031);
nor U5329 (N_5329,N_5017,N_5131);
and U5330 (N_5330,N_5038,N_5179);
and U5331 (N_5331,N_5139,N_5160);
xor U5332 (N_5332,N_5182,N_5142);
nor U5333 (N_5333,N_5033,N_5233);
and U5334 (N_5334,N_5183,N_5073);
nand U5335 (N_5335,N_5105,N_5207);
xnor U5336 (N_5336,N_5056,N_5008);
nand U5337 (N_5337,N_5138,N_5071);
nand U5338 (N_5338,N_5232,N_5036);
nand U5339 (N_5339,N_5100,N_5149);
and U5340 (N_5340,N_5129,N_5093);
nand U5341 (N_5341,N_5145,N_5188);
xnor U5342 (N_5342,N_5225,N_5043);
xor U5343 (N_5343,N_5077,N_5088);
nand U5344 (N_5344,N_5068,N_5229);
nand U5345 (N_5345,N_5010,N_5238);
nor U5346 (N_5346,N_5117,N_5072);
and U5347 (N_5347,N_5214,N_5049);
xor U5348 (N_5348,N_5120,N_5201);
nor U5349 (N_5349,N_5190,N_5165);
xnor U5350 (N_5350,N_5147,N_5021);
xnor U5351 (N_5351,N_5186,N_5212);
nor U5352 (N_5352,N_5082,N_5119);
nand U5353 (N_5353,N_5169,N_5079);
or U5354 (N_5354,N_5039,N_5163);
nor U5355 (N_5355,N_5222,N_5030);
xnor U5356 (N_5356,N_5184,N_5070);
or U5357 (N_5357,N_5239,N_5061);
nor U5358 (N_5358,N_5054,N_5171);
nand U5359 (N_5359,N_5205,N_5202);
nand U5360 (N_5360,N_5064,N_5227);
or U5361 (N_5361,N_5042,N_5213);
nor U5362 (N_5362,N_5164,N_5116);
nor U5363 (N_5363,N_5132,N_5124);
and U5364 (N_5364,N_5065,N_5136);
nor U5365 (N_5365,N_5217,N_5091);
and U5366 (N_5366,N_5080,N_5096);
or U5367 (N_5367,N_5148,N_5248);
nand U5368 (N_5368,N_5081,N_5123);
and U5369 (N_5369,N_5203,N_5195);
nor U5370 (N_5370,N_5241,N_5034);
nand U5371 (N_5371,N_5087,N_5166);
or U5372 (N_5372,N_5059,N_5048);
nor U5373 (N_5373,N_5035,N_5007);
nand U5374 (N_5374,N_5028,N_5185);
or U5375 (N_5375,N_5207,N_5174);
nand U5376 (N_5376,N_5178,N_5063);
nand U5377 (N_5377,N_5094,N_5237);
xnor U5378 (N_5378,N_5219,N_5226);
or U5379 (N_5379,N_5030,N_5052);
nand U5380 (N_5380,N_5171,N_5238);
or U5381 (N_5381,N_5124,N_5080);
and U5382 (N_5382,N_5197,N_5001);
nand U5383 (N_5383,N_5222,N_5099);
xnor U5384 (N_5384,N_5113,N_5221);
and U5385 (N_5385,N_5053,N_5112);
nand U5386 (N_5386,N_5206,N_5216);
or U5387 (N_5387,N_5154,N_5121);
or U5388 (N_5388,N_5166,N_5115);
or U5389 (N_5389,N_5037,N_5020);
xor U5390 (N_5390,N_5006,N_5199);
xor U5391 (N_5391,N_5124,N_5077);
nand U5392 (N_5392,N_5177,N_5184);
or U5393 (N_5393,N_5022,N_5226);
nand U5394 (N_5394,N_5207,N_5093);
or U5395 (N_5395,N_5083,N_5234);
and U5396 (N_5396,N_5050,N_5242);
nand U5397 (N_5397,N_5041,N_5069);
nand U5398 (N_5398,N_5015,N_5001);
and U5399 (N_5399,N_5090,N_5158);
or U5400 (N_5400,N_5232,N_5229);
or U5401 (N_5401,N_5225,N_5081);
xor U5402 (N_5402,N_5090,N_5166);
nand U5403 (N_5403,N_5152,N_5201);
xnor U5404 (N_5404,N_5009,N_5024);
and U5405 (N_5405,N_5242,N_5002);
or U5406 (N_5406,N_5064,N_5010);
nor U5407 (N_5407,N_5046,N_5008);
xor U5408 (N_5408,N_5152,N_5119);
or U5409 (N_5409,N_5214,N_5006);
nand U5410 (N_5410,N_5055,N_5144);
or U5411 (N_5411,N_5005,N_5178);
nor U5412 (N_5412,N_5164,N_5159);
nand U5413 (N_5413,N_5116,N_5103);
and U5414 (N_5414,N_5035,N_5203);
or U5415 (N_5415,N_5104,N_5097);
nor U5416 (N_5416,N_5078,N_5107);
nor U5417 (N_5417,N_5103,N_5018);
nand U5418 (N_5418,N_5091,N_5077);
nand U5419 (N_5419,N_5095,N_5019);
nor U5420 (N_5420,N_5117,N_5130);
nor U5421 (N_5421,N_5085,N_5130);
xor U5422 (N_5422,N_5033,N_5061);
xor U5423 (N_5423,N_5008,N_5061);
nand U5424 (N_5424,N_5192,N_5233);
xor U5425 (N_5425,N_5103,N_5159);
or U5426 (N_5426,N_5178,N_5022);
nor U5427 (N_5427,N_5140,N_5080);
xor U5428 (N_5428,N_5142,N_5144);
nor U5429 (N_5429,N_5235,N_5211);
and U5430 (N_5430,N_5068,N_5025);
and U5431 (N_5431,N_5178,N_5236);
and U5432 (N_5432,N_5185,N_5059);
and U5433 (N_5433,N_5015,N_5111);
xor U5434 (N_5434,N_5127,N_5242);
nand U5435 (N_5435,N_5005,N_5046);
or U5436 (N_5436,N_5113,N_5018);
or U5437 (N_5437,N_5120,N_5019);
nor U5438 (N_5438,N_5125,N_5130);
or U5439 (N_5439,N_5147,N_5131);
and U5440 (N_5440,N_5042,N_5190);
and U5441 (N_5441,N_5225,N_5098);
xnor U5442 (N_5442,N_5123,N_5030);
nor U5443 (N_5443,N_5219,N_5084);
nor U5444 (N_5444,N_5163,N_5113);
and U5445 (N_5445,N_5055,N_5062);
or U5446 (N_5446,N_5215,N_5018);
nand U5447 (N_5447,N_5107,N_5057);
or U5448 (N_5448,N_5217,N_5140);
xor U5449 (N_5449,N_5034,N_5076);
or U5450 (N_5450,N_5196,N_5151);
or U5451 (N_5451,N_5139,N_5015);
or U5452 (N_5452,N_5211,N_5019);
nor U5453 (N_5453,N_5141,N_5122);
xor U5454 (N_5454,N_5034,N_5060);
or U5455 (N_5455,N_5120,N_5200);
nand U5456 (N_5456,N_5215,N_5047);
xnor U5457 (N_5457,N_5060,N_5137);
nor U5458 (N_5458,N_5104,N_5222);
and U5459 (N_5459,N_5071,N_5132);
or U5460 (N_5460,N_5069,N_5031);
nor U5461 (N_5461,N_5061,N_5126);
or U5462 (N_5462,N_5086,N_5063);
nand U5463 (N_5463,N_5009,N_5234);
or U5464 (N_5464,N_5091,N_5192);
xor U5465 (N_5465,N_5144,N_5223);
or U5466 (N_5466,N_5046,N_5187);
xnor U5467 (N_5467,N_5207,N_5230);
or U5468 (N_5468,N_5177,N_5140);
nor U5469 (N_5469,N_5018,N_5144);
nand U5470 (N_5470,N_5237,N_5083);
xnor U5471 (N_5471,N_5020,N_5099);
nand U5472 (N_5472,N_5170,N_5166);
or U5473 (N_5473,N_5068,N_5060);
and U5474 (N_5474,N_5106,N_5040);
nor U5475 (N_5475,N_5015,N_5203);
nand U5476 (N_5476,N_5015,N_5012);
and U5477 (N_5477,N_5133,N_5186);
nor U5478 (N_5478,N_5209,N_5105);
and U5479 (N_5479,N_5102,N_5010);
or U5480 (N_5480,N_5091,N_5206);
xor U5481 (N_5481,N_5180,N_5068);
nor U5482 (N_5482,N_5167,N_5112);
nor U5483 (N_5483,N_5002,N_5246);
nand U5484 (N_5484,N_5132,N_5185);
xnor U5485 (N_5485,N_5087,N_5183);
nor U5486 (N_5486,N_5049,N_5107);
or U5487 (N_5487,N_5249,N_5145);
xor U5488 (N_5488,N_5240,N_5099);
or U5489 (N_5489,N_5116,N_5125);
nor U5490 (N_5490,N_5146,N_5177);
nand U5491 (N_5491,N_5120,N_5189);
xor U5492 (N_5492,N_5233,N_5079);
or U5493 (N_5493,N_5085,N_5121);
and U5494 (N_5494,N_5058,N_5007);
and U5495 (N_5495,N_5122,N_5174);
and U5496 (N_5496,N_5148,N_5009);
or U5497 (N_5497,N_5179,N_5247);
or U5498 (N_5498,N_5076,N_5188);
or U5499 (N_5499,N_5145,N_5217);
nor U5500 (N_5500,N_5306,N_5426);
nand U5501 (N_5501,N_5366,N_5424);
or U5502 (N_5502,N_5312,N_5494);
xnor U5503 (N_5503,N_5288,N_5437);
or U5504 (N_5504,N_5328,N_5290);
nand U5505 (N_5505,N_5287,N_5415);
nor U5506 (N_5506,N_5354,N_5399);
nand U5507 (N_5507,N_5352,N_5431);
and U5508 (N_5508,N_5374,N_5335);
nor U5509 (N_5509,N_5435,N_5360);
or U5510 (N_5510,N_5417,N_5454);
and U5511 (N_5511,N_5301,N_5327);
and U5512 (N_5512,N_5363,N_5378);
and U5513 (N_5513,N_5372,N_5342);
and U5514 (N_5514,N_5331,N_5337);
nand U5515 (N_5515,N_5278,N_5376);
nand U5516 (N_5516,N_5434,N_5392);
and U5517 (N_5517,N_5279,N_5490);
nand U5518 (N_5518,N_5482,N_5457);
nor U5519 (N_5519,N_5493,N_5408);
xor U5520 (N_5520,N_5430,N_5311);
or U5521 (N_5521,N_5438,N_5496);
nor U5522 (N_5522,N_5251,N_5341);
nor U5523 (N_5523,N_5458,N_5345);
or U5524 (N_5524,N_5495,N_5465);
xor U5525 (N_5525,N_5459,N_5250);
or U5526 (N_5526,N_5257,N_5289);
and U5527 (N_5527,N_5461,N_5332);
and U5528 (N_5528,N_5292,N_5322);
or U5529 (N_5529,N_5349,N_5343);
nand U5530 (N_5530,N_5444,N_5281);
nor U5531 (N_5531,N_5375,N_5393);
or U5532 (N_5532,N_5402,N_5272);
nor U5533 (N_5533,N_5260,N_5344);
xor U5534 (N_5534,N_5284,N_5340);
xor U5535 (N_5535,N_5334,N_5268);
nor U5536 (N_5536,N_5478,N_5411);
or U5537 (N_5537,N_5455,N_5462);
nor U5538 (N_5538,N_5373,N_5333);
xnor U5539 (N_5539,N_5271,N_5368);
xor U5540 (N_5540,N_5261,N_5475);
nand U5541 (N_5541,N_5305,N_5471);
and U5542 (N_5542,N_5304,N_5394);
nand U5543 (N_5543,N_5410,N_5385);
or U5544 (N_5544,N_5254,N_5443);
xor U5545 (N_5545,N_5308,N_5329);
nand U5546 (N_5546,N_5266,N_5383);
or U5547 (N_5547,N_5314,N_5416);
xnor U5548 (N_5548,N_5379,N_5295);
and U5549 (N_5549,N_5409,N_5324);
nand U5550 (N_5550,N_5464,N_5473);
or U5551 (N_5551,N_5317,N_5357);
and U5552 (N_5552,N_5286,N_5371);
or U5553 (N_5553,N_5362,N_5369);
nand U5554 (N_5554,N_5316,N_5300);
nand U5555 (N_5555,N_5398,N_5339);
nand U5556 (N_5556,N_5282,N_5449);
and U5557 (N_5557,N_5319,N_5472);
or U5558 (N_5558,N_5309,N_5470);
nor U5559 (N_5559,N_5467,N_5386);
and U5560 (N_5560,N_5441,N_5486);
xnor U5561 (N_5561,N_5291,N_5492);
nand U5562 (N_5562,N_5361,N_5450);
or U5563 (N_5563,N_5320,N_5474);
and U5564 (N_5564,N_5407,N_5401);
nor U5565 (N_5565,N_5265,N_5321);
or U5566 (N_5566,N_5377,N_5428);
nor U5567 (N_5567,N_5405,N_5390);
xor U5568 (N_5568,N_5412,N_5294);
or U5569 (N_5569,N_5420,N_5451);
nand U5570 (N_5570,N_5421,N_5489);
nand U5571 (N_5571,N_5350,N_5269);
and U5572 (N_5572,N_5253,N_5367);
or U5573 (N_5573,N_5487,N_5358);
and U5574 (N_5574,N_5275,N_5262);
or U5575 (N_5575,N_5448,N_5387);
xnor U5576 (N_5576,N_5439,N_5452);
or U5577 (N_5577,N_5299,N_5307);
nor U5578 (N_5578,N_5480,N_5491);
xnor U5579 (N_5579,N_5395,N_5353);
or U5580 (N_5580,N_5280,N_5468);
xnor U5581 (N_5581,N_5274,N_5264);
and U5582 (N_5582,N_5263,N_5298);
nor U5583 (N_5583,N_5380,N_5302);
or U5584 (N_5584,N_5277,N_5330);
and U5585 (N_5585,N_5418,N_5419);
nand U5586 (N_5586,N_5479,N_5303);
and U5587 (N_5587,N_5283,N_5488);
nor U5588 (N_5588,N_5325,N_5436);
xnor U5589 (N_5589,N_5499,N_5469);
nor U5590 (N_5590,N_5453,N_5359);
xnor U5591 (N_5591,N_5466,N_5252);
xor U5592 (N_5592,N_5384,N_5440);
nor U5593 (N_5593,N_5422,N_5351);
and U5594 (N_5594,N_5463,N_5433);
or U5595 (N_5595,N_5397,N_5355);
or U5596 (N_5596,N_5318,N_5323);
and U5597 (N_5597,N_5313,N_5484);
or U5598 (N_5598,N_5365,N_5348);
nand U5599 (N_5599,N_5404,N_5445);
or U5600 (N_5600,N_5273,N_5364);
or U5601 (N_5601,N_5326,N_5481);
or U5602 (N_5602,N_5425,N_5276);
or U5603 (N_5603,N_5406,N_5315);
and U5604 (N_5604,N_5346,N_5270);
xnor U5605 (N_5605,N_5460,N_5356);
and U5606 (N_5606,N_5388,N_5396);
nor U5607 (N_5607,N_5400,N_5423);
nand U5608 (N_5608,N_5442,N_5447);
nor U5609 (N_5609,N_5498,N_5485);
nand U5610 (N_5610,N_5476,N_5293);
or U5611 (N_5611,N_5414,N_5285);
or U5612 (N_5612,N_5258,N_5296);
and U5613 (N_5613,N_5259,N_5370);
xor U5614 (N_5614,N_5429,N_5338);
nand U5615 (N_5615,N_5256,N_5483);
and U5616 (N_5616,N_5310,N_5446);
xnor U5617 (N_5617,N_5255,N_5432);
nor U5618 (N_5618,N_5427,N_5413);
or U5619 (N_5619,N_5297,N_5382);
xor U5620 (N_5620,N_5347,N_5391);
and U5621 (N_5621,N_5456,N_5336);
or U5622 (N_5622,N_5477,N_5381);
nand U5623 (N_5623,N_5267,N_5389);
or U5624 (N_5624,N_5497,N_5403);
xnor U5625 (N_5625,N_5465,N_5335);
nand U5626 (N_5626,N_5315,N_5367);
and U5627 (N_5627,N_5341,N_5254);
and U5628 (N_5628,N_5401,N_5434);
nor U5629 (N_5629,N_5257,N_5462);
or U5630 (N_5630,N_5374,N_5286);
or U5631 (N_5631,N_5300,N_5269);
xor U5632 (N_5632,N_5478,N_5326);
nand U5633 (N_5633,N_5396,N_5465);
nor U5634 (N_5634,N_5403,N_5383);
xnor U5635 (N_5635,N_5307,N_5422);
and U5636 (N_5636,N_5463,N_5288);
and U5637 (N_5637,N_5394,N_5297);
xor U5638 (N_5638,N_5478,N_5300);
and U5639 (N_5639,N_5403,N_5266);
and U5640 (N_5640,N_5434,N_5349);
nor U5641 (N_5641,N_5420,N_5410);
xnor U5642 (N_5642,N_5347,N_5356);
xnor U5643 (N_5643,N_5495,N_5253);
or U5644 (N_5644,N_5362,N_5441);
or U5645 (N_5645,N_5464,N_5401);
xnor U5646 (N_5646,N_5494,N_5468);
or U5647 (N_5647,N_5250,N_5315);
nand U5648 (N_5648,N_5297,N_5262);
xor U5649 (N_5649,N_5495,N_5422);
nor U5650 (N_5650,N_5419,N_5471);
nand U5651 (N_5651,N_5351,N_5392);
nand U5652 (N_5652,N_5292,N_5476);
nor U5653 (N_5653,N_5258,N_5402);
nand U5654 (N_5654,N_5259,N_5278);
nand U5655 (N_5655,N_5324,N_5261);
and U5656 (N_5656,N_5428,N_5404);
nand U5657 (N_5657,N_5334,N_5281);
nor U5658 (N_5658,N_5423,N_5366);
or U5659 (N_5659,N_5252,N_5469);
or U5660 (N_5660,N_5490,N_5336);
xor U5661 (N_5661,N_5488,N_5302);
and U5662 (N_5662,N_5330,N_5407);
and U5663 (N_5663,N_5321,N_5264);
nor U5664 (N_5664,N_5301,N_5367);
and U5665 (N_5665,N_5460,N_5296);
and U5666 (N_5666,N_5447,N_5323);
or U5667 (N_5667,N_5488,N_5498);
nand U5668 (N_5668,N_5284,N_5442);
xnor U5669 (N_5669,N_5443,N_5413);
xnor U5670 (N_5670,N_5441,N_5257);
nor U5671 (N_5671,N_5353,N_5474);
and U5672 (N_5672,N_5377,N_5325);
or U5673 (N_5673,N_5352,N_5417);
nand U5674 (N_5674,N_5400,N_5442);
nor U5675 (N_5675,N_5321,N_5335);
nor U5676 (N_5676,N_5349,N_5478);
xnor U5677 (N_5677,N_5422,N_5444);
nand U5678 (N_5678,N_5267,N_5373);
and U5679 (N_5679,N_5372,N_5258);
or U5680 (N_5680,N_5485,N_5478);
nand U5681 (N_5681,N_5313,N_5396);
xor U5682 (N_5682,N_5449,N_5371);
and U5683 (N_5683,N_5378,N_5468);
nor U5684 (N_5684,N_5308,N_5361);
nand U5685 (N_5685,N_5368,N_5293);
nor U5686 (N_5686,N_5397,N_5426);
xnor U5687 (N_5687,N_5284,N_5251);
nand U5688 (N_5688,N_5488,N_5263);
xor U5689 (N_5689,N_5478,N_5270);
nand U5690 (N_5690,N_5260,N_5294);
nand U5691 (N_5691,N_5481,N_5440);
xor U5692 (N_5692,N_5391,N_5325);
nor U5693 (N_5693,N_5253,N_5327);
and U5694 (N_5694,N_5325,N_5454);
nand U5695 (N_5695,N_5304,N_5337);
nor U5696 (N_5696,N_5347,N_5326);
xnor U5697 (N_5697,N_5277,N_5380);
and U5698 (N_5698,N_5355,N_5428);
nor U5699 (N_5699,N_5452,N_5495);
and U5700 (N_5700,N_5266,N_5329);
or U5701 (N_5701,N_5483,N_5454);
xnor U5702 (N_5702,N_5434,N_5347);
nand U5703 (N_5703,N_5285,N_5389);
nor U5704 (N_5704,N_5478,N_5359);
or U5705 (N_5705,N_5348,N_5341);
nor U5706 (N_5706,N_5413,N_5364);
xnor U5707 (N_5707,N_5428,N_5447);
nand U5708 (N_5708,N_5416,N_5406);
nor U5709 (N_5709,N_5342,N_5493);
xor U5710 (N_5710,N_5433,N_5409);
nor U5711 (N_5711,N_5312,N_5395);
and U5712 (N_5712,N_5377,N_5410);
nand U5713 (N_5713,N_5432,N_5379);
xnor U5714 (N_5714,N_5292,N_5300);
xor U5715 (N_5715,N_5298,N_5291);
nand U5716 (N_5716,N_5391,N_5256);
or U5717 (N_5717,N_5286,N_5457);
nand U5718 (N_5718,N_5325,N_5491);
and U5719 (N_5719,N_5365,N_5298);
and U5720 (N_5720,N_5393,N_5358);
or U5721 (N_5721,N_5291,N_5252);
and U5722 (N_5722,N_5330,N_5496);
or U5723 (N_5723,N_5435,N_5483);
or U5724 (N_5724,N_5438,N_5336);
nand U5725 (N_5725,N_5331,N_5390);
and U5726 (N_5726,N_5433,N_5303);
nand U5727 (N_5727,N_5430,N_5377);
xor U5728 (N_5728,N_5437,N_5314);
or U5729 (N_5729,N_5376,N_5402);
nor U5730 (N_5730,N_5452,N_5301);
or U5731 (N_5731,N_5430,N_5496);
and U5732 (N_5732,N_5261,N_5492);
and U5733 (N_5733,N_5369,N_5292);
xnor U5734 (N_5734,N_5337,N_5402);
or U5735 (N_5735,N_5317,N_5393);
xnor U5736 (N_5736,N_5311,N_5438);
or U5737 (N_5737,N_5317,N_5421);
and U5738 (N_5738,N_5461,N_5453);
xnor U5739 (N_5739,N_5351,N_5492);
xor U5740 (N_5740,N_5329,N_5293);
nand U5741 (N_5741,N_5483,N_5270);
xor U5742 (N_5742,N_5469,N_5449);
xor U5743 (N_5743,N_5363,N_5298);
nor U5744 (N_5744,N_5306,N_5449);
xnor U5745 (N_5745,N_5400,N_5282);
and U5746 (N_5746,N_5474,N_5470);
nor U5747 (N_5747,N_5398,N_5429);
nand U5748 (N_5748,N_5267,N_5416);
and U5749 (N_5749,N_5299,N_5465);
nand U5750 (N_5750,N_5563,N_5616);
xor U5751 (N_5751,N_5705,N_5622);
xnor U5752 (N_5752,N_5517,N_5644);
xor U5753 (N_5753,N_5615,N_5661);
nand U5754 (N_5754,N_5573,N_5701);
xor U5755 (N_5755,N_5691,N_5545);
xor U5756 (N_5756,N_5649,N_5733);
or U5757 (N_5757,N_5544,N_5551);
nor U5758 (N_5758,N_5596,N_5630);
nor U5759 (N_5759,N_5679,N_5654);
nand U5760 (N_5760,N_5674,N_5641);
nor U5761 (N_5761,N_5594,N_5719);
or U5762 (N_5762,N_5739,N_5666);
nor U5763 (N_5763,N_5560,N_5699);
or U5764 (N_5764,N_5547,N_5529);
xor U5765 (N_5765,N_5734,N_5528);
nand U5766 (N_5766,N_5648,N_5640);
xnor U5767 (N_5767,N_5591,N_5673);
and U5768 (N_5768,N_5526,N_5677);
and U5769 (N_5769,N_5741,N_5685);
or U5770 (N_5770,N_5680,N_5735);
xnor U5771 (N_5771,N_5682,N_5521);
or U5772 (N_5772,N_5519,N_5664);
nor U5773 (N_5773,N_5577,N_5540);
nand U5774 (N_5774,N_5610,N_5565);
xor U5775 (N_5775,N_5712,N_5711);
xnor U5776 (N_5776,N_5624,N_5738);
nand U5777 (N_5777,N_5639,N_5609);
and U5778 (N_5778,N_5554,N_5506);
nand U5779 (N_5779,N_5567,N_5709);
nor U5780 (N_5780,N_5672,N_5603);
nor U5781 (N_5781,N_5576,N_5742);
or U5782 (N_5782,N_5636,N_5692);
nor U5783 (N_5783,N_5562,N_5746);
xor U5784 (N_5784,N_5703,N_5555);
nand U5785 (N_5785,N_5611,N_5546);
nor U5786 (N_5786,N_5606,N_5516);
or U5787 (N_5787,N_5539,N_5662);
or U5788 (N_5788,N_5725,N_5524);
and U5789 (N_5789,N_5659,N_5601);
and U5790 (N_5790,N_5627,N_5513);
xnor U5791 (N_5791,N_5541,N_5665);
xor U5792 (N_5792,N_5637,N_5618);
nand U5793 (N_5793,N_5684,N_5652);
xnor U5794 (N_5794,N_5660,N_5718);
and U5795 (N_5795,N_5629,N_5512);
nand U5796 (N_5796,N_5617,N_5749);
nand U5797 (N_5797,N_5579,N_5605);
or U5798 (N_5798,N_5715,N_5503);
and U5799 (N_5799,N_5508,N_5638);
nand U5800 (N_5800,N_5504,N_5568);
or U5801 (N_5801,N_5675,N_5518);
nand U5802 (N_5802,N_5582,N_5628);
xor U5803 (N_5803,N_5595,N_5723);
nand U5804 (N_5804,N_5722,N_5710);
or U5805 (N_5805,N_5570,N_5720);
and U5806 (N_5806,N_5505,N_5693);
or U5807 (N_5807,N_5643,N_5726);
nand U5808 (N_5808,N_5621,N_5553);
or U5809 (N_5809,N_5510,N_5581);
and U5810 (N_5810,N_5729,N_5714);
and U5811 (N_5811,N_5737,N_5696);
nor U5812 (N_5812,N_5588,N_5651);
xnor U5813 (N_5813,N_5676,N_5587);
xor U5814 (N_5814,N_5658,N_5686);
xnor U5815 (N_5815,N_5566,N_5583);
nor U5816 (N_5816,N_5736,N_5557);
or U5817 (N_5817,N_5523,N_5559);
nor U5818 (N_5818,N_5704,N_5571);
and U5819 (N_5819,N_5632,N_5569);
and U5820 (N_5820,N_5647,N_5558);
and U5821 (N_5821,N_5572,N_5602);
or U5822 (N_5822,N_5697,N_5655);
or U5823 (N_5823,N_5748,N_5698);
and U5824 (N_5824,N_5713,N_5717);
xnor U5825 (N_5825,N_5620,N_5597);
nor U5826 (N_5826,N_5730,N_5598);
nand U5827 (N_5827,N_5700,N_5531);
nand U5828 (N_5828,N_5532,N_5538);
nor U5829 (N_5829,N_5599,N_5619);
xnor U5830 (N_5830,N_5515,N_5530);
xnor U5831 (N_5831,N_5653,N_5586);
nand U5832 (N_5832,N_5631,N_5716);
and U5833 (N_5833,N_5668,N_5548);
and U5834 (N_5834,N_5646,N_5642);
or U5835 (N_5835,N_5671,N_5556);
and U5836 (N_5836,N_5575,N_5625);
or U5837 (N_5837,N_5550,N_5614);
or U5838 (N_5838,N_5509,N_5501);
or U5839 (N_5839,N_5747,N_5732);
or U5840 (N_5840,N_5695,N_5689);
nand U5841 (N_5841,N_5543,N_5708);
and U5842 (N_5842,N_5633,N_5525);
and U5843 (N_5843,N_5511,N_5500);
and U5844 (N_5844,N_5650,N_5657);
or U5845 (N_5845,N_5690,N_5694);
nor U5846 (N_5846,N_5549,N_5607);
or U5847 (N_5847,N_5578,N_5635);
or U5848 (N_5848,N_5687,N_5623);
nor U5849 (N_5849,N_5592,N_5502);
xor U5850 (N_5850,N_5744,N_5706);
and U5851 (N_5851,N_5707,N_5634);
xnor U5852 (N_5852,N_5731,N_5561);
nor U5853 (N_5853,N_5537,N_5574);
or U5854 (N_5854,N_5681,N_5678);
nor U5855 (N_5855,N_5584,N_5683);
and U5856 (N_5856,N_5600,N_5663);
or U5857 (N_5857,N_5522,N_5702);
nand U5858 (N_5858,N_5589,N_5743);
xor U5859 (N_5859,N_5740,N_5721);
and U5860 (N_5860,N_5604,N_5608);
nand U5861 (N_5861,N_5527,N_5612);
nand U5862 (N_5862,N_5645,N_5520);
nand U5863 (N_5863,N_5667,N_5552);
nor U5864 (N_5864,N_5580,N_5613);
and U5865 (N_5865,N_5728,N_5533);
nand U5866 (N_5866,N_5656,N_5688);
nand U5867 (N_5867,N_5536,N_5564);
xnor U5868 (N_5868,N_5626,N_5593);
or U5869 (N_5869,N_5727,N_5534);
nand U5870 (N_5870,N_5585,N_5514);
or U5871 (N_5871,N_5507,N_5535);
xnor U5872 (N_5872,N_5669,N_5670);
or U5873 (N_5873,N_5724,N_5745);
and U5874 (N_5874,N_5590,N_5542);
xor U5875 (N_5875,N_5604,N_5502);
nor U5876 (N_5876,N_5566,N_5577);
nand U5877 (N_5877,N_5705,N_5716);
nand U5878 (N_5878,N_5501,N_5640);
xnor U5879 (N_5879,N_5593,N_5571);
nor U5880 (N_5880,N_5535,N_5545);
nand U5881 (N_5881,N_5595,N_5522);
nor U5882 (N_5882,N_5719,N_5515);
nand U5883 (N_5883,N_5510,N_5543);
nand U5884 (N_5884,N_5744,N_5523);
or U5885 (N_5885,N_5676,N_5635);
and U5886 (N_5886,N_5626,N_5611);
and U5887 (N_5887,N_5584,N_5675);
xor U5888 (N_5888,N_5719,N_5675);
xor U5889 (N_5889,N_5530,N_5740);
xor U5890 (N_5890,N_5686,N_5678);
and U5891 (N_5891,N_5669,N_5646);
and U5892 (N_5892,N_5566,N_5606);
nand U5893 (N_5893,N_5538,N_5740);
nor U5894 (N_5894,N_5689,N_5740);
nor U5895 (N_5895,N_5600,N_5554);
xor U5896 (N_5896,N_5636,N_5626);
and U5897 (N_5897,N_5519,N_5721);
nand U5898 (N_5898,N_5549,N_5542);
and U5899 (N_5899,N_5672,N_5746);
or U5900 (N_5900,N_5663,N_5612);
or U5901 (N_5901,N_5626,N_5726);
xnor U5902 (N_5902,N_5698,N_5687);
xnor U5903 (N_5903,N_5692,N_5559);
xor U5904 (N_5904,N_5598,N_5624);
or U5905 (N_5905,N_5709,N_5562);
xnor U5906 (N_5906,N_5518,N_5642);
and U5907 (N_5907,N_5723,N_5668);
and U5908 (N_5908,N_5644,N_5729);
or U5909 (N_5909,N_5503,N_5645);
xor U5910 (N_5910,N_5574,N_5630);
nor U5911 (N_5911,N_5627,N_5541);
or U5912 (N_5912,N_5635,N_5647);
and U5913 (N_5913,N_5661,N_5672);
and U5914 (N_5914,N_5714,N_5597);
xor U5915 (N_5915,N_5591,N_5643);
nand U5916 (N_5916,N_5649,N_5506);
and U5917 (N_5917,N_5711,N_5601);
nor U5918 (N_5918,N_5623,N_5630);
xor U5919 (N_5919,N_5555,N_5620);
or U5920 (N_5920,N_5618,N_5689);
xnor U5921 (N_5921,N_5538,N_5579);
or U5922 (N_5922,N_5588,N_5701);
and U5923 (N_5923,N_5548,N_5618);
nor U5924 (N_5924,N_5694,N_5721);
and U5925 (N_5925,N_5605,N_5698);
or U5926 (N_5926,N_5716,N_5516);
or U5927 (N_5927,N_5562,N_5704);
or U5928 (N_5928,N_5572,N_5584);
or U5929 (N_5929,N_5576,N_5533);
nand U5930 (N_5930,N_5567,N_5579);
and U5931 (N_5931,N_5545,N_5748);
nand U5932 (N_5932,N_5685,N_5715);
and U5933 (N_5933,N_5503,N_5544);
nand U5934 (N_5934,N_5595,N_5530);
nand U5935 (N_5935,N_5589,N_5641);
nor U5936 (N_5936,N_5564,N_5713);
or U5937 (N_5937,N_5720,N_5566);
or U5938 (N_5938,N_5640,N_5616);
or U5939 (N_5939,N_5660,N_5596);
and U5940 (N_5940,N_5531,N_5583);
nand U5941 (N_5941,N_5553,N_5716);
nor U5942 (N_5942,N_5501,N_5528);
and U5943 (N_5943,N_5706,N_5691);
and U5944 (N_5944,N_5639,N_5564);
nor U5945 (N_5945,N_5619,N_5631);
or U5946 (N_5946,N_5709,N_5561);
nand U5947 (N_5947,N_5592,N_5505);
and U5948 (N_5948,N_5599,N_5563);
and U5949 (N_5949,N_5644,N_5555);
nor U5950 (N_5950,N_5506,N_5728);
and U5951 (N_5951,N_5654,N_5636);
xnor U5952 (N_5952,N_5653,N_5583);
nor U5953 (N_5953,N_5668,N_5690);
and U5954 (N_5954,N_5605,N_5725);
nand U5955 (N_5955,N_5574,N_5504);
nor U5956 (N_5956,N_5745,N_5703);
xor U5957 (N_5957,N_5616,N_5686);
or U5958 (N_5958,N_5655,N_5508);
nand U5959 (N_5959,N_5648,N_5712);
and U5960 (N_5960,N_5674,N_5586);
or U5961 (N_5961,N_5718,N_5520);
xnor U5962 (N_5962,N_5652,N_5629);
nor U5963 (N_5963,N_5716,N_5622);
nand U5964 (N_5964,N_5515,N_5717);
or U5965 (N_5965,N_5743,N_5509);
nand U5966 (N_5966,N_5708,N_5695);
nor U5967 (N_5967,N_5590,N_5676);
xor U5968 (N_5968,N_5565,N_5698);
or U5969 (N_5969,N_5593,N_5680);
nor U5970 (N_5970,N_5689,N_5624);
nand U5971 (N_5971,N_5640,N_5741);
xor U5972 (N_5972,N_5510,N_5679);
and U5973 (N_5973,N_5669,N_5536);
nand U5974 (N_5974,N_5501,N_5604);
and U5975 (N_5975,N_5567,N_5501);
nand U5976 (N_5976,N_5673,N_5632);
and U5977 (N_5977,N_5740,N_5706);
nand U5978 (N_5978,N_5566,N_5699);
nand U5979 (N_5979,N_5514,N_5687);
nor U5980 (N_5980,N_5743,N_5710);
nor U5981 (N_5981,N_5598,N_5749);
or U5982 (N_5982,N_5584,N_5581);
and U5983 (N_5983,N_5686,N_5562);
nand U5984 (N_5984,N_5543,N_5595);
and U5985 (N_5985,N_5698,N_5663);
xor U5986 (N_5986,N_5740,N_5517);
xnor U5987 (N_5987,N_5614,N_5606);
xor U5988 (N_5988,N_5727,N_5512);
xor U5989 (N_5989,N_5680,N_5727);
nand U5990 (N_5990,N_5591,N_5692);
nor U5991 (N_5991,N_5598,N_5633);
and U5992 (N_5992,N_5542,N_5508);
nor U5993 (N_5993,N_5581,N_5619);
xnor U5994 (N_5994,N_5727,N_5515);
xnor U5995 (N_5995,N_5699,N_5660);
or U5996 (N_5996,N_5609,N_5588);
xnor U5997 (N_5997,N_5556,N_5577);
and U5998 (N_5998,N_5718,N_5606);
nand U5999 (N_5999,N_5742,N_5698);
xnor U6000 (N_6000,N_5982,N_5943);
nand U6001 (N_6001,N_5938,N_5805);
nand U6002 (N_6002,N_5911,N_5791);
xor U6003 (N_6003,N_5769,N_5903);
and U6004 (N_6004,N_5750,N_5862);
nand U6005 (N_6005,N_5870,N_5865);
xor U6006 (N_6006,N_5919,N_5797);
and U6007 (N_6007,N_5902,N_5780);
nor U6008 (N_6008,N_5840,N_5931);
xnor U6009 (N_6009,N_5951,N_5768);
nand U6010 (N_6010,N_5962,N_5846);
xor U6011 (N_6011,N_5884,N_5896);
or U6012 (N_6012,N_5762,N_5783);
nor U6013 (N_6013,N_5831,N_5756);
nor U6014 (N_6014,N_5970,N_5906);
xor U6015 (N_6015,N_5849,N_5834);
or U6016 (N_6016,N_5787,N_5880);
xor U6017 (N_6017,N_5980,N_5926);
and U6018 (N_6018,N_5814,N_5773);
xnor U6019 (N_6019,N_5810,N_5796);
xnor U6020 (N_6020,N_5795,N_5848);
nand U6021 (N_6021,N_5898,N_5835);
or U6022 (N_6022,N_5905,N_5960);
nor U6023 (N_6023,N_5789,N_5801);
and U6024 (N_6024,N_5895,N_5770);
xor U6025 (N_6025,N_5928,N_5890);
or U6026 (N_6026,N_5864,N_5759);
and U6027 (N_6027,N_5921,N_5851);
xor U6028 (N_6028,N_5843,N_5854);
nor U6029 (N_6029,N_5784,N_5983);
or U6030 (N_6030,N_5996,N_5823);
nor U6031 (N_6031,N_5836,N_5804);
xor U6032 (N_6032,N_5808,N_5965);
or U6033 (N_6033,N_5790,N_5974);
xor U6034 (N_6034,N_5859,N_5763);
nand U6035 (N_6035,N_5986,N_5907);
nor U6036 (N_6036,N_5875,N_5856);
or U6037 (N_6037,N_5803,N_5799);
nor U6038 (N_6038,N_5824,N_5954);
xor U6039 (N_6039,N_5939,N_5866);
nor U6040 (N_6040,N_5874,N_5941);
nor U6041 (N_6041,N_5963,N_5754);
and U6042 (N_6042,N_5984,N_5879);
or U6043 (N_6043,N_5959,N_5872);
nand U6044 (N_6044,N_5782,N_5764);
nor U6045 (N_6045,N_5820,N_5988);
and U6046 (N_6046,N_5881,N_5995);
xor U6047 (N_6047,N_5894,N_5839);
nand U6048 (N_6048,N_5886,N_5976);
nor U6049 (N_6049,N_5969,N_5987);
nor U6050 (N_6050,N_5767,N_5989);
and U6051 (N_6051,N_5927,N_5930);
nand U6052 (N_6052,N_5944,N_5855);
nor U6053 (N_6053,N_5934,N_5793);
and U6054 (N_6054,N_5817,N_5924);
and U6055 (N_6055,N_5788,N_5772);
and U6056 (N_6056,N_5832,N_5792);
and U6057 (N_6057,N_5913,N_5861);
xor U6058 (N_6058,N_5760,N_5920);
nand U6059 (N_6059,N_5776,N_5863);
nor U6060 (N_6060,N_5997,N_5901);
or U6061 (N_6061,N_5915,N_5957);
or U6062 (N_6062,N_5977,N_5758);
and U6063 (N_6063,N_5893,N_5829);
nor U6064 (N_6064,N_5873,N_5936);
nor U6065 (N_6065,N_5830,N_5838);
and U6066 (N_6066,N_5922,N_5892);
nor U6067 (N_6067,N_5806,N_5844);
nand U6068 (N_6068,N_5752,N_5828);
nand U6069 (N_6069,N_5949,N_5994);
xnor U6070 (N_6070,N_5751,N_5955);
xnor U6071 (N_6071,N_5785,N_5798);
or U6072 (N_6072,N_5852,N_5992);
nor U6073 (N_6073,N_5973,N_5871);
xnor U6074 (N_6074,N_5766,N_5757);
nor U6075 (N_6075,N_5860,N_5923);
and U6076 (N_6076,N_5883,N_5937);
nand U6077 (N_6077,N_5775,N_5908);
nor U6078 (N_6078,N_5858,N_5991);
nand U6079 (N_6079,N_5929,N_5825);
nand U6080 (N_6080,N_5826,N_5755);
xnor U6081 (N_6081,N_5940,N_5850);
xnor U6082 (N_6082,N_5947,N_5966);
and U6083 (N_6083,N_5972,N_5952);
xor U6084 (N_6084,N_5765,N_5794);
or U6085 (N_6085,N_5869,N_5771);
xor U6086 (N_6086,N_5916,N_5868);
nand U6087 (N_6087,N_5899,N_5802);
nor U6088 (N_6088,N_5827,N_5847);
nor U6089 (N_6089,N_5819,N_5946);
nor U6090 (N_6090,N_5807,N_5816);
and U6091 (N_6091,N_5956,N_5958);
nand U6092 (N_6092,N_5914,N_5809);
nand U6093 (N_6093,N_5778,N_5761);
nor U6094 (N_6094,N_5878,N_5837);
nor U6095 (N_6095,N_5897,N_5876);
and U6096 (N_6096,N_5910,N_5933);
nor U6097 (N_6097,N_5979,N_5800);
nor U6098 (N_6098,N_5909,N_5822);
nand U6099 (N_6099,N_5888,N_5953);
or U6100 (N_6100,N_5845,N_5912);
xor U6101 (N_6101,N_5999,N_5779);
or U6102 (N_6102,N_5900,N_5981);
and U6103 (N_6103,N_5975,N_5813);
and U6104 (N_6104,N_5998,N_5815);
nor U6105 (N_6105,N_5887,N_5971);
or U6106 (N_6106,N_5867,N_5968);
nand U6107 (N_6107,N_5853,N_5918);
nand U6108 (N_6108,N_5786,N_5993);
and U6109 (N_6109,N_5945,N_5774);
nor U6110 (N_6110,N_5857,N_5882);
or U6111 (N_6111,N_5967,N_5753);
nor U6112 (N_6112,N_5925,N_5889);
and U6113 (N_6113,N_5964,N_5904);
and U6114 (N_6114,N_5833,N_5821);
and U6115 (N_6115,N_5942,N_5811);
or U6116 (N_6116,N_5842,N_5948);
and U6117 (N_6117,N_5841,N_5932);
and U6118 (N_6118,N_5950,N_5990);
or U6119 (N_6119,N_5818,N_5885);
or U6120 (N_6120,N_5961,N_5935);
nor U6121 (N_6121,N_5877,N_5777);
xnor U6122 (N_6122,N_5781,N_5891);
xnor U6123 (N_6123,N_5917,N_5985);
or U6124 (N_6124,N_5812,N_5978);
and U6125 (N_6125,N_5806,N_5888);
xnor U6126 (N_6126,N_5988,N_5752);
nand U6127 (N_6127,N_5997,N_5787);
xor U6128 (N_6128,N_5946,N_5986);
and U6129 (N_6129,N_5908,N_5820);
or U6130 (N_6130,N_5847,N_5785);
xor U6131 (N_6131,N_5829,N_5787);
nand U6132 (N_6132,N_5894,N_5827);
and U6133 (N_6133,N_5795,N_5824);
xor U6134 (N_6134,N_5850,N_5997);
nand U6135 (N_6135,N_5962,N_5842);
nand U6136 (N_6136,N_5770,N_5944);
nor U6137 (N_6137,N_5952,N_5780);
and U6138 (N_6138,N_5852,N_5754);
xnor U6139 (N_6139,N_5868,N_5840);
or U6140 (N_6140,N_5953,N_5777);
or U6141 (N_6141,N_5873,N_5891);
and U6142 (N_6142,N_5986,N_5803);
xnor U6143 (N_6143,N_5830,N_5977);
and U6144 (N_6144,N_5805,N_5849);
xor U6145 (N_6145,N_5766,N_5754);
and U6146 (N_6146,N_5759,N_5927);
or U6147 (N_6147,N_5983,N_5944);
nand U6148 (N_6148,N_5869,N_5753);
and U6149 (N_6149,N_5938,N_5944);
nor U6150 (N_6150,N_5921,N_5819);
or U6151 (N_6151,N_5858,N_5787);
or U6152 (N_6152,N_5993,N_5778);
xnor U6153 (N_6153,N_5848,N_5861);
and U6154 (N_6154,N_5964,N_5760);
and U6155 (N_6155,N_5891,N_5949);
nand U6156 (N_6156,N_5988,N_5877);
xor U6157 (N_6157,N_5794,N_5845);
xnor U6158 (N_6158,N_5807,N_5831);
and U6159 (N_6159,N_5877,N_5959);
and U6160 (N_6160,N_5867,N_5824);
nor U6161 (N_6161,N_5907,N_5873);
and U6162 (N_6162,N_5875,N_5911);
nor U6163 (N_6163,N_5804,N_5952);
and U6164 (N_6164,N_5971,N_5836);
nand U6165 (N_6165,N_5854,N_5985);
nand U6166 (N_6166,N_5851,N_5894);
nor U6167 (N_6167,N_5857,N_5848);
and U6168 (N_6168,N_5992,N_5898);
or U6169 (N_6169,N_5876,N_5890);
xor U6170 (N_6170,N_5868,N_5874);
or U6171 (N_6171,N_5989,N_5768);
or U6172 (N_6172,N_5973,N_5909);
and U6173 (N_6173,N_5918,N_5796);
nor U6174 (N_6174,N_5797,N_5872);
and U6175 (N_6175,N_5862,N_5773);
nor U6176 (N_6176,N_5846,N_5927);
and U6177 (N_6177,N_5988,N_5768);
nor U6178 (N_6178,N_5989,N_5993);
and U6179 (N_6179,N_5885,N_5903);
or U6180 (N_6180,N_5971,N_5758);
xnor U6181 (N_6181,N_5806,N_5819);
and U6182 (N_6182,N_5776,N_5938);
or U6183 (N_6183,N_5898,N_5754);
nor U6184 (N_6184,N_5895,N_5918);
nand U6185 (N_6185,N_5757,N_5856);
nand U6186 (N_6186,N_5814,N_5900);
or U6187 (N_6187,N_5904,N_5816);
and U6188 (N_6188,N_5891,N_5870);
nor U6189 (N_6189,N_5764,N_5979);
or U6190 (N_6190,N_5808,N_5768);
nand U6191 (N_6191,N_5846,N_5837);
nand U6192 (N_6192,N_5981,N_5795);
and U6193 (N_6193,N_5798,N_5937);
xor U6194 (N_6194,N_5825,N_5955);
and U6195 (N_6195,N_5886,N_5917);
nor U6196 (N_6196,N_5919,N_5779);
nor U6197 (N_6197,N_5807,N_5893);
and U6198 (N_6198,N_5789,N_5785);
and U6199 (N_6199,N_5878,N_5822);
or U6200 (N_6200,N_5928,N_5900);
and U6201 (N_6201,N_5875,N_5892);
nor U6202 (N_6202,N_5826,N_5924);
nor U6203 (N_6203,N_5998,N_5914);
and U6204 (N_6204,N_5872,N_5854);
nor U6205 (N_6205,N_5852,N_5918);
and U6206 (N_6206,N_5854,N_5824);
and U6207 (N_6207,N_5946,N_5875);
nor U6208 (N_6208,N_5821,N_5975);
xor U6209 (N_6209,N_5984,N_5816);
xnor U6210 (N_6210,N_5982,N_5923);
and U6211 (N_6211,N_5784,N_5865);
xor U6212 (N_6212,N_5792,N_5786);
and U6213 (N_6213,N_5791,N_5923);
or U6214 (N_6214,N_5825,N_5873);
xnor U6215 (N_6215,N_5750,N_5808);
nand U6216 (N_6216,N_5921,N_5820);
xor U6217 (N_6217,N_5926,N_5960);
nor U6218 (N_6218,N_5966,N_5844);
or U6219 (N_6219,N_5947,N_5847);
or U6220 (N_6220,N_5809,N_5901);
xnor U6221 (N_6221,N_5880,N_5816);
nand U6222 (N_6222,N_5896,N_5929);
and U6223 (N_6223,N_5941,N_5775);
and U6224 (N_6224,N_5932,N_5981);
or U6225 (N_6225,N_5873,N_5957);
and U6226 (N_6226,N_5844,N_5897);
and U6227 (N_6227,N_5874,N_5806);
xnor U6228 (N_6228,N_5860,N_5833);
nor U6229 (N_6229,N_5854,N_5859);
and U6230 (N_6230,N_5977,N_5958);
and U6231 (N_6231,N_5801,N_5921);
and U6232 (N_6232,N_5984,N_5873);
or U6233 (N_6233,N_5807,N_5921);
nor U6234 (N_6234,N_5796,N_5900);
and U6235 (N_6235,N_5966,N_5881);
nand U6236 (N_6236,N_5796,N_5940);
xor U6237 (N_6237,N_5906,N_5765);
xnor U6238 (N_6238,N_5876,N_5950);
nor U6239 (N_6239,N_5905,N_5878);
or U6240 (N_6240,N_5877,N_5969);
and U6241 (N_6241,N_5764,N_5868);
nand U6242 (N_6242,N_5865,N_5889);
xor U6243 (N_6243,N_5808,N_5791);
nor U6244 (N_6244,N_5943,N_5764);
or U6245 (N_6245,N_5835,N_5901);
xnor U6246 (N_6246,N_5885,N_5948);
nand U6247 (N_6247,N_5974,N_5905);
nand U6248 (N_6248,N_5892,N_5889);
or U6249 (N_6249,N_5828,N_5764);
and U6250 (N_6250,N_6012,N_6019);
nor U6251 (N_6251,N_6029,N_6153);
and U6252 (N_6252,N_6237,N_6047);
and U6253 (N_6253,N_6089,N_6204);
and U6254 (N_6254,N_6045,N_6243);
xor U6255 (N_6255,N_6093,N_6172);
nand U6256 (N_6256,N_6130,N_6248);
xor U6257 (N_6257,N_6018,N_6081);
and U6258 (N_6258,N_6039,N_6218);
and U6259 (N_6259,N_6181,N_6139);
xor U6260 (N_6260,N_6215,N_6113);
xor U6261 (N_6261,N_6098,N_6211);
xor U6262 (N_6262,N_6168,N_6155);
nand U6263 (N_6263,N_6049,N_6239);
or U6264 (N_6264,N_6011,N_6111);
or U6265 (N_6265,N_6141,N_6222);
xnor U6266 (N_6266,N_6122,N_6182);
and U6267 (N_6267,N_6213,N_6133);
or U6268 (N_6268,N_6117,N_6107);
and U6269 (N_6269,N_6127,N_6121);
and U6270 (N_6270,N_6235,N_6000);
and U6271 (N_6271,N_6152,N_6007);
or U6272 (N_6272,N_6053,N_6052);
nor U6273 (N_6273,N_6164,N_6224);
nand U6274 (N_6274,N_6175,N_6026);
and U6275 (N_6275,N_6076,N_6203);
xnor U6276 (N_6276,N_6016,N_6171);
and U6277 (N_6277,N_6234,N_6054);
or U6278 (N_6278,N_6085,N_6071);
xnor U6279 (N_6279,N_6021,N_6233);
nand U6280 (N_6280,N_6249,N_6103);
xnor U6281 (N_6281,N_6174,N_6179);
xnor U6282 (N_6282,N_6227,N_6034);
or U6283 (N_6283,N_6009,N_6003);
nor U6284 (N_6284,N_6055,N_6166);
nor U6285 (N_6285,N_6002,N_6046);
or U6286 (N_6286,N_6013,N_6216);
nand U6287 (N_6287,N_6024,N_6092);
xor U6288 (N_6288,N_6229,N_6044);
nor U6289 (N_6289,N_6110,N_6031);
nor U6290 (N_6290,N_6244,N_6058);
nand U6291 (N_6291,N_6005,N_6167);
xnor U6292 (N_6292,N_6095,N_6064);
and U6293 (N_6293,N_6069,N_6073);
and U6294 (N_6294,N_6143,N_6232);
or U6295 (N_6295,N_6096,N_6083);
and U6296 (N_6296,N_6017,N_6150);
or U6297 (N_6297,N_6060,N_6192);
or U6298 (N_6298,N_6033,N_6230);
nand U6299 (N_6299,N_6180,N_6038);
xnor U6300 (N_6300,N_6135,N_6209);
nand U6301 (N_6301,N_6170,N_6032);
or U6302 (N_6302,N_6221,N_6189);
nor U6303 (N_6303,N_6236,N_6088);
xnor U6304 (N_6304,N_6157,N_6128);
or U6305 (N_6305,N_6188,N_6240);
or U6306 (N_6306,N_6165,N_6140);
nor U6307 (N_6307,N_6138,N_6154);
and U6308 (N_6308,N_6100,N_6015);
nand U6309 (N_6309,N_6147,N_6195);
xnor U6310 (N_6310,N_6020,N_6190);
nand U6311 (N_6311,N_6050,N_6087);
xnor U6312 (N_6312,N_6099,N_6148);
nand U6313 (N_6313,N_6177,N_6028);
nor U6314 (N_6314,N_6187,N_6207);
nor U6315 (N_6315,N_6160,N_6198);
nand U6316 (N_6316,N_6059,N_6109);
nand U6317 (N_6317,N_6014,N_6191);
nand U6318 (N_6318,N_6072,N_6084);
nand U6319 (N_6319,N_6242,N_6194);
nand U6320 (N_6320,N_6205,N_6238);
or U6321 (N_6321,N_6066,N_6115);
xor U6322 (N_6322,N_6144,N_6217);
or U6323 (N_6323,N_6247,N_6094);
nor U6324 (N_6324,N_6105,N_6136);
nor U6325 (N_6325,N_6199,N_6056);
nor U6326 (N_6326,N_6036,N_6041);
xnor U6327 (N_6327,N_6178,N_6151);
or U6328 (N_6328,N_6075,N_6163);
and U6329 (N_6329,N_6022,N_6101);
and U6330 (N_6330,N_6008,N_6065);
xor U6331 (N_6331,N_6048,N_6082);
and U6332 (N_6332,N_6061,N_6131);
and U6333 (N_6333,N_6196,N_6219);
or U6334 (N_6334,N_6074,N_6201);
and U6335 (N_6335,N_6057,N_6116);
xor U6336 (N_6336,N_6183,N_6037);
nor U6337 (N_6337,N_6118,N_6114);
nor U6338 (N_6338,N_6120,N_6210);
nor U6339 (N_6339,N_6202,N_6173);
nand U6340 (N_6340,N_6208,N_6245);
and U6341 (N_6341,N_6241,N_6156);
xnor U6342 (N_6342,N_6067,N_6169);
nand U6343 (N_6343,N_6125,N_6142);
and U6344 (N_6344,N_6004,N_6193);
or U6345 (N_6345,N_6112,N_6104);
xor U6346 (N_6346,N_6042,N_6124);
nand U6347 (N_6347,N_6158,N_6149);
xor U6348 (N_6348,N_6030,N_6079);
or U6349 (N_6349,N_6080,N_6223);
or U6350 (N_6350,N_6126,N_6228);
xor U6351 (N_6351,N_6051,N_6123);
or U6352 (N_6352,N_6159,N_6226);
nor U6353 (N_6353,N_6097,N_6197);
and U6354 (N_6354,N_6129,N_6220);
nor U6355 (N_6355,N_6134,N_6090);
nand U6356 (N_6356,N_6027,N_6186);
or U6357 (N_6357,N_6162,N_6001);
or U6358 (N_6358,N_6212,N_6206);
nand U6359 (N_6359,N_6078,N_6108);
nand U6360 (N_6360,N_6185,N_6010);
nor U6361 (N_6361,N_6132,N_6086);
and U6362 (N_6362,N_6035,N_6062);
nand U6363 (N_6363,N_6246,N_6070);
and U6364 (N_6364,N_6145,N_6023);
nand U6365 (N_6365,N_6063,N_6091);
or U6366 (N_6366,N_6040,N_6068);
xor U6367 (N_6367,N_6102,N_6225);
nand U6368 (N_6368,N_6214,N_6025);
or U6369 (N_6369,N_6137,N_6231);
and U6370 (N_6370,N_6200,N_6106);
xor U6371 (N_6371,N_6146,N_6077);
and U6372 (N_6372,N_6043,N_6184);
or U6373 (N_6373,N_6006,N_6176);
nand U6374 (N_6374,N_6161,N_6119);
and U6375 (N_6375,N_6132,N_6179);
or U6376 (N_6376,N_6170,N_6080);
or U6377 (N_6377,N_6085,N_6104);
and U6378 (N_6378,N_6058,N_6156);
nand U6379 (N_6379,N_6046,N_6066);
nand U6380 (N_6380,N_6057,N_6121);
xor U6381 (N_6381,N_6073,N_6121);
nand U6382 (N_6382,N_6160,N_6212);
or U6383 (N_6383,N_6091,N_6179);
nor U6384 (N_6384,N_6219,N_6238);
xor U6385 (N_6385,N_6222,N_6159);
and U6386 (N_6386,N_6079,N_6231);
or U6387 (N_6387,N_6068,N_6157);
xnor U6388 (N_6388,N_6050,N_6237);
nor U6389 (N_6389,N_6135,N_6029);
nor U6390 (N_6390,N_6192,N_6131);
xnor U6391 (N_6391,N_6052,N_6092);
and U6392 (N_6392,N_6020,N_6186);
xor U6393 (N_6393,N_6191,N_6021);
nor U6394 (N_6394,N_6133,N_6037);
nand U6395 (N_6395,N_6051,N_6043);
xor U6396 (N_6396,N_6061,N_6102);
xnor U6397 (N_6397,N_6122,N_6188);
xor U6398 (N_6398,N_6180,N_6139);
nor U6399 (N_6399,N_6004,N_6024);
nand U6400 (N_6400,N_6128,N_6048);
or U6401 (N_6401,N_6204,N_6100);
and U6402 (N_6402,N_6236,N_6094);
nor U6403 (N_6403,N_6191,N_6241);
nand U6404 (N_6404,N_6098,N_6104);
nor U6405 (N_6405,N_6066,N_6093);
or U6406 (N_6406,N_6118,N_6048);
and U6407 (N_6407,N_6119,N_6199);
and U6408 (N_6408,N_6146,N_6162);
and U6409 (N_6409,N_6108,N_6021);
xnor U6410 (N_6410,N_6086,N_6012);
nand U6411 (N_6411,N_6135,N_6030);
or U6412 (N_6412,N_6146,N_6158);
or U6413 (N_6413,N_6159,N_6073);
and U6414 (N_6414,N_6017,N_6020);
nand U6415 (N_6415,N_6126,N_6111);
and U6416 (N_6416,N_6185,N_6056);
nor U6417 (N_6417,N_6048,N_6045);
nand U6418 (N_6418,N_6147,N_6064);
or U6419 (N_6419,N_6066,N_6174);
nor U6420 (N_6420,N_6131,N_6005);
or U6421 (N_6421,N_6078,N_6066);
nor U6422 (N_6422,N_6105,N_6172);
or U6423 (N_6423,N_6244,N_6069);
xor U6424 (N_6424,N_6020,N_6181);
and U6425 (N_6425,N_6098,N_6197);
and U6426 (N_6426,N_6118,N_6220);
nor U6427 (N_6427,N_6220,N_6151);
or U6428 (N_6428,N_6071,N_6028);
and U6429 (N_6429,N_6100,N_6098);
or U6430 (N_6430,N_6239,N_6179);
or U6431 (N_6431,N_6150,N_6065);
nand U6432 (N_6432,N_6233,N_6095);
and U6433 (N_6433,N_6064,N_6123);
xor U6434 (N_6434,N_6147,N_6123);
xnor U6435 (N_6435,N_6241,N_6150);
nand U6436 (N_6436,N_6113,N_6238);
and U6437 (N_6437,N_6048,N_6134);
nor U6438 (N_6438,N_6194,N_6107);
nor U6439 (N_6439,N_6234,N_6224);
or U6440 (N_6440,N_6242,N_6206);
nor U6441 (N_6441,N_6143,N_6028);
or U6442 (N_6442,N_6085,N_6054);
nor U6443 (N_6443,N_6201,N_6129);
xnor U6444 (N_6444,N_6020,N_6059);
and U6445 (N_6445,N_6207,N_6191);
xor U6446 (N_6446,N_6169,N_6154);
nand U6447 (N_6447,N_6029,N_6240);
and U6448 (N_6448,N_6248,N_6145);
or U6449 (N_6449,N_6139,N_6152);
xnor U6450 (N_6450,N_6103,N_6091);
or U6451 (N_6451,N_6209,N_6139);
xor U6452 (N_6452,N_6092,N_6145);
nand U6453 (N_6453,N_6015,N_6138);
nand U6454 (N_6454,N_6240,N_6171);
nand U6455 (N_6455,N_6077,N_6083);
or U6456 (N_6456,N_6191,N_6164);
and U6457 (N_6457,N_6116,N_6202);
nor U6458 (N_6458,N_6102,N_6249);
xor U6459 (N_6459,N_6235,N_6146);
nor U6460 (N_6460,N_6091,N_6112);
nand U6461 (N_6461,N_6196,N_6072);
xor U6462 (N_6462,N_6238,N_6228);
or U6463 (N_6463,N_6002,N_6059);
nor U6464 (N_6464,N_6218,N_6093);
xor U6465 (N_6465,N_6030,N_6144);
and U6466 (N_6466,N_6110,N_6227);
or U6467 (N_6467,N_6099,N_6196);
xor U6468 (N_6468,N_6158,N_6231);
nand U6469 (N_6469,N_6231,N_6092);
or U6470 (N_6470,N_6248,N_6091);
or U6471 (N_6471,N_6155,N_6015);
xor U6472 (N_6472,N_6245,N_6190);
nand U6473 (N_6473,N_6020,N_6225);
nand U6474 (N_6474,N_6181,N_6210);
and U6475 (N_6475,N_6117,N_6032);
nor U6476 (N_6476,N_6226,N_6084);
xnor U6477 (N_6477,N_6187,N_6184);
xor U6478 (N_6478,N_6102,N_6083);
nand U6479 (N_6479,N_6171,N_6208);
xor U6480 (N_6480,N_6202,N_6073);
nand U6481 (N_6481,N_6074,N_6206);
xor U6482 (N_6482,N_6048,N_6092);
nor U6483 (N_6483,N_6050,N_6098);
nand U6484 (N_6484,N_6015,N_6197);
nor U6485 (N_6485,N_6009,N_6142);
nor U6486 (N_6486,N_6026,N_6048);
xor U6487 (N_6487,N_6158,N_6028);
and U6488 (N_6488,N_6093,N_6054);
nor U6489 (N_6489,N_6024,N_6206);
or U6490 (N_6490,N_6084,N_6204);
nor U6491 (N_6491,N_6184,N_6076);
or U6492 (N_6492,N_6167,N_6122);
nor U6493 (N_6493,N_6039,N_6238);
and U6494 (N_6494,N_6031,N_6039);
and U6495 (N_6495,N_6050,N_6052);
xnor U6496 (N_6496,N_6196,N_6248);
or U6497 (N_6497,N_6186,N_6177);
and U6498 (N_6498,N_6015,N_6135);
nand U6499 (N_6499,N_6105,N_6209);
nand U6500 (N_6500,N_6418,N_6273);
xor U6501 (N_6501,N_6319,N_6308);
and U6502 (N_6502,N_6453,N_6457);
nor U6503 (N_6503,N_6439,N_6278);
nand U6504 (N_6504,N_6482,N_6369);
or U6505 (N_6505,N_6326,N_6262);
nand U6506 (N_6506,N_6277,N_6303);
nand U6507 (N_6507,N_6324,N_6259);
and U6508 (N_6508,N_6325,N_6318);
nor U6509 (N_6509,N_6497,N_6274);
nand U6510 (N_6510,N_6357,N_6291);
or U6511 (N_6511,N_6394,N_6359);
nand U6512 (N_6512,N_6282,N_6292);
nor U6513 (N_6513,N_6299,N_6470);
xnor U6514 (N_6514,N_6434,N_6267);
and U6515 (N_6515,N_6428,N_6341);
nor U6516 (N_6516,N_6388,N_6493);
and U6517 (N_6517,N_6446,N_6281);
or U6518 (N_6518,N_6414,N_6276);
nand U6519 (N_6519,N_6403,N_6264);
or U6520 (N_6520,N_6279,N_6290);
nor U6521 (N_6521,N_6419,N_6476);
and U6522 (N_6522,N_6438,N_6338);
and U6523 (N_6523,N_6286,N_6288);
nor U6524 (N_6524,N_6367,N_6484);
nand U6525 (N_6525,N_6390,N_6408);
and U6526 (N_6526,N_6306,N_6405);
nor U6527 (N_6527,N_6348,N_6268);
xor U6528 (N_6528,N_6435,N_6342);
and U6529 (N_6529,N_6383,N_6284);
nand U6530 (N_6530,N_6416,N_6368);
or U6531 (N_6531,N_6411,N_6373);
xor U6532 (N_6532,N_6429,N_6463);
xnor U6533 (N_6533,N_6381,N_6328);
nor U6534 (N_6534,N_6472,N_6375);
and U6535 (N_6535,N_6442,N_6420);
nand U6536 (N_6536,N_6445,N_6321);
xor U6537 (N_6537,N_6467,N_6289);
xor U6538 (N_6538,N_6491,N_6461);
nand U6539 (N_6539,N_6360,N_6347);
and U6540 (N_6540,N_6330,N_6479);
nor U6541 (N_6541,N_6363,N_6293);
or U6542 (N_6542,N_6280,N_6270);
nor U6543 (N_6543,N_6496,N_6258);
nand U6544 (N_6544,N_6460,N_6317);
or U6545 (N_6545,N_6409,N_6404);
nor U6546 (N_6546,N_6354,N_6402);
or U6547 (N_6547,N_6473,N_6331);
nand U6548 (N_6548,N_6349,N_6393);
or U6549 (N_6549,N_6353,N_6287);
nand U6550 (N_6550,N_6485,N_6492);
nor U6551 (N_6551,N_6335,N_6454);
nand U6552 (N_6552,N_6415,N_6423);
nand U6553 (N_6553,N_6437,N_6456);
nor U6554 (N_6554,N_6487,N_6351);
nand U6555 (N_6555,N_6465,N_6451);
xnor U6556 (N_6556,N_6378,N_6413);
nor U6557 (N_6557,N_6361,N_6436);
and U6558 (N_6558,N_6260,N_6355);
and U6559 (N_6559,N_6311,N_6275);
or U6560 (N_6560,N_6327,N_6300);
nor U6561 (N_6561,N_6251,N_6455);
nand U6562 (N_6562,N_6417,N_6399);
nor U6563 (N_6563,N_6400,N_6332);
nand U6564 (N_6564,N_6298,N_6489);
xor U6565 (N_6565,N_6462,N_6395);
xnor U6566 (N_6566,N_6379,N_6250);
or U6567 (N_6567,N_6407,N_6449);
or U6568 (N_6568,N_6350,N_6406);
or U6569 (N_6569,N_6252,N_6385);
xor U6570 (N_6570,N_6310,N_6261);
nor U6571 (N_6571,N_6488,N_6444);
nor U6572 (N_6572,N_6297,N_6458);
or U6573 (N_6573,N_6358,N_6422);
xor U6574 (N_6574,N_6468,N_6471);
nor U6575 (N_6575,N_6389,N_6499);
nor U6576 (N_6576,N_6432,N_6441);
nor U6577 (N_6577,N_6486,N_6380);
and U6578 (N_6578,N_6431,N_6448);
and U6579 (N_6579,N_6440,N_6314);
or U6580 (N_6580,N_6301,N_6313);
nand U6581 (N_6581,N_6447,N_6309);
nor U6582 (N_6582,N_6427,N_6329);
or U6583 (N_6583,N_6269,N_6307);
nor U6584 (N_6584,N_6315,N_6304);
nor U6585 (N_6585,N_6294,N_6494);
and U6586 (N_6586,N_6425,N_6316);
nor U6587 (N_6587,N_6257,N_6424);
and U6588 (N_6588,N_6362,N_6433);
xnor U6589 (N_6589,N_6356,N_6334);
xnor U6590 (N_6590,N_6272,N_6474);
nand U6591 (N_6591,N_6323,N_6490);
xnor U6592 (N_6592,N_6495,N_6285);
and U6593 (N_6593,N_6450,N_6343);
nor U6594 (N_6594,N_6475,N_6478);
nor U6595 (N_6595,N_6371,N_6265);
or U6596 (N_6596,N_6466,N_6372);
nand U6597 (N_6597,N_6421,N_6254);
nand U6598 (N_6598,N_6430,N_6426);
xnor U6599 (N_6599,N_6255,N_6412);
and U6600 (N_6600,N_6480,N_6365);
xor U6601 (N_6601,N_6370,N_6401);
and U6602 (N_6602,N_6392,N_6443);
and U6603 (N_6603,N_6333,N_6377);
nor U6604 (N_6604,N_6398,N_6459);
nand U6605 (N_6605,N_6391,N_6481);
nand U6606 (N_6606,N_6305,N_6410);
nand U6607 (N_6607,N_6376,N_6464);
xor U6608 (N_6608,N_6374,N_6253);
nand U6609 (N_6609,N_6336,N_6295);
or U6610 (N_6610,N_6344,N_6322);
and U6611 (N_6611,N_6366,N_6345);
nand U6612 (N_6612,N_6498,N_6271);
nand U6613 (N_6613,N_6387,N_6256);
or U6614 (N_6614,N_6320,N_6312);
or U6615 (N_6615,N_6452,N_6396);
nand U6616 (N_6616,N_6337,N_6296);
nor U6617 (N_6617,N_6346,N_6302);
or U6618 (N_6618,N_6384,N_6469);
xor U6619 (N_6619,N_6397,N_6283);
nand U6620 (N_6620,N_6483,N_6386);
and U6621 (N_6621,N_6340,N_6339);
xor U6622 (N_6622,N_6364,N_6477);
and U6623 (N_6623,N_6352,N_6382);
and U6624 (N_6624,N_6263,N_6266);
or U6625 (N_6625,N_6342,N_6348);
nand U6626 (N_6626,N_6423,N_6404);
xor U6627 (N_6627,N_6495,N_6251);
and U6628 (N_6628,N_6392,N_6389);
nand U6629 (N_6629,N_6260,N_6432);
xnor U6630 (N_6630,N_6302,N_6476);
and U6631 (N_6631,N_6473,N_6365);
and U6632 (N_6632,N_6268,N_6264);
and U6633 (N_6633,N_6428,N_6463);
nor U6634 (N_6634,N_6455,N_6264);
xor U6635 (N_6635,N_6378,N_6497);
and U6636 (N_6636,N_6298,N_6439);
or U6637 (N_6637,N_6269,N_6427);
nand U6638 (N_6638,N_6375,N_6292);
nor U6639 (N_6639,N_6413,N_6437);
nor U6640 (N_6640,N_6405,N_6382);
nand U6641 (N_6641,N_6341,N_6330);
nand U6642 (N_6642,N_6334,N_6369);
nand U6643 (N_6643,N_6498,N_6407);
nand U6644 (N_6644,N_6302,N_6390);
or U6645 (N_6645,N_6398,N_6382);
or U6646 (N_6646,N_6482,N_6360);
or U6647 (N_6647,N_6355,N_6499);
nand U6648 (N_6648,N_6423,N_6439);
nand U6649 (N_6649,N_6431,N_6474);
and U6650 (N_6650,N_6454,N_6281);
nor U6651 (N_6651,N_6338,N_6369);
or U6652 (N_6652,N_6366,N_6319);
nand U6653 (N_6653,N_6478,N_6427);
or U6654 (N_6654,N_6295,N_6414);
xor U6655 (N_6655,N_6350,N_6458);
nor U6656 (N_6656,N_6364,N_6339);
or U6657 (N_6657,N_6470,N_6255);
nand U6658 (N_6658,N_6362,N_6440);
and U6659 (N_6659,N_6282,N_6459);
and U6660 (N_6660,N_6427,N_6469);
nor U6661 (N_6661,N_6351,N_6344);
or U6662 (N_6662,N_6360,N_6487);
or U6663 (N_6663,N_6395,N_6352);
nor U6664 (N_6664,N_6259,N_6376);
xor U6665 (N_6665,N_6482,N_6341);
or U6666 (N_6666,N_6252,N_6456);
or U6667 (N_6667,N_6406,N_6354);
xor U6668 (N_6668,N_6434,N_6407);
nand U6669 (N_6669,N_6333,N_6356);
nor U6670 (N_6670,N_6406,N_6473);
and U6671 (N_6671,N_6307,N_6361);
nor U6672 (N_6672,N_6255,N_6275);
xnor U6673 (N_6673,N_6375,N_6282);
xor U6674 (N_6674,N_6455,N_6307);
and U6675 (N_6675,N_6480,N_6351);
xnor U6676 (N_6676,N_6458,N_6331);
xor U6677 (N_6677,N_6452,N_6317);
nor U6678 (N_6678,N_6480,N_6471);
and U6679 (N_6679,N_6302,N_6376);
xor U6680 (N_6680,N_6418,N_6371);
nor U6681 (N_6681,N_6477,N_6394);
or U6682 (N_6682,N_6293,N_6388);
or U6683 (N_6683,N_6339,N_6336);
nand U6684 (N_6684,N_6302,N_6339);
or U6685 (N_6685,N_6326,N_6309);
nand U6686 (N_6686,N_6397,N_6294);
xnor U6687 (N_6687,N_6396,N_6422);
xor U6688 (N_6688,N_6439,N_6352);
nand U6689 (N_6689,N_6456,N_6473);
and U6690 (N_6690,N_6281,N_6337);
nor U6691 (N_6691,N_6461,N_6372);
xor U6692 (N_6692,N_6331,N_6469);
and U6693 (N_6693,N_6401,N_6373);
xnor U6694 (N_6694,N_6323,N_6362);
and U6695 (N_6695,N_6464,N_6487);
nand U6696 (N_6696,N_6443,N_6486);
nand U6697 (N_6697,N_6367,N_6401);
nand U6698 (N_6698,N_6317,N_6487);
nor U6699 (N_6699,N_6421,N_6298);
xnor U6700 (N_6700,N_6381,N_6392);
and U6701 (N_6701,N_6424,N_6353);
or U6702 (N_6702,N_6273,N_6451);
nand U6703 (N_6703,N_6481,N_6436);
nor U6704 (N_6704,N_6415,N_6438);
and U6705 (N_6705,N_6259,N_6347);
xor U6706 (N_6706,N_6370,N_6493);
nor U6707 (N_6707,N_6393,N_6354);
nor U6708 (N_6708,N_6434,N_6328);
nor U6709 (N_6709,N_6337,N_6408);
nor U6710 (N_6710,N_6423,N_6459);
nor U6711 (N_6711,N_6314,N_6391);
nand U6712 (N_6712,N_6480,N_6459);
nor U6713 (N_6713,N_6380,N_6455);
xnor U6714 (N_6714,N_6471,N_6372);
xor U6715 (N_6715,N_6437,N_6285);
and U6716 (N_6716,N_6428,N_6447);
nor U6717 (N_6717,N_6328,N_6266);
xnor U6718 (N_6718,N_6478,N_6470);
or U6719 (N_6719,N_6443,N_6339);
nand U6720 (N_6720,N_6335,N_6375);
nor U6721 (N_6721,N_6468,N_6411);
and U6722 (N_6722,N_6265,N_6470);
xnor U6723 (N_6723,N_6288,N_6293);
nor U6724 (N_6724,N_6395,N_6386);
nand U6725 (N_6725,N_6286,N_6337);
xor U6726 (N_6726,N_6433,N_6282);
or U6727 (N_6727,N_6477,N_6254);
nor U6728 (N_6728,N_6398,N_6421);
or U6729 (N_6729,N_6334,N_6252);
and U6730 (N_6730,N_6465,N_6425);
nor U6731 (N_6731,N_6346,N_6366);
nand U6732 (N_6732,N_6320,N_6324);
xnor U6733 (N_6733,N_6318,N_6286);
nor U6734 (N_6734,N_6309,N_6438);
nor U6735 (N_6735,N_6346,N_6258);
xnor U6736 (N_6736,N_6394,N_6436);
or U6737 (N_6737,N_6288,N_6285);
and U6738 (N_6738,N_6407,N_6466);
or U6739 (N_6739,N_6475,N_6491);
nand U6740 (N_6740,N_6462,N_6385);
and U6741 (N_6741,N_6292,N_6278);
or U6742 (N_6742,N_6364,N_6408);
nand U6743 (N_6743,N_6359,N_6357);
or U6744 (N_6744,N_6262,N_6450);
nor U6745 (N_6745,N_6429,N_6273);
xor U6746 (N_6746,N_6411,N_6347);
xnor U6747 (N_6747,N_6368,N_6336);
nor U6748 (N_6748,N_6295,N_6318);
nand U6749 (N_6749,N_6438,N_6412);
nand U6750 (N_6750,N_6654,N_6521);
nor U6751 (N_6751,N_6526,N_6597);
xnor U6752 (N_6752,N_6665,N_6505);
nand U6753 (N_6753,N_6596,N_6686);
or U6754 (N_6754,N_6554,N_6538);
nand U6755 (N_6755,N_6507,N_6684);
or U6756 (N_6756,N_6715,N_6666);
xnor U6757 (N_6757,N_6524,N_6748);
or U6758 (N_6758,N_6576,N_6571);
and U6759 (N_6759,N_6713,N_6503);
and U6760 (N_6760,N_6557,N_6618);
or U6761 (N_6761,N_6559,N_6721);
nand U6762 (N_6762,N_6731,N_6511);
xnor U6763 (N_6763,N_6560,N_6533);
nand U6764 (N_6764,N_6670,N_6709);
xnor U6765 (N_6765,N_6569,N_6616);
xor U6766 (N_6766,N_6733,N_6699);
or U6767 (N_6767,N_6728,N_6707);
xnor U6768 (N_6768,N_6630,N_6712);
nor U6769 (N_6769,N_6517,N_6673);
nand U6770 (N_6770,N_6520,N_6703);
or U6771 (N_6771,N_6598,N_6678);
nand U6772 (N_6772,N_6603,N_6690);
xor U6773 (N_6773,N_6551,N_6504);
nor U6774 (N_6774,N_6529,N_6716);
and U6775 (N_6775,N_6581,N_6516);
and U6776 (N_6776,N_6510,N_6661);
xnor U6777 (N_6777,N_6591,N_6519);
nor U6778 (N_6778,N_6633,N_6583);
or U6779 (N_6779,N_6656,N_6550);
nor U6780 (N_6780,N_6558,N_6736);
and U6781 (N_6781,N_6555,N_6547);
and U6782 (N_6782,N_6613,N_6682);
and U6783 (N_6783,N_6602,N_6582);
nand U6784 (N_6784,N_6626,N_6553);
nand U6785 (N_6785,N_6607,N_6535);
and U6786 (N_6786,N_6580,N_6635);
xor U6787 (N_6787,N_6672,N_6515);
nor U6788 (N_6788,N_6500,N_6564);
nand U6789 (N_6789,N_6586,N_6737);
nor U6790 (N_6790,N_6649,N_6563);
nand U6791 (N_6791,N_6698,N_6729);
nand U6792 (N_6792,N_6567,N_6530);
xnor U6793 (N_6793,N_6719,N_6681);
nand U6794 (N_6794,N_6548,N_6735);
and U6795 (N_6795,N_6701,N_6573);
or U6796 (N_6796,N_6639,N_6549);
or U6797 (N_6797,N_6585,N_6696);
and U6798 (N_6798,N_6627,N_6726);
and U6799 (N_6799,N_6722,N_6570);
or U6800 (N_6800,N_6502,N_6657);
xor U6801 (N_6801,N_6568,N_6590);
xor U6802 (N_6802,N_6695,N_6704);
and U6803 (N_6803,N_6727,N_6501);
xor U6804 (N_6804,N_6622,N_6741);
nor U6805 (N_6805,N_6718,N_6592);
and U6806 (N_6806,N_6546,N_6599);
nor U6807 (N_6807,N_6668,N_6506);
nor U6808 (N_6808,N_6691,N_6653);
nor U6809 (N_6809,N_6562,N_6700);
xor U6810 (N_6810,N_6534,N_6739);
and U6811 (N_6811,N_6693,N_6525);
and U6812 (N_6812,N_6683,N_6615);
nand U6813 (N_6813,N_6646,N_6740);
nor U6814 (N_6814,N_6685,N_6614);
xor U6815 (N_6815,N_6565,N_6621);
nor U6816 (N_6816,N_6705,N_6694);
or U6817 (N_6817,N_6634,N_6746);
nor U6818 (N_6818,N_6522,N_6644);
or U6819 (N_6819,N_6664,N_6566);
and U6820 (N_6820,N_6648,N_6514);
nand U6821 (N_6821,N_6528,N_6738);
nand U6822 (N_6822,N_6620,N_6730);
xor U6823 (N_6823,N_6625,N_6636);
xor U6824 (N_6824,N_6629,N_6643);
nand U6825 (N_6825,N_6542,N_6674);
xor U6826 (N_6826,N_6710,N_6641);
xnor U6827 (N_6827,N_6556,N_6611);
and U6828 (N_6828,N_6714,N_6536);
nor U6829 (N_6829,N_6688,N_6584);
xnor U6830 (N_6830,N_6608,N_6539);
or U6831 (N_6831,N_6744,N_6660);
and U6832 (N_6832,N_6575,N_6724);
and U6833 (N_6833,N_6663,N_6662);
xnor U6834 (N_6834,N_6631,N_6655);
and U6835 (N_6835,N_6689,N_6747);
nor U6836 (N_6836,N_6692,N_6745);
or U6837 (N_6837,N_6593,N_6523);
or U6838 (N_6838,N_6638,N_6509);
xnor U6839 (N_6839,N_6652,N_6679);
xor U6840 (N_6840,N_6601,N_6561);
and U6841 (N_6841,N_6669,N_6732);
nand U6842 (N_6842,N_6574,N_6609);
nand U6843 (N_6843,N_6720,N_6612);
xnor U6844 (N_6844,N_6617,N_6702);
xor U6845 (N_6845,N_6658,N_6578);
and U6846 (N_6846,N_6645,N_6659);
or U6847 (N_6847,N_6640,N_6650);
nor U6848 (N_6848,N_6513,N_6637);
or U6849 (N_6849,N_6734,N_6532);
and U6850 (N_6850,N_6541,N_6687);
nand U6851 (N_6851,N_6671,N_6537);
and U6852 (N_6852,N_6579,N_6743);
nand U6853 (N_6853,N_6647,N_6706);
nand U6854 (N_6854,N_6606,N_6708);
nor U6855 (N_6855,N_6605,N_6623);
nand U6856 (N_6856,N_6600,N_6676);
or U6857 (N_6857,N_6723,N_6572);
or U6858 (N_6858,N_6711,N_6749);
or U6859 (N_6859,N_6589,N_6552);
nand U6860 (N_6860,N_6531,N_6508);
nor U6861 (N_6861,N_6624,N_6651);
xor U6862 (N_6862,N_6540,N_6697);
or U6863 (N_6863,N_6610,N_6545);
or U6864 (N_6864,N_6642,N_6742);
xnor U6865 (N_6865,N_6725,N_6604);
nand U6866 (N_6866,N_6667,N_6675);
nor U6867 (N_6867,N_6588,N_6680);
nand U6868 (N_6868,N_6632,N_6677);
or U6869 (N_6869,N_6594,N_6619);
and U6870 (N_6870,N_6527,N_6544);
or U6871 (N_6871,N_6628,N_6587);
and U6872 (N_6872,N_6717,N_6512);
or U6873 (N_6873,N_6595,N_6543);
and U6874 (N_6874,N_6577,N_6518);
nor U6875 (N_6875,N_6664,N_6722);
xor U6876 (N_6876,N_6632,N_6500);
nor U6877 (N_6877,N_6652,N_6620);
xnor U6878 (N_6878,N_6565,N_6576);
or U6879 (N_6879,N_6530,N_6549);
nor U6880 (N_6880,N_6524,N_6702);
xnor U6881 (N_6881,N_6536,N_6506);
or U6882 (N_6882,N_6568,N_6678);
xor U6883 (N_6883,N_6522,N_6550);
and U6884 (N_6884,N_6562,N_6728);
and U6885 (N_6885,N_6625,N_6546);
nor U6886 (N_6886,N_6710,N_6690);
nor U6887 (N_6887,N_6552,N_6646);
xnor U6888 (N_6888,N_6669,N_6508);
xnor U6889 (N_6889,N_6657,N_6654);
xor U6890 (N_6890,N_6611,N_6538);
or U6891 (N_6891,N_6696,N_6617);
and U6892 (N_6892,N_6680,N_6667);
nand U6893 (N_6893,N_6557,N_6520);
or U6894 (N_6894,N_6553,N_6673);
nor U6895 (N_6895,N_6745,N_6577);
or U6896 (N_6896,N_6543,N_6502);
nand U6897 (N_6897,N_6563,N_6688);
nor U6898 (N_6898,N_6514,N_6529);
xnor U6899 (N_6899,N_6735,N_6672);
nand U6900 (N_6900,N_6678,N_6654);
nand U6901 (N_6901,N_6540,N_6597);
nor U6902 (N_6902,N_6620,N_6539);
nand U6903 (N_6903,N_6654,N_6666);
or U6904 (N_6904,N_6665,N_6675);
xnor U6905 (N_6905,N_6599,N_6721);
or U6906 (N_6906,N_6520,N_6675);
nor U6907 (N_6907,N_6592,N_6681);
and U6908 (N_6908,N_6706,N_6613);
and U6909 (N_6909,N_6713,N_6542);
nand U6910 (N_6910,N_6645,N_6670);
and U6911 (N_6911,N_6595,N_6743);
xor U6912 (N_6912,N_6677,N_6537);
xnor U6913 (N_6913,N_6685,N_6572);
or U6914 (N_6914,N_6713,N_6700);
nor U6915 (N_6915,N_6530,N_6732);
and U6916 (N_6916,N_6529,N_6580);
and U6917 (N_6917,N_6672,N_6599);
nor U6918 (N_6918,N_6553,N_6663);
nand U6919 (N_6919,N_6695,N_6647);
nand U6920 (N_6920,N_6728,N_6717);
or U6921 (N_6921,N_6551,N_6653);
or U6922 (N_6922,N_6744,N_6557);
nor U6923 (N_6923,N_6605,N_6749);
or U6924 (N_6924,N_6653,N_6593);
and U6925 (N_6925,N_6620,N_6607);
nor U6926 (N_6926,N_6605,N_6741);
xor U6927 (N_6927,N_6707,N_6562);
or U6928 (N_6928,N_6569,N_6706);
and U6929 (N_6929,N_6689,N_6526);
xnor U6930 (N_6930,N_6596,N_6520);
nor U6931 (N_6931,N_6738,N_6509);
xnor U6932 (N_6932,N_6581,N_6574);
nand U6933 (N_6933,N_6737,N_6645);
xor U6934 (N_6934,N_6631,N_6729);
or U6935 (N_6935,N_6535,N_6579);
xor U6936 (N_6936,N_6689,N_6609);
nand U6937 (N_6937,N_6727,N_6649);
xor U6938 (N_6938,N_6636,N_6556);
and U6939 (N_6939,N_6554,N_6694);
and U6940 (N_6940,N_6648,N_6703);
nand U6941 (N_6941,N_6565,N_6641);
xor U6942 (N_6942,N_6587,N_6675);
and U6943 (N_6943,N_6632,N_6703);
nand U6944 (N_6944,N_6634,N_6718);
and U6945 (N_6945,N_6604,N_6663);
nor U6946 (N_6946,N_6556,N_6664);
nand U6947 (N_6947,N_6525,N_6629);
xnor U6948 (N_6948,N_6740,N_6608);
nand U6949 (N_6949,N_6730,N_6714);
nor U6950 (N_6950,N_6693,N_6593);
or U6951 (N_6951,N_6525,N_6617);
xnor U6952 (N_6952,N_6651,N_6697);
nor U6953 (N_6953,N_6601,N_6566);
xor U6954 (N_6954,N_6612,N_6576);
nand U6955 (N_6955,N_6720,N_6619);
or U6956 (N_6956,N_6565,N_6595);
or U6957 (N_6957,N_6507,N_6563);
xnor U6958 (N_6958,N_6638,N_6690);
xor U6959 (N_6959,N_6654,N_6615);
nand U6960 (N_6960,N_6683,N_6647);
or U6961 (N_6961,N_6700,N_6711);
and U6962 (N_6962,N_6553,N_6606);
or U6963 (N_6963,N_6749,N_6592);
and U6964 (N_6964,N_6565,N_6626);
and U6965 (N_6965,N_6603,N_6517);
nand U6966 (N_6966,N_6617,N_6503);
xor U6967 (N_6967,N_6747,N_6745);
and U6968 (N_6968,N_6591,N_6737);
and U6969 (N_6969,N_6718,N_6667);
nand U6970 (N_6970,N_6700,N_6620);
and U6971 (N_6971,N_6534,N_6514);
and U6972 (N_6972,N_6529,N_6685);
xor U6973 (N_6973,N_6575,N_6597);
nor U6974 (N_6974,N_6517,N_6534);
and U6975 (N_6975,N_6684,N_6602);
xor U6976 (N_6976,N_6678,N_6666);
nor U6977 (N_6977,N_6530,N_6512);
nand U6978 (N_6978,N_6592,N_6600);
nand U6979 (N_6979,N_6720,N_6635);
and U6980 (N_6980,N_6511,N_6569);
xor U6981 (N_6981,N_6661,N_6736);
xor U6982 (N_6982,N_6644,N_6737);
nand U6983 (N_6983,N_6694,N_6745);
nand U6984 (N_6984,N_6684,N_6594);
and U6985 (N_6985,N_6683,N_6731);
nand U6986 (N_6986,N_6587,N_6520);
or U6987 (N_6987,N_6606,N_6537);
nand U6988 (N_6988,N_6574,N_6535);
nand U6989 (N_6989,N_6669,N_6657);
xor U6990 (N_6990,N_6631,N_6567);
xnor U6991 (N_6991,N_6593,N_6540);
and U6992 (N_6992,N_6575,N_6593);
xnor U6993 (N_6993,N_6715,N_6603);
nand U6994 (N_6994,N_6667,N_6714);
nand U6995 (N_6995,N_6732,N_6646);
or U6996 (N_6996,N_6621,N_6709);
nor U6997 (N_6997,N_6748,N_6554);
or U6998 (N_6998,N_6533,N_6684);
nor U6999 (N_6999,N_6722,N_6658);
nand U7000 (N_7000,N_6871,N_6924);
and U7001 (N_7001,N_6760,N_6930);
nor U7002 (N_7002,N_6759,N_6864);
and U7003 (N_7003,N_6913,N_6780);
and U7004 (N_7004,N_6878,N_6763);
or U7005 (N_7005,N_6807,N_6781);
or U7006 (N_7006,N_6921,N_6764);
xnor U7007 (N_7007,N_6882,N_6755);
nor U7008 (N_7008,N_6783,N_6842);
nand U7009 (N_7009,N_6946,N_6787);
or U7010 (N_7010,N_6928,N_6961);
nor U7011 (N_7011,N_6937,N_6959);
and U7012 (N_7012,N_6813,N_6750);
and U7013 (N_7013,N_6756,N_6911);
and U7014 (N_7014,N_6980,N_6817);
nand U7015 (N_7015,N_6904,N_6966);
and U7016 (N_7016,N_6843,N_6892);
nand U7017 (N_7017,N_6977,N_6916);
or U7018 (N_7018,N_6891,N_6808);
nand U7019 (N_7019,N_6989,N_6987);
nand U7020 (N_7020,N_6971,N_6877);
or U7021 (N_7021,N_6872,N_6758);
or U7022 (N_7022,N_6988,N_6975);
xnor U7023 (N_7023,N_6947,N_6887);
nand U7024 (N_7024,N_6833,N_6849);
xor U7025 (N_7025,N_6770,N_6810);
nand U7026 (N_7026,N_6983,N_6950);
nor U7027 (N_7027,N_6753,N_6830);
nor U7028 (N_7028,N_6822,N_6796);
and U7029 (N_7029,N_6772,N_6968);
xnor U7030 (N_7030,N_6957,N_6844);
nand U7031 (N_7031,N_6859,N_6899);
and U7032 (N_7032,N_6826,N_6841);
nand U7033 (N_7033,N_6769,N_6814);
xnor U7034 (N_7034,N_6985,N_6963);
nor U7035 (N_7035,N_6976,N_6934);
or U7036 (N_7036,N_6837,N_6867);
nor U7037 (N_7037,N_6936,N_6835);
or U7038 (N_7038,N_6854,N_6779);
nand U7039 (N_7039,N_6846,N_6893);
or U7040 (N_7040,N_6803,N_6902);
or U7041 (N_7041,N_6776,N_6819);
or U7042 (N_7042,N_6940,N_6986);
and U7043 (N_7043,N_6852,N_6990);
nand U7044 (N_7044,N_6836,N_6838);
nand U7045 (N_7045,N_6935,N_6782);
xnor U7046 (N_7046,N_6840,N_6905);
xnor U7047 (N_7047,N_6876,N_6806);
or U7048 (N_7048,N_6839,N_6973);
xor U7049 (N_7049,N_6785,N_6927);
nand U7050 (N_7050,N_6829,N_6820);
xnor U7051 (N_7051,N_6944,N_6922);
or U7052 (N_7052,N_6997,N_6790);
nand U7053 (N_7053,N_6926,N_6943);
xnor U7054 (N_7054,N_6789,N_6875);
and U7055 (N_7055,N_6910,N_6920);
and U7056 (N_7056,N_6828,N_6885);
nor U7057 (N_7057,N_6821,N_6898);
or U7058 (N_7058,N_6856,N_6824);
and U7059 (N_7059,N_6771,N_6804);
and U7060 (N_7060,N_6952,N_6886);
and U7061 (N_7061,N_6906,N_6884);
or U7062 (N_7062,N_6818,N_6994);
nor U7063 (N_7063,N_6917,N_6979);
or U7064 (N_7064,N_6896,N_6919);
and U7065 (N_7065,N_6786,N_6880);
xnor U7066 (N_7066,N_6784,N_6909);
nor U7067 (N_7067,N_6802,N_6809);
nand U7068 (N_7068,N_6866,N_6811);
xnor U7069 (N_7069,N_6815,N_6895);
and U7070 (N_7070,N_6834,N_6951);
nor U7071 (N_7071,N_6982,N_6861);
nor U7072 (N_7072,N_6868,N_6949);
or U7073 (N_7073,N_6778,N_6775);
nor U7074 (N_7074,N_6956,N_6967);
xnor U7075 (N_7075,N_6974,N_6798);
nand U7076 (N_7076,N_6825,N_6845);
nor U7077 (N_7077,N_6761,N_6894);
or U7078 (N_7078,N_6766,N_6797);
nand U7079 (N_7079,N_6816,N_6873);
nor U7080 (N_7080,N_6751,N_6870);
xor U7081 (N_7081,N_6792,N_6860);
and U7082 (N_7082,N_6931,N_6794);
nand U7083 (N_7083,N_6903,N_6991);
or U7084 (N_7084,N_6865,N_6915);
or U7085 (N_7085,N_6869,N_6752);
xnor U7086 (N_7086,N_6942,N_6890);
or U7087 (N_7087,N_6847,N_6901);
nand U7088 (N_7088,N_6939,N_6960);
or U7089 (N_7089,N_6791,N_6969);
nor U7090 (N_7090,N_6984,N_6900);
nor U7091 (N_7091,N_6879,N_6954);
xnor U7092 (N_7092,N_6858,N_6805);
nor U7093 (N_7093,N_6995,N_6765);
or U7094 (N_7094,N_6889,N_6981);
or U7095 (N_7095,N_6998,N_6812);
nor U7096 (N_7096,N_6918,N_6863);
nand U7097 (N_7097,N_6774,N_6970);
nor U7098 (N_7098,N_6757,N_6881);
nor U7099 (N_7099,N_6754,N_6912);
nor U7100 (N_7100,N_6925,N_6965);
nor U7101 (N_7101,N_6762,N_6848);
nor U7102 (N_7102,N_6888,N_6862);
nor U7103 (N_7103,N_6923,N_6823);
nand U7104 (N_7104,N_6831,N_6768);
and U7105 (N_7105,N_6874,N_6941);
xor U7106 (N_7106,N_6972,N_6958);
nor U7107 (N_7107,N_6799,N_6999);
and U7108 (N_7108,N_6945,N_6851);
and U7109 (N_7109,N_6948,N_6777);
nand U7110 (N_7110,N_6933,N_6914);
nor U7111 (N_7111,N_6793,N_6907);
and U7112 (N_7112,N_6801,N_6855);
nor U7113 (N_7113,N_6853,N_6832);
nand U7114 (N_7114,N_6827,N_6767);
or U7115 (N_7115,N_6932,N_6788);
nor U7116 (N_7116,N_6850,N_6964);
or U7117 (N_7117,N_6857,N_6929);
xnor U7118 (N_7118,N_6795,N_6996);
or U7119 (N_7119,N_6883,N_6908);
or U7120 (N_7120,N_6955,N_6938);
or U7121 (N_7121,N_6993,N_6953);
xor U7122 (N_7122,N_6962,N_6897);
nor U7123 (N_7123,N_6800,N_6992);
nand U7124 (N_7124,N_6773,N_6978);
nand U7125 (N_7125,N_6975,N_6799);
nand U7126 (N_7126,N_6916,N_6907);
or U7127 (N_7127,N_6997,N_6833);
nand U7128 (N_7128,N_6811,N_6883);
xnor U7129 (N_7129,N_6890,N_6760);
nor U7130 (N_7130,N_6995,N_6968);
nand U7131 (N_7131,N_6970,N_6938);
xor U7132 (N_7132,N_6949,N_6809);
or U7133 (N_7133,N_6832,N_6816);
and U7134 (N_7134,N_6859,N_6949);
or U7135 (N_7135,N_6973,N_6934);
xnor U7136 (N_7136,N_6840,N_6978);
or U7137 (N_7137,N_6893,N_6932);
xor U7138 (N_7138,N_6899,N_6933);
xor U7139 (N_7139,N_6790,N_6988);
nand U7140 (N_7140,N_6956,N_6998);
nand U7141 (N_7141,N_6784,N_6928);
and U7142 (N_7142,N_6845,N_6762);
xnor U7143 (N_7143,N_6812,N_6785);
or U7144 (N_7144,N_6913,N_6993);
nand U7145 (N_7145,N_6750,N_6913);
or U7146 (N_7146,N_6834,N_6877);
xor U7147 (N_7147,N_6960,N_6980);
and U7148 (N_7148,N_6917,N_6974);
nor U7149 (N_7149,N_6760,N_6753);
or U7150 (N_7150,N_6836,N_6958);
nor U7151 (N_7151,N_6881,N_6867);
or U7152 (N_7152,N_6888,N_6925);
nand U7153 (N_7153,N_6981,N_6827);
nor U7154 (N_7154,N_6908,N_6769);
nor U7155 (N_7155,N_6842,N_6864);
nand U7156 (N_7156,N_6868,N_6974);
xor U7157 (N_7157,N_6925,N_6805);
nor U7158 (N_7158,N_6850,N_6982);
or U7159 (N_7159,N_6941,N_6869);
and U7160 (N_7160,N_6883,N_6982);
or U7161 (N_7161,N_6773,N_6952);
nand U7162 (N_7162,N_6800,N_6964);
and U7163 (N_7163,N_6973,N_6791);
and U7164 (N_7164,N_6766,N_6862);
or U7165 (N_7165,N_6886,N_6859);
nand U7166 (N_7166,N_6994,N_6990);
xnor U7167 (N_7167,N_6807,N_6803);
and U7168 (N_7168,N_6890,N_6951);
xor U7169 (N_7169,N_6798,N_6970);
or U7170 (N_7170,N_6900,N_6991);
or U7171 (N_7171,N_6959,N_6877);
nand U7172 (N_7172,N_6872,N_6898);
nand U7173 (N_7173,N_6932,N_6926);
xnor U7174 (N_7174,N_6802,N_6998);
nor U7175 (N_7175,N_6761,N_6980);
nand U7176 (N_7176,N_6992,N_6856);
or U7177 (N_7177,N_6839,N_6901);
nand U7178 (N_7178,N_6941,N_6876);
or U7179 (N_7179,N_6832,N_6964);
nand U7180 (N_7180,N_6803,N_6857);
nand U7181 (N_7181,N_6814,N_6919);
or U7182 (N_7182,N_6872,N_6851);
xor U7183 (N_7183,N_6949,N_6927);
nand U7184 (N_7184,N_6969,N_6787);
or U7185 (N_7185,N_6860,N_6871);
or U7186 (N_7186,N_6976,N_6984);
nand U7187 (N_7187,N_6959,N_6983);
or U7188 (N_7188,N_6770,N_6871);
and U7189 (N_7189,N_6862,N_6934);
nand U7190 (N_7190,N_6854,N_6759);
or U7191 (N_7191,N_6876,N_6865);
nand U7192 (N_7192,N_6755,N_6786);
nor U7193 (N_7193,N_6859,N_6771);
nor U7194 (N_7194,N_6923,N_6941);
xnor U7195 (N_7195,N_6763,N_6781);
nor U7196 (N_7196,N_6906,N_6793);
xnor U7197 (N_7197,N_6886,N_6860);
xnor U7198 (N_7198,N_6773,N_6788);
nor U7199 (N_7199,N_6876,N_6898);
and U7200 (N_7200,N_6976,N_6928);
nor U7201 (N_7201,N_6829,N_6871);
or U7202 (N_7202,N_6968,N_6752);
xor U7203 (N_7203,N_6948,N_6874);
nor U7204 (N_7204,N_6877,N_6763);
nand U7205 (N_7205,N_6881,N_6802);
nand U7206 (N_7206,N_6899,N_6921);
and U7207 (N_7207,N_6922,N_6900);
and U7208 (N_7208,N_6774,N_6844);
xor U7209 (N_7209,N_6905,N_6967);
or U7210 (N_7210,N_6968,N_6813);
and U7211 (N_7211,N_6962,N_6929);
xnor U7212 (N_7212,N_6806,N_6751);
xnor U7213 (N_7213,N_6818,N_6976);
xnor U7214 (N_7214,N_6912,N_6944);
nand U7215 (N_7215,N_6801,N_6847);
nor U7216 (N_7216,N_6988,N_6876);
and U7217 (N_7217,N_6849,N_6975);
or U7218 (N_7218,N_6987,N_6976);
and U7219 (N_7219,N_6962,N_6966);
or U7220 (N_7220,N_6806,N_6836);
nor U7221 (N_7221,N_6977,N_6847);
and U7222 (N_7222,N_6969,N_6929);
nor U7223 (N_7223,N_6914,N_6926);
nor U7224 (N_7224,N_6950,N_6958);
and U7225 (N_7225,N_6754,N_6965);
or U7226 (N_7226,N_6964,N_6973);
and U7227 (N_7227,N_6840,N_6798);
nor U7228 (N_7228,N_6940,N_6774);
nand U7229 (N_7229,N_6990,N_6808);
nor U7230 (N_7230,N_6887,N_6897);
and U7231 (N_7231,N_6942,N_6782);
xnor U7232 (N_7232,N_6850,N_6825);
nor U7233 (N_7233,N_6814,N_6886);
or U7234 (N_7234,N_6939,N_6830);
xnor U7235 (N_7235,N_6772,N_6901);
xnor U7236 (N_7236,N_6834,N_6843);
nor U7237 (N_7237,N_6901,N_6852);
or U7238 (N_7238,N_6830,N_6768);
or U7239 (N_7239,N_6994,N_6914);
or U7240 (N_7240,N_6857,N_6860);
xnor U7241 (N_7241,N_6876,N_6792);
or U7242 (N_7242,N_6976,N_6825);
xnor U7243 (N_7243,N_6810,N_6934);
or U7244 (N_7244,N_6778,N_6945);
and U7245 (N_7245,N_6760,N_6789);
and U7246 (N_7246,N_6912,N_6932);
nor U7247 (N_7247,N_6985,N_6968);
and U7248 (N_7248,N_6911,N_6796);
or U7249 (N_7249,N_6954,N_6930);
nand U7250 (N_7250,N_7193,N_7004);
xnor U7251 (N_7251,N_7035,N_7039);
nor U7252 (N_7252,N_7204,N_7061);
nor U7253 (N_7253,N_7132,N_7099);
xor U7254 (N_7254,N_7086,N_7164);
nor U7255 (N_7255,N_7066,N_7108);
and U7256 (N_7256,N_7024,N_7122);
nand U7257 (N_7257,N_7022,N_7196);
or U7258 (N_7258,N_7092,N_7127);
nor U7259 (N_7259,N_7232,N_7080);
nand U7260 (N_7260,N_7000,N_7117);
nor U7261 (N_7261,N_7089,N_7074);
or U7262 (N_7262,N_7013,N_7238);
xnor U7263 (N_7263,N_7111,N_7212);
nor U7264 (N_7264,N_7175,N_7206);
xnor U7265 (N_7265,N_7056,N_7069);
nor U7266 (N_7266,N_7156,N_7170);
or U7267 (N_7267,N_7037,N_7222);
xnor U7268 (N_7268,N_7186,N_7101);
and U7269 (N_7269,N_7058,N_7046);
nand U7270 (N_7270,N_7059,N_7043);
and U7271 (N_7271,N_7041,N_7235);
and U7272 (N_7272,N_7153,N_7189);
or U7273 (N_7273,N_7230,N_7019);
and U7274 (N_7274,N_7241,N_7246);
nor U7275 (N_7275,N_7050,N_7068);
xnor U7276 (N_7276,N_7105,N_7221);
nor U7277 (N_7277,N_7154,N_7025);
nand U7278 (N_7278,N_7021,N_7178);
nand U7279 (N_7279,N_7208,N_7147);
xnor U7280 (N_7280,N_7009,N_7199);
and U7281 (N_7281,N_7214,N_7016);
xor U7282 (N_7282,N_7187,N_7064);
nor U7283 (N_7283,N_7182,N_7137);
nor U7284 (N_7284,N_7018,N_7093);
nand U7285 (N_7285,N_7073,N_7063);
xor U7286 (N_7286,N_7060,N_7055);
xor U7287 (N_7287,N_7048,N_7242);
or U7288 (N_7288,N_7201,N_7136);
nand U7289 (N_7289,N_7139,N_7076);
or U7290 (N_7290,N_7052,N_7118);
xor U7291 (N_7291,N_7233,N_7142);
nand U7292 (N_7292,N_7245,N_7103);
nand U7293 (N_7293,N_7202,N_7005);
nand U7294 (N_7294,N_7026,N_7038);
nand U7295 (N_7295,N_7166,N_7106);
and U7296 (N_7296,N_7225,N_7240);
nor U7297 (N_7297,N_7091,N_7015);
nand U7298 (N_7298,N_7205,N_7110);
xor U7299 (N_7299,N_7121,N_7044);
or U7300 (N_7300,N_7155,N_7065);
xnor U7301 (N_7301,N_7012,N_7180);
and U7302 (N_7302,N_7095,N_7138);
nor U7303 (N_7303,N_7014,N_7006);
or U7304 (N_7304,N_7023,N_7173);
nor U7305 (N_7305,N_7034,N_7100);
nand U7306 (N_7306,N_7248,N_7070);
xnor U7307 (N_7307,N_7194,N_7010);
xor U7308 (N_7308,N_7145,N_7088);
or U7309 (N_7309,N_7161,N_7042);
xor U7310 (N_7310,N_7033,N_7090);
nor U7311 (N_7311,N_7209,N_7045);
xor U7312 (N_7312,N_7098,N_7215);
nor U7313 (N_7313,N_7031,N_7097);
nor U7314 (N_7314,N_7071,N_7077);
or U7315 (N_7315,N_7211,N_7244);
and U7316 (N_7316,N_7167,N_7231);
nor U7317 (N_7317,N_7247,N_7210);
nor U7318 (N_7318,N_7107,N_7049);
and U7319 (N_7319,N_7133,N_7003);
nand U7320 (N_7320,N_7174,N_7229);
and U7321 (N_7321,N_7002,N_7197);
and U7322 (N_7322,N_7163,N_7219);
nand U7323 (N_7323,N_7085,N_7177);
and U7324 (N_7324,N_7036,N_7113);
nor U7325 (N_7325,N_7216,N_7223);
or U7326 (N_7326,N_7075,N_7029);
and U7327 (N_7327,N_7195,N_7017);
or U7328 (N_7328,N_7078,N_7168);
or U7329 (N_7329,N_7207,N_7109);
nand U7330 (N_7330,N_7179,N_7067);
nor U7331 (N_7331,N_7134,N_7227);
nor U7332 (N_7332,N_7112,N_7082);
or U7333 (N_7333,N_7146,N_7144);
nor U7334 (N_7334,N_7011,N_7084);
nand U7335 (N_7335,N_7081,N_7226);
xor U7336 (N_7336,N_7165,N_7032);
xor U7337 (N_7337,N_7190,N_7028);
nor U7338 (N_7338,N_7143,N_7148);
xor U7339 (N_7339,N_7234,N_7213);
or U7340 (N_7340,N_7237,N_7150);
nor U7341 (N_7341,N_7200,N_7062);
nor U7342 (N_7342,N_7151,N_7191);
xnor U7343 (N_7343,N_7123,N_7169);
and U7344 (N_7344,N_7149,N_7104);
nor U7345 (N_7345,N_7184,N_7158);
nor U7346 (N_7346,N_7124,N_7181);
xnor U7347 (N_7347,N_7102,N_7160);
or U7348 (N_7348,N_7157,N_7188);
or U7349 (N_7349,N_7129,N_7140);
or U7350 (N_7350,N_7083,N_7249);
xnor U7351 (N_7351,N_7220,N_7198);
nand U7352 (N_7352,N_7171,N_7172);
xnor U7353 (N_7353,N_7159,N_7185);
nor U7354 (N_7354,N_7001,N_7125);
xnor U7355 (N_7355,N_7008,N_7126);
and U7356 (N_7356,N_7094,N_7047);
and U7357 (N_7357,N_7053,N_7116);
xor U7358 (N_7358,N_7040,N_7218);
or U7359 (N_7359,N_7176,N_7057);
or U7360 (N_7360,N_7217,N_7072);
xnor U7361 (N_7361,N_7030,N_7224);
nor U7362 (N_7362,N_7114,N_7141);
or U7363 (N_7363,N_7130,N_7228);
or U7364 (N_7364,N_7007,N_7120);
and U7365 (N_7365,N_7027,N_7243);
nor U7366 (N_7366,N_7115,N_7203);
xor U7367 (N_7367,N_7020,N_7162);
and U7368 (N_7368,N_7152,N_7087);
xor U7369 (N_7369,N_7183,N_7192);
and U7370 (N_7370,N_7054,N_7051);
xnor U7371 (N_7371,N_7079,N_7131);
or U7372 (N_7372,N_7239,N_7135);
nor U7373 (N_7373,N_7119,N_7236);
nand U7374 (N_7374,N_7096,N_7128);
nor U7375 (N_7375,N_7153,N_7213);
and U7376 (N_7376,N_7156,N_7008);
or U7377 (N_7377,N_7167,N_7142);
nand U7378 (N_7378,N_7050,N_7013);
and U7379 (N_7379,N_7110,N_7242);
and U7380 (N_7380,N_7140,N_7103);
xnor U7381 (N_7381,N_7136,N_7057);
xnor U7382 (N_7382,N_7157,N_7164);
nand U7383 (N_7383,N_7229,N_7211);
nand U7384 (N_7384,N_7096,N_7009);
nor U7385 (N_7385,N_7137,N_7135);
and U7386 (N_7386,N_7045,N_7212);
xor U7387 (N_7387,N_7059,N_7124);
and U7388 (N_7388,N_7126,N_7022);
xnor U7389 (N_7389,N_7077,N_7115);
xor U7390 (N_7390,N_7043,N_7202);
and U7391 (N_7391,N_7104,N_7192);
or U7392 (N_7392,N_7235,N_7031);
nand U7393 (N_7393,N_7055,N_7214);
nand U7394 (N_7394,N_7067,N_7166);
xor U7395 (N_7395,N_7154,N_7008);
nand U7396 (N_7396,N_7111,N_7234);
nand U7397 (N_7397,N_7048,N_7135);
or U7398 (N_7398,N_7074,N_7130);
nor U7399 (N_7399,N_7059,N_7003);
nand U7400 (N_7400,N_7058,N_7200);
and U7401 (N_7401,N_7013,N_7146);
and U7402 (N_7402,N_7073,N_7177);
or U7403 (N_7403,N_7227,N_7199);
and U7404 (N_7404,N_7094,N_7171);
nand U7405 (N_7405,N_7032,N_7005);
nand U7406 (N_7406,N_7101,N_7167);
nand U7407 (N_7407,N_7175,N_7033);
or U7408 (N_7408,N_7046,N_7041);
and U7409 (N_7409,N_7011,N_7101);
and U7410 (N_7410,N_7142,N_7036);
xnor U7411 (N_7411,N_7047,N_7156);
nand U7412 (N_7412,N_7038,N_7120);
or U7413 (N_7413,N_7205,N_7217);
and U7414 (N_7414,N_7245,N_7147);
or U7415 (N_7415,N_7069,N_7016);
xor U7416 (N_7416,N_7226,N_7165);
and U7417 (N_7417,N_7156,N_7053);
or U7418 (N_7418,N_7079,N_7202);
or U7419 (N_7419,N_7098,N_7139);
xnor U7420 (N_7420,N_7204,N_7003);
nor U7421 (N_7421,N_7232,N_7094);
xnor U7422 (N_7422,N_7240,N_7106);
nand U7423 (N_7423,N_7226,N_7118);
or U7424 (N_7424,N_7181,N_7000);
or U7425 (N_7425,N_7004,N_7106);
and U7426 (N_7426,N_7025,N_7207);
xnor U7427 (N_7427,N_7163,N_7077);
xor U7428 (N_7428,N_7207,N_7064);
and U7429 (N_7429,N_7144,N_7224);
and U7430 (N_7430,N_7157,N_7135);
and U7431 (N_7431,N_7124,N_7171);
nor U7432 (N_7432,N_7026,N_7053);
nand U7433 (N_7433,N_7142,N_7039);
and U7434 (N_7434,N_7033,N_7180);
nand U7435 (N_7435,N_7226,N_7100);
or U7436 (N_7436,N_7131,N_7230);
or U7437 (N_7437,N_7244,N_7161);
or U7438 (N_7438,N_7075,N_7238);
and U7439 (N_7439,N_7186,N_7096);
nand U7440 (N_7440,N_7037,N_7049);
or U7441 (N_7441,N_7051,N_7186);
xnor U7442 (N_7442,N_7136,N_7054);
and U7443 (N_7443,N_7108,N_7145);
xnor U7444 (N_7444,N_7202,N_7222);
nor U7445 (N_7445,N_7183,N_7232);
nor U7446 (N_7446,N_7044,N_7054);
xnor U7447 (N_7447,N_7126,N_7207);
nor U7448 (N_7448,N_7106,N_7080);
or U7449 (N_7449,N_7094,N_7074);
xor U7450 (N_7450,N_7102,N_7186);
nor U7451 (N_7451,N_7168,N_7019);
xor U7452 (N_7452,N_7125,N_7166);
and U7453 (N_7453,N_7130,N_7045);
xnor U7454 (N_7454,N_7046,N_7146);
xor U7455 (N_7455,N_7231,N_7068);
or U7456 (N_7456,N_7057,N_7091);
or U7457 (N_7457,N_7047,N_7035);
and U7458 (N_7458,N_7085,N_7019);
nand U7459 (N_7459,N_7024,N_7030);
nand U7460 (N_7460,N_7049,N_7157);
nor U7461 (N_7461,N_7143,N_7048);
xor U7462 (N_7462,N_7068,N_7180);
nand U7463 (N_7463,N_7148,N_7238);
nor U7464 (N_7464,N_7179,N_7107);
xnor U7465 (N_7465,N_7105,N_7133);
nand U7466 (N_7466,N_7180,N_7048);
or U7467 (N_7467,N_7175,N_7180);
or U7468 (N_7468,N_7034,N_7214);
xor U7469 (N_7469,N_7137,N_7184);
nand U7470 (N_7470,N_7243,N_7164);
nand U7471 (N_7471,N_7012,N_7070);
and U7472 (N_7472,N_7089,N_7179);
nor U7473 (N_7473,N_7177,N_7209);
nand U7474 (N_7474,N_7008,N_7241);
nor U7475 (N_7475,N_7131,N_7111);
nor U7476 (N_7476,N_7006,N_7106);
and U7477 (N_7477,N_7053,N_7091);
nor U7478 (N_7478,N_7196,N_7024);
nor U7479 (N_7479,N_7198,N_7128);
xnor U7480 (N_7480,N_7229,N_7068);
nand U7481 (N_7481,N_7121,N_7081);
nand U7482 (N_7482,N_7182,N_7070);
nand U7483 (N_7483,N_7186,N_7191);
xor U7484 (N_7484,N_7156,N_7169);
nand U7485 (N_7485,N_7038,N_7245);
xnor U7486 (N_7486,N_7211,N_7101);
nand U7487 (N_7487,N_7114,N_7128);
nand U7488 (N_7488,N_7134,N_7084);
or U7489 (N_7489,N_7198,N_7009);
or U7490 (N_7490,N_7011,N_7050);
xor U7491 (N_7491,N_7218,N_7198);
nand U7492 (N_7492,N_7239,N_7030);
or U7493 (N_7493,N_7182,N_7246);
or U7494 (N_7494,N_7110,N_7005);
nor U7495 (N_7495,N_7164,N_7083);
nor U7496 (N_7496,N_7215,N_7176);
xnor U7497 (N_7497,N_7002,N_7113);
and U7498 (N_7498,N_7173,N_7218);
and U7499 (N_7499,N_7244,N_7072);
nand U7500 (N_7500,N_7368,N_7471);
or U7501 (N_7501,N_7295,N_7409);
nand U7502 (N_7502,N_7397,N_7421);
xor U7503 (N_7503,N_7481,N_7458);
and U7504 (N_7504,N_7418,N_7302);
nor U7505 (N_7505,N_7306,N_7489);
nand U7506 (N_7506,N_7322,N_7326);
nand U7507 (N_7507,N_7460,N_7382);
and U7508 (N_7508,N_7420,N_7463);
nor U7509 (N_7509,N_7320,N_7424);
and U7510 (N_7510,N_7318,N_7362);
or U7511 (N_7511,N_7398,N_7276);
nand U7512 (N_7512,N_7499,N_7453);
xor U7513 (N_7513,N_7293,N_7317);
nor U7514 (N_7514,N_7422,N_7256);
or U7515 (N_7515,N_7344,N_7478);
xor U7516 (N_7516,N_7270,N_7430);
xnor U7517 (N_7517,N_7319,N_7253);
and U7518 (N_7518,N_7485,N_7442);
xor U7519 (N_7519,N_7493,N_7267);
and U7520 (N_7520,N_7413,N_7494);
nor U7521 (N_7521,N_7416,N_7364);
and U7522 (N_7522,N_7254,N_7262);
or U7523 (N_7523,N_7432,N_7454);
nor U7524 (N_7524,N_7446,N_7333);
nor U7525 (N_7525,N_7325,N_7323);
or U7526 (N_7526,N_7483,N_7434);
nor U7527 (N_7527,N_7370,N_7404);
nand U7528 (N_7528,N_7451,N_7327);
or U7529 (N_7529,N_7435,N_7415);
xor U7530 (N_7530,N_7329,N_7498);
nor U7531 (N_7531,N_7427,N_7476);
nand U7532 (N_7532,N_7261,N_7285);
and U7533 (N_7533,N_7353,N_7495);
xor U7534 (N_7534,N_7300,N_7426);
nand U7535 (N_7535,N_7341,N_7337);
and U7536 (N_7536,N_7484,N_7252);
nand U7537 (N_7537,N_7265,N_7290);
or U7538 (N_7538,N_7266,N_7393);
or U7539 (N_7539,N_7258,N_7359);
nand U7540 (N_7540,N_7299,N_7473);
or U7541 (N_7541,N_7307,N_7440);
nor U7542 (N_7542,N_7257,N_7355);
nor U7543 (N_7543,N_7277,N_7291);
and U7544 (N_7544,N_7284,N_7330);
or U7545 (N_7545,N_7444,N_7412);
nor U7546 (N_7546,N_7264,N_7487);
or U7547 (N_7547,N_7286,N_7358);
or U7548 (N_7548,N_7271,N_7443);
or U7549 (N_7549,N_7400,N_7305);
xnor U7550 (N_7550,N_7372,N_7376);
and U7551 (N_7551,N_7332,N_7461);
and U7552 (N_7552,N_7439,N_7402);
and U7553 (N_7553,N_7437,N_7380);
nand U7554 (N_7554,N_7312,N_7349);
xor U7555 (N_7555,N_7331,N_7445);
nand U7556 (N_7556,N_7496,N_7470);
xnor U7557 (N_7557,N_7298,N_7260);
nand U7558 (N_7558,N_7351,N_7314);
xnor U7559 (N_7559,N_7449,N_7360);
nand U7560 (N_7560,N_7391,N_7414);
and U7561 (N_7561,N_7396,N_7255);
nor U7562 (N_7562,N_7309,N_7321);
and U7563 (N_7563,N_7450,N_7399);
nor U7564 (N_7564,N_7294,N_7480);
nor U7565 (N_7565,N_7292,N_7388);
or U7566 (N_7566,N_7462,N_7394);
nor U7567 (N_7567,N_7456,N_7328);
nand U7568 (N_7568,N_7386,N_7342);
nor U7569 (N_7569,N_7410,N_7259);
nand U7570 (N_7570,N_7310,N_7269);
xnor U7571 (N_7571,N_7308,N_7459);
xnor U7572 (N_7572,N_7275,N_7346);
or U7573 (N_7573,N_7369,N_7385);
or U7574 (N_7574,N_7490,N_7296);
nand U7575 (N_7575,N_7303,N_7497);
or U7576 (N_7576,N_7316,N_7288);
nand U7577 (N_7577,N_7441,N_7345);
and U7578 (N_7578,N_7488,N_7313);
xnor U7579 (N_7579,N_7374,N_7447);
and U7580 (N_7580,N_7395,N_7468);
and U7581 (N_7581,N_7407,N_7373);
nor U7582 (N_7582,N_7315,N_7352);
or U7583 (N_7583,N_7336,N_7401);
xnor U7584 (N_7584,N_7465,N_7281);
nor U7585 (N_7585,N_7477,N_7278);
nand U7586 (N_7586,N_7438,N_7452);
nand U7587 (N_7587,N_7340,N_7455);
nand U7588 (N_7588,N_7387,N_7492);
xor U7589 (N_7589,N_7289,N_7486);
nand U7590 (N_7590,N_7475,N_7287);
or U7591 (N_7591,N_7464,N_7384);
and U7592 (N_7592,N_7301,N_7390);
xnor U7593 (N_7593,N_7457,N_7363);
nor U7594 (N_7594,N_7466,N_7403);
nand U7595 (N_7595,N_7392,N_7425);
nand U7596 (N_7596,N_7389,N_7405);
and U7597 (N_7597,N_7448,N_7304);
or U7598 (N_7598,N_7263,N_7311);
or U7599 (N_7599,N_7274,N_7338);
or U7600 (N_7600,N_7371,N_7423);
nand U7601 (N_7601,N_7431,N_7354);
and U7602 (N_7602,N_7279,N_7429);
and U7603 (N_7603,N_7361,N_7377);
xnor U7604 (N_7604,N_7335,N_7365);
and U7605 (N_7605,N_7268,N_7357);
nand U7606 (N_7606,N_7283,N_7280);
nor U7607 (N_7607,N_7273,N_7297);
or U7608 (N_7608,N_7428,N_7350);
nor U7609 (N_7609,N_7367,N_7324);
or U7610 (N_7610,N_7343,N_7282);
xnor U7611 (N_7611,N_7436,N_7491);
nor U7612 (N_7612,N_7479,N_7381);
nor U7613 (N_7613,N_7366,N_7482);
nand U7614 (N_7614,N_7411,N_7339);
and U7615 (N_7615,N_7467,N_7379);
xor U7616 (N_7616,N_7347,N_7469);
and U7617 (N_7617,N_7272,N_7433);
nand U7618 (N_7618,N_7408,N_7417);
and U7619 (N_7619,N_7334,N_7378);
nor U7620 (N_7620,N_7472,N_7356);
nand U7621 (N_7621,N_7375,N_7419);
nand U7622 (N_7622,N_7474,N_7406);
or U7623 (N_7623,N_7348,N_7251);
nand U7624 (N_7624,N_7383,N_7250);
nor U7625 (N_7625,N_7274,N_7435);
nand U7626 (N_7626,N_7390,N_7304);
and U7627 (N_7627,N_7358,N_7393);
nand U7628 (N_7628,N_7319,N_7411);
xor U7629 (N_7629,N_7364,N_7262);
and U7630 (N_7630,N_7322,N_7407);
nor U7631 (N_7631,N_7394,N_7431);
xnor U7632 (N_7632,N_7367,N_7375);
nand U7633 (N_7633,N_7478,N_7460);
nor U7634 (N_7634,N_7252,N_7300);
and U7635 (N_7635,N_7477,N_7329);
nand U7636 (N_7636,N_7353,N_7435);
and U7637 (N_7637,N_7375,N_7405);
nor U7638 (N_7638,N_7432,N_7331);
xnor U7639 (N_7639,N_7257,N_7322);
nand U7640 (N_7640,N_7335,N_7466);
nor U7641 (N_7641,N_7359,N_7321);
nand U7642 (N_7642,N_7400,N_7299);
xor U7643 (N_7643,N_7309,N_7437);
and U7644 (N_7644,N_7453,N_7383);
xor U7645 (N_7645,N_7428,N_7330);
or U7646 (N_7646,N_7385,N_7485);
xor U7647 (N_7647,N_7269,N_7458);
xor U7648 (N_7648,N_7263,N_7278);
and U7649 (N_7649,N_7343,N_7397);
or U7650 (N_7650,N_7453,N_7312);
nand U7651 (N_7651,N_7498,N_7377);
nand U7652 (N_7652,N_7352,N_7307);
xor U7653 (N_7653,N_7283,N_7435);
and U7654 (N_7654,N_7278,N_7422);
nand U7655 (N_7655,N_7395,N_7472);
xor U7656 (N_7656,N_7444,N_7375);
nor U7657 (N_7657,N_7354,N_7264);
nor U7658 (N_7658,N_7361,N_7499);
nor U7659 (N_7659,N_7316,N_7278);
xor U7660 (N_7660,N_7301,N_7380);
xnor U7661 (N_7661,N_7391,N_7445);
nor U7662 (N_7662,N_7432,N_7327);
nor U7663 (N_7663,N_7482,N_7392);
nor U7664 (N_7664,N_7432,N_7319);
or U7665 (N_7665,N_7393,N_7276);
nor U7666 (N_7666,N_7453,N_7491);
or U7667 (N_7667,N_7416,N_7288);
or U7668 (N_7668,N_7484,N_7286);
or U7669 (N_7669,N_7412,N_7359);
nand U7670 (N_7670,N_7303,N_7494);
xnor U7671 (N_7671,N_7446,N_7383);
nand U7672 (N_7672,N_7477,N_7387);
and U7673 (N_7673,N_7433,N_7457);
nand U7674 (N_7674,N_7268,N_7468);
nand U7675 (N_7675,N_7321,N_7443);
nor U7676 (N_7676,N_7445,N_7413);
or U7677 (N_7677,N_7273,N_7290);
nand U7678 (N_7678,N_7366,N_7383);
xnor U7679 (N_7679,N_7416,N_7266);
xor U7680 (N_7680,N_7368,N_7485);
nor U7681 (N_7681,N_7343,N_7408);
nand U7682 (N_7682,N_7304,N_7435);
and U7683 (N_7683,N_7425,N_7365);
nand U7684 (N_7684,N_7277,N_7292);
xor U7685 (N_7685,N_7460,N_7367);
nor U7686 (N_7686,N_7361,N_7258);
xor U7687 (N_7687,N_7453,N_7403);
xor U7688 (N_7688,N_7271,N_7450);
or U7689 (N_7689,N_7359,N_7405);
xnor U7690 (N_7690,N_7464,N_7491);
or U7691 (N_7691,N_7474,N_7431);
and U7692 (N_7692,N_7346,N_7441);
nand U7693 (N_7693,N_7250,N_7274);
nor U7694 (N_7694,N_7455,N_7459);
xnor U7695 (N_7695,N_7321,N_7363);
xor U7696 (N_7696,N_7254,N_7329);
xnor U7697 (N_7697,N_7441,N_7272);
xnor U7698 (N_7698,N_7396,N_7375);
xnor U7699 (N_7699,N_7291,N_7428);
nand U7700 (N_7700,N_7393,N_7259);
and U7701 (N_7701,N_7292,N_7483);
or U7702 (N_7702,N_7327,N_7470);
xnor U7703 (N_7703,N_7340,N_7433);
xor U7704 (N_7704,N_7285,N_7478);
xor U7705 (N_7705,N_7343,N_7429);
nor U7706 (N_7706,N_7323,N_7483);
xnor U7707 (N_7707,N_7356,N_7259);
nor U7708 (N_7708,N_7271,N_7351);
xnor U7709 (N_7709,N_7334,N_7252);
or U7710 (N_7710,N_7265,N_7421);
and U7711 (N_7711,N_7340,N_7374);
nor U7712 (N_7712,N_7342,N_7473);
nand U7713 (N_7713,N_7397,N_7326);
nand U7714 (N_7714,N_7446,N_7269);
or U7715 (N_7715,N_7484,N_7325);
nand U7716 (N_7716,N_7290,N_7261);
nand U7717 (N_7717,N_7386,N_7286);
or U7718 (N_7718,N_7289,N_7389);
and U7719 (N_7719,N_7427,N_7294);
nand U7720 (N_7720,N_7383,N_7373);
nand U7721 (N_7721,N_7428,N_7298);
nand U7722 (N_7722,N_7452,N_7419);
and U7723 (N_7723,N_7499,N_7424);
or U7724 (N_7724,N_7292,N_7452);
nand U7725 (N_7725,N_7492,N_7364);
xnor U7726 (N_7726,N_7260,N_7489);
nand U7727 (N_7727,N_7498,N_7292);
nand U7728 (N_7728,N_7317,N_7321);
nor U7729 (N_7729,N_7343,N_7437);
nand U7730 (N_7730,N_7423,N_7472);
and U7731 (N_7731,N_7254,N_7318);
xor U7732 (N_7732,N_7349,N_7379);
nor U7733 (N_7733,N_7479,N_7462);
and U7734 (N_7734,N_7412,N_7498);
xor U7735 (N_7735,N_7370,N_7360);
nand U7736 (N_7736,N_7439,N_7395);
or U7737 (N_7737,N_7403,N_7431);
and U7738 (N_7738,N_7480,N_7271);
nand U7739 (N_7739,N_7282,N_7355);
or U7740 (N_7740,N_7393,N_7449);
nand U7741 (N_7741,N_7275,N_7342);
xnor U7742 (N_7742,N_7325,N_7467);
and U7743 (N_7743,N_7431,N_7375);
and U7744 (N_7744,N_7303,N_7388);
or U7745 (N_7745,N_7414,N_7389);
nand U7746 (N_7746,N_7328,N_7444);
nand U7747 (N_7747,N_7307,N_7387);
xnor U7748 (N_7748,N_7343,N_7430);
and U7749 (N_7749,N_7373,N_7368);
nor U7750 (N_7750,N_7749,N_7652);
and U7751 (N_7751,N_7735,N_7502);
nand U7752 (N_7752,N_7513,N_7514);
nand U7753 (N_7753,N_7686,N_7679);
or U7754 (N_7754,N_7542,N_7661);
nand U7755 (N_7755,N_7741,N_7729);
nand U7756 (N_7756,N_7706,N_7575);
xor U7757 (N_7757,N_7731,N_7659);
and U7758 (N_7758,N_7628,N_7733);
and U7759 (N_7759,N_7690,N_7693);
xor U7760 (N_7760,N_7521,N_7527);
or U7761 (N_7761,N_7534,N_7543);
xnor U7762 (N_7762,N_7503,N_7717);
xnor U7763 (N_7763,N_7562,N_7650);
nand U7764 (N_7764,N_7639,N_7589);
nand U7765 (N_7765,N_7538,N_7605);
or U7766 (N_7766,N_7746,N_7703);
nor U7767 (N_7767,N_7501,N_7546);
or U7768 (N_7768,N_7643,N_7663);
xor U7769 (N_7769,N_7636,N_7713);
nor U7770 (N_7770,N_7736,N_7582);
and U7771 (N_7771,N_7657,N_7545);
and U7772 (N_7772,N_7518,N_7596);
nor U7773 (N_7773,N_7645,N_7539);
or U7774 (N_7774,N_7553,N_7547);
nor U7775 (N_7775,N_7620,N_7675);
nand U7776 (N_7776,N_7555,N_7550);
xor U7777 (N_7777,N_7603,N_7525);
and U7778 (N_7778,N_7611,N_7588);
and U7779 (N_7779,N_7610,N_7597);
or U7780 (N_7780,N_7642,N_7532);
xnor U7781 (N_7781,N_7601,N_7725);
and U7782 (N_7782,N_7508,N_7609);
nor U7783 (N_7783,N_7646,N_7738);
or U7784 (N_7784,N_7530,N_7608);
nor U7785 (N_7785,N_7578,N_7549);
xnor U7786 (N_7786,N_7590,N_7627);
xnor U7787 (N_7787,N_7685,N_7535);
nand U7788 (N_7788,N_7612,N_7580);
or U7789 (N_7789,N_7629,N_7734);
nand U7790 (N_7790,N_7699,N_7574);
or U7791 (N_7791,N_7509,N_7592);
or U7792 (N_7792,N_7737,N_7747);
xor U7793 (N_7793,N_7533,N_7520);
xor U7794 (N_7794,N_7709,N_7585);
nand U7795 (N_7795,N_7651,N_7587);
xor U7796 (N_7796,N_7656,N_7724);
nand U7797 (N_7797,N_7682,N_7640);
nor U7798 (N_7798,N_7564,N_7678);
or U7799 (N_7799,N_7625,N_7722);
xor U7800 (N_7800,N_7654,N_7743);
xnor U7801 (N_7801,N_7568,N_7701);
xor U7802 (N_7802,N_7666,N_7674);
nor U7803 (N_7803,N_7698,N_7524);
nor U7804 (N_7804,N_7565,N_7669);
and U7805 (N_7805,N_7576,N_7660);
nor U7806 (N_7806,N_7710,N_7551);
nor U7807 (N_7807,N_7536,N_7544);
and U7808 (N_7808,N_7632,N_7711);
and U7809 (N_7809,N_7558,N_7563);
nor U7810 (N_7810,N_7680,N_7500);
nand U7811 (N_7811,N_7619,N_7623);
nor U7812 (N_7812,N_7617,N_7740);
and U7813 (N_7813,N_7606,N_7649);
nand U7814 (N_7814,N_7707,N_7664);
nor U7815 (N_7815,N_7705,N_7655);
xor U7816 (N_7816,N_7677,N_7630);
and U7817 (N_7817,N_7591,N_7571);
nand U7818 (N_7818,N_7505,N_7604);
or U7819 (N_7819,N_7579,N_7519);
or U7820 (N_7820,N_7621,N_7613);
xnor U7821 (N_7821,N_7607,N_7692);
xor U7822 (N_7822,N_7511,N_7648);
nand U7823 (N_7823,N_7522,N_7572);
or U7824 (N_7824,N_7715,N_7531);
xnor U7825 (N_7825,N_7665,N_7566);
nor U7826 (N_7826,N_7593,N_7644);
and U7827 (N_7827,N_7714,N_7581);
nor U7828 (N_7828,N_7559,N_7723);
nand U7829 (N_7829,N_7742,N_7673);
xnor U7830 (N_7830,N_7569,N_7622);
nand U7831 (N_7831,N_7744,N_7681);
or U7832 (N_7832,N_7689,N_7694);
xnor U7833 (N_7833,N_7634,N_7626);
and U7834 (N_7834,N_7616,N_7584);
nand U7835 (N_7835,N_7517,N_7577);
or U7836 (N_7836,N_7583,N_7662);
nor U7837 (N_7837,N_7702,N_7510);
or U7838 (N_7838,N_7688,N_7515);
and U7839 (N_7839,N_7599,N_7700);
nand U7840 (N_7840,N_7719,N_7618);
xor U7841 (N_7841,N_7529,N_7516);
xor U7842 (N_7842,N_7560,N_7614);
and U7843 (N_7843,N_7586,N_7602);
nand U7844 (N_7844,N_7507,N_7670);
nand U7845 (N_7845,N_7720,N_7540);
nor U7846 (N_7846,N_7667,N_7615);
nor U7847 (N_7847,N_7541,N_7552);
nor U7848 (N_7848,N_7697,N_7647);
nand U7849 (N_7849,N_7668,N_7671);
and U7850 (N_7850,N_7537,N_7637);
nand U7851 (N_7851,N_7745,N_7716);
or U7852 (N_7852,N_7696,N_7570);
nand U7853 (N_7853,N_7676,N_7635);
and U7854 (N_7854,N_7573,N_7730);
or U7855 (N_7855,N_7561,N_7684);
nor U7856 (N_7856,N_7732,N_7641);
and U7857 (N_7857,N_7557,N_7658);
xor U7858 (N_7858,N_7726,N_7523);
nand U7859 (N_7859,N_7653,N_7512);
or U7860 (N_7860,N_7506,N_7718);
nor U7861 (N_7861,N_7739,N_7554);
nand U7862 (N_7862,N_7595,N_7598);
or U7863 (N_7863,N_7526,N_7748);
or U7864 (N_7864,N_7633,N_7691);
xnor U7865 (N_7865,N_7638,N_7594);
and U7866 (N_7866,N_7721,N_7528);
or U7867 (N_7867,N_7600,N_7631);
or U7868 (N_7868,N_7708,N_7683);
and U7869 (N_7869,N_7672,N_7712);
and U7870 (N_7870,N_7548,N_7687);
or U7871 (N_7871,N_7504,N_7695);
and U7872 (N_7872,N_7727,N_7728);
nor U7873 (N_7873,N_7624,N_7556);
and U7874 (N_7874,N_7704,N_7567);
xnor U7875 (N_7875,N_7562,N_7666);
xor U7876 (N_7876,N_7604,N_7719);
and U7877 (N_7877,N_7566,N_7547);
xor U7878 (N_7878,N_7578,N_7532);
and U7879 (N_7879,N_7637,N_7730);
and U7880 (N_7880,N_7614,N_7577);
xnor U7881 (N_7881,N_7613,N_7567);
nand U7882 (N_7882,N_7544,N_7609);
and U7883 (N_7883,N_7640,N_7656);
nor U7884 (N_7884,N_7536,N_7568);
or U7885 (N_7885,N_7728,N_7676);
nand U7886 (N_7886,N_7717,N_7573);
xnor U7887 (N_7887,N_7680,N_7631);
nand U7888 (N_7888,N_7682,N_7576);
and U7889 (N_7889,N_7733,N_7649);
and U7890 (N_7890,N_7639,N_7689);
nor U7891 (N_7891,N_7678,N_7714);
and U7892 (N_7892,N_7527,N_7629);
or U7893 (N_7893,N_7563,N_7628);
and U7894 (N_7894,N_7575,N_7744);
nor U7895 (N_7895,N_7659,N_7644);
xnor U7896 (N_7896,N_7595,N_7532);
and U7897 (N_7897,N_7631,N_7581);
xor U7898 (N_7898,N_7735,N_7582);
nor U7899 (N_7899,N_7540,N_7681);
nor U7900 (N_7900,N_7635,N_7572);
nand U7901 (N_7901,N_7617,N_7599);
nor U7902 (N_7902,N_7599,N_7639);
nor U7903 (N_7903,N_7739,N_7548);
nor U7904 (N_7904,N_7648,N_7739);
or U7905 (N_7905,N_7705,N_7507);
nor U7906 (N_7906,N_7576,N_7681);
or U7907 (N_7907,N_7523,N_7568);
and U7908 (N_7908,N_7550,N_7564);
nor U7909 (N_7909,N_7663,N_7725);
xor U7910 (N_7910,N_7621,N_7683);
nor U7911 (N_7911,N_7667,N_7507);
xor U7912 (N_7912,N_7670,N_7506);
and U7913 (N_7913,N_7544,N_7747);
and U7914 (N_7914,N_7629,N_7737);
xnor U7915 (N_7915,N_7725,N_7742);
nor U7916 (N_7916,N_7620,N_7562);
nand U7917 (N_7917,N_7672,N_7637);
and U7918 (N_7918,N_7701,N_7738);
xnor U7919 (N_7919,N_7660,N_7573);
and U7920 (N_7920,N_7732,N_7538);
nor U7921 (N_7921,N_7552,N_7588);
or U7922 (N_7922,N_7653,N_7623);
xor U7923 (N_7923,N_7739,N_7655);
xnor U7924 (N_7924,N_7711,N_7735);
or U7925 (N_7925,N_7674,N_7745);
xnor U7926 (N_7926,N_7730,N_7646);
xnor U7927 (N_7927,N_7562,N_7524);
xnor U7928 (N_7928,N_7663,N_7526);
xor U7929 (N_7929,N_7590,N_7518);
and U7930 (N_7930,N_7663,N_7684);
and U7931 (N_7931,N_7530,N_7640);
or U7932 (N_7932,N_7707,N_7674);
or U7933 (N_7933,N_7541,N_7725);
and U7934 (N_7934,N_7565,N_7749);
nor U7935 (N_7935,N_7635,N_7665);
and U7936 (N_7936,N_7611,N_7747);
nand U7937 (N_7937,N_7623,N_7534);
nor U7938 (N_7938,N_7606,N_7590);
nor U7939 (N_7939,N_7507,N_7641);
and U7940 (N_7940,N_7617,N_7510);
and U7941 (N_7941,N_7504,N_7734);
xor U7942 (N_7942,N_7569,N_7725);
nor U7943 (N_7943,N_7551,N_7696);
xnor U7944 (N_7944,N_7723,N_7592);
xor U7945 (N_7945,N_7560,N_7642);
nor U7946 (N_7946,N_7536,N_7714);
xor U7947 (N_7947,N_7500,N_7588);
xor U7948 (N_7948,N_7520,N_7644);
or U7949 (N_7949,N_7724,N_7741);
and U7950 (N_7950,N_7746,N_7735);
and U7951 (N_7951,N_7623,N_7564);
or U7952 (N_7952,N_7603,N_7618);
xnor U7953 (N_7953,N_7545,N_7541);
or U7954 (N_7954,N_7541,N_7727);
xnor U7955 (N_7955,N_7740,N_7706);
nor U7956 (N_7956,N_7576,N_7549);
or U7957 (N_7957,N_7742,N_7534);
nor U7958 (N_7958,N_7642,N_7656);
nand U7959 (N_7959,N_7561,N_7708);
xnor U7960 (N_7960,N_7701,N_7528);
or U7961 (N_7961,N_7724,N_7539);
nor U7962 (N_7962,N_7559,N_7636);
xnor U7963 (N_7963,N_7697,N_7615);
and U7964 (N_7964,N_7747,N_7671);
nand U7965 (N_7965,N_7697,N_7620);
nand U7966 (N_7966,N_7528,N_7556);
and U7967 (N_7967,N_7635,N_7685);
nand U7968 (N_7968,N_7540,N_7532);
nand U7969 (N_7969,N_7564,N_7533);
nand U7970 (N_7970,N_7724,N_7516);
xor U7971 (N_7971,N_7620,N_7636);
and U7972 (N_7972,N_7531,N_7614);
nand U7973 (N_7973,N_7538,N_7588);
xor U7974 (N_7974,N_7589,N_7718);
nand U7975 (N_7975,N_7652,N_7677);
or U7976 (N_7976,N_7677,N_7657);
nand U7977 (N_7977,N_7666,N_7721);
nand U7978 (N_7978,N_7602,N_7711);
and U7979 (N_7979,N_7579,N_7598);
nand U7980 (N_7980,N_7609,N_7646);
nor U7981 (N_7981,N_7657,N_7739);
or U7982 (N_7982,N_7661,N_7543);
nand U7983 (N_7983,N_7658,N_7696);
xnor U7984 (N_7984,N_7591,N_7505);
xnor U7985 (N_7985,N_7688,N_7563);
or U7986 (N_7986,N_7667,N_7561);
or U7987 (N_7987,N_7704,N_7691);
nor U7988 (N_7988,N_7625,N_7686);
and U7989 (N_7989,N_7714,N_7583);
xnor U7990 (N_7990,N_7640,N_7602);
xnor U7991 (N_7991,N_7637,N_7707);
and U7992 (N_7992,N_7678,N_7654);
or U7993 (N_7993,N_7649,N_7581);
or U7994 (N_7994,N_7713,N_7702);
xor U7995 (N_7995,N_7672,N_7625);
and U7996 (N_7996,N_7587,N_7635);
nand U7997 (N_7997,N_7637,N_7518);
nor U7998 (N_7998,N_7614,N_7616);
nor U7999 (N_7999,N_7626,N_7503);
and U8000 (N_8000,N_7896,N_7899);
xor U8001 (N_8001,N_7811,N_7763);
xnor U8002 (N_8002,N_7879,N_7978);
xnor U8003 (N_8003,N_7860,N_7838);
xnor U8004 (N_8004,N_7801,N_7847);
or U8005 (N_8005,N_7928,N_7891);
xnor U8006 (N_8006,N_7881,N_7994);
nand U8007 (N_8007,N_7775,N_7766);
nor U8008 (N_8008,N_7772,N_7981);
and U8009 (N_8009,N_7950,N_7855);
and U8010 (N_8010,N_7780,N_7826);
nand U8011 (N_8011,N_7751,N_7823);
xnor U8012 (N_8012,N_7784,N_7959);
xor U8013 (N_8013,N_7869,N_7874);
xnor U8014 (N_8014,N_7791,N_7863);
nor U8015 (N_8015,N_7974,N_7979);
and U8016 (N_8016,N_7888,N_7931);
nor U8017 (N_8017,N_7967,N_7902);
or U8018 (N_8018,N_7901,N_7827);
and U8019 (N_8019,N_7969,N_7854);
and U8020 (N_8020,N_7929,N_7880);
or U8021 (N_8021,N_7982,N_7940);
nand U8022 (N_8022,N_7819,N_7794);
xnor U8023 (N_8023,N_7996,N_7988);
or U8024 (N_8024,N_7870,N_7760);
xnor U8025 (N_8025,N_7927,N_7814);
nand U8026 (N_8026,N_7900,N_7764);
nand U8027 (N_8027,N_7799,N_7924);
nand U8028 (N_8028,N_7807,N_7951);
or U8029 (N_8029,N_7970,N_7804);
or U8030 (N_8030,N_7808,N_7973);
nor U8031 (N_8031,N_7977,N_7935);
and U8032 (N_8032,N_7786,N_7972);
nand U8033 (N_8033,N_7858,N_7865);
nor U8034 (N_8034,N_7803,N_7939);
nand U8035 (N_8035,N_7904,N_7948);
or U8036 (N_8036,N_7806,N_7839);
xor U8037 (N_8037,N_7933,N_7975);
nand U8038 (N_8038,N_7836,N_7882);
and U8039 (N_8039,N_7923,N_7862);
and U8040 (N_8040,N_7918,N_7831);
or U8041 (N_8041,N_7800,N_7779);
or U8042 (N_8042,N_7774,N_7825);
and U8043 (N_8043,N_7944,N_7966);
and U8044 (N_8044,N_7943,N_7828);
xnor U8045 (N_8045,N_7818,N_7890);
nor U8046 (N_8046,N_7897,N_7946);
xor U8047 (N_8047,N_7752,N_7873);
or U8048 (N_8048,N_7952,N_7958);
and U8049 (N_8049,N_7983,N_7954);
and U8050 (N_8050,N_7905,N_7914);
or U8051 (N_8051,N_7930,N_7817);
or U8052 (N_8052,N_7945,N_7856);
xnor U8053 (N_8053,N_7908,N_7789);
nor U8054 (N_8054,N_7991,N_7842);
and U8055 (N_8055,N_7999,N_7909);
xnor U8056 (N_8056,N_7877,N_7989);
or U8057 (N_8057,N_7898,N_7833);
xnor U8058 (N_8058,N_7990,N_7859);
xnor U8059 (N_8059,N_7997,N_7797);
nor U8060 (N_8060,N_7802,N_7926);
or U8061 (N_8061,N_7867,N_7956);
and U8062 (N_8062,N_7987,N_7916);
nor U8063 (N_8063,N_7915,N_7850);
xnor U8064 (N_8064,N_7822,N_7750);
nor U8065 (N_8065,N_7947,N_7864);
nand U8066 (N_8066,N_7984,N_7913);
xnor U8067 (N_8067,N_7821,N_7871);
xnor U8068 (N_8068,N_7887,N_7875);
or U8069 (N_8069,N_7942,N_7770);
or U8070 (N_8070,N_7921,N_7995);
or U8071 (N_8071,N_7773,N_7851);
nand U8072 (N_8072,N_7816,N_7798);
and U8073 (N_8073,N_7829,N_7776);
and U8074 (N_8074,N_7853,N_7980);
nand U8075 (N_8075,N_7998,N_7761);
nand U8076 (N_8076,N_7815,N_7992);
and U8077 (N_8077,N_7961,N_7755);
nor U8078 (N_8078,N_7976,N_7759);
nor U8079 (N_8079,N_7957,N_7837);
and U8080 (N_8080,N_7894,N_7883);
xor U8081 (N_8081,N_7872,N_7778);
or U8082 (N_8082,N_7937,N_7846);
nor U8083 (N_8083,N_7765,N_7812);
and U8084 (N_8084,N_7895,N_7925);
nor U8085 (N_8085,N_7968,N_7841);
xor U8086 (N_8086,N_7889,N_7767);
nand U8087 (N_8087,N_7849,N_7790);
nand U8088 (N_8088,N_7886,N_7920);
or U8089 (N_8089,N_7844,N_7787);
nand U8090 (N_8090,N_7885,N_7960);
and U8091 (N_8091,N_7820,N_7932);
xor U8092 (N_8092,N_7758,N_7936);
nand U8093 (N_8093,N_7852,N_7906);
nor U8094 (N_8094,N_7771,N_7795);
xor U8095 (N_8095,N_7965,N_7805);
xor U8096 (N_8096,N_7949,N_7986);
xnor U8097 (N_8097,N_7917,N_7830);
xnor U8098 (N_8098,N_7971,N_7832);
and U8099 (N_8099,N_7907,N_7962);
xnor U8100 (N_8100,N_7753,N_7964);
nor U8101 (N_8101,N_7824,N_7985);
nor U8102 (N_8102,N_7868,N_7754);
xnor U8103 (N_8103,N_7963,N_7878);
and U8104 (N_8104,N_7861,N_7892);
nand U8105 (N_8105,N_7835,N_7876);
nand U8106 (N_8106,N_7938,N_7922);
and U8107 (N_8107,N_7783,N_7809);
or U8108 (N_8108,N_7893,N_7813);
nor U8109 (N_8109,N_7785,N_7781);
xor U8110 (N_8110,N_7792,N_7941);
and U8111 (N_8111,N_7911,N_7843);
nand U8112 (N_8112,N_7840,N_7834);
or U8113 (N_8113,N_7884,N_7912);
xnor U8114 (N_8114,N_7793,N_7768);
xnor U8115 (N_8115,N_7810,N_7782);
nor U8116 (N_8116,N_7777,N_7953);
nor U8117 (N_8117,N_7993,N_7955);
xor U8118 (N_8118,N_7769,N_7757);
nor U8119 (N_8119,N_7857,N_7903);
nand U8120 (N_8120,N_7796,N_7756);
or U8121 (N_8121,N_7788,N_7762);
xnor U8122 (N_8122,N_7848,N_7934);
nand U8123 (N_8123,N_7845,N_7910);
and U8124 (N_8124,N_7866,N_7919);
xor U8125 (N_8125,N_7807,N_7848);
nor U8126 (N_8126,N_7995,N_7868);
xnor U8127 (N_8127,N_7914,N_7781);
nand U8128 (N_8128,N_7879,N_7951);
nor U8129 (N_8129,N_7839,N_7969);
nand U8130 (N_8130,N_7865,N_7957);
nor U8131 (N_8131,N_7764,N_7854);
nor U8132 (N_8132,N_7870,N_7984);
nand U8133 (N_8133,N_7994,N_7988);
or U8134 (N_8134,N_7895,N_7778);
nand U8135 (N_8135,N_7851,N_7899);
xor U8136 (N_8136,N_7940,N_7976);
nand U8137 (N_8137,N_7794,N_7998);
or U8138 (N_8138,N_7833,N_7927);
or U8139 (N_8139,N_7826,N_7880);
xor U8140 (N_8140,N_7881,N_7924);
nor U8141 (N_8141,N_7794,N_7906);
and U8142 (N_8142,N_7763,N_7767);
and U8143 (N_8143,N_7868,N_7932);
nand U8144 (N_8144,N_7817,N_7954);
nand U8145 (N_8145,N_7968,N_7990);
or U8146 (N_8146,N_7795,N_7892);
nand U8147 (N_8147,N_7928,N_7772);
nor U8148 (N_8148,N_7892,N_7821);
and U8149 (N_8149,N_7993,N_7808);
xor U8150 (N_8150,N_7963,N_7959);
nor U8151 (N_8151,N_7936,N_7980);
and U8152 (N_8152,N_7864,N_7865);
nand U8153 (N_8153,N_7928,N_7943);
or U8154 (N_8154,N_7996,N_7919);
xnor U8155 (N_8155,N_7794,N_7974);
and U8156 (N_8156,N_7911,N_7833);
and U8157 (N_8157,N_7961,N_7796);
and U8158 (N_8158,N_7892,N_7851);
xnor U8159 (N_8159,N_7878,N_7791);
xnor U8160 (N_8160,N_7821,N_7926);
and U8161 (N_8161,N_7794,N_7797);
nor U8162 (N_8162,N_7946,N_7916);
or U8163 (N_8163,N_7885,N_7795);
xnor U8164 (N_8164,N_7945,N_7920);
and U8165 (N_8165,N_7961,N_7875);
xnor U8166 (N_8166,N_7905,N_7889);
nor U8167 (N_8167,N_7831,N_7897);
and U8168 (N_8168,N_7889,N_7982);
and U8169 (N_8169,N_7925,N_7964);
and U8170 (N_8170,N_7848,N_7969);
nand U8171 (N_8171,N_7857,N_7986);
or U8172 (N_8172,N_7854,N_7828);
and U8173 (N_8173,N_7759,N_7932);
nor U8174 (N_8174,N_7811,N_7807);
or U8175 (N_8175,N_7820,N_7810);
or U8176 (N_8176,N_7839,N_7890);
nand U8177 (N_8177,N_7932,N_7837);
xnor U8178 (N_8178,N_7947,N_7912);
nand U8179 (N_8179,N_7753,N_7891);
or U8180 (N_8180,N_7995,N_7950);
nand U8181 (N_8181,N_7898,N_7870);
nand U8182 (N_8182,N_7844,N_7974);
nor U8183 (N_8183,N_7964,N_7847);
or U8184 (N_8184,N_7930,N_7870);
or U8185 (N_8185,N_7772,N_7915);
nor U8186 (N_8186,N_7883,N_7845);
nor U8187 (N_8187,N_7971,N_7970);
xor U8188 (N_8188,N_7842,N_7861);
or U8189 (N_8189,N_7832,N_7997);
and U8190 (N_8190,N_7796,N_7887);
xnor U8191 (N_8191,N_7841,N_7760);
nor U8192 (N_8192,N_7785,N_7911);
nand U8193 (N_8193,N_7895,N_7828);
nor U8194 (N_8194,N_7978,N_7845);
and U8195 (N_8195,N_7875,N_7842);
xor U8196 (N_8196,N_7872,N_7891);
or U8197 (N_8197,N_7926,N_7859);
xor U8198 (N_8198,N_7949,N_7856);
nand U8199 (N_8199,N_7891,N_7949);
nor U8200 (N_8200,N_7982,N_7943);
and U8201 (N_8201,N_7781,N_7960);
nor U8202 (N_8202,N_7982,N_7862);
xor U8203 (N_8203,N_7840,N_7810);
and U8204 (N_8204,N_7761,N_7855);
nand U8205 (N_8205,N_7879,N_7964);
and U8206 (N_8206,N_7868,N_7846);
and U8207 (N_8207,N_7782,N_7999);
xor U8208 (N_8208,N_7920,N_7990);
or U8209 (N_8209,N_7830,N_7941);
and U8210 (N_8210,N_7894,N_7770);
or U8211 (N_8211,N_7930,N_7952);
xnor U8212 (N_8212,N_7799,N_7905);
nor U8213 (N_8213,N_7990,N_7974);
nor U8214 (N_8214,N_7796,N_7856);
or U8215 (N_8215,N_7858,N_7751);
xor U8216 (N_8216,N_7831,N_7816);
nand U8217 (N_8217,N_7945,N_7873);
and U8218 (N_8218,N_7870,N_7917);
and U8219 (N_8219,N_7759,N_7999);
xnor U8220 (N_8220,N_7951,N_7943);
or U8221 (N_8221,N_7982,N_7822);
xor U8222 (N_8222,N_7865,N_7874);
nand U8223 (N_8223,N_7882,N_7821);
nand U8224 (N_8224,N_7775,N_7959);
and U8225 (N_8225,N_7795,N_7766);
or U8226 (N_8226,N_7838,N_7805);
nor U8227 (N_8227,N_7759,N_7845);
nand U8228 (N_8228,N_7792,N_7926);
and U8229 (N_8229,N_7777,N_7965);
nand U8230 (N_8230,N_7888,N_7968);
and U8231 (N_8231,N_7784,N_7756);
xor U8232 (N_8232,N_7968,N_7796);
nand U8233 (N_8233,N_7953,N_7924);
nand U8234 (N_8234,N_7868,N_7763);
nand U8235 (N_8235,N_7971,N_7851);
and U8236 (N_8236,N_7785,N_7960);
nand U8237 (N_8237,N_7775,N_7807);
or U8238 (N_8238,N_7993,N_7786);
xor U8239 (N_8239,N_7889,N_7979);
nor U8240 (N_8240,N_7935,N_7808);
nand U8241 (N_8241,N_7978,N_7896);
nor U8242 (N_8242,N_7818,N_7987);
and U8243 (N_8243,N_7970,N_7925);
xor U8244 (N_8244,N_7947,N_7750);
nor U8245 (N_8245,N_7984,N_7824);
xnor U8246 (N_8246,N_7969,N_7917);
or U8247 (N_8247,N_7922,N_7842);
or U8248 (N_8248,N_7856,N_7932);
nor U8249 (N_8249,N_7907,N_7900);
nand U8250 (N_8250,N_8124,N_8071);
xor U8251 (N_8251,N_8165,N_8099);
and U8252 (N_8252,N_8239,N_8152);
and U8253 (N_8253,N_8035,N_8241);
nor U8254 (N_8254,N_8063,N_8129);
nand U8255 (N_8255,N_8147,N_8174);
or U8256 (N_8256,N_8108,N_8137);
and U8257 (N_8257,N_8172,N_8224);
or U8258 (N_8258,N_8185,N_8150);
and U8259 (N_8259,N_8193,N_8164);
or U8260 (N_8260,N_8131,N_8000);
nor U8261 (N_8261,N_8092,N_8078);
nand U8262 (N_8262,N_8113,N_8168);
nand U8263 (N_8263,N_8076,N_8018);
xor U8264 (N_8264,N_8153,N_8187);
or U8265 (N_8265,N_8162,N_8097);
nor U8266 (N_8266,N_8114,N_8080);
and U8267 (N_8267,N_8064,N_8013);
or U8268 (N_8268,N_8049,N_8221);
and U8269 (N_8269,N_8149,N_8095);
nand U8270 (N_8270,N_8236,N_8121);
nor U8271 (N_8271,N_8040,N_8222);
and U8272 (N_8272,N_8161,N_8214);
or U8273 (N_8273,N_8183,N_8053);
nand U8274 (N_8274,N_8192,N_8186);
nand U8275 (N_8275,N_8085,N_8034);
xor U8276 (N_8276,N_8238,N_8247);
and U8277 (N_8277,N_8144,N_8138);
nor U8278 (N_8278,N_8205,N_8202);
nand U8279 (N_8279,N_8115,N_8022);
nor U8280 (N_8280,N_8096,N_8154);
and U8281 (N_8281,N_8079,N_8216);
or U8282 (N_8282,N_8060,N_8048);
nand U8283 (N_8283,N_8190,N_8191);
xor U8284 (N_8284,N_8234,N_8180);
xnor U8285 (N_8285,N_8089,N_8188);
nand U8286 (N_8286,N_8225,N_8005);
xnor U8287 (N_8287,N_8014,N_8036);
nand U8288 (N_8288,N_8201,N_8230);
nand U8289 (N_8289,N_8133,N_8056);
xnor U8290 (N_8290,N_8066,N_8118);
nor U8291 (N_8291,N_8226,N_8062);
nor U8292 (N_8292,N_8041,N_8123);
or U8293 (N_8293,N_8102,N_8173);
or U8294 (N_8294,N_8128,N_8110);
nand U8295 (N_8295,N_8098,N_8002);
xor U8296 (N_8296,N_8194,N_8126);
xor U8297 (N_8297,N_8181,N_8227);
or U8298 (N_8298,N_8101,N_8052);
nor U8299 (N_8299,N_8009,N_8196);
nor U8300 (N_8300,N_8015,N_8065);
xor U8301 (N_8301,N_8011,N_8215);
and U8302 (N_8302,N_8231,N_8037);
nand U8303 (N_8303,N_8244,N_8004);
nor U8304 (N_8304,N_8045,N_8033);
or U8305 (N_8305,N_8130,N_8090);
or U8306 (N_8306,N_8019,N_8136);
xor U8307 (N_8307,N_8243,N_8142);
or U8308 (N_8308,N_8182,N_8039);
xor U8309 (N_8309,N_8167,N_8135);
xnor U8310 (N_8310,N_8209,N_8184);
and U8311 (N_8311,N_8139,N_8074);
nand U8312 (N_8312,N_8070,N_8237);
xnor U8313 (N_8313,N_8158,N_8017);
xnor U8314 (N_8314,N_8051,N_8067);
or U8315 (N_8315,N_8068,N_8169);
nor U8316 (N_8316,N_8111,N_8246);
nand U8317 (N_8317,N_8020,N_8151);
and U8318 (N_8318,N_8025,N_8116);
nand U8319 (N_8319,N_8177,N_8054);
nand U8320 (N_8320,N_8106,N_8103);
nand U8321 (N_8321,N_8105,N_8026);
and U8322 (N_8322,N_8204,N_8178);
or U8323 (N_8323,N_8044,N_8038);
xor U8324 (N_8324,N_8094,N_8240);
nor U8325 (N_8325,N_8117,N_8175);
nor U8326 (N_8326,N_8072,N_8112);
or U8327 (N_8327,N_8145,N_8132);
xor U8328 (N_8328,N_8200,N_8248);
xor U8329 (N_8329,N_8213,N_8061);
nand U8330 (N_8330,N_8206,N_8077);
and U8331 (N_8331,N_8107,N_8197);
and U8332 (N_8332,N_8219,N_8104);
and U8333 (N_8333,N_8125,N_8143);
nor U8334 (N_8334,N_8083,N_8228);
or U8335 (N_8335,N_8203,N_8134);
nand U8336 (N_8336,N_8127,N_8028);
or U8337 (N_8337,N_8050,N_8159);
or U8338 (N_8338,N_8058,N_8043);
xnor U8339 (N_8339,N_8171,N_8001);
nand U8340 (N_8340,N_8047,N_8086);
and U8341 (N_8341,N_8176,N_8082);
and U8342 (N_8342,N_8217,N_8208);
xnor U8343 (N_8343,N_8235,N_8008);
and U8344 (N_8344,N_8223,N_8218);
xnor U8345 (N_8345,N_8032,N_8093);
nor U8346 (N_8346,N_8030,N_8024);
nand U8347 (N_8347,N_8179,N_8109);
xor U8348 (N_8348,N_8245,N_8091);
nor U8349 (N_8349,N_8211,N_8199);
xor U8350 (N_8350,N_8046,N_8189);
or U8351 (N_8351,N_8170,N_8055);
xnor U8352 (N_8352,N_8073,N_8003);
and U8353 (N_8353,N_8232,N_8119);
nor U8354 (N_8354,N_8023,N_8195);
and U8355 (N_8355,N_8029,N_8057);
and U8356 (N_8356,N_8087,N_8075);
and U8357 (N_8357,N_8081,N_8146);
nor U8358 (N_8358,N_8198,N_8156);
nor U8359 (N_8359,N_8016,N_8031);
nand U8360 (N_8360,N_8042,N_8212);
nor U8361 (N_8361,N_8021,N_8207);
nand U8362 (N_8362,N_8084,N_8166);
and U8363 (N_8363,N_8233,N_8100);
nand U8364 (N_8364,N_8242,N_8140);
or U8365 (N_8365,N_8229,N_8160);
nor U8366 (N_8366,N_8210,N_8012);
xor U8367 (N_8367,N_8157,N_8148);
nand U8368 (N_8368,N_8006,N_8155);
and U8369 (N_8369,N_8010,N_8122);
xnor U8370 (N_8370,N_8069,N_8249);
and U8371 (N_8371,N_8141,N_8088);
nand U8372 (N_8372,N_8007,N_8163);
nand U8373 (N_8373,N_8059,N_8220);
nand U8374 (N_8374,N_8120,N_8027);
nand U8375 (N_8375,N_8176,N_8096);
and U8376 (N_8376,N_8231,N_8244);
nor U8377 (N_8377,N_8145,N_8019);
or U8378 (N_8378,N_8242,N_8041);
and U8379 (N_8379,N_8216,N_8157);
xnor U8380 (N_8380,N_8188,N_8017);
or U8381 (N_8381,N_8071,N_8048);
nand U8382 (N_8382,N_8208,N_8126);
or U8383 (N_8383,N_8112,N_8046);
nand U8384 (N_8384,N_8016,N_8208);
nor U8385 (N_8385,N_8067,N_8101);
nor U8386 (N_8386,N_8044,N_8191);
nand U8387 (N_8387,N_8036,N_8047);
nor U8388 (N_8388,N_8163,N_8229);
xor U8389 (N_8389,N_8070,N_8235);
and U8390 (N_8390,N_8198,N_8073);
or U8391 (N_8391,N_8015,N_8159);
nor U8392 (N_8392,N_8197,N_8210);
or U8393 (N_8393,N_8168,N_8211);
and U8394 (N_8394,N_8226,N_8160);
nor U8395 (N_8395,N_8243,N_8093);
xor U8396 (N_8396,N_8120,N_8001);
nor U8397 (N_8397,N_8232,N_8009);
and U8398 (N_8398,N_8242,N_8070);
or U8399 (N_8399,N_8230,N_8221);
or U8400 (N_8400,N_8047,N_8045);
xnor U8401 (N_8401,N_8088,N_8106);
nand U8402 (N_8402,N_8058,N_8123);
nor U8403 (N_8403,N_8185,N_8124);
or U8404 (N_8404,N_8172,N_8242);
or U8405 (N_8405,N_8224,N_8182);
nand U8406 (N_8406,N_8137,N_8157);
xor U8407 (N_8407,N_8221,N_8194);
nand U8408 (N_8408,N_8053,N_8218);
or U8409 (N_8409,N_8031,N_8070);
xnor U8410 (N_8410,N_8150,N_8044);
nor U8411 (N_8411,N_8174,N_8127);
xnor U8412 (N_8412,N_8239,N_8211);
nand U8413 (N_8413,N_8231,N_8104);
nand U8414 (N_8414,N_8101,N_8054);
and U8415 (N_8415,N_8194,N_8116);
nor U8416 (N_8416,N_8206,N_8194);
and U8417 (N_8417,N_8045,N_8228);
or U8418 (N_8418,N_8184,N_8211);
xor U8419 (N_8419,N_8173,N_8120);
nand U8420 (N_8420,N_8124,N_8233);
xor U8421 (N_8421,N_8137,N_8152);
nor U8422 (N_8422,N_8089,N_8011);
or U8423 (N_8423,N_8143,N_8224);
xnor U8424 (N_8424,N_8155,N_8150);
xnor U8425 (N_8425,N_8231,N_8092);
or U8426 (N_8426,N_8200,N_8184);
nor U8427 (N_8427,N_8192,N_8246);
nor U8428 (N_8428,N_8222,N_8014);
xor U8429 (N_8429,N_8097,N_8095);
or U8430 (N_8430,N_8240,N_8117);
xnor U8431 (N_8431,N_8238,N_8234);
nor U8432 (N_8432,N_8120,N_8000);
nor U8433 (N_8433,N_8198,N_8166);
and U8434 (N_8434,N_8038,N_8136);
xnor U8435 (N_8435,N_8066,N_8021);
xnor U8436 (N_8436,N_8045,N_8098);
and U8437 (N_8437,N_8180,N_8193);
and U8438 (N_8438,N_8034,N_8057);
xor U8439 (N_8439,N_8230,N_8209);
or U8440 (N_8440,N_8186,N_8121);
nand U8441 (N_8441,N_8224,N_8236);
xor U8442 (N_8442,N_8152,N_8202);
nor U8443 (N_8443,N_8116,N_8216);
xnor U8444 (N_8444,N_8155,N_8232);
nor U8445 (N_8445,N_8146,N_8205);
xor U8446 (N_8446,N_8023,N_8177);
and U8447 (N_8447,N_8028,N_8189);
nor U8448 (N_8448,N_8094,N_8024);
and U8449 (N_8449,N_8030,N_8228);
or U8450 (N_8450,N_8204,N_8048);
or U8451 (N_8451,N_8071,N_8013);
nor U8452 (N_8452,N_8166,N_8139);
or U8453 (N_8453,N_8176,N_8188);
xor U8454 (N_8454,N_8067,N_8215);
or U8455 (N_8455,N_8121,N_8016);
or U8456 (N_8456,N_8249,N_8132);
xnor U8457 (N_8457,N_8015,N_8110);
nor U8458 (N_8458,N_8131,N_8053);
xor U8459 (N_8459,N_8089,N_8224);
nand U8460 (N_8460,N_8068,N_8186);
nor U8461 (N_8461,N_8042,N_8140);
xor U8462 (N_8462,N_8023,N_8163);
or U8463 (N_8463,N_8176,N_8195);
nor U8464 (N_8464,N_8165,N_8035);
and U8465 (N_8465,N_8162,N_8023);
nand U8466 (N_8466,N_8106,N_8002);
xor U8467 (N_8467,N_8019,N_8174);
xnor U8468 (N_8468,N_8003,N_8023);
or U8469 (N_8469,N_8196,N_8021);
xor U8470 (N_8470,N_8232,N_8094);
and U8471 (N_8471,N_8119,N_8245);
nor U8472 (N_8472,N_8101,N_8120);
nand U8473 (N_8473,N_8203,N_8052);
nor U8474 (N_8474,N_8042,N_8244);
and U8475 (N_8475,N_8010,N_8011);
nand U8476 (N_8476,N_8160,N_8047);
and U8477 (N_8477,N_8116,N_8018);
xor U8478 (N_8478,N_8216,N_8243);
xnor U8479 (N_8479,N_8161,N_8219);
xnor U8480 (N_8480,N_8145,N_8242);
or U8481 (N_8481,N_8201,N_8060);
and U8482 (N_8482,N_8229,N_8134);
nand U8483 (N_8483,N_8176,N_8141);
nor U8484 (N_8484,N_8197,N_8190);
nand U8485 (N_8485,N_8216,N_8093);
nor U8486 (N_8486,N_8158,N_8047);
xor U8487 (N_8487,N_8164,N_8073);
nand U8488 (N_8488,N_8210,N_8193);
xnor U8489 (N_8489,N_8235,N_8005);
nand U8490 (N_8490,N_8089,N_8019);
nand U8491 (N_8491,N_8014,N_8247);
or U8492 (N_8492,N_8036,N_8164);
or U8493 (N_8493,N_8232,N_8111);
nor U8494 (N_8494,N_8144,N_8073);
or U8495 (N_8495,N_8187,N_8081);
and U8496 (N_8496,N_8063,N_8047);
and U8497 (N_8497,N_8145,N_8130);
and U8498 (N_8498,N_8004,N_8005);
or U8499 (N_8499,N_8110,N_8184);
nor U8500 (N_8500,N_8412,N_8388);
and U8501 (N_8501,N_8491,N_8423);
xor U8502 (N_8502,N_8276,N_8429);
nor U8503 (N_8503,N_8393,N_8335);
nor U8504 (N_8504,N_8366,N_8382);
nand U8505 (N_8505,N_8442,N_8403);
nand U8506 (N_8506,N_8496,N_8258);
and U8507 (N_8507,N_8375,N_8309);
nand U8508 (N_8508,N_8401,N_8459);
xor U8509 (N_8509,N_8386,N_8292);
nand U8510 (N_8510,N_8457,N_8436);
or U8511 (N_8511,N_8390,N_8415);
xnor U8512 (N_8512,N_8367,N_8354);
xnor U8513 (N_8513,N_8279,N_8325);
nand U8514 (N_8514,N_8339,N_8431);
nor U8515 (N_8515,N_8322,N_8396);
xor U8516 (N_8516,N_8263,N_8448);
nand U8517 (N_8517,N_8430,N_8348);
xor U8518 (N_8518,N_8266,N_8372);
and U8519 (N_8519,N_8444,N_8418);
nor U8520 (N_8520,N_8398,N_8499);
xnor U8521 (N_8521,N_8482,N_8338);
and U8522 (N_8522,N_8283,N_8441);
and U8523 (N_8523,N_8282,N_8397);
or U8524 (N_8524,N_8460,N_8255);
nor U8525 (N_8525,N_8288,N_8497);
and U8526 (N_8526,N_8356,N_8463);
and U8527 (N_8527,N_8410,N_8449);
nand U8528 (N_8528,N_8378,N_8387);
xnor U8529 (N_8529,N_8296,N_8456);
nand U8530 (N_8530,N_8370,N_8297);
xor U8531 (N_8531,N_8329,N_8452);
nand U8532 (N_8532,N_8307,N_8399);
nand U8533 (N_8533,N_8473,N_8477);
or U8534 (N_8534,N_8392,N_8351);
and U8535 (N_8535,N_8250,N_8349);
or U8536 (N_8536,N_8376,N_8394);
nor U8537 (N_8537,N_8285,N_8373);
or U8538 (N_8538,N_8346,N_8336);
nand U8539 (N_8539,N_8293,N_8432);
and U8540 (N_8540,N_8280,N_8369);
and U8541 (N_8541,N_8332,N_8414);
nor U8542 (N_8542,N_8271,N_8467);
and U8543 (N_8543,N_8284,N_8486);
nand U8544 (N_8544,N_8447,N_8357);
nor U8545 (N_8545,N_8433,N_8417);
and U8546 (N_8546,N_8440,N_8313);
xor U8547 (N_8547,N_8331,N_8384);
or U8548 (N_8548,N_8303,N_8438);
xor U8549 (N_8549,N_8321,N_8278);
nor U8550 (N_8550,N_8466,N_8264);
and U8551 (N_8551,N_8379,N_8454);
nand U8552 (N_8552,N_8419,N_8330);
xnor U8553 (N_8553,N_8352,N_8395);
nand U8554 (N_8554,N_8317,N_8341);
xor U8555 (N_8555,N_8295,N_8286);
or U8556 (N_8556,N_8406,N_8474);
or U8557 (N_8557,N_8385,N_8408);
or U8558 (N_8558,N_8480,N_8362);
nand U8559 (N_8559,N_8298,N_8475);
xnor U8560 (N_8560,N_8453,N_8261);
nor U8561 (N_8561,N_8306,N_8450);
nor U8562 (N_8562,N_8363,N_8377);
xor U8563 (N_8563,N_8439,N_8407);
nor U8564 (N_8564,N_8365,N_8305);
xor U8565 (N_8565,N_8492,N_8358);
nand U8566 (N_8566,N_8424,N_8257);
xnor U8567 (N_8567,N_8252,N_8490);
nand U8568 (N_8568,N_8402,N_8316);
xnor U8569 (N_8569,N_8371,N_8471);
nand U8570 (N_8570,N_8272,N_8267);
and U8571 (N_8571,N_8333,N_8485);
nor U8572 (N_8572,N_8269,N_8484);
nor U8573 (N_8573,N_8327,N_8312);
and U8574 (N_8574,N_8347,N_8380);
nand U8575 (N_8575,N_8302,N_8355);
or U8576 (N_8576,N_8319,N_8479);
xor U8577 (N_8577,N_8400,N_8361);
nand U8578 (N_8578,N_8451,N_8287);
nor U8579 (N_8579,N_8254,N_8478);
nor U8580 (N_8580,N_8334,N_8294);
nand U8581 (N_8581,N_8462,N_8498);
or U8582 (N_8582,N_8290,N_8311);
nor U8583 (N_8583,N_8323,N_8353);
nor U8584 (N_8584,N_8445,N_8281);
xor U8585 (N_8585,N_8315,N_8337);
or U8586 (N_8586,N_8262,N_8383);
nand U8587 (N_8587,N_8318,N_8324);
nand U8588 (N_8588,N_8320,N_8259);
and U8589 (N_8589,N_8268,N_8344);
or U8590 (N_8590,N_8273,N_8340);
nor U8591 (N_8591,N_8308,N_8472);
or U8592 (N_8592,N_8343,N_8304);
xor U8593 (N_8593,N_8291,N_8469);
xor U8594 (N_8594,N_8251,N_8435);
xor U8595 (N_8595,N_8404,N_8494);
or U8596 (N_8596,N_8416,N_8381);
nand U8597 (N_8597,N_8481,N_8487);
or U8598 (N_8598,N_8277,N_8265);
or U8599 (N_8599,N_8405,N_8326);
xor U8600 (N_8600,N_8443,N_8495);
nor U8601 (N_8601,N_8256,N_8270);
nand U8602 (N_8602,N_8488,N_8458);
nor U8603 (N_8603,N_8425,N_8300);
nor U8604 (N_8604,N_8374,N_8391);
and U8605 (N_8605,N_8476,N_8428);
nand U8606 (N_8606,N_8389,N_8253);
nand U8607 (N_8607,N_8470,N_8345);
xnor U8608 (N_8608,N_8350,N_8489);
and U8609 (N_8609,N_8420,N_8411);
or U8610 (N_8610,N_8328,N_8422);
nor U8611 (N_8611,N_8299,N_8434);
and U8612 (N_8612,N_8342,N_8289);
or U8613 (N_8613,N_8360,N_8301);
or U8614 (N_8614,N_8409,N_8455);
nand U8615 (N_8615,N_8465,N_8461);
or U8616 (N_8616,N_8437,N_8274);
nand U8617 (N_8617,N_8310,N_8483);
xor U8618 (N_8618,N_8464,N_8468);
xnor U8619 (N_8619,N_8364,N_8427);
or U8620 (N_8620,N_8493,N_8413);
and U8621 (N_8621,N_8446,N_8368);
and U8622 (N_8622,N_8275,N_8359);
or U8623 (N_8623,N_8426,N_8421);
nor U8624 (N_8624,N_8314,N_8260);
nor U8625 (N_8625,N_8476,N_8344);
xnor U8626 (N_8626,N_8394,N_8314);
nor U8627 (N_8627,N_8425,N_8282);
nand U8628 (N_8628,N_8443,N_8354);
nor U8629 (N_8629,N_8330,N_8392);
and U8630 (N_8630,N_8353,N_8428);
xor U8631 (N_8631,N_8327,N_8389);
nor U8632 (N_8632,N_8463,N_8349);
xor U8633 (N_8633,N_8259,N_8395);
nand U8634 (N_8634,N_8353,N_8264);
nor U8635 (N_8635,N_8356,N_8460);
and U8636 (N_8636,N_8459,N_8285);
nand U8637 (N_8637,N_8376,N_8300);
or U8638 (N_8638,N_8466,N_8405);
nor U8639 (N_8639,N_8324,N_8339);
or U8640 (N_8640,N_8250,N_8446);
xnor U8641 (N_8641,N_8361,N_8350);
or U8642 (N_8642,N_8323,N_8423);
nor U8643 (N_8643,N_8499,N_8408);
nand U8644 (N_8644,N_8315,N_8318);
or U8645 (N_8645,N_8282,N_8320);
nor U8646 (N_8646,N_8417,N_8331);
or U8647 (N_8647,N_8347,N_8359);
nor U8648 (N_8648,N_8350,N_8385);
or U8649 (N_8649,N_8450,N_8305);
nand U8650 (N_8650,N_8272,N_8310);
xnor U8651 (N_8651,N_8358,N_8399);
xor U8652 (N_8652,N_8268,N_8428);
or U8653 (N_8653,N_8259,N_8427);
and U8654 (N_8654,N_8300,N_8307);
nand U8655 (N_8655,N_8267,N_8419);
or U8656 (N_8656,N_8449,N_8367);
and U8657 (N_8657,N_8459,N_8383);
or U8658 (N_8658,N_8407,N_8358);
or U8659 (N_8659,N_8350,N_8309);
nand U8660 (N_8660,N_8304,N_8367);
or U8661 (N_8661,N_8431,N_8403);
nand U8662 (N_8662,N_8393,N_8315);
or U8663 (N_8663,N_8481,N_8384);
and U8664 (N_8664,N_8376,N_8378);
nand U8665 (N_8665,N_8302,N_8485);
nand U8666 (N_8666,N_8325,N_8430);
nand U8667 (N_8667,N_8354,N_8391);
nor U8668 (N_8668,N_8255,N_8414);
nor U8669 (N_8669,N_8476,N_8327);
or U8670 (N_8670,N_8322,N_8457);
nor U8671 (N_8671,N_8474,N_8329);
nand U8672 (N_8672,N_8493,N_8481);
nor U8673 (N_8673,N_8273,N_8443);
or U8674 (N_8674,N_8350,N_8317);
or U8675 (N_8675,N_8433,N_8480);
xnor U8676 (N_8676,N_8475,N_8395);
and U8677 (N_8677,N_8281,N_8375);
or U8678 (N_8678,N_8495,N_8316);
nor U8679 (N_8679,N_8257,N_8486);
and U8680 (N_8680,N_8340,N_8492);
nand U8681 (N_8681,N_8494,N_8458);
nor U8682 (N_8682,N_8273,N_8274);
xnor U8683 (N_8683,N_8280,N_8260);
or U8684 (N_8684,N_8318,N_8305);
nor U8685 (N_8685,N_8483,N_8291);
nand U8686 (N_8686,N_8390,N_8387);
xor U8687 (N_8687,N_8406,N_8440);
xnor U8688 (N_8688,N_8434,N_8341);
and U8689 (N_8689,N_8364,N_8316);
and U8690 (N_8690,N_8322,N_8492);
and U8691 (N_8691,N_8295,N_8375);
nand U8692 (N_8692,N_8292,N_8425);
xor U8693 (N_8693,N_8391,N_8301);
nor U8694 (N_8694,N_8409,N_8456);
xnor U8695 (N_8695,N_8299,N_8425);
nor U8696 (N_8696,N_8465,N_8346);
nand U8697 (N_8697,N_8259,N_8336);
nor U8698 (N_8698,N_8279,N_8347);
and U8699 (N_8699,N_8348,N_8477);
nor U8700 (N_8700,N_8377,N_8289);
and U8701 (N_8701,N_8474,N_8318);
or U8702 (N_8702,N_8489,N_8319);
nor U8703 (N_8703,N_8458,N_8472);
xor U8704 (N_8704,N_8452,N_8436);
or U8705 (N_8705,N_8273,N_8260);
nand U8706 (N_8706,N_8388,N_8492);
nor U8707 (N_8707,N_8279,N_8337);
nand U8708 (N_8708,N_8284,N_8386);
nand U8709 (N_8709,N_8446,N_8479);
and U8710 (N_8710,N_8283,N_8258);
nor U8711 (N_8711,N_8421,N_8255);
nand U8712 (N_8712,N_8327,N_8293);
nor U8713 (N_8713,N_8388,N_8422);
xnor U8714 (N_8714,N_8402,N_8344);
nand U8715 (N_8715,N_8456,N_8402);
or U8716 (N_8716,N_8423,N_8429);
and U8717 (N_8717,N_8430,N_8307);
and U8718 (N_8718,N_8400,N_8320);
nand U8719 (N_8719,N_8371,N_8402);
nor U8720 (N_8720,N_8468,N_8299);
nand U8721 (N_8721,N_8485,N_8336);
or U8722 (N_8722,N_8364,N_8308);
or U8723 (N_8723,N_8487,N_8276);
and U8724 (N_8724,N_8415,N_8312);
xor U8725 (N_8725,N_8468,N_8264);
nand U8726 (N_8726,N_8425,N_8418);
and U8727 (N_8727,N_8273,N_8257);
or U8728 (N_8728,N_8272,N_8359);
nor U8729 (N_8729,N_8496,N_8432);
nor U8730 (N_8730,N_8321,N_8387);
or U8731 (N_8731,N_8288,N_8457);
nand U8732 (N_8732,N_8412,N_8298);
nor U8733 (N_8733,N_8255,N_8304);
and U8734 (N_8734,N_8288,N_8483);
nor U8735 (N_8735,N_8381,N_8349);
xnor U8736 (N_8736,N_8484,N_8305);
or U8737 (N_8737,N_8403,N_8260);
xor U8738 (N_8738,N_8379,N_8469);
or U8739 (N_8739,N_8321,N_8406);
xnor U8740 (N_8740,N_8474,N_8384);
xor U8741 (N_8741,N_8341,N_8250);
nand U8742 (N_8742,N_8294,N_8459);
or U8743 (N_8743,N_8420,N_8415);
xnor U8744 (N_8744,N_8401,N_8476);
or U8745 (N_8745,N_8369,N_8449);
xnor U8746 (N_8746,N_8381,N_8360);
and U8747 (N_8747,N_8341,N_8308);
nand U8748 (N_8748,N_8274,N_8430);
or U8749 (N_8749,N_8399,N_8299);
nand U8750 (N_8750,N_8546,N_8558);
or U8751 (N_8751,N_8608,N_8643);
or U8752 (N_8752,N_8710,N_8619);
or U8753 (N_8753,N_8574,N_8629);
or U8754 (N_8754,N_8731,N_8718);
nand U8755 (N_8755,N_8585,N_8715);
and U8756 (N_8756,N_8571,N_8651);
nand U8757 (N_8757,N_8527,N_8559);
or U8758 (N_8758,N_8600,N_8696);
or U8759 (N_8759,N_8662,N_8632);
and U8760 (N_8760,N_8598,N_8602);
or U8761 (N_8761,N_8562,N_8576);
nand U8762 (N_8762,N_8513,N_8644);
xor U8763 (N_8763,N_8594,N_8508);
xnor U8764 (N_8764,N_8541,N_8504);
nor U8765 (N_8765,N_8523,N_8519);
nor U8766 (N_8766,N_8698,N_8742);
and U8767 (N_8767,N_8590,N_8681);
nor U8768 (N_8768,N_8617,N_8635);
nand U8769 (N_8769,N_8631,N_8645);
xor U8770 (N_8770,N_8653,N_8704);
xnor U8771 (N_8771,N_8621,N_8539);
or U8772 (N_8772,N_8609,N_8737);
and U8773 (N_8773,N_8568,N_8693);
or U8774 (N_8774,N_8599,N_8553);
xnor U8775 (N_8775,N_8666,N_8663);
and U8776 (N_8776,N_8616,N_8569);
nor U8777 (N_8777,N_8642,N_8531);
nand U8778 (N_8778,N_8661,N_8684);
and U8779 (N_8779,N_8687,N_8689);
nand U8780 (N_8780,N_8591,N_8540);
or U8781 (N_8781,N_8507,N_8564);
nand U8782 (N_8782,N_8575,N_8589);
nand U8783 (N_8783,N_8528,N_8677);
xnor U8784 (N_8784,N_8727,N_8695);
nor U8785 (N_8785,N_8669,N_8622);
xor U8786 (N_8786,N_8694,N_8554);
or U8787 (N_8787,N_8724,N_8707);
nand U8788 (N_8788,N_8510,N_8530);
nor U8789 (N_8789,N_8538,N_8665);
or U8790 (N_8790,N_8518,N_8536);
and U8791 (N_8791,N_8676,N_8570);
or U8792 (N_8792,N_8537,N_8650);
nand U8793 (N_8793,N_8579,N_8683);
or U8794 (N_8794,N_8743,N_8603);
or U8795 (N_8795,N_8521,N_8713);
nand U8796 (N_8796,N_8675,N_8514);
xor U8797 (N_8797,N_8620,N_8749);
nor U8798 (N_8798,N_8601,N_8702);
nor U8799 (N_8799,N_8748,N_8655);
nor U8800 (N_8800,N_8592,N_8593);
or U8801 (N_8801,N_8506,N_8596);
and U8802 (N_8802,N_8691,N_8744);
and U8803 (N_8803,N_8573,N_8646);
or U8804 (N_8804,N_8685,N_8544);
xnor U8805 (N_8805,N_8734,N_8723);
and U8806 (N_8806,N_8709,N_8517);
and U8807 (N_8807,N_8630,N_8648);
and U8808 (N_8808,N_8658,N_8726);
or U8809 (N_8809,N_8548,N_8736);
or U8810 (N_8810,N_8706,N_8674);
nor U8811 (N_8811,N_8740,N_8595);
and U8812 (N_8812,N_8529,N_8547);
nor U8813 (N_8813,N_8533,N_8522);
xnor U8814 (N_8814,N_8636,N_8634);
nor U8815 (N_8815,N_8668,N_8584);
and U8816 (N_8816,N_8586,N_8543);
nor U8817 (N_8817,N_8515,N_8690);
xnor U8818 (N_8818,N_8664,N_8625);
nor U8819 (N_8819,N_8733,N_8532);
xor U8820 (N_8820,N_8587,N_8534);
nand U8821 (N_8821,N_8561,N_8551);
and U8822 (N_8822,N_8500,N_8671);
nor U8823 (N_8823,N_8652,N_8745);
nand U8824 (N_8824,N_8607,N_8626);
and U8825 (N_8825,N_8699,N_8667);
or U8826 (N_8826,N_8509,N_8720);
nor U8827 (N_8827,N_8552,N_8578);
or U8828 (N_8828,N_8739,N_8638);
and U8829 (N_8829,N_8612,N_8682);
nor U8830 (N_8830,N_8679,N_8660);
xnor U8831 (N_8831,N_8588,N_8728);
nor U8832 (N_8832,N_8637,N_8633);
xnor U8833 (N_8833,N_8639,N_8566);
or U8834 (N_8834,N_8673,N_8716);
xor U8835 (N_8835,N_8618,N_8557);
nor U8836 (N_8836,N_8567,N_8501);
nor U8837 (N_8837,N_8511,N_8611);
xor U8838 (N_8838,N_8697,N_8725);
or U8839 (N_8839,N_8613,N_8678);
nand U8840 (N_8840,N_8746,N_8657);
xor U8841 (N_8841,N_8555,N_8605);
nor U8842 (N_8842,N_8708,N_8512);
or U8843 (N_8843,N_8714,N_8535);
or U8844 (N_8844,N_8692,N_8542);
xnor U8845 (N_8845,N_8525,N_8526);
or U8846 (N_8846,N_8717,N_8701);
or U8847 (N_8847,N_8721,N_8516);
nand U8848 (N_8848,N_8628,N_8577);
or U8849 (N_8849,N_8583,N_8623);
or U8850 (N_8850,N_8520,N_8641);
nand U8851 (N_8851,N_8560,N_8680);
and U8852 (N_8852,N_8703,N_8700);
and U8853 (N_8853,N_8670,N_8624);
xnor U8854 (N_8854,N_8615,N_8572);
or U8855 (N_8855,N_8705,N_8741);
nor U8856 (N_8856,N_8565,N_8604);
nor U8857 (N_8857,N_8719,N_8581);
xor U8858 (N_8858,N_8580,N_8505);
nand U8859 (N_8859,N_8627,N_8549);
and U8860 (N_8860,N_8647,N_8640);
and U8861 (N_8861,N_8656,N_8672);
nor U8862 (N_8862,N_8556,N_8606);
nor U8863 (N_8863,N_8735,N_8503);
xor U8864 (N_8864,N_8610,N_8688);
xnor U8865 (N_8865,N_8738,N_8729);
nor U8866 (N_8866,N_8524,N_8582);
xnor U8867 (N_8867,N_8732,N_8614);
xor U8868 (N_8868,N_8550,N_8545);
nor U8869 (N_8869,N_8649,N_8502);
or U8870 (N_8870,N_8711,N_8712);
nand U8871 (N_8871,N_8747,N_8686);
nand U8872 (N_8872,N_8730,N_8563);
nand U8873 (N_8873,N_8722,N_8659);
nor U8874 (N_8874,N_8597,N_8654);
nand U8875 (N_8875,N_8559,N_8668);
xnor U8876 (N_8876,N_8527,N_8612);
nor U8877 (N_8877,N_8503,N_8571);
and U8878 (N_8878,N_8693,N_8731);
and U8879 (N_8879,N_8540,N_8663);
xnor U8880 (N_8880,N_8589,N_8698);
or U8881 (N_8881,N_8647,N_8675);
or U8882 (N_8882,N_8562,N_8627);
xor U8883 (N_8883,N_8510,N_8728);
xnor U8884 (N_8884,N_8514,N_8527);
and U8885 (N_8885,N_8668,N_8536);
and U8886 (N_8886,N_8531,N_8708);
or U8887 (N_8887,N_8606,N_8535);
and U8888 (N_8888,N_8746,N_8547);
nor U8889 (N_8889,N_8517,N_8554);
xor U8890 (N_8890,N_8667,N_8736);
or U8891 (N_8891,N_8733,N_8634);
and U8892 (N_8892,N_8714,N_8597);
xor U8893 (N_8893,N_8673,N_8612);
or U8894 (N_8894,N_8726,N_8620);
xor U8895 (N_8895,N_8519,N_8729);
or U8896 (N_8896,N_8714,N_8568);
nor U8897 (N_8897,N_8576,N_8503);
nor U8898 (N_8898,N_8616,N_8544);
nor U8899 (N_8899,N_8643,N_8588);
xor U8900 (N_8900,N_8572,N_8689);
nor U8901 (N_8901,N_8584,N_8579);
xnor U8902 (N_8902,N_8520,N_8692);
nand U8903 (N_8903,N_8515,N_8509);
nor U8904 (N_8904,N_8748,N_8719);
or U8905 (N_8905,N_8589,N_8563);
xor U8906 (N_8906,N_8624,N_8681);
or U8907 (N_8907,N_8651,N_8643);
nor U8908 (N_8908,N_8681,N_8728);
or U8909 (N_8909,N_8728,N_8676);
and U8910 (N_8910,N_8577,N_8659);
or U8911 (N_8911,N_8534,N_8547);
nand U8912 (N_8912,N_8707,N_8674);
and U8913 (N_8913,N_8641,N_8559);
nor U8914 (N_8914,N_8557,N_8625);
or U8915 (N_8915,N_8568,N_8539);
and U8916 (N_8916,N_8558,N_8606);
and U8917 (N_8917,N_8615,N_8595);
nor U8918 (N_8918,N_8638,N_8612);
nor U8919 (N_8919,N_8678,N_8662);
nand U8920 (N_8920,N_8515,N_8672);
xnor U8921 (N_8921,N_8725,N_8560);
and U8922 (N_8922,N_8599,N_8569);
and U8923 (N_8923,N_8700,N_8677);
nand U8924 (N_8924,N_8639,N_8613);
nor U8925 (N_8925,N_8570,N_8672);
and U8926 (N_8926,N_8671,N_8538);
and U8927 (N_8927,N_8556,N_8695);
nor U8928 (N_8928,N_8679,N_8646);
nor U8929 (N_8929,N_8596,N_8607);
xnor U8930 (N_8930,N_8529,N_8570);
nor U8931 (N_8931,N_8541,N_8735);
or U8932 (N_8932,N_8723,N_8602);
and U8933 (N_8933,N_8542,N_8615);
xor U8934 (N_8934,N_8602,N_8742);
xor U8935 (N_8935,N_8597,N_8598);
nor U8936 (N_8936,N_8569,N_8551);
nand U8937 (N_8937,N_8538,N_8716);
nand U8938 (N_8938,N_8592,N_8601);
or U8939 (N_8939,N_8523,N_8629);
nand U8940 (N_8940,N_8599,N_8666);
xor U8941 (N_8941,N_8597,N_8653);
xnor U8942 (N_8942,N_8641,N_8576);
nand U8943 (N_8943,N_8517,N_8628);
nor U8944 (N_8944,N_8633,N_8627);
and U8945 (N_8945,N_8642,N_8538);
nor U8946 (N_8946,N_8709,N_8569);
nor U8947 (N_8947,N_8635,N_8654);
nor U8948 (N_8948,N_8540,N_8595);
or U8949 (N_8949,N_8739,N_8732);
xnor U8950 (N_8950,N_8747,N_8645);
nor U8951 (N_8951,N_8615,N_8552);
nor U8952 (N_8952,N_8574,N_8612);
nand U8953 (N_8953,N_8563,N_8512);
and U8954 (N_8954,N_8697,N_8689);
nor U8955 (N_8955,N_8580,N_8721);
xnor U8956 (N_8956,N_8693,N_8502);
nand U8957 (N_8957,N_8714,N_8582);
or U8958 (N_8958,N_8731,N_8537);
and U8959 (N_8959,N_8516,N_8565);
and U8960 (N_8960,N_8581,N_8661);
and U8961 (N_8961,N_8599,N_8525);
nor U8962 (N_8962,N_8631,N_8604);
nand U8963 (N_8963,N_8626,N_8743);
xnor U8964 (N_8964,N_8577,N_8716);
nor U8965 (N_8965,N_8716,N_8623);
nor U8966 (N_8966,N_8745,N_8551);
nor U8967 (N_8967,N_8586,N_8682);
nand U8968 (N_8968,N_8696,N_8632);
or U8969 (N_8969,N_8612,N_8743);
xnor U8970 (N_8970,N_8671,N_8630);
or U8971 (N_8971,N_8719,N_8569);
and U8972 (N_8972,N_8557,N_8705);
xor U8973 (N_8973,N_8704,N_8712);
nor U8974 (N_8974,N_8529,N_8561);
xnor U8975 (N_8975,N_8657,N_8558);
xor U8976 (N_8976,N_8533,N_8526);
or U8977 (N_8977,N_8558,N_8711);
nand U8978 (N_8978,N_8692,N_8557);
xnor U8979 (N_8979,N_8690,N_8659);
and U8980 (N_8980,N_8606,N_8599);
or U8981 (N_8981,N_8669,N_8738);
xnor U8982 (N_8982,N_8520,N_8634);
xnor U8983 (N_8983,N_8667,N_8644);
nor U8984 (N_8984,N_8591,N_8563);
xor U8985 (N_8985,N_8718,N_8620);
xor U8986 (N_8986,N_8603,N_8523);
and U8987 (N_8987,N_8504,N_8695);
xnor U8988 (N_8988,N_8509,N_8593);
xnor U8989 (N_8989,N_8629,N_8592);
xnor U8990 (N_8990,N_8690,N_8563);
xor U8991 (N_8991,N_8644,N_8635);
nor U8992 (N_8992,N_8589,N_8500);
nand U8993 (N_8993,N_8598,N_8590);
nor U8994 (N_8994,N_8625,N_8549);
or U8995 (N_8995,N_8642,N_8529);
xnor U8996 (N_8996,N_8733,N_8685);
nand U8997 (N_8997,N_8661,N_8595);
nand U8998 (N_8998,N_8687,N_8571);
nand U8999 (N_8999,N_8615,N_8681);
nor U9000 (N_9000,N_8943,N_8761);
xor U9001 (N_9001,N_8757,N_8929);
nor U9002 (N_9002,N_8884,N_8835);
xor U9003 (N_9003,N_8842,N_8856);
or U9004 (N_9004,N_8877,N_8866);
nand U9005 (N_9005,N_8807,N_8926);
nor U9006 (N_9006,N_8852,N_8887);
and U9007 (N_9007,N_8933,N_8939);
xnor U9008 (N_9008,N_8799,N_8966);
nor U9009 (N_9009,N_8876,N_8774);
nor U9010 (N_9010,N_8947,N_8973);
nor U9011 (N_9011,N_8821,N_8851);
nand U9012 (N_9012,N_8843,N_8989);
nand U9013 (N_9013,N_8932,N_8861);
nand U9014 (N_9014,N_8996,N_8840);
nor U9015 (N_9015,N_8896,N_8764);
xor U9016 (N_9016,N_8829,N_8894);
or U9017 (N_9017,N_8971,N_8809);
nand U9018 (N_9018,N_8936,N_8916);
and U9019 (N_9019,N_8953,N_8776);
xnor U9020 (N_9020,N_8862,N_8899);
nor U9021 (N_9021,N_8766,N_8830);
nand U9022 (N_9022,N_8880,N_8981);
and U9023 (N_9023,N_8778,N_8907);
and U9024 (N_9024,N_8962,N_8858);
or U9025 (N_9025,N_8920,N_8883);
nor U9026 (N_9026,N_8906,N_8972);
and U9027 (N_9027,N_8760,N_8976);
xor U9028 (N_9028,N_8863,N_8758);
nand U9029 (N_9029,N_8984,N_8847);
nand U9030 (N_9030,N_8754,N_8955);
nor U9031 (N_9031,N_8762,N_8811);
and U9032 (N_9032,N_8922,N_8796);
and U9033 (N_9033,N_8849,N_8923);
nand U9034 (N_9034,N_8779,N_8871);
and U9035 (N_9035,N_8781,N_8833);
nand U9036 (N_9036,N_8794,N_8759);
xor U9037 (N_9037,N_8820,N_8803);
nand U9038 (N_9038,N_8870,N_8927);
and U9039 (N_9039,N_8788,N_8879);
or U9040 (N_9040,N_8959,N_8804);
xor U9041 (N_9041,N_8853,N_8948);
or U9042 (N_9042,N_8928,N_8914);
or U9043 (N_9043,N_8956,N_8752);
nand U9044 (N_9044,N_8957,N_8991);
xnor U9045 (N_9045,N_8841,N_8898);
and U9046 (N_9046,N_8911,N_8944);
xnor U9047 (N_9047,N_8934,N_8812);
nor U9048 (N_9048,N_8867,N_8753);
nor U9049 (N_9049,N_8980,N_8949);
xor U9050 (N_9050,N_8931,N_8825);
nor U9051 (N_9051,N_8924,N_8831);
and U9052 (N_9052,N_8838,N_8945);
xnor U9053 (N_9053,N_8773,N_8782);
xnor U9054 (N_9054,N_8768,N_8897);
nand U9055 (N_9055,N_8937,N_8791);
or U9056 (N_9056,N_8913,N_8793);
and U9057 (N_9057,N_8816,N_8965);
and U9058 (N_9058,N_8941,N_8942);
and U9059 (N_9059,N_8848,N_8817);
and U9060 (N_9060,N_8969,N_8795);
nand U9061 (N_9061,N_8977,N_8946);
nand U9062 (N_9062,N_8872,N_8818);
and U9063 (N_9063,N_8868,N_8987);
nor U9064 (N_9064,N_8901,N_8893);
nand U9065 (N_9065,N_8772,N_8952);
and U9066 (N_9066,N_8822,N_8990);
xnor U9067 (N_9067,N_8988,N_8846);
nand U9068 (N_9068,N_8968,N_8792);
nor U9069 (N_9069,N_8921,N_8802);
nand U9070 (N_9070,N_8910,N_8892);
nand U9071 (N_9071,N_8967,N_8850);
or U9072 (N_9072,N_8881,N_8854);
or U9073 (N_9073,N_8763,N_8915);
xnor U9074 (N_9074,N_8983,N_8889);
and U9075 (N_9075,N_8951,N_8930);
xnor U9076 (N_9076,N_8978,N_8828);
or U9077 (N_9077,N_8909,N_8813);
nand U9078 (N_9078,N_8998,N_8823);
nor U9079 (N_9079,N_8860,N_8903);
and U9080 (N_9080,N_8827,N_8751);
and U9081 (N_9081,N_8912,N_8770);
and U9082 (N_9082,N_8891,N_8940);
xnor U9083 (N_9083,N_8785,N_8985);
or U9084 (N_9084,N_8886,N_8874);
and U9085 (N_9085,N_8771,N_8885);
or U9086 (N_9086,N_8982,N_8784);
and U9087 (N_9087,N_8800,N_8750);
xor U9088 (N_9088,N_8904,N_8780);
nand U9089 (N_9089,N_8900,N_8986);
or U9090 (N_9090,N_8805,N_8859);
or U9091 (N_9091,N_8918,N_8993);
nor U9092 (N_9092,N_8826,N_8875);
or U9093 (N_9093,N_8855,N_8975);
nand U9094 (N_9094,N_8890,N_8865);
or U9095 (N_9095,N_8790,N_8869);
nand U9096 (N_9096,N_8837,N_8919);
and U9097 (N_9097,N_8767,N_8864);
xor U9098 (N_9098,N_8834,N_8797);
xnor U9099 (N_9099,N_8765,N_8958);
xnor U9100 (N_9100,N_8756,N_8895);
xnor U9101 (N_9101,N_8992,N_8783);
or U9102 (N_9102,N_8777,N_8964);
xor U9103 (N_9103,N_8801,N_8938);
nor U9104 (N_9104,N_8974,N_8775);
nand U9105 (N_9105,N_8857,N_8836);
and U9106 (N_9106,N_8832,N_8917);
xnor U9107 (N_9107,N_8873,N_8960);
nand U9108 (N_9108,N_8970,N_8839);
nand U9109 (N_9109,N_8814,N_8824);
and U9110 (N_9110,N_8999,N_8888);
or U9111 (N_9111,N_8819,N_8815);
and U9112 (N_9112,N_8844,N_8979);
nand U9113 (N_9113,N_8954,N_8997);
nand U9114 (N_9114,N_8905,N_8769);
and U9115 (N_9115,N_8798,N_8908);
nand U9116 (N_9116,N_8935,N_8882);
xor U9117 (N_9117,N_8808,N_8950);
or U9118 (N_9118,N_8925,N_8755);
xnor U9119 (N_9119,N_8963,N_8806);
nand U9120 (N_9120,N_8878,N_8994);
nand U9121 (N_9121,N_8995,N_8902);
xor U9122 (N_9122,N_8961,N_8810);
xor U9123 (N_9123,N_8786,N_8787);
xor U9124 (N_9124,N_8845,N_8789);
or U9125 (N_9125,N_8820,N_8971);
nor U9126 (N_9126,N_8833,N_8827);
and U9127 (N_9127,N_8957,N_8847);
xor U9128 (N_9128,N_8778,N_8785);
nand U9129 (N_9129,N_8939,N_8844);
nand U9130 (N_9130,N_8770,N_8874);
or U9131 (N_9131,N_8825,N_8815);
or U9132 (N_9132,N_8886,N_8803);
nor U9133 (N_9133,N_8851,N_8799);
nor U9134 (N_9134,N_8863,N_8962);
xnor U9135 (N_9135,N_8986,N_8941);
and U9136 (N_9136,N_8929,N_8813);
or U9137 (N_9137,N_8891,N_8785);
nor U9138 (N_9138,N_8900,N_8854);
nand U9139 (N_9139,N_8903,N_8955);
nand U9140 (N_9140,N_8766,N_8842);
or U9141 (N_9141,N_8814,N_8976);
or U9142 (N_9142,N_8876,N_8892);
or U9143 (N_9143,N_8866,N_8807);
nor U9144 (N_9144,N_8936,N_8857);
or U9145 (N_9145,N_8753,N_8904);
nand U9146 (N_9146,N_8773,N_8841);
nor U9147 (N_9147,N_8889,N_8980);
nand U9148 (N_9148,N_8928,N_8750);
or U9149 (N_9149,N_8995,N_8857);
or U9150 (N_9150,N_8822,N_8942);
nor U9151 (N_9151,N_8931,N_8873);
nand U9152 (N_9152,N_8986,N_8859);
nand U9153 (N_9153,N_8998,N_8925);
xor U9154 (N_9154,N_8774,N_8888);
and U9155 (N_9155,N_8961,N_8898);
xor U9156 (N_9156,N_8842,N_8966);
xor U9157 (N_9157,N_8811,N_8998);
xnor U9158 (N_9158,N_8776,N_8988);
nor U9159 (N_9159,N_8882,N_8992);
or U9160 (N_9160,N_8924,N_8874);
or U9161 (N_9161,N_8985,N_8784);
xnor U9162 (N_9162,N_8813,N_8791);
nand U9163 (N_9163,N_8838,N_8970);
nor U9164 (N_9164,N_8946,N_8871);
xor U9165 (N_9165,N_8870,N_8881);
and U9166 (N_9166,N_8868,N_8791);
and U9167 (N_9167,N_8959,N_8854);
nor U9168 (N_9168,N_8828,N_8965);
xnor U9169 (N_9169,N_8929,N_8805);
and U9170 (N_9170,N_8754,N_8794);
or U9171 (N_9171,N_8996,N_8946);
nor U9172 (N_9172,N_8762,N_8806);
or U9173 (N_9173,N_8789,N_8993);
and U9174 (N_9174,N_8933,N_8916);
or U9175 (N_9175,N_8846,N_8831);
or U9176 (N_9176,N_8971,N_8817);
nor U9177 (N_9177,N_8818,N_8996);
and U9178 (N_9178,N_8756,N_8845);
nand U9179 (N_9179,N_8971,N_8950);
and U9180 (N_9180,N_8786,N_8874);
xnor U9181 (N_9181,N_8842,N_8825);
and U9182 (N_9182,N_8801,N_8862);
and U9183 (N_9183,N_8979,N_8810);
or U9184 (N_9184,N_8952,N_8846);
or U9185 (N_9185,N_8850,N_8857);
nand U9186 (N_9186,N_8965,N_8827);
and U9187 (N_9187,N_8902,N_8967);
and U9188 (N_9188,N_8792,N_8776);
nand U9189 (N_9189,N_8904,N_8993);
or U9190 (N_9190,N_8814,N_8863);
xnor U9191 (N_9191,N_8798,N_8906);
and U9192 (N_9192,N_8809,N_8886);
nand U9193 (N_9193,N_8941,N_8912);
nand U9194 (N_9194,N_8877,N_8922);
nor U9195 (N_9195,N_8889,N_8864);
or U9196 (N_9196,N_8781,N_8910);
xor U9197 (N_9197,N_8910,N_8996);
or U9198 (N_9198,N_8750,N_8984);
and U9199 (N_9199,N_8799,N_8931);
nor U9200 (N_9200,N_8761,N_8762);
nand U9201 (N_9201,N_8848,N_8900);
nor U9202 (N_9202,N_8792,N_8938);
nand U9203 (N_9203,N_8961,N_8813);
nor U9204 (N_9204,N_8843,N_8897);
xnor U9205 (N_9205,N_8825,N_8847);
nor U9206 (N_9206,N_8880,N_8958);
xor U9207 (N_9207,N_8788,N_8817);
xor U9208 (N_9208,N_8904,N_8859);
xnor U9209 (N_9209,N_8831,N_8856);
nor U9210 (N_9210,N_8910,N_8978);
or U9211 (N_9211,N_8853,N_8922);
or U9212 (N_9212,N_8801,N_8864);
nor U9213 (N_9213,N_8936,N_8940);
nor U9214 (N_9214,N_8776,N_8840);
nor U9215 (N_9215,N_8794,N_8851);
nand U9216 (N_9216,N_8875,N_8876);
nand U9217 (N_9217,N_8975,N_8769);
or U9218 (N_9218,N_8884,N_8845);
nor U9219 (N_9219,N_8760,N_8966);
or U9220 (N_9220,N_8778,N_8842);
or U9221 (N_9221,N_8879,N_8776);
xnor U9222 (N_9222,N_8853,N_8855);
nor U9223 (N_9223,N_8925,N_8863);
xor U9224 (N_9224,N_8783,N_8935);
nor U9225 (N_9225,N_8776,N_8823);
or U9226 (N_9226,N_8885,N_8968);
nand U9227 (N_9227,N_8892,N_8995);
nor U9228 (N_9228,N_8786,N_8938);
or U9229 (N_9229,N_8798,N_8933);
and U9230 (N_9230,N_8971,N_8822);
and U9231 (N_9231,N_8779,N_8920);
and U9232 (N_9232,N_8871,N_8851);
nand U9233 (N_9233,N_8791,N_8776);
or U9234 (N_9234,N_8798,N_8967);
nor U9235 (N_9235,N_8855,N_8984);
nand U9236 (N_9236,N_8884,N_8858);
nand U9237 (N_9237,N_8855,N_8969);
xor U9238 (N_9238,N_8900,N_8984);
nor U9239 (N_9239,N_8754,N_8775);
nand U9240 (N_9240,N_8781,N_8987);
nor U9241 (N_9241,N_8990,N_8869);
xor U9242 (N_9242,N_8893,N_8959);
xor U9243 (N_9243,N_8933,N_8856);
and U9244 (N_9244,N_8858,N_8909);
nor U9245 (N_9245,N_8973,N_8954);
xor U9246 (N_9246,N_8957,N_8761);
nor U9247 (N_9247,N_8785,N_8896);
and U9248 (N_9248,N_8830,N_8811);
and U9249 (N_9249,N_8861,N_8834);
or U9250 (N_9250,N_9030,N_9208);
or U9251 (N_9251,N_9157,N_9243);
nor U9252 (N_9252,N_9086,N_9131);
nand U9253 (N_9253,N_9223,N_9107);
xnor U9254 (N_9254,N_9117,N_9127);
and U9255 (N_9255,N_9144,N_9244);
nor U9256 (N_9256,N_9162,N_9077);
and U9257 (N_9257,N_9067,N_9133);
or U9258 (N_9258,N_9129,N_9089);
and U9259 (N_9259,N_9147,N_9036);
xnor U9260 (N_9260,N_9024,N_9109);
or U9261 (N_9261,N_9006,N_9193);
or U9262 (N_9262,N_9183,N_9059);
and U9263 (N_9263,N_9200,N_9022);
nand U9264 (N_9264,N_9111,N_9085);
or U9265 (N_9265,N_9199,N_9161);
xnor U9266 (N_9266,N_9222,N_9105);
nor U9267 (N_9267,N_9171,N_9217);
xnor U9268 (N_9268,N_9230,N_9078);
nand U9269 (N_9269,N_9040,N_9181);
nor U9270 (N_9270,N_9075,N_9150);
and U9271 (N_9271,N_9155,N_9239);
xnor U9272 (N_9272,N_9080,N_9095);
xor U9273 (N_9273,N_9233,N_9003);
xnor U9274 (N_9274,N_9084,N_9009);
or U9275 (N_9275,N_9151,N_9143);
xor U9276 (N_9276,N_9015,N_9098);
nand U9277 (N_9277,N_9055,N_9113);
or U9278 (N_9278,N_9179,N_9247);
xor U9279 (N_9279,N_9163,N_9033);
or U9280 (N_9280,N_9092,N_9178);
nand U9281 (N_9281,N_9156,N_9206);
nor U9282 (N_9282,N_9068,N_9031);
and U9283 (N_9283,N_9212,N_9007);
or U9284 (N_9284,N_9173,N_9096);
nand U9285 (N_9285,N_9081,N_9130);
or U9286 (N_9286,N_9210,N_9041);
nand U9287 (N_9287,N_9017,N_9184);
or U9288 (N_9288,N_9194,N_9083);
and U9289 (N_9289,N_9176,N_9014);
nand U9290 (N_9290,N_9240,N_9225);
xor U9291 (N_9291,N_9160,N_9189);
or U9292 (N_9292,N_9056,N_9191);
and U9293 (N_9293,N_9182,N_9100);
xnor U9294 (N_9294,N_9020,N_9216);
xor U9295 (N_9295,N_9069,N_9112);
nand U9296 (N_9296,N_9220,N_9044);
nand U9297 (N_9297,N_9049,N_9221);
xor U9298 (N_9298,N_9241,N_9146);
nor U9299 (N_9299,N_9246,N_9001);
or U9300 (N_9300,N_9185,N_9042);
and U9301 (N_9301,N_9238,N_9126);
xor U9302 (N_9302,N_9013,N_9242);
or U9303 (N_9303,N_9115,N_9101);
and U9304 (N_9304,N_9145,N_9187);
nor U9305 (N_9305,N_9180,N_9093);
xnor U9306 (N_9306,N_9087,N_9123);
xor U9307 (N_9307,N_9211,N_9153);
xor U9308 (N_9308,N_9065,N_9139);
xor U9309 (N_9309,N_9154,N_9201);
nand U9310 (N_9310,N_9032,N_9116);
nand U9311 (N_9311,N_9121,N_9004);
or U9312 (N_9312,N_9213,N_9076);
and U9313 (N_9313,N_9029,N_9026);
nand U9314 (N_9314,N_9064,N_9237);
or U9315 (N_9315,N_9063,N_9158);
xor U9316 (N_9316,N_9088,N_9197);
or U9317 (N_9317,N_9023,N_9052);
or U9318 (N_9318,N_9079,N_9008);
or U9319 (N_9319,N_9054,N_9224);
xor U9320 (N_9320,N_9227,N_9051);
or U9321 (N_9321,N_9012,N_9019);
and U9322 (N_9322,N_9128,N_9120);
nor U9323 (N_9323,N_9166,N_9053);
and U9324 (N_9324,N_9057,N_9122);
xor U9325 (N_9325,N_9164,N_9226);
nand U9326 (N_9326,N_9021,N_9207);
and U9327 (N_9327,N_9205,N_9025);
nor U9328 (N_9328,N_9090,N_9110);
nor U9329 (N_9329,N_9136,N_9050);
nor U9330 (N_9330,N_9167,N_9066);
nor U9331 (N_9331,N_9249,N_9231);
or U9332 (N_9332,N_9070,N_9074);
xnor U9333 (N_9333,N_9135,N_9060);
xor U9334 (N_9334,N_9152,N_9010);
and U9335 (N_9335,N_9132,N_9235);
or U9336 (N_9336,N_9005,N_9228);
xnor U9337 (N_9337,N_9138,N_9037);
nor U9338 (N_9338,N_9236,N_9097);
xnor U9339 (N_9339,N_9114,N_9035);
nor U9340 (N_9340,N_9104,N_9232);
nor U9341 (N_9341,N_9108,N_9141);
nor U9342 (N_9342,N_9245,N_9218);
or U9343 (N_9343,N_9028,N_9018);
or U9344 (N_9344,N_9140,N_9198);
nand U9345 (N_9345,N_9048,N_9124);
or U9346 (N_9346,N_9142,N_9177);
and U9347 (N_9347,N_9190,N_9102);
or U9348 (N_9348,N_9188,N_9172);
and U9349 (N_9349,N_9195,N_9094);
xnor U9350 (N_9350,N_9165,N_9073);
nor U9351 (N_9351,N_9168,N_9215);
or U9352 (N_9352,N_9192,N_9034);
or U9353 (N_9353,N_9134,N_9038);
xnor U9354 (N_9354,N_9118,N_9062);
xor U9355 (N_9355,N_9082,N_9248);
or U9356 (N_9356,N_9027,N_9186);
and U9357 (N_9357,N_9203,N_9169);
nor U9358 (N_9358,N_9175,N_9209);
xor U9359 (N_9359,N_9047,N_9000);
nor U9360 (N_9360,N_9043,N_9148);
nand U9361 (N_9361,N_9099,N_9071);
nand U9362 (N_9362,N_9174,N_9196);
and U9363 (N_9363,N_9072,N_9125);
nor U9364 (N_9364,N_9002,N_9011);
xor U9365 (N_9365,N_9229,N_9106);
xor U9366 (N_9366,N_9119,N_9214);
xnor U9367 (N_9367,N_9234,N_9159);
nor U9368 (N_9368,N_9046,N_9045);
nand U9369 (N_9369,N_9149,N_9058);
nand U9370 (N_9370,N_9202,N_9016);
nand U9371 (N_9371,N_9137,N_9170);
xor U9372 (N_9372,N_9219,N_9204);
nand U9373 (N_9373,N_9091,N_9061);
xnor U9374 (N_9374,N_9039,N_9103);
nor U9375 (N_9375,N_9212,N_9023);
and U9376 (N_9376,N_9244,N_9104);
nor U9377 (N_9377,N_9060,N_9038);
and U9378 (N_9378,N_9138,N_9173);
xnor U9379 (N_9379,N_9120,N_9213);
nor U9380 (N_9380,N_9172,N_9142);
xor U9381 (N_9381,N_9184,N_9119);
and U9382 (N_9382,N_9192,N_9068);
nand U9383 (N_9383,N_9230,N_9035);
or U9384 (N_9384,N_9146,N_9089);
nor U9385 (N_9385,N_9114,N_9136);
xnor U9386 (N_9386,N_9145,N_9131);
and U9387 (N_9387,N_9199,N_9244);
and U9388 (N_9388,N_9065,N_9134);
nor U9389 (N_9389,N_9007,N_9176);
or U9390 (N_9390,N_9114,N_9041);
or U9391 (N_9391,N_9136,N_9139);
or U9392 (N_9392,N_9215,N_9142);
xor U9393 (N_9393,N_9178,N_9091);
nand U9394 (N_9394,N_9011,N_9140);
xnor U9395 (N_9395,N_9134,N_9007);
nand U9396 (N_9396,N_9208,N_9171);
or U9397 (N_9397,N_9064,N_9199);
and U9398 (N_9398,N_9135,N_9132);
xor U9399 (N_9399,N_9141,N_9146);
nand U9400 (N_9400,N_9000,N_9095);
nand U9401 (N_9401,N_9210,N_9099);
nand U9402 (N_9402,N_9060,N_9052);
and U9403 (N_9403,N_9012,N_9174);
and U9404 (N_9404,N_9120,N_9090);
nor U9405 (N_9405,N_9114,N_9202);
nor U9406 (N_9406,N_9195,N_9118);
nor U9407 (N_9407,N_9126,N_9122);
nor U9408 (N_9408,N_9116,N_9120);
and U9409 (N_9409,N_9121,N_9235);
nor U9410 (N_9410,N_9157,N_9038);
or U9411 (N_9411,N_9204,N_9140);
nand U9412 (N_9412,N_9043,N_9125);
or U9413 (N_9413,N_9062,N_9144);
or U9414 (N_9414,N_9246,N_9025);
xnor U9415 (N_9415,N_9101,N_9111);
or U9416 (N_9416,N_9018,N_9201);
or U9417 (N_9417,N_9076,N_9063);
xnor U9418 (N_9418,N_9219,N_9139);
or U9419 (N_9419,N_9074,N_9239);
nand U9420 (N_9420,N_9163,N_9242);
and U9421 (N_9421,N_9107,N_9073);
or U9422 (N_9422,N_9065,N_9026);
xnor U9423 (N_9423,N_9002,N_9010);
or U9424 (N_9424,N_9101,N_9061);
xnor U9425 (N_9425,N_9133,N_9194);
nand U9426 (N_9426,N_9152,N_9094);
xnor U9427 (N_9427,N_9225,N_9193);
xor U9428 (N_9428,N_9029,N_9056);
nand U9429 (N_9429,N_9195,N_9072);
nand U9430 (N_9430,N_9062,N_9210);
nor U9431 (N_9431,N_9049,N_9147);
and U9432 (N_9432,N_9078,N_9054);
nand U9433 (N_9433,N_9014,N_9108);
nand U9434 (N_9434,N_9032,N_9205);
nand U9435 (N_9435,N_9198,N_9076);
nand U9436 (N_9436,N_9075,N_9151);
nor U9437 (N_9437,N_9064,N_9004);
xnor U9438 (N_9438,N_9209,N_9204);
nor U9439 (N_9439,N_9047,N_9243);
nor U9440 (N_9440,N_9090,N_9228);
xor U9441 (N_9441,N_9078,N_9169);
xor U9442 (N_9442,N_9028,N_9234);
or U9443 (N_9443,N_9093,N_9221);
or U9444 (N_9444,N_9211,N_9125);
xnor U9445 (N_9445,N_9013,N_9195);
xnor U9446 (N_9446,N_9146,N_9081);
xnor U9447 (N_9447,N_9130,N_9105);
xor U9448 (N_9448,N_9201,N_9028);
and U9449 (N_9449,N_9105,N_9114);
nor U9450 (N_9450,N_9051,N_9243);
or U9451 (N_9451,N_9119,N_9211);
xor U9452 (N_9452,N_9155,N_9227);
and U9453 (N_9453,N_9008,N_9119);
or U9454 (N_9454,N_9054,N_9036);
xnor U9455 (N_9455,N_9155,N_9240);
nor U9456 (N_9456,N_9058,N_9102);
xor U9457 (N_9457,N_9216,N_9231);
and U9458 (N_9458,N_9044,N_9148);
nor U9459 (N_9459,N_9055,N_9119);
nor U9460 (N_9460,N_9150,N_9192);
nand U9461 (N_9461,N_9105,N_9091);
xor U9462 (N_9462,N_9017,N_9083);
nand U9463 (N_9463,N_9038,N_9145);
nand U9464 (N_9464,N_9185,N_9038);
nand U9465 (N_9465,N_9204,N_9154);
xor U9466 (N_9466,N_9129,N_9228);
nand U9467 (N_9467,N_9077,N_9033);
and U9468 (N_9468,N_9249,N_9107);
or U9469 (N_9469,N_9019,N_9194);
nand U9470 (N_9470,N_9207,N_9076);
nor U9471 (N_9471,N_9166,N_9112);
xor U9472 (N_9472,N_9110,N_9146);
xor U9473 (N_9473,N_9180,N_9193);
and U9474 (N_9474,N_9155,N_9055);
nand U9475 (N_9475,N_9139,N_9094);
nor U9476 (N_9476,N_9174,N_9130);
xor U9477 (N_9477,N_9135,N_9179);
or U9478 (N_9478,N_9078,N_9235);
nand U9479 (N_9479,N_9208,N_9056);
or U9480 (N_9480,N_9017,N_9132);
nand U9481 (N_9481,N_9149,N_9209);
and U9482 (N_9482,N_9157,N_9179);
nand U9483 (N_9483,N_9042,N_9066);
or U9484 (N_9484,N_9052,N_9236);
nor U9485 (N_9485,N_9173,N_9232);
or U9486 (N_9486,N_9059,N_9057);
and U9487 (N_9487,N_9247,N_9014);
nand U9488 (N_9488,N_9022,N_9174);
and U9489 (N_9489,N_9142,N_9171);
xor U9490 (N_9490,N_9077,N_9236);
and U9491 (N_9491,N_9164,N_9139);
nor U9492 (N_9492,N_9110,N_9046);
and U9493 (N_9493,N_9174,N_9024);
xor U9494 (N_9494,N_9080,N_9058);
and U9495 (N_9495,N_9158,N_9217);
xnor U9496 (N_9496,N_9026,N_9206);
xor U9497 (N_9497,N_9125,N_9228);
nand U9498 (N_9498,N_9008,N_9156);
or U9499 (N_9499,N_9230,N_9179);
xnor U9500 (N_9500,N_9318,N_9290);
or U9501 (N_9501,N_9310,N_9431);
xnor U9502 (N_9502,N_9333,N_9287);
nor U9503 (N_9503,N_9373,N_9281);
nand U9504 (N_9504,N_9383,N_9384);
or U9505 (N_9505,N_9399,N_9276);
nor U9506 (N_9506,N_9482,N_9327);
nand U9507 (N_9507,N_9291,N_9320);
or U9508 (N_9508,N_9269,N_9491);
and U9509 (N_9509,N_9423,N_9270);
xor U9510 (N_9510,N_9346,N_9317);
nand U9511 (N_9511,N_9430,N_9350);
and U9512 (N_9512,N_9449,N_9378);
or U9513 (N_9513,N_9274,N_9465);
xor U9514 (N_9514,N_9481,N_9324);
nand U9515 (N_9515,N_9377,N_9397);
or U9516 (N_9516,N_9389,N_9447);
nor U9517 (N_9517,N_9288,N_9370);
or U9518 (N_9518,N_9425,N_9341);
and U9519 (N_9519,N_9296,N_9480);
and U9520 (N_9520,N_9354,N_9405);
nand U9521 (N_9521,N_9454,N_9263);
nand U9522 (N_9522,N_9474,N_9371);
nor U9523 (N_9523,N_9294,N_9466);
nand U9524 (N_9524,N_9305,N_9437);
nand U9525 (N_9525,N_9266,N_9435);
xnor U9526 (N_9526,N_9470,N_9469);
or U9527 (N_9527,N_9395,N_9368);
or U9528 (N_9528,N_9391,N_9301);
xor U9529 (N_9529,N_9388,N_9485);
or U9530 (N_9530,N_9467,N_9306);
nor U9531 (N_9531,N_9277,N_9256);
or U9532 (N_9532,N_9259,N_9250);
nand U9533 (N_9533,N_9451,N_9366);
and U9534 (N_9534,N_9392,N_9353);
nor U9535 (N_9535,N_9311,N_9359);
nand U9536 (N_9536,N_9462,N_9261);
or U9537 (N_9537,N_9351,N_9442);
xor U9538 (N_9538,N_9369,N_9381);
nand U9539 (N_9539,N_9441,N_9468);
xor U9540 (N_9540,N_9387,N_9448);
nor U9541 (N_9541,N_9475,N_9326);
or U9542 (N_9542,N_9495,N_9477);
or U9543 (N_9543,N_9415,N_9499);
xor U9544 (N_9544,N_9494,N_9459);
nand U9545 (N_9545,N_9408,N_9367);
or U9546 (N_9546,N_9283,N_9444);
and U9547 (N_9547,N_9410,N_9409);
and U9548 (N_9548,N_9406,N_9349);
nor U9549 (N_9549,N_9260,N_9411);
nand U9550 (N_9550,N_9362,N_9376);
nor U9551 (N_9551,N_9461,N_9292);
and U9552 (N_9552,N_9315,N_9487);
or U9553 (N_9553,N_9360,N_9489);
nor U9554 (N_9554,N_9355,N_9471);
xor U9555 (N_9555,N_9286,N_9404);
nor U9556 (N_9556,N_9476,N_9329);
and U9557 (N_9557,N_9325,N_9330);
or U9558 (N_9558,N_9450,N_9338);
nor U9559 (N_9559,N_9356,N_9314);
or U9560 (N_9560,N_9284,N_9342);
and U9561 (N_9561,N_9251,N_9420);
nor U9562 (N_9562,N_9297,N_9374);
nor U9563 (N_9563,N_9335,N_9394);
xor U9564 (N_9564,N_9272,N_9257);
xnor U9565 (N_9565,N_9344,N_9337);
or U9566 (N_9566,N_9278,N_9303);
nand U9567 (N_9567,N_9414,N_9336);
or U9568 (N_9568,N_9357,N_9304);
nor U9569 (N_9569,N_9427,N_9426);
nand U9570 (N_9570,N_9352,N_9340);
and U9571 (N_9571,N_9438,N_9280);
or U9572 (N_9572,N_9400,N_9460);
nor U9573 (N_9573,N_9416,N_9348);
or U9574 (N_9574,N_9456,N_9363);
xnor U9575 (N_9575,N_9419,N_9273);
nand U9576 (N_9576,N_9453,N_9434);
nand U9577 (N_9577,N_9464,N_9380);
nor U9578 (N_9578,N_9253,N_9439);
or U9579 (N_9579,N_9428,N_9275);
nor U9580 (N_9580,N_9396,N_9421);
or U9581 (N_9581,N_9417,N_9254);
xnor U9582 (N_9582,N_9331,N_9322);
and U9583 (N_9583,N_9379,N_9401);
xor U9584 (N_9584,N_9312,N_9293);
and U9585 (N_9585,N_9497,N_9299);
xor U9586 (N_9586,N_9265,N_9473);
xnor U9587 (N_9587,N_9267,N_9484);
nand U9588 (N_9588,N_9262,N_9343);
or U9589 (N_9589,N_9295,N_9289);
nand U9590 (N_9590,N_9279,N_9339);
nor U9591 (N_9591,N_9308,N_9334);
or U9592 (N_9592,N_9316,N_9486);
nor U9593 (N_9593,N_9463,N_9358);
nor U9594 (N_9594,N_9398,N_9422);
xnor U9595 (N_9595,N_9255,N_9307);
nand U9596 (N_9596,N_9418,N_9424);
and U9597 (N_9597,N_9385,N_9492);
xnor U9598 (N_9598,N_9490,N_9302);
xor U9599 (N_9599,N_9319,N_9403);
nand U9600 (N_9600,N_9372,N_9432);
nor U9601 (N_9601,N_9361,N_9298);
nand U9602 (N_9602,N_9382,N_9323);
and U9603 (N_9603,N_9445,N_9429);
or U9604 (N_9604,N_9282,N_9375);
nand U9605 (N_9605,N_9455,N_9321);
and U9606 (N_9606,N_9271,N_9402);
and U9607 (N_9607,N_9443,N_9390);
nand U9608 (N_9608,N_9436,N_9258);
or U9609 (N_9609,N_9364,N_9413);
nand U9610 (N_9610,N_9300,N_9393);
xor U9611 (N_9611,N_9483,N_9252);
nor U9612 (N_9612,N_9478,N_9386);
and U9613 (N_9613,N_9264,N_9496);
xnor U9614 (N_9614,N_9440,N_9328);
xor U9615 (N_9615,N_9452,N_9365);
and U9616 (N_9616,N_9347,N_9412);
nor U9617 (N_9617,N_9309,N_9268);
nand U9618 (N_9618,N_9433,N_9458);
or U9619 (N_9619,N_9285,N_9313);
or U9620 (N_9620,N_9407,N_9446);
xnor U9621 (N_9621,N_9479,N_9345);
and U9622 (N_9622,N_9457,N_9332);
xnor U9623 (N_9623,N_9488,N_9493);
nor U9624 (N_9624,N_9472,N_9498);
and U9625 (N_9625,N_9370,N_9389);
xnor U9626 (N_9626,N_9301,N_9453);
and U9627 (N_9627,N_9441,N_9266);
nor U9628 (N_9628,N_9284,N_9426);
or U9629 (N_9629,N_9486,N_9423);
xor U9630 (N_9630,N_9324,N_9417);
and U9631 (N_9631,N_9332,N_9251);
nor U9632 (N_9632,N_9465,N_9300);
nor U9633 (N_9633,N_9307,N_9435);
or U9634 (N_9634,N_9261,N_9315);
nor U9635 (N_9635,N_9491,N_9378);
xor U9636 (N_9636,N_9305,N_9496);
nor U9637 (N_9637,N_9285,N_9346);
or U9638 (N_9638,N_9341,N_9354);
and U9639 (N_9639,N_9318,N_9337);
or U9640 (N_9640,N_9315,N_9422);
and U9641 (N_9641,N_9420,N_9399);
xnor U9642 (N_9642,N_9331,N_9467);
xnor U9643 (N_9643,N_9298,N_9483);
xnor U9644 (N_9644,N_9251,N_9399);
nor U9645 (N_9645,N_9405,N_9340);
or U9646 (N_9646,N_9454,N_9443);
xor U9647 (N_9647,N_9408,N_9435);
nor U9648 (N_9648,N_9357,N_9256);
nor U9649 (N_9649,N_9277,N_9284);
and U9650 (N_9650,N_9364,N_9457);
nor U9651 (N_9651,N_9251,N_9263);
nor U9652 (N_9652,N_9353,N_9283);
nor U9653 (N_9653,N_9312,N_9445);
or U9654 (N_9654,N_9470,N_9404);
and U9655 (N_9655,N_9494,N_9404);
nor U9656 (N_9656,N_9284,N_9298);
or U9657 (N_9657,N_9443,N_9299);
nor U9658 (N_9658,N_9386,N_9256);
nand U9659 (N_9659,N_9394,N_9321);
or U9660 (N_9660,N_9412,N_9296);
nor U9661 (N_9661,N_9316,N_9382);
nand U9662 (N_9662,N_9486,N_9256);
xor U9663 (N_9663,N_9419,N_9413);
xnor U9664 (N_9664,N_9374,N_9325);
nor U9665 (N_9665,N_9441,N_9398);
nor U9666 (N_9666,N_9264,N_9431);
nor U9667 (N_9667,N_9289,N_9335);
and U9668 (N_9668,N_9461,N_9421);
nor U9669 (N_9669,N_9399,N_9441);
xor U9670 (N_9670,N_9344,N_9291);
nand U9671 (N_9671,N_9366,N_9388);
nand U9672 (N_9672,N_9381,N_9422);
nand U9673 (N_9673,N_9288,N_9331);
nor U9674 (N_9674,N_9264,N_9406);
xor U9675 (N_9675,N_9445,N_9355);
or U9676 (N_9676,N_9298,N_9335);
and U9677 (N_9677,N_9443,N_9333);
xnor U9678 (N_9678,N_9460,N_9490);
nand U9679 (N_9679,N_9256,N_9388);
xor U9680 (N_9680,N_9483,N_9280);
and U9681 (N_9681,N_9259,N_9486);
xnor U9682 (N_9682,N_9404,N_9455);
and U9683 (N_9683,N_9489,N_9449);
nor U9684 (N_9684,N_9275,N_9414);
or U9685 (N_9685,N_9433,N_9492);
xnor U9686 (N_9686,N_9457,N_9355);
or U9687 (N_9687,N_9287,N_9448);
and U9688 (N_9688,N_9461,N_9449);
or U9689 (N_9689,N_9289,N_9427);
or U9690 (N_9690,N_9443,N_9267);
or U9691 (N_9691,N_9305,N_9435);
nor U9692 (N_9692,N_9272,N_9490);
or U9693 (N_9693,N_9473,N_9465);
nor U9694 (N_9694,N_9332,N_9484);
xor U9695 (N_9695,N_9340,N_9323);
nor U9696 (N_9696,N_9467,N_9436);
xnor U9697 (N_9697,N_9273,N_9329);
nand U9698 (N_9698,N_9310,N_9432);
nand U9699 (N_9699,N_9432,N_9257);
or U9700 (N_9700,N_9463,N_9285);
and U9701 (N_9701,N_9253,N_9343);
xnor U9702 (N_9702,N_9295,N_9422);
and U9703 (N_9703,N_9384,N_9487);
and U9704 (N_9704,N_9423,N_9275);
and U9705 (N_9705,N_9267,N_9269);
and U9706 (N_9706,N_9275,N_9348);
and U9707 (N_9707,N_9409,N_9419);
or U9708 (N_9708,N_9406,N_9391);
or U9709 (N_9709,N_9368,N_9388);
or U9710 (N_9710,N_9380,N_9402);
nor U9711 (N_9711,N_9331,N_9419);
and U9712 (N_9712,N_9416,N_9352);
nor U9713 (N_9713,N_9427,N_9264);
xor U9714 (N_9714,N_9317,N_9377);
or U9715 (N_9715,N_9348,N_9458);
xor U9716 (N_9716,N_9296,N_9299);
xor U9717 (N_9717,N_9273,N_9381);
xnor U9718 (N_9718,N_9294,N_9255);
or U9719 (N_9719,N_9336,N_9476);
nand U9720 (N_9720,N_9250,N_9437);
xnor U9721 (N_9721,N_9417,N_9400);
and U9722 (N_9722,N_9282,N_9409);
nor U9723 (N_9723,N_9251,N_9326);
nor U9724 (N_9724,N_9380,N_9447);
and U9725 (N_9725,N_9432,N_9408);
nand U9726 (N_9726,N_9254,N_9479);
and U9727 (N_9727,N_9495,N_9304);
and U9728 (N_9728,N_9370,N_9441);
xnor U9729 (N_9729,N_9483,N_9372);
or U9730 (N_9730,N_9357,N_9467);
and U9731 (N_9731,N_9300,N_9450);
and U9732 (N_9732,N_9433,N_9491);
xnor U9733 (N_9733,N_9480,N_9342);
xor U9734 (N_9734,N_9479,N_9336);
and U9735 (N_9735,N_9269,N_9371);
nor U9736 (N_9736,N_9273,N_9494);
nand U9737 (N_9737,N_9267,N_9356);
nor U9738 (N_9738,N_9437,N_9348);
xor U9739 (N_9739,N_9495,N_9415);
and U9740 (N_9740,N_9475,N_9456);
nand U9741 (N_9741,N_9440,N_9475);
xnor U9742 (N_9742,N_9304,N_9307);
nor U9743 (N_9743,N_9400,N_9255);
xnor U9744 (N_9744,N_9366,N_9273);
nand U9745 (N_9745,N_9454,N_9270);
xnor U9746 (N_9746,N_9294,N_9400);
nand U9747 (N_9747,N_9262,N_9363);
nor U9748 (N_9748,N_9316,N_9469);
nor U9749 (N_9749,N_9301,N_9288);
xor U9750 (N_9750,N_9549,N_9602);
or U9751 (N_9751,N_9717,N_9741);
xor U9752 (N_9752,N_9556,N_9583);
nor U9753 (N_9753,N_9662,N_9560);
xor U9754 (N_9754,N_9572,N_9707);
or U9755 (N_9755,N_9704,N_9621);
or U9756 (N_9756,N_9608,N_9604);
and U9757 (N_9757,N_9618,N_9656);
and U9758 (N_9758,N_9641,N_9558);
nor U9759 (N_9759,N_9748,N_9696);
or U9760 (N_9760,N_9702,N_9647);
or U9761 (N_9761,N_9642,N_9567);
xor U9762 (N_9762,N_9650,N_9694);
nor U9763 (N_9763,N_9512,N_9588);
and U9764 (N_9764,N_9659,N_9526);
nand U9765 (N_9765,N_9522,N_9534);
nor U9766 (N_9766,N_9569,N_9657);
xnor U9767 (N_9767,N_9668,N_9601);
nor U9768 (N_9768,N_9630,N_9614);
or U9769 (N_9769,N_9518,N_9557);
xnor U9770 (N_9770,N_9686,N_9563);
nand U9771 (N_9771,N_9735,N_9637);
xor U9772 (N_9772,N_9672,N_9680);
xnor U9773 (N_9773,N_9509,N_9628);
or U9774 (N_9774,N_9718,N_9689);
and U9775 (N_9775,N_9503,N_9548);
nor U9776 (N_9776,N_9624,N_9597);
and U9777 (N_9777,N_9559,N_9594);
and U9778 (N_9778,N_9673,N_9681);
nor U9779 (N_9779,N_9653,N_9623);
xnor U9780 (N_9780,N_9543,N_9660);
xnor U9781 (N_9781,N_9606,N_9613);
and U9782 (N_9782,N_9734,N_9574);
nor U9783 (N_9783,N_9540,N_9609);
nand U9784 (N_9784,N_9538,N_9579);
nand U9785 (N_9785,N_9706,N_9690);
nand U9786 (N_9786,N_9622,N_9733);
or U9787 (N_9787,N_9721,N_9545);
and U9788 (N_9788,N_9573,N_9697);
nand U9789 (N_9789,N_9737,N_9670);
or U9790 (N_9790,N_9646,N_9555);
nand U9791 (N_9791,N_9727,N_9716);
nor U9792 (N_9792,N_9577,N_9546);
nor U9793 (N_9793,N_9654,N_9644);
and U9794 (N_9794,N_9500,N_9698);
nand U9795 (N_9795,N_9519,N_9695);
nor U9796 (N_9796,N_9677,N_9714);
nand U9797 (N_9797,N_9539,N_9591);
nor U9798 (N_9798,N_9515,N_9638);
nor U9799 (N_9799,N_9523,N_9732);
xnor U9800 (N_9800,N_9554,N_9729);
and U9801 (N_9801,N_9575,N_9631);
nand U9802 (N_9802,N_9535,N_9612);
nor U9803 (N_9803,N_9617,N_9730);
or U9804 (N_9804,N_9626,N_9521);
xnor U9805 (N_9805,N_9731,N_9705);
nand U9806 (N_9806,N_9517,N_9634);
nor U9807 (N_9807,N_9562,N_9611);
or U9808 (N_9808,N_9683,N_9699);
nand U9809 (N_9809,N_9635,N_9658);
xnor U9810 (N_9810,N_9675,N_9599);
and U9811 (N_9811,N_9568,N_9736);
or U9812 (N_9812,N_9506,N_9629);
nand U9813 (N_9813,N_9537,N_9516);
or U9814 (N_9814,N_9655,N_9640);
nand U9815 (N_9815,N_9615,N_9708);
nand U9816 (N_9816,N_9723,N_9595);
or U9817 (N_9817,N_9596,N_9649);
nor U9818 (N_9818,N_9715,N_9528);
nand U9819 (N_9819,N_9620,N_9520);
nor U9820 (N_9820,N_9607,N_9603);
nor U9821 (N_9821,N_9711,N_9643);
or U9822 (N_9822,N_9710,N_9645);
nor U9823 (N_9823,N_9738,N_9712);
or U9824 (N_9824,N_9542,N_9527);
nand U9825 (N_9825,N_9501,N_9532);
or U9826 (N_9826,N_9525,N_9692);
and U9827 (N_9827,N_9616,N_9605);
and U9828 (N_9828,N_9553,N_9669);
nand U9829 (N_9829,N_9740,N_9584);
nand U9830 (N_9830,N_9744,N_9693);
or U9831 (N_9831,N_9587,N_9508);
or U9832 (N_9832,N_9747,N_9749);
and U9833 (N_9833,N_9578,N_9739);
nand U9834 (N_9834,N_9514,N_9565);
nor U9835 (N_9835,N_9724,N_9592);
nand U9836 (N_9836,N_9585,N_9665);
or U9837 (N_9837,N_9671,N_9722);
nand U9838 (N_9838,N_9719,N_9726);
or U9839 (N_9839,N_9651,N_9700);
xor U9840 (N_9840,N_9510,N_9627);
and U9841 (N_9841,N_9610,N_9652);
and U9842 (N_9842,N_9505,N_9561);
or U9843 (N_9843,N_9502,N_9511);
xor U9844 (N_9844,N_9709,N_9600);
nor U9845 (N_9845,N_9582,N_9661);
and U9846 (N_9846,N_9691,N_9728);
nand U9847 (N_9847,N_9685,N_9536);
xnor U9848 (N_9848,N_9552,N_9566);
xor U9849 (N_9849,N_9678,N_9586);
nor U9850 (N_9850,N_9720,N_9581);
xor U9851 (N_9851,N_9674,N_9570);
or U9852 (N_9852,N_9551,N_9632);
nand U9853 (N_9853,N_9713,N_9663);
and U9854 (N_9854,N_9701,N_9667);
xnor U9855 (N_9855,N_9666,N_9745);
nor U9856 (N_9856,N_9746,N_9625);
nor U9857 (N_9857,N_9580,N_9513);
nand U9858 (N_9858,N_9639,N_9619);
nand U9859 (N_9859,N_9593,N_9633);
nor U9860 (N_9860,N_9725,N_9598);
nor U9861 (N_9861,N_9504,N_9571);
xor U9862 (N_9862,N_9531,N_9544);
nand U9863 (N_9863,N_9590,N_9529);
nand U9864 (N_9864,N_9648,N_9576);
nand U9865 (N_9865,N_9530,N_9507);
nor U9866 (N_9866,N_9742,N_9687);
nor U9867 (N_9867,N_9564,N_9533);
nand U9868 (N_9868,N_9589,N_9524);
nand U9869 (N_9869,N_9636,N_9541);
nand U9870 (N_9870,N_9664,N_9676);
and U9871 (N_9871,N_9547,N_9743);
nand U9872 (N_9872,N_9688,N_9682);
or U9873 (N_9873,N_9703,N_9550);
nand U9874 (N_9874,N_9684,N_9679);
or U9875 (N_9875,N_9655,N_9742);
nor U9876 (N_9876,N_9734,N_9520);
and U9877 (N_9877,N_9653,N_9519);
and U9878 (N_9878,N_9580,N_9601);
or U9879 (N_9879,N_9619,N_9713);
xor U9880 (N_9880,N_9521,N_9693);
or U9881 (N_9881,N_9587,N_9736);
or U9882 (N_9882,N_9595,N_9627);
and U9883 (N_9883,N_9500,N_9679);
nor U9884 (N_9884,N_9724,N_9561);
nor U9885 (N_9885,N_9705,N_9646);
nor U9886 (N_9886,N_9611,N_9721);
xnor U9887 (N_9887,N_9653,N_9521);
or U9888 (N_9888,N_9643,N_9513);
nand U9889 (N_9889,N_9739,N_9695);
and U9890 (N_9890,N_9730,N_9618);
nand U9891 (N_9891,N_9696,N_9554);
and U9892 (N_9892,N_9534,N_9661);
xnor U9893 (N_9893,N_9608,N_9621);
xnor U9894 (N_9894,N_9684,N_9553);
or U9895 (N_9895,N_9624,N_9748);
nor U9896 (N_9896,N_9655,N_9569);
nand U9897 (N_9897,N_9733,N_9627);
nand U9898 (N_9898,N_9638,N_9649);
xnor U9899 (N_9899,N_9745,N_9646);
nand U9900 (N_9900,N_9698,N_9704);
nand U9901 (N_9901,N_9542,N_9618);
and U9902 (N_9902,N_9518,N_9520);
or U9903 (N_9903,N_9673,N_9652);
and U9904 (N_9904,N_9684,N_9700);
nand U9905 (N_9905,N_9557,N_9511);
or U9906 (N_9906,N_9537,N_9745);
nand U9907 (N_9907,N_9557,N_9534);
and U9908 (N_9908,N_9549,N_9645);
and U9909 (N_9909,N_9684,N_9749);
nor U9910 (N_9910,N_9577,N_9571);
nor U9911 (N_9911,N_9726,N_9621);
nor U9912 (N_9912,N_9696,N_9611);
nor U9913 (N_9913,N_9665,N_9618);
or U9914 (N_9914,N_9506,N_9691);
and U9915 (N_9915,N_9748,N_9529);
and U9916 (N_9916,N_9591,N_9558);
or U9917 (N_9917,N_9591,N_9513);
or U9918 (N_9918,N_9613,N_9519);
or U9919 (N_9919,N_9551,N_9510);
and U9920 (N_9920,N_9703,N_9674);
xor U9921 (N_9921,N_9591,N_9749);
nand U9922 (N_9922,N_9717,N_9567);
nor U9923 (N_9923,N_9622,N_9722);
nand U9924 (N_9924,N_9669,N_9718);
nor U9925 (N_9925,N_9702,N_9686);
nand U9926 (N_9926,N_9568,N_9544);
or U9927 (N_9927,N_9588,N_9591);
xnor U9928 (N_9928,N_9641,N_9533);
nand U9929 (N_9929,N_9550,N_9549);
nor U9930 (N_9930,N_9577,N_9619);
and U9931 (N_9931,N_9560,N_9627);
nand U9932 (N_9932,N_9687,N_9661);
nand U9933 (N_9933,N_9540,N_9565);
nand U9934 (N_9934,N_9646,N_9700);
or U9935 (N_9935,N_9637,N_9586);
and U9936 (N_9936,N_9640,N_9734);
and U9937 (N_9937,N_9648,N_9536);
nor U9938 (N_9938,N_9707,N_9501);
nor U9939 (N_9939,N_9630,N_9514);
xor U9940 (N_9940,N_9649,N_9530);
nand U9941 (N_9941,N_9603,N_9538);
nand U9942 (N_9942,N_9618,N_9505);
nor U9943 (N_9943,N_9683,N_9541);
and U9944 (N_9944,N_9666,N_9660);
nor U9945 (N_9945,N_9502,N_9652);
and U9946 (N_9946,N_9685,N_9593);
nor U9947 (N_9947,N_9670,N_9538);
xor U9948 (N_9948,N_9643,N_9695);
xnor U9949 (N_9949,N_9573,N_9522);
nand U9950 (N_9950,N_9688,N_9706);
nand U9951 (N_9951,N_9519,N_9578);
nand U9952 (N_9952,N_9563,N_9559);
nand U9953 (N_9953,N_9737,N_9680);
xor U9954 (N_9954,N_9560,N_9666);
nor U9955 (N_9955,N_9671,N_9512);
or U9956 (N_9956,N_9536,N_9680);
xor U9957 (N_9957,N_9692,N_9682);
nor U9958 (N_9958,N_9519,N_9545);
nor U9959 (N_9959,N_9641,N_9704);
or U9960 (N_9960,N_9705,N_9522);
nor U9961 (N_9961,N_9624,N_9721);
nor U9962 (N_9962,N_9744,N_9553);
and U9963 (N_9963,N_9627,N_9619);
nor U9964 (N_9964,N_9651,N_9608);
xor U9965 (N_9965,N_9649,N_9503);
nand U9966 (N_9966,N_9568,N_9533);
nand U9967 (N_9967,N_9619,N_9720);
and U9968 (N_9968,N_9663,N_9636);
xor U9969 (N_9969,N_9543,N_9506);
nor U9970 (N_9970,N_9573,N_9597);
or U9971 (N_9971,N_9684,N_9734);
and U9972 (N_9972,N_9599,N_9571);
xor U9973 (N_9973,N_9631,N_9589);
or U9974 (N_9974,N_9543,N_9712);
and U9975 (N_9975,N_9551,N_9515);
and U9976 (N_9976,N_9577,N_9668);
or U9977 (N_9977,N_9688,N_9552);
nand U9978 (N_9978,N_9648,N_9746);
and U9979 (N_9979,N_9567,N_9617);
and U9980 (N_9980,N_9502,N_9670);
nand U9981 (N_9981,N_9599,N_9602);
and U9982 (N_9982,N_9637,N_9595);
nor U9983 (N_9983,N_9664,N_9712);
nand U9984 (N_9984,N_9680,N_9671);
nand U9985 (N_9985,N_9540,N_9654);
and U9986 (N_9986,N_9731,N_9632);
xor U9987 (N_9987,N_9709,N_9748);
or U9988 (N_9988,N_9671,N_9664);
nand U9989 (N_9989,N_9723,N_9542);
nor U9990 (N_9990,N_9679,N_9535);
nor U9991 (N_9991,N_9622,N_9563);
xnor U9992 (N_9992,N_9575,N_9648);
and U9993 (N_9993,N_9581,N_9570);
and U9994 (N_9994,N_9513,N_9735);
nand U9995 (N_9995,N_9736,N_9685);
and U9996 (N_9996,N_9673,N_9671);
and U9997 (N_9997,N_9716,N_9692);
xor U9998 (N_9998,N_9575,N_9580);
nand U9999 (N_9999,N_9652,N_9625);
or U10000 (N_10000,N_9821,N_9785);
and U10001 (N_10001,N_9844,N_9774);
and U10002 (N_10002,N_9971,N_9803);
xnor U10003 (N_10003,N_9851,N_9984);
nand U10004 (N_10004,N_9980,N_9827);
and U10005 (N_10005,N_9962,N_9881);
nand U10006 (N_10006,N_9887,N_9903);
and U10007 (N_10007,N_9752,N_9798);
nor U10008 (N_10008,N_9869,N_9852);
xnor U10009 (N_10009,N_9922,N_9890);
nor U10010 (N_10010,N_9975,N_9812);
nand U10011 (N_10011,N_9983,N_9907);
nand U10012 (N_10012,N_9856,N_9918);
nor U10013 (N_10013,N_9895,N_9846);
or U10014 (N_10014,N_9837,N_9986);
nor U10015 (N_10015,N_9875,N_9835);
nand U10016 (N_10016,N_9843,N_9972);
nor U10017 (N_10017,N_9896,N_9863);
and U10018 (N_10018,N_9860,N_9910);
and U10019 (N_10019,N_9911,N_9782);
xor U10020 (N_10020,N_9871,N_9955);
or U10021 (N_10021,N_9943,N_9964);
nor U10022 (N_10022,N_9909,N_9938);
nand U10023 (N_10023,N_9832,N_9839);
and U10024 (N_10024,N_9865,N_9781);
or U10025 (N_10025,N_9829,N_9770);
nand U10026 (N_10026,N_9768,N_9796);
and U10027 (N_10027,N_9967,N_9797);
nand U10028 (N_10028,N_9959,N_9961);
xor U10029 (N_10029,N_9892,N_9914);
xor U10030 (N_10030,N_9998,N_9969);
and U10031 (N_10031,N_9970,N_9762);
and U10032 (N_10032,N_9826,N_9883);
or U10033 (N_10033,N_9816,N_9989);
nor U10034 (N_10034,N_9756,N_9953);
and U10035 (N_10035,N_9800,N_9951);
and U10036 (N_10036,N_9985,N_9791);
nand U10037 (N_10037,N_9999,N_9857);
and U10038 (N_10038,N_9849,N_9947);
nand U10039 (N_10039,N_9927,N_9818);
and U10040 (N_10040,N_9765,N_9870);
nor U10041 (N_10041,N_9926,N_9993);
and U10042 (N_10042,N_9994,N_9793);
or U10043 (N_10043,N_9976,N_9919);
nand U10044 (N_10044,N_9758,N_9861);
and U10045 (N_10045,N_9982,N_9995);
and U10046 (N_10046,N_9804,N_9834);
nor U10047 (N_10047,N_9990,N_9991);
or U10048 (N_10048,N_9905,N_9815);
nor U10049 (N_10049,N_9935,N_9788);
nor U10050 (N_10050,N_9862,N_9924);
nor U10051 (N_10051,N_9965,N_9992);
or U10052 (N_10052,N_9802,N_9946);
xor U10053 (N_10053,N_9787,N_9866);
nand U10054 (N_10054,N_9928,N_9878);
xor U10055 (N_10055,N_9831,N_9859);
xor U10056 (N_10056,N_9894,N_9784);
and U10057 (N_10057,N_9763,N_9987);
or U10058 (N_10058,N_9819,N_9886);
nor U10059 (N_10059,N_9900,N_9840);
and U10060 (N_10060,N_9941,N_9957);
or U10061 (N_10061,N_9944,N_9855);
nand U10062 (N_10062,N_9810,N_9902);
nand U10063 (N_10063,N_9974,N_9950);
and U10064 (N_10064,N_9917,N_9814);
and U10065 (N_10065,N_9889,N_9772);
nor U10066 (N_10066,N_9934,N_9897);
or U10067 (N_10067,N_9868,N_9874);
or U10068 (N_10068,N_9932,N_9916);
and U10069 (N_10069,N_9963,N_9966);
or U10070 (N_10070,N_9931,N_9755);
and U10071 (N_10071,N_9759,N_9915);
nor U10072 (N_10072,N_9939,N_9873);
nand U10073 (N_10073,N_9766,N_9893);
or U10074 (N_10074,N_9925,N_9771);
xor U10075 (N_10075,N_9754,N_9808);
and U10076 (N_10076,N_9960,N_9958);
nand U10077 (N_10077,N_9833,N_9864);
or U10078 (N_10078,N_9809,N_9945);
or U10079 (N_10079,N_9923,N_9811);
or U10080 (N_10080,N_9979,N_9876);
or U10081 (N_10081,N_9799,N_9776);
or U10082 (N_10082,N_9820,N_9930);
xnor U10083 (N_10083,N_9978,N_9805);
nand U10084 (N_10084,N_9764,N_9845);
or U10085 (N_10085,N_9801,N_9822);
and U10086 (N_10086,N_9778,N_9806);
nand U10087 (N_10087,N_9828,N_9948);
and U10088 (N_10088,N_9882,N_9906);
xnor U10089 (N_10089,N_9981,N_9968);
nor U10090 (N_10090,N_9977,N_9901);
nand U10091 (N_10091,N_9920,N_9854);
xor U10092 (N_10092,N_9973,N_9807);
nor U10093 (N_10093,N_9952,N_9792);
and U10094 (N_10094,N_9879,N_9988);
nand U10095 (N_10095,N_9779,N_9954);
and U10096 (N_10096,N_9767,N_9753);
or U10097 (N_10097,N_9997,N_9929);
or U10098 (N_10098,N_9817,N_9761);
and U10099 (N_10099,N_9850,N_9780);
nand U10100 (N_10100,N_9830,N_9841);
nor U10101 (N_10101,N_9933,N_9912);
nor U10102 (N_10102,N_9885,N_9777);
and U10103 (N_10103,N_9775,N_9956);
and U10104 (N_10104,N_9888,N_9872);
and U10105 (N_10105,N_9773,N_9904);
and U10106 (N_10106,N_9853,N_9838);
nor U10107 (N_10107,N_9790,N_9823);
nor U10108 (N_10108,N_9842,N_9750);
or U10109 (N_10109,N_9908,N_9751);
xor U10110 (N_10110,N_9891,N_9913);
or U10111 (N_10111,N_9936,N_9940);
xor U10112 (N_10112,N_9847,N_9813);
xnor U10113 (N_10113,N_9880,N_9789);
nand U10114 (N_10114,N_9783,N_9848);
nor U10115 (N_10115,N_9836,N_9858);
nor U10116 (N_10116,N_9824,N_9884);
and U10117 (N_10117,N_9949,N_9942);
or U10118 (N_10118,N_9899,N_9825);
and U10119 (N_10119,N_9898,N_9795);
nor U10120 (N_10120,N_9877,N_9937);
and U10121 (N_10121,N_9757,N_9996);
xnor U10122 (N_10122,N_9867,N_9921);
nand U10123 (N_10123,N_9794,N_9769);
or U10124 (N_10124,N_9760,N_9786);
xor U10125 (N_10125,N_9848,N_9844);
nand U10126 (N_10126,N_9865,N_9774);
nand U10127 (N_10127,N_9750,N_9988);
xnor U10128 (N_10128,N_9993,N_9836);
nand U10129 (N_10129,N_9900,N_9839);
nand U10130 (N_10130,N_9895,N_9870);
and U10131 (N_10131,N_9807,N_9875);
nand U10132 (N_10132,N_9974,N_9806);
xor U10133 (N_10133,N_9806,N_9884);
nand U10134 (N_10134,N_9950,N_9911);
xnor U10135 (N_10135,N_9904,N_9842);
xor U10136 (N_10136,N_9780,N_9845);
nor U10137 (N_10137,N_9776,N_9970);
nor U10138 (N_10138,N_9894,N_9787);
nand U10139 (N_10139,N_9851,N_9793);
and U10140 (N_10140,N_9858,N_9866);
nor U10141 (N_10141,N_9928,N_9812);
and U10142 (N_10142,N_9974,N_9831);
xnor U10143 (N_10143,N_9933,N_9986);
and U10144 (N_10144,N_9917,N_9856);
or U10145 (N_10145,N_9943,N_9958);
xnor U10146 (N_10146,N_9996,N_9970);
xor U10147 (N_10147,N_9885,N_9958);
nand U10148 (N_10148,N_9751,N_9777);
xor U10149 (N_10149,N_9772,N_9890);
and U10150 (N_10150,N_9897,N_9930);
xor U10151 (N_10151,N_9795,N_9800);
and U10152 (N_10152,N_9927,N_9827);
nor U10153 (N_10153,N_9954,N_9990);
xnor U10154 (N_10154,N_9811,N_9834);
nand U10155 (N_10155,N_9908,N_9943);
nand U10156 (N_10156,N_9947,N_9920);
nor U10157 (N_10157,N_9950,N_9908);
nand U10158 (N_10158,N_9922,N_9875);
or U10159 (N_10159,N_9990,N_9876);
nand U10160 (N_10160,N_9912,N_9968);
or U10161 (N_10161,N_9858,N_9887);
or U10162 (N_10162,N_9932,N_9806);
nor U10163 (N_10163,N_9797,N_9989);
nand U10164 (N_10164,N_9878,N_9818);
xnor U10165 (N_10165,N_9815,N_9801);
or U10166 (N_10166,N_9873,N_9918);
nand U10167 (N_10167,N_9774,N_9834);
or U10168 (N_10168,N_9848,N_9798);
xnor U10169 (N_10169,N_9842,N_9783);
or U10170 (N_10170,N_9955,N_9872);
nor U10171 (N_10171,N_9998,N_9838);
or U10172 (N_10172,N_9782,N_9972);
nor U10173 (N_10173,N_9781,N_9867);
xnor U10174 (N_10174,N_9938,N_9848);
nand U10175 (N_10175,N_9765,N_9994);
nor U10176 (N_10176,N_9790,N_9753);
xnor U10177 (N_10177,N_9990,N_9862);
and U10178 (N_10178,N_9928,N_9917);
and U10179 (N_10179,N_9922,N_9955);
or U10180 (N_10180,N_9907,N_9815);
and U10181 (N_10181,N_9995,N_9965);
or U10182 (N_10182,N_9936,N_9968);
nor U10183 (N_10183,N_9818,N_9948);
nand U10184 (N_10184,N_9970,N_9808);
nor U10185 (N_10185,N_9873,N_9778);
and U10186 (N_10186,N_9796,N_9968);
xor U10187 (N_10187,N_9973,N_9958);
or U10188 (N_10188,N_9869,N_9839);
nor U10189 (N_10189,N_9983,N_9872);
nor U10190 (N_10190,N_9893,N_9800);
nor U10191 (N_10191,N_9864,N_9903);
nor U10192 (N_10192,N_9980,N_9924);
or U10193 (N_10193,N_9869,N_9972);
and U10194 (N_10194,N_9783,N_9773);
nand U10195 (N_10195,N_9941,N_9870);
xnor U10196 (N_10196,N_9895,N_9757);
and U10197 (N_10197,N_9816,N_9822);
xor U10198 (N_10198,N_9885,N_9908);
and U10199 (N_10199,N_9846,N_9950);
nor U10200 (N_10200,N_9994,N_9831);
xor U10201 (N_10201,N_9992,N_9814);
xnor U10202 (N_10202,N_9833,N_9866);
or U10203 (N_10203,N_9934,N_9907);
nand U10204 (N_10204,N_9956,N_9869);
or U10205 (N_10205,N_9954,N_9867);
or U10206 (N_10206,N_9884,N_9956);
nor U10207 (N_10207,N_9924,N_9893);
nand U10208 (N_10208,N_9756,N_9820);
and U10209 (N_10209,N_9990,N_9984);
and U10210 (N_10210,N_9933,N_9786);
nand U10211 (N_10211,N_9974,N_9759);
and U10212 (N_10212,N_9933,N_9914);
or U10213 (N_10213,N_9934,N_9988);
or U10214 (N_10214,N_9956,N_9970);
xor U10215 (N_10215,N_9920,N_9754);
or U10216 (N_10216,N_9944,N_9891);
nand U10217 (N_10217,N_9987,N_9816);
or U10218 (N_10218,N_9909,N_9831);
or U10219 (N_10219,N_9757,N_9758);
xnor U10220 (N_10220,N_9851,N_9838);
or U10221 (N_10221,N_9889,N_9900);
nand U10222 (N_10222,N_9760,N_9987);
or U10223 (N_10223,N_9907,N_9911);
or U10224 (N_10224,N_9982,N_9943);
nor U10225 (N_10225,N_9796,N_9995);
nor U10226 (N_10226,N_9915,N_9801);
nor U10227 (N_10227,N_9998,N_9940);
nand U10228 (N_10228,N_9957,N_9859);
xor U10229 (N_10229,N_9893,N_9870);
nand U10230 (N_10230,N_9888,N_9941);
or U10231 (N_10231,N_9767,N_9778);
nor U10232 (N_10232,N_9826,N_9995);
xnor U10233 (N_10233,N_9807,N_9797);
xnor U10234 (N_10234,N_9795,N_9783);
nand U10235 (N_10235,N_9997,N_9931);
or U10236 (N_10236,N_9779,N_9842);
nand U10237 (N_10237,N_9950,N_9823);
and U10238 (N_10238,N_9928,N_9763);
nand U10239 (N_10239,N_9772,N_9800);
or U10240 (N_10240,N_9805,N_9904);
xnor U10241 (N_10241,N_9990,N_9951);
nor U10242 (N_10242,N_9756,N_9776);
or U10243 (N_10243,N_9918,N_9802);
and U10244 (N_10244,N_9782,N_9846);
or U10245 (N_10245,N_9956,N_9930);
and U10246 (N_10246,N_9832,N_9928);
or U10247 (N_10247,N_9996,N_9819);
xor U10248 (N_10248,N_9822,N_9868);
nor U10249 (N_10249,N_9777,N_9967);
or U10250 (N_10250,N_10133,N_10019);
nand U10251 (N_10251,N_10249,N_10151);
and U10252 (N_10252,N_10193,N_10211);
or U10253 (N_10253,N_10238,N_10165);
nand U10254 (N_10254,N_10218,N_10173);
nor U10255 (N_10255,N_10206,N_10061);
xnor U10256 (N_10256,N_10091,N_10145);
nand U10257 (N_10257,N_10236,N_10096);
nor U10258 (N_10258,N_10106,N_10052);
nand U10259 (N_10259,N_10045,N_10202);
xor U10260 (N_10260,N_10198,N_10121);
xor U10261 (N_10261,N_10079,N_10178);
nor U10262 (N_10262,N_10036,N_10018);
or U10263 (N_10263,N_10186,N_10187);
and U10264 (N_10264,N_10053,N_10060);
xnor U10265 (N_10265,N_10093,N_10111);
or U10266 (N_10266,N_10188,N_10190);
and U10267 (N_10267,N_10203,N_10110);
nand U10268 (N_10268,N_10023,N_10022);
or U10269 (N_10269,N_10210,N_10137);
or U10270 (N_10270,N_10102,N_10179);
nor U10271 (N_10271,N_10195,N_10062);
and U10272 (N_10272,N_10055,N_10153);
and U10273 (N_10273,N_10215,N_10118);
nand U10274 (N_10274,N_10016,N_10072);
nand U10275 (N_10275,N_10152,N_10004);
nand U10276 (N_10276,N_10013,N_10054);
nand U10277 (N_10277,N_10124,N_10191);
nand U10278 (N_10278,N_10039,N_10162);
nand U10279 (N_10279,N_10122,N_10189);
or U10280 (N_10280,N_10107,N_10135);
or U10281 (N_10281,N_10014,N_10158);
nor U10282 (N_10282,N_10081,N_10119);
nand U10283 (N_10283,N_10012,N_10205);
or U10284 (N_10284,N_10174,N_10083);
and U10285 (N_10285,N_10000,N_10046);
and U10286 (N_10286,N_10037,N_10015);
or U10287 (N_10287,N_10235,N_10047);
nand U10288 (N_10288,N_10168,N_10155);
xor U10289 (N_10289,N_10177,N_10194);
or U10290 (N_10290,N_10148,N_10108);
and U10291 (N_10291,N_10007,N_10138);
and U10292 (N_10292,N_10200,N_10078);
or U10293 (N_10293,N_10059,N_10149);
xor U10294 (N_10294,N_10084,N_10204);
nor U10295 (N_10295,N_10243,N_10146);
or U10296 (N_10296,N_10025,N_10051);
xor U10297 (N_10297,N_10058,N_10031);
or U10298 (N_10298,N_10089,N_10160);
and U10299 (N_10299,N_10224,N_10131);
nand U10300 (N_10300,N_10132,N_10134);
or U10301 (N_10301,N_10150,N_10244);
nor U10302 (N_10302,N_10049,N_10073);
or U10303 (N_10303,N_10112,N_10097);
and U10304 (N_10304,N_10127,N_10065);
xor U10305 (N_10305,N_10011,N_10085);
xor U10306 (N_10306,N_10183,N_10209);
nor U10307 (N_10307,N_10067,N_10050);
nor U10308 (N_10308,N_10038,N_10092);
nand U10309 (N_10309,N_10114,N_10010);
nand U10310 (N_10310,N_10229,N_10120);
nand U10311 (N_10311,N_10199,N_10136);
nor U10312 (N_10312,N_10175,N_10113);
nand U10313 (N_10313,N_10032,N_10139);
nand U10314 (N_10314,N_10170,N_10233);
xor U10315 (N_10315,N_10003,N_10094);
or U10316 (N_10316,N_10125,N_10234);
xnor U10317 (N_10317,N_10217,N_10157);
and U10318 (N_10318,N_10213,N_10242);
and U10319 (N_10319,N_10180,N_10185);
xor U10320 (N_10320,N_10220,N_10212);
nor U10321 (N_10321,N_10129,N_10245);
or U10322 (N_10322,N_10115,N_10237);
nand U10323 (N_10323,N_10192,N_10164);
nor U10324 (N_10324,N_10028,N_10239);
and U10325 (N_10325,N_10071,N_10208);
and U10326 (N_10326,N_10247,N_10227);
nand U10327 (N_10327,N_10095,N_10020);
nand U10328 (N_10328,N_10057,N_10116);
xor U10329 (N_10329,N_10090,N_10214);
nand U10330 (N_10330,N_10098,N_10163);
nor U10331 (N_10331,N_10222,N_10197);
or U10332 (N_10332,N_10216,N_10104);
nand U10333 (N_10333,N_10117,N_10040);
xor U10334 (N_10334,N_10169,N_10063);
and U10335 (N_10335,N_10142,N_10017);
and U10336 (N_10336,N_10140,N_10033);
nor U10337 (N_10337,N_10184,N_10147);
nand U10338 (N_10338,N_10029,N_10221);
xnor U10339 (N_10339,N_10042,N_10126);
nor U10340 (N_10340,N_10248,N_10172);
nand U10341 (N_10341,N_10064,N_10026);
nor U10342 (N_10342,N_10034,N_10002);
or U10343 (N_10343,N_10167,N_10070);
xor U10344 (N_10344,N_10182,N_10075);
or U10345 (N_10345,N_10066,N_10207);
and U10346 (N_10346,N_10056,N_10144);
or U10347 (N_10347,N_10009,N_10035);
nor U10348 (N_10348,N_10099,N_10044);
or U10349 (N_10349,N_10231,N_10080);
nor U10350 (N_10350,N_10006,N_10219);
nand U10351 (N_10351,N_10109,N_10001);
nand U10352 (N_10352,N_10100,N_10086);
xor U10353 (N_10353,N_10069,N_10230);
nor U10354 (N_10354,N_10008,N_10176);
nor U10355 (N_10355,N_10024,N_10128);
and U10356 (N_10356,N_10005,N_10068);
nor U10357 (N_10357,N_10027,N_10043);
nor U10358 (N_10358,N_10166,N_10076);
or U10359 (N_10359,N_10077,N_10226);
nand U10360 (N_10360,N_10130,N_10223);
nand U10361 (N_10361,N_10228,N_10082);
and U10362 (N_10362,N_10041,N_10156);
nand U10363 (N_10363,N_10141,N_10087);
xnor U10364 (N_10364,N_10181,N_10030);
nand U10365 (N_10365,N_10105,N_10225);
nor U10366 (N_10366,N_10201,N_10171);
or U10367 (N_10367,N_10101,N_10240);
nand U10368 (N_10368,N_10048,N_10088);
and U10369 (N_10369,N_10161,N_10246);
or U10370 (N_10370,N_10143,N_10074);
and U10371 (N_10371,N_10123,N_10232);
or U10372 (N_10372,N_10196,N_10154);
xnor U10373 (N_10373,N_10103,N_10159);
xnor U10374 (N_10374,N_10241,N_10021);
and U10375 (N_10375,N_10051,N_10140);
xor U10376 (N_10376,N_10154,N_10166);
and U10377 (N_10377,N_10239,N_10016);
nor U10378 (N_10378,N_10165,N_10052);
xnor U10379 (N_10379,N_10076,N_10115);
xor U10380 (N_10380,N_10168,N_10225);
xnor U10381 (N_10381,N_10067,N_10167);
xnor U10382 (N_10382,N_10006,N_10164);
nor U10383 (N_10383,N_10227,N_10142);
nand U10384 (N_10384,N_10222,N_10239);
or U10385 (N_10385,N_10240,N_10040);
or U10386 (N_10386,N_10130,N_10242);
xnor U10387 (N_10387,N_10001,N_10243);
and U10388 (N_10388,N_10192,N_10010);
nand U10389 (N_10389,N_10230,N_10136);
nand U10390 (N_10390,N_10211,N_10202);
nor U10391 (N_10391,N_10143,N_10138);
and U10392 (N_10392,N_10117,N_10000);
or U10393 (N_10393,N_10070,N_10140);
or U10394 (N_10394,N_10073,N_10000);
nor U10395 (N_10395,N_10086,N_10087);
nand U10396 (N_10396,N_10013,N_10043);
and U10397 (N_10397,N_10193,N_10170);
nor U10398 (N_10398,N_10039,N_10160);
nor U10399 (N_10399,N_10239,N_10080);
nand U10400 (N_10400,N_10126,N_10015);
nand U10401 (N_10401,N_10032,N_10017);
nand U10402 (N_10402,N_10203,N_10003);
xor U10403 (N_10403,N_10182,N_10188);
and U10404 (N_10404,N_10187,N_10108);
nor U10405 (N_10405,N_10095,N_10143);
and U10406 (N_10406,N_10060,N_10087);
and U10407 (N_10407,N_10028,N_10228);
or U10408 (N_10408,N_10051,N_10056);
xnor U10409 (N_10409,N_10036,N_10200);
nor U10410 (N_10410,N_10174,N_10245);
nor U10411 (N_10411,N_10144,N_10005);
and U10412 (N_10412,N_10023,N_10115);
nand U10413 (N_10413,N_10109,N_10069);
xor U10414 (N_10414,N_10076,N_10202);
nor U10415 (N_10415,N_10153,N_10197);
and U10416 (N_10416,N_10108,N_10132);
nor U10417 (N_10417,N_10142,N_10185);
xor U10418 (N_10418,N_10116,N_10007);
nand U10419 (N_10419,N_10103,N_10055);
nor U10420 (N_10420,N_10207,N_10148);
xor U10421 (N_10421,N_10246,N_10081);
or U10422 (N_10422,N_10220,N_10103);
and U10423 (N_10423,N_10066,N_10141);
nor U10424 (N_10424,N_10022,N_10015);
and U10425 (N_10425,N_10072,N_10070);
or U10426 (N_10426,N_10046,N_10173);
nand U10427 (N_10427,N_10004,N_10082);
xnor U10428 (N_10428,N_10002,N_10036);
xnor U10429 (N_10429,N_10065,N_10244);
or U10430 (N_10430,N_10030,N_10117);
nand U10431 (N_10431,N_10005,N_10239);
nand U10432 (N_10432,N_10177,N_10066);
and U10433 (N_10433,N_10024,N_10188);
xor U10434 (N_10434,N_10075,N_10005);
or U10435 (N_10435,N_10200,N_10153);
and U10436 (N_10436,N_10160,N_10069);
xor U10437 (N_10437,N_10066,N_10087);
nand U10438 (N_10438,N_10123,N_10239);
xor U10439 (N_10439,N_10026,N_10077);
or U10440 (N_10440,N_10085,N_10249);
and U10441 (N_10441,N_10182,N_10176);
xnor U10442 (N_10442,N_10109,N_10114);
and U10443 (N_10443,N_10217,N_10006);
nand U10444 (N_10444,N_10106,N_10111);
or U10445 (N_10445,N_10165,N_10170);
nor U10446 (N_10446,N_10049,N_10037);
or U10447 (N_10447,N_10107,N_10007);
nand U10448 (N_10448,N_10143,N_10077);
or U10449 (N_10449,N_10186,N_10094);
nand U10450 (N_10450,N_10127,N_10047);
xnor U10451 (N_10451,N_10199,N_10109);
xor U10452 (N_10452,N_10245,N_10150);
and U10453 (N_10453,N_10218,N_10128);
nand U10454 (N_10454,N_10010,N_10211);
nand U10455 (N_10455,N_10116,N_10198);
xor U10456 (N_10456,N_10146,N_10129);
or U10457 (N_10457,N_10213,N_10171);
nor U10458 (N_10458,N_10161,N_10226);
nor U10459 (N_10459,N_10084,N_10221);
nor U10460 (N_10460,N_10107,N_10044);
nor U10461 (N_10461,N_10099,N_10071);
and U10462 (N_10462,N_10163,N_10232);
and U10463 (N_10463,N_10157,N_10023);
or U10464 (N_10464,N_10001,N_10159);
or U10465 (N_10465,N_10198,N_10223);
xnor U10466 (N_10466,N_10070,N_10024);
nand U10467 (N_10467,N_10019,N_10043);
xor U10468 (N_10468,N_10092,N_10239);
and U10469 (N_10469,N_10218,N_10031);
xor U10470 (N_10470,N_10024,N_10203);
and U10471 (N_10471,N_10175,N_10189);
nor U10472 (N_10472,N_10060,N_10135);
and U10473 (N_10473,N_10110,N_10141);
nor U10474 (N_10474,N_10141,N_10019);
xor U10475 (N_10475,N_10132,N_10237);
and U10476 (N_10476,N_10192,N_10122);
xor U10477 (N_10477,N_10006,N_10016);
nand U10478 (N_10478,N_10139,N_10070);
nand U10479 (N_10479,N_10158,N_10177);
and U10480 (N_10480,N_10231,N_10215);
xor U10481 (N_10481,N_10026,N_10223);
nor U10482 (N_10482,N_10069,N_10031);
or U10483 (N_10483,N_10180,N_10127);
nand U10484 (N_10484,N_10011,N_10125);
xnor U10485 (N_10485,N_10187,N_10099);
or U10486 (N_10486,N_10225,N_10093);
nand U10487 (N_10487,N_10061,N_10147);
xnor U10488 (N_10488,N_10063,N_10038);
nand U10489 (N_10489,N_10029,N_10081);
and U10490 (N_10490,N_10086,N_10073);
nand U10491 (N_10491,N_10007,N_10068);
or U10492 (N_10492,N_10070,N_10075);
or U10493 (N_10493,N_10203,N_10141);
nand U10494 (N_10494,N_10105,N_10133);
nand U10495 (N_10495,N_10058,N_10143);
or U10496 (N_10496,N_10170,N_10221);
nand U10497 (N_10497,N_10088,N_10234);
nor U10498 (N_10498,N_10035,N_10079);
xnor U10499 (N_10499,N_10239,N_10150);
nor U10500 (N_10500,N_10434,N_10485);
nand U10501 (N_10501,N_10402,N_10420);
nor U10502 (N_10502,N_10289,N_10353);
nand U10503 (N_10503,N_10340,N_10424);
xor U10504 (N_10504,N_10323,N_10268);
or U10505 (N_10505,N_10443,N_10326);
and U10506 (N_10506,N_10380,N_10331);
or U10507 (N_10507,N_10445,N_10429);
nand U10508 (N_10508,N_10479,N_10266);
xnor U10509 (N_10509,N_10361,N_10314);
nand U10510 (N_10510,N_10334,N_10294);
or U10511 (N_10511,N_10469,N_10405);
or U10512 (N_10512,N_10437,N_10349);
nor U10513 (N_10513,N_10292,N_10282);
nand U10514 (N_10514,N_10387,N_10254);
or U10515 (N_10515,N_10275,N_10465);
nand U10516 (N_10516,N_10423,N_10286);
nand U10517 (N_10517,N_10304,N_10371);
nor U10518 (N_10518,N_10398,N_10298);
xor U10519 (N_10519,N_10311,N_10263);
and U10520 (N_10520,N_10438,N_10478);
xnor U10521 (N_10521,N_10290,N_10394);
or U10522 (N_10522,N_10396,N_10346);
or U10523 (N_10523,N_10494,N_10372);
nor U10524 (N_10524,N_10354,N_10252);
nor U10525 (N_10525,N_10301,N_10368);
or U10526 (N_10526,N_10337,N_10255);
nand U10527 (N_10527,N_10392,N_10457);
and U10528 (N_10528,N_10381,N_10377);
xor U10529 (N_10529,N_10273,N_10393);
xnor U10530 (N_10530,N_10484,N_10345);
nand U10531 (N_10531,N_10476,N_10364);
and U10532 (N_10532,N_10447,N_10446);
and U10533 (N_10533,N_10285,N_10335);
xnor U10534 (N_10534,N_10497,N_10473);
nand U10535 (N_10535,N_10365,N_10369);
xor U10536 (N_10536,N_10449,N_10343);
or U10537 (N_10537,N_10297,N_10336);
nand U10538 (N_10538,N_10448,N_10281);
nor U10539 (N_10539,N_10270,N_10436);
nor U10540 (N_10540,N_10356,N_10302);
nor U10541 (N_10541,N_10486,N_10403);
xnor U10542 (N_10542,N_10458,N_10459);
nor U10543 (N_10543,N_10407,N_10262);
nor U10544 (N_10544,N_10491,N_10385);
and U10545 (N_10545,N_10279,N_10333);
and U10546 (N_10546,N_10330,N_10303);
nand U10547 (N_10547,N_10462,N_10341);
nor U10548 (N_10548,N_10451,N_10428);
and U10549 (N_10549,N_10439,N_10492);
xor U10550 (N_10550,N_10350,N_10321);
nor U10551 (N_10551,N_10362,N_10375);
nand U10552 (N_10552,N_10430,N_10278);
nor U10553 (N_10553,N_10418,N_10253);
xor U10554 (N_10554,N_10296,N_10440);
and U10555 (N_10555,N_10284,N_10342);
or U10556 (N_10556,N_10426,N_10419);
xor U10557 (N_10557,N_10348,N_10363);
nor U10558 (N_10558,N_10338,N_10299);
or U10559 (N_10559,N_10318,N_10455);
nand U10560 (N_10560,N_10312,N_10373);
and U10561 (N_10561,N_10260,N_10495);
xor U10562 (N_10562,N_10376,N_10325);
and U10563 (N_10563,N_10425,N_10309);
nor U10564 (N_10564,N_10322,N_10374);
nand U10565 (N_10565,N_10251,N_10499);
nor U10566 (N_10566,N_10327,N_10306);
nor U10567 (N_10567,N_10307,N_10489);
nor U10568 (N_10568,N_10295,N_10267);
nor U10569 (N_10569,N_10366,N_10328);
or U10570 (N_10570,N_10432,N_10280);
and U10571 (N_10571,N_10422,N_10498);
or U10572 (N_10572,N_10315,N_10468);
or U10573 (N_10573,N_10488,N_10287);
xor U10574 (N_10574,N_10355,N_10378);
nor U10575 (N_10575,N_10258,N_10433);
xor U10576 (N_10576,N_10388,N_10256);
nor U10577 (N_10577,N_10347,N_10480);
or U10578 (N_10578,N_10308,N_10397);
nand U10579 (N_10579,N_10300,N_10379);
nand U10580 (N_10580,N_10409,N_10305);
nand U10581 (N_10581,N_10454,N_10319);
and U10582 (N_10582,N_10435,N_10259);
nor U10583 (N_10583,N_10481,N_10370);
xnor U10584 (N_10584,N_10310,N_10464);
nand U10585 (N_10585,N_10264,N_10483);
or U10586 (N_10586,N_10400,N_10271);
nand U10587 (N_10587,N_10269,N_10367);
or U10588 (N_10588,N_10444,N_10399);
nand U10589 (N_10589,N_10329,N_10412);
and U10590 (N_10590,N_10415,N_10416);
or U10591 (N_10591,N_10389,N_10274);
and U10592 (N_10592,N_10339,N_10357);
xor U10593 (N_10593,N_10391,N_10261);
nand U10594 (N_10594,N_10472,N_10490);
and U10595 (N_10595,N_10360,N_10466);
nor U10596 (N_10596,N_10324,N_10293);
xnor U10597 (N_10597,N_10452,N_10450);
nor U10598 (N_10598,N_10283,N_10471);
xnor U10599 (N_10599,N_10320,N_10272);
or U10600 (N_10600,N_10250,N_10413);
or U10601 (N_10601,N_10359,N_10441);
nor U10602 (N_10602,N_10474,N_10404);
xnor U10603 (N_10603,N_10410,N_10401);
xnor U10604 (N_10604,N_10383,N_10386);
nand U10605 (N_10605,N_10358,N_10442);
and U10606 (N_10606,N_10390,N_10291);
or U10607 (N_10607,N_10431,N_10384);
or U10608 (N_10608,N_10352,N_10487);
nand U10609 (N_10609,N_10493,N_10421);
xnor U10610 (N_10610,N_10276,N_10313);
and U10611 (N_10611,N_10496,N_10317);
nand U10612 (N_10612,N_10257,N_10414);
nand U10613 (N_10613,N_10477,N_10288);
or U10614 (N_10614,N_10408,N_10467);
nand U10615 (N_10615,N_10427,N_10316);
and U10616 (N_10616,N_10332,N_10411);
xnor U10617 (N_10617,N_10406,N_10475);
or U10618 (N_10618,N_10395,N_10456);
or U10619 (N_10619,N_10482,N_10382);
nor U10620 (N_10620,N_10453,N_10460);
nand U10621 (N_10621,N_10265,N_10351);
and U10622 (N_10622,N_10417,N_10344);
nand U10623 (N_10623,N_10461,N_10463);
nor U10624 (N_10624,N_10277,N_10470);
or U10625 (N_10625,N_10304,N_10444);
nor U10626 (N_10626,N_10439,N_10485);
nor U10627 (N_10627,N_10338,N_10270);
xor U10628 (N_10628,N_10408,N_10407);
nor U10629 (N_10629,N_10375,N_10441);
or U10630 (N_10630,N_10391,N_10390);
nor U10631 (N_10631,N_10357,N_10414);
nor U10632 (N_10632,N_10483,N_10444);
nor U10633 (N_10633,N_10367,N_10309);
or U10634 (N_10634,N_10258,N_10322);
and U10635 (N_10635,N_10269,N_10271);
or U10636 (N_10636,N_10434,N_10498);
nand U10637 (N_10637,N_10417,N_10263);
and U10638 (N_10638,N_10413,N_10350);
xnor U10639 (N_10639,N_10376,N_10269);
or U10640 (N_10640,N_10324,N_10453);
nand U10641 (N_10641,N_10294,N_10250);
and U10642 (N_10642,N_10368,N_10390);
and U10643 (N_10643,N_10313,N_10373);
xnor U10644 (N_10644,N_10417,N_10410);
and U10645 (N_10645,N_10496,N_10300);
and U10646 (N_10646,N_10360,N_10296);
nor U10647 (N_10647,N_10322,N_10341);
nand U10648 (N_10648,N_10298,N_10320);
or U10649 (N_10649,N_10481,N_10311);
nor U10650 (N_10650,N_10299,N_10250);
and U10651 (N_10651,N_10483,N_10261);
or U10652 (N_10652,N_10277,N_10397);
nand U10653 (N_10653,N_10361,N_10328);
or U10654 (N_10654,N_10258,N_10340);
or U10655 (N_10655,N_10424,N_10254);
nor U10656 (N_10656,N_10422,N_10476);
nand U10657 (N_10657,N_10445,N_10398);
and U10658 (N_10658,N_10498,N_10329);
xnor U10659 (N_10659,N_10393,N_10346);
nor U10660 (N_10660,N_10287,N_10302);
nand U10661 (N_10661,N_10291,N_10259);
nand U10662 (N_10662,N_10280,N_10439);
nor U10663 (N_10663,N_10305,N_10274);
xor U10664 (N_10664,N_10376,N_10430);
and U10665 (N_10665,N_10321,N_10383);
or U10666 (N_10666,N_10395,N_10252);
and U10667 (N_10667,N_10258,N_10286);
or U10668 (N_10668,N_10487,N_10466);
nor U10669 (N_10669,N_10377,N_10394);
or U10670 (N_10670,N_10354,N_10373);
nand U10671 (N_10671,N_10421,N_10255);
and U10672 (N_10672,N_10465,N_10324);
xnor U10673 (N_10673,N_10266,N_10382);
xnor U10674 (N_10674,N_10329,N_10449);
and U10675 (N_10675,N_10292,N_10342);
xnor U10676 (N_10676,N_10256,N_10281);
or U10677 (N_10677,N_10429,N_10298);
xnor U10678 (N_10678,N_10384,N_10332);
nand U10679 (N_10679,N_10312,N_10298);
nor U10680 (N_10680,N_10268,N_10360);
or U10681 (N_10681,N_10262,N_10413);
xnor U10682 (N_10682,N_10343,N_10283);
nand U10683 (N_10683,N_10368,N_10436);
and U10684 (N_10684,N_10294,N_10379);
or U10685 (N_10685,N_10274,N_10430);
xnor U10686 (N_10686,N_10315,N_10422);
nand U10687 (N_10687,N_10256,N_10468);
or U10688 (N_10688,N_10497,N_10456);
and U10689 (N_10689,N_10440,N_10399);
nand U10690 (N_10690,N_10439,N_10476);
nand U10691 (N_10691,N_10305,N_10422);
or U10692 (N_10692,N_10377,N_10281);
xor U10693 (N_10693,N_10427,N_10293);
and U10694 (N_10694,N_10267,N_10371);
and U10695 (N_10695,N_10277,N_10394);
or U10696 (N_10696,N_10410,N_10363);
nor U10697 (N_10697,N_10465,N_10422);
xnor U10698 (N_10698,N_10306,N_10295);
nand U10699 (N_10699,N_10483,N_10299);
nor U10700 (N_10700,N_10411,N_10296);
or U10701 (N_10701,N_10435,N_10423);
nor U10702 (N_10702,N_10423,N_10465);
or U10703 (N_10703,N_10349,N_10320);
nand U10704 (N_10704,N_10485,N_10319);
xnor U10705 (N_10705,N_10480,N_10445);
nand U10706 (N_10706,N_10299,N_10405);
and U10707 (N_10707,N_10428,N_10256);
xor U10708 (N_10708,N_10352,N_10404);
nand U10709 (N_10709,N_10251,N_10274);
nor U10710 (N_10710,N_10276,N_10453);
xor U10711 (N_10711,N_10384,N_10441);
nand U10712 (N_10712,N_10312,N_10313);
and U10713 (N_10713,N_10406,N_10437);
nor U10714 (N_10714,N_10319,N_10313);
and U10715 (N_10715,N_10391,N_10465);
and U10716 (N_10716,N_10342,N_10289);
xor U10717 (N_10717,N_10322,N_10309);
xnor U10718 (N_10718,N_10367,N_10396);
xnor U10719 (N_10719,N_10306,N_10359);
nand U10720 (N_10720,N_10468,N_10473);
or U10721 (N_10721,N_10343,N_10432);
and U10722 (N_10722,N_10497,N_10355);
nor U10723 (N_10723,N_10488,N_10259);
nand U10724 (N_10724,N_10254,N_10466);
nor U10725 (N_10725,N_10415,N_10430);
and U10726 (N_10726,N_10309,N_10347);
nor U10727 (N_10727,N_10448,N_10337);
and U10728 (N_10728,N_10306,N_10354);
nor U10729 (N_10729,N_10351,N_10289);
and U10730 (N_10730,N_10254,N_10255);
nand U10731 (N_10731,N_10299,N_10400);
and U10732 (N_10732,N_10289,N_10495);
nand U10733 (N_10733,N_10355,N_10360);
nor U10734 (N_10734,N_10406,N_10364);
xor U10735 (N_10735,N_10462,N_10377);
xnor U10736 (N_10736,N_10347,N_10326);
nor U10737 (N_10737,N_10273,N_10488);
or U10738 (N_10738,N_10448,N_10476);
and U10739 (N_10739,N_10349,N_10343);
nor U10740 (N_10740,N_10270,N_10494);
nor U10741 (N_10741,N_10368,N_10287);
nand U10742 (N_10742,N_10468,N_10318);
xor U10743 (N_10743,N_10339,N_10341);
nor U10744 (N_10744,N_10301,N_10428);
nor U10745 (N_10745,N_10299,N_10491);
and U10746 (N_10746,N_10317,N_10458);
and U10747 (N_10747,N_10388,N_10450);
xnor U10748 (N_10748,N_10385,N_10489);
xor U10749 (N_10749,N_10449,N_10471);
or U10750 (N_10750,N_10647,N_10620);
xor U10751 (N_10751,N_10655,N_10571);
nand U10752 (N_10752,N_10684,N_10728);
or U10753 (N_10753,N_10521,N_10694);
xnor U10754 (N_10754,N_10656,N_10695);
xor U10755 (N_10755,N_10675,N_10651);
or U10756 (N_10756,N_10543,N_10729);
xor U10757 (N_10757,N_10631,N_10668);
or U10758 (N_10758,N_10744,N_10642);
or U10759 (N_10759,N_10560,N_10511);
xor U10760 (N_10760,N_10507,N_10649);
nand U10761 (N_10761,N_10673,N_10606);
nor U10762 (N_10762,N_10514,N_10699);
nand U10763 (N_10763,N_10632,N_10567);
nor U10764 (N_10764,N_10731,N_10563);
or U10765 (N_10765,N_10679,N_10584);
or U10766 (N_10766,N_10696,N_10628);
nand U10767 (N_10767,N_10671,N_10739);
and U10768 (N_10768,N_10509,N_10541);
nand U10769 (N_10769,N_10549,N_10515);
nand U10770 (N_10770,N_10539,N_10624);
and U10771 (N_10771,N_10576,N_10503);
xnor U10772 (N_10772,N_10715,N_10702);
nor U10773 (N_10773,N_10627,N_10733);
nand U10774 (N_10774,N_10551,N_10657);
xnor U10775 (N_10775,N_10603,N_10634);
xnor U10776 (N_10776,N_10615,N_10597);
nand U10777 (N_10777,N_10542,N_10552);
nor U10778 (N_10778,N_10504,N_10536);
xor U10779 (N_10779,N_10566,N_10550);
and U10780 (N_10780,N_10516,N_10578);
and U10781 (N_10781,N_10686,N_10609);
and U10782 (N_10782,N_10710,N_10742);
nor U10783 (N_10783,N_10640,N_10723);
and U10784 (N_10784,N_10681,N_10625);
and U10785 (N_10785,N_10582,N_10749);
nor U10786 (N_10786,N_10594,N_10724);
nor U10787 (N_10787,N_10577,N_10535);
nor U10788 (N_10788,N_10557,N_10730);
xnor U10789 (N_10789,N_10639,N_10689);
nor U10790 (N_10790,N_10717,N_10687);
and U10791 (N_10791,N_10741,N_10526);
or U10792 (N_10792,N_10545,N_10643);
and U10793 (N_10793,N_10629,N_10585);
nor U10794 (N_10794,N_10532,N_10646);
nor U10795 (N_10795,N_10623,N_10579);
nor U10796 (N_10796,N_10604,N_10562);
or U10797 (N_10797,N_10709,N_10570);
nand U10798 (N_10798,N_10700,N_10547);
nor U10799 (N_10799,N_10569,N_10559);
and U10800 (N_10800,N_10630,N_10614);
xnor U10801 (N_10801,N_10540,N_10645);
nor U10802 (N_10802,N_10678,N_10591);
and U10803 (N_10803,N_10564,N_10574);
and U10804 (N_10804,N_10530,N_10572);
nand U10805 (N_10805,N_10711,N_10590);
xnor U10806 (N_10806,N_10661,N_10602);
and U10807 (N_10807,N_10667,N_10708);
or U10808 (N_10808,N_10683,N_10748);
and U10809 (N_10809,N_10593,N_10722);
xor U10810 (N_10810,N_10621,N_10666);
xor U10811 (N_10811,N_10662,N_10519);
or U10812 (N_10812,N_10523,N_10727);
or U10813 (N_10813,N_10619,N_10644);
or U10814 (N_10814,N_10726,N_10537);
or U10815 (N_10815,N_10600,N_10586);
nor U10816 (N_10816,N_10589,N_10598);
or U10817 (N_10817,N_10654,N_10725);
and U10818 (N_10818,N_10738,N_10510);
xnor U10819 (N_10819,N_10529,N_10554);
xnor U10820 (N_10820,N_10613,N_10608);
nand U10821 (N_10821,N_10743,N_10565);
nand U10822 (N_10822,N_10525,N_10553);
xnor U10823 (N_10823,N_10713,N_10735);
nor U10824 (N_10824,N_10605,N_10622);
nor U10825 (N_10825,N_10517,N_10610);
nand U10826 (N_10826,N_10659,N_10534);
or U10827 (N_10827,N_10538,N_10527);
and U10828 (N_10828,N_10693,N_10658);
and U10829 (N_10829,N_10531,N_10664);
xor U10830 (N_10830,N_10670,N_10692);
nand U10831 (N_10831,N_10719,N_10601);
xnor U10832 (N_10832,N_10502,N_10583);
and U10833 (N_10833,N_10618,N_10555);
xor U10834 (N_10834,N_10690,N_10611);
xnor U10835 (N_10835,N_10691,N_10703);
nand U10836 (N_10836,N_10716,N_10500);
and U10837 (N_10837,N_10513,N_10704);
xnor U10838 (N_10838,N_10718,N_10740);
nand U10839 (N_10839,N_10669,N_10665);
xor U10840 (N_10840,N_10677,N_10501);
or U10841 (N_10841,N_10746,N_10524);
nor U10842 (N_10842,N_10548,N_10546);
or U10843 (N_10843,N_10637,N_10592);
xor U10844 (N_10844,N_10544,N_10573);
xor U10845 (N_10845,N_10745,N_10626);
nand U10846 (N_10846,N_10561,N_10732);
and U10847 (N_10847,N_10558,N_10580);
xor U10848 (N_10848,N_10688,N_10672);
and U10849 (N_10849,N_10505,N_10706);
xnor U10850 (N_10850,N_10641,N_10697);
nand U10851 (N_10851,N_10648,N_10701);
and U10852 (N_10852,N_10721,N_10714);
xnor U10853 (N_10853,N_10650,N_10734);
nor U10854 (N_10854,N_10680,N_10674);
and U10855 (N_10855,N_10633,N_10612);
nand U10856 (N_10856,N_10581,N_10506);
or U10857 (N_10857,N_10705,N_10682);
and U10858 (N_10858,N_10660,N_10663);
and U10859 (N_10859,N_10522,N_10607);
and U10860 (N_10860,N_10617,N_10595);
or U10861 (N_10861,N_10638,N_10747);
or U10862 (N_10862,N_10712,N_10653);
and U10863 (N_10863,N_10588,N_10599);
nor U10864 (N_10864,N_10575,N_10568);
xnor U10865 (N_10865,N_10587,N_10685);
nor U10866 (N_10866,N_10698,N_10520);
or U10867 (N_10867,N_10512,N_10707);
nor U10868 (N_10868,N_10676,N_10556);
nand U10869 (N_10869,N_10508,N_10720);
or U10870 (N_10870,N_10616,N_10736);
nor U10871 (N_10871,N_10533,N_10737);
nor U10872 (N_10872,N_10518,N_10652);
nor U10873 (N_10873,N_10636,N_10596);
and U10874 (N_10874,N_10635,N_10528);
nand U10875 (N_10875,N_10745,N_10631);
and U10876 (N_10876,N_10545,N_10584);
and U10877 (N_10877,N_10731,N_10713);
xor U10878 (N_10878,N_10674,N_10527);
nor U10879 (N_10879,N_10558,N_10711);
xor U10880 (N_10880,N_10693,N_10679);
nand U10881 (N_10881,N_10556,N_10740);
and U10882 (N_10882,N_10740,N_10582);
nand U10883 (N_10883,N_10564,N_10678);
nand U10884 (N_10884,N_10623,N_10663);
nor U10885 (N_10885,N_10582,N_10686);
xor U10886 (N_10886,N_10527,N_10549);
xnor U10887 (N_10887,N_10715,N_10704);
xor U10888 (N_10888,N_10675,N_10662);
and U10889 (N_10889,N_10515,N_10676);
and U10890 (N_10890,N_10743,N_10664);
nor U10891 (N_10891,N_10547,N_10641);
or U10892 (N_10892,N_10624,N_10746);
xnor U10893 (N_10893,N_10650,N_10738);
and U10894 (N_10894,N_10628,N_10606);
nor U10895 (N_10895,N_10666,N_10712);
and U10896 (N_10896,N_10586,N_10658);
nand U10897 (N_10897,N_10589,N_10699);
and U10898 (N_10898,N_10647,N_10679);
and U10899 (N_10899,N_10704,N_10618);
or U10900 (N_10900,N_10577,N_10573);
nand U10901 (N_10901,N_10548,N_10733);
xor U10902 (N_10902,N_10574,N_10523);
nor U10903 (N_10903,N_10556,N_10561);
nor U10904 (N_10904,N_10593,N_10543);
nor U10905 (N_10905,N_10544,N_10650);
or U10906 (N_10906,N_10538,N_10682);
xnor U10907 (N_10907,N_10698,N_10631);
and U10908 (N_10908,N_10748,N_10676);
or U10909 (N_10909,N_10673,N_10675);
and U10910 (N_10910,N_10697,N_10648);
nand U10911 (N_10911,N_10652,N_10724);
or U10912 (N_10912,N_10614,N_10646);
or U10913 (N_10913,N_10558,N_10645);
nand U10914 (N_10914,N_10738,N_10543);
nor U10915 (N_10915,N_10681,N_10624);
nor U10916 (N_10916,N_10682,N_10666);
nand U10917 (N_10917,N_10578,N_10649);
nor U10918 (N_10918,N_10606,N_10503);
or U10919 (N_10919,N_10541,N_10647);
xnor U10920 (N_10920,N_10544,N_10552);
xnor U10921 (N_10921,N_10618,N_10615);
and U10922 (N_10922,N_10533,N_10562);
nor U10923 (N_10923,N_10575,N_10635);
nand U10924 (N_10924,N_10540,N_10733);
or U10925 (N_10925,N_10597,N_10662);
and U10926 (N_10926,N_10631,N_10502);
nand U10927 (N_10927,N_10624,N_10540);
nor U10928 (N_10928,N_10695,N_10634);
nor U10929 (N_10929,N_10727,N_10689);
or U10930 (N_10930,N_10517,N_10690);
nor U10931 (N_10931,N_10621,N_10550);
and U10932 (N_10932,N_10670,N_10583);
xor U10933 (N_10933,N_10650,N_10502);
or U10934 (N_10934,N_10626,N_10522);
nor U10935 (N_10935,N_10649,N_10607);
nand U10936 (N_10936,N_10644,N_10503);
or U10937 (N_10937,N_10546,N_10578);
nor U10938 (N_10938,N_10580,N_10616);
nor U10939 (N_10939,N_10500,N_10743);
nand U10940 (N_10940,N_10677,N_10592);
and U10941 (N_10941,N_10726,N_10634);
nand U10942 (N_10942,N_10730,N_10508);
xor U10943 (N_10943,N_10535,N_10695);
xor U10944 (N_10944,N_10663,N_10747);
nor U10945 (N_10945,N_10563,N_10517);
and U10946 (N_10946,N_10519,N_10714);
nor U10947 (N_10947,N_10732,N_10563);
nand U10948 (N_10948,N_10565,N_10590);
nand U10949 (N_10949,N_10669,N_10682);
nor U10950 (N_10950,N_10664,N_10716);
xnor U10951 (N_10951,N_10662,N_10640);
nor U10952 (N_10952,N_10543,N_10658);
and U10953 (N_10953,N_10727,N_10554);
nor U10954 (N_10954,N_10574,N_10698);
nor U10955 (N_10955,N_10629,N_10611);
nand U10956 (N_10956,N_10647,N_10639);
nand U10957 (N_10957,N_10652,N_10699);
nand U10958 (N_10958,N_10574,N_10732);
nand U10959 (N_10959,N_10523,N_10564);
xor U10960 (N_10960,N_10554,N_10505);
xor U10961 (N_10961,N_10596,N_10534);
xnor U10962 (N_10962,N_10541,N_10656);
or U10963 (N_10963,N_10540,N_10686);
nor U10964 (N_10964,N_10707,N_10588);
nor U10965 (N_10965,N_10571,N_10746);
nand U10966 (N_10966,N_10737,N_10698);
or U10967 (N_10967,N_10569,N_10530);
nor U10968 (N_10968,N_10500,N_10711);
nand U10969 (N_10969,N_10643,N_10632);
or U10970 (N_10970,N_10726,N_10617);
xor U10971 (N_10971,N_10621,N_10532);
or U10972 (N_10972,N_10591,N_10739);
xnor U10973 (N_10973,N_10513,N_10706);
and U10974 (N_10974,N_10706,N_10675);
xor U10975 (N_10975,N_10674,N_10591);
nand U10976 (N_10976,N_10525,N_10712);
nand U10977 (N_10977,N_10530,N_10693);
nor U10978 (N_10978,N_10592,N_10538);
or U10979 (N_10979,N_10658,N_10657);
and U10980 (N_10980,N_10543,N_10649);
nor U10981 (N_10981,N_10741,N_10609);
nand U10982 (N_10982,N_10671,N_10702);
nor U10983 (N_10983,N_10600,N_10557);
xor U10984 (N_10984,N_10625,N_10597);
or U10985 (N_10985,N_10616,N_10526);
nand U10986 (N_10986,N_10576,N_10537);
xnor U10987 (N_10987,N_10651,N_10566);
nand U10988 (N_10988,N_10582,N_10563);
nand U10989 (N_10989,N_10509,N_10651);
nor U10990 (N_10990,N_10541,N_10710);
xnor U10991 (N_10991,N_10734,N_10564);
nand U10992 (N_10992,N_10725,N_10555);
and U10993 (N_10993,N_10630,N_10599);
and U10994 (N_10994,N_10514,N_10542);
xor U10995 (N_10995,N_10508,N_10676);
and U10996 (N_10996,N_10606,N_10675);
or U10997 (N_10997,N_10587,N_10675);
and U10998 (N_10998,N_10694,N_10597);
or U10999 (N_10999,N_10704,N_10632);
nand U11000 (N_11000,N_10988,N_10809);
xnor U11001 (N_11001,N_10885,N_10787);
or U11002 (N_11002,N_10996,N_10991);
nand U11003 (N_11003,N_10810,N_10755);
nand U11004 (N_11004,N_10928,N_10877);
nand U11005 (N_11005,N_10980,N_10857);
and U11006 (N_11006,N_10802,N_10976);
nand U11007 (N_11007,N_10927,N_10785);
or U11008 (N_11008,N_10845,N_10938);
and U11009 (N_11009,N_10948,N_10925);
and U11010 (N_11010,N_10812,N_10935);
or U11011 (N_11011,N_10933,N_10867);
nand U11012 (N_11012,N_10796,N_10889);
nor U11013 (N_11013,N_10997,N_10825);
and U11014 (N_11014,N_10972,N_10816);
or U11015 (N_11015,N_10828,N_10945);
nand U11016 (N_11016,N_10846,N_10890);
or U11017 (N_11017,N_10773,N_10932);
or U11018 (N_11018,N_10999,N_10758);
or U11019 (N_11019,N_10908,N_10987);
nor U11020 (N_11020,N_10793,N_10887);
xnor U11021 (N_11021,N_10841,N_10926);
and U11022 (N_11022,N_10818,N_10788);
nand U11023 (N_11023,N_10916,N_10849);
or U11024 (N_11024,N_10803,N_10778);
and U11025 (N_11025,N_10993,N_10865);
xnor U11026 (N_11026,N_10878,N_10899);
nand U11027 (N_11027,N_10943,N_10963);
or U11028 (N_11028,N_10995,N_10921);
nand U11029 (N_11029,N_10880,N_10941);
xnor U11030 (N_11030,N_10859,N_10842);
or U11031 (N_11031,N_10897,N_10750);
or U11032 (N_11032,N_10962,N_10836);
xnor U11033 (N_11033,N_10811,N_10918);
nand U11034 (N_11034,N_10807,N_10754);
or U11035 (N_11035,N_10798,N_10886);
nand U11036 (N_11036,N_10762,N_10990);
and U11037 (N_11037,N_10830,N_10883);
and U11038 (N_11038,N_10923,N_10879);
xor U11039 (N_11039,N_10871,N_10874);
nand U11040 (N_11040,N_10847,N_10806);
nand U11041 (N_11041,N_10882,N_10780);
nor U11042 (N_11042,N_10786,N_10982);
xor U11043 (N_11043,N_10813,N_10979);
nor U11044 (N_11044,N_10794,N_10821);
nand U11045 (N_11045,N_10912,N_10784);
and U11046 (N_11046,N_10770,N_10872);
nand U11047 (N_11047,N_10946,N_10992);
or U11048 (N_11048,N_10957,N_10851);
and U11049 (N_11049,N_10985,N_10920);
and U11050 (N_11050,N_10833,N_10792);
or U11051 (N_11051,N_10757,N_10984);
nand U11052 (N_11052,N_10856,N_10815);
xnor U11053 (N_11053,N_10902,N_10969);
or U11054 (N_11054,N_10771,N_10804);
and U11055 (N_11055,N_10903,N_10817);
xor U11056 (N_11056,N_10937,N_10942);
or U11057 (N_11057,N_10966,N_10983);
and U11058 (N_11058,N_10834,N_10853);
xor U11059 (N_11059,N_10873,N_10958);
and U11060 (N_11060,N_10860,N_10753);
nand U11061 (N_11061,N_10869,N_10961);
nor U11062 (N_11062,N_10881,N_10892);
nand U11063 (N_11063,N_10866,N_10783);
nand U11064 (N_11064,N_10875,N_10954);
xnor U11065 (N_11065,N_10823,N_10930);
or U11066 (N_11066,N_10952,N_10953);
nand U11067 (N_11067,N_10947,N_10863);
and U11068 (N_11068,N_10781,N_10968);
or U11069 (N_11069,N_10894,N_10905);
and U11070 (N_11070,N_10766,N_10919);
nor U11071 (N_11071,N_10805,N_10837);
or U11072 (N_11072,N_10751,N_10975);
or U11073 (N_11073,N_10955,N_10852);
nor U11074 (N_11074,N_10900,N_10964);
nor U11075 (N_11075,N_10765,N_10752);
nand U11076 (N_11076,N_10824,N_10891);
xor U11077 (N_11077,N_10826,N_10858);
nor U11078 (N_11078,N_10904,N_10864);
and U11079 (N_11079,N_10876,N_10949);
xor U11080 (N_11080,N_10772,N_10967);
and U11081 (N_11081,N_10978,N_10782);
nand U11082 (N_11082,N_10795,N_10769);
or U11083 (N_11083,N_10831,N_10909);
nor U11084 (N_11084,N_10922,N_10801);
nor U11085 (N_11085,N_10848,N_10832);
nand U11086 (N_11086,N_10819,N_10888);
nor U11087 (N_11087,N_10977,N_10763);
nand U11088 (N_11088,N_10911,N_10767);
and U11089 (N_11089,N_10861,N_10965);
or U11090 (N_11090,N_10915,N_10989);
or U11091 (N_11091,N_10956,N_10971);
xor U11092 (N_11092,N_10973,N_10940);
or U11093 (N_11093,N_10854,N_10814);
and U11094 (N_11094,N_10862,N_10820);
nand U11095 (N_11095,N_10827,N_10843);
or U11096 (N_11096,N_10808,N_10931);
xor U11097 (N_11097,N_10774,N_10907);
and U11098 (N_11098,N_10756,N_10776);
nor U11099 (N_11099,N_10944,N_10775);
nand U11100 (N_11100,N_10893,N_10896);
and U11101 (N_11101,N_10924,N_10768);
or U11102 (N_11102,N_10764,N_10901);
nor U11103 (N_11103,N_10790,N_10855);
and U11104 (N_11104,N_10981,N_10910);
and U11105 (N_11105,N_10950,N_10986);
nor U11106 (N_11106,N_10759,N_10898);
nor U11107 (N_11107,N_10914,N_10951);
and U11108 (N_11108,N_10936,N_10791);
nor U11109 (N_11109,N_10917,N_10829);
or U11110 (N_11110,N_10838,N_10929);
xnor U11111 (N_11111,N_10974,N_10913);
and U11112 (N_11112,N_10959,N_10870);
nor U11113 (N_11113,N_10970,N_10998);
nand U11114 (N_11114,N_10760,N_10939);
or U11115 (N_11115,N_10840,N_10895);
xor U11116 (N_11116,N_10850,N_10835);
xnor U11117 (N_11117,N_10800,N_10822);
or U11118 (N_11118,N_10839,N_10761);
nand U11119 (N_11119,N_10868,N_10934);
nor U11120 (N_11120,N_10844,N_10994);
and U11121 (N_11121,N_10789,N_10777);
or U11122 (N_11122,N_10884,N_10799);
nor U11123 (N_11123,N_10906,N_10797);
nand U11124 (N_11124,N_10960,N_10779);
nand U11125 (N_11125,N_10857,N_10853);
or U11126 (N_11126,N_10777,N_10925);
nand U11127 (N_11127,N_10858,N_10779);
nand U11128 (N_11128,N_10934,N_10802);
nor U11129 (N_11129,N_10783,N_10957);
nand U11130 (N_11130,N_10903,N_10994);
xnor U11131 (N_11131,N_10926,N_10868);
xnor U11132 (N_11132,N_10931,N_10880);
xnor U11133 (N_11133,N_10927,N_10827);
nand U11134 (N_11134,N_10972,N_10835);
nand U11135 (N_11135,N_10766,N_10856);
xor U11136 (N_11136,N_10929,N_10794);
nor U11137 (N_11137,N_10908,N_10909);
or U11138 (N_11138,N_10994,N_10864);
nand U11139 (N_11139,N_10896,N_10960);
nand U11140 (N_11140,N_10963,N_10828);
xnor U11141 (N_11141,N_10975,N_10873);
nand U11142 (N_11142,N_10885,N_10795);
and U11143 (N_11143,N_10855,N_10764);
or U11144 (N_11144,N_10759,N_10810);
nand U11145 (N_11145,N_10762,N_10944);
and U11146 (N_11146,N_10807,N_10809);
and U11147 (N_11147,N_10949,N_10797);
or U11148 (N_11148,N_10821,N_10884);
or U11149 (N_11149,N_10961,N_10776);
or U11150 (N_11150,N_10884,N_10832);
nand U11151 (N_11151,N_10827,N_10846);
or U11152 (N_11152,N_10956,N_10892);
nand U11153 (N_11153,N_10909,N_10766);
xnor U11154 (N_11154,N_10968,N_10773);
and U11155 (N_11155,N_10875,N_10758);
or U11156 (N_11156,N_10906,N_10899);
nor U11157 (N_11157,N_10947,N_10897);
nand U11158 (N_11158,N_10921,N_10811);
and U11159 (N_11159,N_10947,N_10890);
nand U11160 (N_11160,N_10976,N_10885);
xor U11161 (N_11161,N_10869,N_10819);
xor U11162 (N_11162,N_10952,N_10980);
and U11163 (N_11163,N_10822,N_10994);
nand U11164 (N_11164,N_10767,N_10989);
or U11165 (N_11165,N_10978,N_10861);
nor U11166 (N_11166,N_10799,N_10773);
xor U11167 (N_11167,N_10921,N_10964);
or U11168 (N_11168,N_10991,N_10902);
and U11169 (N_11169,N_10890,N_10807);
xor U11170 (N_11170,N_10942,N_10751);
nor U11171 (N_11171,N_10764,N_10935);
or U11172 (N_11172,N_10888,N_10850);
nor U11173 (N_11173,N_10897,N_10778);
xor U11174 (N_11174,N_10998,N_10809);
xor U11175 (N_11175,N_10977,N_10865);
nor U11176 (N_11176,N_10828,N_10852);
or U11177 (N_11177,N_10768,N_10901);
nand U11178 (N_11178,N_10995,N_10998);
nor U11179 (N_11179,N_10783,N_10752);
xnor U11180 (N_11180,N_10991,N_10756);
and U11181 (N_11181,N_10990,N_10892);
xnor U11182 (N_11182,N_10825,N_10976);
nor U11183 (N_11183,N_10859,N_10998);
xor U11184 (N_11184,N_10849,N_10909);
xnor U11185 (N_11185,N_10867,N_10907);
or U11186 (N_11186,N_10892,N_10913);
nand U11187 (N_11187,N_10827,N_10833);
and U11188 (N_11188,N_10796,N_10911);
and U11189 (N_11189,N_10950,N_10907);
xor U11190 (N_11190,N_10847,N_10990);
nor U11191 (N_11191,N_10910,N_10847);
nor U11192 (N_11192,N_10843,N_10859);
nand U11193 (N_11193,N_10913,N_10933);
and U11194 (N_11194,N_10964,N_10840);
nand U11195 (N_11195,N_10766,N_10803);
or U11196 (N_11196,N_10944,N_10822);
xnor U11197 (N_11197,N_10872,N_10920);
nand U11198 (N_11198,N_10911,N_10895);
and U11199 (N_11199,N_10905,N_10838);
nor U11200 (N_11200,N_10906,N_10852);
and U11201 (N_11201,N_10969,N_10931);
xnor U11202 (N_11202,N_10895,N_10975);
and U11203 (N_11203,N_10773,N_10755);
xnor U11204 (N_11204,N_10983,N_10947);
and U11205 (N_11205,N_10770,N_10871);
xor U11206 (N_11206,N_10818,N_10952);
nor U11207 (N_11207,N_10954,N_10860);
or U11208 (N_11208,N_10899,N_10990);
nor U11209 (N_11209,N_10865,N_10912);
nand U11210 (N_11210,N_10992,N_10901);
and U11211 (N_11211,N_10939,N_10864);
xor U11212 (N_11212,N_10990,N_10988);
or U11213 (N_11213,N_10962,N_10964);
nand U11214 (N_11214,N_10998,N_10925);
nand U11215 (N_11215,N_10918,N_10997);
and U11216 (N_11216,N_10759,N_10772);
and U11217 (N_11217,N_10921,N_10827);
or U11218 (N_11218,N_10767,N_10838);
xor U11219 (N_11219,N_10874,N_10996);
and U11220 (N_11220,N_10780,N_10880);
or U11221 (N_11221,N_10797,N_10819);
nand U11222 (N_11222,N_10977,N_10786);
xor U11223 (N_11223,N_10858,N_10979);
nand U11224 (N_11224,N_10760,N_10968);
nor U11225 (N_11225,N_10844,N_10775);
xor U11226 (N_11226,N_10916,N_10894);
xor U11227 (N_11227,N_10978,N_10827);
xnor U11228 (N_11228,N_10832,N_10757);
nand U11229 (N_11229,N_10751,N_10919);
nor U11230 (N_11230,N_10811,N_10781);
and U11231 (N_11231,N_10946,N_10822);
or U11232 (N_11232,N_10778,N_10980);
nor U11233 (N_11233,N_10998,N_10957);
xor U11234 (N_11234,N_10833,N_10800);
or U11235 (N_11235,N_10983,N_10784);
and U11236 (N_11236,N_10834,N_10815);
xor U11237 (N_11237,N_10813,N_10791);
nor U11238 (N_11238,N_10873,N_10892);
xor U11239 (N_11239,N_10847,N_10751);
and U11240 (N_11240,N_10814,N_10932);
nand U11241 (N_11241,N_10827,N_10866);
or U11242 (N_11242,N_10773,N_10852);
nor U11243 (N_11243,N_10875,N_10843);
nand U11244 (N_11244,N_10900,N_10871);
nor U11245 (N_11245,N_10837,N_10856);
and U11246 (N_11246,N_10826,N_10754);
xor U11247 (N_11247,N_10994,N_10855);
or U11248 (N_11248,N_10965,N_10853);
or U11249 (N_11249,N_10894,N_10941);
nand U11250 (N_11250,N_11222,N_11228);
and U11251 (N_11251,N_11115,N_11138);
and U11252 (N_11252,N_11140,N_11245);
xnor U11253 (N_11253,N_11061,N_11049);
nand U11254 (N_11254,N_11105,N_11167);
and U11255 (N_11255,N_11082,N_11178);
nand U11256 (N_11256,N_11176,N_11186);
nand U11257 (N_11257,N_11204,N_11032);
or U11258 (N_11258,N_11196,N_11109);
xnor U11259 (N_11259,N_11103,N_11119);
xnor U11260 (N_11260,N_11041,N_11120);
xnor U11261 (N_11261,N_11183,N_11084);
and U11262 (N_11262,N_11135,N_11189);
or U11263 (N_11263,N_11174,N_11063);
nor U11264 (N_11264,N_11158,N_11062);
and U11265 (N_11265,N_11170,N_11034);
or U11266 (N_11266,N_11166,N_11152);
and U11267 (N_11267,N_11190,N_11066);
nand U11268 (N_11268,N_11089,N_11142);
or U11269 (N_11269,N_11132,N_11141);
nor U11270 (N_11270,N_11097,N_11203);
xor U11271 (N_11271,N_11235,N_11100);
nand U11272 (N_11272,N_11005,N_11215);
xnor U11273 (N_11273,N_11056,N_11159);
or U11274 (N_11274,N_11013,N_11187);
and U11275 (N_11275,N_11127,N_11087);
nor U11276 (N_11276,N_11217,N_11216);
nand U11277 (N_11277,N_11081,N_11059);
xor U11278 (N_11278,N_11018,N_11210);
xnor U11279 (N_11279,N_11126,N_11072);
xnor U11280 (N_11280,N_11038,N_11171);
nand U11281 (N_11281,N_11133,N_11150);
nand U11282 (N_11282,N_11104,N_11108);
or U11283 (N_11283,N_11016,N_11212);
xnor U11284 (N_11284,N_11071,N_11244);
or U11285 (N_11285,N_11099,N_11191);
nand U11286 (N_11286,N_11045,N_11101);
nand U11287 (N_11287,N_11157,N_11147);
and U11288 (N_11288,N_11019,N_11047);
or U11289 (N_11289,N_11113,N_11060);
or U11290 (N_11290,N_11236,N_11232);
or U11291 (N_11291,N_11202,N_11207);
or U11292 (N_11292,N_11226,N_11035);
xor U11293 (N_11293,N_11246,N_11114);
nor U11294 (N_11294,N_11012,N_11181);
and U11295 (N_11295,N_11007,N_11078);
nand U11296 (N_11296,N_11095,N_11242);
and U11297 (N_11297,N_11224,N_11052);
or U11298 (N_11298,N_11117,N_11090);
xnor U11299 (N_11299,N_11091,N_11205);
or U11300 (N_11300,N_11000,N_11233);
xnor U11301 (N_11301,N_11102,N_11065);
xnor U11302 (N_11302,N_11198,N_11029);
and U11303 (N_11303,N_11163,N_11179);
xnor U11304 (N_11304,N_11249,N_11192);
or U11305 (N_11305,N_11037,N_11083);
nor U11306 (N_11306,N_11031,N_11027);
nor U11307 (N_11307,N_11200,N_11055);
nand U11308 (N_11308,N_11220,N_11214);
and U11309 (N_11309,N_11057,N_11094);
nor U11310 (N_11310,N_11014,N_11046);
nand U11311 (N_11311,N_11042,N_11088);
xnor U11312 (N_11312,N_11177,N_11161);
or U11313 (N_11313,N_11173,N_11002);
and U11314 (N_11314,N_11107,N_11172);
nor U11315 (N_11315,N_11069,N_11098);
nand U11316 (N_11316,N_11118,N_11247);
and U11317 (N_11317,N_11243,N_11051);
and U11318 (N_11318,N_11143,N_11086);
and U11319 (N_11319,N_11129,N_11064);
or U11320 (N_11320,N_11036,N_11006);
or U11321 (N_11321,N_11128,N_11206);
nor U11322 (N_11322,N_11225,N_11015);
xnor U11323 (N_11323,N_11221,N_11112);
and U11324 (N_11324,N_11044,N_11239);
xnor U11325 (N_11325,N_11218,N_11154);
nand U11326 (N_11326,N_11054,N_11085);
or U11327 (N_11327,N_11164,N_11134);
nand U11328 (N_11328,N_11155,N_11076);
nand U11329 (N_11329,N_11223,N_11211);
or U11330 (N_11330,N_11110,N_11208);
nand U11331 (N_11331,N_11197,N_11025);
and U11332 (N_11332,N_11003,N_11195);
xor U11333 (N_11333,N_11162,N_11106);
nand U11334 (N_11334,N_11023,N_11009);
or U11335 (N_11335,N_11093,N_11080);
or U11336 (N_11336,N_11017,N_11010);
xnor U11337 (N_11337,N_11182,N_11043);
and U11338 (N_11338,N_11096,N_11053);
nor U11339 (N_11339,N_11030,N_11169);
nor U11340 (N_11340,N_11048,N_11149);
and U11341 (N_11341,N_11122,N_11160);
or U11342 (N_11342,N_11240,N_11227);
or U11343 (N_11343,N_11201,N_11146);
or U11344 (N_11344,N_11008,N_11073);
nand U11345 (N_11345,N_11153,N_11230);
or U11346 (N_11346,N_11028,N_11168);
and U11347 (N_11347,N_11131,N_11213);
nand U11348 (N_11348,N_11123,N_11021);
xnor U11349 (N_11349,N_11199,N_11185);
and U11350 (N_11350,N_11039,N_11180);
nor U11351 (N_11351,N_11022,N_11175);
or U11352 (N_11352,N_11151,N_11001);
nand U11353 (N_11353,N_11116,N_11184);
xnor U11354 (N_11354,N_11011,N_11156);
nor U11355 (N_11355,N_11241,N_11231);
and U11356 (N_11356,N_11033,N_11075);
nor U11357 (N_11357,N_11004,N_11229);
and U11358 (N_11358,N_11070,N_11024);
nand U11359 (N_11359,N_11194,N_11219);
nand U11360 (N_11360,N_11248,N_11136);
nor U11361 (N_11361,N_11209,N_11040);
nor U11362 (N_11362,N_11137,N_11188);
xor U11363 (N_11363,N_11079,N_11068);
nor U11364 (N_11364,N_11125,N_11050);
nor U11365 (N_11365,N_11074,N_11067);
or U11366 (N_11366,N_11139,N_11026);
nand U11367 (N_11367,N_11058,N_11121);
nor U11368 (N_11368,N_11124,N_11144);
or U11369 (N_11369,N_11237,N_11077);
nor U11370 (N_11370,N_11020,N_11092);
and U11371 (N_11371,N_11238,N_11165);
nand U11372 (N_11372,N_11193,N_11111);
nand U11373 (N_11373,N_11148,N_11234);
and U11374 (N_11374,N_11145,N_11130);
and U11375 (N_11375,N_11080,N_11186);
and U11376 (N_11376,N_11074,N_11073);
xnor U11377 (N_11377,N_11010,N_11211);
xor U11378 (N_11378,N_11027,N_11216);
xnor U11379 (N_11379,N_11240,N_11146);
xnor U11380 (N_11380,N_11168,N_11103);
nand U11381 (N_11381,N_11125,N_11231);
nand U11382 (N_11382,N_11011,N_11194);
or U11383 (N_11383,N_11243,N_11028);
and U11384 (N_11384,N_11116,N_11185);
nand U11385 (N_11385,N_11035,N_11125);
or U11386 (N_11386,N_11225,N_11198);
and U11387 (N_11387,N_11125,N_11157);
nand U11388 (N_11388,N_11105,N_11196);
xor U11389 (N_11389,N_11062,N_11222);
and U11390 (N_11390,N_11155,N_11210);
nand U11391 (N_11391,N_11161,N_11000);
or U11392 (N_11392,N_11224,N_11226);
xnor U11393 (N_11393,N_11134,N_11152);
and U11394 (N_11394,N_11222,N_11058);
or U11395 (N_11395,N_11199,N_11092);
xnor U11396 (N_11396,N_11159,N_11130);
and U11397 (N_11397,N_11056,N_11091);
or U11398 (N_11398,N_11130,N_11146);
nor U11399 (N_11399,N_11130,N_11135);
nand U11400 (N_11400,N_11119,N_11037);
nand U11401 (N_11401,N_11097,N_11063);
and U11402 (N_11402,N_11061,N_11136);
and U11403 (N_11403,N_11100,N_11052);
nand U11404 (N_11404,N_11080,N_11135);
nor U11405 (N_11405,N_11014,N_11103);
and U11406 (N_11406,N_11188,N_11210);
xnor U11407 (N_11407,N_11196,N_11000);
nand U11408 (N_11408,N_11231,N_11035);
nand U11409 (N_11409,N_11016,N_11210);
nor U11410 (N_11410,N_11229,N_11123);
nand U11411 (N_11411,N_11107,N_11184);
xor U11412 (N_11412,N_11101,N_11013);
and U11413 (N_11413,N_11106,N_11163);
and U11414 (N_11414,N_11016,N_11144);
nor U11415 (N_11415,N_11161,N_11178);
or U11416 (N_11416,N_11210,N_11184);
nand U11417 (N_11417,N_11096,N_11060);
and U11418 (N_11418,N_11068,N_11157);
nand U11419 (N_11419,N_11085,N_11153);
and U11420 (N_11420,N_11151,N_11142);
or U11421 (N_11421,N_11094,N_11153);
nand U11422 (N_11422,N_11246,N_11128);
or U11423 (N_11423,N_11092,N_11226);
nand U11424 (N_11424,N_11132,N_11076);
xor U11425 (N_11425,N_11157,N_11110);
xnor U11426 (N_11426,N_11047,N_11235);
xnor U11427 (N_11427,N_11060,N_11065);
nand U11428 (N_11428,N_11105,N_11235);
nand U11429 (N_11429,N_11019,N_11017);
or U11430 (N_11430,N_11165,N_11019);
xor U11431 (N_11431,N_11070,N_11000);
nor U11432 (N_11432,N_11024,N_11092);
nor U11433 (N_11433,N_11157,N_11078);
and U11434 (N_11434,N_11017,N_11096);
and U11435 (N_11435,N_11197,N_11195);
or U11436 (N_11436,N_11114,N_11199);
nand U11437 (N_11437,N_11093,N_11127);
nand U11438 (N_11438,N_11249,N_11133);
or U11439 (N_11439,N_11206,N_11075);
or U11440 (N_11440,N_11196,N_11080);
nor U11441 (N_11441,N_11125,N_11167);
and U11442 (N_11442,N_11185,N_11084);
nor U11443 (N_11443,N_11136,N_11092);
and U11444 (N_11444,N_11108,N_11143);
and U11445 (N_11445,N_11200,N_11205);
nand U11446 (N_11446,N_11248,N_11196);
or U11447 (N_11447,N_11105,N_11074);
or U11448 (N_11448,N_11205,N_11225);
nor U11449 (N_11449,N_11212,N_11083);
nor U11450 (N_11450,N_11144,N_11008);
nor U11451 (N_11451,N_11248,N_11182);
xor U11452 (N_11452,N_11212,N_11224);
nand U11453 (N_11453,N_11039,N_11174);
xnor U11454 (N_11454,N_11032,N_11242);
and U11455 (N_11455,N_11160,N_11151);
or U11456 (N_11456,N_11144,N_11046);
or U11457 (N_11457,N_11087,N_11149);
and U11458 (N_11458,N_11064,N_11215);
nand U11459 (N_11459,N_11093,N_11075);
and U11460 (N_11460,N_11229,N_11013);
or U11461 (N_11461,N_11214,N_11225);
or U11462 (N_11462,N_11066,N_11151);
nor U11463 (N_11463,N_11246,N_11169);
xnor U11464 (N_11464,N_11239,N_11157);
nor U11465 (N_11465,N_11083,N_11141);
or U11466 (N_11466,N_11197,N_11085);
xnor U11467 (N_11467,N_11208,N_11023);
nand U11468 (N_11468,N_11039,N_11082);
nor U11469 (N_11469,N_11047,N_11112);
and U11470 (N_11470,N_11025,N_11177);
and U11471 (N_11471,N_11199,N_11094);
and U11472 (N_11472,N_11130,N_11060);
xor U11473 (N_11473,N_11059,N_11029);
nand U11474 (N_11474,N_11182,N_11013);
xnor U11475 (N_11475,N_11202,N_11126);
or U11476 (N_11476,N_11071,N_11135);
nand U11477 (N_11477,N_11190,N_11036);
nand U11478 (N_11478,N_11113,N_11242);
nand U11479 (N_11479,N_11153,N_11049);
nand U11480 (N_11480,N_11079,N_11040);
xor U11481 (N_11481,N_11224,N_11141);
nor U11482 (N_11482,N_11029,N_11193);
and U11483 (N_11483,N_11046,N_11160);
xor U11484 (N_11484,N_11249,N_11185);
nor U11485 (N_11485,N_11167,N_11119);
nand U11486 (N_11486,N_11219,N_11093);
or U11487 (N_11487,N_11003,N_11249);
nand U11488 (N_11488,N_11018,N_11236);
and U11489 (N_11489,N_11045,N_11190);
nor U11490 (N_11490,N_11063,N_11212);
nor U11491 (N_11491,N_11040,N_11183);
or U11492 (N_11492,N_11070,N_11087);
nand U11493 (N_11493,N_11164,N_11138);
nand U11494 (N_11494,N_11195,N_11133);
nand U11495 (N_11495,N_11227,N_11096);
nand U11496 (N_11496,N_11069,N_11143);
and U11497 (N_11497,N_11228,N_11185);
and U11498 (N_11498,N_11218,N_11213);
xnor U11499 (N_11499,N_11161,N_11022);
nand U11500 (N_11500,N_11304,N_11390);
nand U11501 (N_11501,N_11345,N_11455);
nor U11502 (N_11502,N_11473,N_11258);
and U11503 (N_11503,N_11404,N_11291);
nor U11504 (N_11504,N_11446,N_11443);
nand U11505 (N_11505,N_11391,N_11471);
and U11506 (N_11506,N_11482,N_11268);
xnor U11507 (N_11507,N_11269,N_11309);
nand U11508 (N_11508,N_11299,N_11419);
nor U11509 (N_11509,N_11479,N_11340);
and U11510 (N_11510,N_11481,N_11463);
and U11511 (N_11511,N_11396,N_11312);
and U11512 (N_11512,N_11460,N_11461);
xnor U11513 (N_11513,N_11397,N_11431);
nand U11514 (N_11514,N_11410,N_11470);
xnor U11515 (N_11515,N_11282,N_11284);
xor U11516 (N_11516,N_11307,N_11469);
or U11517 (N_11517,N_11358,N_11322);
and U11518 (N_11518,N_11294,N_11475);
nand U11519 (N_11519,N_11256,N_11306);
nor U11520 (N_11520,N_11462,N_11350);
or U11521 (N_11521,N_11428,N_11454);
xor U11522 (N_11522,N_11491,N_11417);
nand U11523 (N_11523,N_11476,N_11383);
nand U11524 (N_11524,N_11363,N_11495);
or U11525 (N_11525,N_11361,N_11347);
xor U11526 (N_11526,N_11381,N_11285);
nand U11527 (N_11527,N_11400,N_11424);
xor U11528 (N_11528,N_11368,N_11278);
xor U11529 (N_11529,N_11448,N_11364);
nand U11530 (N_11530,N_11274,N_11300);
and U11531 (N_11531,N_11366,N_11423);
or U11532 (N_11532,N_11490,N_11377);
nand U11533 (N_11533,N_11498,N_11408);
nor U11534 (N_11534,N_11324,N_11385);
or U11535 (N_11535,N_11326,N_11459);
xor U11536 (N_11536,N_11320,N_11325);
and U11537 (N_11537,N_11430,N_11394);
and U11538 (N_11538,N_11360,N_11365);
and U11539 (N_11539,N_11316,N_11254);
xnor U11540 (N_11540,N_11250,N_11323);
and U11541 (N_11541,N_11327,N_11338);
or U11542 (N_11542,N_11499,N_11331);
or U11543 (N_11543,N_11418,N_11493);
xor U11544 (N_11544,N_11378,N_11429);
nand U11545 (N_11545,N_11382,N_11478);
nand U11546 (N_11546,N_11287,N_11319);
and U11547 (N_11547,N_11439,N_11421);
and U11548 (N_11548,N_11405,N_11295);
and U11549 (N_11549,N_11388,N_11356);
or U11550 (N_11550,N_11355,N_11348);
nand U11551 (N_11551,N_11346,N_11426);
xnor U11552 (N_11552,N_11275,N_11286);
nor U11553 (N_11553,N_11341,N_11477);
nand U11554 (N_11554,N_11296,N_11425);
xnor U11555 (N_11555,N_11450,N_11487);
nor U11556 (N_11556,N_11456,N_11317);
or U11557 (N_11557,N_11472,N_11276);
or U11558 (N_11558,N_11465,N_11466);
and U11559 (N_11559,N_11259,N_11467);
nand U11560 (N_11560,N_11483,N_11384);
xor U11561 (N_11561,N_11442,N_11395);
nand U11562 (N_11562,N_11464,N_11281);
xnor U11563 (N_11563,N_11370,N_11451);
nand U11564 (N_11564,N_11313,N_11449);
xor U11565 (N_11565,N_11335,N_11349);
and U11566 (N_11566,N_11270,N_11399);
and U11567 (N_11567,N_11412,N_11458);
or U11568 (N_11568,N_11272,N_11407);
or U11569 (N_11569,N_11387,N_11271);
or U11570 (N_11570,N_11415,N_11436);
nor U11571 (N_11571,N_11416,N_11301);
or U11572 (N_11572,N_11380,N_11497);
nor U11573 (N_11573,N_11367,N_11265);
xnor U11574 (N_11574,N_11432,N_11289);
or U11575 (N_11575,N_11392,N_11283);
nand U11576 (N_11576,N_11266,N_11264);
or U11577 (N_11577,N_11371,N_11357);
nand U11578 (N_11578,N_11305,N_11343);
xor U11579 (N_11579,N_11318,N_11336);
or U11580 (N_11580,N_11420,N_11488);
nor U11581 (N_11581,N_11376,N_11393);
xor U11582 (N_11582,N_11311,N_11411);
and U11583 (N_11583,N_11257,N_11330);
nand U11584 (N_11584,N_11457,N_11386);
or U11585 (N_11585,N_11310,N_11292);
nor U11586 (N_11586,N_11298,N_11337);
and U11587 (N_11587,N_11444,N_11277);
nor U11588 (N_11588,N_11260,N_11433);
and U11589 (N_11589,N_11342,N_11369);
or U11590 (N_11590,N_11372,N_11303);
xnor U11591 (N_11591,N_11315,N_11445);
or U11592 (N_11592,N_11288,N_11252);
xnor U11593 (N_11593,N_11374,N_11362);
nor U11594 (N_11594,N_11486,N_11263);
nor U11595 (N_11595,N_11496,N_11402);
xor U11596 (N_11596,N_11489,N_11261);
and U11597 (N_11597,N_11353,N_11302);
xnor U11598 (N_11598,N_11447,N_11406);
or U11599 (N_11599,N_11437,N_11293);
or U11600 (N_11600,N_11438,N_11422);
nand U11601 (N_11601,N_11440,N_11297);
nand U11602 (N_11602,N_11480,N_11255);
and U11603 (N_11603,N_11262,N_11494);
nor U11604 (N_11604,N_11414,N_11441);
nor U11605 (N_11605,N_11329,N_11492);
nor U11606 (N_11606,N_11339,N_11452);
xnor U11607 (N_11607,N_11333,N_11375);
nand U11608 (N_11608,N_11427,N_11398);
or U11609 (N_11609,N_11379,N_11321);
xnor U11610 (N_11610,N_11290,N_11332);
or U11611 (N_11611,N_11314,N_11453);
and U11612 (N_11612,N_11485,N_11308);
or U11613 (N_11613,N_11403,N_11344);
nand U11614 (N_11614,N_11251,N_11389);
xor U11615 (N_11615,N_11413,N_11474);
nor U11616 (N_11616,N_11401,N_11354);
and U11617 (N_11617,N_11373,N_11328);
and U11618 (N_11618,N_11253,N_11434);
nor U11619 (N_11619,N_11334,N_11468);
or U11620 (N_11620,N_11484,N_11352);
nand U11621 (N_11621,N_11267,N_11273);
nand U11622 (N_11622,N_11359,N_11435);
nand U11623 (N_11623,N_11279,N_11409);
or U11624 (N_11624,N_11280,N_11351);
or U11625 (N_11625,N_11358,N_11490);
nor U11626 (N_11626,N_11479,N_11432);
nor U11627 (N_11627,N_11356,N_11275);
or U11628 (N_11628,N_11383,N_11366);
xor U11629 (N_11629,N_11272,N_11304);
nor U11630 (N_11630,N_11268,N_11381);
nand U11631 (N_11631,N_11333,N_11407);
nor U11632 (N_11632,N_11440,N_11436);
or U11633 (N_11633,N_11355,N_11396);
nand U11634 (N_11634,N_11329,N_11376);
and U11635 (N_11635,N_11419,N_11402);
nor U11636 (N_11636,N_11265,N_11472);
or U11637 (N_11637,N_11414,N_11301);
nor U11638 (N_11638,N_11468,N_11478);
or U11639 (N_11639,N_11367,N_11425);
nand U11640 (N_11640,N_11417,N_11431);
or U11641 (N_11641,N_11496,N_11446);
nand U11642 (N_11642,N_11423,N_11492);
xnor U11643 (N_11643,N_11327,N_11487);
and U11644 (N_11644,N_11433,N_11412);
nor U11645 (N_11645,N_11330,N_11287);
nor U11646 (N_11646,N_11473,N_11323);
or U11647 (N_11647,N_11416,N_11479);
nor U11648 (N_11648,N_11269,N_11492);
or U11649 (N_11649,N_11488,N_11424);
xor U11650 (N_11650,N_11454,N_11276);
or U11651 (N_11651,N_11463,N_11365);
or U11652 (N_11652,N_11274,N_11269);
nand U11653 (N_11653,N_11434,N_11331);
xor U11654 (N_11654,N_11311,N_11362);
xor U11655 (N_11655,N_11314,N_11317);
xnor U11656 (N_11656,N_11465,N_11475);
xor U11657 (N_11657,N_11431,N_11344);
nand U11658 (N_11658,N_11273,N_11415);
nor U11659 (N_11659,N_11288,N_11465);
or U11660 (N_11660,N_11416,N_11434);
nand U11661 (N_11661,N_11343,N_11386);
nor U11662 (N_11662,N_11272,N_11271);
nand U11663 (N_11663,N_11284,N_11432);
xor U11664 (N_11664,N_11418,N_11365);
xor U11665 (N_11665,N_11348,N_11349);
nand U11666 (N_11666,N_11471,N_11359);
nor U11667 (N_11667,N_11427,N_11403);
xor U11668 (N_11668,N_11258,N_11478);
and U11669 (N_11669,N_11340,N_11262);
and U11670 (N_11670,N_11423,N_11299);
or U11671 (N_11671,N_11302,N_11392);
nand U11672 (N_11672,N_11441,N_11348);
nand U11673 (N_11673,N_11411,N_11490);
nand U11674 (N_11674,N_11343,N_11347);
or U11675 (N_11675,N_11446,N_11265);
nor U11676 (N_11676,N_11436,N_11405);
nor U11677 (N_11677,N_11343,N_11383);
or U11678 (N_11678,N_11461,N_11414);
nor U11679 (N_11679,N_11312,N_11329);
nor U11680 (N_11680,N_11364,N_11438);
nor U11681 (N_11681,N_11396,N_11491);
and U11682 (N_11682,N_11436,N_11312);
nand U11683 (N_11683,N_11266,N_11392);
or U11684 (N_11684,N_11404,N_11334);
nand U11685 (N_11685,N_11499,N_11275);
or U11686 (N_11686,N_11418,N_11444);
nor U11687 (N_11687,N_11252,N_11420);
nor U11688 (N_11688,N_11350,N_11438);
nor U11689 (N_11689,N_11396,N_11254);
nor U11690 (N_11690,N_11470,N_11471);
nor U11691 (N_11691,N_11316,N_11485);
xnor U11692 (N_11692,N_11415,N_11360);
nor U11693 (N_11693,N_11288,N_11474);
xor U11694 (N_11694,N_11345,N_11452);
xnor U11695 (N_11695,N_11379,N_11429);
or U11696 (N_11696,N_11394,N_11440);
xnor U11697 (N_11697,N_11430,N_11490);
nor U11698 (N_11698,N_11482,N_11439);
or U11699 (N_11699,N_11301,N_11322);
and U11700 (N_11700,N_11321,N_11415);
or U11701 (N_11701,N_11415,N_11461);
and U11702 (N_11702,N_11368,N_11443);
nor U11703 (N_11703,N_11353,N_11493);
and U11704 (N_11704,N_11356,N_11358);
xor U11705 (N_11705,N_11314,N_11402);
nand U11706 (N_11706,N_11256,N_11370);
xnor U11707 (N_11707,N_11476,N_11266);
or U11708 (N_11708,N_11349,N_11326);
nand U11709 (N_11709,N_11358,N_11452);
or U11710 (N_11710,N_11281,N_11414);
and U11711 (N_11711,N_11275,N_11412);
or U11712 (N_11712,N_11346,N_11308);
nand U11713 (N_11713,N_11415,N_11399);
or U11714 (N_11714,N_11383,N_11370);
nor U11715 (N_11715,N_11254,N_11493);
or U11716 (N_11716,N_11421,N_11498);
or U11717 (N_11717,N_11475,N_11467);
nand U11718 (N_11718,N_11261,N_11364);
or U11719 (N_11719,N_11280,N_11481);
nor U11720 (N_11720,N_11323,N_11364);
and U11721 (N_11721,N_11345,N_11264);
xnor U11722 (N_11722,N_11261,N_11451);
and U11723 (N_11723,N_11393,N_11370);
nor U11724 (N_11724,N_11388,N_11382);
or U11725 (N_11725,N_11348,N_11304);
xor U11726 (N_11726,N_11335,N_11404);
and U11727 (N_11727,N_11329,N_11355);
nand U11728 (N_11728,N_11310,N_11315);
or U11729 (N_11729,N_11408,N_11274);
nand U11730 (N_11730,N_11418,N_11255);
xnor U11731 (N_11731,N_11344,N_11389);
nand U11732 (N_11732,N_11310,N_11323);
xnor U11733 (N_11733,N_11450,N_11362);
or U11734 (N_11734,N_11309,N_11282);
and U11735 (N_11735,N_11330,N_11335);
nor U11736 (N_11736,N_11413,N_11462);
or U11737 (N_11737,N_11447,N_11391);
nor U11738 (N_11738,N_11382,N_11340);
and U11739 (N_11739,N_11279,N_11438);
or U11740 (N_11740,N_11368,N_11454);
xor U11741 (N_11741,N_11494,N_11445);
nor U11742 (N_11742,N_11403,N_11387);
nor U11743 (N_11743,N_11261,N_11267);
nor U11744 (N_11744,N_11382,N_11353);
xnor U11745 (N_11745,N_11446,N_11485);
or U11746 (N_11746,N_11451,N_11391);
and U11747 (N_11747,N_11382,N_11269);
and U11748 (N_11748,N_11399,N_11374);
or U11749 (N_11749,N_11422,N_11369);
nor U11750 (N_11750,N_11610,N_11590);
nand U11751 (N_11751,N_11551,N_11674);
or U11752 (N_11752,N_11742,N_11648);
nor U11753 (N_11753,N_11646,N_11608);
nand U11754 (N_11754,N_11740,N_11552);
or U11755 (N_11755,N_11593,N_11591);
and U11756 (N_11756,N_11626,N_11620);
xnor U11757 (N_11757,N_11654,N_11549);
or U11758 (N_11758,N_11666,N_11669);
or U11759 (N_11759,N_11685,N_11525);
and U11760 (N_11760,N_11566,N_11625);
and U11761 (N_11761,N_11747,N_11511);
xor U11762 (N_11762,N_11731,N_11718);
and U11763 (N_11763,N_11540,N_11616);
nor U11764 (N_11764,N_11746,N_11567);
nor U11765 (N_11765,N_11678,N_11658);
or U11766 (N_11766,N_11596,N_11673);
or U11767 (N_11767,N_11519,N_11505);
or U11768 (N_11768,N_11638,N_11690);
or U11769 (N_11769,N_11529,N_11576);
nand U11770 (N_11770,N_11691,N_11619);
nand U11771 (N_11771,N_11513,N_11521);
nor U11772 (N_11772,N_11657,N_11595);
nand U11773 (N_11773,N_11688,N_11649);
or U11774 (N_11774,N_11635,N_11680);
nor U11775 (N_11775,N_11631,N_11651);
and U11776 (N_11776,N_11642,N_11719);
and U11777 (N_11777,N_11526,N_11583);
or U11778 (N_11778,N_11530,N_11588);
nand U11779 (N_11779,N_11737,N_11641);
nor U11780 (N_11780,N_11681,N_11512);
or U11781 (N_11781,N_11655,N_11546);
or U11782 (N_11782,N_11736,N_11697);
or U11783 (N_11783,N_11507,N_11671);
or U11784 (N_11784,N_11533,N_11621);
and U11785 (N_11785,N_11598,N_11689);
nand U11786 (N_11786,N_11677,N_11545);
nor U11787 (N_11787,N_11729,N_11716);
xnor U11788 (N_11788,N_11713,N_11502);
or U11789 (N_11789,N_11650,N_11696);
and U11790 (N_11790,N_11693,N_11587);
and U11791 (N_11791,N_11615,N_11622);
or U11792 (N_11792,N_11532,N_11647);
nor U11793 (N_11793,N_11535,N_11633);
xnor U11794 (N_11794,N_11701,N_11692);
nand U11795 (N_11795,N_11748,N_11714);
nor U11796 (N_11796,N_11732,N_11599);
xor U11797 (N_11797,N_11738,N_11522);
or U11798 (N_11798,N_11561,N_11634);
or U11799 (N_11799,N_11554,N_11664);
or U11800 (N_11800,N_11703,N_11605);
xor U11801 (N_11801,N_11594,N_11679);
and U11802 (N_11802,N_11668,N_11727);
or U11803 (N_11803,N_11744,N_11543);
xor U11804 (N_11804,N_11699,N_11580);
xor U11805 (N_11805,N_11506,N_11672);
and U11806 (N_11806,N_11745,N_11501);
nor U11807 (N_11807,N_11702,N_11636);
or U11808 (N_11808,N_11667,N_11710);
or U11809 (N_11809,N_11534,N_11720);
xor U11810 (N_11810,N_11508,N_11589);
and U11811 (N_11811,N_11586,N_11739);
nor U11812 (N_11812,N_11575,N_11640);
and U11813 (N_11813,N_11541,N_11618);
nand U11814 (N_11814,N_11565,N_11538);
and U11815 (N_11815,N_11694,N_11707);
or U11816 (N_11816,N_11527,N_11523);
and U11817 (N_11817,N_11609,N_11539);
nand U11818 (N_11818,N_11728,N_11741);
nand U11819 (N_11819,N_11695,N_11581);
nand U11820 (N_11820,N_11706,N_11717);
nand U11821 (N_11821,N_11684,N_11601);
and U11822 (N_11822,N_11686,N_11724);
nor U11823 (N_11823,N_11733,N_11687);
or U11824 (N_11824,N_11569,N_11544);
nand U11825 (N_11825,N_11585,N_11711);
xnor U11826 (N_11826,N_11571,N_11570);
and U11827 (N_11827,N_11725,N_11553);
nor U11828 (N_11828,N_11662,N_11564);
and U11829 (N_11829,N_11698,N_11584);
and U11830 (N_11830,N_11579,N_11665);
and U11831 (N_11831,N_11645,N_11602);
xnor U11832 (N_11832,N_11573,N_11557);
xor U11833 (N_11833,N_11700,N_11524);
or U11834 (N_11834,N_11516,N_11604);
or U11835 (N_11835,N_11542,N_11574);
and U11836 (N_11836,N_11734,N_11749);
and U11837 (N_11837,N_11709,N_11600);
nand U11838 (N_11838,N_11517,N_11556);
nand U11839 (N_11839,N_11632,N_11722);
and U11840 (N_11840,N_11676,N_11659);
nand U11841 (N_11841,N_11572,N_11726);
nor U11842 (N_11842,N_11509,N_11504);
nor U11843 (N_11843,N_11675,N_11550);
nor U11844 (N_11844,N_11653,N_11612);
xnor U11845 (N_11845,N_11627,N_11560);
nor U11846 (N_11846,N_11682,N_11515);
xor U11847 (N_11847,N_11558,N_11643);
or U11848 (N_11848,N_11568,N_11656);
or U11849 (N_11849,N_11639,N_11628);
or U11850 (N_11850,N_11624,N_11563);
nor U11851 (N_11851,N_11528,N_11537);
nor U11852 (N_11852,N_11547,N_11730);
nor U11853 (N_11853,N_11644,N_11518);
nor U11854 (N_11854,N_11712,N_11661);
xnor U11855 (N_11855,N_11531,N_11660);
or U11856 (N_11856,N_11652,N_11670);
and U11857 (N_11857,N_11510,N_11611);
or U11858 (N_11858,N_11708,N_11577);
nand U11859 (N_11859,N_11613,N_11559);
nand U11860 (N_11860,N_11723,N_11603);
nand U11861 (N_11861,N_11629,N_11743);
nor U11862 (N_11862,N_11623,N_11637);
nand U11863 (N_11863,N_11597,N_11555);
nor U11864 (N_11864,N_11630,N_11614);
or U11865 (N_11865,N_11607,N_11520);
nor U11866 (N_11866,N_11500,N_11592);
or U11867 (N_11867,N_11715,N_11663);
xor U11868 (N_11868,N_11514,N_11606);
or U11869 (N_11869,N_11548,N_11503);
nand U11870 (N_11870,N_11562,N_11683);
nand U11871 (N_11871,N_11536,N_11582);
and U11872 (N_11872,N_11578,N_11617);
nor U11873 (N_11873,N_11705,N_11735);
xnor U11874 (N_11874,N_11704,N_11721);
nand U11875 (N_11875,N_11708,N_11568);
or U11876 (N_11876,N_11640,N_11618);
nor U11877 (N_11877,N_11739,N_11663);
nor U11878 (N_11878,N_11710,N_11730);
or U11879 (N_11879,N_11523,N_11696);
nor U11880 (N_11880,N_11548,N_11500);
or U11881 (N_11881,N_11679,N_11619);
xnor U11882 (N_11882,N_11598,N_11607);
nand U11883 (N_11883,N_11611,N_11676);
nand U11884 (N_11884,N_11500,N_11740);
and U11885 (N_11885,N_11580,N_11711);
or U11886 (N_11886,N_11626,N_11695);
xor U11887 (N_11887,N_11564,N_11665);
nand U11888 (N_11888,N_11576,N_11748);
and U11889 (N_11889,N_11708,N_11524);
and U11890 (N_11890,N_11689,N_11519);
or U11891 (N_11891,N_11507,N_11720);
nand U11892 (N_11892,N_11602,N_11624);
or U11893 (N_11893,N_11703,N_11546);
and U11894 (N_11894,N_11609,N_11613);
nor U11895 (N_11895,N_11748,N_11695);
nand U11896 (N_11896,N_11611,N_11565);
or U11897 (N_11897,N_11702,N_11503);
nor U11898 (N_11898,N_11618,N_11647);
and U11899 (N_11899,N_11590,N_11521);
nor U11900 (N_11900,N_11722,N_11618);
and U11901 (N_11901,N_11664,N_11566);
nor U11902 (N_11902,N_11623,N_11715);
xor U11903 (N_11903,N_11701,N_11647);
or U11904 (N_11904,N_11525,N_11635);
xor U11905 (N_11905,N_11541,N_11744);
xnor U11906 (N_11906,N_11573,N_11662);
xor U11907 (N_11907,N_11566,N_11503);
xnor U11908 (N_11908,N_11677,N_11524);
xnor U11909 (N_11909,N_11744,N_11721);
xnor U11910 (N_11910,N_11691,N_11553);
nand U11911 (N_11911,N_11524,N_11633);
xor U11912 (N_11912,N_11739,N_11601);
or U11913 (N_11913,N_11513,N_11533);
and U11914 (N_11914,N_11685,N_11712);
or U11915 (N_11915,N_11526,N_11740);
nand U11916 (N_11916,N_11748,N_11698);
or U11917 (N_11917,N_11709,N_11657);
and U11918 (N_11918,N_11661,N_11514);
nor U11919 (N_11919,N_11544,N_11657);
or U11920 (N_11920,N_11744,N_11600);
xor U11921 (N_11921,N_11504,N_11709);
nor U11922 (N_11922,N_11542,N_11546);
and U11923 (N_11923,N_11550,N_11519);
or U11924 (N_11924,N_11509,N_11701);
nand U11925 (N_11925,N_11581,N_11627);
xnor U11926 (N_11926,N_11560,N_11655);
nand U11927 (N_11927,N_11658,N_11732);
and U11928 (N_11928,N_11643,N_11736);
and U11929 (N_11929,N_11741,N_11718);
and U11930 (N_11930,N_11737,N_11619);
or U11931 (N_11931,N_11699,N_11560);
nor U11932 (N_11932,N_11749,N_11705);
xor U11933 (N_11933,N_11585,N_11678);
and U11934 (N_11934,N_11636,N_11607);
nand U11935 (N_11935,N_11579,N_11703);
nand U11936 (N_11936,N_11716,N_11567);
and U11937 (N_11937,N_11723,N_11648);
nor U11938 (N_11938,N_11742,N_11636);
nand U11939 (N_11939,N_11647,N_11596);
and U11940 (N_11940,N_11528,N_11650);
or U11941 (N_11941,N_11644,N_11666);
xor U11942 (N_11942,N_11728,N_11720);
and U11943 (N_11943,N_11549,N_11643);
xnor U11944 (N_11944,N_11719,N_11621);
or U11945 (N_11945,N_11567,N_11592);
and U11946 (N_11946,N_11607,N_11649);
nand U11947 (N_11947,N_11536,N_11674);
nand U11948 (N_11948,N_11653,N_11633);
nor U11949 (N_11949,N_11501,N_11538);
or U11950 (N_11950,N_11522,N_11689);
xor U11951 (N_11951,N_11745,N_11687);
xor U11952 (N_11952,N_11728,N_11711);
xnor U11953 (N_11953,N_11716,N_11727);
and U11954 (N_11954,N_11538,N_11560);
and U11955 (N_11955,N_11708,N_11737);
and U11956 (N_11956,N_11693,N_11545);
nand U11957 (N_11957,N_11714,N_11710);
nor U11958 (N_11958,N_11716,N_11694);
or U11959 (N_11959,N_11746,N_11713);
nand U11960 (N_11960,N_11687,N_11631);
and U11961 (N_11961,N_11627,N_11533);
and U11962 (N_11962,N_11606,N_11749);
nor U11963 (N_11963,N_11571,N_11555);
nor U11964 (N_11964,N_11509,N_11612);
xor U11965 (N_11965,N_11721,N_11597);
or U11966 (N_11966,N_11514,N_11682);
nor U11967 (N_11967,N_11552,N_11637);
nand U11968 (N_11968,N_11503,N_11553);
nand U11969 (N_11969,N_11673,N_11551);
xnor U11970 (N_11970,N_11583,N_11573);
nand U11971 (N_11971,N_11729,N_11565);
and U11972 (N_11972,N_11640,N_11511);
or U11973 (N_11973,N_11688,N_11554);
nor U11974 (N_11974,N_11588,N_11511);
or U11975 (N_11975,N_11627,N_11543);
xnor U11976 (N_11976,N_11607,N_11554);
nor U11977 (N_11977,N_11690,N_11539);
xor U11978 (N_11978,N_11519,N_11685);
or U11979 (N_11979,N_11568,N_11682);
nand U11980 (N_11980,N_11522,N_11577);
nand U11981 (N_11981,N_11681,N_11553);
and U11982 (N_11982,N_11624,N_11590);
nor U11983 (N_11983,N_11504,N_11680);
nor U11984 (N_11984,N_11579,N_11560);
or U11985 (N_11985,N_11732,N_11727);
nand U11986 (N_11986,N_11627,N_11591);
and U11987 (N_11987,N_11575,N_11626);
xnor U11988 (N_11988,N_11693,N_11582);
and U11989 (N_11989,N_11693,N_11666);
xnor U11990 (N_11990,N_11717,N_11610);
nor U11991 (N_11991,N_11522,N_11583);
xor U11992 (N_11992,N_11660,N_11748);
xor U11993 (N_11993,N_11615,N_11677);
nand U11994 (N_11994,N_11611,N_11735);
nor U11995 (N_11995,N_11509,N_11613);
xor U11996 (N_11996,N_11565,N_11519);
or U11997 (N_11997,N_11748,N_11669);
nand U11998 (N_11998,N_11525,N_11642);
nand U11999 (N_11999,N_11720,N_11741);
nor U12000 (N_12000,N_11776,N_11873);
xor U12001 (N_12001,N_11866,N_11962);
nor U12002 (N_12002,N_11771,N_11763);
xor U12003 (N_12003,N_11770,N_11757);
xor U12004 (N_12004,N_11943,N_11826);
nor U12005 (N_12005,N_11912,N_11931);
xor U12006 (N_12006,N_11813,N_11819);
and U12007 (N_12007,N_11842,N_11977);
or U12008 (N_12008,N_11894,N_11801);
nand U12009 (N_12009,N_11955,N_11809);
or U12010 (N_12010,N_11818,N_11996);
xor U12011 (N_12011,N_11859,N_11998);
or U12012 (N_12012,N_11768,N_11885);
nor U12013 (N_12013,N_11803,N_11775);
nor U12014 (N_12014,N_11862,N_11880);
nand U12015 (N_12015,N_11877,N_11995);
or U12016 (N_12016,N_11758,N_11753);
nand U12017 (N_12017,N_11934,N_11805);
nand U12018 (N_12018,N_11889,N_11863);
and U12019 (N_12019,N_11944,N_11975);
xnor U12020 (N_12020,N_11825,N_11923);
xnor U12021 (N_12021,N_11917,N_11864);
nand U12022 (N_12022,N_11905,N_11856);
nor U12023 (N_12023,N_11807,N_11903);
or U12024 (N_12024,N_11848,N_11781);
or U12025 (N_12025,N_11844,N_11900);
nand U12026 (N_12026,N_11761,N_11953);
xor U12027 (N_12027,N_11854,N_11867);
nor U12028 (N_12028,N_11847,N_11790);
nor U12029 (N_12029,N_11766,N_11893);
nor U12030 (N_12030,N_11796,N_11780);
or U12031 (N_12031,N_11872,N_11891);
nand U12032 (N_12032,N_11840,N_11993);
xnor U12033 (N_12033,N_11817,N_11957);
nor U12034 (N_12034,N_11942,N_11828);
nor U12035 (N_12035,N_11846,N_11978);
or U12036 (N_12036,N_11956,N_11890);
nand U12037 (N_12037,N_11835,N_11952);
xnor U12038 (N_12038,N_11858,N_11986);
nor U12039 (N_12039,N_11969,N_11836);
or U12040 (N_12040,N_11999,N_11839);
nor U12041 (N_12041,N_11811,N_11950);
nand U12042 (N_12042,N_11800,N_11751);
nand U12043 (N_12043,N_11786,N_11970);
nor U12044 (N_12044,N_11794,N_11795);
nor U12045 (N_12045,N_11868,N_11982);
nand U12046 (N_12046,N_11849,N_11887);
nand U12047 (N_12047,N_11783,N_11935);
xnor U12048 (N_12048,N_11874,N_11870);
nor U12049 (N_12049,N_11876,N_11968);
and U12050 (N_12050,N_11997,N_11940);
or U12051 (N_12051,N_11991,N_11829);
or U12052 (N_12052,N_11762,N_11971);
xnor U12053 (N_12053,N_11861,N_11875);
or U12054 (N_12054,N_11960,N_11926);
nor U12055 (N_12055,N_11941,N_11901);
or U12056 (N_12056,N_11785,N_11949);
nor U12057 (N_12057,N_11884,N_11904);
xor U12058 (N_12058,N_11895,N_11908);
or U12059 (N_12059,N_11898,N_11979);
nor U12060 (N_12060,N_11888,N_11883);
xor U12061 (N_12061,N_11812,N_11920);
and U12062 (N_12062,N_11967,N_11922);
xor U12063 (N_12063,N_11911,N_11853);
nor U12064 (N_12064,N_11871,N_11851);
nand U12065 (N_12065,N_11906,N_11937);
xor U12066 (N_12066,N_11850,N_11981);
xor U12067 (N_12067,N_11965,N_11929);
xnor U12068 (N_12068,N_11769,N_11983);
nor U12069 (N_12069,N_11837,N_11928);
and U12070 (N_12070,N_11930,N_11966);
xnor U12071 (N_12071,N_11984,N_11860);
nand U12072 (N_12072,N_11834,N_11881);
nor U12073 (N_12073,N_11907,N_11841);
nor U12074 (N_12074,N_11852,N_11821);
nor U12075 (N_12075,N_11782,N_11961);
and U12076 (N_12076,N_11886,N_11985);
nor U12077 (N_12077,N_11815,N_11857);
nor U12078 (N_12078,N_11750,N_11914);
nand U12079 (N_12079,N_11987,N_11994);
nand U12080 (N_12080,N_11779,N_11838);
nand U12081 (N_12081,N_11820,N_11958);
and U12082 (N_12082,N_11963,N_11802);
nand U12083 (N_12083,N_11992,N_11772);
nor U12084 (N_12084,N_11973,N_11899);
nand U12085 (N_12085,N_11804,N_11869);
or U12086 (N_12086,N_11946,N_11927);
or U12087 (N_12087,N_11959,N_11787);
xnor U12088 (N_12088,N_11988,N_11916);
or U12089 (N_12089,N_11806,N_11948);
nor U12090 (N_12090,N_11831,N_11845);
nand U12091 (N_12091,N_11755,N_11990);
or U12092 (N_12092,N_11767,N_11756);
nor U12093 (N_12093,N_11760,N_11823);
and U12094 (N_12094,N_11824,N_11855);
nand U12095 (N_12095,N_11925,N_11915);
nor U12096 (N_12096,N_11936,N_11897);
nor U12097 (N_12097,N_11843,N_11777);
and U12098 (N_12098,N_11814,N_11788);
nor U12099 (N_12099,N_11933,N_11910);
and U12100 (N_12100,N_11919,N_11810);
xnor U12101 (N_12101,N_11798,N_11939);
nor U12102 (N_12102,N_11980,N_11951);
nor U12103 (N_12103,N_11865,N_11827);
or U12104 (N_12104,N_11879,N_11808);
xor U12105 (N_12105,N_11882,N_11833);
or U12106 (N_12106,N_11759,N_11792);
nor U12107 (N_12107,N_11902,N_11972);
xor U12108 (N_12108,N_11945,N_11764);
or U12109 (N_12109,N_11832,N_11896);
xor U12110 (N_12110,N_11752,N_11892);
nor U12111 (N_12111,N_11964,N_11947);
and U12112 (N_12112,N_11932,N_11822);
or U12113 (N_12113,N_11954,N_11989);
or U12114 (N_12114,N_11974,N_11765);
xnor U12115 (N_12115,N_11784,N_11913);
nand U12116 (N_12116,N_11789,N_11921);
xor U12117 (N_12117,N_11938,N_11924);
or U12118 (N_12118,N_11816,N_11976);
or U12119 (N_12119,N_11791,N_11793);
and U12120 (N_12120,N_11754,N_11830);
and U12121 (N_12121,N_11797,N_11773);
nor U12122 (N_12122,N_11799,N_11909);
or U12123 (N_12123,N_11778,N_11918);
xnor U12124 (N_12124,N_11878,N_11774);
nor U12125 (N_12125,N_11969,N_11990);
nor U12126 (N_12126,N_11885,N_11924);
or U12127 (N_12127,N_11841,N_11979);
or U12128 (N_12128,N_11952,N_11792);
xor U12129 (N_12129,N_11784,N_11891);
or U12130 (N_12130,N_11799,N_11856);
nor U12131 (N_12131,N_11860,N_11934);
or U12132 (N_12132,N_11801,N_11843);
nor U12133 (N_12133,N_11977,N_11953);
xor U12134 (N_12134,N_11937,N_11835);
nand U12135 (N_12135,N_11773,N_11976);
nand U12136 (N_12136,N_11914,N_11815);
nand U12137 (N_12137,N_11840,N_11863);
nor U12138 (N_12138,N_11896,N_11943);
and U12139 (N_12139,N_11897,N_11929);
xor U12140 (N_12140,N_11993,N_11878);
or U12141 (N_12141,N_11906,N_11889);
nand U12142 (N_12142,N_11803,N_11982);
or U12143 (N_12143,N_11766,N_11954);
xor U12144 (N_12144,N_11894,N_11762);
nand U12145 (N_12145,N_11914,N_11978);
or U12146 (N_12146,N_11875,N_11977);
or U12147 (N_12147,N_11935,N_11943);
nand U12148 (N_12148,N_11830,N_11945);
nand U12149 (N_12149,N_11852,N_11835);
xnor U12150 (N_12150,N_11886,N_11846);
and U12151 (N_12151,N_11898,N_11992);
and U12152 (N_12152,N_11916,N_11943);
nor U12153 (N_12153,N_11916,N_11904);
nor U12154 (N_12154,N_11792,N_11995);
and U12155 (N_12155,N_11944,N_11818);
and U12156 (N_12156,N_11968,N_11939);
nor U12157 (N_12157,N_11912,N_11795);
nor U12158 (N_12158,N_11913,N_11802);
nor U12159 (N_12159,N_11943,N_11824);
xor U12160 (N_12160,N_11945,N_11906);
xnor U12161 (N_12161,N_11887,N_11802);
xnor U12162 (N_12162,N_11853,N_11875);
nor U12163 (N_12163,N_11944,N_11817);
xor U12164 (N_12164,N_11847,N_11838);
or U12165 (N_12165,N_11857,N_11961);
nand U12166 (N_12166,N_11993,N_11839);
and U12167 (N_12167,N_11953,N_11836);
xnor U12168 (N_12168,N_11931,N_11908);
and U12169 (N_12169,N_11988,N_11799);
nor U12170 (N_12170,N_11991,N_11763);
or U12171 (N_12171,N_11798,N_11946);
and U12172 (N_12172,N_11836,N_11856);
or U12173 (N_12173,N_11984,N_11883);
nand U12174 (N_12174,N_11969,N_11826);
xnor U12175 (N_12175,N_11831,N_11805);
nor U12176 (N_12176,N_11873,N_11979);
and U12177 (N_12177,N_11958,N_11796);
nand U12178 (N_12178,N_11768,N_11794);
nand U12179 (N_12179,N_11891,N_11762);
nand U12180 (N_12180,N_11774,N_11779);
xnor U12181 (N_12181,N_11941,N_11851);
and U12182 (N_12182,N_11853,N_11840);
and U12183 (N_12183,N_11960,N_11759);
xor U12184 (N_12184,N_11823,N_11839);
xor U12185 (N_12185,N_11752,N_11952);
and U12186 (N_12186,N_11922,N_11915);
nor U12187 (N_12187,N_11998,N_11793);
xor U12188 (N_12188,N_11995,N_11814);
nand U12189 (N_12189,N_11850,N_11998);
or U12190 (N_12190,N_11947,N_11806);
nand U12191 (N_12191,N_11772,N_11874);
nand U12192 (N_12192,N_11971,N_11805);
and U12193 (N_12193,N_11828,N_11799);
nand U12194 (N_12194,N_11845,N_11755);
or U12195 (N_12195,N_11762,N_11789);
and U12196 (N_12196,N_11789,N_11969);
nand U12197 (N_12197,N_11943,N_11754);
or U12198 (N_12198,N_11782,N_11945);
or U12199 (N_12199,N_11994,N_11951);
and U12200 (N_12200,N_11828,N_11975);
nor U12201 (N_12201,N_11844,N_11877);
or U12202 (N_12202,N_11885,N_11954);
nand U12203 (N_12203,N_11935,N_11759);
and U12204 (N_12204,N_11883,N_11776);
xor U12205 (N_12205,N_11898,N_11983);
nand U12206 (N_12206,N_11794,N_11992);
nor U12207 (N_12207,N_11927,N_11789);
nor U12208 (N_12208,N_11921,N_11814);
and U12209 (N_12209,N_11811,N_11995);
nand U12210 (N_12210,N_11925,N_11968);
and U12211 (N_12211,N_11908,N_11758);
nand U12212 (N_12212,N_11954,N_11975);
xor U12213 (N_12213,N_11820,N_11999);
or U12214 (N_12214,N_11808,N_11892);
xnor U12215 (N_12215,N_11916,N_11933);
or U12216 (N_12216,N_11845,N_11820);
or U12217 (N_12217,N_11812,N_11918);
or U12218 (N_12218,N_11986,N_11769);
xnor U12219 (N_12219,N_11974,N_11862);
or U12220 (N_12220,N_11754,N_11880);
nand U12221 (N_12221,N_11993,N_11851);
xor U12222 (N_12222,N_11825,N_11800);
or U12223 (N_12223,N_11795,N_11979);
or U12224 (N_12224,N_11915,N_11865);
nor U12225 (N_12225,N_11774,N_11867);
or U12226 (N_12226,N_11792,N_11870);
nand U12227 (N_12227,N_11914,N_11880);
nand U12228 (N_12228,N_11824,N_11947);
nor U12229 (N_12229,N_11927,N_11910);
and U12230 (N_12230,N_11934,N_11782);
and U12231 (N_12231,N_11864,N_11846);
xor U12232 (N_12232,N_11812,N_11786);
nand U12233 (N_12233,N_11762,N_11857);
xor U12234 (N_12234,N_11898,N_11753);
nand U12235 (N_12235,N_11780,N_11911);
nor U12236 (N_12236,N_11754,N_11774);
xor U12237 (N_12237,N_11831,N_11769);
nand U12238 (N_12238,N_11763,N_11923);
or U12239 (N_12239,N_11760,N_11886);
xor U12240 (N_12240,N_11998,N_11821);
and U12241 (N_12241,N_11751,N_11778);
nand U12242 (N_12242,N_11848,N_11807);
or U12243 (N_12243,N_11882,N_11946);
nand U12244 (N_12244,N_11877,N_11750);
nor U12245 (N_12245,N_11980,N_11777);
xor U12246 (N_12246,N_11995,N_11886);
or U12247 (N_12247,N_11981,N_11823);
xor U12248 (N_12248,N_11879,N_11790);
nand U12249 (N_12249,N_11916,N_11761);
nor U12250 (N_12250,N_12091,N_12003);
nand U12251 (N_12251,N_12238,N_12190);
and U12252 (N_12252,N_12147,N_12048);
or U12253 (N_12253,N_12224,N_12028);
nor U12254 (N_12254,N_12000,N_12053);
or U12255 (N_12255,N_12121,N_12183);
or U12256 (N_12256,N_12089,N_12115);
xor U12257 (N_12257,N_12150,N_12067);
xor U12258 (N_12258,N_12239,N_12002);
nand U12259 (N_12259,N_12023,N_12022);
nand U12260 (N_12260,N_12018,N_12200);
nand U12261 (N_12261,N_12029,N_12016);
xnor U12262 (N_12262,N_12164,N_12216);
and U12263 (N_12263,N_12045,N_12013);
or U12264 (N_12264,N_12055,N_12214);
nand U12265 (N_12265,N_12155,N_12123);
and U12266 (N_12266,N_12176,N_12059);
nand U12267 (N_12267,N_12163,N_12170);
and U12268 (N_12268,N_12187,N_12156);
nand U12269 (N_12269,N_12021,N_12161);
nand U12270 (N_12270,N_12052,N_12241);
nand U12271 (N_12271,N_12042,N_12116);
and U12272 (N_12272,N_12202,N_12084);
or U12273 (N_12273,N_12014,N_12112);
or U12274 (N_12274,N_12092,N_12087);
or U12275 (N_12275,N_12093,N_12247);
xor U12276 (N_12276,N_12127,N_12001);
or U12277 (N_12277,N_12213,N_12064);
nor U12278 (N_12278,N_12026,N_12151);
xor U12279 (N_12279,N_12160,N_12005);
nand U12280 (N_12280,N_12038,N_12119);
or U12281 (N_12281,N_12143,N_12065);
or U12282 (N_12282,N_12074,N_12061);
and U12283 (N_12283,N_12148,N_12072);
nor U12284 (N_12284,N_12110,N_12204);
or U12285 (N_12285,N_12228,N_12129);
xor U12286 (N_12286,N_12144,N_12120);
xnor U12287 (N_12287,N_12167,N_12025);
nor U12288 (N_12288,N_12237,N_12236);
and U12289 (N_12289,N_12106,N_12232);
and U12290 (N_12290,N_12073,N_12166);
nand U12291 (N_12291,N_12139,N_12173);
xnor U12292 (N_12292,N_12113,N_12231);
xnor U12293 (N_12293,N_12015,N_12230);
nand U12294 (N_12294,N_12149,N_12062);
and U12295 (N_12295,N_12128,N_12098);
nand U12296 (N_12296,N_12162,N_12208);
nor U12297 (N_12297,N_12101,N_12180);
nor U12298 (N_12298,N_12184,N_12096);
xnor U12299 (N_12299,N_12192,N_12117);
or U12300 (N_12300,N_12217,N_12068);
xor U12301 (N_12301,N_12248,N_12218);
nor U12302 (N_12302,N_12194,N_12080);
and U12303 (N_12303,N_12070,N_12057);
and U12304 (N_12304,N_12032,N_12234);
nand U12305 (N_12305,N_12078,N_12165);
nand U12306 (N_12306,N_12246,N_12227);
nor U12307 (N_12307,N_12069,N_12186);
xor U12308 (N_12308,N_12036,N_12223);
xor U12309 (N_12309,N_12040,N_12229);
or U12310 (N_12310,N_12024,N_12125);
xnor U12311 (N_12311,N_12108,N_12090);
or U12312 (N_12312,N_12138,N_12196);
or U12313 (N_12313,N_12221,N_12034);
and U12314 (N_12314,N_12066,N_12046);
xnor U12315 (N_12315,N_12235,N_12142);
xor U12316 (N_12316,N_12243,N_12136);
nor U12317 (N_12317,N_12118,N_12222);
xnor U12318 (N_12318,N_12153,N_12010);
and U12319 (N_12319,N_12175,N_12104);
nor U12320 (N_12320,N_12076,N_12085);
xor U12321 (N_12321,N_12158,N_12178);
and U12322 (N_12322,N_12111,N_12205);
xor U12323 (N_12323,N_12134,N_12097);
xnor U12324 (N_12324,N_12033,N_12191);
nand U12325 (N_12325,N_12009,N_12159);
or U12326 (N_12326,N_12242,N_12049);
or U12327 (N_12327,N_12219,N_12198);
nand U12328 (N_12328,N_12177,N_12195);
and U12329 (N_12329,N_12203,N_12006);
nor U12330 (N_12330,N_12051,N_12233);
nor U12331 (N_12331,N_12041,N_12100);
and U12332 (N_12332,N_12210,N_12133);
xnor U12333 (N_12333,N_12109,N_12044);
nor U12334 (N_12334,N_12030,N_12249);
xor U12335 (N_12335,N_12193,N_12172);
or U12336 (N_12336,N_12019,N_12215);
xor U12337 (N_12337,N_12012,N_12095);
and U12338 (N_12338,N_12075,N_12056);
nand U12339 (N_12339,N_12082,N_12154);
nand U12340 (N_12340,N_12169,N_12152);
nor U12341 (N_12341,N_12037,N_12088);
xnor U12342 (N_12342,N_12102,N_12181);
nor U12343 (N_12343,N_12114,N_12188);
and U12344 (N_12344,N_12131,N_12086);
or U12345 (N_12345,N_12043,N_12124);
xor U12346 (N_12346,N_12206,N_12058);
xor U12347 (N_12347,N_12212,N_12081);
nand U12348 (N_12348,N_12211,N_12107);
or U12349 (N_12349,N_12050,N_12197);
xnor U12350 (N_12350,N_12105,N_12199);
nor U12351 (N_12351,N_12027,N_12054);
or U12352 (N_12352,N_12244,N_12225);
nand U12353 (N_12353,N_12245,N_12035);
nor U12354 (N_12354,N_12007,N_12189);
nor U12355 (N_12355,N_12132,N_12174);
or U12356 (N_12356,N_12240,N_12226);
xnor U12357 (N_12357,N_12071,N_12039);
or U12358 (N_12358,N_12135,N_12145);
nand U12359 (N_12359,N_12182,N_12141);
nand U12360 (N_12360,N_12122,N_12063);
and U12361 (N_12361,N_12004,N_12094);
or U12362 (N_12362,N_12103,N_12171);
nand U12363 (N_12363,N_12130,N_12126);
or U12364 (N_12364,N_12220,N_12031);
and U12365 (N_12365,N_12146,N_12168);
or U12366 (N_12366,N_12047,N_12185);
nor U12367 (N_12367,N_12209,N_12060);
and U12368 (N_12368,N_12207,N_12077);
nor U12369 (N_12369,N_12008,N_12011);
or U12370 (N_12370,N_12017,N_12099);
nand U12371 (N_12371,N_12137,N_12020);
and U12372 (N_12372,N_12083,N_12157);
or U12373 (N_12373,N_12179,N_12201);
nand U12374 (N_12374,N_12140,N_12079);
or U12375 (N_12375,N_12049,N_12187);
nand U12376 (N_12376,N_12023,N_12041);
xor U12377 (N_12377,N_12224,N_12236);
nand U12378 (N_12378,N_12097,N_12016);
or U12379 (N_12379,N_12116,N_12064);
and U12380 (N_12380,N_12133,N_12017);
or U12381 (N_12381,N_12204,N_12230);
nand U12382 (N_12382,N_12048,N_12130);
nand U12383 (N_12383,N_12129,N_12010);
xor U12384 (N_12384,N_12012,N_12228);
nor U12385 (N_12385,N_12094,N_12021);
or U12386 (N_12386,N_12047,N_12142);
nand U12387 (N_12387,N_12129,N_12122);
nand U12388 (N_12388,N_12156,N_12076);
nor U12389 (N_12389,N_12197,N_12032);
or U12390 (N_12390,N_12206,N_12123);
or U12391 (N_12391,N_12053,N_12221);
and U12392 (N_12392,N_12058,N_12147);
nand U12393 (N_12393,N_12097,N_12064);
xor U12394 (N_12394,N_12132,N_12093);
xnor U12395 (N_12395,N_12207,N_12182);
nor U12396 (N_12396,N_12128,N_12243);
xor U12397 (N_12397,N_12079,N_12073);
nand U12398 (N_12398,N_12131,N_12216);
or U12399 (N_12399,N_12097,N_12248);
and U12400 (N_12400,N_12098,N_12214);
and U12401 (N_12401,N_12078,N_12096);
and U12402 (N_12402,N_12118,N_12072);
and U12403 (N_12403,N_12147,N_12243);
nor U12404 (N_12404,N_12079,N_12180);
nand U12405 (N_12405,N_12194,N_12051);
nor U12406 (N_12406,N_12159,N_12093);
nand U12407 (N_12407,N_12087,N_12198);
and U12408 (N_12408,N_12198,N_12243);
xnor U12409 (N_12409,N_12147,N_12036);
nand U12410 (N_12410,N_12195,N_12156);
xnor U12411 (N_12411,N_12178,N_12085);
xor U12412 (N_12412,N_12187,N_12172);
and U12413 (N_12413,N_12070,N_12205);
or U12414 (N_12414,N_12082,N_12052);
nand U12415 (N_12415,N_12028,N_12125);
or U12416 (N_12416,N_12200,N_12064);
nor U12417 (N_12417,N_12009,N_12123);
nor U12418 (N_12418,N_12099,N_12061);
nand U12419 (N_12419,N_12047,N_12062);
nand U12420 (N_12420,N_12244,N_12246);
nor U12421 (N_12421,N_12162,N_12136);
nand U12422 (N_12422,N_12189,N_12030);
nor U12423 (N_12423,N_12127,N_12100);
nand U12424 (N_12424,N_12041,N_12204);
xor U12425 (N_12425,N_12084,N_12075);
nor U12426 (N_12426,N_12082,N_12053);
xor U12427 (N_12427,N_12119,N_12237);
xor U12428 (N_12428,N_12073,N_12153);
nor U12429 (N_12429,N_12076,N_12153);
nor U12430 (N_12430,N_12215,N_12234);
and U12431 (N_12431,N_12080,N_12021);
nor U12432 (N_12432,N_12102,N_12070);
or U12433 (N_12433,N_12200,N_12096);
nand U12434 (N_12434,N_12045,N_12157);
nand U12435 (N_12435,N_12169,N_12091);
and U12436 (N_12436,N_12130,N_12120);
xor U12437 (N_12437,N_12056,N_12243);
or U12438 (N_12438,N_12032,N_12164);
nor U12439 (N_12439,N_12228,N_12105);
or U12440 (N_12440,N_12235,N_12132);
nand U12441 (N_12441,N_12220,N_12051);
or U12442 (N_12442,N_12089,N_12170);
or U12443 (N_12443,N_12201,N_12146);
or U12444 (N_12444,N_12061,N_12100);
nand U12445 (N_12445,N_12182,N_12161);
xnor U12446 (N_12446,N_12023,N_12190);
or U12447 (N_12447,N_12102,N_12031);
and U12448 (N_12448,N_12012,N_12009);
or U12449 (N_12449,N_12120,N_12088);
and U12450 (N_12450,N_12195,N_12148);
nor U12451 (N_12451,N_12018,N_12117);
or U12452 (N_12452,N_12216,N_12018);
nand U12453 (N_12453,N_12101,N_12104);
xnor U12454 (N_12454,N_12027,N_12076);
and U12455 (N_12455,N_12236,N_12027);
or U12456 (N_12456,N_12209,N_12128);
xnor U12457 (N_12457,N_12058,N_12149);
xnor U12458 (N_12458,N_12179,N_12219);
nand U12459 (N_12459,N_12196,N_12063);
or U12460 (N_12460,N_12058,N_12057);
xnor U12461 (N_12461,N_12073,N_12185);
xor U12462 (N_12462,N_12208,N_12064);
nor U12463 (N_12463,N_12074,N_12037);
and U12464 (N_12464,N_12230,N_12196);
nor U12465 (N_12465,N_12237,N_12123);
nand U12466 (N_12466,N_12174,N_12234);
and U12467 (N_12467,N_12174,N_12165);
xnor U12468 (N_12468,N_12013,N_12160);
xor U12469 (N_12469,N_12041,N_12171);
nand U12470 (N_12470,N_12098,N_12245);
nor U12471 (N_12471,N_12140,N_12108);
xnor U12472 (N_12472,N_12085,N_12237);
xnor U12473 (N_12473,N_12231,N_12123);
or U12474 (N_12474,N_12217,N_12130);
or U12475 (N_12475,N_12096,N_12230);
or U12476 (N_12476,N_12123,N_12165);
or U12477 (N_12477,N_12231,N_12117);
nand U12478 (N_12478,N_12238,N_12221);
or U12479 (N_12479,N_12235,N_12204);
and U12480 (N_12480,N_12093,N_12092);
xor U12481 (N_12481,N_12051,N_12008);
nand U12482 (N_12482,N_12194,N_12104);
and U12483 (N_12483,N_12034,N_12017);
or U12484 (N_12484,N_12248,N_12104);
nand U12485 (N_12485,N_12229,N_12087);
and U12486 (N_12486,N_12104,N_12070);
or U12487 (N_12487,N_12116,N_12225);
or U12488 (N_12488,N_12073,N_12000);
nand U12489 (N_12489,N_12207,N_12060);
xor U12490 (N_12490,N_12248,N_12040);
xor U12491 (N_12491,N_12022,N_12089);
or U12492 (N_12492,N_12122,N_12194);
or U12493 (N_12493,N_12199,N_12235);
and U12494 (N_12494,N_12045,N_12069);
xor U12495 (N_12495,N_12172,N_12221);
nand U12496 (N_12496,N_12035,N_12106);
or U12497 (N_12497,N_12112,N_12051);
nand U12498 (N_12498,N_12210,N_12075);
and U12499 (N_12499,N_12006,N_12246);
nor U12500 (N_12500,N_12286,N_12478);
nor U12501 (N_12501,N_12393,N_12490);
xnor U12502 (N_12502,N_12333,N_12385);
xor U12503 (N_12503,N_12399,N_12284);
and U12504 (N_12504,N_12459,N_12384);
nand U12505 (N_12505,N_12252,N_12376);
xor U12506 (N_12506,N_12398,N_12499);
xor U12507 (N_12507,N_12288,N_12415);
nor U12508 (N_12508,N_12268,N_12367);
nand U12509 (N_12509,N_12479,N_12368);
nand U12510 (N_12510,N_12295,N_12339);
and U12511 (N_12511,N_12451,N_12462);
nand U12512 (N_12512,N_12424,N_12299);
nor U12513 (N_12513,N_12388,N_12470);
xor U12514 (N_12514,N_12400,N_12441);
and U12515 (N_12515,N_12468,N_12342);
nor U12516 (N_12516,N_12392,N_12485);
or U12517 (N_12517,N_12366,N_12317);
nand U12518 (N_12518,N_12464,N_12395);
xnor U12519 (N_12519,N_12403,N_12313);
or U12520 (N_12520,N_12463,N_12316);
and U12521 (N_12521,N_12251,N_12359);
nand U12522 (N_12522,N_12259,N_12473);
and U12523 (N_12523,N_12417,N_12484);
or U12524 (N_12524,N_12477,N_12454);
or U12525 (N_12525,N_12364,N_12496);
nand U12526 (N_12526,N_12371,N_12282);
nor U12527 (N_12527,N_12419,N_12353);
or U12528 (N_12528,N_12446,N_12324);
and U12529 (N_12529,N_12455,N_12370);
and U12530 (N_12530,N_12476,N_12276);
nor U12531 (N_12531,N_12264,N_12332);
or U12532 (N_12532,N_12495,N_12378);
nor U12533 (N_12533,N_12326,N_12278);
and U12534 (N_12534,N_12412,N_12297);
xor U12535 (N_12535,N_12414,N_12443);
xor U12536 (N_12536,N_12408,N_12287);
or U12537 (N_12537,N_12480,N_12271);
and U12538 (N_12538,N_12449,N_12289);
and U12539 (N_12539,N_12290,N_12380);
and U12540 (N_12540,N_12323,N_12272);
nor U12541 (N_12541,N_12291,N_12306);
nand U12542 (N_12542,N_12281,N_12255);
nand U12543 (N_12543,N_12337,N_12314);
xnor U12544 (N_12544,N_12283,N_12302);
nor U12545 (N_12545,N_12347,N_12257);
xnor U12546 (N_12546,N_12475,N_12487);
nand U12547 (N_12547,N_12350,N_12433);
or U12548 (N_12548,N_12311,N_12394);
and U12549 (N_12549,N_12429,N_12354);
xor U12550 (N_12550,N_12352,N_12423);
nor U12551 (N_12551,N_12386,N_12457);
or U12552 (N_12552,N_12253,N_12439);
nor U12553 (N_12553,N_12325,N_12355);
nor U12554 (N_12554,N_12292,N_12497);
and U12555 (N_12555,N_12312,N_12461);
xnor U12556 (N_12556,N_12488,N_12307);
nor U12557 (N_12557,N_12327,N_12343);
nand U12558 (N_12558,N_12374,N_12447);
xnor U12559 (N_12559,N_12465,N_12258);
xnor U12560 (N_12560,N_12358,N_12407);
and U12561 (N_12561,N_12469,N_12310);
or U12562 (N_12562,N_12472,N_12425);
nand U12563 (N_12563,N_12466,N_12340);
xnor U12564 (N_12564,N_12309,N_12360);
and U12565 (N_12565,N_12390,N_12345);
or U12566 (N_12566,N_12491,N_12349);
or U12567 (N_12567,N_12260,N_12351);
and U12568 (N_12568,N_12361,N_12494);
nor U12569 (N_12569,N_12274,N_12492);
nand U12570 (N_12570,N_12438,N_12334);
nand U12571 (N_12571,N_12305,N_12256);
or U12572 (N_12572,N_12450,N_12448);
nand U12573 (N_12573,N_12250,N_12432);
or U12574 (N_12574,N_12382,N_12319);
or U12575 (N_12575,N_12406,N_12320);
nor U12576 (N_12576,N_12372,N_12262);
and U12577 (N_12577,N_12265,N_12318);
nand U12578 (N_12578,N_12445,N_12338);
nand U12579 (N_12579,N_12263,N_12254);
xnor U12580 (N_12580,N_12467,N_12402);
nor U12581 (N_12581,N_12270,N_12301);
and U12582 (N_12582,N_12267,N_12421);
and U12583 (N_12583,N_12346,N_12269);
nand U12584 (N_12584,N_12315,N_12296);
or U12585 (N_12585,N_12357,N_12391);
nand U12586 (N_12586,N_12280,N_12308);
and U12587 (N_12587,N_12452,N_12275);
or U12588 (N_12588,N_12303,N_12277);
nand U12589 (N_12589,N_12434,N_12498);
nor U12590 (N_12590,N_12413,N_12397);
and U12591 (N_12591,N_12437,N_12293);
nand U12592 (N_12592,N_12389,N_12428);
or U12593 (N_12593,N_12369,N_12365);
or U12594 (N_12594,N_12362,N_12440);
and U12595 (N_12595,N_12427,N_12481);
or U12596 (N_12596,N_12294,N_12273);
nand U12597 (N_12597,N_12336,N_12279);
and U12598 (N_12598,N_12266,N_12411);
xnor U12599 (N_12599,N_12404,N_12416);
nand U12600 (N_12600,N_12330,N_12379);
nor U12601 (N_12601,N_12341,N_12298);
and U12602 (N_12602,N_12456,N_12261);
nand U12603 (N_12603,N_12442,N_12285);
nor U12604 (N_12604,N_12483,N_12344);
nand U12605 (N_12605,N_12486,N_12410);
nor U12606 (N_12606,N_12348,N_12363);
nor U12607 (N_12607,N_12375,N_12460);
or U12608 (N_12608,N_12482,N_12471);
xnor U12609 (N_12609,N_12381,N_12458);
xor U12610 (N_12610,N_12444,N_12489);
nand U12611 (N_12611,N_12418,N_12328);
nor U12612 (N_12612,N_12383,N_12453);
and U12613 (N_12613,N_12356,N_12331);
and U12614 (N_12614,N_12430,N_12300);
nor U12615 (N_12615,N_12321,N_12377);
or U12616 (N_12616,N_12387,N_12322);
nand U12617 (N_12617,N_12401,N_12409);
nand U12618 (N_12618,N_12435,N_12304);
nand U12619 (N_12619,N_12474,N_12405);
or U12620 (N_12620,N_12329,N_12426);
and U12621 (N_12621,N_12396,N_12335);
xor U12622 (N_12622,N_12436,N_12431);
nor U12623 (N_12623,N_12420,N_12373);
or U12624 (N_12624,N_12422,N_12493);
and U12625 (N_12625,N_12318,N_12282);
or U12626 (N_12626,N_12263,N_12346);
and U12627 (N_12627,N_12308,N_12452);
nor U12628 (N_12628,N_12431,N_12368);
or U12629 (N_12629,N_12263,N_12407);
and U12630 (N_12630,N_12343,N_12271);
nand U12631 (N_12631,N_12268,N_12250);
nor U12632 (N_12632,N_12469,N_12485);
nor U12633 (N_12633,N_12281,N_12494);
nor U12634 (N_12634,N_12354,N_12299);
nor U12635 (N_12635,N_12464,N_12317);
xnor U12636 (N_12636,N_12377,N_12329);
or U12637 (N_12637,N_12430,N_12356);
nand U12638 (N_12638,N_12477,N_12466);
nand U12639 (N_12639,N_12312,N_12327);
or U12640 (N_12640,N_12359,N_12476);
or U12641 (N_12641,N_12483,N_12414);
and U12642 (N_12642,N_12314,N_12431);
nand U12643 (N_12643,N_12324,N_12309);
or U12644 (N_12644,N_12385,N_12349);
xor U12645 (N_12645,N_12404,N_12347);
nor U12646 (N_12646,N_12448,N_12364);
and U12647 (N_12647,N_12369,N_12344);
or U12648 (N_12648,N_12420,N_12486);
nor U12649 (N_12649,N_12282,N_12485);
and U12650 (N_12650,N_12434,N_12396);
nor U12651 (N_12651,N_12424,N_12417);
xnor U12652 (N_12652,N_12274,N_12406);
nor U12653 (N_12653,N_12319,N_12341);
and U12654 (N_12654,N_12342,N_12412);
nor U12655 (N_12655,N_12483,N_12443);
nand U12656 (N_12656,N_12412,N_12321);
and U12657 (N_12657,N_12484,N_12258);
and U12658 (N_12658,N_12266,N_12386);
nor U12659 (N_12659,N_12275,N_12397);
xnor U12660 (N_12660,N_12366,N_12255);
nor U12661 (N_12661,N_12289,N_12384);
and U12662 (N_12662,N_12282,N_12302);
and U12663 (N_12663,N_12409,N_12370);
nor U12664 (N_12664,N_12268,N_12320);
or U12665 (N_12665,N_12325,N_12388);
nand U12666 (N_12666,N_12331,N_12493);
or U12667 (N_12667,N_12279,N_12496);
or U12668 (N_12668,N_12381,N_12471);
nand U12669 (N_12669,N_12301,N_12496);
or U12670 (N_12670,N_12349,N_12321);
nand U12671 (N_12671,N_12362,N_12418);
xor U12672 (N_12672,N_12358,N_12313);
and U12673 (N_12673,N_12432,N_12460);
and U12674 (N_12674,N_12374,N_12484);
or U12675 (N_12675,N_12468,N_12304);
nand U12676 (N_12676,N_12256,N_12321);
or U12677 (N_12677,N_12331,N_12409);
nor U12678 (N_12678,N_12295,N_12425);
xnor U12679 (N_12679,N_12471,N_12441);
and U12680 (N_12680,N_12283,N_12487);
nor U12681 (N_12681,N_12491,N_12417);
or U12682 (N_12682,N_12378,N_12272);
nand U12683 (N_12683,N_12415,N_12346);
or U12684 (N_12684,N_12407,N_12456);
nor U12685 (N_12685,N_12275,N_12430);
xnor U12686 (N_12686,N_12351,N_12470);
nor U12687 (N_12687,N_12429,N_12409);
nor U12688 (N_12688,N_12300,N_12325);
nand U12689 (N_12689,N_12262,N_12472);
xor U12690 (N_12690,N_12318,N_12385);
nand U12691 (N_12691,N_12395,N_12471);
xnor U12692 (N_12692,N_12359,N_12294);
nand U12693 (N_12693,N_12260,N_12432);
nor U12694 (N_12694,N_12258,N_12471);
nor U12695 (N_12695,N_12394,N_12425);
and U12696 (N_12696,N_12418,N_12375);
nand U12697 (N_12697,N_12468,N_12264);
nor U12698 (N_12698,N_12297,N_12421);
nand U12699 (N_12699,N_12345,N_12321);
nand U12700 (N_12700,N_12493,N_12421);
xor U12701 (N_12701,N_12485,N_12268);
or U12702 (N_12702,N_12294,N_12384);
or U12703 (N_12703,N_12478,N_12262);
nor U12704 (N_12704,N_12456,N_12350);
nor U12705 (N_12705,N_12418,N_12434);
xnor U12706 (N_12706,N_12333,N_12302);
or U12707 (N_12707,N_12303,N_12272);
xor U12708 (N_12708,N_12400,N_12312);
and U12709 (N_12709,N_12377,N_12395);
nor U12710 (N_12710,N_12471,N_12385);
or U12711 (N_12711,N_12386,N_12419);
or U12712 (N_12712,N_12461,N_12491);
and U12713 (N_12713,N_12291,N_12483);
or U12714 (N_12714,N_12299,N_12437);
and U12715 (N_12715,N_12268,N_12417);
nand U12716 (N_12716,N_12483,N_12250);
nand U12717 (N_12717,N_12492,N_12438);
or U12718 (N_12718,N_12420,N_12349);
xor U12719 (N_12719,N_12423,N_12453);
xor U12720 (N_12720,N_12444,N_12319);
or U12721 (N_12721,N_12417,N_12498);
and U12722 (N_12722,N_12322,N_12427);
and U12723 (N_12723,N_12303,N_12300);
or U12724 (N_12724,N_12294,N_12391);
nand U12725 (N_12725,N_12267,N_12253);
nand U12726 (N_12726,N_12349,N_12378);
and U12727 (N_12727,N_12413,N_12401);
or U12728 (N_12728,N_12360,N_12359);
and U12729 (N_12729,N_12473,N_12433);
nor U12730 (N_12730,N_12488,N_12303);
and U12731 (N_12731,N_12362,N_12459);
or U12732 (N_12732,N_12410,N_12293);
xnor U12733 (N_12733,N_12495,N_12274);
nand U12734 (N_12734,N_12418,N_12289);
or U12735 (N_12735,N_12316,N_12446);
or U12736 (N_12736,N_12341,N_12327);
xor U12737 (N_12737,N_12428,N_12286);
nor U12738 (N_12738,N_12301,N_12394);
nor U12739 (N_12739,N_12392,N_12422);
and U12740 (N_12740,N_12353,N_12378);
nand U12741 (N_12741,N_12257,N_12317);
and U12742 (N_12742,N_12327,N_12305);
nand U12743 (N_12743,N_12319,N_12388);
nand U12744 (N_12744,N_12354,N_12379);
nand U12745 (N_12745,N_12410,N_12471);
nand U12746 (N_12746,N_12430,N_12413);
and U12747 (N_12747,N_12414,N_12418);
xnor U12748 (N_12748,N_12330,N_12262);
and U12749 (N_12749,N_12458,N_12384);
nand U12750 (N_12750,N_12680,N_12558);
nand U12751 (N_12751,N_12728,N_12557);
nor U12752 (N_12752,N_12582,N_12565);
xor U12753 (N_12753,N_12539,N_12605);
and U12754 (N_12754,N_12516,N_12703);
and U12755 (N_12755,N_12650,N_12567);
nand U12756 (N_12756,N_12690,N_12723);
nand U12757 (N_12757,N_12736,N_12664);
and U12758 (N_12758,N_12523,N_12684);
and U12759 (N_12759,N_12720,N_12520);
nor U12760 (N_12760,N_12503,N_12697);
nand U12761 (N_12761,N_12578,N_12666);
and U12762 (N_12762,N_12575,N_12584);
nor U12763 (N_12763,N_12544,N_12733);
nor U12764 (N_12764,N_12505,N_12502);
and U12765 (N_12765,N_12564,N_12695);
xor U12766 (N_12766,N_12670,N_12726);
or U12767 (N_12767,N_12563,N_12541);
or U12768 (N_12768,N_12731,N_12708);
xnor U12769 (N_12769,N_12629,N_12514);
and U12770 (N_12770,N_12644,N_12626);
and U12771 (N_12771,N_12643,N_12727);
nor U12772 (N_12772,N_12694,N_12685);
or U12773 (N_12773,N_12509,N_12618);
xnor U12774 (N_12774,N_12746,N_12531);
and U12775 (N_12775,N_12621,N_12552);
and U12776 (N_12776,N_12663,N_12589);
or U12777 (N_12777,N_12638,N_12637);
and U12778 (N_12778,N_12607,N_12594);
or U12779 (N_12779,N_12586,N_12702);
nand U12780 (N_12780,N_12732,N_12507);
and U12781 (N_12781,N_12616,N_12554);
nor U12782 (N_12782,N_12660,N_12566);
or U12783 (N_12783,N_12742,N_12500);
or U12784 (N_12784,N_12639,N_12611);
and U12785 (N_12785,N_12669,N_12654);
and U12786 (N_12786,N_12590,N_12546);
or U12787 (N_12787,N_12615,N_12622);
nand U12788 (N_12788,N_12549,N_12625);
xnor U12789 (N_12789,N_12508,N_12667);
nor U12790 (N_12790,N_12653,N_12530);
xor U12791 (N_12791,N_12588,N_12630);
or U12792 (N_12792,N_12698,N_12619);
or U12793 (N_12793,N_12574,N_12691);
nor U12794 (N_12794,N_12512,N_12572);
or U12795 (N_12795,N_12674,N_12741);
xor U12796 (N_12796,N_12592,N_12604);
nor U12797 (N_12797,N_12749,N_12526);
or U12798 (N_12798,N_12717,N_12540);
nand U12799 (N_12799,N_12632,N_12562);
nor U12800 (N_12800,N_12581,N_12597);
nor U12801 (N_12801,N_12662,N_12614);
or U12802 (N_12802,N_12744,N_12709);
nand U12803 (N_12803,N_12510,N_12647);
or U12804 (N_12804,N_12529,N_12601);
nand U12805 (N_12805,N_12722,N_12532);
and U12806 (N_12806,N_12687,N_12704);
xor U12807 (N_12807,N_12633,N_12699);
or U12808 (N_12808,N_12547,N_12679);
nor U12809 (N_12809,N_12583,N_12515);
nand U12810 (N_12810,N_12671,N_12655);
nand U12811 (N_12811,N_12545,N_12620);
xnor U12812 (N_12812,N_12714,N_12683);
xnor U12813 (N_12813,N_12623,N_12646);
xor U12814 (N_12814,N_12740,N_12580);
or U12815 (N_12815,N_12738,N_12561);
and U12816 (N_12816,N_12715,N_12606);
nand U12817 (N_12817,N_12729,N_12628);
or U12818 (N_12818,N_12617,N_12656);
xnor U12819 (N_12819,N_12577,N_12706);
or U12820 (N_12820,N_12593,N_12745);
and U12821 (N_12821,N_12718,N_12689);
nand U12822 (N_12822,N_12686,N_12665);
and U12823 (N_12823,N_12652,N_12737);
nand U12824 (N_12824,N_12692,N_12521);
xor U12825 (N_12825,N_12672,N_12658);
nand U12826 (N_12826,N_12570,N_12524);
and U12827 (N_12827,N_12525,N_12591);
nand U12828 (N_12828,N_12705,N_12513);
and U12829 (N_12829,N_12624,N_12579);
and U12830 (N_12830,N_12556,N_12645);
and U12831 (N_12831,N_12668,N_12700);
or U12832 (N_12832,N_12518,N_12719);
xor U12833 (N_12833,N_12576,N_12634);
nand U12834 (N_12834,N_12504,N_12543);
nor U12835 (N_12835,N_12641,N_12598);
nor U12836 (N_12836,N_12678,N_12747);
nor U12837 (N_12837,N_12560,N_12610);
and U12838 (N_12838,N_12511,N_12675);
or U12839 (N_12839,N_12551,N_12535);
nand U12840 (N_12840,N_12676,N_12609);
or U12841 (N_12841,N_12627,N_12724);
and U12842 (N_12842,N_12534,N_12651);
nor U12843 (N_12843,N_12648,N_12613);
nor U12844 (N_12844,N_12555,N_12542);
or U12845 (N_12845,N_12519,N_12501);
nor U12846 (N_12846,N_12677,N_12710);
nor U12847 (N_12847,N_12571,N_12587);
or U12848 (N_12848,N_12734,N_12713);
or U12849 (N_12849,N_12585,N_12748);
and U12850 (N_12850,N_12596,N_12735);
nand U12851 (N_12851,N_12640,N_12527);
and U12852 (N_12852,N_12716,N_12707);
xnor U12853 (N_12853,N_12661,N_12536);
nand U12854 (N_12854,N_12612,N_12506);
or U12855 (N_12855,N_12642,N_12600);
xnor U12856 (N_12856,N_12693,N_12649);
or U12857 (N_12857,N_12673,N_12659);
nor U12858 (N_12858,N_12559,N_12635);
xor U12859 (N_12859,N_12568,N_12599);
xnor U12860 (N_12860,N_12631,N_12553);
nand U12861 (N_12861,N_12712,N_12602);
and U12862 (N_12862,N_12701,N_12743);
xnor U12863 (N_12863,N_12682,N_12608);
and U12864 (N_12864,N_12711,N_12688);
or U12865 (N_12865,N_12533,N_12517);
or U12866 (N_12866,N_12636,N_12569);
nand U12867 (N_12867,N_12522,N_12595);
xor U12868 (N_12868,N_12603,N_12725);
nor U12869 (N_12869,N_12721,N_12696);
nor U12870 (N_12870,N_12538,N_12730);
nor U12871 (N_12871,N_12573,N_12537);
nor U12872 (N_12872,N_12528,N_12681);
or U12873 (N_12873,N_12548,N_12550);
or U12874 (N_12874,N_12739,N_12657);
and U12875 (N_12875,N_12568,N_12630);
nand U12876 (N_12876,N_12704,N_12540);
nor U12877 (N_12877,N_12611,N_12714);
and U12878 (N_12878,N_12587,N_12683);
xor U12879 (N_12879,N_12653,N_12741);
and U12880 (N_12880,N_12509,N_12520);
xnor U12881 (N_12881,N_12666,N_12595);
xor U12882 (N_12882,N_12645,N_12646);
nor U12883 (N_12883,N_12604,N_12524);
nor U12884 (N_12884,N_12656,N_12638);
nand U12885 (N_12885,N_12639,N_12575);
or U12886 (N_12886,N_12666,N_12622);
nor U12887 (N_12887,N_12743,N_12591);
and U12888 (N_12888,N_12529,N_12621);
and U12889 (N_12889,N_12708,N_12701);
nand U12890 (N_12890,N_12690,N_12682);
nand U12891 (N_12891,N_12701,N_12506);
or U12892 (N_12892,N_12702,N_12517);
xor U12893 (N_12893,N_12676,N_12502);
xor U12894 (N_12894,N_12722,N_12530);
or U12895 (N_12895,N_12562,N_12527);
xnor U12896 (N_12896,N_12576,N_12505);
xnor U12897 (N_12897,N_12511,N_12725);
nor U12898 (N_12898,N_12511,N_12583);
nor U12899 (N_12899,N_12569,N_12719);
and U12900 (N_12900,N_12714,N_12571);
xnor U12901 (N_12901,N_12666,N_12582);
or U12902 (N_12902,N_12594,N_12729);
nand U12903 (N_12903,N_12576,N_12555);
nor U12904 (N_12904,N_12730,N_12633);
nand U12905 (N_12905,N_12655,N_12628);
and U12906 (N_12906,N_12668,N_12549);
nor U12907 (N_12907,N_12523,N_12515);
or U12908 (N_12908,N_12689,N_12612);
nor U12909 (N_12909,N_12532,N_12601);
xor U12910 (N_12910,N_12642,N_12704);
xor U12911 (N_12911,N_12564,N_12635);
nand U12912 (N_12912,N_12741,N_12536);
nor U12913 (N_12913,N_12631,N_12685);
or U12914 (N_12914,N_12735,N_12636);
and U12915 (N_12915,N_12635,N_12622);
nor U12916 (N_12916,N_12506,N_12623);
xnor U12917 (N_12917,N_12648,N_12524);
nor U12918 (N_12918,N_12596,N_12545);
nor U12919 (N_12919,N_12628,N_12653);
nor U12920 (N_12920,N_12595,N_12524);
xnor U12921 (N_12921,N_12659,N_12617);
xnor U12922 (N_12922,N_12510,N_12666);
xor U12923 (N_12923,N_12736,N_12502);
xor U12924 (N_12924,N_12653,N_12503);
nor U12925 (N_12925,N_12554,N_12737);
or U12926 (N_12926,N_12595,N_12646);
nand U12927 (N_12927,N_12598,N_12678);
and U12928 (N_12928,N_12509,N_12697);
or U12929 (N_12929,N_12523,N_12543);
xor U12930 (N_12930,N_12730,N_12620);
xnor U12931 (N_12931,N_12554,N_12543);
nand U12932 (N_12932,N_12505,N_12643);
xnor U12933 (N_12933,N_12547,N_12564);
nor U12934 (N_12934,N_12502,N_12536);
nand U12935 (N_12935,N_12675,N_12534);
or U12936 (N_12936,N_12638,N_12663);
or U12937 (N_12937,N_12512,N_12650);
xnor U12938 (N_12938,N_12719,N_12703);
nand U12939 (N_12939,N_12673,N_12539);
xor U12940 (N_12940,N_12546,N_12705);
or U12941 (N_12941,N_12554,N_12671);
and U12942 (N_12942,N_12635,N_12674);
nand U12943 (N_12943,N_12616,N_12574);
or U12944 (N_12944,N_12665,N_12518);
nand U12945 (N_12945,N_12644,N_12732);
and U12946 (N_12946,N_12745,N_12638);
xnor U12947 (N_12947,N_12712,N_12634);
nor U12948 (N_12948,N_12625,N_12648);
xnor U12949 (N_12949,N_12606,N_12534);
or U12950 (N_12950,N_12653,N_12542);
xnor U12951 (N_12951,N_12508,N_12576);
nor U12952 (N_12952,N_12744,N_12584);
nand U12953 (N_12953,N_12625,N_12731);
xor U12954 (N_12954,N_12622,N_12531);
nor U12955 (N_12955,N_12509,N_12582);
nand U12956 (N_12956,N_12590,N_12577);
nor U12957 (N_12957,N_12541,N_12687);
nand U12958 (N_12958,N_12644,N_12522);
xor U12959 (N_12959,N_12695,N_12738);
nand U12960 (N_12960,N_12686,N_12620);
or U12961 (N_12961,N_12625,N_12525);
nor U12962 (N_12962,N_12508,N_12682);
nand U12963 (N_12963,N_12604,N_12570);
xnor U12964 (N_12964,N_12725,N_12684);
or U12965 (N_12965,N_12506,N_12731);
or U12966 (N_12966,N_12742,N_12650);
nor U12967 (N_12967,N_12542,N_12514);
xnor U12968 (N_12968,N_12640,N_12668);
and U12969 (N_12969,N_12583,N_12537);
and U12970 (N_12970,N_12674,N_12587);
nor U12971 (N_12971,N_12601,N_12593);
nand U12972 (N_12972,N_12692,N_12621);
and U12973 (N_12973,N_12660,N_12545);
xnor U12974 (N_12974,N_12615,N_12580);
and U12975 (N_12975,N_12676,N_12733);
xnor U12976 (N_12976,N_12696,N_12649);
xnor U12977 (N_12977,N_12666,N_12643);
xnor U12978 (N_12978,N_12641,N_12737);
and U12979 (N_12979,N_12618,N_12520);
nor U12980 (N_12980,N_12600,N_12724);
xor U12981 (N_12981,N_12578,N_12641);
nand U12982 (N_12982,N_12723,N_12579);
and U12983 (N_12983,N_12550,N_12668);
xnor U12984 (N_12984,N_12689,N_12513);
xor U12985 (N_12985,N_12642,N_12592);
xnor U12986 (N_12986,N_12550,N_12631);
nand U12987 (N_12987,N_12526,N_12586);
nand U12988 (N_12988,N_12508,N_12648);
or U12989 (N_12989,N_12647,N_12544);
nor U12990 (N_12990,N_12659,N_12671);
or U12991 (N_12991,N_12564,N_12738);
xnor U12992 (N_12992,N_12559,N_12655);
nor U12993 (N_12993,N_12698,N_12662);
and U12994 (N_12994,N_12730,N_12631);
nor U12995 (N_12995,N_12593,N_12589);
nand U12996 (N_12996,N_12651,N_12726);
and U12997 (N_12997,N_12706,N_12651);
nand U12998 (N_12998,N_12700,N_12675);
xor U12999 (N_12999,N_12619,N_12519);
or U13000 (N_13000,N_12894,N_12988);
and U13001 (N_13001,N_12828,N_12990);
and U13002 (N_13002,N_12935,N_12998);
nand U13003 (N_13003,N_12964,N_12987);
xnor U13004 (N_13004,N_12941,N_12889);
nor U13005 (N_13005,N_12875,N_12816);
xor U13006 (N_13006,N_12837,N_12933);
nand U13007 (N_13007,N_12824,N_12829);
and U13008 (N_13008,N_12939,N_12975);
or U13009 (N_13009,N_12836,N_12916);
or U13010 (N_13010,N_12831,N_12902);
nand U13011 (N_13011,N_12764,N_12968);
nand U13012 (N_13012,N_12761,N_12995);
or U13013 (N_13013,N_12900,N_12843);
xnor U13014 (N_13014,N_12912,N_12890);
nand U13015 (N_13015,N_12910,N_12810);
nand U13016 (N_13016,N_12946,N_12842);
xor U13017 (N_13017,N_12788,N_12940);
xor U13018 (N_13018,N_12880,N_12781);
or U13019 (N_13019,N_12770,N_12906);
xor U13020 (N_13020,N_12814,N_12758);
and U13021 (N_13021,N_12957,N_12978);
nor U13022 (N_13022,N_12963,N_12895);
xor U13023 (N_13023,N_12898,N_12942);
xor U13024 (N_13024,N_12918,N_12999);
nor U13025 (N_13025,N_12974,N_12773);
xor U13026 (N_13026,N_12982,N_12896);
nand U13027 (N_13027,N_12769,N_12780);
and U13028 (N_13028,N_12838,N_12822);
nor U13029 (N_13029,N_12930,N_12751);
nand U13030 (N_13030,N_12911,N_12960);
and U13031 (N_13031,N_12803,N_12871);
nand U13032 (N_13032,N_12864,N_12955);
nand U13033 (N_13033,N_12887,N_12983);
xnor U13034 (N_13034,N_12791,N_12779);
xnor U13035 (N_13035,N_12905,N_12782);
and U13036 (N_13036,N_12937,N_12823);
nor U13037 (N_13037,N_12841,N_12818);
or U13038 (N_13038,N_12771,N_12966);
xor U13039 (N_13039,N_12899,N_12929);
nand U13040 (N_13040,N_12932,N_12945);
or U13041 (N_13041,N_12952,N_12976);
or U13042 (N_13042,N_12830,N_12931);
and U13043 (N_13043,N_12778,N_12949);
and U13044 (N_13044,N_12756,N_12926);
or U13045 (N_13045,N_12868,N_12969);
nand U13046 (N_13046,N_12921,N_12877);
nor U13047 (N_13047,N_12884,N_12762);
or U13048 (N_13048,N_12844,N_12786);
nor U13049 (N_13049,N_12792,N_12907);
or U13050 (N_13050,N_12821,N_12938);
and U13051 (N_13051,N_12768,N_12919);
nand U13052 (N_13052,N_12790,N_12794);
and U13053 (N_13053,N_12886,N_12853);
and U13054 (N_13054,N_12973,N_12971);
xor U13055 (N_13055,N_12840,N_12909);
and U13056 (N_13056,N_12981,N_12878);
nand U13057 (N_13057,N_12994,N_12901);
nand U13058 (N_13058,N_12904,N_12867);
or U13059 (N_13059,N_12846,N_12860);
nand U13060 (N_13060,N_12834,N_12857);
and U13061 (N_13061,N_12908,N_12950);
nor U13062 (N_13062,N_12760,N_12953);
xor U13063 (N_13063,N_12977,N_12859);
xor U13064 (N_13064,N_12783,N_12980);
xor U13065 (N_13065,N_12934,N_12839);
or U13066 (N_13066,N_12806,N_12811);
xor U13067 (N_13067,N_12766,N_12797);
or U13068 (N_13068,N_12777,N_12984);
nand U13069 (N_13069,N_12928,N_12925);
or U13070 (N_13070,N_12956,N_12826);
or U13071 (N_13071,N_12775,N_12845);
or U13072 (N_13072,N_12865,N_12776);
and U13073 (N_13073,N_12858,N_12936);
nand U13074 (N_13074,N_12892,N_12870);
or U13075 (N_13075,N_12827,N_12787);
nor U13076 (N_13076,N_12804,N_12789);
xnor U13077 (N_13077,N_12863,N_12913);
or U13078 (N_13078,N_12753,N_12873);
or U13079 (N_13079,N_12833,N_12813);
nand U13080 (N_13080,N_12820,N_12874);
xor U13081 (N_13081,N_12798,N_12817);
nand U13082 (N_13082,N_12832,N_12799);
or U13083 (N_13083,N_12883,N_12989);
and U13084 (N_13084,N_12772,N_12914);
nor U13085 (N_13085,N_12855,N_12954);
nor U13086 (N_13086,N_12847,N_12888);
and U13087 (N_13087,N_12872,N_12805);
nand U13088 (N_13088,N_12991,N_12767);
nand U13089 (N_13089,N_12763,N_12948);
or U13090 (N_13090,N_12915,N_12996);
and U13091 (N_13091,N_12795,N_12757);
and U13092 (N_13092,N_12849,N_12986);
nor U13093 (N_13093,N_12961,N_12951);
nor U13094 (N_13094,N_12882,N_12759);
xor U13095 (N_13095,N_12881,N_12851);
xor U13096 (N_13096,N_12774,N_12862);
xnor U13097 (N_13097,N_12924,N_12812);
nor U13098 (N_13098,N_12885,N_12807);
or U13099 (N_13099,N_12808,N_12835);
and U13100 (N_13100,N_12785,N_12848);
and U13101 (N_13101,N_12819,N_12893);
or U13102 (N_13102,N_12943,N_12869);
nor U13103 (N_13103,N_12972,N_12861);
xor U13104 (N_13104,N_12962,N_12917);
xor U13105 (N_13105,N_12796,N_12997);
and U13106 (N_13106,N_12755,N_12866);
or U13107 (N_13107,N_12927,N_12947);
nor U13108 (N_13108,N_12754,N_12944);
or U13109 (N_13109,N_12992,N_12876);
or U13110 (N_13110,N_12802,N_12879);
or U13111 (N_13111,N_12852,N_12897);
nand U13112 (N_13112,N_12815,N_12801);
nand U13113 (N_13113,N_12922,N_12979);
nor U13114 (N_13114,N_12850,N_12800);
nor U13115 (N_13115,N_12923,N_12958);
nand U13116 (N_13116,N_12765,N_12809);
nand U13117 (N_13117,N_12920,N_12993);
nand U13118 (N_13118,N_12967,N_12891);
xor U13119 (N_13119,N_12752,N_12825);
and U13120 (N_13120,N_12970,N_12985);
and U13121 (N_13121,N_12854,N_12965);
or U13122 (N_13122,N_12856,N_12750);
nor U13123 (N_13123,N_12959,N_12903);
or U13124 (N_13124,N_12793,N_12784);
nor U13125 (N_13125,N_12927,N_12832);
or U13126 (N_13126,N_12977,N_12816);
and U13127 (N_13127,N_12857,N_12914);
nor U13128 (N_13128,N_12997,N_12766);
nor U13129 (N_13129,N_12773,N_12785);
xor U13130 (N_13130,N_12913,N_12808);
nor U13131 (N_13131,N_12791,N_12761);
nand U13132 (N_13132,N_12776,N_12924);
xnor U13133 (N_13133,N_12768,N_12961);
or U13134 (N_13134,N_12936,N_12752);
or U13135 (N_13135,N_12788,N_12833);
nor U13136 (N_13136,N_12778,N_12943);
nand U13137 (N_13137,N_12984,N_12869);
nand U13138 (N_13138,N_12994,N_12968);
and U13139 (N_13139,N_12756,N_12818);
and U13140 (N_13140,N_12807,N_12957);
or U13141 (N_13141,N_12794,N_12883);
nand U13142 (N_13142,N_12912,N_12861);
and U13143 (N_13143,N_12793,N_12898);
and U13144 (N_13144,N_12911,N_12863);
or U13145 (N_13145,N_12983,N_12879);
nand U13146 (N_13146,N_12995,N_12778);
or U13147 (N_13147,N_12940,N_12958);
and U13148 (N_13148,N_12995,N_12855);
nor U13149 (N_13149,N_12987,N_12795);
xnor U13150 (N_13150,N_12793,N_12805);
and U13151 (N_13151,N_12890,N_12801);
or U13152 (N_13152,N_12776,N_12751);
nor U13153 (N_13153,N_12929,N_12833);
xor U13154 (N_13154,N_12792,N_12824);
nand U13155 (N_13155,N_12825,N_12971);
nand U13156 (N_13156,N_12853,N_12762);
xor U13157 (N_13157,N_12763,N_12803);
and U13158 (N_13158,N_12860,N_12755);
nor U13159 (N_13159,N_12767,N_12947);
nor U13160 (N_13160,N_12907,N_12969);
nand U13161 (N_13161,N_12847,N_12944);
nor U13162 (N_13162,N_12811,N_12892);
nor U13163 (N_13163,N_12863,N_12972);
nor U13164 (N_13164,N_12908,N_12898);
nor U13165 (N_13165,N_12852,N_12946);
or U13166 (N_13166,N_12825,N_12875);
and U13167 (N_13167,N_12800,N_12997);
and U13168 (N_13168,N_12810,N_12797);
or U13169 (N_13169,N_12822,N_12803);
and U13170 (N_13170,N_12904,N_12771);
and U13171 (N_13171,N_12864,N_12757);
nor U13172 (N_13172,N_12953,N_12924);
or U13173 (N_13173,N_12926,N_12767);
and U13174 (N_13174,N_12877,N_12911);
nor U13175 (N_13175,N_12906,N_12894);
nor U13176 (N_13176,N_12908,N_12762);
xor U13177 (N_13177,N_12768,N_12819);
xnor U13178 (N_13178,N_12821,N_12999);
nand U13179 (N_13179,N_12939,N_12814);
and U13180 (N_13180,N_12958,N_12985);
nand U13181 (N_13181,N_12888,N_12952);
and U13182 (N_13182,N_12760,N_12890);
or U13183 (N_13183,N_12890,N_12851);
or U13184 (N_13184,N_12988,N_12863);
xor U13185 (N_13185,N_12794,N_12916);
xnor U13186 (N_13186,N_12851,N_12786);
xor U13187 (N_13187,N_12860,N_12803);
nor U13188 (N_13188,N_12980,N_12769);
nor U13189 (N_13189,N_12864,N_12831);
and U13190 (N_13190,N_12951,N_12865);
nor U13191 (N_13191,N_12832,N_12902);
nor U13192 (N_13192,N_12920,N_12819);
xnor U13193 (N_13193,N_12760,N_12955);
and U13194 (N_13194,N_12998,N_12761);
or U13195 (N_13195,N_12785,N_12908);
xor U13196 (N_13196,N_12997,N_12866);
nor U13197 (N_13197,N_12769,N_12927);
or U13198 (N_13198,N_12992,N_12917);
or U13199 (N_13199,N_12801,N_12894);
nand U13200 (N_13200,N_12967,N_12849);
and U13201 (N_13201,N_12780,N_12887);
nor U13202 (N_13202,N_12789,N_12890);
nand U13203 (N_13203,N_12793,N_12895);
or U13204 (N_13204,N_12996,N_12767);
xnor U13205 (N_13205,N_12917,N_12889);
or U13206 (N_13206,N_12918,N_12769);
or U13207 (N_13207,N_12943,N_12865);
xor U13208 (N_13208,N_12753,N_12981);
or U13209 (N_13209,N_12971,N_12985);
and U13210 (N_13210,N_12989,N_12878);
and U13211 (N_13211,N_12870,N_12786);
nor U13212 (N_13212,N_12956,N_12785);
xnor U13213 (N_13213,N_12759,N_12829);
nor U13214 (N_13214,N_12758,N_12823);
and U13215 (N_13215,N_12887,N_12966);
and U13216 (N_13216,N_12834,N_12971);
xnor U13217 (N_13217,N_12831,N_12822);
or U13218 (N_13218,N_12992,N_12919);
nor U13219 (N_13219,N_12979,N_12831);
and U13220 (N_13220,N_12933,N_12904);
xnor U13221 (N_13221,N_12829,N_12898);
nor U13222 (N_13222,N_12965,N_12940);
or U13223 (N_13223,N_12786,N_12853);
nand U13224 (N_13224,N_12768,N_12783);
nor U13225 (N_13225,N_12884,N_12816);
and U13226 (N_13226,N_12982,N_12886);
nand U13227 (N_13227,N_12888,N_12912);
and U13228 (N_13228,N_12867,N_12926);
xnor U13229 (N_13229,N_12991,N_12958);
and U13230 (N_13230,N_12908,N_12843);
nor U13231 (N_13231,N_12769,N_12992);
or U13232 (N_13232,N_12881,N_12886);
or U13233 (N_13233,N_12919,N_12968);
or U13234 (N_13234,N_12821,N_12769);
and U13235 (N_13235,N_12940,N_12836);
nand U13236 (N_13236,N_12873,N_12771);
xnor U13237 (N_13237,N_12868,N_12872);
or U13238 (N_13238,N_12751,N_12892);
or U13239 (N_13239,N_12874,N_12865);
nand U13240 (N_13240,N_12803,N_12771);
and U13241 (N_13241,N_12960,N_12835);
nor U13242 (N_13242,N_12757,N_12974);
xnor U13243 (N_13243,N_12995,N_12754);
xnor U13244 (N_13244,N_12969,N_12945);
or U13245 (N_13245,N_12978,N_12833);
xnor U13246 (N_13246,N_12918,N_12803);
and U13247 (N_13247,N_12832,N_12795);
nor U13248 (N_13248,N_12975,N_12879);
or U13249 (N_13249,N_12765,N_12934);
and U13250 (N_13250,N_13201,N_13109);
nor U13251 (N_13251,N_13077,N_13079);
nand U13252 (N_13252,N_13125,N_13126);
or U13253 (N_13253,N_13247,N_13103);
or U13254 (N_13254,N_13135,N_13165);
or U13255 (N_13255,N_13214,N_13147);
nor U13256 (N_13256,N_13166,N_13243);
nand U13257 (N_13257,N_13001,N_13118);
or U13258 (N_13258,N_13073,N_13024);
nor U13259 (N_13259,N_13014,N_13074);
nand U13260 (N_13260,N_13102,N_13233);
nand U13261 (N_13261,N_13101,N_13167);
or U13262 (N_13262,N_13041,N_13042);
nand U13263 (N_13263,N_13010,N_13211);
and U13264 (N_13264,N_13168,N_13016);
or U13265 (N_13265,N_13098,N_13054);
and U13266 (N_13266,N_13129,N_13008);
nor U13267 (N_13267,N_13195,N_13113);
nand U13268 (N_13268,N_13203,N_13178);
and U13269 (N_13269,N_13163,N_13065);
nand U13270 (N_13270,N_13090,N_13157);
nand U13271 (N_13271,N_13036,N_13022);
nor U13272 (N_13272,N_13087,N_13068);
nand U13273 (N_13273,N_13116,N_13064);
nand U13274 (N_13274,N_13249,N_13177);
and U13275 (N_13275,N_13207,N_13197);
nor U13276 (N_13276,N_13175,N_13111);
nor U13277 (N_13277,N_13245,N_13217);
xor U13278 (N_13278,N_13162,N_13239);
nand U13279 (N_13279,N_13152,N_13134);
and U13280 (N_13280,N_13131,N_13194);
and U13281 (N_13281,N_13170,N_13023);
nor U13282 (N_13282,N_13062,N_13019);
nand U13283 (N_13283,N_13212,N_13055);
or U13284 (N_13284,N_13048,N_13185);
or U13285 (N_13285,N_13080,N_13060);
or U13286 (N_13286,N_13138,N_13000);
xnor U13287 (N_13287,N_13198,N_13226);
nand U13288 (N_13288,N_13063,N_13104);
nor U13289 (N_13289,N_13121,N_13150);
nand U13290 (N_13290,N_13066,N_13047);
xor U13291 (N_13291,N_13037,N_13058);
nor U13292 (N_13292,N_13230,N_13221);
and U13293 (N_13293,N_13199,N_13137);
nand U13294 (N_13294,N_13020,N_13021);
nand U13295 (N_13295,N_13205,N_13200);
and U13296 (N_13296,N_13049,N_13191);
nand U13297 (N_13297,N_13088,N_13210);
xnor U13298 (N_13298,N_13108,N_13144);
and U13299 (N_13299,N_13114,N_13035);
and U13300 (N_13300,N_13120,N_13218);
and U13301 (N_13301,N_13061,N_13181);
nand U13302 (N_13302,N_13159,N_13187);
or U13303 (N_13303,N_13220,N_13034);
and U13304 (N_13304,N_13209,N_13133);
or U13305 (N_13305,N_13161,N_13228);
nand U13306 (N_13306,N_13190,N_13117);
nor U13307 (N_13307,N_13004,N_13172);
nand U13308 (N_13308,N_13011,N_13017);
or U13309 (N_13309,N_13127,N_13240);
or U13310 (N_13310,N_13174,N_13204);
or U13311 (N_13311,N_13069,N_13094);
or U13312 (N_13312,N_13176,N_13160);
or U13313 (N_13313,N_13151,N_13100);
nor U13314 (N_13314,N_13189,N_13179);
nor U13315 (N_13315,N_13095,N_13208);
nand U13316 (N_13316,N_13012,N_13216);
or U13317 (N_13317,N_13028,N_13196);
nor U13318 (N_13318,N_13076,N_13026);
nand U13319 (N_13319,N_13231,N_13043);
or U13320 (N_13320,N_13033,N_13132);
or U13321 (N_13321,N_13053,N_13072);
xnor U13322 (N_13322,N_13219,N_13171);
or U13323 (N_13323,N_13097,N_13139);
or U13324 (N_13324,N_13070,N_13227);
nand U13325 (N_13325,N_13237,N_13156);
or U13326 (N_13326,N_13025,N_13099);
and U13327 (N_13327,N_13009,N_13248);
nand U13328 (N_13328,N_13224,N_13141);
and U13329 (N_13329,N_13184,N_13059);
nand U13330 (N_13330,N_13164,N_13078);
nor U13331 (N_13331,N_13182,N_13091);
nand U13332 (N_13332,N_13155,N_13051);
xor U13333 (N_13333,N_13232,N_13085);
and U13334 (N_13334,N_13083,N_13096);
and U13335 (N_13335,N_13031,N_13056);
and U13336 (N_13336,N_13112,N_13192);
and U13337 (N_13337,N_13006,N_13110);
and U13338 (N_13338,N_13046,N_13235);
and U13339 (N_13339,N_13044,N_13119);
and U13340 (N_13340,N_13149,N_13222);
nand U13341 (N_13341,N_13032,N_13081);
xnor U13342 (N_13342,N_13052,N_13234);
nor U13343 (N_13343,N_13115,N_13169);
xor U13344 (N_13344,N_13093,N_13084);
nand U13345 (N_13345,N_13158,N_13107);
and U13346 (N_13346,N_13106,N_13071);
or U13347 (N_13347,N_13246,N_13213);
xor U13348 (N_13348,N_13050,N_13173);
or U13349 (N_13349,N_13193,N_13153);
xor U13350 (N_13350,N_13154,N_13105);
xor U13351 (N_13351,N_13242,N_13236);
xor U13352 (N_13352,N_13123,N_13206);
nand U13353 (N_13353,N_13244,N_13030);
xnor U13354 (N_13354,N_13003,N_13186);
nor U13355 (N_13355,N_13045,N_13027);
or U13356 (N_13356,N_13075,N_13124);
xnor U13357 (N_13357,N_13140,N_13223);
nand U13358 (N_13358,N_13146,N_13183);
xor U13359 (N_13359,N_13241,N_13130);
or U13360 (N_13360,N_13180,N_13142);
nor U13361 (N_13361,N_13143,N_13018);
or U13362 (N_13362,N_13148,N_13215);
or U13363 (N_13363,N_13002,N_13089);
and U13364 (N_13364,N_13122,N_13225);
nor U13365 (N_13365,N_13188,N_13039);
or U13366 (N_13366,N_13007,N_13145);
nand U13367 (N_13367,N_13082,N_13013);
or U13368 (N_13368,N_13005,N_13128);
nor U13369 (N_13369,N_13092,N_13057);
nor U13370 (N_13370,N_13229,N_13202);
nor U13371 (N_13371,N_13015,N_13038);
nor U13372 (N_13372,N_13238,N_13136);
and U13373 (N_13373,N_13040,N_13029);
or U13374 (N_13374,N_13067,N_13086);
nand U13375 (N_13375,N_13109,N_13156);
nor U13376 (N_13376,N_13104,N_13086);
nand U13377 (N_13377,N_13060,N_13002);
xor U13378 (N_13378,N_13116,N_13199);
and U13379 (N_13379,N_13055,N_13029);
nand U13380 (N_13380,N_13045,N_13100);
nor U13381 (N_13381,N_13098,N_13108);
and U13382 (N_13382,N_13163,N_13028);
nor U13383 (N_13383,N_13128,N_13022);
and U13384 (N_13384,N_13249,N_13087);
or U13385 (N_13385,N_13142,N_13213);
and U13386 (N_13386,N_13060,N_13035);
xor U13387 (N_13387,N_13210,N_13171);
xnor U13388 (N_13388,N_13201,N_13025);
nor U13389 (N_13389,N_13023,N_13101);
or U13390 (N_13390,N_13052,N_13053);
nor U13391 (N_13391,N_13094,N_13239);
and U13392 (N_13392,N_13140,N_13058);
nor U13393 (N_13393,N_13078,N_13165);
xor U13394 (N_13394,N_13229,N_13220);
nor U13395 (N_13395,N_13115,N_13225);
or U13396 (N_13396,N_13183,N_13205);
xnor U13397 (N_13397,N_13095,N_13140);
or U13398 (N_13398,N_13154,N_13050);
nor U13399 (N_13399,N_13109,N_13202);
and U13400 (N_13400,N_13077,N_13053);
xor U13401 (N_13401,N_13158,N_13245);
or U13402 (N_13402,N_13181,N_13117);
nor U13403 (N_13403,N_13101,N_13135);
nand U13404 (N_13404,N_13176,N_13206);
nor U13405 (N_13405,N_13138,N_13242);
or U13406 (N_13406,N_13240,N_13198);
and U13407 (N_13407,N_13089,N_13197);
and U13408 (N_13408,N_13045,N_13052);
nand U13409 (N_13409,N_13106,N_13159);
nand U13410 (N_13410,N_13043,N_13182);
and U13411 (N_13411,N_13110,N_13072);
nor U13412 (N_13412,N_13045,N_13241);
xnor U13413 (N_13413,N_13096,N_13232);
nand U13414 (N_13414,N_13234,N_13163);
and U13415 (N_13415,N_13168,N_13126);
nand U13416 (N_13416,N_13116,N_13030);
nor U13417 (N_13417,N_13199,N_13192);
nor U13418 (N_13418,N_13191,N_13178);
xor U13419 (N_13419,N_13102,N_13037);
nor U13420 (N_13420,N_13015,N_13055);
xor U13421 (N_13421,N_13092,N_13072);
or U13422 (N_13422,N_13119,N_13159);
and U13423 (N_13423,N_13248,N_13051);
or U13424 (N_13424,N_13041,N_13023);
nand U13425 (N_13425,N_13222,N_13069);
nand U13426 (N_13426,N_13229,N_13203);
nand U13427 (N_13427,N_13167,N_13083);
nor U13428 (N_13428,N_13211,N_13142);
nand U13429 (N_13429,N_13166,N_13195);
nor U13430 (N_13430,N_13191,N_13018);
or U13431 (N_13431,N_13083,N_13114);
nand U13432 (N_13432,N_13072,N_13203);
and U13433 (N_13433,N_13192,N_13123);
or U13434 (N_13434,N_13168,N_13046);
nand U13435 (N_13435,N_13013,N_13106);
nand U13436 (N_13436,N_13115,N_13153);
or U13437 (N_13437,N_13154,N_13091);
or U13438 (N_13438,N_13168,N_13100);
nor U13439 (N_13439,N_13245,N_13233);
xnor U13440 (N_13440,N_13033,N_13194);
nand U13441 (N_13441,N_13002,N_13219);
xor U13442 (N_13442,N_13036,N_13085);
xor U13443 (N_13443,N_13225,N_13083);
nor U13444 (N_13444,N_13244,N_13208);
and U13445 (N_13445,N_13116,N_13140);
nand U13446 (N_13446,N_13047,N_13010);
and U13447 (N_13447,N_13176,N_13199);
and U13448 (N_13448,N_13205,N_13089);
nor U13449 (N_13449,N_13030,N_13155);
nand U13450 (N_13450,N_13013,N_13104);
and U13451 (N_13451,N_13214,N_13030);
and U13452 (N_13452,N_13011,N_13061);
and U13453 (N_13453,N_13094,N_13002);
nor U13454 (N_13454,N_13118,N_13177);
and U13455 (N_13455,N_13104,N_13019);
nand U13456 (N_13456,N_13001,N_13055);
xnor U13457 (N_13457,N_13233,N_13236);
nand U13458 (N_13458,N_13215,N_13247);
or U13459 (N_13459,N_13180,N_13217);
nand U13460 (N_13460,N_13080,N_13219);
and U13461 (N_13461,N_13228,N_13159);
nand U13462 (N_13462,N_13236,N_13050);
or U13463 (N_13463,N_13245,N_13050);
xnor U13464 (N_13464,N_13218,N_13175);
nand U13465 (N_13465,N_13204,N_13111);
nand U13466 (N_13466,N_13077,N_13085);
nand U13467 (N_13467,N_13011,N_13070);
nor U13468 (N_13468,N_13093,N_13237);
nand U13469 (N_13469,N_13212,N_13201);
xor U13470 (N_13470,N_13165,N_13208);
xnor U13471 (N_13471,N_13179,N_13099);
nor U13472 (N_13472,N_13104,N_13112);
and U13473 (N_13473,N_13006,N_13100);
and U13474 (N_13474,N_13135,N_13117);
and U13475 (N_13475,N_13247,N_13145);
and U13476 (N_13476,N_13111,N_13211);
xnor U13477 (N_13477,N_13039,N_13049);
xnor U13478 (N_13478,N_13076,N_13120);
nand U13479 (N_13479,N_13059,N_13068);
nor U13480 (N_13480,N_13058,N_13069);
xor U13481 (N_13481,N_13066,N_13034);
and U13482 (N_13482,N_13073,N_13157);
and U13483 (N_13483,N_13122,N_13174);
nand U13484 (N_13484,N_13214,N_13235);
or U13485 (N_13485,N_13023,N_13230);
nor U13486 (N_13486,N_13239,N_13207);
and U13487 (N_13487,N_13198,N_13179);
nor U13488 (N_13488,N_13037,N_13018);
and U13489 (N_13489,N_13164,N_13133);
nor U13490 (N_13490,N_13176,N_13184);
or U13491 (N_13491,N_13200,N_13120);
xor U13492 (N_13492,N_13015,N_13185);
and U13493 (N_13493,N_13215,N_13198);
or U13494 (N_13494,N_13164,N_13141);
nand U13495 (N_13495,N_13055,N_13083);
xnor U13496 (N_13496,N_13202,N_13098);
nand U13497 (N_13497,N_13192,N_13149);
xor U13498 (N_13498,N_13046,N_13125);
nor U13499 (N_13499,N_13246,N_13185);
and U13500 (N_13500,N_13371,N_13447);
and U13501 (N_13501,N_13404,N_13491);
nor U13502 (N_13502,N_13322,N_13439);
or U13503 (N_13503,N_13428,N_13300);
and U13504 (N_13504,N_13457,N_13389);
nand U13505 (N_13505,N_13263,N_13286);
and U13506 (N_13506,N_13272,N_13476);
xnor U13507 (N_13507,N_13383,N_13398);
or U13508 (N_13508,N_13477,N_13352);
nand U13509 (N_13509,N_13358,N_13429);
nor U13510 (N_13510,N_13258,N_13334);
or U13511 (N_13511,N_13379,N_13408);
nand U13512 (N_13512,N_13285,N_13327);
nand U13513 (N_13513,N_13472,N_13329);
and U13514 (N_13514,N_13259,N_13435);
xor U13515 (N_13515,N_13335,N_13475);
and U13516 (N_13516,N_13438,N_13431);
nor U13517 (N_13517,N_13448,N_13490);
or U13518 (N_13518,N_13316,N_13461);
and U13519 (N_13519,N_13416,N_13267);
nor U13520 (N_13520,N_13305,N_13264);
nor U13521 (N_13521,N_13410,N_13463);
nor U13522 (N_13522,N_13310,N_13271);
and U13523 (N_13523,N_13455,N_13366);
and U13524 (N_13524,N_13433,N_13406);
nor U13525 (N_13525,N_13464,N_13283);
xor U13526 (N_13526,N_13466,N_13434);
nand U13527 (N_13527,N_13426,N_13260);
and U13528 (N_13528,N_13391,N_13284);
nand U13529 (N_13529,N_13384,N_13498);
and U13530 (N_13530,N_13486,N_13360);
nand U13531 (N_13531,N_13301,N_13478);
and U13532 (N_13532,N_13397,N_13456);
or U13533 (N_13533,N_13315,N_13320);
nor U13534 (N_13534,N_13376,N_13390);
nand U13535 (N_13535,N_13417,N_13324);
xnor U13536 (N_13536,N_13295,N_13276);
nor U13537 (N_13537,N_13338,N_13446);
nand U13538 (N_13538,N_13350,N_13370);
or U13539 (N_13539,N_13251,N_13441);
nor U13540 (N_13540,N_13344,N_13458);
xnor U13541 (N_13541,N_13277,N_13420);
xor U13542 (N_13542,N_13396,N_13336);
xnor U13543 (N_13543,N_13402,N_13467);
nand U13544 (N_13544,N_13373,N_13422);
and U13545 (N_13545,N_13400,N_13432);
or U13546 (N_13546,N_13298,N_13293);
xor U13547 (N_13547,N_13484,N_13311);
xor U13548 (N_13548,N_13321,N_13265);
xor U13549 (N_13549,N_13330,N_13489);
nand U13550 (N_13550,N_13362,N_13473);
and U13551 (N_13551,N_13280,N_13262);
or U13552 (N_13552,N_13436,N_13407);
nand U13553 (N_13553,N_13409,N_13314);
or U13554 (N_13554,N_13303,N_13392);
and U13555 (N_13555,N_13480,N_13325);
or U13556 (N_13556,N_13361,N_13288);
and U13557 (N_13557,N_13382,N_13424);
xor U13558 (N_13558,N_13318,N_13340);
nor U13559 (N_13559,N_13412,N_13430);
nor U13560 (N_13560,N_13359,N_13339);
xor U13561 (N_13561,N_13306,N_13401);
or U13562 (N_13562,N_13375,N_13282);
nand U13563 (N_13563,N_13343,N_13469);
or U13564 (N_13564,N_13348,N_13481);
nor U13565 (N_13565,N_13421,N_13452);
and U13566 (N_13566,N_13483,N_13419);
xnor U13567 (N_13567,N_13323,N_13427);
or U13568 (N_13568,N_13440,N_13257);
or U13569 (N_13569,N_13279,N_13395);
nor U13570 (N_13570,N_13291,N_13328);
and U13571 (N_13571,N_13363,N_13281);
nand U13572 (N_13572,N_13368,N_13333);
xor U13573 (N_13573,N_13474,N_13462);
or U13574 (N_13574,N_13380,N_13250);
nor U13575 (N_13575,N_13302,N_13270);
and U13576 (N_13576,N_13304,N_13425);
nor U13577 (N_13577,N_13274,N_13387);
or U13578 (N_13578,N_13308,N_13442);
or U13579 (N_13579,N_13256,N_13471);
or U13580 (N_13580,N_13444,N_13485);
nand U13581 (N_13581,N_13253,N_13292);
nand U13582 (N_13582,N_13351,N_13492);
nor U13583 (N_13583,N_13299,N_13342);
or U13584 (N_13584,N_13495,N_13346);
or U13585 (N_13585,N_13399,N_13414);
or U13586 (N_13586,N_13355,N_13273);
nor U13587 (N_13587,N_13468,N_13347);
xor U13588 (N_13588,N_13411,N_13294);
or U13589 (N_13589,N_13287,N_13369);
nor U13590 (N_13590,N_13364,N_13415);
nand U13591 (N_13591,N_13367,N_13496);
and U13592 (N_13592,N_13307,N_13393);
and U13593 (N_13593,N_13377,N_13365);
xor U13594 (N_13594,N_13296,N_13488);
and U13595 (N_13595,N_13261,N_13317);
nand U13596 (N_13596,N_13494,N_13413);
or U13597 (N_13597,N_13482,N_13297);
and U13598 (N_13598,N_13449,N_13266);
nand U13599 (N_13599,N_13451,N_13386);
and U13600 (N_13600,N_13269,N_13443);
nand U13601 (N_13601,N_13312,N_13354);
and U13602 (N_13602,N_13337,N_13453);
nor U13603 (N_13603,N_13385,N_13313);
or U13604 (N_13604,N_13372,N_13278);
and U13605 (N_13605,N_13331,N_13405);
xnor U13606 (N_13606,N_13499,N_13357);
nand U13607 (N_13607,N_13319,N_13374);
or U13608 (N_13608,N_13487,N_13356);
xor U13609 (N_13609,N_13309,N_13454);
or U13610 (N_13610,N_13378,N_13403);
nor U13611 (N_13611,N_13341,N_13275);
and U13612 (N_13612,N_13290,N_13445);
nor U13613 (N_13613,N_13459,N_13252);
or U13614 (N_13614,N_13381,N_13349);
nand U13615 (N_13615,N_13388,N_13289);
or U13616 (N_13616,N_13493,N_13418);
xnor U13617 (N_13617,N_13254,N_13450);
xnor U13618 (N_13618,N_13470,N_13268);
xor U13619 (N_13619,N_13497,N_13255);
and U13620 (N_13620,N_13437,N_13423);
xor U13621 (N_13621,N_13479,N_13353);
xnor U13622 (N_13622,N_13345,N_13332);
nor U13623 (N_13623,N_13465,N_13460);
and U13624 (N_13624,N_13326,N_13394);
and U13625 (N_13625,N_13375,N_13316);
nor U13626 (N_13626,N_13299,N_13277);
and U13627 (N_13627,N_13306,N_13305);
nor U13628 (N_13628,N_13275,N_13327);
and U13629 (N_13629,N_13444,N_13307);
nand U13630 (N_13630,N_13347,N_13272);
nand U13631 (N_13631,N_13433,N_13400);
nor U13632 (N_13632,N_13366,N_13277);
xnor U13633 (N_13633,N_13314,N_13265);
xor U13634 (N_13634,N_13450,N_13335);
and U13635 (N_13635,N_13432,N_13489);
and U13636 (N_13636,N_13469,N_13271);
and U13637 (N_13637,N_13254,N_13465);
nand U13638 (N_13638,N_13401,N_13489);
nand U13639 (N_13639,N_13261,N_13276);
nor U13640 (N_13640,N_13424,N_13361);
nand U13641 (N_13641,N_13318,N_13397);
xnor U13642 (N_13642,N_13258,N_13398);
and U13643 (N_13643,N_13295,N_13476);
or U13644 (N_13644,N_13327,N_13351);
xnor U13645 (N_13645,N_13480,N_13395);
nand U13646 (N_13646,N_13251,N_13317);
or U13647 (N_13647,N_13369,N_13379);
and U13648 (N_13648,N_13380,N_13419);
nor U13649 (N_13649,N_13259,N_13288);
or U13650 (N_13650,N_13410,N_13327);
xnor U13651 (N_13651,N_13442,N_13491);
xnor U13652 (N_13652,N_13437,N_13331);
xor U13653 (N_13653,N_13376,N_13454);
and U13654 (N_13654,N_13497,N_13330);
xor U13655 (N_13655,N_13297,N_13292);
xnor U13656 (N_13656,N_13473,N_13333);
and U13657 (N_13657,N_13411,N_13270);
xnor U13658 (N_13658,N_13422,N_13309);
and U13659 (N_13659,N_13267,N_13440);
xor U13660 (N_13660,N_13457,N_13291);
xnor U13661 (N_13661,N_13356,N_13320);
or U13662 (N_13662,N_13393,N_13351);
nand U13663 (N_13663,N_13478,N_13434);
or U13664 (N_13664,N_13461,N_13306);
or U13665 (N_13665,N_13420,N_13334);
or U13666 (N_13666,N_13332,N_13344);
xor U13667 (N_13667,N_13424,N_13329);
nand U13668 (N_13668,N_13256,N_13326);
or U13669 (N_13669,N_13439,N_13415);
xor U13670 (N_13670,N_13302,N_13477);
xnor U13671 (N_13671,N_13448,N_13459);
xnor U13672 (N_13672,N_13297,N_13497);
xor U13673 (N_13673,N_13268,N_13322);
and U13674 (N_13674,N_13440,N_13284);
nand U13675 (N_13675,N_13379,N_13362);
nor U13676 (N_13676,N_13455,N_13388);
and U13677 (N_13677,N_13348,N_13336);
nand U13678 (N_13678,N_13422,N_13455);
or U13679 (N_13679,N_13402,N_13421);
and U13680 (N_13680,N_13276,N_13477);
and U13681 (N_13681,N_13477,N_13373);
nand U13682 (N_13682,N_13359,N_13405);
or U13683 (N_13683,N_13345,N_13409);
nor U13684 (N_13684,N_13258,N_13364);
nand U13685 (N_13685,N_13409,N_13406);
and U13686 (N_13686,N_13470,N_13392);
and U13687 (N_13687,N_13447,N_13265);
and U13688 (N_13688,N_13404,N_13358);
nand U13689 (N_13689,N_13452,N_13415);
xor U13690 (N_13690,N_13292,N_13499);
xnor U13691 (N_13691,N_13393,N_13314);
nand U13692 (N_13692,N_13283,N_13390);
or U13693 (N_13693,N_13410,N_13311);
xor U13694 (N_13694,N_13402,N_13444);
and U13695 (N_13695,N_13261,N_13284);
xnor U13696 (N_13696,N_13313,N_13352);
nand U13697 (N_13697,N_13309,N_13398);
and U13698 (N_13698,N_13409,N_13273);
xor U13699 (N_13699,N_13311,N_13477);
and U13700 (N_13700,N_13389,N_13329);
xnor U13701 (N_13701,N_13330,N_13450);
xnor U13702 (N_13702,N_13330,N_13409);
or U13703 (N_13703,N_13255,N_13352);
and U13704 (N_13704,N_13384,N_13360);
xnor U13705 (N_13705,N_13346,N_13472);
nor U13706 (N_13706,N_13353,N_13369);
nor U13707 (N_13707,N_13324,N_13353);
nand U13708 (N_13708,N_13420,N_13465);
xor U13709 (N_13709,N_13459,N_13389);
or U13710 (N_13710,N_13272,N_13457);
xor U13711 (N_13711,N_13342,N_13458);
or U13712 (N_13712,N_13343,N_13363);
or U13713 (N_13713,N_13330,N_13364);
or U13714 (N_13714,N_13460,N_13296);
or U13715 (N_13715,N_13450,N_13444);
and U13716 (N_13716,N_13472,N_13466);
nor U13717 (N_13717,N_13495,N_13402);
or U13718 (N_13718,N_13354,N_13435);
xor U13719 (N_13719,N_13311,N_13308);
nor U13720 (N_13720,N_13425,N_13376);
or U13721 (N_13721,N_13495,N_13445);
xor U13722 (N_13722,N_13445,N_13359);
nand U13723 (N_13723,N_13274,N_13438);
xnor U13724 (N_13724,N_13278,N_13410);
and U13725 (N_13725,N_13421,N_13292);
and U13726 (N_13726,N_13281,N_13406);
xor U13727 (N_13727,N_13379,N_13411);
and U13728 (N_13728,N_13460,N_13269);
and U13729 (N_13729,N_13372,N_13407);
nor U13730 (N_13730,N_13417,N_13426);
and U13731 (N_13731,N_13440,N_13324);
and U13732 (N_13732,N_13406,N_13332);
or U13733 (N_13733,N_13256,N_13330);
and U13734 (N_13734,N_13477,N_13452);
nand U13735 (N_13735,N_13319,N_13471);
xor U13736 (N_13736,N_13495,N_13268);
nand U13737 (N_13737,N_13319,N_13259);
nor U13738 (N_13738,N_13387,N_13333);
nor U13739 (N_13739,N_13452,N_13404);
and U13740 (N_13740,N_13314,N_13279);
and U13741 (N_13741,N_13433,N_13334);
or U13742 (N_13742,N_13438,N_13261);
or U13743 (N_13743,N_13441,N_13486);
nor U13744 (N_13744,N_13255,N_13262);
nand U13745 (N_13745,N_13347,N_13391);
nand U13746 (N_13746,N_13425,N_13308);
and U13747 (N_13747,N_13470,N_13407);
nor U13748 (N_13748,N_13434,N_13326);
xor U13749 (N_13749,N_13483,N_13387);
or U13750 (N_13750,N_13577,N_13727);
nor U13751 (N_13751,N_13503,N_13535);
and U13752 (N_13752,N_13624,N_13643);
xnor U13753 (N_13753,N_13629,N_13572);
xor U13754 (N_13754,N_13670,N_13743);
nor U13755 (N_13755,N_13518,N_13730);
nor U13756 (N_13756,N_13693,N_13704);
nand U13757 (N_13757,N_13640,N_13563);
nor U13758 (N_13758,N_13610,N_13548);
nand U13759 (N_13759,N_13644,N_13722);
nor U13760 (N_13760,N_13666,N_13595);
xnor U13761 (N_13761,N_13502,N_13632);
and U13762 (N_13762,N_13700,N_13663);
and U13763 (N_13763,N_13559,N_13635);
nor U13764 (N_13764,N_13534,N_13618);
nand U13765 (N_13765,N_13708,N_13584);
nand U13766 (N_13766,N_13556,N_13542);
nand U13767 (N_13767,N_13639,N_13701);
nor U13768 (N_13768,N_13593,N_13723);
nand U13769 (N_13769,N_13519,N_13672);
nor U13770 (N_13770,N_13637,N_13516);
nand U13771 (N_13771,N_13552,N_13575);
nor U13772 (N_13772,N_13605,N_13737);
and U13773 (N_13773,N_13716,N_13689);
nand U13774 (N_13774,N_13523,N_13719);
xnor U13775 (N_13775,N_13718,N_13697);
nand U13776 (N_13776,N_13735,N_13705);
xor U13777 (N_13777,N_13696,N_13597);
xnor U13778 (N_13778,N_13564,N_13504);
and U13779 (N_13779,N_13538,N_13527);
xor U13780 (N_13780,N_13550,N_13617);
nor U13781 (N_13781,N_13533,N_13684);
and U13782 (N_13782,N_13678,N_13698);
and U13783 (N_13783,N_13553,N_13611);
or U13784 (N_13784,N_13603,N_13565);
xnor U13785 (N_13785,N_13626,N_13540);
nor U13786 (N_13786,N_13671,N_13668);
and U13787 (N_13787,N_13537,N_13561);
or U13788 (N_13788,N_13745,N_13649);
nor U13789 (N_13789,N_13622,N_13562);
nor U13790 (N_13790,N_13739,N_13501);
nand U13791 (N_13791,N_13638,N_13586);
or U13792 (N_13792,N_13583,N_13692);
nor U13793 (N_13793,N_13608,N_13582);
and U13794 (N_13794,N_13709,N_13529);
nor U13795 (N_13795,N_13526,N_13683);
nor U13796 (N_13796,N_13657,N_13660);
xnor U13797 (N_13797,N_13620,N_13713);
and U13798 (N_13798,N_13733,N_13512);
or U13799 (N_13799,N_13742,N_13513);
or U13800 (N_13800,N_13659,N_13728);
nand U13801 (N_13801,N_13568,N_13715);
or U13802 (N_13802,N_13546,N_13569);
or U13803 (N_13803,N_13566,N_13601);
and U13804 (N_13804,N_13645,N_13514);
nor U13805 (N_13805,N_13604,N_13656);
and U13806 (N_13806,N_13675,N_13686);
or U13807 (N_13807,N_13658,N_13636);
and U13808 (N_13808,N_13500,N_13746);
xor U13809 (N_13809,N_13695,N_13647);
nand U13810 (N_13810,N_13631,N_13613);
and U13811 (N_13811,N_13541,N_13736);
or U13812 (N_13812,N_13623,N_13633);
nand U13813 (N_13813,N_13574,N_13655);
or U13814 (N_13814,N_13691,N_13600);
and U13815 (N_13815,N_13654,N_13676);
nor U13816 (N_13816,N_13625,N_13641);
or U13817 (N_13817,N_13560,N_13594);
xor U13818 (N_13818,N_13528,N_13525);
nor U13819 (N_13819,N_13521,N_13734);
and U13820 (N_13820,N_13615,N_13576);
nand U13821 (N_13821,N_13724,N_13642);
or U13822 (N_13822,N_13619,N_13509);
and U13823 (N_13823,N_13581,N_13726);
nand U13824 (N_13824,N_13515,N_13703);
nand U13825 (N_13825,N_13628,N_13585);
and U13826 (N_13826,N_13662,N_13598);
and U13827 (N_13827,N_13589,N_13711);
nor U13828 (N_13828,N_13580,N_13749);
and U13829 (N_13829,N_13681,N_13536);
xor U13830 (N_13830,N_13543,N_13731);
or U13831 (N_13831,N_13524,N_13511);
nand U13832 (N_13832,N_13721,N_13707);
nand U13833 (N_13833,N_13591,N_13549);
or U13834 (N_13834,N_13532,N_13522);
and U13835 (N_13835,N_13680,N_13720);
or U13836 (N_13836,N_13510,N_13621);
nand U13837 (N_13837,N_13652,N_13612);
and U13838 (N_13838,N_13587,N_13682);
or U13839 (N_13839,N_13599,N_13725);
xor U13840 (N_13840,N_13554,N_13741);
or U13841 (N_13841,N_13596,N_13664);
nand U13842 (N_13842,N_13714,N_13505);
or U13843 (N_13843,N_13588,N_13571);
and U13844 (N_13844,N_13517,N_13602);
nand U13845 (N_13845,N_13740,N_13531);
xor U13846 (N_13846,N_13558,N_13627);
nor U13847 (N_13847,N_13732,N_13673);
and U13848 (N_13848,N_13699,N_13653);
nand U13849 (N_13849,N_13573,N_13606);
or U13850 (N_13850,N_13747,N_13661);
nand U13851 (N_13851,N_13687,N_13557);
nor U13852 (N_13852,N_13646,N_13551);
xor U13853 (N_13853,N_13545,N_13729);
and U13854 (N_13854,N_13578,N_13690);
xor U13855 (N_13855,N_13634,N_13555);
nand U13856 (N_13856,N_13674,N_13570);
nor U13857 (N_13857,N_13607,N_13579);
xor U13858 (N_13858,N_13669,N_13539);
or U13859 (N_13859,N_13520,N_13508);
xor U13860 (N_13860,N_13544,N_13665);
and U13861 (N_13861,N_13614,N_13738);
nand U13862 (N_13862,N_13677,N_13706);
xor U13863 (N_13863,N_13744,N_13609);
and U13864 (N_13864,N_13507,N_13748);
or U13865 (N_13865,N_13650,N_13616);
xor U13866 (N_13866,N_13530,N_13651);
nand U13867 (N_13867,N_13710,N_13688);
or U13868 (N_13868,N_13630,N_13712);
nor U13869 (N_13869,N_13567,N_13702);
and U13870 (N_13870,N_13694,N_13590);
or U13871 (N_13871,N_13685,N_13648);
nor U13872 (N_13872,N_13592,N_13667);
and U13873 (N_13873,N_13717,N_13506);
nor U13874 (N_13874,N_13679,N_13547);
and U13875 (N_13875,N_13538,N_13700);
nor U13876 (N_13876,N_13527,N_13569);
or U13877 (N_13877,N_13695,N_13719);
nor U13878 (N_13878,N_13634,N_13638);
or U13879 (N_13879,N_13705,N_13528);
nand U13880 (N_13880,N_13671,N_13585);
nor U13881 (N_13881,N_13532,N_13625);
nand U13882 (N_13882,N_13532,N_13659);
and U13883 (N_13883,N_13540,N_13700);
nor U13884 (N_13884,N_13688,N_13518);
nor U13885 (N_13885,N_13716,N_13737);
or U13886 (N_13886,N_13651,N_13683);
nand U13887 (N_13887,N_13523,N_13641);
nor U13888 (N_13888,N_13740,N_13587);
and U13889 (N_13889,N_13727,N_13668);
nor U13890 (N_13890,N_13551,N_13629);
nand U13891 (N_13891,N_13747,N_13689);
nor U13892 (N_13892,N_13632,N_13566);
nand U13893 (N_13893,N_13609,N_13543);
nor U13894 (N_13894,N_13506,N_13697);
or U13895 (N_13895,N_13629,N_13525);
and U13896 (N_13896,N_13554,N_13688);
xnor U13897 (N_13897,N_13733,N_13735);
xnor U13898 (N_13898,N_13507,N_13509);
and U13899 (N_13899,N_13666,N_13535);
and U13900 (N_13900,N_13701,N_13662);
and U13901 (N_13901,N_13608,N_13575);
or U13902 (N_13902,N_13612,N_13650);
nand U13903 (N_13903,N_13625,N_13622);
and U13904 (N_13904,N_13514,N_13738);
or U13905 (N_13905,N_13565,N_13747);
and U13906 (N_13906,N_13639,N_13678);
nand U13907 (N_13907,N_13614,N_13729);
nor U13908 (N_13908,N_13571,N_13600);
nor U13909 (N_13909,N_13631,N_13743);
nor U13910 (N_13910,N_13596,N_13747);
xor U13911 (N_13911,N_13719,N_13529);
nand U13912 (N_13912,N_13542,N_13675);
and U13913 (N_13913,N_13645,N_13508);
nand U13914 (N_13914,N_13551,N_13604);
xnor U13915 (N_13915,N_13733,N_13589);
nand U13916 (N_13916,N_13502,N_13722);
or U13917 (N_13917,N_13704,N_13567);
and U13918 (N_13918,N_13583,N_13569);
and U13919 (N_13919,N_13500,N_13709);
nand U13920 (N_13920,N_13600,N_13550);
xnor U13921 (N_13921,N_13598,N_13553);
nor U13922 (N_13922,N_13529,N_13516);
nor U13923 (N_13923,N_13622,N_13519);
xor U13924 (N_13924,N_13629,N_13671);
nand U13925 (N_13925,N_13572,N_13506);
nand U13926 (N_13926,N_13565,N_13679);
nand U13927 (N_13927,N_13592,N_13597);
or U13928 (N_13928,N_13661,N_13554);
and U13929 (N_13929,N_13685,N_13700);
nor U13930 (N_13930,N_13702,N_13699);
nand U13931 (N_13931,N_13679,N_13563);
or U13932 (N_13932,N_13569,N_13680);
nand U13933 (N_13933,N_13583,N_13545);
or U13934 (N_13934,N_13703,N_13742);
nand U13935 (N_13935,N_13724,N_13685);
xnor U13936 (N_13936,N_13507,N_13512);
and U13937 (N_13937,N_13716,N_13707);
and U13938 (N_13938,N_13619,N_13693);
and U13939 (N_13939,N_13530,N_13580);
nand U13940 (N_13940,N_13638,N_13615);
or U13941 (N_13941,N_13542,N_13557);
nand U13942 (N_13942,N_13682,N_13617);
nand U13943 (N_13943,N_13659,N_13651);
xor U13944 (N_13944,N_13637,N_13691);
and U13945 (N_13945,N_13613,N_13502);
nor U13946 (N_13946,N_13654,N_13519);
xor U13947 (N_13947,N_13736,N_13732);
and U13948 (N_13948,N_13583,N_13686);
or U13949 (N_13949,N_13596,N_13501);
or U13950 (N_13950,N_13560,N_13529);
nor U13951 (N_13951,N_13545,N_13659);
xor U13952 (N_13952,N_13743,N_13576);
or U13953 (N_13953,N_13700,N_13683);
nand U13954 (N_13954,N_13719,N_13574);
nor U13955 (N_13955,N_13719,N_13614);
or U13956 (N_13956,N_13590,N_13601);
or U13957 (N_13957,N_13595,N_13568);
or U13958 (N_13958,N_13745,N_13601);
nand U13959 (N_13959,N_13593,N_13685);
nand U13960 (N_13960,N_13510,N_13624);
nor U13961 (N_13961,N_13505,N_13738);
nand U13962 (N_13962,N_13526,N_13517);
nor U13963 (N_13963,N_13655,N_13641);
and U13964 (N_13964,N_13545,N_13530);
and U13965 (N_13965,N_13669,N_13668);
nand U13966 (N_13966,N_13592,N_13680);
and U13967 (N_13967,N_13502,N_13600);
nor U13968 (N_13968,N_13637,N_13522);
xnor U13969 (N_13969,N_13689,N_13552);
nor U13970 (N_13970,N_13673,N_13692);
and U13971 (N_13971,N_13561,N_13533);
xnor U13972 (N_13972,N_13596,N_13580);
nand U13973 (N_13973,N_13690,N_13564);
nor U13974 (N_13974,N_13594,N_13638);
nand U13975 (N_13975,N_13735,N_13597);
nand U13976 (N_13976,N_13734,N_13700);
nand U13977 (N_13977,N_13552,N_13634);
nor U13978 (N_13978,N_13629,N_13719);
and U13979 (N_13979,N_13509,N_13540);
xnor U13980 (N_13980,N_13504,N_13749);
xor U13981 (N_13981,N_13505,N_13668);
or U13982 (N_13982,N_13569,N_13666);
or U13983 (N_13983,N_13664,N_13539);
and U13984 (N_13984,N_13542,N_13695);
nor U13985 (N_13985,N_13583,N_13508);
xnor U13986 (N_13986,N_13704,N_13686);
nor U13987 (N_13987,N_13645,N_13653);
or U13988 (N_13988,N_13526,N_13702);
or U13989 (N_13989,N_13518,N_13662);
nor U13990 (N_13990,N_13646,N_13624);
nand U13991 (N_13991,N_13655,N_13658);
and U13992 (N_13992,N_13692,N_13668);
nor U13993 (N_13993,N_13607,N_13747);
xor U13994 (N_13994,N_13530,N_13635);
nor U13995 (N_13995,N_13642,N_13739);
xnor U13996 (N_13996,N_13556,N_13662);
or U13997 (N_13997,N_13649,N_13551);
or U13998 (N_13998,N_13748,N_13611);
nand U13999 (N_13999,N_13703,N_13724);
nor U14000 (N_14000,N_13912,N_13803);
xor U14001 (N_14001,N_13913,N_13962);
or U14002 (N_14002,N_13874,N_13951);
xor U14003 (N_14003,N_13753,N_13885);
or U14004 (N_14004,N_13918,N_13869);
and U14005 (N_14005,N_13788,N_13910);
or U14006 (N_14006,N_13833,N_13886);
nand U14007 (N_14007,N_13937,N_13996);
or U14008 (N_14008,N_13783,N_13888);
or U14009 (N_14009,N_13938,N_13959);
nor U14010 (N_14010,N_13855,N_13802);
nand U14011 (N_14011,N_13778,N_13840);
or U14012 (N_14012,N_13862,N_13870);
and U14013 (N_14013,N_13814,N_13812);
and U14014 (N_14014,N_13828,N_13752);
nand U14015 (N_14015,N_13851,N_13977);
or U14016 (N_14016,N_13807,N_13923);
nor U14017 (N_14017,N_13971,N_13976);
nor U14018 (N_14018,N_13901,N_13932);
xnor U14019 (N_14019,N_13956,N_13924);
and U14020 (N_14020,N_13944,N_13772);
nand U14021 (N_14021,N_13825,N_13804);
xor U14022 (N_14022,N_13769,N_13800);
or U14023 (N_14023,N_13987,N_13794);
or U14024 (N_14024,N_13782,N_13751);
and U14025 (N_14025,N_13877,N_13968);
nand U14026 (N_14026,N_13993,N_13879);
nor U14027 (N_14027,N_13907,N_13835);
and U14028 (N_14028,N_13758,N_13767);
and U14029 (N_14029,N_13922,N_13984);
xor U14030 (N_14030,N_13942,N_13954);
and U14031 (N_14031,N_13775,N_13820);
or U14032 (N_14032,N_13891,N_13936);
or U14033 (N_14033,N_13921,N_13982);
nand U14034 (N_14034,N_13784,N_13860);
and U14035 (N_14035,N_13945,N_13779);
or U14036 (N_14036,N_13990,N_13836);
xor U14037 (N_14037,N_13989,N_13952);
or U14038 (N_14038,N_13899,N_13955);
nor U14039 (N_14039,N_13830,N_13792);
nor U14040 (N_14040,N_13897,N_13997);
nand U14041 (N_14041,N_13981,N_13750);
nor U14042 (N_14042,N_13791,N_13966);
or U14043 (N_14043,N_13768,N_13796);
or U14044 (N_14044,N_13838,N_13960);
xor U14045 (N_14045,N_13928,N_13893);
and U14046 (N_14046,N_13905,N_13946);
xnor U14047 (N_14047,N_13809,N_13980);
nor U14048 (N_14048,N_13866,N_13849);
nand U14049 (N_14049,N_13858,N_13850);
or U14050 (N_14050,N_13843,N_13777);
nor U14051 (N_14051,N_13931,N_13771);
nor U14052 (N_14052,N_13839,N_13801);
xnor U14053 (N_14053,N_13822,N_13949);
xor U14054 (N_14054,N_13881,N_13995);
nor U14055 (N_14055,N_13765,N_13917);
and U14056 (N_14056,N_13821,N_13842);
or U14057 (N_14057,N_13759,N_13834);
nand U14058 (N_14058,N_13762,N_13941);
or U14059 (N_14059,N_13785,N_13857);
nor U14060 (N_14060,N_13974,N_13754);
nor U14061 (N_14061,N_13887,N_13882);
nand U14062 (N_14062,N_13983,N_13914);
nor U14063 (N_14063,N_13873,N_13756);
nor U14064 (N_14064,N_13818,N_13935);
nor U14065 (N_14065,N_13805,N_13985);
nor U14066 (N_14066,N_13972,N_13832);
nand U14067 (N_14067,N_13790,N_13911);
and U14068 (N_14068,N_13797,N_13880);
nor U14069 (N_14069,N_13831,N_13950);
xor U14070 (N_14070,N_13898,N_13806);
nand U14071 (N_14071,N_13871,N_13894);
xnor U14072 (N_14072,N_13763,N_13861);
and U14073 (N_14073,N_13813,N_13808);
nor U14074 (N_14074,N_13902,N_13979);
nor U14075 (N_14075,N_13789,N_13991);
and U14076 (N_14076,N_13815,N_13852);
nand U14077 (N_14077,N_13927,N_13774);
and U14078 (N_14078,N_13998,N_13930);
nand U14079 (N_14079,N_13780,N_13837);
nand U14080 (N_14080,N_13863,N_13773);
xor U14081 (N_14081,N_13761,N_13817);
or U14082 (N_14082,N_13865,N_13957);
and U14083 (N_14083,N_13967,N_13755);
xnor U14084 (N_14084,N_13848,N_13829);
nor U14085 (N_14085,N_13940,N_13764);
or U14086 (N_14086,N_13963,N_13823);
nand U14087 (N_14087,N_13856,N_13859);
xnor U14088 (N_14088,N_13845,N_13846);
xnor U14089 (N_14089,N_13994,N_13776);
and U14090 (N_14090,N_13841,N_13884);
nand U14091 (N_14091,N_13770,N_13889);
or U14092 (N_14092,N_13975,N_13915);
or U14093 (N_14093,N_13819,N_13872);
nand U14094 (N_14094,N_13986,N_13757);
nor U14095 (N_14095,N_13875,N_13916);
nand U14096 (N_14096,N_13929,N_13903);
nor U14097 (N_14097,N_13925,N_13908);
nor U14098 (N_14098,N_13933,N_13799);
nor U14099 (N_14099,N_13795,N_13958);
or U14100 (N_14100,N_13853,N_13793);
xor U14101 (N_14101,N_13939,N_13854);
nand U14102 (N_14102,N_13798,N_13892);
nor U14103 (N_14103,N_13787,N_13827);
and U14104 (N_14104,N_13847,N_13781);
nor U14105 (N_14105,N_13978,N_13896);
xor U14106 (N_14106,N_13906,N_13878);
nor U14107 (N_14107,N_13867,N_13973);
xor U14108 (N_14108,N_13826,N_13948);
nor U14109 (N_14109,N_13970,N_13919);
and U14110 (N_14110,N_13965,N_13864);
and U14111 (N_14111,N_13883,N_13876);
or U14112 (N_14112,N_13824,N_13934);
or U14113 (N_14113,N_13816,N_13811);
and U14114 (N_14114,N_13766,N_13943);
nor U14115 (N_14115,N_13900,N_13810);
and U14116 (N_14116,N_13844,N_13895);
xnor U14117 (N_14117,N_13890,N_13992);
xor U14118 (N_14118,N_13920,N_13868);
and U14119 (N_14119,N_13904,N_13953);
nand U14120 (N_14120,N_13786,N_13988);
and U14121 (N_14121,N_13964,N_13926);
nor U14122 (N_14122,N_13760,N_13961);
nand U14123 (N_14123,N_13909,N_13947);
or U14124 (N_14124,N_13969,N_13999);
nor U14125 (N_14125,N_13984,N_13990);
xor U14126 (N_14126,N_13797,N_13953);
xnor U14127 (N_14127,N_13942,N_13781);
xnor U14128 (N_14128,N_13967,N_13795);
or U14129 (N_14129,N_13988,N_13907);
or U14130 (N_14130,N_13963,N_13792);
xor U14131 (N_14131,N_13910,N_13939);
and U14132 (N_14132,N_13873,N_13931);
and U14133 (N_14133,N_13819,N_13761);
xor U14134 (N_14134,N_13756,N_13830);
and U14135 (N_14135,N_13962,N_13859);
nand U14136 (N_14136,N_13822,N_13871);
nand U14137 (N_14137,N_13933,N_13754);
nand U14138 (N_14138,N_13991,N_13847);
nand U14139 (N_14139,N_13817,N_13994);
and U14140 (N_14140,N_13869,N_13814);
xor U14141 (N_14141,N_13943,N_13970);
nand U14142 (N_14142,N_13878,N_13829);
or U14143 (N_14143,N_13753,N_13919);
xnor U14144 (N_14144,N_13981,N_13830);
nor U14145 (N_14145,N_13934,N_13884);
and U14146 (N_14146,N_13755,N_13960);
nand U14147 (N_14147,N_13935,N_13860);
nor U14148 (N_14148,N_13972,N_13969);
or U14149 (N_14149,N_13814,N_13825);
nand U14150 (N_14150,N_13773,N_13801);
nor U14151 (N_14151,N_13885,N_13948);
nand U14152 (N_14152,N_13875,N_13907);
or U14153 (N_14153,N_13966,N_13977);
and U14154 (N_14154,N_13964,N_13985);
nor U14155 (N_14155,N_13790,N_13937);
nand U14156 (N_14156,N_13926,N_13880);
nand U14157 (N_14157,N_13937,N_13926);
or U14158 (N_14158,N_13777,N_13955);
or U14159 (N_14159,N_13906,N_13784);
nor U14160 (N_14160,N_13873,N_13764);
nand U14161 (N_14161,N_13956,N_13895);
and U14162 (N_14162,N_13878,N_13840);
nand U14163 (N_14163,N_13883,N_13994);
nor U14164 (N_14164,N_13750,N_13779);
nand U14165 (N_14165,N_13893,N_13919);
and U14166 (N_14166,N_13842,N_13999);
or U14167 (N_14167,N_13908,N_13932);
nor U14168 (N_14168,N_13754,N_13788);
xor U14169 (N_14169,N_13981,N_13855);
or U14170 (N_14170,N_13849,N_13945);
xor U14171 (N_14171,N_13925,N_13873);
and U14172 (N_14172,N_13840,N_13904);
nand U14173 (N_14173,N_13894,N_13880);
xor U14174 (N_14174,N_13812,N_13876);
xnor U14175 (N_14175,N_13867,N_13966);
nor U14176 (N_14176,N_13834,N_13922);
nor U14177 (N_14177,N_13855,N_13973);
xor U14178 (N_14178,N_13767,N_13989);
and U14179 (N_14179,N_13786,N_13876);
and U14180 (N_14180,N_13842,N_13925);
nor U14181 (N_14181,N_13841,N_13787);
nand U14182 (N_14182,N_13859,N_13968);
nand U14183 (N_14183,N_13836,N_13772);
nand U14184 (N_14184,N_13855,N_13896);
and U14185 (N_14185,N_13793,N_13800);
nand U14186 (N_14186,N_13952,N_13772);
nor U14187 (N_14187,N_13865,N_13963);
or U14188 (N_14188,N_13798,N_13976);
and U14189 (N_14189,N_13855,N_13990);
xnor U14190 (N_14190,N_13785,N_13913);
xor U14191 (N_14191,N_13947,N_13778);
nor U14192 (N_14192,N_13805,N_13825);
nor U14193 (N_14193,N_13976,N_13845);
nor U14194 (N_14194,N_13974,N_13780);
nor U14195 (N_14195,N_13790,N_13797);
xor U14196 (N_14196,N_13858,N_13821);
nand U14197 (N_14197,N_13956,N_13974);
and U14198 (N_14198,N_13918,N_13901);
nand U14199 (N_14199,N_13858,N_13771);
and U14200 (N_14200,N_13990,N_13789);
or U14201 (N_14201,N_13897,N_13803);
nand U14202 (N_14202,N_13889,N_13792);
nor U14203 (N_14203,N_13770,N_13956);
nor U14204 (N_14204,N_13780,N_13941);
nand U14205 (N_14205,N_13970,N_13924);
nand U14206 (N_14206,N_13977,N_13817);
and U14207 (N_14207,N_13758,N_13944);
or U14208 (N_14208,N_13842,N_13819);
nor U14209 (N_14209,N_13927,N_13840);
nor U14210 (N_14210,N_13756,N_13894);
nand U14211 (N_14211,N_13838,N_13773);
xnor U14212 (N_14212,N_13879,N_13901);
nand U14213 (N_14213,N_13943,N_13822);
nand U14214 (N_14214,N_13841,N_13891);
nor U14215 (N_14215,N_13937,N_13777);
xor U14216 (N_14216,N_13765,N_13793);
xnor U14217 (N_14217,N_13893,N_13830);
xor U14218 (N_14218,N_13864,N_13773);
xnor U14219 (N_14219,N_13775,N_13900);
nand U14220 (N_14220,N_13943,N_13782);
or U14221 (N_14221,N_13751,N_13780);
xor U14222 (N_14222,N_13965,N_13931);
and U14223 (N_14223,N_13969,N_13792);
nand U14224 (N_14224,N_13819,N_13921);
xnor U14225 (N_14225,N_13921,N_13895);
xnor U14226 (N_14226,N_13900,N_13785);
and U14227 (N_14227,N_13896,N_13875);
and U14228 (N_14228,N_13873,N_13888);
and U14229 (N_14229,N_13826,N_13999);
xor U14230 (N_14230,N_13805,N_13925);
and U14231 (N_14231,N_13875,N_13767);
and U14232 (N_14232,N_13852,N_13961);
xnor U14233 (N_14233,N_13773,N_13849);
nor U14234 (N_14234,N_13891,N_13849);
or U14235 (N_14235,N_13993,N_13921);
or U14236 (N_14236,N_13855,N_13778);
and U14237 (N_14237,N_13825,N_13925);
nor U14238 (N_14238,N_13785,N_13834);
nand U14239 (N_14239,N_13943,N_13999);
nand U14240 (N_14240,N_13963,N_13874);
xnor U14241 (N_14241,N_13793,N_13840);
nor U14242 (N_14242,N_13993,N_13848);
nor U14243 (N_14243,N_13871,N_13785);
xnor U14244 (N_14244,N_13891,N_13961);
or U14245 (N_14245,N_13912,N_13916);
nand U14246 (N_14246,N_13834,N_13799);
nor U14247 (N_14247,N_13853,N_13884);
or U14248 (N_14248,N_13971,N_13753);
nor U14249 (N_14249,N_13981,N_13899);
or U14250 (N_14250,N_14118,N_14207);
and U14251 (N_14251,N_14248,N_14180);
and U14252 (N_14252,N_14129,N_14206);
nor U14253 (N_14253,N_14212,N_14196);
nor U14254 (N_14254,N_14140,N_14186);
xor U14255 (N_14255,N_14053,N_14015);
nand U14256 (N_14256,N_14117,N_14052);
nand U14257 (N_14257,N_14193,N_14225);
nor U14258 (N_14258,N_14145,N_14181);
xor U14259 (N_14259,N_14146,N_14008);
xor U14260 (N_14260,N_14203,N_14184);
xnor U14261 (N_14261,N_14169,N_14183);
and U14262 (N_14262,N_14096,N_14107);
nand U14263 (N_14263,N_14137,N_14004);
and U14264 (N_14264,N_14006,N_14178);
or U14265 (N_14265,N_14036,N_14219);
and U14266 (N_14266,N_14158,N_14094);
and U14267 (N_14267,N_14019,N_14204);
and U14268 (N_14268,N_14182,N_14127);
nor U14269 (N_14269,N_14024,N_14039);
nor U14270 (N_14270,N_14033,N_14194);
and U14271 (N_14271,N_14133,N_14195);
and U14272 (N_14272,N_14075,N_14043);
xnor U14273 (N_14273,N_14081,N_14233);
or U14274 (N_14274,N_14162,N_14110);
xor U14275 (N_14275,N_14112,N_14073);
nand U14276 (N_14276,N_14022,N_14124);
nand U14277 (N_14277,N_14243,N_14234);
nand U14278 (N_14278,N_14001,N_14235);
or U14279 (N_14279,N_14069,N_14210);
and U14280 (N_14280,N_14037,N_14168);
or U14281 (N_14281,N_14097,N_14047);
xor U14282 (N_14282,N_14027,N_14056);
nand U14283 (N_14283,N_14163,N_14211);
nand U14284 (N_14284,N_14170,N_14177);
and U14285 (N_14285,N_14029,N_14084);
and U14286 (N_14286,N_14061,N_14245);
and U14287 (N_14287,N_14165,N_14172);
nor U14288 (N_14288,N_14093,N_14231);
or U14289 (N_14289,N_14202,N_14166);
nand U14290 (N_14290,N_14223,N_14188);
or U14291 (N_14291,N_14201,N_14040);
nor U14292 (N_14292,N_14190,N_14200);
xnor U14293 (N_14293,N_14011,N_14142);
nand U14294 (N_14294,N_14007,N_14123);
and U14295 (N_14295,N_14078,N_14113);
and U14296 (N_14296,N_14108,N_14173);
xnor U14297 (N_14297,N_14059,N_14000);
xor U14298 (N_14298,N_14130,N_14187);
and U14299 (N_14299,N_14134,N_14208);
xor U14300 (N_14300,N_14189,N_14085);
nor U14301 (N_14301,N_14109,N_14236);
nand U14302 (N_14302,N_14159,N_14218);
nand U14303 (N_14303,N_14077,N_14128);
nor U14304 (N_14304,N_14242,N_14222);
or U14305 (N_14305,N_14119,N_14063);
and U14306 (N_14306,N_14216,N_14106);
xnor U14307 (N_14307,N_14126,N_14065);
nand U14308 (N_14308,N_14054,N_14164);
nand U14309 (N_14309,N_14066,N_14148);
and U14310 (N_14310,N_14080,N_14224);
nor U14311 (N_14311,N_14012,N_14105);
and U14312 (N_14312,N_14215,N_14030);
and U14313 (N_14313,N_14227,N_14149);
or U14314 (N_14314,N_14120,N_14074);
nand U14315 (N_14315,N_14082,N_14152);
nand U14316 (N_14316,N_14171,N_14249);
and U14317 (N_14317,N_14192,N_14246);
nand U14318 (N_14318,N_14197,N_14028);
or U14319 (N_14319,N_14135,N_14035);
nand U14320 (N_14320,N_14088,N_14092);
and U14321 (N_14321,N_14115,N_14016);
nand U14322 (N_14322,N_14018,N_14058);
or U14323 (N_14323,N_14083,N_14221);
and U14324 (N_14324,N_14101,N_14090);
xnor U14325 (N_14325,N_14241,N_14021);
xnor U14326 (N_14326,N_14157,N_14167);
nor U14327 (N_14327,N_14174,N_14034);
and U14328 (N_14328,N_14091,N_14114);
nand U14329 (N_14329,N_14220,N_14104);
nand U14330 (N_14330,N_14232,N_14214);
and U14331 (N_14331,N_14139,N_14055);
xnor U14332 (N_14332,N_14098,N_14199);
xor U14333 (N_14333,N_14051,N_14138);
nand U14334 (N_14334,N_14057,N_14244);
xor U14335 (N_14335,N_14031,N_14156);
nand U14336 (N_14336,N_14064,N_14131);
xnor U14337 (N_14337,N_14005,N_14143);
nand U14338 (N_14338,N_14191,N_14238);
nand U14339 (N_14339,N_14089,N_14025);
and U14340 (N_14340,N_14002,N_14239);
and U14341 (N_14341,N_14032,N_14237);
nand U14342 (N_14342,N_14072,N_14155);
or U14343 (N_14343,N_14229,N_14044);
nor U14344 (N_14344,N_14151,N_14185);
nand U14345 (N_14345,N_14003,N_14099);
nor U14346 (N_14346,N_14111,N_14086);
xor U14347 (N_14347,N_14042,N_14020);
nor U14348 (N_14348,N_14160,N_14147);
nor U14349 (N_14349,N_14103,N_14010);
xor U14350 (N_14350,N_14049,N_14121);
and U14351 (N_14351,N_14017,N_14013);
and U14352 (N_14352,N_14050,N_14213);
nor U14353 (N_14353,N_14247,N_14048);
nor U14354 (N_14354,N_14023,N_14045);
nor U14355 (N_14355,N_14041,N_14009);
nand U14356 (N_14356,N_14209,N_14154);
nand U14357 (N_14357,N_14076,N_14240);
xor U14358 (N_14358,N_14161,N_14144);
xor U14359 (N_14359,N_14150,N_14141);
and U14360 (N_14360,N_14132,N_14116);
nor U14361 (N_14361,N_14176,N_14095);
or U14362 (N_14362,N_14228,N_14179);
xnor U14363 (N_14363,N_14100,N_14087);
and U14364 (N_14364,N_14067,N_14136);
and U14365 (N_14365,N_14046,N_14060);
and U14366 (N_14366,N_14062,N_14026);
or U14367 (N_14367,N_14079,N_14230);
xnor U14368 (N_14368,N_14071,N_14014);
and U14369 (N_14369,N_14070,N_14068);
xnor U14370 (N_14370,N_14038,N_14175);
xnor U14371 (N_14371,N_14122,N_14125);
xnor U14372 (N_14372,N_14198,N_14217);
nor U14373 (N_14373,N_14205,N_14102);
nor U14374 (N_14374,N_14153,N_14226);
nand U14375 (N_14375,N_14133,N_14050);
and U14376 (N_14376,N_14100,N_14226);
nand U14377 (N_14377,N_14195,N_14161);
xnor U14378 (N_14378,N_14231,N_14071);
or U14379 (N_14379,N_14189,N_14016);
nor U14380 (N_14380,N_14152,N_14186);
nor U14381 (N_14381,N_14186,N_14200);
nand U14382 (N_14382,N_14248,N_14050);
nand U14383 (N_14383,N_14152,N_14206);
nand U14384 (N_14384,N_14241,N_14100);
xor U14385 (N_14385,N_14131,N_14150);
nor U14386 (N_14386,N_14002,N_14186);
nor U14387 (N_14387,N_14234,N_14100);
nor U14388 (N_14388,N_14038,N_14013);
nor U14389 (N_14389,N_14058,N_14094);
nor U14390 (N_14390,N_14129,N_14189);
nand U14391 (N_14391,N_14129,N_14124);
or U14392 (N_14392,N_14208,N_14174);
and U14393 (N_14393,N_14046,N_14218);
xor U14394 (N_14394,N_14226,N_14099);
nor U14395 (N_14395,N_14126,N_14231);
nand U14396 (N_14396,N_14181,N_14024);
xor U14397 (N_14397,N_14125,N_14186);
and U14398 (N_14398,N_14203,N_14200);
xor U14399 (N_14399,N_14114,N_14189);
nor U14400 (N_14400,N_14068,N_14119);
nor U14401 (N_14401,N_14031,N_14017);
nand U14402 (N_14402,N_14121,N_14241);
xor U14403 (N_14403,N_14176,N_14009);
or U14404 (N_14404,N_14229,N_14090);
nor U14405 (N_14405,N_14135,N_14210);
nand U14406 (N_14406,N_14087,N_14109);
nor U14407 (N_14407,N_14175,N_14099);
or U14408 (N_14408,N_14064,N_14194);
nor U14409 (N_14409,N_14173,N_14059);
nor U14410 (N_14410,N_14167,N_14067);
and U14411 (N_14411,N_14219,N_14099);
and U14412 (N_14412,N_14088,N_14056);
and U14413 (N_14413,N_14166,N_14010);
nor U14414 (N_14414,N_14069,N_14029);
nor U14415 (N_14415,N_14146,N_14160);
and U14416 (N_14416,N_14063,N_14073);
or U14417 (N_14417,N_14116,N_14249);
and U14418 (N_14418,N_14070,N_14081);
and U14419 (N_14419,N_14197,N_14072);
xor U14420 (N_14420,N_14026,N_14092);
nor U14421 (N_14421,N_14194,N_14044);
and U14422 (N_14422,N_14216,N_14082);
and U14423 (N_14423,N_14130,N_14156);
or U14424 (N_14424,N_14033,N_14096);
and U14425 (N_14425,N_14010,N_14192);
and U14426 (N_14426,N_14219,N_14230);
nor U14427 (N_14427,N_14081,N_14134);
nor U14428 (N_14428,N_14059,N_14161);
and U14429 (N_14429,N_14207,N_14068);
nor U14430 (N_14430,N_14177,N_14182);
xnor U14431 (N_14431,N_14140,N_14093);
nor U14432 (N_14432,N_14001,N_14089);
and U14433 (N_14433,N_14212,N_14160);
xnor U14434 (N_14434,N_14202,N_14012);
and U14435 (N_14435,N_14154,N_14196);
xnor U14436 (N_14436,N_14015,N_14019);
and U14437 (N_14437,N_14104,N_14135);
nand U14438 (N_14438,N_14138,N_14223);
nand U14439 (N_14439,N_14110,N_14057);
or U14440 (N_14440,N_14164,N_14077);
and U14441 (N_14441,N_14161,N_14039);
xor U14442 (N_14442,N_14076,N_14094);
xor U14443 (N_14443,N_14044,N_14098);
nor U14444 (N_14444,N_14110,N_14071);
or U14445 (N_14445,N_14060,N_14082);
xnor U14446 (N_14446,N_14028,N_14092);
xor U14447 (N_14447,N_14241,N_14103);
nand U14448 (N_14448,N_14128,N_14093);
or U14449 (N_14449,N_14116,N_14162);
and U14450 (N_14450,N_14121,N_14197);
and U14451 (N_14451,N_14072,N_14007);
nand U14452 (N_14452,N_14247,N_14078);
and U14453 (N_14453,N_14112,N_14204);
nand U14454 (N_14454,N_14197,N_14099);
xor U14455 (N_14455,N_14123,N_14091);
xor U14456 (N_14456,N_14157,N_14112);
and U14457 (N_14457,N_14218,N_14081);
nor U14458 (N_14458,N_14115,N_14241);
nand U14459 (N_14459,N_14128,N_14244);
xnor U14460 (N_14460,N_14247,N_14144);
xnor U14461 (N_14461,N_14220,N_14193);
nand U14462 (N_14462,N_14226,N_14172);
or U14463 (N_14463,N_14185,N_14041);
xor U14464 (N_14464,N_14154,N_14182);
nand U14465 (N_14465,N_14219,N_14105);
nand U14466 (N_14466,N_14185,N_14081);
xor U14467 (N_14467,N_14012,N_14074);
xnor U14468 (N_14468,N_14071,N_14103);
nor U14469 (N_14469,N_14230,N_14189);
nor U14470 (N_14470,N_14224,N_14169);
nor U14471 (N_14471,N_14096,N_14158);
nor U14472 (N_14472,N_14158,N_14176);
and U14473 (N_14473,N_14173,N_14134);
nor U14474 (N_14474,N_14021,N_14132);
and U14475 (N_14475,N_14044,N_14169);
xor U14476 (N_14476,N_14098,N_14093);
xor U14477 (N_14477,N_14084,N_14190);
nor U14478 (N_14478,N_14214,N_14004);
nor U14479 (N_14479,N_14001,N_14000);
and U14480 (N_14480,N_14236,N_14001);
nor U14481 (N_14481,N_14180,N_14118);
and U14482 (N_14482,N_14102,N_14095);
or U14483 (N_14483,N_14051,N_14071);
and U14484 (N_14484,N_14028,N_14240);
or U14485 (N_14485,N_14140,N_14152);
and U14486 (N_14486,N_14086,N_14143);
and U14487 (N_14487,N_14033,N_14007);
and U14488 (N_14488,N_14059,N_14145);
nand U14489 (N_14489,N_14132,N_14150);
nor U14490 (N_14490,N_14231,N_14209);
xor U14491 (N_14491,N_14173,N_14113);
nor U14492 (N_14492,N_14244,N_14214);
nor U14493 (N_14493,N_14246,N_14158);
xor U14494 (N_14494,N_14024,N_14200);
nand U14495 (N_14495,N_14205,N_14246);
nor U14496 (N_14496,N_14030,N_14164);
nand U14497 (N_14497,N_14064,N_14155);
or U14498 (N_14498,N_14004,N_14179);
and U14499 (N_14499,N_14142,N_14176);
nand U14500 (N_14500,N_14482,N_14479);
nand U14501 (N_14501,N_14318,N_14453);
and U14502 (N_14502,N_14351,N_14327);
nand U14503 (N_14503,N_14358,N_14276);
nand U14504 (N_14504,N_14348,N_14362);
or U14505 (N_14505,N_14277,N_14308);
or U14506 (N_14506,N_14379,N_14259);
nand U14507 (N_14507,N_14490,N_14408);
and U14508 (N_14508,N_14400,N_14406);
and U14509 (N_14509,N_14294,N_14491);
nand U14510 (N_14510,N_14427,N_14366);
and U14511 (N_14511,N_14342,N_14316);
nor U14512 (N_14512,N_14412,N_14429);
and U14513 (N_14513,N_14452,N_14465);
xnor U14514 (N_14514,N_14459,N_14369);
and U14515 (N_14515,N_14317,N_14447);
and U14516 (N_14516,N_14493,N_14338);
nand U14517 (N_14517,N_14468,N_14345);
nand U14518 (N_14518,N_14344,N_14486);
and U14519 (N_14519,N_14270,N_14446);
nand U14520 (N_14520,N_14315,N_14293);
and U14521 (N_14521,N_14395,N_14332);
or U14522 (N_14522,N_14314,N_14291);
nand U14523 (N_14523,N_14497,N_14492);
and U14524 (N_14524,N_14435,N_14456);
nor U14525 (N_14525,N_14470,N_14454);
nor U14526 (N_14526,N_14361,N_14378);
xnor U14527 (N_14527,N_14352,N_14487);
or U14528 (N_14528,N_14495,N_14275);
or U14529 (N_14529,N_14305,N_14271);
and U14530 (N_14530,N_14250,N_14449);
xor U14531 (N_14531,N_14444,N_14476);
or U14532 (N_14532,N_14253,N_14407);
or U14533 (N_14533,N_14460,N_14295);
or U14534 (N_14534,N_14373,N_14343);
nor U14535 (N_14535,N_14335,N_14274);
nor U14536 (N_14536,N_14310,N_14448);
nand U14537 (N_14537,N_14334,N_14442);
xor U14538 (N_14538,N_14419,N_14304);
xor U14539 (N_14539,N_14363,N_14463);
xor U14540 (N_14540,N_14328,N_14356);
or U14541 (N_14541,N_14282,N_14404);
or U14542 (N_14542,N_14273,N_14477);
xor U14543 (N_14543,N_14472,N_14471);
nand U14544 (N_14544,N_14360,N_14371);
nand U14545 (N_14545,N_14415,N_14322);
nor U14546 (N_14546,N_14279,N_14397);
nand U14547 (N_14547,N_14498,N_14422);
and U14548 (N_14548,N_14300,N_14451);
xnor U14549 (N_14549,N_14414,N_14473);
nand U14550 (N_14550,N_14287,N_14394);
and U14551 (N_14551,N_14264,N_14417);
xor U14552 (N_14552,N_14433,N_14278);
and U14553 (N_14553,N_14461,N_14496);
xnor U14554 (N_14554,N_14464,N_14261);
and U14555 (N_14555,N_14354,N_14483);
xnor U14556 (N_14556,N_14313,N_14268);
nand U14557 (N_14557,N_14372,N_14269);
or U14558 (N_14558,N_14386,N_14330);
nand U14559 (N_14559,N_14481,N_14413);
nand U14560 (N_14560,N_14382,N_14396);
or U14561 (N_14561,N_14280,N_14485);
xor U14562 (N_14562,N_14381,N_14474);
or U14563 (N_14563,N_14391,N_14309);
nand U14564 (N_14564,N_14387,N_14475);
xnor U14565 (N_14565,N_14263,N_14290);
xnor U14566 (N_14566,N_14462,N_14445);
and U14567 (N_14567,N_14424,N_14288);
xor U14568 (N_14568,N_14323,N_14331);
xor U14569 (N_14569,N_14302,N_14306);
nand U14570 (N_14570,N_14311,N_14458);
and U14571 (N_14571,N_14385,N_14421);
nand U14572 (N_14572,N_14281,N_14376);
or U14573 (N_14573,N_14409,N_14437);
or U14574 (N_14574,N_14283,N_14254);
xnor U14575 (N_14575,N_14252,N_14455);
and U14576 (N_14576,N_14499,N_14368);
and U14577 (N_14577,N_14426,N_14402);
nand U14578 (N_14578,N_14301,N_14430);
and U14579 (N_14579,N_14440,N_14267);
nor U14580 (N_14580,N_14494,N_14398);
xnor U14581 (N_14581,N_14292,N_14325);
and U14582 (N_14582,N_14457,N_14340);
nand U14583 (N_14583,N_14296,N_14367);
xnor U14584 (N_14584,N_14262,N_14346);
nor U14585 (N_14585,N_14489,N_14389);
xnor U14586 (N_14586,N_14319,N_14392);
nand U14587 (N_14587,N_14380,N_14403);
and U14588 (N_14588,N_14467,N_14436);
nand U14589 (N_14589,N_14434,N_14307);
nor U14590 (N_14590,N_14439,N_14298);
and U14591 (N_14591,N_14480,N_14370);
nand U14592 (N_14592,N_14388,N_14347);
and U14593 (N_14593,N_14355,N_14425);
or U14594 (N_14594,N_14410,N_14450);
nor U14595 (N_14595,N_14272,N_14432);
nor U14596 (N_14596,N_14350,N_14420);
nor U14597 (N_14597,N_14365,N_14341);
xor U14598 (N_14598,N_14329,N_14423);
or U14599 (N_14599,N_14375,N_14258);
or U14600 (N_14600,N_14321,N_14349);
nor U14601 (N_14601,N_14405,N_14286);
xnor U14602 (N_14602,N_14357,N_14303);
and U14603 (N_14603,N_14390,N_14256);
or U14604 (N_14604,N_14384,N_14443);
nand U14605 (N_14605,N_14393,N_14377);
nor U14606 (N_14606,N_14320,N_14484);
or U14607 (N_14607,N_14428,N_14339);
xor U14608 (N_14608,N_14359,N_14326);
nand U14609 (N_14609,N_14399,N_14364);
or U14610 (N_14610,N_14431,N_14469);
or U14611 (N_14611,N_14488,N_14441);
xnor U14612 (N_14612,N_14255,N_14289);
xor U14613 (N_14613,N_14478,N_14257);
nor U14614 (N_14614,N_14266,N_14401);
xor U14615 (N_14615,N_14260,N_14333);
nand U14616 (N_14616,N_14312,N_14265);
and U14617 (N_14617,N_14418,N_14324);
or U14618 (N_14618,N_14383,N_14299);
or U14619 (N_14619,N_14438,N_14251);
or U14620 (N_14620,N_14337,N_14336);
or U14621 (N_14621,N_14284,N_14285);
nor U14622 (N_14622,N_14353,N_14416);
or U14623 (N_14623,N_14297,N_14374);
or U14624 (N_14624,N_14411,N_14466);
nand U14625 (N_14625,N_14387,N_14474);
or U14626 (N_14626,N_14285,N_14369);
and U14627 (N_14627,N_14353,N_14276);
nand U14628 (N_14628,N_14298,N_14456);
nor U14629 (N_14629,N_14264,N_14254);
nor U14630 (N_14630,N_14260,N_14486);
and U14631 (N_14631,N_14261,N_14257);
and U14632 (N_14632,N_14356,N_14265);
and U14633 (N_14633,N_14406,N_14499);
nor U14634 (N_14634,N_14447,N_14340);
nand U14635 (N_14635,N_14407,N_14477);
and U14636 (N_14636,N_14303,N_14392);
and U14637 (N_14637,N_14421,N_14377);
nor U14638 (N_14638,N_14269,N_14494);
nor U14639 (N_14639,N_14368,N_14332);
xor U14640 (N_14640,N_14252,N_14263);
nand U14641 (N_14641,N_14290,N_14450);
and U14642 (N_14642,N_14285,N_14358);
nor U14643 (N_14643,N_14351,N_14494);
nand U14644 (N_14644,N_14324,N_14277);
or U14645 (N_14645,N_14269,N_14429);
and U14646 (N_14646,N_14264,N_14432);
xnor U14647 (N_14647,N_14418,N_14389);
nand U14648 (N_14648,N_14475,N_14358);
nand U14649 (N_14649,N_14498,N_14468);
and U14650 (N_14650,N_14268,N_14456);
nand U14651 (N_14651,N_14382,N_14367);
and U14652 (N_14652,N_14324,N_14331);
nor U14653 (N_14653,N_14442,N_14351);
or U14654 (N_14654,N_14312,N_14385);
nand U14655 (N_14655,N_14312,N_14420);
or U14656 (N_14656,N_14400,N_14366);
nor U14657 (N_14657,N_14421,N_14478);
nor U14658 (N_14658,N_14335,N_14475);
or U14659 (N_14659,N_14252,N_14405);
nand U14660 (N_14660,N_14420,N_14446);
and U14661 (N_14661,N_14295,N_14321);
and U14662 (N_14662,N_14314,N_14422);
or U14663 (N_14663,N_14470,N_14354);
or U14664 (N_14664,N_14275,N_14440);
or U14665 (N_14665,N_14283,N_14449);
xnor U14666 (N_14666,N_14467,N_14442);
or U14667 (N_14667,N_14463,N_14422);
nand U14668 (N_14668,N_14265,N_14424);
xor U14669 (N_14669,N_14269,N_14441);
nand U14670 (N_14670,N_14473,N_14372);
xor U14671 (N_14671,N_14447,N_14475);
or U14672 (N_14672,N_14326,N_14263);
nand U14673 (N_14673,N_14368,N_14361);
nand U14674 (N_14674,N_14377,N_14484);
nand U14675 (N_14675,N_14399,N_14420);
and U14676 (N_14676,N_14493,N_14455);
xnor U14677 (N_14677,N_14485,N_14318);
nor U14678 (N_14678,N_14452,N_14347);
nand U14679 (N_14679,N_14404,N_14325);
nand U14680 (N_14680,N_14327,N_14322);
and U14681 (N_14681,N_14483,N_14352);
xnor U14682 (N_14682,N_14337,N_14459);
nor U14683 (N_14683,N_14316,N_14420);
nor U14684 (N_14684,N_14486,N_14325);
or U14685 (N_14685,N_14274,N_14425);
or U14686 (N_14686,N_14464,N_14283);
or U14687 (N_14687,N_14384,N_14298);
or U14688 (N_14688,N_14318,N_14351);
xor U14689 (N_14689,N_14301,N_14319);
or U14690 (N_14690,N_14344,N_14435);
or U14691 (N_14691,N_14279,N_14490);
xnor U14692 (N_14692,N_14294,N_14470);
nor U14693 (N_14693,N_14345,N_14318);
xnor U14694 (N_14694,N_14474,N_14261);
and U14695 (N_14695,N_14301,N_14311);
and U14696 (N_14696,N_14436,N_14268);
xnor U14697 (N_14697,N_14283,N_14381);
xnor U14698 (N_14698,N_14297,N_14336);
xnor U14699 (N_14699,N_14387,N_14308);
xnor U14700 (N_14700,N_14334,N_14272);
and U14701 (N_14701,N_14406,N_14346);
nor U14702 (N_14702,N_14336,N_14374);
and U14703 (N_14703,N_14454,N_14324);
or U14704 (N_14704,N_14348,N_14326);
or U14705 (N_14705,N_14365,N_14427);
or U14706 (N_14706,N_14282,N_14403);
nand U14707 (N_14707,N_14285,N_14480);
xnor U14708 (N_14708,N_14343,N_14487);
nand U14709 (N_14709,N_14378,N_14325);
and U14710 (N_14710,N_14342,N_14385);
or U14711 (N_14711,N_14374,N_14483);
nand U14712 (N_14712,N_14424,N_14468);
and U14713 (N_14713,N_14399,N_14320);
nor U14714 (N_14714,N_14484,N_14290);
nand U14715 (N_14715,N_14260,N_14491);
nor U14716 (N_14716,N_14347,N_14424);
or U14717 (N_14717,N_14307,N_14437);
or U14718 (N_14718,N_14273,N_14311);
nand U14719 (N_14719,N_14320,N_14418);
nor U14720 (N_14720,N_14346,N_14289);
nand U14721 (N_14721,N_14362,N_14470);
xor U14722 (N_14722,N_14301,N_14428);
nand U14723 (N_14723,N_14363,N_14452);
xor U14724 (N_14724,N_14442,N_14383);
and U14725 (N_14725,N_14347,N_14340);
or U14726 (N_14726,N_14291,N_14342);
or U14727 (N_14727,N_14300,N_14372);
or U14728 (N_14728,N_14409,N_14412);
or U14729 (N_14729,N_14375,N_14374);
and U14730 (N_14730,N_14359,N_14320);
nor U14731 (N_14731,N_14303,N_14438);
and U14732 (N_14732,N_14463,N_14393);
nand U14733 (N_14733,N_14296,N_14283);
nor U14734 (N_14734,N_14393,N_14409);
or U14735 (N_14735,N_14419,N_14329);
xnor U14736 (N_14736,N_14382,N_14485);
or U14737 (N_14737,N_14274,N_14400);
or U14738 (N_14738,N_14371,N_14476);
or U14739 (N_14739,N_14348,N_14451);
nor U14740 (N_14740,N_14251,N_14479);
nor U14741 (N_14741,N_14458,N_14326);
and U14742 (N_14742,N_14374,N_14421);
xor U14743 (N_14743,N_14251,N_14330);
or U14744 (N_14744,N_14416,N_14471);
nor U14745 (N_14745,N_14402,N_14416);
and U14746 (N_14746,N_14470,N_14390);
and U14747 (N_14747,N_14275,N_14374);
nor U14748 (N_14748,N_14433,N_14439);
nand U14749 (N_14749,N_14391,N_14308);
nor U14750 (N_14750,N_14722,N_14572);
nand U14751 (N_14751,N_14670,N_14749);
or U14752 (N_14752,N_14720,N_14564);
xor U14753 (N_14753,N_14519,N_14625);
xnor U14754 (N_14754,N_14695,N_14736);
nor U14755 (N_14755,N_14568,N_14712);
nor U14756 (N_14756,N_14616,N_14643);
nand U14757 (N_14757,N_14733,N_14567);
nand U14758 (N_14758,N_14613,N_14558);
xnor U14759 (N_14759,N_14543,N_14660);
nand U14760 (N_14760,N_14620,N_14619);
xnor U14761 (N_14761,N_14718,N_14627);
nor U14762 (N_14762,N_14688,N_14582);
and U14763 (N_14763,N_14632,N_14601);
or U14764 (N_14764,N_14645,N_14525);
and U14765 (N_14765,N_14624,N_14524);
nor U14766 (N_14766,N_14500,N_14520);
and U14767 (N_14767,N_14518,N_14631);
nand U14768 (N_14768,N_14596,N_14679);
xor U14769 (N_14769,N_14605,N_14606);
and U14770 (N_14770,N_14553,N_14581);
or U14771 (N_14771,N_14686,N_14570);
xnor U14772 (N_14772,N_14717,N_14549);
nor U14773 (N_14773,N_14653,N_14563);
nor U14774 (N_14774,N_14639,N_14650);
and U14775 (N_14775,N_14589,N_14710);
and U14776 (N_14776,N_14723,N_14566);
or U14777 (N_14777,N_14622,N_14742);
and U14778 (N_14778,N_14636,N_14647);
nor U14779 (N_14779,N_14635,N_14740);
xor U14780 (N_14780,N_14552,N_14547);
nor U14781 (N_14781,N_14676,N_14732);
xnor U14782 (N_14782,N_14593,N_14548);
nor U14783 (N_14783,N_14697,N_14687);
or U14784 (N_14784,N_14557,N_14704);
nor U14785 (N_14785,N_14554,N_14578);
nor U14786 (N_14786,N_14611,N_14725);
or U14787 (N_14787,N_14692,N_14514);
and U14788 (N_14788,N_14661,N_14538);
nand U14789 (N_14789,N_14745,N_14714);
or U14790 (N_14790,N_14560,N_14509);
nand U14791 (N_14791,N_14516,N_14609);
or U14792 (N_14792,N_14556,N_14706);
nand U14793 (N_14793,N_14536,N_14668);
nor U14794 (N_14794,N_14671,N_14565);
xor U14795 (N_14795,N_14610,N_14672);
xor U14796 (N_14796,N_14727,N_14708);
xor U14797 (N_14797,N_14510,N_14511);
and U14798 (N_14798,N_14662,N_14642);
nor U14799 (N_14799,N_14512,N_14615);
xor U14800 (N_14800,N_14654,N_14598);
nor U14801 (N_14801,N_14637,N_14734);
nand U14802 (N_14802,N_14562,N_14646);
and U14803 (N_14803,N_14731,N_14663);
nor U14804 (N_14804,N_14729,N_14638);
nand U14805 (N_14805,N_14588,N_14528);
nand U14806 (N_14806,N_14630,N_14621);
xor U14807 (N_14807,N_14701,N_14657);
nor U14808 (N_14808,N_14623,N_14537);
nor U14809 (N_14809,N_14575,N_14644);
and U14810 (N_14810,N_14608,N_14721);
or U14811 (N_14811,N_14684,N_14693);
nor U14812 (N_14812,N_14594,N_14705);
xnor U14813 (N_14813,N_14612,N_14571);
or U14814 (N_14814,N_14689,N_14604);
nor U14815 (N_14815,N_14651,N_14599);
or U14816 (N_14816,N_14685,N_14585);
or U14817 (N_14817,N_14741,N_14673);
and U14818 (N_14818,N_14590,N_14664);
nand U14819 (N_14819,N_14707,N_14675);
nor U14820 (N_14820,N_14607,N_14517);
and U14821 (N_14821,N_14711,N_14600);
nor U14822 (N_14822,N_14534,N_14529);
nor U14823 (N_14823,N_14658,N_14559);
nand U14824 (N_14824,N_14508,N_14713);
nand U14825 (N_14825,N_14505,N_14503);
and U14826 (N_14826,N_14592,N_14730);
nor U14827 (N_14827,N_14545,N_14602);
nand U14828 (N_14828,N_14540,N_14738);
and U14829 (N_14829,N_14546,N_14580);
xnor U14830 (N_14830,N_14587,N_14649);
nand U14831 (N_14831,N_14666,N_14515);
and U14832 (N_14832,N_14677,N_14641);
nand U14833 (N_14833,N_14735,N_14678);
or U14834 (N_14834,N_14655,N_14682);
nand U14835 (N_14835,N_14542,N_14665);
and U14836 (N_14836,N_14586,N_14617);
and U14837 (N_14837,N_14577,N_14696);
xor U14838 (N_14838,N_14699,N_14522);
or U14839 (N_14839,N_14691,N_14541);
or U14840 (N_14840,N_14523,N_14539);
and U14841 (N_14841,N_14561,N_14573);
and U14842 (N_14842,N_14583,N_14614);
nor U14843 (N_14843,N_14555,N_14640);
nand U14844 (N_14844,N_14648,N_14504);
nor U14845 (N_14845,N_14702,N_14501);
or U14846 (N_14846,N_14674,N_14719);
and U14847 (N_14847,N_14737,N_14739);
xnor U14848 (N_14848,N_14574,N_14634);
and U14849 (N_14849,N_14579,N_14629);
and U14850 (N_14850,N_14506,N_14703);
and U14851 (N_14851,N_14544,N_14507);
or U14852 (N_14852,N_14533,N_14680);
nand U14853 (N_14853,N_14633,N_14597);
xor U14854 (N_14854,N_14716,N_14527);
xnor U14855 (N_14855,N_14550,N_14532);
nor U14856 (N_14856,N_14683,N_14748);
nor U14857 (N_14857,N_14569,N_14698);
nor U14858 (N_14858,N_14628,N_14694);
nor U14859 (N_14859,N_14530,N_14743);
xnor U14860 (N_14860,N_14513,N_14521);
nand U14861 (N_14861,N_14744,N_14656);
xnor U14862 (N_14862,N_14709,N_14576);
and U14863 (N_14863,N_14584,N_14591);
nor U14864 (N_14864,N_14502,N_14603);
nand U14865 (N_14865,N_14746,N_14595);
and U14866 (N_14866,N_14728,N_14700);
nor U14867 (N_14867,N_14531,N_14526);
and U14868 (N_14868,N_14659,N_14724);
and U14869 (N_14869,N_14669,N_14690);
nor U14870 (N_14870,N_14618,N_14681);
and U14871 (N_14871,N_14535,N_14747);
nor U14872 (N_14872,N_14551,N_14652);
xor U14873 (N_14873,N_14726,N_14626);
and U14874 (N_14874,N_14667,N_14715);
nor U14875 (N_14875,N_14598,N_14600);
nor U14876 (N_14876,N_14582,N_14567);
or U14877 (N_14877,N_14710,N_14622);
or U14878 (N_14878,N_14643,N_14627);
xnor U14879 (N_14879,N_14537,N_14659);
or U14880 (N_14880,N_14529,N_14721);
and U14881 (N_14881,N_14727,N_14688);
nor U14882 (N_14882,N_14597,N_14628);
or U14883 (N_14883,N_14590,N_14562);
nand U14884 (N_14884,N_14654,N_14579);
or U14885 (N_14885,N_14664,N_14673);
and U14886 (N_14886,N_14608,N_14527);
nand U14887 (N_14887,N_14526,N_14608);
xnor U14888 (N_14888,N_14587,N_14664);
nand U14889 (N_14889,N_14721,N_14694);
nor U14890 (N_14890,N_14724,N_14701);
nand U14891 (N_14891,N_14668,N_14501);
nand U14892 (N_14892,N_14683,N_14516);
xor U14893 (N_14893,N_14671,N_14531);
and U14894 (N_14894,N_14678,N_14690);
nand U14895 (N_14895,N_14548,N_14572);
or U14896 (N_14896,N_14708,N_14530);
or U14897 (N_14897,N_14613,N_14505);
nand U14898 (N_14898,N_14666,N_14733);
or U14899 (N_14899,N_14588,N_14514);
xor U14900 (N_14900,N_14569,N_14689);
xor U14901 (N_14901,N_14664,N_14504);
nand U14902 (N_14902,N_14733,N_14618);
nand U14903 (N_14903,N_14500,N_14678);
or U14904 (N_14904,N_14697,N_14540);
or U14905 (N_14905,N_14604,N_14568);
nor U14906 (N_14906,N_14522,N_14573);
or U14907 (N_14907,N_14615,N_14651);
nor U14908 (N_14908,N_14656,N_14625);
nor U14909 (N_14909,N_14725,N_14628);
nor U14910 (N_14910,N_14554,N_14583);
nand U14911 (N_14911,N_14730,N_14673);
nor U14912 (N_14912,N_14586,N_14612);
or U14913 (N_14913,N_14720,N_14584);
or U14914 (N_14914,N_14615,N_14515);
or U14915 (N_14915,N_14717,N_14696);
nand U14916 (N_14916,N_14533,N_14739);
and U14917 (N_14917,N_14516,N_14534);
nor U14918 (N_14918,N_14652,N_14558);
or U14919 (N_14919,N_14584,N_14747);
nor U14920 (N_14920,N_14645,N_14562);
nor U14921 (N_14921,N_14648,N_14616);
nor U14922 (N_14922,N_14698,N_14682);
xor U14923 (N_14923,N_14621,N_14743);
xor U14924 (N_14924,N_14534,N_14668);
and U14925 (N_14925,N_14617,N_14548);
and U14926 (N_14926,N_14719,N_14652);
xnor U14927 (N_14927,N_14652,N_14554);
and U14928 (N_14928,N_14616,N_14546);
nand U14929 (N_14929,N_14623,N_14515);
nor U14930 (N_14930,N_14722,N_14664);
or U14931 (N_14931,N_14578,N_14513);
nor U14932 (N_14932,N_14616,N_14529);
xnor U14933 (N_14933,N_14543,N_14608);
and U14934 (N_14934,N_14560,N_14528);
nand U14935 (N_14935,N_14507,N_14698);
or U14936 (N_14936,N_14554,N_14597);
xnor U14937 (N_14937,N_14739,N_14744);
nor U14938 (N_14938,N_14749,N_14741);
or U14939 (N_14939,N_14519,N_14671);
xnor U14940 (N_14940,N_14660,N_14625);
nor U14941 (N_14941,N_14686,N_14618);
or U14942 (N_14942,N_14699,N_14674);
and U14943 (N_14943,N_14523,N_14673);
and U14944 (N_14944,N_14675,N_14588);
or U14945 (N_14945,N_14618,N_14517);
nand U14946 (N_14946,N_14577,N_14507);
or U14947 (N_14947,N_14577,N_14724);
or U14948 (N_14948,N_14538,N_14734);
xor U14949 (N_14949,N_14605,N_14709);
and U14950 (N_14950,N_14637,N_14538);
or U14951 (N_14951,N_14510,N_14585);
xor U14952 (N_14952,N_14715,N_14676);
nand U14953 (N_14953,N_14551,N_14555);
xnor U14954 (N_14954,N_14567,N_14601);
and U14955 (N_14955,N_14537,N_14641);
nand U14956 (N_14956,N_14583,N_14720);
or U14957 (N_14957,N_14747,N_14675);
nand U14958 (N_14958,N_14648,N_14682);
xor U14959 (N_14959,N_14633,N_14695);
xor U14960 (N_14960,N_14540,N_14598);
and U14961 (N_14961,N_14557,N_14581);
nor U14962 (N_14962,N_14508,N_14576);
or U14963 (N_14963,N_14700,N_14663);
nand U14964 (N_14964,N_14661,N_14726);
xnor U14965 (N_14965,N_14534,N_14607);
xor U14966 (N_14966,N_14725,N_14683);
and U14967 (N_14967,N_14691,N_14593);
or U14968 (N_14968,N_14622,N_14537);
or U14969 (N_14969,N_14526,N_14535);
and U14970 (N_14970,N_14683,N_14656);
nor U14971 (N_14971,N_14669,N_14644);
nand U14972 (N_14972,N_14622,N_14684);
nand U14973 (N_14973,N_14727,N_14512);
nand U14974 (N_14974,N_14513,N_14717);
or U14975 (N_14975,N_14565,N_14743);
and U14976 (N_14976,N_14707,N_14609);
nor U14977 (N_14977,N_14721,N_14688);
nand U14978 (N_14978,N_14570,N_14534);
nand U14979 (N_14979,N_14649,N_14596);
nand U14980 (N_14980,N_14573,N_14517);
xor U14981 (N_14981,N_14621,N_14508);
nand U14982 (N_14982,N_14542,N_14537);
nor U14983 (N_14983,N_14733,N_14668);
xnor U14984 (N_14984,N_14652,N_14724);
xor U14985 (N_14985,N_14543,N_14531);
xor U14986 (N_14986,N_14565,N_14526);
nor U14987 (N_14987,N_14719,N_14684);
or U14988 (N_14988,N_14664,N_14597);
xnor U14989 (N_14989,N_14597,N_14552);
and U14990 (N_14990,N_14705,N_14718);
nor U14991 (N_14991,N_14748,N_14650);
and U14992 (N_14992,N_14519,N_14539);
xnor U14993 (N_14993,N_14697,N_14685);
or U14994 (N_14994,N_14575,N_14525);
nor U14995 (N_14995,N_14568,N_14589);
nor U14996 (N_14996,N_14745,N_14660);
or U14997 (N_14997,N_14523,N_14571);
or U14998 (N_14998,N_14573,N_14553);
nand U14999 (N_14999,N_14654,N_14707);
nand U15000 (N_15000,N_14947,N_14810);
nand U15001 (N_15001,N_14765,N_14866);
and U15002 (N_15002,N_14987,N_14753);
nor U15003 (N_15003,N_14931,N_14876);
nand U15004 (N_15004,N_14760,N_14880);
xor U15005 (N_15005,N_14871,N_14813);
or U15006 (N_15006,N_14892,N_14878);
nand U15007 (N_15007,N_14982,N_14814);
xor U15008 (N_15008,N_14988,N_14824);
xor U15009 (N_15009,N_14903,N_14833);
or U15010 (N_15010,N_14811,N_14963);
or U15011 (N_15011,N_14964,N_14948);
nand U15012 (N_15012,N_14972,N_14818);
or U15013 (N_15013,N_14804,N_14795);
and U15014 (N_15014,N_14797,N_14845);
nor U15015 (N_15015,N_14999,N_14887);
nor U15016 (N_15016,N_14959,N_14904);
and U15017 (N_15017,N_14957,N_14994);
and U15018 (N_15018,N_14942,N_14946);
nand U15019 (N_15019,N_14862,N_14874);
nor U15020 (N_15020,N_14756,N_14881);
or U15021 (N_15021,N_14956,N_14897);
nand U15022 (N_15022,N_14925,N_14981);
and U15023 (N_15023,N_14846,N_14825);
nor U15024 (N_15024,N_14870,N_14777);
or U15025 (N_15025,N_14997,N_14858);
or U15026 (N_15026,N_14784,N_14754);
xor U15027 (N_15027,N_14791,N_14782);
and U15028 (N_15028,N_14940,N_14938);
and U15029 (N_15029,N_14960,N_14885);
or U15030 (N_15030,N_14884,N_14785);
nand U15031 (N_15031,N_14879,N_14776);
nand U15032 (N_15032,N_14848,N_14816);
nand U15033 (N_15033,N_14886,N_14829);
and U15034 (N_15034,N_14830,N_14986);
and U15035 (N_15035,N_14826,N_14828);
or U15036 (N_15036,N_14869,N_14751);
and U15037 (N_15037,N_14872,N_14775);
nor U15038 (N_15038,N_14928,N_14930);
xor U15039 (N_15039,N_14953,N_14805);
nand U15040 (N_15040,N_14801,N_14839);
or U15041 (N_15041,N_14958,N_14978);
and U15042 (N_15042,N_14841,N_14757);
and U15043 (N_15043,N_14853,N_14922);
nor U15044 (N_15044,N_14888,N_14821);
nand U15045 (N_15045,N_14789,N_14819);
nor U15046 (N_15046,N_14788,N_14900);
and U15047 (N_15047,N_14771,N_14979);
nor U15048 (N_15048,N_14950,N_14837);
nand U15049 (N_15049,N_14995,N_14923);
or U15050 (N_15050,N_14914,N_14926);
nand U15051 (N_15051,N_14889,N_14907);
xor U15052 (N_15052,N_14913,N_14910);
xnor U15053 (N_15053,N_14792,N_14898);
nor U15054 (N_15054,N_14967,N_14865);
nor U15055 (N_15055,N_14807,N_14762);
nor U15056 (N_15056,N_14873,N_14920);
and U15057 (N_15057,N_14779,N_14932);
nand U15058 (N_15058,N_14750,N_14875);
nor U15059 (N_15059,N_14850,N_14847);
or U15060 (N_15060,N_14844,N_14970);
or U15061 (N_15061,N_14935,N_14838);
xnor U15062 (N_15062,N_14803,N_14780);
and U15063 (N_15063,N_14835,N_14796);
nor U15064 (N_15064,N_14759,N_14790);
xnor U15065 (N_15065,N_14993,N_14998);
nor U15066 (N_15066,N_14962,N_14961);
and U15067 (N_15067,N_14919,N_14764);
xnor U15068 (N_15068,N_14768,N_14868);
nand U15069 (N_15069,N_14799,N_14894);
nor U15070 (N_15070,N_14831,N_14761);
nor U15071 (N_15071,N_14895,N_14763);
xor U15072 (N_15072,N_14990,N_14849);
xnor U15073 (N_15073,N_14783,N_14980);
nor U15074 (N_15074,N_14944,N_14859);
nor U15075 (N_15075,N_14773,N_14798);
nor U15076 (N_15076,N_14854,N_14933);
xor U15077 (N_15077,N_14808,N_14971);
xnor U15078 (N_15078,N_14817,N_14815);
nor U15079 (N_15079,N_14857,N_14832);
and U15080 (N_15080,N_14916,N_14812);
nor U15081 (N_15081,N_14943,N_14851);
xor U15082 (N_15082,N_14823,N_14758);
or U15083 (N_15083,N_14794,N_14766);
xnor U15084 (N_15084,N_14840,N_14772);
or U15085 (N_15085,N_14767,N_14977);
nand U15086 (N_15086,N_14770,N_14861);
xnor U15087 (N_15087,N_14882,N_14856);
nor U15088 (N_15088,N_14774,N_14852);
nand U15089 (N_15089,N_14806,N_14755);
xnor U15090 (N_15090,N_14929,N_14954);
xnor U15091 (N_15091,N_14842,N_14949);
xor U15092 (N_15092,N_14924,N_14968);
and U15093 (N_15093,N_14905,N_14834);
and U15094 (N_15094,N_14915,N_14951);
nor U15095 (N_15095,N_14996,N_14778);
nor U15096 (N_15096,N_14975,N_14786);
nand U15097 (N_15097,N_14827,N_14867);
or U15098 (N_15098,N_14802,N_14860);
and U15099 (N_15099,N_14941,N_14917);
nand U15100 (N_15100,N_14985,N_14793);
xor U15101 (N_15101,N_14974,N_14965);
nor U15102 (N_15102,N_14787,N_14939);
or U15103 (N_15103,N_14890,N_14800);
or U15104 (N_15104,N_14991,N_14912);
nand U15105 (N_15105,N_14983,N_14901);
nor U15106 (N_15106,N_14966,N_14936);
or U15107 (N_15107,N_14836,N_14896);
xor U15108 (N_15108,N_14911,N_14822);
nand U15109 (N_15109,N_14937,N_14863);
nor U15110 (N_15110,N_14976,N_14781);
nor U15111 (N_15111,N_14769,N_14952);
xnor U15112 (N_15112,N_14877,N_14945);
or U15113 (N_15113,N_14992,N_14820);
nand U15114 (N_15114,N_14908,N_14984);
and U15115 (N_15115,N_14909,N_14752);
nand U15116 (N_15116,N_14891,N_14955);
and U15117 (N_15117,N_14969,N_14899);
and U15118 (N_15118,N_14918,N_14883);
nand U15119 (N_15119,N_14906,N_14927);
and U15120 (N_15120,N_14893,N_14855);
and U15121 (N_15121,N_14809,N_14934);
xnor U15122 (N_15122,N_14902,N_14864);
xor U15123 (N_15123,N_14989,N_14843);
xor U15124 (N_15124,N_14921,N_14973);
or U15125 (N_15125,N_14981,N_14771);
nand U15126 (N_15126,N_14888,N_14857);
or U15127 (N_15127,N_14795,N_14939);
nor U15128 (N_15128,N_14790,N_14811);
and U15129 (N_15129,N_14779,N_14964);
nor U15130 (N_15130,N_14861,N_14896);
nor U15131 (N_15131,N_14795,N_14821);
nand U15132 (N_15132,N_14827,N_14947);
and U15133 (N_15133,N_14956,N_14772);
nor U15134 (N_15134,N_14846,N_14954);
nand U15135 (N_15135,N_14810,N_14939);
nand U15136 (N_15136,N_14937,N_14861);
or U15137 (N_15137,N_14968,N_14993);
or U15138 (N_15138,N_14831,N_14935);
nand U15139 (N_15139,N_14841,N_14839);
or U15140 (N_15140,N_14820,N_14859);
nand U15141 (N_15141,N_14757,N_14872);
nor U15142 (N_15142,N_14977,N_14876);
or U15143 (N_15143,N_14778,N_14905);
xor U15144 (N_15144,N_14843,N_14927);
and U15145 (N_15145,N_14884,N_14818);
nand U15146 (N_15146,N_14844,N_14988);
nand U15147 (N_15147,N_14972,N_14807);
and U15148 (N_15148,N_14845,N_14907);
or U15149 (N_15149,N_14924,N_14912);
and U15150 (N_15150,N_14948,N_14988);
xor U15151 (N_15151,N_14756,N_14785);
nand U15152 (N_15152,N_14833,N_14800);
and U15153 (N_15153,N_14770,N_14862);
nand U15154 (N_15154,N_14801,N_14937);
nor U15155 (N_15155,N_14796,N_14816);
or U15156 (N_15156,N_14823,N_14806);
nand U15157 (N_15157,N_14837,N_14912);
xor U15158 (N_15158,N_14830,N_14909);
nor U15159 (N_15159,N_14896,N_14860);
xnor U15160 (N_15160,N_14865,N_14764);
nor U15161 (N_15161,N_14769,N_14829);
and U15162 (N_15162,N_14935,N_14883);
nand U15163 (N_15163,N_14953,N_14846);
or U15164 (N_15164,N_14963,N_14961);
xnor U15165 (N_15165,N_14970,N_14918);
nor U15166 (N_15166,N_14981,N_14923);
and U15167 (N_15167,N_14906,N_14845);
xnor U15168 (N_15168,N_14902,N_14994);
and U15169 (N_15169,N_14770,N_14961);
and U15170 (N_15170,N_14765,N_14798);
xor U15171 (N_15171,N_14794,N_14777);
and U15172 (N_15172,N_14922,N_14846);
nor U15173 (N_15173,N_14823,N_14944);
or U15174 (N_15174,N_14923,N_14855);
nor U15175 (N_15175,N_14797,N_14994);
nand U15176 (N_15176,N_14879,N_14853);
xor U15177 (N_15177,N_14831,N_14947);
or U15178 (N_15178,N_14790,N_14965);
nor U15179 (N_15179,N_14758,N_14799);
or U15180 (N_15180,N_14934,N_14823);
or U15181 (N_15181,N_14992,N_14942);
nand U15182 (N_15182,N_14998,N_14859);
nand U15183 (N_15183,N_14928,N_14884);
nor U15184 (N_15184,N_14919,N_14779);
nor U15185 (N_15185,N_14808,N_14822);
nand U15186 (N_15186,N_14963,N_14799);
or U15187 (N_15187,N_14912,N_14868);
and U15188 (N_15188,N_14907,N_14934);
nand U15189 (N_15189,N_14801,N_14930);
or U15190 (N_15190,N_14807,N_14914);
nor U15191 (N_15191,N_14797,N_14895);
nand U15192 (N_15192,N_14823,N_14876);
and U15193 (N_15193,N_14816,N_14754);
nor U15194 (N_15194,N_14968,N_14783);
nor U15195 (N_15195,N_14953,N_14893);
xor U15196 (N_15196,N_14856,N_14871);
nand U15197 (N_15197,N_14942,N_14913);
or U15198 (N_15198,N_14832,N_14806);
nor U15199 (N_15199,N_14810,N_14856);
and U15200 (N_15200,N_14825,N_14909);
nand U15201 (N_15201,N_14779,N_14996);
nor U15202 (N_15202,N_14856,N_14763);
nand U15203 (N_15203,N_14875,N_14946);
nand U15204 (N_15204,N_14911,N_14756);
nor U15205 (N_15205,N_14980,N_14757);
nor U15206 (N_15206,N_14946,N_14800);
nor U15207 (N_15207,N_14998,N_14894);
xor U15208 (N_15208,N_14775,N_14905);
xor U15209 (N_15209,N_14861,N_14753);
or U15210 (N_15210,N_14927,N_14907);
nand U15211 (N_15211,N_14751,N_14793);
or U15212 (N_15212,N_14961,N_14888);
and U15213 (N_15213,N_14988,N_14782);
xnor U15214 (N_15214,N_14853,N_14898);
nor U15215 (N_15215,N_14907,N_14911);
or U15216 (N_15216,N_14897,N_14934);
and U15217 (N_15217,N_14956,N_14763);
nand U15218 (N_15218,N_14966,N_14845);
or U15219 (N_15219,N_14899,N_14987);
and U15220 (N_15220,N_14896,N_14945);
or U15221 (N_15221,N_14907,N_14827);
and U15222 (N_15222,N_14840,N_14831);
nand U15223 (N_15223,N_14794,N_14775);
xnor U15224 (N_15224,N_14816,N_14788);
or U15225 (N_15225,N_14837,N_14926);
and U15226 (N_15226,N_14925,N_14784);
nand U15227 (N_15227,N_14880,N_14779);
xnor U15228 (N_15228,N_14820,N_14928);
xnor U15229 (N_15229,N_14854,N_14844);
and U15230 (N_15230,N_14853,N_14924);
and U15231 (N_15231,N_14856,N_14863);
and U15232 (N_15232,N_14752,N_14844);
xnor U15233 (N_15233,N_14901,N_14900);
xnor U15234 (N_15234,N_14844,N_14782);
xnor U15235 (N_15235,N_14953,N_14820);
nor U15236 (N_15236,N_14895,N_14875);
nor U15237 (N_15237,N_14956,N_14979);
or U15238 (N_15238,N_14921,N_14761);
and U15239 (N_15239,N_14791,N_14960);
or U15240 (N_15240,N_14825,N_14924);
or U15241 (N_15241,N_14993,N_14992);
xnor U15242 (N_15242,N_14778,N_14903);
xnor U15243 (N_15243,N_14944,N_14896);
nor U15244 (N_15244,N_14795,N_14955);
and U15245 (N_15245,N_14932,N_14900);
nand U15246 (N_15246,N_14797,N_14767);
nor U15247 (N_15247,N_14969,N_14832);
nand U15248 (N_15248,N_14761,N_14983);
nand U15249 (N_15249,N_14865,N_14830);
nor U15250 (N_15250,N_15220,N_15233);
or U15251 (N_15251,N_15105,N_15123);
xor U15252 (N_15252,N_15031,N_15141);
and U15253 (N_15253,N_15111,N_15249);
and U15254 (N_15254,N_15160,N_15051);
nor U15255 (N_15255,N_15043,N_15113);
xnor U15256 (N_15256,N_15029,N_15005);
nand U15257 (N_15257,N_15138,N_15247);
and U15258 (N_15258,N_15140,N_15144);
or U15259 (N_15259,N_15053,N_15107);
xnor U15260 (N_15260,N_15042,N_15012);
and U15261 (N_15261,N_15061,N_15040);
nor U15262 (N_15262,N_15095,N_15030);
or U15263 (N_15263,N_15189,N_15203);
xor U15264 (N_15264,N_15121,N_15198);
or U15265 (N_15265,N_15013,N_15208);
xnor U15266 (N_15266,N_15148,N_15245);
or U15267 (N_15267,N_15163,N_15204);
nand U15268 (N_15268,N_15026,N_15136);
nand U15269 (N_15269,N_15178,N_15210);
and U15270 (N_15270,N_15033,N_15060);
and U15271 (N_15271,N_15032,N_15096);
nand U15272 (N_15272,N_15244,N_15122);
and U15273 (N_15273,N_15231,N_15175);
xnor U15274 (N_15274,N_15084,N_15226);
nand U15275 (N_15275,N_15248,N_15078);
nor U15276 (N_15276,N_15024,N_15117);
nor U15277 (N_15277,N_15213,N_15212);
nand U15278 (N_15278,N_15080,N_15237);
and U15279 (N_15279,N_15034,N_15156);
or U15280 (N_15280,N_15018,N_15225);
or U15281 (N_15281,N_15015,N_15159);
xnor U15282 (N_15282,N_15151,N_15157);
or U15283 (N_15283,N_15194,N_15181);
nand U15284 (N_15284,N_15197,N_15041);
xnor U15285 (N_15285,N_15147,N_15154);
or U15286 (N_15286,N_15008,N_15146);
or U15287 (N_15287,N_15093,N_15073);
nor U15288 (N_15288,N_15118,N_15236);
or U15289 (N_15289,N_15150,N_15007);
xor U15290 (N_15290,N_15082,N_15097);
and U15291 (N_15291,N_15149,N_15223);
nand U15292 (N_15292,N_15172,N_15224);
or U15293 (N_15293,N_15188,N_15038);
nor U15294 (N_15294,N_15011,N_15170);
nor U15295 (N_15295,N_15062,N_15191);
xnor U15296 (N_15296,N_15202,N_15173);
or U15297 (N_15297,N_15109,N_15063);
nor U15298 (N_15298,N_15165,N_15186);
or U15299 (N_15299,N_15081,N_15099);
and U15300 (N_15300,N_15079,N_15126);
and U15301 (N_15301,N_15166,N_15006);
nand U15302 (N_15302,N_15240,N_15091);
xnor U15303 (N_15303,N_15027,N_15153);
and U15304 (N_15304,N_15075,N_15068);
or U15305 (N_15305,N_15124,N_15211);
and U15306 (N_15306,N_15180,N_15171);
nand U15307 (N_15307,N_15127,N_15025);
nor U15308 (N_15308,N_15137,N_15217);
nor U15309 (N_15309,N_15241,N_15059);
xnor U15310 (N_15310,N_15066,N_15065);
nor U15311 (N_15311,N_15064,N_15047);
nand U15312 (N_15312,N_15087,N_15108);
and U15313 (N_15313,N_15182,N_15021);
and U15314 (N_15314,N_15176,N_15139);
xnor U15315 (N_15315,N_15056,N_15052);
nand U15316 (N_15316,N_15114,N_15207);
xnor U15317 (N_15317,N_15116,N_15243);
xor U15318 (N_15318,N_15106,N_15125);
xor U15319 (N_15319,N_15199,N_15049);
and U15320 (N_15320,N_15179,N_15045);
nand U15321 (N_15321,N_15002,N_15238);
nor U15322 (N_15322,N_15057,N_15094);
or U15323 (N_15323,N_15090,N_15155);
xor U15324 (N_15324,N_15221,N_15129);
nand U15325 (N_15325,N_15169,N_15101);
nand U15326 (N_15326,N_15162,N_15209);
nand U15327 (N_15327,N_15227,N_15077);
nand U15328 (N_15328,N_15201,N_15130);
and U15329 (N_15329,N_15083,N_15067);
or U15330 (N_15330,N_15103,N_15229);
xnor U15331 (N_15331,N_15119,N_15177);
or U15332 (N_15332,N_15164,N_15196);
nor U15333 (N_15333,N_15192,N_15016);
and U15334 (N_15334,N_15086,N_15216);
nor U15335 (N_15335,N_15167,N_15133);
or U15336 (N_15336,N_15131,N_15037);
or U15337 (N_15337,N_15023,N_15168);
xor U15338 (N_15338,N_15242,N_15036);
xnor U15339 (N_15339,N_15158,N_15035);
nor U15340 (N_15340,N_15054,N_15050);
and U15341 (N_15341,N_15115,N_15152);
and U15342 (N_15342,N_15222,N_15058);
xor U15343 (N_15343,N_15074,N_15219);
and U15344 (N_15344,N_15184,N_15234);
and U15345 (N_15345,N_15132,N_15142);
or U15346 (N_15346,N_15104,N_15190);
nand U15347 (N_15347,N_15000,N_15088);
nand U15348 (N_15348,N_15183,N_15102);
nand U15349 (N_15349,N_15112,N_15001);
or U15350 (N_15350,N_15143,N_15218);
nor U15351 (N_15351,N_15174,N_15230);
or U15352 (N_15352,N_15246,N_15200);
xnor U15353 (N_15353,N_15135,N_15003);
xnor U15354 (N_15354,N_15044,N_15134);
nor U15355 (N_15355,N_15009,N_15206);
nor U15356 (N_15356,N_15070,N_15092);
nor U15357 (N_15357,N_15017,N_15185);
or U15358 (N_15358,N_15071,N_15214);
nor U15359 (N_15359,N_15193,N_15039);
xnor U15360 (N_15360,N_15076,N_15069);
xor U15361 (N_15361,N_15014,N_15089);
and U15362 (N_15362,N_15195,N_15120);
nor U15363 (N_15363,N_15055,N_15239);
and U15364 (N_15364,N_15128,N_15019);
nor U15365 (N_15365,N_15010,N_15228);
or U15366 (N_15366,N_15187,N_15046);
nand U15367 (N_15367,N_15028,N_15048);
or U15368 (N_15368,N_15085,N_15161);
nor U15369 (N_15369,N_15072,N_15145);
and U15370 (N_15370,N_15100,N_15235);
nand U15371 (N_15371,N_15232,N_15215);
xor U15372 (N_15372,N_15004,N_15110);
and U15373 (N_15373,N_15205,N_15022);
nor U15374 (N_15374,N_15098,N_15020);
nand U15375 (N_15375,N_15136,N_15104);
and U15376 (N_15376,N_15158,N_15034);
and U15377 (N_15377,N_15109,N_15235);
or U15378 (N_15378,N_15128,N_15144);
xnor U15379 (N_15379,N_15053,N_15159);
xor U15380 (N_15380,N_15010,N_15056);
or U15381 (N_15381,N_15220,N_15227);
xor U15382 (N_15382,N_15027,N_15178);
nor U15383 (N_15383,N_15247,N_15192);
xor U15384 (N_15384,N_15085,N_15014);
and U15385 (N_15385,N_15242,N_15009);
or U15386 (N_15386,N_15069,N_15241);
and U15387 (N_15387,N_15053,N_15015);
nor U15388 (N_15388,N_15083,N_15114);
or U15389 (N_15389,N_15066,N_15053);
and U15390 (N_15390,N_15211,N_15017);
and U15391 (N_15391,N_15216,N_15138);
or U15392 (N_15392,N_15063,N_15180);
xor U15393 (N_15393,N_15069,N_15122);
nand U15394 (N_15394,N_15140,N_15194);
nor U15395 (N_15395,N_15055,N_15187);
xnor U15396 (N_15396,N_15104,N_15096);
or U15397 (N_15397,N_15247,N_15069);
and U15398 (N_15398,N_15200,N_15169);
xor U15399 (N_15399,N_15201,N_15116);
nor U15400 (N_15400,N_15112,N_15046);
or U15401 (N_15401,N_15194,N_15040);
or U15402 (N_15402,N_15132,N_15218);
nor U15403 (N_15403,N_15147,N_15043);
and U15404 (N_15404,N_15062,N_15018);
and U15405 (N_15405,N_15117,N_15111);
nor U15406 (N_15406,N_15014,N_15142);
nand U15407 (N_15407,N_15113,N_15015);
xor U15408 (N_15408,N_15028,N_15243);
nor U15409 (N_15409,N_15022,N_15019);
nor U15410 (N_15410,N_15165,N_15214);
nand U15411 (N_15411,N_15058,N_15078);
and U15412 (N_15412,N_15189,N_15186);
or U15413 (N_15413,N_15047,N_15053);
nand U15414 (N_15414,N_15107,N_15105);
nand U15415 (N_15415,N_15009,N_15073);
or U15416 (N_15416,N_15081,N_15044);
xor U15417 (N_15417,N_15041,N_15011);
or U15418 (N_15418,N_15002,N_15055);
xor U15419 (N_15419,N_15054,N_15195);
and U15420 (N_15420,N_15094,N_15109);
nor U15421 (N_15421,N_15054,N_15247);
and U15422 (N_15422,N_15088,N_15092);
xnor U15423 (N_15423,N_15044,N_15169);
nor U15424 (N_15424,N_15070,N_15145);
and U15425 (N_15425,N_15057,N_15231);
and U15426 (N_15426,N_15083,N_15155);
and U15427 (N_15427,N_15144,N_15050);
nor U15428 (N_15428,N_15061,N_15172);
nor U15429 (N_15429,N_15177,N_15212);
nand U15430 (N_15430,N_15084,N_15179);
or U15431 (N_15431,N_15013,N_15016);
nor U15432 (N_15432,N_15135,N_15089);
nand U15433 (N_15433,N_15149,N_15238);
or U15434 (N_15434,N_15106,N_15085);
or U15435 (N_15435,N_15034,N_15041);
or U15436 (N_15436,N_15118,N_15237);
xor U15437 (N_15437,N_15088,N_15127);
nand U15438 (N_15438,N_15154,N_15101);
xnor U15439 (N_15439,N_15239,N_15214);
nand U15440 (N_15440,N_15032,N_15027);
and U15441 (N_15441,N_15162,N_15201);
or U15442 (N_15442,N_15187,N_15224);
xnor U15443 (N_15443,N_15116,N_15162);
and U15444 (N_15444,N_15196,N_15015);
nand U15445 (N_15445,N_15003,N_15128);
and U15446 (N_15446,N_15168,N_15225);
nor U15447 (N_15447,N_15078,N_15175);
or U15448 (N_15448,N_15228,N_15035);
and U15449 (N_15449,N_15005,N_15055);
nand U15450 (N_15450,N_15119,N_15224);
nand U15451 (N_15451,N_15105,N_15116);
or U15452 (N_15452,N_15236,N_15205);
xnor U15453 (N_15453,N_15121,N_15004);
nand U15454 (N_15454,N_15149,N_15192);
or U15455 (N_15455,N_15198,N_15184);
xnor U15456 (N_15456,N_15225,N_15088);
or U15457 (N_15457,N_15237,N_15207);
xnor U15458 (N_15458,N_15028,N_15167);
nand U15459 (N_15459,N_15179,N_15203);
and U15460 (N_15460,N_15234,N_15193);
nand U15461 (N_15461,N_15109,N_15032);
nor U15462 (N_15462,N_15193,N_15015);
and U15463 (N_15463,N_15001,N_15079);
and U15464 (N_15464,N_15077,N_15087);
or U15465 (N_15465,N_15201,N_15037);
nor U15466 (N_15466,N_15155,N_15085);
nand U15467 (N_15467,N_15010,N_15006);
nor U15468 (N_15468,N_15213,N_15121);
and U15469 (N_15469,N_15065,N_15038);
and U15470 (N_15470,N_15249,N_15099);
and U15471 (N_15471,N_15185,N_15090);
nor U15472 (N_15472,N_15065,N_15027);
xnor U15473 (N_15473,N_15023,N_15242);
nor U15474 (N_15474,N_15003,N_15241);
and U15475 (N_15475,N_15044,N_15159);
xnor U15476 (N_15476,N_15143,N_15095);
xor U15477 (N_15477,N_15027,N_15173);
xnor U15478 (N_15478,N_15101,N_15129);
xnor U15479 (N_15479,N_15181,N_15225);
nor U15480 (N_15480,N_15183,N_15178);
nor U15481 (N_15481,N_15079,N_15178);
xnor U15482 (N_15482,N_15026,N_15183);
nand U15483 (N_15483,N_15100,N_15106);
or U15484 (N_15484,N_15205,N_15157);
nand U15485 (N_15485,N_15220,N_15186);
xnor U15486 (N_15486,N_15141,N_15238);
or U15487 (N_15487,N_15010,N_15115);
or U15488 (N_15488,N_15173,N_15138);
xnor U15489 (N_15489,N_15210,N_15175);
or U15490 (N_15490,N_15180,N_15106);
or U15491 (N_15491,N_15151,N_15229);
nand U15492 (N_15492,N_15051,N_15026);
and U15493 (N_15493,N_15171,N_15024);
or U15494 (N_15494,N_15174,N_15009);
or U15495 (N_15495,N_15148,N_15019);
or U15496 (N_15496,N_15244,N_15019);
and U15497 (N_15497,N_15102,N_15081);
and U15498 (N_15498,N_15005,N_15203);
and U15499 (N_15499,N_15067,N_15149);
and U15500 (N_15500,N_15431,N_15483);
or U15501 (N_15501,N_15450,N_15463);
or U15502 (N_15502,N_15268,N_15347);
or U15503 (N_15503,N_15465,N_15321);
xor U15504 (N_15504,N_15399,N_15289);
xnor U15505 (N_15505,N_15446,N_15477);
and U15506 (N_15506,N_15495,N_15479);
xnor U15507 (N_15507,N_15439,N_15382);
xnor U15508 (N_15508,N_15354,N_15294);
nand U15509 (N_15509,N_15422,N_15389);
and U15510 (N_15510,N_15307,N_15361);
nor U15511 (N_15511,N_15337,N_15468);
nor U15512 (N_15512,N_15310,N_15251);
xnor U15513 (N_15513,N_15488,N_15323);
nor U15514 (N_15514,N_15425,N_15279);
nand U15515 (N_15515,N_15257,N_15408);
xnor U15516 (N_15516,N_15349,N_15386);
or U15517 (N_15517,N_15394,N_15281);
nor U15518 (N_15518,N_15403,N_15442);
and U15519 (N_15519,N_15340,N_15447);
xnor U15520 (N_15520,N_15401,N_15271);
nand U15521 (N_15521,N_15316,N_15493);
nor U15522 (N_15522,N_15381,N_15370);
or U15523 (N_15523,N_15319,N_15306);
and U15524 (N_15524,N_15313,N_15376);
or U15525 (N_15525,N_15464,N_15371);
xnor U15526 (N_15526,N_15411,N_15402);
nand U15527 (N_15527,N_15405,N_15496);
nor U15528 (N_15528,N_15288,N_15482);
nor U15529 (N_15529,N_15259,N_15264);
nand U15530 (N_15530,N_15476,N_15303);
nor U15531 (N_15531,N_15364,N_15322);
nand U15532 (N_15532,N_15406,N_15462);
and U15533 (N_15533,N_15338,N_15404);
xor U15534 (N_15534,N_15395,N_15430);
xor U15535 (N_15535,N_15398,N_15345);
and U15536 (N_15536,N_15481,N_15416);
nor U15537 (N_15537,N_15365,N_15284);
nand U15538 (N_15538,N_15350,N_15261);
nand U15539 (N_15539,N_15419,N_15254);
xor U15540 (N_15540,N_15317,N_15384);
nand U15541 (N_15541,N_15308,N_15418);
nor U15542 (N_15542,N_15454,N_15369);
nand U15543 (N_15543,N_15469,N_15429);
xnor U15544 (N_15544,N_15388,N_15258);
or U15545 (N_15545,N_15285,N_15426);
nor U15546 (N_15546,N_15491,N_15435);
and U15547 (N_15547,N_15353,N_15278);
and U15548 (N_15548,N_15461,N_15359);
or U15549 (N_15549,N_15295,N_15330);
nor U15550 (N_15550,N_15453,N_15357);
nor U15551 (N_15551,N_15383,N_15414);
nand U15552 (N_15552,N_15451,N_15352);
nand U15553 (N_15553,N_15324,N_15390);
or U15554 (N_15554,N_15309,N_15333);
xnor U15555 (N_15555,N_15356,N_15282);
xor U15556 (N_15556,N_15360,N_15328);
nand U15557 (N_15557,N_15253,N_15332);
or U15558 (N_15558,N_15252,N_15343);
and U15559 (N_15559,N_15272,N_15397);
xor U15560 (N_15560,N_15448,N_15470);
or U15561 (N_15561,N_15346,N_15298);
nand U15562 (N_15562,N_15485,N_15291);
or U15563 (N_15563,N_15366,N_15471);
or U15564 (N_15564,N_15250,N_15409);
or U15565 (N_15565,N_15391,N_15262);
and U15566 (N_15566,N_15320,N_15339);
xor U15567 (N_15567,N_15296,N_15396);
xnor U15568 (N_15568,N_15355,N_15270);
nand U15569 (N_15569,N_15457,N_15445);
and U15570 (N_15570,N_15400,N_15276);
or U15571 (N_15571,N_15292,N_15334);
nor U15572 (N_15572,N_15368,N_15379);
and U15573 (N_15573,N_15466,N_15274);
xnor U15574 (N_15574,N_15428,N_15312);
or U15575 (N_15575,N_15331,N_15283);
xor U15576 (N_15576,N_15421,N_15255);
or U15577 (N_15577,N_15437,N_15266);
xor U15578 (N_15578,N_15311,N_15256);
or U15579 (N_15579,N_15275,N_15458);
nor U15580 (N_15580,N_15412,N_15377);
and U15581 (N_15581,N_15325,N_15499);
or U15582 (N_15582,N_15456,N_15287);
or U15583 (N_15583,N_15314,N_15263);
and U15584 (N_15584,N_15489,N_15375);
and U15585 (N_15585,N_15480,N_15304);
nand U15586 (N_15586,N_15392,N_15351);
and U15587 (N_15587,N_15497,N_15486);
xnor U15588 (N_15588,N_15348,N_15424);
nor U15589 (N_15589,N_15452,N_15417);
or U15590 (N_15590,N_15344,N_15433);
nand U15591 (N_15591,N_15380,N_15387);
or U15592 (N_15592,N_15420,N_15478);
and U15593 (N_15593,N_15449,N_15362);
nor U15594 (N_15594,N_15363,N_15441);
or U15595 (N_15595,N_15372,N_15455);
nor U15596 (N_15596,N_15329,N_15293);
nor U15597 (N_15597,N_15413,N_15286);
and U15598 (N_15598,N_15335,N_15280);
and U15599 (N_15599,N_15297,N_15300);
nor U15600 (N_15600,N_15487,N_15277);
xor U15601 (N_15601,N_15438,N_15326);
and U15602 (N_15602,N_15459,N_15367);
nor U15603 (N_15603,N_15494,N_15474);
nand U15604 (N_15604,N_15436,N_15305);
nand U15605 (N_15605,N_15341,N_15327);
xnor U15606 (N_15606,N_15434,N_15336);
or U15607 (N_15607,N_15440,N_15269);
and U15608 (N_15608,N_15315,N_15265);
xnor U15609 (N_15609,N_15498,N_15267);
nor U15610 (N_15610,N_15410,N_15473);
and U15611 (N_15611,N_15472,N_15427);
and U15612 (N_15612,N_15318,N_15385);
nand U15613 (N_15613,N_15415,N_15467);
nand U15614 (N_15614,N_15378,N_15423);
and U15615 (N_15615,N_15393,N_15490);
nand U15616 (N_15616,N_15302,N_15443);
and U15617 (N_15617,N_15299,N_15374);
or U15618 (N_15618,N_15373,N_15290);
nor U15619 (N_15619,N_15460,N_15260);
nand U15620 (N_15620,N_15444,N_15342);
or U15621 (N_15621,N_15301,N_15407);
and U15622 (N_15622,N_15475,N_15484);
and U15623 (N_15623,N_15273,N_15358);
xor U15624 (N_15624,N_15492,N_15432);
or U15625 (N_15625,N_15461,N_15262);
and U15626 (N_15626,N_15355,N_15377);
xnor U15627 (N_15627,N_15350,N_15449);
and U15628 (N_15628,N_15438,N_15354);
nand U15629 (N_15629,N_15325,N_15479);
and U15630 (N_15630,N_15292,N_15327);
or U15631 (N_15631,N_15417,N_15363);
xor U15632 (N_15632,N_15367,N_15463);
xnor U15633 (N_15633,N_15335,N_15438);
nand U15634 (N_15634,N_15296,N_15389);
or U15635 (N_15635,N_15419,N_15494);
nand U15636 (N_15636,N_15279,N_15465);
nor U15637 (N_15637,N_15464,N_15431);
nor U15638 (N_15638,N_15358,N_15270);
nor U15639 (N_15639,N_15437,N_15332);
and U15640 (N_15640,N_15423,N_15365);
and U15641 (N_15641,N_15285,N_15390);
nand U15642 (N_15642,N_15282,N_15447);
or U15643 (N_15643,N_15261,N_15272);
nor U15644 (N_15644,N_15332,N_15382);
nor U15645 (N_15645,N_15444,N_15347);
nor U15646 (N_15646,N_15323,N_15469);
nor U15647 (N_15647,N_15462,N_15454);
nand U15648 (N_15648,N_15294,N_15338);
or U15649 (N_15649,N_15389,N_15476);
nand U15650 (N_15650,N_15374,N_15333);
xor U15651 (N_15651,N_15300,N_15334);
xor U15652 (N_15652,N_15496,N_15381);
or U15653 (N_15653,N_15370,N_15309);
xor U15654 (N_15654,N_15384,N_15350);
nand U15655 (N_15655,N_15413,N_15447);
nand U15656 (N_15656,N_15317,N_15395);
or U15657 (N_15657,N_15490,N_15291);
nor U15658 (N_15658,N_15284,N_15312);
xor U15659 (N_15659,N_15448,N_15368);
xnor U15660 (N_15660,N_15404,N_15440);
and U15661 (N_15661,N_15470,N_15491);
nand U15662 (N_15662,N_15449,N_15308);
nand U15663 (N_15663,N_15428,N_15260);
and U15664 (N_15664,N_15471,N_15308);
nor U15665 (N_15665,N_15300,N_15304);
or U15666 (N_15666,N_15480,N_15466);
nor U15667 (N_15667,N_15311,N_15473);
or U15668 (N_15668,N_15263,N_15305);
xnor U15669 (N_15669,N_15256,N_15353);
or U15670 (N_15670,N_15319,N_15285);
xor U15671 (N_15671,N_15355,N_15381);
or U15672 (N_15672,N_15376,N_15440);
nor U15673 (N_15673,N_15426,N_15262);
xnor U15674 (N_15674,N_15328,N_15393);
and U15675 (N_15675,N_15329,N_15379);
nor U15676 (N_15676,N_15489,N_15459);
or U15677 (N_15677,N_15470,N_15287);
nor U15678 (N_15678,N_15498,N_15449);
nand U15679 (N_15679,N_15398,N_15265);
and U15680 (N_15680,N_15432,N_15277);
xor U15681 (N_15681,N_15497,N_15358);
nand U15682 (N_15682,N_15254,N_15258);
nor U15683 (N_15683,N_15413,N_15451);
nor U15684 (N_15684,N_15313,N_15355);
or U15685 (N_15685,N_15456,N_15264);
or U15686 (N_15686,N_15365,N_15390);
nand U15687 (N_15687,N_15296,N_15266);
nand U15688 (N_15688,N_15458,N_15445);
xor U15689 (N_15689,N_15273,N_15302);
xor U15690 (N_15690,N_15474,N_15440);
and U15691 (N_15691,N_15270,N_15350);
or U15692 (N_15692,N_15361,N_15401);
nand U15693 (N_15693,N_15480,N_15373);
or U15694 (N_15694,N_15458,N_15276);
xor U15695 (N_15695,N_15452,N_15453);
and U15696 (N_15696,N_15456,N_15436);
or U15697 (N_15697,N_15455,N_15486);
nor U15698 (N_15698,N_15487,N_15422);
xnor U15699 (N_15699,N_15343,N_15491);
nand U15700 (N_15700,N_15354,N_15335);
and U15701 (N_15701,N_15423,N_15401);
xnor U15702 (N_15702,N_15413,N_15433);
nor U15703 (N_15703,N_15475,N_15415);
xnor U15704 (N_15704,N_15355,N_15416);
xor U15705 (N_15705,N_15387,N_15326);
or U15706 (N_15706,N_15456,N_15434);
or U15707 (N_15707,N_15304,N_15329);
or U15708 (N_15708,N_15464,N_15256);
or U15709 (N_15709,N_15491,N_15308);
or U15710 (N_15710,N_15498,N_15262);
and U15711 (N_15711,N_15476,N_15385);
and U15712 (N_15712,N_15384,N_15431);
xnor U15713 (N_15713,N_15308,N_15349);
nor U15714 (N_15714,N_15472,N_15447);
nand U15715 (N_15715,N_15273,N_15297);
and U15716 (N_15716,N_15408,N_15450);
nor U15717 (N_15717,N_15352,N_15446);
nor U15718 (N_15718,N_15388,N_15491);
xor U15719 (N_15719,N_15287,N_15415);
or U15720 (N_15720,N_15339,N_15314);
or U15721 (N_15721,N_15484,N_15301);
and U15722 (N_15722,N_15349,N_15317);
nor U15723 (N_15723,N_15392,N_15463);
or U15724 (N_15724,N_15364,N_15301);
and U15725 (N_15725,N_15289,N_15253);
nand U15726 (N_15726,N_15436,N_15444);
nor U15727 (N_15727,N_15336,N_15252);
nor U15728 (N_15728,N_15397,N_15493);
or U15729 (N_15729,N_15252,N_15453);
xnor U15730 (N_15730,N_15340,N_15309);
nand U15731 (N_15731,N_15262,N_15278);
xor U15732 (N_15732,N_15331,N_15288);
or U15733 (N_15733,N_15307,N_15455);
nand U15734 (N_15734,N_15280,N_15396);
or U15735 (N_15735,N_15325,N_15250);
xnor U15736 (N_15736,N_15334,N_15288);
nor U15737 (N_15737,N_15292,N_15452);
nor U15738 (N_15738,N_15430,N_15489);
and U15739 (N_15739,N_15400,N_15281);
and U15740 (N_15740,N_15341,N_15376);
xor U15741 (N_15741,N_15402,N_15333);
and U15742 (N_15742,N_15413,N_15485);
nand U15743 (N_15743,N_15335,N_15386);
xnor U15744 (N_15744,N_15449,N_15440);
and U15745 (N_15745,N_15287,N_15276);
and U15746 (N_15746,N_15327,N_15294);
xor U15747 (N_15747,N_15312,N_15466);
nor U15748 (N_15748,N_15462,N_15379);
xor U15749 (N_15749,N_15398,N_15491);
nor U15750 (N_15750,N_15642,N_15617);
and U15751 (N_15751,N_15718,N_15512);
nor U15752 (N_15752,N_15604,N_15634);
xor U15753 (N_15753,N_15656,N_15662);
or U15754 (N_15754,N_15686,N_15585);
xnor U15755 (N_15755,N_15500,N_15707);
xnor U15756 (N_15756,N_15513,N_15599);
nor U15757 (N_15757,N_15511,N_15545);
nor U15758 (N_15758,N_15678,N_15597);
xnor U15759 (N_15759,N_15529,N_15616);
xor U15760 (N_15760,N_15677,N_15539);
or U15761 (N_15761,N_15552,N_15659);
nand U15762 (N_15762,N_15622,N_15679);
nor U15763 (N_15763,N_15544,N_15701);
nor U15764 (N_15764,N_15525,N_15609);
nor U15765 (N_15765,N_15613,N_15533);
nor U15766 (N_15766,N_15692,N_15726);
nor U15767 (N_15767,N_15700,N_15565);
and U15768 (N_15768,N_15652,N_15605);
nand U15769 (N_15769,N_15637,N_15504);
nor U15770 (N_15770,N_15651,N_15671);
xor U15771 (N_15771,N_15577,N_15509);
nor U15772 (N_15772,N_15543,N_15653);
xor U15773 (N_15773,N_15703,N_15748);
and U15774 (N_15774,N_15550,N_15635);
and U15775 (N_15775,N_15666,N_15714);
or U15776 (N_15776,N_15591,N_15719);
nand U15777 (N_15777,N_15636,N_15625);
and U15778 (N_15778,N_15689,N_15628);
or U15779 (N_15779,N_15670,N_15621);
or U15780 (N_15780,N_15615,N_15515);
nor U15781 (N_15781,N_15696,N_15502);
nand U15782 (N_15782,N_15590,N_15744);
and U15783 (N_15783,N_15594,N_15580);
xor U15784 (N_15784,N_15734,N_15669);
and U15785 (N_15785,N_15732,N_15655);
nor U15786 (N_15786,N_15535,N_15595);
and U15787 (N_15787,N_15610,N_15606);
and U15788 (N_15788,N_15747,N_15521);
xnor U15789 (N_15789,N_15690,N_15680);
nand U15790 (N_15790,N_15537,N_15534);
nor U15791 (N_15791,N_15568,N_15508);
nand U15792 (N_15792,N_15742,N_15694);
xnor U15793 (N_15793,N_15522,N_15728);
xor U15794 (N_15794,N_15560,N_15675);
xnor U15795 (N_15795,N_15695,N_15576);
xnor U15796 (N_15796,N_15586,N_15654);
or U15797 (N_15797,N_15598,N_15731);
nand U15798 (N_15798,N_15602,N_15710);
nand U15799 (N_15799,N_15561,N_15667);
xnor U15800 (N_15800,N_15526,N_15640);
xnor U15801 (N_15801,N_15608,N_15517);
xnor U15802 (N_15802,N_15743,N_15601);
nor U15803 (N_15803,N_15519,N_15660);
and U15804 (N_15804,N_15623,N_15709);
nor U15805 (N_15805,N_15717,N_15574);
and U15806 (N_15806,N_15548,N_15518);
xnor U15807 (N_15807,N_15739,N_15647);
or U15808 (N_15808,N_15596,N_15632);
nor U15809 (N_15809,N_15600,N_15638);
or U15810 (N_15810,N_15672,N_15564);
and U15811 (N_15811,N_15722,N_15566);
nor U15812 (N_15812,N_15614,N_15557);
xor U15813 (N_15813,N_15639,N_15658);
nor U15814 (N_15814,N_15661,N_15501);
or U15815 (N_15815,N_15746,N_15620);
nand U15816 (N_15816,N_15546,N_15573);
nand U15817 (N_15817,N_15749,N_15611);
or U15818 (N_15818,N_15674,N_15527);
nand U15819 (N_15819,N_15542,N_15551);
or U15820 (N_15820,N_15730,N_15740);
or U15821 (N_15821,N_15698,N_15607);
and U15822 (N_15822,N_15741,N_15558);
nand U15823 (N_15823,N_15587,N_15688);
nor U15824 (N_15824,N_15725,N_15673);
nor U15825 (N_15825,N_15584,N_15592);
or U15826 (N_15826,N_15650,N_15531);
and U15827 (N_15827,N_15721,N_15588);
or U15828 (N_15828,N_15704,N_15645);
nand U15829 (N_15829,N_15676,N_15745);
nand U15830 (N_15830,N_15699,N_15593);
or U15831 (N_15831,N_15540,N_15603);
nor U15832 (N_15832,N_15729,N_15559);
nor U15833 (N_15833,N_15624,N_15716);
or U15834 (N_15834,N_15668,N_15570);
nand U15835 (N_15835,N_15554,N_15644);
and U15836 (N_15836,N_15618,N_15530);
and U15837 (N_15837,N_15643,N_15578);
xor U15838 (N_15838,N_15646,N_15631);
nor U15839 (N_15839,N_15708,N_15663);
nand U15840 (N_15840,N_15702,N_15626);
or U15841 (N_15841,N_15507,N_15735);
nand U15842 (N_15842,N_15664,N_15524);
xor U15843 (N_15843,N_15629,N_15555);
and U15844 (N_15844,N_15736,N_15583);
nor U15845 (N_15845,N_15589,N_15723);
xor U15846 (N_15846,N_15681,N_15612);
nor U15847 (N_15847,N_15541,N_15506);
or U15848 (N_15848,N_15579,N_15581);
nor U15849 (N_15849,N_15549,N_15569);
xor U15850 (N_15850,N_15505,N_15737);
nand U15851 (N_15851,N_15538,N_15532);
or U15852 (N_15852,N_15682,N_15503);
xor U15853 (N_15853,N_15619,N_15571);
or U15854 (N_15854,N_15691,N_15516);
nor U15855 (N_15855,N_15724,N_15657);
nand U15856 (N_15856,N_15633,N_15711);
and U15857 (N_15857,N_15713,N_15697);
or U15858 (N_15858,N_15572,N_15553);
nor U15859 (N_15859,N_15720,N_15738);
nor U15860 (N_15860,N_15733,N_15665);
or U15861 (N_15861,N_15582,N_15684);
xor U15862 (N_15862,N_15693,N_15514);
or U15863 (N_15863,N_15712,N_15706);
nand U15864 (N_15864,N_15649,N_15510);
nand U15865 (N_15865,N_15648,N_15547);
and U15866 (N_15866,N_15520,N_15641);
nor U15867 (N_15867,N_15536,N_15528);
nand U15868 (N_15868,N_15727,N_15563);
xor U15869 (N_15869,N_15575,N_15523);
and U15870 (N_15870,N_15685,N_15567);
or U15871 (N_15871,N_15627,N_15683);
nor U15872 (N_15872,N_15630,N_15687);
nor U15873 (N_15873,N_15705,N_15556);
and U15874 (N_15874,N_15562,N_15715);
nand U15875 (N_15875,N_15637,N_15663);
or U15876 (N_15876,N_15634,N_15513);
xnor U15877 (N_15877,N_15584,N_15513);
xnor U15878 (N_15878,N_15660,N_15525);
and U15879 (N_15879,N_15542,N_15662);
xor U15880 (N_15880,N_15749,N_15654);
nor U15881 (N_15881,N_15512,N_15749);
and U15882 (N_15882,N_15703,N_15530);
xnor U15883 (N_15883,N_15720,N_15500);
or U15884 (N_15884,N_15583,N_15734);
nor U15885 (N_15885,N_15668,N_15545);
or U15886 (N_15886,N_15740,N_15643);
nand U15887 (N_15887,N_15561,N_15542);
or U15888 (N_15888,N_15532,N_15635);
or U15889 (N_15889,N_15731,N_15721);
xor U15890 (N_15890,N_15695,N_15580);
or U15891 (N_15891,N_15731,N_15689);
and U15892 (N_15892,N_15552,N_15551);
nor U15893 (N_15893,N_15676,N_15585);
or U15894 (N_15894,N_15594,N_15717);
or U15895 (N_15895,N_15695,N_15503);
nor U15896 (N_15896,N_15722,N_15657);
or U15897 (N_15897,N_15578,N_15695);
or U15898 (N_15898,N_15729,N_15722);
xor U15899 (N_15899,N_15722,N_15737);
nand U15900 (N_15900,N_15676,N_15552);
xnor U15901 (N_15901,N_15663,N_15737);
xor U15902 (N_15902,N_15593,N_15601);
or U15903 (N_15903,N_15718,N_15504);
xor U15904 (N_15904,N_15608,N_15658);
nor U15905 (N_15905,N_15568,N_15546);
and U15906 (N_15906,N_15599,N_15580);
nor U15907 (N_15907,N_15588,N_15524);
and U15908 (N_15908,N_15526,N_15653);
nor U15909 (N_15909,N_15564,N_15634);
xor U15910 (N_15910,N_15514,N_15546);
or U15911 (N_15911,N_15617,N_15574);
xnor U15912 (N_15912,N_15594,N_15518);
nand U15913 (N_15913,N_15561,N_15610);
xnor U15914 (N_15914,N_15748,N_15694);
or U15915 (N_15915,N_15713,N_15709);
xor U15916 (N_15916,N_15516,N_15613);
xnor U15917 (N_15917,N_15548,N_15618);
and U15918 (N_15918,N_15617,N_15544);
and U15919 (N_15919,N_15556,N_15719);
nor U15920 (N_15920,N_15638,N_15636);
and U15921 (N_15921,N_15537,N_15691);
and U15922 (N_15922,N_15525,N_15529);
or U15923 (N_15923,N_15698,N_15510);
nor U15924 (N_15924,N_15604,N_15534);
xor U15925 (N_15925,N_15525,N_15734);
nor U15926 (N_15926,N_15631,N_15679);
and U15927 (N_15927,N_15669,N_15587);
and U15928 (N_15928,N_15611,N_15710);
or U15929 (N_15929,N_15617,N_15523);
nand U15930 (N_15930,N_15519,N_15529);
and U15931 (N_15931,N_15739,N_15511);
nand U15932 (N_15932,N_15607,N_15516);
or U15933 (N_15933,N_15600,N_15598);
and U15934 (N_15934,N_15642,N_15733);
and U15935 (N_15935,N_15741,N_15586);
or U15936 (N_15936,N_15546,N_15702);
and U15937 (N_15937,N_15729,N_15726);
or U15938 (N_15938,N_15669,N_15511);
nor U15939 (N_15939,N_15723,N_15695);
nor U15940 (N_15940,N_15702,N_15743);
nor U15941 (N_15941,N_15622,N_15705);
and U15942 (N_15942,N_15685,N_15699);
xor U15943 (N_15943,N_15657,N_15645);
xor U15944 (N_15944,N_15529,N_15524);
nor U15945 (N_15945,N_15690,N_15577);
xnor U15946 (N_15946,N_15634,N_15557);
xnor U15947 (N_15947,N_15626,N_15659);
and U15948 (N_15948,N_15548,N_15601);
nor U15949 (N_15949,N_15661,N_15705);
and U15950 (N_15950,N_15641,N_15708);
nand U15951 (N_15951,N_15739,N_15665);
xor U15952 (N_15952,N_15639,N_15529);
and U15953 (N_15953,N_15508,N_15577);
or U15954 (N_15954,N_15603,N_15579);
nor U15955 (N_15955,N_15621,N_15529);
xor U15956 (N_15956,N_15623,N_15705);
nand U15957 (N_15957,N_15512,N_15568);
xor U15958 (N_15958,N_15660,N_15688);
nand U15959 (N_15959,N_15559,N_15635);
or U15960 (N_15960,N_15534,N_15601);
or U15961 (N_15961,N_15713,N_15729);
nor U15962 (N_15962,N_15518,N_15666);
nor U15963 (N_15963,N_15682,N_15603);
xnor U15964 (N_15964,N_15582,N_15514);
nand U15965 (N_15965,N_15620,N_15735);
nand U15966 (N_15966,N_15698,N_15628);
xnor U15967 (N_15967,N_15561,N_15694);
xnor U15968 (N_15968,N_15658,N_15726);
nor U15969 (N_15969,N_15720,N_15529);
nand U15970 (N_15970,N_15623,N_15602);
xor U15971 (N_15971,N_15521,N_15729);
nor U15972 (N_15972,N_15678,N_15649);
and U15973 (N_15973,N_15724,N_15531);
nor U15974 (N_15974,N_15594,N_15621);
nand U15975 (N_15975,N_15632,N_15541);
nor U15976 (N_15976,N_15511,N_15662);
or U15977 (N_15977,N_15736,N_15509);
nor U15978 (N_15978,N_15716,N_15634);
and U15979 (N_15979,N_15714,N_15665);
and U15980 (N_15980,N_15744,N_15617);
nor U15981 (N_15981,N_15691,N_15625);
xor U15982 (N_15982,N_15667,N_15746);
or U15983 (N_15983,N_15557,N_15519);
xor U15984 (N_15984,N_15523,N_15737);
nand U15985 (N_15985,N_15519,N_15601);
xor U15986 (N_15986,N_15553,N_15660);
and U15987 (N_15987,N_15553,N_15516);
nor U15988 (N_15988,N_15690,N_15692);
and U15989 (N_15989,N_15659,N_15593);
and U15990 (N_15990,N_15702,N_15733);
and U15991 (N_15991,N_15590,N_15670);
nor U15992 (N_15992,N_15526,N_15572);
nand U15993 (N_15993,N_15662,N_15592);
xor U15994 (N_15994,N_15721,N_15655);
xor U15995 (N_15995,N_15739,N_15689);
xnor U15996 (N_15996,N_15724,N_15551);
xnor U15997 (N_15997,N_15698,N_15648);
or U15998 (N_15998,N_15513,N_15525);
nor U15999 (N_15999,N_15637,N_15626);
nand U16000 (N_16000,N_15827,N_15829);
nand U16001 (N_16001,N_15835,N_15886);
and U16002 (N_16002,N_15962,N_15864);
nand U16003 (N_16003,N_15927,N_15969);
xor U16004 (N_16004,N_15921,N_15970);
and U16005 (N_16005,N_15910,N_15803);
nor U16006 (N_16006,N_15841,N_15865);
and U16007 (N_16007,N_15906,N_15791);
nor U16008 (N_16008,N_15901,N_15909);
and U16009 (N_16009,N_15982,N_15957);
xnor U16010 (N_16010,N_15917,N_15805);
or U16011 (N_16011,N_15937,N_15920);
xor U16012 (N_16012,N_15875,N_15898);
xor U16013 (N_16013,N_15944,N_15911);
nor U16014 (N_16014,N_15833,N_15936);
nand U16015 (N_16015,N_15961,N_15767);
or U16016 (N_16016,N_15928,N_15776);
nor U16017 (N_16017,N_15879,N_15996);
nand U16018 (N_16018,N_15950,N_15770);
or U16019 (N_16019,N_15856,N_15849);
or U16020 (N_16020,N_15801,N_15787);
nor U16021 (N_16021,N_15765,N_15907);
nand U16022 (N_16022,N_15860,N_15857);
nand U16023 (N_16023,N_15812,N_15868);
and U16024 (N_16024,N_15793,N_15929);
xnor U16025 (N_16025,N_15878,N_15756);
xnor U16026 (N_16026,N_15940,N_15795);
nor U16027 (N_16027,N_15843,N_15932);
nor U16028 (N_16028,N_15968,N_15834);
nand U16029 (N_16029,N_15766,N_15863);
or U16030 (N_16030,N_15895,N_15983);
or U16031 (N_16031,N_15882,N_15903);
nor U16032 (N_16032,N_15930,N_15771);
nand U16033 (N_16033,N_15897,N_15811);
and U16034 (N_16034,N_15781,N_15995);
nor U16035 (N_16035,N_15991,N_15981);
xor U16036 (N_16036,N_15872,N_15783);
and U16037 (N_16037,N_15926,N_15855);
nor U16038 (N_16038,N_15816,N_15777);
nand U16039 (N_16039,N_15925,N_15974);
nand U16040 (N_16040,N_15847,N_15821);
xnor U16041 (N_16041,N_15956,N_15946);
nor U16042 (N_16042,N_15867,N_15818);
xor U16043 (N_16043,N_15858,N_15804);
nor U16044 (N_16044,N_15922,N_15892);
or U16045 (N_16045,N_15785,N_15820);
and U16046 (N_16046,N_15825,N_15914);
nand U16047 (N_16047,N_15992,N_15784);
or U16048 (N_16048,N_15758,N_15837);
or U16049 (N_16049,N_15966,N_15848);
xor U16050 (N_16050,N_15989,N_15819);
or U16051 (N_16051,N_15838,N_15964);
xor U16052 (N_16052,N_15953,N_15931);
xnor U16053 (N_16053,N_15845,N_15952);
nand U16054 (N_16054,N_15870,N_15902);
nand U16055 (N_16055,N_15792,N_15822);
nand U16056 (N_16056,N_15800,N_15891);
nor U16057 (N_16057,N_15852,N_15808);
or U16058 (N_16058,N_15880,N_15762);
xor U16059 (N_16059,N_15994,N_15814);
xor U16060 (N_16060,N_15876,N_15883);
and U16061 (N_16061,N_15862,N_15918);
xnor U16062 (N_16062,N_15809,N_15951);
or U16063 (N_16063,N_15881,N_15761);
xor U16064 (N_16064,N_15802,N_15960);
or U16065 (N_16065,N_15993,N_15851);
or U16066 (N_16066,N_15861,N_15884);
and U16067 (N_16067,N_15775,N_15810);
or U16068 (N_16068,N_15839,N_15939);
or U16069 (N_16069,N_15885,N_15840);
and U16070 (N_16070,N_15997,N_15943);
nor U16071 (N_16071,N_15975,N_15831);
xor U16072 (N_16072,N_15899,N_15817);
nand U16073 (N_16073,N_15807,N_15972);
xnor U16074 (N_16074,N_15958,N_15913);
xor U16075 (N_16075,N_15873,N_15798);
or U16076 (N_16076,N_15824,N_15912);
nand U16077 (N_16077,N_15977,N_15947);
and U16078 (N_16078,N_15985,N_15769);
or U16079 (N_16079,N_15751,N_15768);
and U16080 (N_16080,N_15967,N_15763);
nor U16081 (N_16081,N_15905,N_15774);
xnor U16082 (N_16082,N_15780,N_15850);
or U16083 (N_16083,N_15945,N_15755);
nor U16084 (N_16084,N_15908,N_15904);
and U16085 (N_16085,N_15887,N_15806);
nor U16086 (N_16086,N_15978,N_15934);
nor U16087 (N_16087,N_15797,N_15773);
xor U16088 (N_16088,N_15836,N_15789);
nand U16089 (N_16089,N_15890,N_15955);
or U16090 (N_16090,N_15853,N_15764);
and U16091 (N_16091,N_15894,N_15832);
xnor U16092 (N_16092,N_15933,N_15772);
and U16093 (N_16093,N_15971,N_15782);
and U16094 (N_16094,N_15778,N_15854);
nand U16095 (N_16095,N_15828,N_15842);
nand U16096 (N_16096,N_15916,N_15889);
and U16097 (N_16097,N_15924,N_15794);
nor U16098 (N_16098,N_15893,N_15900);
or U16099 (N_16099,N_15796,N_15757);
nor U16100 (N_16100,N_15986,N_15874);
and U16101 (N_16101,N_15759,N_15919);
and U16102 (N_16102,N_15813,N_15990);
nor U16103 (N_16103,N_15790,N_15941);
or U16104 (N_16104,N_15753,N_15999);
xor U16105 (N_16105,N_15976,N_15866);
or U16106 (N_16106,N_15954,N_15844);
and U16107 (N_16107,N_15869,N_15760);
and U16108 (N_16108,N_15799,N_15750);
nand U16109 (N_16109,N_15754,N_15923);
nand U16110 (N_16110,N_15959,N_15938);
nor U16111 (N_16111,N_15871,N_15752);
nor U16112 (N_16112,N_15987,N_15942);
nor U16113 (N_16113,N_15973,N_15965);
xor U16114 (N_16114,N_15979,N_15815);
and U16115 (N_16115,N_15963,N_15859);
xnor U16116 (N_16116,N_15915,N_15896);
nor U16117 (N_16117,N_15846,N_15786);
xnor U16118 (N_16118,N_15823,N_15830);
and U16119 (N_16119,N_15826,N_15980);
nand U16120 (N_16120,N_15988,N_15877);
xnor U16121 (N_16121,N_15984,N_15949);
or U16122 (N_16122,N_15948,N_15998);
nand U16123 (N_16123,N_15779,N_15935);
nor U16124 (N_16124,N_15888,N_15788);
nand U16125 (N_16125,N_15939,N_15962);
or U16126 (N_16126,N_15820,N_15755);
or U16127 (N_16127,N_15977,N_15796);
xnor U16128 (N_16128,N_15881,N_15982);
nor U16129 (N_16129,N_15989,N_15866);
and U16130 (N_16130,N_15863,N_15964);
and U16131 (N_16131,N_15848,N_15916);
or U16132 (N_16132,N_15912,N_15983);
nor U16133 (N_16133,N_15761,N_15864);
and U16134 (N_16134,N_15819,N_15795);
nand U16135 (N_16135,N_15930,N_15974);
and U16136 (N_16136,N_15806,N_15873);
xnor U16137 (N_16137,N_15998,N_15867);
nor U16138 (N_16138,N_15871,N_15844);
nand U16139 (N_16139,N_15978,N_15896);
and U16140 (N_16140,N_15918,N_15994);
xor U16141 (N_16141,N_15979,N_15985);
xnor U16142 (N_16142,N_15797,N_15770);
nor U16143 (N_16143,N_15916,N_15951);
nor U16144 (N_16144,N_15851,N_15939);
xnor U16145 (N_16145,N_15881,N_15827);
or U16146 (N_16146,N_15962,N_15930);
nor U16147 (N_16147,N_15784,N_15756);
nand U16148 (N_16148,N_15945,N_15814);
or U16149 (N_16149,N_15989,N_15887);
xnor U16150 (N_16150,N_15958,N_15767);
nor U16151 (N_16151,N_15810,N_15786);
nor U16152 (N_16152,N_15777,N_15795);
and U16153 (N_16153,N_15971,N_15915);
nor U16154 (N_16154,N_15807,N_15948);
and U16155 (N_16155,N_15761,N_15974);
or U16156 (N_16156,N_15770,N_15957);
or U16157 (N_16157,N_15752,N_15800);
nand U16158 (N_16158,N_15955,N_15760);
nand U16159 (N_16159,N_15893,N_15834);
or U16160 (N_16160,N_15866,N_15823);
or U16161 (N_16161,N_15791,N_15892);
nand U16162 (N_16162,N_15837,N_15914);
or U16163 (N_16163,N_15819,N_15912);
nand U16164 (N_16164,N_15920,N_15767);
xnor U16165 (N_16165,N_15820,N_15985);
xnor U16166 (N_16166,N_15977,N_15958);
xnor U16167 (N_16167,N_15764,N_15750);
nand U16168 (N_16168,N_15769,N_15795);
nand U16169 (N_16169,N_15871,N_15904);
nand U16170 (N_16170,N_15767,N_15823);
and U16171 (N_16171,N_15943,N_15813);
nand U16172 (N_16172,N_15901,N_15950);
xnor U16173 (N_16173,N_15941,N_15944);
nor U16174 (N_16174,N_15993,N_15862);
and U16175 (N_16175,N_15902,N_15777);
xnor U16176 (N_16176,N_15962,N_15915);
nand U16177 (N_16177,N_15928,N_15851);
or U16178 (N_16178,N_15819,N_15997);
nor U16179 (N_16179,N_15980,N_15804);
xor U16180 (N_16180,N_15909,N_15898);
xnor U16181 (N_16181,N_15802,N_15957);
nor U16182 (N_16182,N_15784,N_15866);
xnor U16183 (N_16183,N_15877,N_15861);
and U16184 (N_16184,N_15896,N_15878);
nand U16185 (N_16185,N_15784,N_15975);
xor U16186 (N_16186,N_15866,N_15916);
xnor U16187 (N_16187,N_15996,N_15931);
nor U16188 (N_16188,N_15847,N_15825);
nand U16189 (N_16189,N_15996,N_15962);
nand U16190 (N_16190,N_15835,N_15933);
or U16191 (N_16191,N_15762,N_15794);
or U16192 (N_16192,N_15913,N_15865);
nand U16193 (N_16193,N_15810,N_15849);
and U16194 (N_16194,N_15754,N_15851);
nor U16195 (N_16195,N_15972,N_15844);
nor U16196 (N_16196,N_15968,N_15814);
nor U16197 (N_16197,N_15904,N_15812);
nor U16198 (N_16198,N_15867,N_15797);
xnor U16199 (N_16199,N_15916,N_15752);
nand U16200 (N_16200,N_15796,N_15798);
nand U16201 (N_16201,N_15760,N_15766);
and U16202 (N_16202,N_15988,N_15751);
xor U16203 (N_16203,N_15854,N_15979);
nor U16204 (N_16204,N_15761,N_15779);
or U16205 (N_16205,N_15788,N_15785);
or U16206 (N_16206,N_15841,N_15973);
nor U16207 (N_16207,N_15826,N_15943);
nor U16208 (N_16208,N_15886,N_15752);
nand U16209 (N_16209,N_15801,N_15860);
and U16210 (N_16210,N_15881,N_15889);
and U16211 (N_16211,N_15889,N_15861);
xor U16212 (N_16212,N_15893,N_15866);
nand U16213 (N_16213,N_15793,N_15774);
or U16214 (N_16214,N_15763,N_15975);
or U16215 (N_16215,N_15973,N_15826);
or U16216 (N_16216,N_15836,N_15839);
nor U16217 (N_16217,N_15852,N_15903);
nor U16218 (N_16218,N_15902,N_15834);
nand U16219 (N_16219,N_15846,N_15764);
and U16220 (N_16220,N_15918,N_15783);
xnor U16221 (N_16221,N_15805,N_15862);
nand U16222 (N_16222,N_15787,N_15906);
and U16223 (N_16223,N_15943,N_15791);
and U16224 (N_16224,N_15829,N_15905);
nor U16225 (N_16225,N_15974,N_15794);
nor U16226 (N_16226,N_15879,N_15800);
and U16227 (N_16227,N_15845,N_15765);
nor U16228 (N_16228,N_15899,N_15862);
or U16229 (N_16229,N_15763,N_15930);
nor U16230 (N_16230,N_15978,N_15988);
and U16231 (N_16231,N_15757,N_15999);
nand U16232 (N_16232,N_15848,N_15758);
nor U16233 (N_16233,N_15813,N_15867);
and U16234 (N_16234,N_15953,N_15867);
xor U16235 (N_16235,N_15791,N_15921);
and U16236 (N_16236,N_15895,N_15955);
nand U16237 (N_16237,N_15852,N_15995);
xnor U16238 (N_16238,N_15830,N_15884);
xnor U16239 (N_16239,N_15952,N_15770);
or U16240 (N_16240,N_15786,N_15949);
or U16241 (N_16241,N_15754,N_15868);
or U16242 (N_16242,N_15784,N_15765);
nand U16243 (N_16243,N_15847,N_15998);
nor U16244 (N_16244,N_15971,N_15881);
or U16245 (N_16245,N_15817,N_15861);
nand U16246 (N_16246,N_15874,N_15898);
nand U16247 (N_16247,N_15976,N_15906);
nand U16248 (N_16248,N_15808,N_15976);
xor U16249 (N_16249,N_15894,N_15826);
and U16250 (N_16250,N_16131,N_16206);
nor U16251 (N_16251,N_16134,N_16077);
nor U16252 (N_16252,N_16031,N_16071);
nand U16253 (N_16253,N_16147,N_16098);
nand U16254 (N_16254,N_16014,N_16075);
nand U16255 (N_16255,N_16101,N_16142);
and U16256 (N_16256,N_16180,N_16029);
xnor U16257 (N_16257,N_16128,N_16230);
nand U16258 (N_16258,N_16070,N_16048);
nor U16259 (N_16259,N_16249,N_16172);
or U16260 (N_16260,N_16239,N_16084);
nor U16261 (N_16261,N_16212,N_16137);
nor U16262 (N_16262,N_16190,N_16138);
or U16263 (N_16263,N_16245,N_16205);
nand U16264 (N_16264,N_16114,N_16069);
nand U16265 (N_16265,N_16129,N_16220);
or U16266 (N_16266,N_16167,N_16100);
and U16267 (N_16267,N_16174,N_16045);
nand U16268 (N_16268,N_16079,N_16231);
nor U16269 (N_16269,N_16235,N_16015);
or U16270 (N_16270,N_16112,N_16052);
xor U16271 (N_16271,N_16103,N_16182);
xor U16272 (N_16272,N_16140,N_16021);
xnor U16273 (N_16273,N_16153,N_16189);
xnor U16274 (N_16274,N_16003,N_16081);
nor U16275 (N_16275,N_16166,N_16169);
nor U16276 (N_16276,N_16120,N_16043);
and U16277 (N_16277,N_16159,N_16096);
xnor U16278 (N_16278,N_16049,N_16030);
nand U16279 (N_16279,N_16177,N_16121);
or U16280 (N_16280,N_16032,N_16025);
nor U16281 (N_16281,N_16179,N_16068);
or U16282 (N_16282,N_16173,N_16204);
xor U16283 (N_16283,N_16028,N_16006);
xor U16284 (N_16284,N_16203,N_16136);
and U16285 (N_16285,N_16132,N_16171);
nand U16286 (N_16286,N_16082,N_16165);
and U16287 (N_16287,N_16067,N_16026);
nor U16288 (N_16288,N_16144,N_16020);
xnor U16289 (N_16289,N_16073,N_16095);
nand U16290 (N_16290,N_16023,N_16091);
nand U16291 (N_16291,N_16184,N_16200);
nor U16292 (N_16292,N_16024,N_16139);
nand U16293 (N_16293,N_16018,N_16149);
xnor U16294 (N_16294,N_16234,N_16115);
or U16295 (N_16295,N_16001,N_16141);
nor U16296 (N_16296,N_16150,N_16085);
and U16297 (N_16297,N_16053,N_16090);
nand U16298 (N_16298,N_16010,N_16219);
and U16299 (N_16299,N_16016,N_16221);
or U16300 (N_16300,N_16197,N_16229);
xor U16301 (N_16301,N_16034,N_16154);
xnor U16302 (N_16302,N_16074,N_16248);
xor U16303 (N_16303,N_16185,N_16145);
xor U16304 (N_16304,N_16099,N_16004);
xor U16305 (N_16305,N_16218,N_16041);
or U16306 (N_16306,N_16046,N_16164);
nor U16307 (N_16307,N_16093,N_16056);
xnor U16308 (N_16308,N_16163,N_16040);
nor U16309 (N_16309,N_16247,N_16201);
nand U16310 (N_16310,N_16155,N_16186);
and U16311 (N_16311,N_16094,N_16176);
xnor U16312 (N_16312,N_16215,N_16236);
nand U16313 (N_16313,N_16119,N_16035);
and U16314 (N_16314,N_16047,N_16207);
or U16315 (N_16315,N_16042,N_16113);
or U16316 (N_16316,N_16143,N_16228);
nor U16317 (N_16317,N_16156,N_16037);
or U16318 (N_16318,N_16017,N_16187);
nor U16319 (N_16319,N_16102,N_16213);
nand U16320 (N_16320,N_16214,N_16122);
nand U16321 (N_16321,N_16243,N_16022);
nand U16322 (N_16322,N_16244,N_16192);
nand U16323 (N_16323,N_16124,N_16088);
nor U16324 (N_16324,N_16011,N_16060);
and U16325 (N_16325,N_16237,N_16111);
or U16326 (N_16326,N_16216,N_16118);
nor U16327 (N_16327,N_16133,N_16196);
nand U16328 (N_16328,N_16036,N_16123);
or U16329 (N_16329,N_16202,N_16027);
nor U16330 (N_16330,N_16193,N_16058);
nor U16331 (N_16331,N_16066,N_16242);
xor U16332 (N_16332,N_16227,N_16086);
or U16333 (N_16333,N_16157,N_16199);
and U16334 (N_16334,N_16125,N_16054);
nand U16335 (N_16335,N_16208,N_16151);
and U16336 (N_16336,N_16033,N_16050);
or U16337 (N_16337,N_16222,N_16183);
nor U16338 (N_16338,N_16059,N_16209);
or U16339 (N_16339,N_16065,N_16051);
and U16340 (N_16340,N_16224,N_16062);
and U16341 (N_16341,N_16000,N_16195);
xnor U16342 (N_16342,N_16170,N_16063);
nor U16343 (N_16343,N_16083,N_16191);
nand U16344 (N_16344,N_16104,N_16080);
nand U16345 (N_16345,N_16148,N_16109);
nand U16346 (N_16346,N_16130,N_16097);
nor U16347 (N_16347,N_16108,N_16013);
xnor U16348 (N_16348,N_16117,N_16226);
or U16349 (N_16349,N_16188,N_16044);
nand U16350 (N_16350,N_16232,N_16039);
or U16351 (N_16351,N_16152,N_16076);
nand U16352 (N_16352,N_16211,N_16246);
nand U16353 (N_16353,N_16110,N_16061);
and U16354 (N_16354,N_16064,N_16233);
nand U16355 (N_16355,N_16005,N_16168);
and U16356 (N_16356,N_16106,N_16092);
and U16357 (N_16357,N_16009,N_16238);
xnor U16358 (N_16358,N_16105,N_16087);
xnor U16359 (N_16359,N_16116,N_16135);
xor U16360 (N_16360,N_16240,N_16162);
or U16361 (N_16361,N_16038,N_16078);
nor U16362 (N_16362,N_16223,N_16007);
xnor U16363 (N_16363,N_16055,N_16126);
or U16364 (N_16364,N_16161,N_16057);
xnor U16365 (N_16365,N_16012,N_16146);
or U16366 (N_16366,N_16241,N_16072);
nor U16367 (N_16367,N_16194,N_16160);
or U16368 (N_16368,N_16178,N_16008);
nor U16369 (N_16369,N_16175,N_16019);
and U16370 (N_16370,N_16181,N_16217);
nand U16371 (N_16371,N_16127,N_16158);
or U16372 (N_16372,N_16002,N_16089);
nor U16373 (N_16373,N_16210,N_16107);
nor U16374 (N_16374,N_16198,N_16225);
nor U16375 (N_16375,N_16055,N_16242);
and U16376 (N_16376,N_16018,N_16246);
and U16377 (N_16377,N_16223,N_16138);
nand U16378 (N_16378,N_16205,N_16097);
xnor U16379 (N_16379,N_16098,N_16183);
nand U16380 (N_16380,N_16189,N_16249);
xor U16381 (N_16381,N_16054,N_16140);
nor U16382 (N_16382,N_16181,N_16047);
nand U16383 (N_16383,N_16184,N_16063);
nand U16384 (N_16384,N_16213,N_16243);
xor U16385 (N_16385,N_16198,N_16099);
xor U16386 (N_16386,N_16125,N_16011);
and U16387 (N_16387,N_16092,N_16105);
nor U16388 (N_16388,N_16131,N_16057);
xnor U16389 (N_16389,N_16245,N_16036);
nand U16390 (N_16390,N_16081,N_16009);
or U16391 (N_16391,N_16163,N_16086);
nand U16392 (N_16392,N_16100,N_16093);
nor U16393 (N_16393,N_16020,N_16047);
xnor U16394 (N_16394,N_16069,N_16138);
nand U16395 (N_16395,N_16105,N_16039);
nand U16396 (N_16396,N_16162,N_16191);
xor U16397 (N_16397,N_16064,N_16074);
xnor U16398 (N_16398,N_16054,N_16082);
nor U16399 (N_16399,N_16042,N_16115);
and U16400 (N_16400,N_16189,N_16216);
xnor U16401 (N_16401,N_16230,N_16138);
or U16402 (N_16402,N_16143,N_16064);
nand U16403 (N_16403,N_16020,N_16053);
and U16404 (N_16404,N_16193,N_16083);
and U16405 (N_16405,N_16136,N_16056);
or U16406 (N_16406,N_16244,N_16214);
and U16407 (N_16407,N_16022,N_16042);
or U16408 (N_16408,N_16179,N_16082);
and U16409 (N_16409,N_16040,N_16175);
and U16410 (N_16410,N_16112,N_16119);
nand U16411 (N_16411,N_16054,N_16241);
or U16412 (N_16412,N_16206,N_16226);
or U16413 (N_16413,N_16128,N_16119);
nand U16414 (N_16414,N_16069,N_16063);
and U16415 (N_16415,N_16196,N_16130);
nand U16416 (N_16416,N_16004,N_16084);
nor U16417 (N_16417,N_16213,N_16153);
nor U16418 (N_16418,N_16173,N_16112);
xnor U16419 (N_16419,N_16197,N_16188);
xnor U16420 (N_16420,N_16210,N_16213);
and U16421 (N_16421,N_16120,N_16168);
or U16422 (N_16422,N_16212,N_16054);
nand U16423 (N_16423,N_16151,N_16162);
nor U16424 (N_16424,N_16107,N_16211);
and U16425 (N_16425,N_16030,N_16158);
nor U16426 (N_16426,N_16210,N_16039);
xnor U16427 (N_16427,N_16063,N_16125);
nor U16428 (N_16428,N_16031,N_16013);
nand U16429 (N_16429,N_16086,N_16032);
xnor U16430 (N_16430,N_16216,N_16182);
nand U16431 (N_16431,N_16092,N_16147);
and U16432 (N_16432,N_16083,N_16120);
and U16433 (N_16433,N_16221,N_16064);
and U16434 (N_16434,N_16010,N_16069);
nor U16435 (N_16435,N_16104,N_16068);
nor U16436 (N_16436,N_16175,N_16003);
xor U16437 (N_16437,N_16206,N_16154);
nor U16438 (N_16438,N_16192,N_16101);
or U16439 (N_16439,N_16225,N_16206);
and U16440 (N_16440,N_16166,N_16048);
xor U16441 (N_16441,N_16015,N_16239);
and U16442 (N_16442,N_16027,N_16052);
and U16443 (N_16443,N_16217,N_16022);
or U16444 (N_16444,N_16150,N_16213);
or U16445 (N_16445,N_16163,N_16196);
nand U16446 (N_16446,N_16241,N_16122);
or U16447 (N_16447,N_16117,N_16051);
xnor U16448 (N_16448,N_16171,N_16210);
nand U16449 (N_16449,N_16093,N_16111);
and U16450 (N_16450,N_16002,N_16185);
nand U16451 (N_16451,N_16064,N_16098);
or U16452 (N_16452,N_16015,N_16082);
nor U16453 (N_16453,N_16087,N_16215);
nand U16454 (N_16454,N_16094,N_16169);
xnor U16455 (N_16455,N_16076,N_16227);
nor U16456 (N_16456,N_16196,N_16030);
or U16457 (N_16457,N_16025,N_16199);
or U16458 (N_16458,N_16186,N_16193);
nand U16459 (N_16459,N_16247,N_16181);
nand U16460 (N_16460,N_16203,N_16039);
and U16461 (N_16461,N_16152,N_16249);
or U16462 (N_16462,N_16102,N_16249);
nand U16463 (N_16463,N_16148,N_16233);
nor U16464 (N_16464,N_16081,N_16086);
nand U16465 (N_16465,N_16072,N_16156);
xnor U16466 (N_16466,N_16215,N_16066);
and U16467 (N_16467,N_16185,N_16117);
nand U16468 (N_16468,N_16200,N_16004);
and U16469 (N_16469,N_16179,N_16132);
or U16470 (N_16470,N_16024,N_16022);
nor U16471 (N_16471,N_16124,N_16015);
nor U16472 (N_16472,N_16120,N_16030);
nand U16473 (N_16473,N_16054,N_16147);
nand U16474 (N_16474,N_16142,N_16155);
or U16475 (N_16475,N_16019,N_16027);
xor U16476 (N_16476,N_16155,N_16024);
or U16477 (N_16477,N_16214,N_16106);
nand U16478 (N_16478,N_16033,N_16163);
and U16479 (N_16479,N_16019,N_16140);
nand U16480 (N_16480,N_16034,N_16175);
xor U16481 (N_16481,N_16195,N_16057);
nand U16482 (N_16482,N_16090,N_16244);
nand U16483 (N_16483,N_16007,N_16146);
nand U16484 (N_16484,N_16098,N_16149);
or U16485 (N_16485,N_16141,N_16040);
and U16486 (N_16486,N_16025,N_16214);
xnor U16487 (N_16487,N_16040,N_16162);
or U16488 (N_16488,N_16133,N_16113);
nand U16489 (N_16489,N_16005,N_16103);
nand U16490 (N_16490,N_16083,N_16109);
nand U16491 (N_16491,N_16145,N_16209);
xnor U16492 (N_16492,N_16114,N_16150);
or U16493 (N_16493,N_16177,N_16025);
nand U16494 (N_16494,N_16019,N_16218);
or U16495 (N_16495,N_16073,N_16211);
or U16496 (N_16496,N_16221,N_16236);
and U16497 (N_16497,N_16249,N_16231);
or U16498 (N_16498,N_16209,N_16081);
or U16499 (N_16499,N_16130,N_16109);
xor U16500 (N_16500,N_16259,N_16417);
xor U16501 (N_16501,N_16418,N_16467);
xnor U16502 (N_16502,N_16356,N_16340);
nor U16503 (N_16503,N_16354,N_16473);
nand U16504 (N_16504,N_16435,N_16364);
xor U16505 (N_16505,N_16292,N_16271);
xnor U16506 (N_16506,N_16460,N_16266);
xor U16507 (N_16507,N_16253,N_16365);
or U16508 (N_16508,N_16496,N_16286);
or U16509 (N_16509,N_16359,N_16319);
nand U16510 (N_16510,N_16396,N_16475);
nor U16511 (N_16511,N_16442,N_16438);
and U16512 (N_16512,N_16350,N_16274);
and U16513 (N_16513,N_16324,N_16293);
and U16514 (N_16514,N_16411,N_16329);
nand U16515 (N_16515,N_16287,N_16269);
and U16516 (N_16516,N_16343,N_16332);
nand U16517 (N_16517,N_16457,N_16300);
or U16518 (N_16518,N_16255,N_16497);
nor U16519 (N_16519,N_16367,N_16372);
nand U16520 (N_16520,N_16419,N_16488);
and U16521 (N_16521,N_16303,N_16478);
xnor U16522 (N_16522,N_16377,N_16291);
and U16523 (N_16523,N_16495,N_16383);
and U16524 (N_16524,N_16304,N_16339);
nand U16525 (N_16525,N_16443,N_16468);
nand U16526 (N_16526,N_16470,N_16407);
nor U16527 (N_16527,N_16426,N_16281);
nand U16528 (N_16528,N_16301,N_16391);
nand U16529 (N_16529,N_16461,N_16427);
nor U16530 (N_16530,N_16278,N_16494);
nor U16531 (N_16531,N_16412,N_16401);
nor U16532 (N_16532,N_16260,N_16450);
nor U16533 (N_16533,N_16378,N_16375);
and U16534 (N_16534,N_16446,N_16344);
nand U16535 (N_16535,N_16346,N_16380);
xnor U16536 (N_16536,N_16342,N_16465);
nor U16537 (N_16537,N_16430,N_16458);
or U16538 (N_16538,N_16361,N_16369);
nor U16539 (N_16539,N_16313,N_16479);
or U16540 (N_16540,N_16400,N_16327);
or U16541 (N_16541,N_16337,N_16405);
nor U16542 (N_16542,N_16431,N_16257);
and U16543 (N_16543,N_16408,N_16492);
and U16544 (N_16544,N_16394,N_16264);
xnor U16545 (N_16545,N_16472,N_16330);
nand U16546 (N_16546,N_16444,N_16403);
or U16547 (N_16547,N_16314,N_16452);
nand U16548 (N_16548,N_16288,N_16261);
nand U16549 (N_16549,N_16353,N_16273);
and U16550 (N_16550,N_16390,N_16366);
xor U16551 (N_16551,N_16285,N_16393);
nor U16552 (N_16552,N_16421,N_16316);
nand U16553 (N_16553,N_16436,N_16429);
nand U16554 (N_16554,N_16480,N_16335);
and U16555 (N_16555,N_16382,N_16282);
nand U16556 (N_16556,N_16432,N_16311);
or U16557 (N_16557,N_16464,N_16381);
or U16558 (N_16558,N_16357,N_16491);
nand U16559 (N_16559,N_16395,N_16306);
nand U16560 (N_16560,N_16466,N_16425);
and U16561 (N_16561,N_16420,N_16456);
nor U16562 (N_16562,N_16331,N_16374);
nor U16563 (N_16563,N_16320,N_16336);
xor U16564 (N_16564,N_16447,N_16485);
xor U16565 (N_16565,N_16379,N_16424);
nand U16566 (N_16566,N_16453,N_16258);
or U16567 (N_16567,N_16422,N_16414);
nor U16568 (N_16568,N_16317,N_16323);
nor U16569 (N_16569,N_16384,N_16371);
xnor U16570 (N_16570,N_16283,N_16462);
nor U16571 (N_16571,N_16370,N_16284);
nor U16572 (N_16572,N_16388,N_16402);
xnor U16573 (N_16573,N_16347,N_16483);
nand U16574 (N_16574,N_16275,N_16309);
nor U16575 (N_16575,N_16252,N_16268);
nand U16576 (N_16576,N_16410,N_16459);
and U16577 (N_16577,N_16310,N_16302);
nand U16578 (N_16578,N_16416,N_16440);
xor U16579 (N_16579,N_16349,N_16318);
and U16580 (N_16580,N_16277,N_16263);
nand U16581 (N_16581,N_16490,N_16368);
nor U16582 (N_16582,N_16308,N_16451);
xnor U16583 (N_16583,N_16376,N_16305);
or U16584 (N_16584,N_16386,N_16471);
and U16585 (N_16585,N_16299,N_16449);
nand U16586 (N_16586,N_16295,N_16423);
or U16587 (N_16587,N_16437,N_16250);
and U16588 (N_16588,N_16404,N_16294);
or U16589 (N_16589,N_16351,N_16279);
nand U16590 (N_16590,N_16441,N_16481);
or U16591 (N_16591,N_16484,N_16433);
or U16592 (N_16592,N_16262,N_16315);
and U16593 (N_16593,N_16476,N_16265);
and U16594 (N_16594,N_16358,N_16341);
xnor U16595 (N_16595,N_16387,N_16307);
or U16596 (N_16596,N_16463,N_16454);
nand U16597 (N_16597,N_16321,N_16270);
nor U16598 (N_16598,N_16486,N_16493);
nand U16599 (N_16599,N_16498,N_16333);
or U16600 (N_16600,N_16334,N_16413);
or U16601 (N_16601,N_16428,N_16363);
or U16602 (N_16602,N_16297,N_16397);
and U16603 (N_16603,N_16352,N_16322);
or U16604 (N_16604,N_16434,N_16398);
or U16605 (N_16605,N_16469,N_16373);
nor U16606 (N_16606,N_16276,N_16360);
nand U16607 (N_16607,N_16477,N_16455);
xor U16608 (N_16608,N_16312,N_16362);
nor U16609 (N_16609,N_16256,N_16474);
xnor U16610 (N_16610,N_16448,N_16348);
or U16611 (N_16611,N_16325,N_16482);
or U16612 (N_16612,N_16298,N_16415);
nor U16613 (N_16613,N_16489,N_16326);
nor U16614 (N_16614,N_16392,N_16487);
xor U16615 (N_16615,N_16289,N_16272);
and U16616 (N_16616,N_16385,N_16399);
nor U16617 (N_16617,N_16254,N_16290);
and U16618 (N_16618,N_16251,N_16355);
or U16619 (N_16619,N_16328,N_16267);
nor U16620 (N_16620,N_16406,N_16338);
nand U16621 (N_16621,N_16296,N_16499);
nand U16622 (N_16622,N_16345,N_16280);
nand U16623 (N_16623,N_16409,N_16389);
nor U16624 (N_16624,N_16445,N_16439);
or U16625 (N_16625,N_16276,N_16404);
and U16626 (N_16626,N_16368,N_16403);
and U16627 (N_16627,N_16499,N_16367);
nor U16628 (N_16628,N_16470,N_16398);
xor U16629 (N_16629,N_16364,N_16368);
nand U16630 (N_16630,N_16283,N_16491);
and U16631 (N_16631,N_16420,N_16351);
xor U16632 (N_16632,N_16490,N_16287);
xnor U16633 (N_16633,N_16375,N_16300);
nand U16634 (N_16634,N_16401,N_16380);
and U16635 (N_16635,N_16461,N_16362);
nor U16636 (N_16636,N_16394,N_16438);
nand U16637 (N_16637,N_16430,N_16291);
and U16638 (N_16638,N_16424,N_16290);
nand U16639 (N_16639,N_16307,N_16404);
and U16640 (N_16640,N_16378,N_16428);
or U16641 (N_16641,N_16329,N_16439);
nor U16642 (N_16642,N_16447,N_16436);
nand U16643 (N_16643,N_16432,N_16403);
and U16644 (N_16644,N_16488,N_16399);
nand U16645 (N_16645,N_16325,N_16320);
or U16646 (N_16646,N_16384,N_16485);
and U16647 (N_16647,N_16253,N_16452);
or U16648 (N_16648,N_16373,N_16358);
nor U16649 (N_16649,N_16414,N_16440);
or U16650 (N_16650,N_16430,N_16344);
or U16651 (N_16651,N_16301,N_16367);
xnor U16652 (N_16652,N_16454,N_16325);
nor U16653 (N_16653,N_16277,N_16273);
or U16654 (N_16654,N_16273,N_16325);
xnor U16655 (N_16655,N_16453,N_16490);
nand U16656 (N_16656,N_16499,N_16357);
nor U16657 (N_16657,N_16264,N_16321);
nor U16658 (N_16658,N_16374,N_16372);
nand U16659 (N_16659,N_16290,N_16253);
or U16660 (N_16660,N_16320,N_16266);
or U16661 (N_16661,N_16481,N_16361);
and U16662 (N_16662,N_16289,N_16431);
xor U16663 (N_16663,N_16425,N_16460);
nand U16664 (N_16664,N_16467,N_16334);
xnor U16665 (N_16665,N_16318,N_16467);
or U16666 (N_16666,N_16288,N_16333);
nor U16667 (N_16667,N_16455,N_16483);
nand U16668 (N_16668,N_16473,N_16466);
or U16669 (N_16669,N_16369,N_16338);
nand U16670 (N_16670,N_16411,N_16412);
and U16671 (N_16671,N_16281,N_16324);
or U16672 (N_16672,N_16392,N_16478);
nand U16673 (N_16673,N_16357,N_16289);
xnor U16674 (N_16674,N_16327,N_16309);
and U16675 (N_16675,N_16471,N_16370);
xor U16676 (N_16676,N_16461,N_16331);
nand U16677 (N_16677,N_16343,N_16442);
xor U16678 (N_16678,N_16490,N_16346);
nand U16679 (N_16679,N_16302,N_16402);
or U16680 (N_16680,N_16363,N_16426);
or U16681 (N_16681,N_16439,N_16428);
xor U16682 (N_16682,N_16396,N_16306);
or U16683 (N_16683,N_16276,N_16375);
nor U16684 (N_16684,N_16447,N_16318);
and U16685 (N_16685,N_16370,N_16305);
xnor U16686 (N_16686,N_16470,N_16454);
nor U16687 (N_16687,N_16309,N_16267);
and U16688 (N_16688,N_16314,N_16485);
xnor U16689 (N_16689,N_16376,N_16355);
or U16690 (N_16690,N_16252,N_16463);
nand U16691 (N_16691,N_16338,N_16290);
nand U16692 (N_16692,N_16481,N_16411);
or U16693 (N_16693,N_16300,N_16406);
nand U16694 (N_16694,N_16489,N_16332);
and U16695 (N_16695,N_16277,N_16313);
nand U16696 (N_16696,N_16300,N_16270);
or U16697 (N_16697,N_16483,N_16392);
xor U16698 (N_16698,N_16325,N_16258);
nor U16699 (N_16699,N_16447,N_16411);
or U16700 (N_16700,N_16440,N_16441);
nand U16701 (N_16701,N_16319,N_16470);
or U16702 (N_16702,N_16456,N_16380);
and U16703 (N_16703,N_16301,N_16281);
nand U16704 (N_16704,N_16439,N_16295);
xor U16705 (N_16705,N_16466,N_16307);
nand U16706 (N_16706,N_16418,N_16358);
xnor U16707 (N_16707,N_16363,N_16403);
and U16708 (N_16708,N_16416,N_16276);
xnor U16709 (N_16709,N_16257,N_16267);
and U16710 (N_16710,N_16432,N_16316);
or U16711 (N_16711,N_16339,N_16349);
and U16712 (N_16712,N_16299,N_16440);
or U16713 (N_16713,N_16375,N_16397);
nor U16714 (N_16714,N_16396,N_16313);
xnor U16715 (N_16715,N_16414,N_16408);
nor U16716 (N_16716,N_16494,N_16449);
or U16717 (N_16717,N_16322,N_16362);
and U16718 (N_16718,N_16464,N_16254);
nand U16719 (N_16719,N_16292,N_16486);
nand U16720 (N_16720,N_16461,N_16364);
xor U16721 (N_16721,N_16359,N_16336);
xor U16722 (N_16722,N_16454,N_16362);
nor U16723 (N_16723,N_16434,N_16392);
or U16724 (N_16724,N_16330,N_16451);
or U16725 (N_16725,N_16283,N_16427);
and U16726 (N_16726,N_16464,N_16410);
nor U16727 (N_16727,N_16405,N_16471);
and U16728 (N_16728,N_16413,N_16484);
and U16729 (N_16729,N_16473,N_16362);
or U16730 (N_16730,N_16437,N_16460);
or U16731 (N_16731,N_16250,N_16383);
or U16732 (N_16732,N_16491,N_16479);
or U16733 (N_16733,N_16268,N_16478);
nand U16734 (N_16734,N_16419,N_16456);
nand U16735 (N_16735,N_16438,N_16298);
and U16736 (N_16736,N_16278,N_16270);
nand U16737 (N_16737,N_16258,N_16261);
or U16738 (N_16738,N_16259,N_16276);
nor U16739 (N_16739,N_16386,N_16423);
nand U16740 (N_16740,N_16327,N_16412);
or U16741 (N_16741,N_16389,N_16290);
nand U16742 (N_16742,N_16406,N_16462);
or U16743 (N_16743,N_16275,N_16449);
or U16744 (N_16744,N_16411,N_16486);
or U16745 (N_16745,N_16265,N_16288);
nor U16746 (N_16746,N_16446,N_16314);
nand U16747 (N_16747,N_16488,N_16278);
xor U16748 (N_16748,N_16395,N_16371);
nand U16749 (N_16749,N_16334,N_16385);
or U16750 (N_16750,N_16603,N_16588);
xnor U16751 (N_16751,N_16531,N_16734);
and U16752 (N_16752,N_16727,N_16606);
and U16753 (N_16753,N_16513,N_16635);
or U16754 (N_16754,N_16672,N_16520);
and U16755 (N_16755,N_16579,N_16655);
and U16756 (N_16756,N_16534,N_16566);
or U16757 (N_16757,N_16512,N_16597);
and U16758 (N_16758,N_16506,N_16742);
and U16759 (N_16759,N_16505,N_16714);
or U16760 (N_16760,N_16563,N_16712);
and U16761 (N_16761,N_16745,N_16674);
and U16762 (N_16762,N_16695,N_16507);
or U16763 (N_16763,N_16542,N_16717);
nand U16764 (N_16764,N_16673,N_16740);
nand U16765 (N_16765,N_16592,N_16509);
and U16766 (N_16766,N_16687,N_16557);
or U16767 (N_16767,N_16646,N_16639);
or U16768 (N_16768,N_16739,N_16692);
or U16769 (N_16769,N_16500,N_16626);
nor U16770 (N_16770,N_16558,N_16684);
nor U16771 (N_16771,N_16590,N_16641);
nor U16772 (N_16772,N_16665,N_16585);
and U16773 (N_16773,N_16627,N_16724);
nand U16774 (N_16774,N_16525,N_16581);
nand U16775 (N_16775,N_16618,N_16586);
xnor U16776 (N_16776,N_16656,N_16686);
and U16777 (N_16777,N_16689,N_16600);
xnor U16778 (N_16778,N_16722,N_16576);
and U16779 (N_16779,N_16501,N_16616);
or U16780 (N_16780,N_16544,N_16620);
or U16781 (N_16781,N_16749,N_16550);
nand U16782 (N_16782,N_16703,N_16669);
nor U16783 (N_16783,N_16659,N_16571);
or U16784 (N_16784,N_16664,N_16624);
and U16785 (N_16785,N_16637,N_16629);
xnor U16786 (N_16786,N_16691,N_16632);
or U16787 (N_16787,N_16631,N_16747);
nand U16788 (N_16788,N_16733,N_16519);
nor U16789 (N_16789,N_16560,N_16741);
xnor U16790 (N_16790,N_16526,N_16660);
or U16791 (N_16791,N_16678,N_16716);
nor U16792 (N_16792,N_16648,N_16685);
nand U16793 (N_16793,N_16683,N_16723);
xnor U16794 (N_16794,N_16698,N_16577);
xor U16795 (N_16795,N_16562,N_16622);
nand U16796 (N_16796,N_16609,N_16652);
xor U16797 (N_16797,N_16688,N_16559);
nor U16798 (N_16798,N_16662,N_16548);
and U16799 (N_16799,N_16575,N_16748);
or U16800 (N_16800,N_16541,N_16667);
or U16801 (N_16801,N_16574,N_16681);
and U16802 (N_16802,N_16569,N_16601);
nor U16803 (N_16803,N_16702,N_16595);
and U16804 (N_16804,N_16682,N_16538);
xor U16805 (N_16805,N_16602,N_16584);
or U16806 (N_16806,N_16605,N_16532);
and U16807 (N_16807,N_16504,N_16556);
and U16808 (N_16808,N_16552,N_16594);
xnor U16809 (N_16809,N_16720,N_16610);
or U16810 (N_16810,N_16738,N_16697);
xnor U16811 (N_16811,N_16516,N_16679);
and U16812 (N_16812,N_16699,N_16589);
or U16813 (N_16813,N_16546,N_16653);
nand U16814 (N_16814,N_16708,N_16670);
or U16815 (N_16815,N_16643,N_16677);
nand U16816 (N_16816,N_16573,N_16715);
nand U16817 (N_16817,N_16539,N_16729);
or U16818 (N_16818,N_16568,N_16718);
xnor U16819 (N_16819,N_16696,N_16613);
xor U16820 (N_16820,N_16528,N_16651);
or U16821 (N_16821,N_16658,N_16680);
nand U16822 (N_16822,N_16580,N_16731);
and U16823 (N_16823,N_16649,N_16617);
xnor U16824 (N_16824,N_16633,N_16654);
and U16825 (N_16825,N_16628,N_16604);
nand U16826 (N_16826,N_16510,N_16529);
and U16827 (N_16827,N_16650,N_16675);
nor U16828 (N_16828,N_16593,N_16543);
nand U16829 (N_16829,N_16721,N_16511);
and U16830 (N_16830,N_16596,N_16707);
and U16831 (N_16831,N_16554,N_16582);
or U16832 (N_16832,N_16640,N_16694);
or U16833 (N_16833,N_16737,N_16732);
and U16834 (N_16834,N_16561,N_16636);
nand U16835 (N_16835,N_16551,N_16713);
xnor U16836 (N_16836,N_16705,N_16527);
nor U16837 (N_16837,N_16564,N_16710);
nor U16838 (N_16838,N_16502,N_16642);
and U16839 (N_16839,N_16522,N_16608);
nor U16840 (N_16840,N_16701,N_16518);
nor U16841 (N_16841,N_16693,N_16621);
or U16842 (N_16842,N_16517,N_16666);
nand U16843 (N_16843,N_16700,N_16630);
and U16844 (N_16844,N_16508,N_16545);
nor U16845 (N_16845,N_16725,N_16587);
nor U16846 (N_16846,N_16578,N_16570);
xor U16847 (N_16847,N_16521,N_16547);
nor U16848 (N_16848,N_16555,N_16524);
nand U16849 (N_16849,N_16549,N_16668);
or U16850 (N_16850,N_16535,N_16634);
nand U16851 (N_16851,N_16644,N_16623);
nand U16852 (N_16852,N_16598,N_16638);
or U16853 (N_16853,N_16583,N_16619);
nand U16854 (N_16854,N_16661,N_16530);
nand U16855 (N_16855,N_16746,N_16704);
and U16856 (N_16856,N_16515,N_16663);
xor U16857 (N_16857,N_16514,N_16503);
and U16858 (N_16858,N_16726,N_16743);
and U16859 (N_16859,N_16567,N_16599);
and U16860 (N_16860,N_16565,N_16706);
and U16861 (N_16861,N_16533,N_16728);
or U16862 (N_16862,N_16536,N_16553);
xnor U16863 (N_16863,N_16671,N_16657);
xnor U16864 (N_16864,N_16537,N_16719);
or U16865 (N_16865,N_16625,N_16647);
or U16866 (N_16866,N_16736,N_16591);
nand U16867 (N_16867,N_16709,N_16611);
or U16868 (N_16868,N_16645,N_16615);
or U16869 (N_16869,N_16523,N_16711);
nand U16870 (N_16870,N_16730,N_16735);
nand U16871 (N_16871,N_16614,N_16572);
xnor U16872 (N_16872,N_16607,N_16690);
xor U16873 (N_16873,N_16612,N_16540);
nor U16874 (N_16874,N_16744,N_16676);
and U16875 (N_16875,N_16591,N_16584);
nor U16876 (N_16876,N_16608,N_16540);
nand U16877 (N_16877,N_16719,N_16630);
nand U16878 (N_16878,N_16543,N_16723);
xnor U16879 (N_16879,N_16506,N_16550);
nand U16880 (N_16880,N_16522,N_16602);
nor U16881 (N_16881,N_16696,N_16650);
xnor U16882 (N_16882,N_16607,N_16559);
nor U16883 (N_16883,N_16576,N_16687);
nor U16884 (N_16884,N_16647,N_16502);
or U16885 (N_16885,N_16526,N_16588);
xnor U16886 (N_16886,N_16744,N_16693);
or U16887 (N_16887,N_16737,N_16676);
and U16888 (N_16888,N_16734,N_16513);
and U16889 (N_16889,N_16693,N_16612);
or U16890 (N_16890,N_16687,N_16592);
or U16891 (N_16891,N_16529,N_16644);
xnor U16892 (N_16892,N_16582,N_16542);
nor U16893 (N_16893,N_16664,N_16627);
nor U16894 (N_16894,N_16673,N_16549);
xnor U16895 (N_16895,N_16632,N_16548);
nor U16896 (N_16896,N_16526,N_16585);
nor U16897 (N_16897,N_16511,N_16684);
nand U16898 (N_16898,N_16644,N_16537);
or U16899 (N_16899,N_16619,N_16629);
xor U16900 (N_16900,N_16512,N_16605);
and U16901 (N_16901,N_16556,N_16732);
nand U16902 (N_16902,N_16561,N_16556);
or U16903 (N_16903,N_16541,N_16526);
nor U16904 (N_16904,N_16702,N_16740);
nand U16905 (N_16905,N_16544,N_16613);
xnor U16906 (N_16906,N_16624,N_16702);
or U16907 (N_16907,N_16500,N_16510);
or U16908 (N_16908,N_16708,N_16667);
xor U16909 (N_16909,N_16578,N_16571);
nand U16910 (N_16910,N_16748,N_16696);
nor U16911 (N_16911,N_16664,N_16638);
or U16912 (N_16912,N_16557,N_16543);
xnor U16913 (N_16913,N_16538,N_16679);
and U16914 (N_16914,N_16746,N_16637);
nand U16915 (N_16915,N_16680,N_16673);
or U16916 (N_16916,N_16572,N_16657);
nor U16917 (N_16917,N_16534,N_16554);
nor U16918 (N_16918,N_16579,N_16568);
nand U16919 (N_16919,N_16590,N_16538);
nor U16920 (N_16920,N_16569,N_16678);
nand U16921 (N_16921,N_16587,N_16574);
nand U16922 (N_16922,N_16694,N_16513);
xor U16923 (N_16923,N_16724,N_16682);
nor U16924 (N_16924,N_16604,N_16595);
and U16925 (N_16925,N_16584,N_16509);
or U16926 (N_16926,N_16666,N_16544);
xor U16927 (N_16927,N_16700,N_16549);
and U16928 (N_16928,N_16621,N_16577);
and U16929 (N_16929,N_16628,N_16582);
xnor U16930 (N_16930,N_16645,N_16722);
nand U16931 (N_16931,N_16528,N_16605);
nor U16932 (N_16932,N_16732,N_16739);
and U16933 (N_16933,N_16682,N_16610);
xnor U16934 (N_16934,N_16675,N_16606);
nor U16935 (N_16935,N_16623,N_16656);
nor U16936 (N_16936,N_16667,N_16723);
or U16937 (N_16937,N_16592,N_16538);
nand U16938 (N_16938,N_16564,N_16619);
or U16939 (N_16939,N_16653,N_16687);
or U16940 (N_16940,N_16597,N_16509);
and U16941 (N_16941,N_16725,N_16701);
and U16942 (N_16942,N_16578,N_16560);
or U16943 (N_16943,N_16672,N_16616);
and U16944 (N_16944,N_16605,N_16731);
xnor U16945 (N_16945,N_16679,N_16657);
and U16946 (N_16946,N_16745,N_16691);
nor U16947 (N_16947,N_16745,N_16553);
nand U16948 (N_16948,N_16719,N_16728);
xnor U16949 (N_16949,N_16585,N_16674);
nand U16950 (N_16950,N_16665,N_16592);
xnor U16951 (N_16951,N_16541,N_16651);
nor U16952 (N_16952,N_16605,N_16539);
or U16953 (N_16953,N_16688,N_16509);
and U16954 (N_16954,N_16668,N_16648);
nor U16955 (N_16955,N_16632,N_16506);
nor U16956 (N_16956,N_16709,N_16695);
or U16957 (N_16957,N_16685,N_16654);
and U16958 (N_16958,N_16550,N_16627);
nor U16959 (N_16959,N_16694,N_16500);
xnor U16960 (N_16960,N_16626,N_16674);
and U16961 (N_16961,N_16736,N_16739);
nor U16962 (N_16962,N_16545,N_16739);
nand U16963 (N_16963,N_16538,N_16685);
and U16964 (N_16964,N_16609,N_16612);
or U16965 (N_16965,N_16713,N_16681);
or U16966 (N_16966,N_16590,N_16743);
and U16967 (N_16967,N_16606,N_16580);
nor U16968 (N_16968,N_16511,N_16661);
nand U16969 (N_16969,N_16576,N_16645);
nor U16970 (N_16970,N_16550,N_16511);
and U16971 (N_16971,N_16720,N_16717);
nor U16972 (N_16972,N_16663,N_16526);
xor U16973 (N_16973,N_16629,N_16581);
nor U16974 (N_16974,N_16554,N_16530);
or U16975 (N_16975,N_16733,N_16704);
and U16976 (N_16976,N_16720,N_16748);
or U16977 (N_16977,N_16657,N_16686);
and U16978 (N_16978,N_16536,N_16586);
nand U16979 (N_16979,N_16626,N_16715);
and U16980 (N_16980,N_16571,N_16703);
nand U16981 (N_16981,N_16685,N_16580);
nor U16982 (N_16982,N_16618,N_16691);
or U16983 (N_16983,N_16542,N_16590);
or U16984 (N_16984,N_16538,N_16580);
and U16985 (N_16985,N_16674,N_16605);
nor U16986 (N_16986,N_16581,N_16671);
nor U16987 (N_16987,N_16578,N_16692);
nor U16988 (N_16988,N_16634,N_16709);
nor U16989 (N_16989,N_16610,N_16705);
nand U16990 (N_16990,N_16570,N_16705);
or U16991 (N_16991,N_16730,N_16737);
nand U16992 (N_16992,N_16707,N_16549);
nor U16993 (N_16993,N_16680,N_16728);
nor U16994 (N_16994,N_16535,N_16709);
and U16995 (N_16995,N_16507,N_16679);
or U16996 (N_16996,N_16642,N_16559);
nand U16997 (N_16997,N_16520,N_16630);
xor U16998 (N_16998,N_16702,N_16638);
nand U16999 (N_16999,N_16611,N_16620);
and U17000 (N_17000,N_16991,N_16837);
or U17001 (N_17001,N_16851,N_16882);
or U17002 (N_17002,N_16914,N_16905);
nor U17003 (N_17003,N_16907,N_16951);
or U17004 (N_17004,N_16777,N_16885);
nor U17005 (N_17005,N_16989,N_16829);
nand U17006 (N_17006,N_16821,N_16852);
and U17007 (N_17007,N_16874,N_16976);
xor U17008 (N_17008,N_16759,N_16928);
nand U17009 (N_17009,N_16795,N_16940);
xor U17010 (N_17010,N_16901,N_16854);
xnor U17011 (N_17011,N_16835,N_16938);
nor U17012 (N_17012,N_16894,N_16988);
xor U17013 (N_17013,N_16983,N_16809);
nand U17014 (N_17014,N_16958,N_16955);
xor U17015 (N_17015,N_16784,N_16872);
nand U17016 (N_17016,N_16847,N_16825);
or U17017 (N_17017,N_16814,N_16838);
nand U17018 (N_17018,N_16915,N_16775);
nor U17019 (N_17019,N_16933,N_16819);
nand U17020 (N_17020,N_16880,N_16945);
nor U17021 (N_17021,N_16798,N_16956);
nor U17022 (N_17022,N_16879,N_16753);
nand U17023 (N_17023,N_16927,N_16785);
or U17024 (N_17024,N_16779,N_16985);
nor U17025 (N_17025,N_16817,N_16808);
or U17026 (N_17026,N_16805,N_16974);
nand U17027 (N_17027,N_16755,N_16815);
and U17028 (N_17028,N_16919,N_16754);
or U17029 (N_17029,N_16833,N_16950);
xor U17030 (N_17030,N_16920,N_16972);
nand U17031 (N_17031,N_16865,N_16922);
or U17032 (N_17032,N_16776,N_16994);
and U17033 (N_17033,N_16918,N_16890);
and U17034 (N_17034,N_16772,N_16791);
and U17035 (N_17035,N_16900,N_16960);
or U17036 (N_17036,N_16813,N_16869);
nor U17037 (N_17037,N_16782,N_16886);
xor U17038 (N_17038,N_16980,N_16926);
nor U17039 (N_17039,N_16966,N_16764);
and U17040 (N_17040,N_16765,N_16923);
or U17041 (N_17041,N_16816,N_16771);
nor U17042 (N_17042,N_16987,N_16954);
nand U17043 (N_17043,N_16868,N_16939);
or U17044 (N_17044,N_16977,N_16761);
nand U17045 (N_17045,N_16892,N_16902);
xor U17046 (N_17046,N_16799,N_16936);
xnor U17047 (N_17047,N_16864,N_16778);
or U17048 (N_17048,N_16909,N_16804);
nor U17049 (N_17049,N_16946,N_16986);
and U17050 (N_17050,N_16858,N_16971);
nor U17051 (N_17051,N_16783,N_16766);
xnor U17052 (N_17052,N_16916,N_16959);
xor U17053 (N_17053,N_16937,N_16999);
and U17054 (N_17054,N_16982,N_16873);
nor U17055 (N_17055,N_16803,N_16820);
xnor U17056 (N_17056,N_16877,N_16767);
and U17057 (N_17057,N_16859,N_16929);
nor U17058 (N_17058,N_16881,N_16866);
nor U17059 (N_17059,N_16963,N_16786);
or U17060 (N_17060,N_16893,N_16981);
nand U17061 (N_17061,N_16921,N_16850);
xnor U17062 (N_17062,N_16973,N_16952);
and U17063 (N_17063,N_16830,N_16789);
and U17064 (N_17064,N_16912,N_16845);
and U17065 (N_17065,N_16811,N_16968);
and U17066 (N_17066,N_16796,N_16773);
nand U17067 (N_17067,N_16787,N_16870);
nand U17068 (N_17068,N_16806,N_16895);
and U17069 (N_17069,N_16975,N_16997);
nor U17070 (N_17070,N_16807,N_16843);
nand U17071 (N_17071,N_16832,N_16910);
nand U17072 (N_17072,N_16935,N_16941);
nand U17073 (N_17073,N_16883,N_16948);
nand U17074 (N_17074,N_16932,N_16797);
xnor U17075 (N_17075,N_16792,N_16762);
nor U17076 (N_17076,N_16908,N_16993);
and U17077 (N_17077,N_16824,N_16949);
or U17078 (N_17078,N_16970,N_16943);
nand U17079 (N_17079,N_16758,N_16889);
or U17080 (N_17080,N_16842,N_16930);
nand U17081 (N_17081,N_16800,N_16917);
nand U17082 (N_17082,N_16757,N_16978);
or U17083 (N_17083,N_16995,N_16760);
xnor U17084 (N_17084,N_16992,N_16961);
xor U17085 (N_17085,N_16867,N_16823);
nor U17086 (N_17086,N_16840,N_16953);
and U17087 (N_17087,N_16887,N_16876);
and U17088 (N_17088,N_16856,N_16860);
or U17089 (N_17089,N_16898,N_16841);
xnor U17090 (N_17090,N_16770,N_16944);
xor U17091 (N_17091,N_16810,N_16878);
nand U17092 (N_17092,N_16861,N_16855);
or U17093 (N_17093,N_16844,N_16931);
or U17094 (N_17094,N_16793,N_16990);
nand U17095 (N_17095,N_16768,N_16863);
nor U17096 (N_17096,N_16846,N_16903);
nand U17097 (N_17097,N_16862,N_16853);
nor U17098 (N_17098,N_16947,N_16834);
nor U17099 (N_17099,N_16964,N_16871);
nor U17100 (N_17100,N_16801,N_16848);
and U17101 (N_17101,N_16774,N_16812);
nand U17102 (N_17102,N_16996,N_16788);
or U17103 (N_17103,N_16924,N_16934);
nor U17104 (N_17104,N_16899,N_16969);
nand U17105 (N_17105,N_16828,N_16849);
xnor U17106 (N_17106,N_16818,N_16911);
and U17107 (N_17107,N_16884,N_16790);
and U17108 (N_17108,N_16802,N_16984);
xnor U17109 (N_17109,N_16836,N_16752);
and U17110 (N_17110,N_16962,N_16857);
xnor U17111 (N_17111,N_16780,N_16875);
nor U17112 (N_17112,N_16998,N_16794);
and U17113 (N_17113,N_16957,N_16979);
and U17114 (N_17114,N_16826,N_16831);
nor U17115 (N_17115,N_16763,N_16942);
xnor U17116 (N_17116,N_16897,N_16925);
nand U17117 (N_17117,N_16891,N_16750);
and U17118 (N_17118,N_16781,N_16827);
nor U17119 (N_17119,N_16839,N_16906);
nand U17120 (N_17120,N_16756,N_16751);
or U17121 (N_17121,N_16967,N_16769);
nor U17122 (N_17122,N_16888,N_16965);
nand U17123 (N_17123,N_16822,N_16913);
and U17124 (N_17124,N_16904,N_16896);
or U17125 (N_17125,N_16970,N_16888);
or U17126 (N_17126,N_16833,N_16852);
xor U17127 (N_17127,N_16956,N_16851);
or U17128 (N_17128,N_16820,N_16899);
xnor U17129 (N_17129,N_16868,N_16836);
nand U17130 (N_17130,N_16814,N_16828);
or U17131 (N_17131,N_16897,N_16885);
nor U17132 (N_17132,N_16857,N_16922);
or U17133 (N_17133,N_16817,N_16784);
or U17134 (N_17134,N_16981,N_16967);
nor U17135 (N_17135,N_16798,N_16953);
xor U17136 (N_17136,N_16775,N_16863);
xor U17137 (N_17137,N_16826,N_16960);
nor U17138 (N_17138,N_16900,N_16764);
nand U17139 (N_17139,N_16872,N_16793);
and U17140 (N_17140,N_16785,N_16932);
and U17141 (N_17141,N_16966,N_16911);
nand U17142 (N_17142,N_16919,N_16774);
or U17143 (N_17143,N_16960,N_16843);
nor U17144 (N_17144,N_16791,N_16927);
xnor U17145 (N_17145,N_16769,N_16981);
and U17146 (N_17146,N_16787,N_16951);
nor U17147 (N_17147,N_16877,N_16776);
nand U17148 (N_17148,N_16936,N_16912);
nor U17149 (N_17149,N_16829,N_16971);
nor U17150 (N_17150,N_16942,N_16774);
and U17151 (N_17151,N_16866,N_16908);
nor U17152 (N_17152,N_16954,N_16949);
nor U17153 (N_17153,N_16761,N_16880);
and U17154 (N_17154,N_16822,N_16763);
xnor U17155 (N_17155,N_16850,N_16824);
nor U17156 (N_17156,N_16781,N_16830);
xnor U17157 (N_17157,N_16884,N_16791);
or U17158 (N_17158,N_16802,N_16796);
nand U17159 (N_17159,N_16878,N_16945);
and U17160 (N_17160,N_16877,N_16987);
or U17161 (N_17161,N_16947,N_16760);
and U17162 (N_17162,N_16852,N_16854);
nand U17163 (N_17163,N_16870,N_16766);
nand U17164 (N_17164,N_16895,N_16979);
or U17165 (N_17165,N_16853,N_16842);
and U17166 (N_17166,N_16863,N_16841);
nor U17167 (N_17167,N_16982,N_16976);
nor U17168 (N_17168,N_16756,N_16785);
nand U17169 (N_17169,N_16859,N_16771);
and U17170 (N_17170,N_16812,N_16890);
xnor U17171 (N_17171,N_16913,N_16875);
and U17172 (N_17172,N_16918,N_16878);
nor U17173 (N_17173,N_16892,N_16937);
or U17174 (N_17174,N_16863,N_16946);
nand U17175 (N_17175,N_16861,N_16987);
nor U17176 (N_17176,N_16882,N_16784);
and U17177 (N_17177,N_16971,N_16770);
nand U17178 (N_17178,N_16905,N_16978);
nor U17179 (N_17179,N_16961,N_16801);
and U17180 (N_17180,N_16901,N_16858);
nor U17181 (N_17181,N_16917,N_16818);
and U17182 (N_17182,N_16911,N_16808);
or U17183 (N_17183,N_16967,N_16933);
xnor U17184 (N_17184,N_16853,N_16803);
or U17185 (N_17185,N_16774,N_16799);
nor U17186 (N_17186,N_16951,N_16784);
nor U17187 (N_17187,N_16939,N_16828);
xor U17188 (N_17188,N_16905,N_16866);
or U17189 (N_17189,N_16942,N_16925);
or U17190 (N_17190,N_16781,N_16809);
and U17191 (N_17191,N_16834,N_16941);
nor U17192 (N_17192,N_16798,N_16976);
or U17193 (N_17193,N_16879,N_16811);
nor U17194 (N_17194,N_16868,N_16941);
nand U17195 (N_17195,N_16797,N_16956);
xor U17196 (N_17196,N_16793,N_16751);
nor U17197 (N_17197,N_16950,N_16946);
and U17198 (N_17198,N_16792,N_16980);
and U17199 (N_17199,N_16799,N_16865);
or U17200 (N_17200,N_16796,N_16772);
or U17201 (N_17201,N_16831,N_16829);
and U17202 (N_17202,N_16965,N_16758);
nand U17203 (N_17203,N_16780,N_16965);
and U17204 (N_17204,N_16996,N_16791);
and U17205 (N_17205,N_16755,N_16955);
nand U17206 (N_17206,N_16834,N_16976);
or U17207 (N_17207,N_16874,N_16999);
or U17208 (N_17208,N_16943,N_16852);
xor U17209 (N_17209,N_16847,N_16930);
xor U17210 (N_17210,N_16957,N_16836);
or U17211 (N_17211,N_16874,N_16833);
nor U17212 (N_17212,N_16881,N_16790);
or U17213 (N_17213,N_16986,N_16780);
and U17214 (N_17214,N_16879,N_16844);
or U17215 (N_17215,N_16851,N_16886);
xor U17216 (N_17216,N_16825,N_16798);
nor U17217 (N_17217,N_16985,N_16919);
and U17218 (N_17218,N_16816,N_16948);
nor U17219 (N_17219,N_16851,N_16885);
or U17220 (N_17220,N_16868,N_16753);
and U17221 (N_17221,N_16779,N_16752);
nand U17222 (N_17222,N_16813,N_16877);
or U17223 (N_17223,N_16756,N_16984);
and U17224 (N_17224,N_16834,N_16888);
or U17225 (N_17225,N_16752,N_16815);
and U17226 (N_17226,N_16790,N_16848);
nand U17227 (N_17227,N_16831,N_16907);
nand U17228 (N_17228,N_16926,N_16868);
nor U17229 (N_17229,N_16912,N_16969);
and U17230 (N_17230,N_16928,N_16899);
or U17231 (N_17231,N_16908,N_16758);
xor U17232 (N_17232,N_16847,N_16751);
and U17233 (N_17233,N_16954,N_16913);
nor U17234 (N_17234,N_16859,N_16831);
or U17235 (N_17235,N_16812,N_16993);
xor U17236 (N_17236,N_16941,N_16840);
nand U17237 (N_17237,N_16764,N_16792);
xor U17238 (N_17238,N_16822,N_16771);
xor U17239 (N_17239,N_16865,N_16894);
nor U17240 (N_17240,N_16994,N_16964);
xor U17241 (N_17241,N_16753,N_16775);
xor U17242 (N_17242,N_16796,N_16880);
and U17243 (N_17243,N_16786,N_16911);
nor U17244 (N_17244,N_16997,N_16771);
xnor U17245 (N_17245,N_16922,N_16917);
nor U17246 (N_17246,N_16834,N_16868);
or U17247 (N_17247,N_16870,N_16894);
nor U17248 (N_17248,N_16937,N_16907);
nand U17249 (N_17249,N_16963,N_16839);
nor U17250 (N_17250,N_17012,N_17135);
and U17251 (N_17251,N_17030,N_17022);
or U17252 (N_17252,N_17039,N_17128);
nor U17253 (N_17253,N_17049,N_17242);
nand U17254 (N_17254,N_17051,N_17183);
or U17255 (N_17255,N_17021,N_17087);
xor U17256 (N_17256,N_17155,N_17052);
or U17257 (N_17257,N_17102,N_17129);
nand U17258 (N_17258,N_17216,N_17248);
nand U17259 (N_17259,N_17027,N_17240);
xor U17260 (N_17260,N_17145,N_17215);
nor U17261 (N_17261,N_17076,N_17222);
and U17262 (N_17262,N_17169,N_17034);
xor U17263 (N_17263,N_17032,N_17249);
nand U17264 (N_17264,N_17127,N_17223);
or U17265 (N_17265,N_17098,N_17139);
or U17266 (N_17266,N_17202,N_17028);
nor U17267 (N_17267,N_17175,N_17066);
and U17268 (N_17268,N_17208,N_17213);
and U17269 (N_17269,N_17130,N_17020);
xor U17270 (N_17270,N_17109,N_17173);
or U17271 (N_17271,N_17064,N_17042);
nand U17272 (N_17272,N_17225,N_17170);
and U17273 (N_17273,N_17118,N_17189);
nand U17274 (N_17274,N_17153,N_17245);
or U17275 (N_17275,N_17138,N_17046);
and U17276 (N_17276,N_17069,N_17158);
xor U17277 (N_17277,N_17044,N_17013);
xnor U17278 (N_17278,N_17017,N_17073);
and U17279 (N_17279,N_17195,N_17119);
and U17280 (N_17280,N_17019,N_17234);
xor U17281 (N_17281,N_17081,N_17162);
nor U17282 (N_17282,N_17115,N_17241);
xor U17283 (N_17283,N_17203,N_17116);
and U17284 (N_17284,N_17220,N_17057);
or U17285 (N_17285,N_17065,N_17163);
or U17286 (N_17286,N_17210,N_17229);
nand U17287 (N_17287,N_17078,N_17071);
xor U17288 (N_17288,N_17094,N_17205);
xor U17289 (N_17289,N_17089,N_17166);
xnor U17290 (N_17290,N_17218,N_17141);
nor U17291 (N_17291,N_17113,N_17157);
or U17292 (N_17292,N_17137,N_17001);
or U17293 (N_17293,N_17181,N_17111);
nand U17294 (N_17294,N_17201,N_17146);
and U17295 (N_17295,N_17009,N_17231);
xor U17296 (N_17296,N_17077,N_17184);
and U17297 (N_17297,N_17041,N_17165);
nor U17298 (N_17298,N_17082,N_17004);
xnor U17299 (N_17299,N_17151,N_17054);
and U17300 (N_17300,N_17075,N_17024);
or U17301 (N_17301,N_17136,N_17230);
and U17302 (N_17302,N_17095,N_17224);
or U17303 (N_17303,N_17209,N_17148);
and U17304 (N_17304,N_17172,N_17226);
nor U17305 (N_17305,N_17010,N_17074);
and U17306 (N_17306,N_17134,N_17038);
xnor U17307 (N_17307,N_17047,N_17025);
nor U17308 (N_17308,N_17164,N_17133);
xnor U17309 (N_17309,N_17238,N_17015);
xnor U17310 (N_17310,N_17110,N_17221);
xnor U17311 (N_17311,N_17171,N_17011);
xnor U17312 (N_17312,N_17217,N_17100);
and U17313 (N_17313,N_17131,N_17000);
xnor U17314 (N_17314,N_17103,N_17033);
xor U17315 (N_17315,N_17232,N_17228);
xnor U17316 (N_17316,N_17104,N_17026);
xor U17317 (N_17317,N_17187,N_17114);
xnor U17318 (N_17318,N_17008,N_17196);
xnor U17319 (N_17319,N_17006,N_17227);
or U17320 (N_17320,N_17186,N_17126);
xnor U17321 (N_17321,N_17177,N_17058);
xor U17322 (N_17322,N_17150,N_17096);
nand U17323 (N_17323,N_17043,N_17197);
nand U17324 (N_17324,N_17093,N_17191);
and U17325 (N_17325,N_17085,N_17056);
and U17326 (N_17326,N_17045,N_17060);
nand U17327 (N_17327,N_17239,N_17036);
and U17328 (N_17328,N_17003,N_17244);
nor U17329 (N_17329,N_17160,N_17031);
nand U17330 (N_17330,N_17178,N_17080);
and U17331 (N_17331,N_17007,N_17117);
or U17332 (N_17332,N_17053,N_17108);
xnor U17333 (N_17333,N_17105,N_17237);
nor U17334 (N_17334,N_17088,N_17005);
or U17335 (N_17335,N_17067,N_17040);
nand U17336 (N_17336,N_17243,N_17185);
xnor U17337 (N_17337,N_17192,N_17207);
xor U17338 (N_17338,N_17143,N_17188);
nand U17339 (N_17339,N_17091,N_17159);
and U17340 (N_17340,N_17206,N_17048);
or U17341 (N_17341,N_17016,N_17101);
or U17342 (N_17342,N_17132,N_17023);
nor U17343 (N_17343,N_17063,N_17092);
and U17344 (N_17344,N_17122,N_17140);
nand U17345 (N_17345,N_17125,N_17212);
or U17346 (N_17346,N_17083,N_17154);
nand U17347 (N_17347,N_17142,N_17193);
nor U17348 (N_17348,N_17084,N_17182);
nand U17349 (N_17349,N_17097,N_17214);
nand U17350 (N_17350,N_17070,N_17180);
or U17351 (N_17351,N_17176,N_17121);
nand U17352 (N_17352,N_17200,N_17194);
and U17353 (N_17353,N_17090,N_17029);
and U17354 (N_17354,N_17247,N_17035);
xor U17355 (N_17355,N_17168,N_17002);
and U17356 (N_17356,N_17219,N_17161);
nor U17357 (N_17357,N_17068,N_17152);
nor U17358 (N_17358,N_17112,N_17086);
or U17359 (N_17359,N_17072,N_17179);
nand U17360 (N_17360,N_17199,N_17149);
or U17361 (N_17361,N_17156,N_17211);
or U17362 (N_17362,N_17235,N_17167);
nand U17363 (N_17363,N_17079,N_17147);
nand U17364 (N_17364,N_17120,N_17014);
nor U17365 (N_17365,N_17059,N_17061);
xnor U17366 (N_17366,N_17124,N_17107);
nor U17367 (N_17367,N_17144,N_17204);
and U17368 (N_17368,N_17062,N_17174);
and U17369 (N_17369,N_17037,N_17018);
and U17370 (N_17370,N_17123,N_17190);
xor U17371 (N_17371,N_17236,N_17233);
and U17372 (N_17372,N_17055,N_17246);
and U17373 (N_17373,N_17099,N_17106);
xnor U17374 (N_17374,N_17198,N_17050);
xnor U17375 (N_17375,N_17189,N_17201);
xnor U17376 (N_17376,N_17143,N_17035);
nor U17377 (N_17377,N_17227,N_17180);
or U17378 (N_17378,N_17164,N_17066);
or U17379 (N_17379,N_17133,N_17143);
and U17380 (N_17380,N_17242,N_17100);
and U17381 (N_17381,N_17043,N_17131);
xor U17382 (N_17382,N_17038,N_17159);
nor U17383 (N_17383,N_17245,N_17179);
xor U17384 (N_17384,N_17101,N_17032);
nor U17385 (N_17385,N_17137,N_17083);
xnor U17386 (N_17386,N_17054,N_17190);
nor U17387 (N_17387,N_17037,N_17008);
nor U17388 (N_17388,N_17049,N_17139);
and U17389 (N_17389,N_17219,N_17016);
nor U17390 (N_17390,N_17182,N_17045);
nor U17391 (N_17391,N_17011,N_17090);
nor U17392 (N_17392,N_17006,N_17206);
or U17393 (N_17393,N_17191,N_17119);
or U17394 (N_17394,N_17025,N_17152);
nand U17395 (N_17395,N_17068,N_17069);
or U17396 (N_17396,N_17077,N_17230);
xor U17397 (N_17397,N_17025,N_17098);
and U17398 (N_17398,N_17055,N_17058);
xnor U17399 (N_17399,N_17082,N_17197);
xnor U17400 (N_17400,N_17013,N_17017);
xnor U17401 (N_17401,N_17131,N_17127);
or U17402 (N_17402,N_17178,N_17243);
xnor U17403 (N_17403,N_17112,N_17047);
nand U17404 (N_17404,N_17232,N_17217);
and U17405 (N_17405,N_17169,N_17090);
or U17406 (N_17406,N_17048,N_17181);
nor U17407 (N_17407,N_17153,N_17055);
nand U17408 (N_17408,N_17036,N_17024);
and U17409 (N_17409,N_17113,N_17078);
nand U17410 (N_17410,N_17094,N_17163);
and U17411 (N_17411,N_17087,N_17047);
nor U17412 (N_17412,N_17128,N_17202);
and U17413 (N_17413,N_17248,N_17176);
xnor U17414 (N_17414,N_17036,N_17049);
and U17415 (N_17415,N_17185,N_17127);
xnor U17416 (N_17416,N_17172,N_17168);
or U17417 (N_17417,N_17111,N_17065);
or U17418 (N_17418,N_17089,N_17053);
nand U17419 (N_17419,N_17224,N_17006);
or U17420 (N_17420,N_17104,N_17129);
or U17421 (N_17421,N_17049,N_17020);
and U17422 (N_17422,N_17206,N_17111);
nand U17423 (N_17423,N_17178,N_17238);
nor U17424 (N_17424,N_17160,N_17123);
and U17425 (N_17425,N_17037,N_17177);
nor U17426 (N_17426,N_17159,N_17081);
xor U17427 (N_17427,N_17094,N_17010);
nor U17428 (N_17428,N_17134,N_17086);
nor U17429 (N_17429,N_17046,N_17121);
xnor U17430 (N_17430,N_17068,N_17053);
or U17431 (N_17431,N_17032,N_17045);
and U17432 (N_17432,N_17079,N_17220);
or U17433 (N_17433,N_17155,N_17013);
nand U17434 (N_17434,N_17215,N_17210);
xor U17435 (N_17435,N_17018,N_17147);
or U17436 (N_17436,N_17072,N_17221);
or U17437 (N_17437,N_17105,N_17249);
and U17438 (N_17438,N_17119,N_17113);
nor U17439 (N_17439,N_17236,N_17218);
nand U17440 (N_17440,N_17119,N_17050);
xnor U17441 (N_17441,N_17210,N_17114);
nor U17442 (N_17442,N_17132,N_17042);
and U17443 (N_17443,N_17083,N_17097);
nor U17444 (N_17444,N_17068,N_17073);
xnor U17445 (N_17445,N_17132,N_17171);
and U17446 (N_17446,N_17201,N_17119);
nand U17447 (N_17447,N_17174,N_17240);
nor U17448 (N_17448,N_17170,N_17146);
or U17449 (N_17449,N_17011,N_17065);
nand U17450 (N_17450,N_17206,N_17001);
or U17451 (N_17451,N_17009,N_17111);
and U17452 (N_17452,N_17057,N_17110);
and U17453 (N_17453,N_17211,N_17019);
xor U17454 (N_17454,N_17049,N_17088);
nand U17455 (N_17455,N_17133,N_17220);
or U17456 (N_17456,N_17151,N_17100);
and U17457 (N_17457,N_17193,N_17150);
xor U17458 (N_17458,N_17033,N_17086);
nor U17459 (N_17459,N_17069,N_17227);
or U17460 (N_17460,N_17057,N_17213);
nand U17461 (N_17461,N_17229,N_17240);
xnor U17462 (N_17462,N_17130,N_17161);
or U17463 (N_17463,N_17197,N_17168);
and U17464 (N_17464,N_17006,N_17011);
nor U17465 (N_17465,N_17240,N_17202);
or U17466 (N_17466,N_17102,N_17105);
nand U17467 (N_17467,N_17079,N_17121);
xnor U17468 (N_17468,N_17167,N_17176);
xor U17469 (N_17469,N_17047,N_17224);
xor U17470 (N_17470,N_17229,N_17004);
or U17471 (N_17471,N_17226,N_17220);
xnor U17472 (N_17472,N_17001,N_17200);
nor U17473 (N_17473,N_17173,N_17162);
and U17474 (N_17474,N_17064,N_17084);
nor U17475 (N_17475,N_17067,N_17058);
and U17476 (N_17476,N_17235,N_17017);
xor U17477 (N_17477,N_17241,N_17055);
or U17478 (N_17478,N_17122,N_17060);
nand U17479 (N_17479,N_17035,N_17118);
nor U17480 (N_17480,N_17190,N_17110);
or U17481 (N_17481,N_17225,N_17150);
nand U17482 (N_17482,N_17236,N_17131);
and U17483 (N_17483,N_17232,N_17050);
xor U17484 (N_17484,N_17126,N_17165);
nor U17485 (N_17485,N_17184,N_17048);
or U17486 (N_17486,N_17191,N_17018);
nand U17487 (N_17487,N_17035,N_17094);
nor U17488 (N_17488,N_17191,N_17189);
nor U17489 (N_17489,N_17231,N_17230);
xnor U17490 (N_17490,N_17195,N_17173);
and U17491 (N_17491,N_17109,N_17202);
nor U17492 (N_17492,N_17016,N_17222);
xnor U17493 (N_17493,N_17239,N_17001);
and U17494 (N_17494,N_17203,N_17220);
xnor U17495 (N_17495,N_17014,N_17078);
nor U17496 (N_17496,N_17146,N_17218);
and U17497 (N_17497,N_17058,N_17207);
nor U17498 (N_17498,N_17031,N_17193);
and U17499 (N_17499,N_17003,N_17128);
nand U17500 (N_17500,N_17354,N_17250);
xnor U17501 (N_17501,N_17465,N_17456);
and U17502 (N_17502,N_17454,N_17450);
nand U17503 (N_17503,N_17378,N_17269);
and U17504 (N_17504,N_17424,N_17471);
nor U17505 (N_17505,N_17265,N_17444);
and U17506 (N_17506,N_17253,N_17370);
and U17507 (N_17507,N_17286,N_17305);
nor U17508 (N_17508,N_17473,N_17469);
or U17509 (N_17509,N_17458,N_17295);
nand U17510 (N_17510,N_17492,N_17396);
nor U17511 (N_17511,N_17292,N_17393);
xor U17512 (N_17512,N_17421,N_17383);
or U17513 (N_17513,N_17470,N_17384);
or U17514 (N_17514,N_17419,N_17400);
and U17515 (N_17515,N_17280,N_17441);
or U17516 (N_17516,N_17316,N_17308);
nand U17517 (N_17517,N_17344,N_17272);
nor U17518 (N_17518,N_17498,N_17382);
nor U17519 (N_17519,N_17323,N_17379);
nor U17520 (N_17520,N_17255,N_17477);
and U17521 (N_17521,N_17392,N_17472);
nor U17522 (N_17522,N_17281,N_17432);
xnor U17523 (N_17523,N_17417,N_17282);
or U17524 (N_17524,N_17436,N_17274);
nor U17525 (N_17525,N_17495,N_17414);
or U17526 (N_17526,N_17452,N_17412);
nor U17527 (N_17527,N_17277,N_17434);
nor U17528 (N_17528,N_17307,N_17343);
nor U17529 (N_17529,N_17461,N_17349);
xnor U17530 (N_17530,N_17331,N_17332);
nand U17531 (N_17531,N_17351,N_17363);
xor U17532 (N_17532,N_17499,N_17481);
xnor U17533 (N_17533,N_17480,N_17496);
or U17534 (N_17534,N_17294,N_17321);
nand U17535 (N_17535,N_17468,N_17401);
and U17536 (N_17536,N_17494,N_17445);
or U17537 (N_17537,N_17488,N_17447);
nand U17538 (N_17538,N_17389,N_17365);
or U17539 (N_17539,N_17448,N_17273);
and U17540 (N_17540,N_17303,N_17267);
nand U17541 (N_17541,N_17395,N_17446);
and U17542 (N_17542,N_17313,N_17487);
nor U17543 (N_17543,N_17275,N_17324);
nand U17544 (N_17544,N_17301,N_17466);
xor U17545 (N_17545,N_17300,N_17359);
and U17546 (N_17546,N_17264,N_17404);
xor U17547 (N_17547,N_17356,N_17254);
nand U17548 (N_17548,N_17362,N_17266);
nand U17549 (N_17549,N_17296,N_17398);
and U17550 (N_17550,N_17260,N_17352);
nor U17551 (N_17551,N_17475,N_17262);
or U17552 (N_17552,N_17263,N_17346);
xor U17553 (N_17553,N_17437,N_17416);
and U17554 (N_17554,N_17491,N_17338);
and U17555 (N_17555,N_17426,N_17345);
nand U17556 (N_17556,N_17459,N_17304);
and U17557 (N_17557,N_17408,N_17328);
nand U17558 (N_17558,N_17259,N_17413);
and U17559 (N_17559,N_17283,N_17369);
nand U17560 (N_17560,N_17339,N_17411);
nand U17561 (N_17561,N_17371,N_17479);
nor U17562 (N_17562,N_17478,N_17460);
xnor U17563 (N_17563,N_17427,N_17486);
and U17564 (N_17564,N_17415,N_17299);
nand U17565 (N_17565,N_17329,N_17409);
nor U17566 (N_17566,N_17422,N_17287);
and U17567 (N_17567,N_17435,N_17336);
nor U17568 (N_17568,N_17256,N_17315);
nand U17569 (N_17569,N_17333,N_17355);
nand U17570 (N_17570,N_17350,N_17317);
nor U17571 (N_17571,N_17407,N_17402);
nand U17572 (N_17572,N_17399,N_17364);
or U17573 (N_17573,N_17368,N_17453);
nor U17574 (N_17574,N_17467,N_17387);
or U17575 (N_17575,N_17386,N_17482);
nor U17576 (N_17576,N_17463,N_17335);
and U17577 (N_17577,N_17373,N_17360);
xnor U17578 (N_17578,N_17455,N_17429);
and U17579 (N_17579,N_17464,N_17289);
xor U17580 (N_17580,N_17391,N_17439);
or U17581 (N_17581,N_17377,N_17366);
nand U17582 (N_17582,N_17457,N_17276);
or U17583 (N_17583,N_17462,N_17476);
and U17584 (N_17584,N_17372,N_17306);
or U17585 (N_17585,N_17340,N_17293);
xor U17586 (N_17586,N_17497,N_17290);
nand U17587 (N_17587,N_17385,N_17381);
nor U17588 (N_17588,N_17490,N_17403);
or U17589 (N_17589,N_17291,N_17430);
nor U17590 (N_17590,N_17374,N_17285);
nor U17591 (N_17591,N_17442,N_17251);
nand U17592 (N_17592,N_17440,N_17341);
nand U17593 (N_17593,N_17493,N_17320);
or U17594 (N_17594,N_17347,N_17376);
nand U17595 (N_17595,N_17268,N_17357);
or U17596 (N_17596,N_17258,N_17438);
or U17597 (N_17597,N_17375,N_17394);
and U17598 (N_17598,N_17428,N_17367);
nand U17599 (N_17599,N_17330,N_17325);
or U17600 (N_17600,N_17342,N_17443);
nand U17601 (N_17601,N_17353,N_17390);
xor U17602 (N_17602,N_17314,N_17326);
xnor U17603 (N_17603,N_17334,N_17271);
nor U17604 (N_17604,N_17406,N_17278);
nor U17605 (N_17605,N_17319,N_17405);
and U17606 (N_17606,N_17483,N_17397);
and U17607 (N_17607,N_17425,N_17358);
nor U17608 (N_17608,N_17252,N_17431);
nor U17609 (N_17609,N_17474,N_17302);
xnor U17610 (N_17610,N_17348,N_17284);
nor U17611 (N_17611,N_17257,N_17418);
nand U17612 (N_17612,N_17451,N_17485);
or U17613 (N_17613,N_17449,N_17288);
nor U17614 (N_17614,N_17361,N_17311);
and U17615 (N_17615,N_17279,N_17484);
nand U17616 (N_17616,N_17310,N_17309);
nand U17617 (N_17617,N_17489,N_17337);
nor U17618 (N_17618,N_17297,N_17423);
xor U17619 (N_17619,N_17327,N_17312);
and U17620 (N_17620,N_17388,N_17261);
nand U17621 (N_17621,N_17322,N_17318);
xnor U17622 (N_17622,N_17298,N_17420);
xor U17623 (N_17623,N_17433,N_17380);
nor U17624 (N_17624,N_17270,N_17410);
or U17625 (N_17625,N_17308,N_17492);
nand U17626 (N_17626,N_17366,N_17419);
and U17627 (N_17627,N_17493,N_17436);
and U17628 (N_17628,N_17316,N_17453);
nand U17629 (N_17629,N_17269,N_17393);
nor U17630 (N_17630,N_17334,N_17456);
and U17631 (N_17631,N_17443,N_17253);
or U17632 (N_17632,N_17453,N_17372);
xor U17633 (N_17633,N_17472,N_17276);
xor U17634 (N_17634,N_17427,N_17293);
xnor U17635 (N_17635,N_17498,N_17385);
nor U17636 (N_17636,N_17497,N_17282);
or U17637 (N_17637,N_17342,N_17338);
nor U17638 (N_17638,N_17341,N_17427);
nand U17639 (N_17639,N_17345,N_17288);
nand U17640 (N_17640,N_17413,N_17455);
xor U17641 (N_17641,N_17325,N_17495);
and U17642 (N_17642,N_17312,N_17398);
nor U17643 (N_17643,N_17256,N_17486);
xor U17644 (N_17644,N_17354,N_17347);
xnor U17645 (N_17645,N_17278,N_17340);
nor U17646 (N_17646,N_17290,N_17263);
or U17647 (N_17647,N_17452,N_17363);
xor U17648 (N_17648,N_17401,N_17322);
nand U17649 (N_17649,N_17485,N_17359);
nand U17650 (N_17650,N_17407,N_17317);
and U17651 (N_17651,N_17452,N_17364);
nor U17652 (N_17652,N_17258,N_17415);
nand U17653 (N_17653,N_17364,N_17421);
nand U17654 (N_17654,N_17334,N_17402);
or U17655 (N_17655,N_17400,N_17366);
xnor U17656 (N_17656,N_17389,N_17256);
nor U17657 (N_17657,N_17468,N_17476);
or U17658 (N_17658,N_17304,N_17254);
nor U17659 (N_17659,N_17319,N_17410);
nor U17660 (N_17660,N_17407,N_17281);
xnor U17661 (N_17661,N_17426,N_17251);
nand U17662 (N_17662,N_17255,N_17376);
xor U17663 (N_17663,N_17306,N_17309);
nor U17664 (N_17664,N_17398,N_17453);
nor U17665 (N_17665,N_17463,N_17254);
xnor U17666 (N_17666,N_17400,N_17271);
and U17667 (N_17667,N_17467,N_17357);
nand U17668 (N_17668,N_17373,N_17344);
nor U17669 (N_17669,N_17416,N_17402);
or U17670 (N_17670,N_17493,N_17447);
and U17671 (N_17671,N_17269,N_17288);
or U17672 (N_17672,N_17427,N_17394);
nor U17673 (N_17673,N_17281,N_17318);
nand U17674 (N_17674,N_17361,N_17320);
xor U17675 (N_17675,N_17411,N_17427);
and U17676 (N_17676,N_17351,N_17308);
xor U17677 (N_17677,N_17435,N_17342);
nor U17678 (N_17678,N_17445,N_17396);
xor U17679 (N_17679,N_17478,N_17273);
and U17680 (N_17680,N_17492,N_17285);
and U17681 (N_17681,N_17474,N_17301);
nand U17682 (N_17682,N_17315,N_17355);
and U17683 (N_17683,N_17352,N_17274);
or U17684 (N_17684,N_17448,N_17400);
and U17685 (N_17685,N_17467,N_17457);
and U17686 (N_17686,N_17400,N_17287);
nand U17687 (N_17687,N_17341,N_17255);
or U17688 (N_17688,N_17426,N_17454);
nor U17689 (N_17689,N_17326,N_17373);
and U17690 (N_17690,N_17274,N_17485);
nor U17691 (N_17691,N_17328,N_17472);
nand U17692 (N_17692,N_17379,N_17387);
nor U17693 (N_17693,N_17260,N_17358);
nand U17694 (N_17694,N_17254,N_17370);
and U17695 (N_17695,N_17335,N_17468);
or U17696 (N_17696,N_17387,N_17275);
or U17697 (N_17697,N_17385,N_17343);
nand U17698 (N_17698,N_17432,N_17472);
and U17699 (N_17699,N_17489,N_17446);
xnor U17700 (N_17700,N_17332,N_17456);
nor U17701 (N_17701,N_17478,N_17268);
nand U17702 (N_17702,N_17267,N_17409);
and U17703 (N_17703,N_17428,N_17304);
nand U17704 (N_17704,N_17416,N_17275);
xnor U17705 (N_17705,N_17494,N_17357);
nand U17706 (N_17706,N_17359,N_17419);
nor U17707 (N_17707,N_17464,N_17250);
nand U17708 (N_17708,N_17476,N_17491);
and U17709 (N_17709,N_17426,N_17276);
xnor U17710 (N_17710,N_17490,N_17330);
xnor U17711 (N_17711,N_17331,N_17388);
or U17712 (N_17712,N_17309,N_17491);
nand U17713 (N_17713,N_17320,N_17461);
or U17714 (N_17714,N_17259,N_17400);
nor U17715 (N_17715,N_17467,N_17393);
and U17716 (N_17716,N_17465,N_17452);
and U17717 (N_17717,N_17257,N_17319);
nor U17718 (N_17718,N_17303,N_17310);
or U17719 (N_17719,N_17482,N_17450);
or U17720 (N_17720,N_17297,N_17411);
and U17721 (N_17721,N_17355,N_17496);
nor U17722 (N_17722,N_17477,N_17389);
or U17723 (N_17723,N_17451,N_17499);
xnor U17724 (N_17724,N_17271,N_17401);
xor U17725 (N_17725,N_17496,N_17294);
xnor U17726 (N_17726,N_17261,N_17366);
or U17727 (N_17727,N_17441,N_17322);
and U17728 (N_17728,N_17494,N_17465);
xor U17729 (N_17729,N_17290,N_17430);
xnor U17730 (N_17730,N_17416,N_17397);
and U17731 (N_17731,N_17411,N_17274);
nor U17732 (N_17732,N_17448,N_17362);
or U17733 (N_17733,N_17441,N_17298);
and U17734 (N_17734,N_17310,N_17271);
and U17735 (N_17735,N_17464,N_17304);
xnor U17736 (N_17736,N_17264,N_17316);
or U17737 (N_17737,N_17267,N_17444);
nor U17738 (N_17738,N_17495,N_17487);
and U17739 (N_17739,N_17470,N_17486);
nand U17740 (N_17740,N_17366,N_17397);
xnor U17741 (N_17741,N_17480,N_17400);
and U17742 (N_17742,N_17347,N_17455);
or U17743 (N_17743,N_17414,N_17487);
xnor U17744 (N_17744,N_17375,N_17425);
xnor U17745 (N_17745,N_17424,N_17434);
nor U17746 (N_17746,N_17409,N_17320);
nor U17747 (N_17747,N_17367,N_17475);
xor U17748 (N_17748,N_17353,N_17405);
nor U17749 (N_17749,N_17360,N_17418);
xor U17750 (N_17750,N_17620,N_17614);
and U17751 (N_17751,N_17519,N_17668);
nand U17752 (N_17752,N_17683,N_17549);
nand U17753 (N_17753,N_17730,N_17587);
or U17754 (N_17754,N_17676,N_17702);
or U17755 (N_17755,N_17563,N_17667);
xnor U17756 (N_17756,N_17705,N_17719);
nand U17757 (N_17757,N_17707,N_17593);
nand U17758 (N_17758,N_17728,N_17746);
nor U17759 (N_17759,N_17712,N_17565);
and U17760 (N_17760,N_17529,N_17694);
and U17761 (N_17761,N_17557,N_17555);
and U17762 (N_17762,N_17535,N_17713);
or U17763 (N_17763,N_17742,N_17546);
and U17764 (N_17764,N_17633,N_17560);
xor U17765 (N_17765,N_17640,N_17604);
nor U17766 (N_17766,N_17580,N_17714);
or U17767 (N_17767,N_17570,N_17630);
nor U17768 (N_17768,N_17654,N_17637);
nor U17769 (N_17769,N_17509,N_17603);
or U17770 (N_17770,N_17720,N_17748);
and U17771 (N_17771,N_17679,N_17513);
or U17772 (N_17772,N_17581,N_17692);
and U17773 (N_17773,N_17652,N_17599);
or U17774 (N_17774,N_17698,N_17624);
and U17775 (N_17775,N_17503,N_17611);
nor U17776 (N_17776,N_17569,N_17735);
or U17777 (N_17777,N_17699,N_17558);
xnor U17778 (N_17778,N_17635,N_17533);
nand U17779 (N_17779,N_17512,N_17553);
xor U17780 (N_17780,N_17726,N_17677);
or U17781 (N_17781,N_17596,N_17650);
and U17782 (N_17782,N_17615,N_17592);
nor U17783 (N_17783,N_17693,N_17623);
or U17784 (N_17784,N_17724,N_17554);
nand U17785 (N_17785,N_17551,N_17669);
and U17786 (N_17786,N_17566,N_17528);
or U17787 (N_17787,N_17643,N_17734);
or U17788 (N_17788,N_17638,N_17515);
or U17789 (N_17789,N_17722,N_17556);
nor U17790 (N_17790,N_17506,N_17542);
xor U17791 (N_17791,N_17612,N_17656);
or U17792 (N_17792,N_17745,N_17664);
and U17793 (N_17793,N_17514,N_17576);
nor U17794 (N_17794,N_17508,N_17625);
nor U17795 (N_17795,N_17736,N_17718);
and U17796 (N_17796,N_17696,N_17744);
nor U17797 (N_17797,N_17559,N_17572);
and U17798 (N_17798,N_17544,N_17573);
or U17799 (N_17799,N_17579,N_17715);
and U17800 (N_17800,N_17629,N_17657);
nand U17801 (N_17801,N_17740,N_17627);
xnor U17802 (N_17802,N_17685,N_17541);
nand U17803 (N_17803,N_17649,N_17500);
nand U17804 (N_17804,N_17723,N_17590);
nor U17805 (N_17805,N_17504,N_17710);
and U17806 (N_17806,N_17716,N_17527);
xnor U17807 (N_17807,N_17648,N_17636);
or U17808 (N_17808,N_17682,N_17700);
nor U17809 (N_17809,N_17586,N_17507);
nand U17810 (N_17810,N_17647,N_17601);
xor U17811 (N_17811,N_17727,N_17626);
nor U17812 (N_17812,N_17536,N_17532);
or U17813 (N_17813,N_17521,N_17721);
and U17814 (N_17814,N_17680,N_17518);
and U17815 (N_17815,N_17608,N_17659);
xor U17816 (N_17816,N_17562,N_17591);
and U17817 (N_17817,N_17645,N_17741);
nor U17818 (N_17818,N_17660,N_17609);
nor U17819 (N_17819,N_17522,N_17709);
nor U17820 (N_17820,N_17725,N_17689);
nand U17821 (N_17821,N_17749,N_17585);
nor U17822 (N_17822,N_17545,N_17665);
and U17823 (N_17823,N_17670,N_17589);
nor U17824 (N_17824,N_17524,N_17594);
or U17825 (N_17825,N_17731,N_17534);
or U17826 (N_17826,N_17733,N_17617);
or U17827 (N_17827,N_17540,N_17738);
or U17828 (N_17828,N_17543,N_17703);
nor U17829 (N_17829,N_17684,N_17711);
or U17830 (N_17830,N_17662,N_17675);
xor U17831 (N_17831,N_17516,N_17550);
and U17832 (N_17832,N_17678,N_17653);
and U17833 (N_17833,N_17747,N_17538);
and U17834 (N_17834,N_17697,N_17732);
xor U17835 (N_17835,N_17578,N_17681);
xor U17836 (N_17836,N_17686,N_17666);
and U17837 (N_17837,N_17517,N_17598);
or U17838 (N_17838,N_17690,N_17523);
nor U17839 (N_17839,N_17704,N_17505);
nor U17840 (N_17840,N_17717,N_17634);
nor U17841 (N_17841,N_17618,N_17671);
xnor U17842 (N_17842,N_17537,N_17530);
and U17843 (N_17843,N_17701,N_17520);
or U17844 (N_17844,N_17691,N_17502);
nand U17845 (N_17845,N_17687,N_17561);
and U17846 (N_17846,N_17641,N_17577);
and U17847 (N_17847,N_17632,N_17607);
or U17848 (N_17848,N_17695,N_17597);
nand U17849 (N_17849,N_17595,N_17673);
nor U17850 (N_17850,N_17511,N_17525);
and U17851 (N_17851,N_17574,N_17583);
and U17852 (N_17852,N_17552,N_17743);
xor U17853 (N_17853,N_17688,N_17622);
nor U17854 (N_17854,N_17588,N_17606);
xor U17855 (N_17855,N_17661,N_17584);
or U17856 (N_17856,N_17658,N_17628);
xor U17857 (N_17857,N_17605,N_17616);
or U17858 (N_17858,N_17600,N_17674);
xor U17859 (N_17859,N_17663,N_17610);
nand U17860 (N_17860,N_17655,N_17501);
nand U17861 (N_17861,N_17526,N_17729);
or U17862 (N_17862,N_17646,N_17737);
or U17863 (N_17863,N_17539,N_17639);
nor U17864 (N_17864,N_17708,N_17621);
nand U17865 (N_17865,N_17510,N_17531);
nand U17866 (N_17866,N_17571,N_17547);
and U17867 (N_17867,N_17739,N_17619);
or U17868 (N_17868,N_17567,N_17582);
and U17869 (N_17869,N_17548,N_17672);
nand U17870 (N_17870,N_17706,N_17575);
or U17871 (N_17871,N_17631,N_17568);
or U17872 (N_17872,N_17644,N_17613);
xor U17873 (N_17873,N_17642,N_17651);
and U17874 (N_17874,N_17564,N_17602);
xor U17875 (N_17875,N_17520,N_17721);
and U17876 (N_17876,N_17518,N_17674);
nor U17877 (N_17877,N_17648,N_17538);
or U17878 (N_17878,N_17674,N_17731);
nor U17879 (N_17879,N_17648,N_17738);
xor U17880 (N_17880,N_17626,N_17514);
or U17881 (N_17881,N_17721,N_17611);
nand U17882 (N_17882,N_17566,N_17641);
xor U17883 (N_17883,N_17513,N_17515);
nor U17884 (N_17884,N_17672,N_17730);
xor U17885 (N_17885,N_17697,N_17639);
nor U17886 (N_17886,N_17532,N_17666);
or U17887 (N_17887,N_17587,N_17600);
and U17888 (N_17888,N_17590,N_17530);
and U17889 (N_17889,N_17604,N_17526);
xnor U17890 (N_17890,N_17726,N_17685);
xnor U17891 (N_17891,N_17564,N_17574);
nand U17892 (N_17892,N_17549,N_17657);
nor U17893 (N_17893,N_17735,N_17561);
or U17894 (N_17894,N_17595,N_17672);
and U17895 (N_17895,N_17657,N_17531);
nor U17896 (N_17896,N_17615,N_17600);
nor U17897 (N_17897,N_17670,N_17569);
nand U17898 (N_17898,N_17643,N_17581);
nor U17899 (N_17899,N_17596,N_17610);
nor U17900 (N_17900,N_17623,N_17604);
nand U17901 (N_17901,N_17556,N_17516);
xnor U17902 (N_17902,N_17629,N_17691);
nor U17903 (N_17903,N_17730,N_17516);
nand U17904 (N_17904,N_17728,N_17656);
or U17905 (N_17905,N_17665,N_17671);
xnor U17906 (N_17906,N_17569,N_17697);
nand U17907 (N_17907,N_17626,N_17647);
or U17908 (N_17908,N_17654,N_17513);
nand U17909 (N_17909,N_17567,N_17649);
nand U17910 (N_17910,N_17565,N_17589);
xnor U17911 (N_17911,N_17603,N_17540);
and U17912 (N_17912,N_17665,N_17566);
nand U17913 (N_17913,N_17608,N_17741);
nor U17914 (N_17914,N_17562,N_17523);
nand U17915 (N_17915,N_17709,N_17513);
and U17916 (N_17916,N_17526,N_17732);
and U17917 (N_17917,N_17662,N_17734);
and U17918 (N_17918,N_17740,N_17648);
and U17919 (N_17919,N_17605,N_17563);
xor U17920 (N_17920,N_17501,N_17709);
and U17921 (N_17921,N_17508,N_17532);
or U17922 (N_17922,N_17521,N_17511);
xnor U17923 (N_17923,N_17634,N_17609);
xnor U17924 (N_17924,N_17578,N_17722);
nand U17925 (N_17925,N_17590,N_17686);
or U17926 (N_17926,N_17651,N_17538);
or U17927 (N_17927,N_17671,N_17666);
nand U17928 (N_17928,N_17506,N_17508);
nor U17929 (N_17929,N_17532,N_17590);
or U17930 (N_17930,N_17685,N_17552);
and U17931 (N_17931,N_17609,N_17683);
and U17932 (N_17932,N_17513,N_17564);
nand U17933 (N_17933,N_17747,N_17604);
nor U17934 (N_17934,N_17531,N_17616);
and U17935 (N_17935,N_17611,N_17725);
or U17936 (N_17936,N_17709,N_17740);
nand U17937 (N_17937,N_17633,N_17550);
and U17938 (N_17938,N_17737,N_17594);
xor U17939 (N_17939,N_17533,N_17577);
or U17940 (N_17940,N_17588,N_17501);
and U17941 (N_17941,N_17578,N_17536);
nand U17942 (N_17942,N_17708,N_17589);
or U17943 (N_17943,N_17523,N_17598);
nor U17944 (N_17944,N_17663,N_17500);
nor U17945 (N_17945,N_17609,N_17547);
xnor U17946 (N_17946,N_17725,N_17547);
nand U17947 (N_17947,N_17615,N_17695);
xnor U17948 (N_17948,N_17530,N_17500);
xnor U17949 (N_17949,N_17714,N_17541);
or U17950 (N_17950,N_17573,N_17686);
or U17951 (N_17951,N_17677,N_17585);
nand U17952 (N_17952,N_17650,N_17739);
and U17953 (N_17953,N_17745,N_17669);
nand U17954 (N_17954,N_17731,N_17690);
nor U17955 (N_17955,N_17587,N_17689);
nand U17956 (N_17956,N_17657,N_17512);
and U17957 (N_17957,N_17580,N_17719);
nor U17958 (N_17958,N_17512,N_17695);
xor U17959 (N_17959,N_17554,N_17618);
xor U17960 (N_17960,N_17671,N_17663);
and U17961 (N_17961,N_17746,N_17736);
nor U17962 (N_17962,N_17551,N_17737);
xor U17963 (N_17963,N_17688,N_17643);
xor U17964 (N_17964,N_17574,N_17719);
nor U17965 (N_17965,N_17539,N_17633);
and U17966 (N_17966,N_17649,N_17515);
nand U17967 (N_17967,N_17537,N_17508);
and U17968 (N_17968,N_17533,N_17529);
or U17969 (N_17969,N_17579,N_17512);
xor U17970 (N_17970,N_17555,N_17655);
xnor U17971 (N_17971,N_17504,N_17523);
nand U17972 (N_17972,N_17700,N_17534);
and U17973 (N_17973,N_17650,N_17705);
or U17974 (N_17974,N_17655,N_17508);
or U17975 (N_17975,N_17649,N_17716);
or U17976 (N_17976,N_17615,N_17731);
nor U17977 (N_17977,N_17680,N_17719);
nand U17978 (N_17978,N_17733,N_17526);
nand U17979 (N_17979,N_17699,N_17636);
and U17980 (N_17980,N_17603,N_17713);
and U17981 (N_17981,N_17610,N_17711);
nor U17982 (N_17982,N_17606,N_17597);
nand U17983 (N_17983,N_17592,N_17525);
or U17984 (N_17984,N_17593,N_17506);
nor U17985 (N_17985,N_17590,N_17556);
xnor U17986 (N_17986,N_17625,N_17587);
nand U17987 (N_17987,N_17608,N_17647);
nor U17988 (N_17988,N_17582,N_17664);
xor U17989 (N_17989,N_17536,N_17646);
or U17990 (N_17990,N_17558,N_17717);
nand U17991 (N_17991,N_17571,N_17624);
xor U17992 (N_17992,N_17613,N_17710);
or U17993 (N_17993,N_17612,N_17538);
xnor U17994 (N_17994,N_17744,N_17702);
and U17995 (N_17995,N_17655,N_17617);
xnor U17996 (N_17996,N_17602,N_17546);
xor U17997 (N_17997,N_17644,N_17670);
and U17998 (N_17998,N_17588,N_17703);
nor U17999 (N_17999,N_17636,N_17733);
nand U18000 (N_18000,N_17977,N_17901);
and U18001 (N_18001,N_17939,N_17862);
xor U18002 (N_18002,N_17954,N_17842);
or U18003 (N_18003,N_17777,N_17763);
and U18004 (N_18004,N_17983,N_17941);
nor U18005 (N_18005,N_17803,N_17887);
nand U18006 (N_18006,N_17867,N_17990);
and U18007 (N_18007,N_17973,N_17899);
and U18008 (N_18008,N_17856,N_17995);
and U18009 (N_18009,N_17795,N_17761);
and U18010 (N_18010,N_17970,N_17979);
xnor U18011 (N_18011,N_17923,N_17894);
or U18012 (N_18012,N_17787,N_17888);
xnor U18013 (N_18013,N_17846,N_17804);
nor U18014 (N_18014,N_17785,N_17934);
or U18015 (N_18015,N_17929,N_17854);
xnor U18016 (N_18016,N_17840,N_17988);
or U18017 (N_18017,N_17764,N_17776);
or U18018 (N_18018,N_17869,N_17806);
xor U18019 (N_18019,N_17930,N_17823);
nand U18020 (N_18020,N_17808,N_17768);
nand U18021 (N_18021,N_17865,N_17841);
nand U18022 (N_18022,N_17965,N_17826);
xor U18023 (N_18023,N_17922,N_17896);
and U18024 (N_18024,N_17851,N_17817);
nor U18025 (N_18025,N_17998,N_17883);
xnor U18026 (N_18026,N_17871,N_17953);
nand U18027 (N_18027,N_17760,N_17882);
xnor U18028 (N_18028,N_17945,N_17868);
or U18029 (N_18029,N_17982,N_17994);
or U18030 (N_18030,N_17984,N_17928);
xor U18031 (N_18031,N_17890,N_17786);
nor U18032 (N_18032,N_17799,N_17821);
nor U18033 (N_18033,N_17835,N_17946);
nor U18034 (N_18034,N_17989,N_17766);
nand U18035 (N_18035,N_17809,N_17937);
and U18036 (N_18036,N_17900,N_17770);
xnor U18037 (N_18037,N_17872,N_17828);
xor U18038 (N_18038,N_17911,N_17791);
xor U18039 (N_18039,N_17903,N_17978);
and U18040 (N_18040,N_17825,N_17950);
nand U18041 (N_18041,N_17788,N_17794);
nand U18042 (N_18042,N_17811,N_17783);
xor U18043 (N_18043,N_17962,N_17792);
and U18044 (N_18044,N_17782,N_17836);
nor U18045 (N_18045,N_17762,N_17975);
and U18046 (N_18046,N_17885,N_17765);
or U18047 (N_18047,N_17798,N_17891);
nand U18048 (N_18048,N_17845,N_17963);
or U18049 (N_18049,N_17848,N_17834);
xor U18050 (N_18050,N_17912,N_17844);
xor U18051 (N_18051,N_17832,N_17754);
and U18052 (N_18052,N_17820,N_17933);
xnor U18053 (N_18053,N_17905,N_17801);
or U18054 (N_18054,N_17897,N_17926);
and U18055 (N_18055,N_17757,N_17910);
or U18056 (N_18056,N_17952,N_17898);
xor U18057 (N_18057,N_17864,N_17827);
and U18058 (N_18058,N_17987,N_17857);
and U18059 (N_18059,N_17949,N_17895);
nor U18060 (N_18060,N_17824,N_17815);
or U18061 (N_18061,N_17847,N_17784);
xnor U18062 (N_18062,N_17751,N_17893);
nand U18063 (N_18063,N_17920,N_17956);
and U18064 (N_18064,N_17948,N_17800);
nor U18065 (N_18065,N_17813,N_17843);
xnor U18066 (N_18066,N_17860,N_17951);
nor U18067 (N_18067,N_17886,N_17914);
nor U18068 (N_18068,N_17859,N_17902);
xnor U18069 (N_18069,N_17810,N_17773);
and U18070 (N_18070,N_17924,N_17992);
or U18071 (N_18071,N_17942,N_17972);
or U18072 (N_18072,N_17879,N_17974);
nor U18073 (N_18073,N_17779,N_17781);
nand U18074 (N_18074,N_17932,N_17793);
nor U18075 (N_18075,N_17822,N_17993);
or U18076 (N_18076,N_17818,N_17907);
nor U18077 (N_18077,N_17919,N_17837);
nor U18078 (N_18078,N_17797,N_17904);
xor U18079 (N_18079,N_17936,N_17796);
xnor U18080 (N_18080,N_17812,N_17816);
nor U18081 (N_18081,N_17753,N_17935);
and U18082 (N_18082,N_17940,N_17976);
nor U18083 (N_18083,N_17927,N_17913);
or U18084 (N_18084,N_17971,N_17789);
and U18085 (N_18085,N_17985,N_17968);
nor U18086 (N_18086,N_17780,N_17833);
nand U18087 (N_18087,N_17986,N_17839);
nor U18088 (N_18088,N_17866,N_17829);
xnor U18089 (N_18089,N_17955,N_17991);
or U18090 (N_18090,N_17997,N_17755);
and U18091 (N_18091,N_17878,N_17858);
and U18092 (N_18092,N_17908,N_17831);
or U18093 (N_18093,N_17850,N_17855);
nand U18094 (N_18094,N_17756,N_17915);
nand U18095 (N_18095,N_17964,N_17774);
nor U18096 (N_18096,N_17958,N_17759);
nor U18097 (N_18097,N_17790,N_17875);
nor U18098 (N_18098,N_17769,N_17959);
and U18099 (N_18099,N_17961,N_17876);
and U18100 (N_18100,N_17778,N_17931);
nand U18101 (N_18101,N_17758,N_17830);
nand U18102 (N_18102,N_17767,N_17916);
or U18103 (N_18103,N_17750,N_17999);
nand U18104 (N_18104,N_17892,N_17957);
nand U18105 (N_18105,N_17960,N_17925);
and U18106 (N_18106,N_17863,N_17881);
and U18107 (N_18107,N_17772,N_17861);
nand U18108 (N_18108,N_17967,N_17807);
or U18109 (N_18109,N_17996,N_17943);
nor U18110 (N_18110,N_17814,N_17771);
xnor U18111 (N_18111,N_17873,N_17938);
and U18112 (N_18112,N_17838,N_17918);
or U18113 (N_18113,N_17880,N_17947);
nand U18114 (N_18114,N_17802,N_17980);
nand U18115 (N_18115,N_17853,N_17981);
and U18116 (N_18116,N_17921,N_17909);
and U18117 (N_18117,N_17805,N_17849);
nand U18118 (N_18118,N_17966,N_17917);
and U18119 (N_18119,N_17944,N_17852);
nor U18120 (N_18120,N_17870,N_17906);
or U18121 (N_18121,N_17874,N_17752);
nor U18122 (N_18122,N_17819,N_17884);
xor U18123 (N_18123,N_17877,N_17889);
xnor U18124 (N_18124,N_17969,N_17775);
or U18125 (N_18125,N_17947,N_17850);
nor U18126 (N_18126,N_17986,N_17954);
xnor U18127 (N_18127,N_17879,N_17859);
xnor U18128 (N_18128,N_17750,N_17954);
or U18129 (N_18129,N_17763,N_17962);
nand U18130 (N_18130,N_17796,N_17807);
xnor U18131 (N_18131,N_17768,N_17962);
or U18132 (N_18132,N_17923,N_17762);
xnor U18133 (N_18133,N_17765,N_17783);
nand U18134 (N_18134,N_17880,N_17827);
or U18135 (N_18135,N_17869,N_17886);
and U18136 (N_18136,N_17954,N_17977);
or U18137 (N_18137,N_17779,N_17875);
nor U18138 (N_18138,N_17754,N_17931);
nand U18139 (N_18139,N_17821,N_17823);
xnor U18140 (N_18140,N_17812,N_17903);
and U18141 (N_18141,N_17814,N_17844);
or U18142 (N_18142,N_17862,N_17881);
nand U18143 (N_18143,N_17800,N_17861);
nor U18144 (N_18144,N_17956,N_17963);
or U18145 (N_18145,N_17784,N_17991);
or U18146 (N_18146,N_17788,N_17816);
nand U18147 (N_18147,N_17910,N_17960);
and U18148 (N_18148,N_17928,N_17956);
nand U18149 (N_18149,N_17888,N_17858);
nand U18150 (N_18150,N_17765,N_17899);
nor U18151 (N_18151,N_17854,N_17792);
nand U18152 (N_18152,N_17811,N_17779);
or U18153 (N_18153,N_17761,N_17833);
nand U18154 (N_18154,N_17777,N_17789);
nor U18155 (N_18155,N_17925,N_17853);
and U18156 (N_18156,N_17890,N_17881);
nand U18157 (N_18157,N_17958,N_17919);
and U18158 (N_18158,N_17952,N_17891);
and U18159 (N_18159,N_17989,N_17871);
nor U18160 (N_18160,N_17881,N_17891);
nor U18161 (N_18161,N_17938,N_17976);
nand U18162 (N_18162,N_17907,N_17755);
and U18163 (N_18163,N_17881,N_17889);
or U18164 (N_18164,N_17879,N_17804);
nand U18165 (N_18165,N_17825,N_17848);
and U18166 (N_18166,N_17777,N_17802);
or U18167 (N_18167,N_17799,N_17985);
nor U18168 (N_18168,N_17933,N_17864);
or U18169 (N_18169,N_17932,N_17938);
xnor U18170 (N_18170,N_17992,N_17840);
nor U18171 (N_18171,N_17977,N_17944);
nand U18172 (N_18172,N_17812,N_17947);
nand U18173 (N_18173,N_17858,N_17861);
nand U18174 (N_18174,N_17993,N_17909);
xnor U18175 (N_18175,N_17759,N_17878);
xor U18176 (N_18176,N_17930,N_17765);
xnor U18177 (N_18177,N_17988,N_17972);
nor U18178 (N_18178,N_17805,N_17942);
xnor U18179 (N_18179,N_17868,N_17859);
nor U18180 (N_18180,N_17941,N_17915);
xnor U18181 (N_18181,N_17921,N_17757);
or U18182 (N_18182,N_17881,N_17783);
and U18183 (N_18183,N_17974,N_17918);
nor U18184 (N_18184,N_17827,N_17823);
or U18185 (N_18185,N_17967,N_17896);
and U18186 (N_18186,N_17873,N_17843);
and U18187 (N_18187,N_17830,N_17909);
or U18188 (N_18188,N_17862,N_17765);
nor U18189 (N_18189,N_17994,N_17995);
nor U18190 (N_18190,N_17960,N_17767);
nor U18191 (N_18191,N_17913,N_17903);
and U18192 (N_18192,N_17860,N_17807);
xor U18193 (N_18193,N_17820,N_17936);
and U18194 (N_18194,N_17797,N_17944);
nor U18195 (N_18195,N_17857,N_17996);
xnor U18196 (N_18196,N_17947,N_17755);
xnor U18197 (N_18197,N_17930,N_17912);
nor U18198 (N_18198,N_17966,N_17804);
xor U18199 (N_18199,N_17766,N_17888);
or U18200 (N_18200,N_17854,N_17945);
nand U18201 (N_18201,N_17905,N_17939);
nor U18202 (N_18202,N_17870,N_17818);
xor U18203 (N_18203,N_17751,N_17968);
and U18204 (N_18204,N_17822,N_17996);
xnor U18205 (N_18205,N_17949,N_17921);
xor U18206 (N_18206,N_17968,N_17804);
and U18207 (N_18207,N_17988,N_17857);
and U18208 (N_18208,N_17999,N_17934);
and U18209 (N_18209,N_17976,N_17816);
nor U18210 (N_18210,N_17792,N_17832);
nor U18211 (N_18211,N_17871,N_17774);
nor U18212 (N_18212,N_17836,N_17780);
and U18213 (N_18213,N_17854,N_17788);
or U18214 (N_18214,N_17767,N_17974);
xor U18215 (N_18215,N_17786,N_17768);
or U18216 (N_18216,N_17887,N_17797);
xnor U18217 (N_18217,N_17755,N_17819);
and U18218 (N_18218,N_17826,N_17996);
or U18219 (N_18219,N_17886,N_17758);
xor U18220 (N_18220,N_17873,N_17937);
or U18221 (N_18221,N_17889,N_17948);
or U18222 (N_18222,N_17812,N_17918);
or U18223 (N_18223,N_17922,N_17994);
nor U18224 (N_18224,N_17864,N_17879);
nand U18225 (N_18225,N_17814,N_17858);
xnor U18226 (N_18226,N_17890,N_17759);
and U18227 (N_18227,N_17842,N_17767);
xor U18228 (N_18228,N_17993,N_17821);
nor U18229 (N_18229,N_17843,N_17875);
nor U18230 (N_18230,N_17886,N_17821);
nor U18231 (N_18231,N_17863,N_17756);
and U18232 (N_18232,N_17905,N_17984);
nand U18233 (N_18233,N_17974,N_17793);
nand U18234 (N_18234,N_17891,N_17899);
xor U18235 (N_18235,N_17939,N_17823);
nor U18236 (N_18236,N_17885,N_17767);
nand U18237 (N_18237,N_17823,N_17997);
and U18238 (N_18238,N_17810,N_17947);
nand U18239 (N_18239,N_17953,N_17979);
nor U18240 (N_18240,N_17948,N_17835);
nor U18241 (N_18241,N_17977,N_17873);
nor U18242 (N_18242,N_17825,N_17904);
xnor U18243 (N_18243,N_17842,N_17804);
xor U18244 (N_18244,N_17925,N_17901);
nor U18245 (N_18245,N_17971,N_17990);
or U18246 (N_18246,N_17825,N_17869);
xor U18247 (N_18247,N_17910,N_17859);
or U18248 (N_18248,N_17864,N_17819);
or U18249 (N_18249,N_17956,N_17812);
xor U18250 (N_18250,N_18096,N_18089);
xnor U18251 (N_18251,N_18194,N_18233);
xor U18252 (N_18252,N_18205,N_18164);
and U18253 (N_18253,N_18245,N_18163);
xnor U18254 (N_18254,N_18017,N_18062);
nand U18255 (N_18255,N_18003,N_18171);
and U18256 (N_18256,N_18015,N_18151);
xor U18257 (N_18257,N_18204,N_18021);
nand U18258 (N_18258,N_18074,N_18182);
xor U18259 (N_18259,N_18020,N_18119);
and U18260 (N_18260,N_18192,N_18046);
xor U18261 (N_18261,N_18161,N_18183);
nand U18262 (N_18262,N_18061,N_18219);
or U18263 (N_18263,N_18208,N_18110);
nand U18264 (N_18264,N_18092,N_18044);
nor U18265 (N_18265,N_18107,N_18083);
xor U18266 (N_18266,N_18090,N_18075);
xor U18267 (N_18267,N_18162,N_18141);
xnor U18268 (N_18268,N_18035,N_18060);
or U18269 (N_18269,N_18034,N_18196);
or U18270 (N_18270,N_18180,N_18124);
xor U18271 (N_18271,N_18023,N_18167);
nor U18272 (N_18272,N_18033,N_18159);
xor U18273 (N_18273,N_18117,N_18127);
nand U18274 (N_18274,N_18169,N_18104);
nor U18275 (N_18275,N_18174,N_18047);
or U18276 (N_18276,N_18160,N_18239);
nand U18277 (N_18277,N_18009,N_18248);
and U18278 (N_18278,N_18108,N_18246);
and U18279 (N_18279,N_18229,N_18105);
or U18280 (N_18280,N_18059,N_18038);
xor U18281 (N_18281,N_18008,N_18101);
xnor U18282 (N_18282,N_18150,N_18066);
or U18283 (N_18283,N_18184,N_18113);
or U18284 (N_18284,N_18014,N_18050);
nor U18285 (N_18285,N_18069,N_18098);
nor U18286 (N_18286,N_18048,N_18027);
nand U18287 (N_18287,N_18200,N_18057);
nor U18288 (N_18288,N_18199,N_18129);
nand U18289 (N_18289,N_18157,N_18191);
and U18290 (N_18290,N_18138,N_18122);
xnor U18291 (N_18291,N_18018,N_18187);
or U18292 (N_18292,N_18095,N_18243);
and U18293 (N_18293,N_18242,N_18140);
nand U18294 (N_18294,N_18212,N_18185);
nand U18295 (N_18295,N_18002,N_18128);
xnor U18296 (N_18296,N_18210,N_18207);
xnor U18297 (N_18297,N_18081,N_18173);
nor U18298 (N_18298,N_18147,N_18211);
and U18299 (N_18299,N_18158,N_18247);
and U18300 (N_18300,N_18218,N_18225);
nand U18301 (N_18301,N_18143,N_18209);
and U18302 (N_18302,N_18244,N_18206);
or U18303 (N_18303,N_18001,N_18077);
nor U18304 (N_18304,N_18026,N_18178);
nor U18305 (N_18305,N_18176,N_18220);
nor U18306 (N_18306,N_18013,N_18030);
xnor U18307 (N_18307,N_18088,N_18112);
nor U18308 (N_18308,N_18045,N_18168);
nand U18309 (N_18309,N_18231,N_18053);
nand U18310 (N_18310,N_18146,N_18007);
and U18311 (N_18311,N_18041,N_18132);
or U18312 (N_18312,N_18067,N_18100);
nand U18313 (N_18313,N_18238,N_18118);
nand U18314 (N_18314,N_18072,N_18234);
nor U18315 (N_18315,N_18106,N_18135);
and U18316 (N_18316,N_18042,N_18097);
xnor U18317 (N_18317,N_18010,N_18224);
and U18318 (N_18318,N_18094,N_18006);
nand U18319 (N_18319,N_18198,N_18149);
nand U18320 (N_18320,N_18188,N_18070);
nand U18321 (N_18321,N_18079,N_18040);
or U18322 (N_18322,N_18121,N_18133);
nor U18323 (N_18323,N_18156,N_18103);
nand U18324 (N_18324,N_18093,N_18043);
or U18325 (N_18325,N_18226,N_18091);
or U18326 (N_18326,N_18123,N_18087);
xor U18327 (N_18327,N_18202,N_18189);
or U18328 (N_18328,N_18011,N_18148);
xor U18329 (N_18329,N_18181,N_18086);
and U18330 (N_18330,N_18214,N_18022);
or U18331 (N_18331,N_18137,N_18049);
xor U18332 (N_18332,N_18222,N_18058);
nand U18333 (N_18333,N_18249,N_18177);
nor U18334 (N_18334,N_18170,N_18029);
nor U18335 (N_18335,N_18068,N_18175);
and U18336 (N_18336,N_18223,N_18145);
nor U18337 (N_18337,N_18024,N_18134);
nand U18338 (N_18338,N_18165,N_18172);
nor U18339 (N_18339,N_18080,N_18203);
xor U18340 (N_18340,N_18102,N_18126);
nand U18341 (N_18341,N_18115,N_18000);
or U18342 (N_18342,N_18099,N_18028);
and U18343 (N_18343,N_18216,N_18085);
xor U18344 (N_18344,N_18213,N_18193);
nand U18345 (N_18345,N_18051,N_18144);
and U18346 (N_18346,N_18078,N_18195);
and U18347 (N_18347,N_18237,N_18082);
or U18348 (N_18348,N_18120,N_18032);
nor U18349 (N_18349,N_18139,N_18004);
nor U18350 (N_18350,N_18227,N_18215);
xor U18351 (N_18351,N_18240,N_18073);
nand U18352 (N_18352,N_18036,N_18190);
nand U18353 (N_18353,N_18063,N_18025);
nand U18354 (N_18354,N_18201,N_18056);
nor U18355 (N_18355,N_18019,N_18031);
xor U18356 (N_18356,N_18065,N_18241);
or U18357 (N_18357,N_18071,N_18114);
and U18358 (N_18358,N_18230,N_18186);
nor U18359 (N_18359,N_18084,N_18054);
or U18360 (N_18360,N_18037,N_18109);
xnor U18361 (N_18361,N_18005,N_18136);
xor U18362 (N_18362,N_18064,N_18197);
or U18363 (N_18363,N_18076,N_18235);
xor U18364 (N_18364,N_18221,N_18131);
and U18365 (N_18365,N_18142,N_18012);
or U18366 (N_18366,N_18052,N_18217);
or U18367 (N_18367,N_18179,N_18152);
or U18368 (N_18368,N_18116,N_18228);
or U18369 (N_18369,N_18125,N_18154);
and U18370 (N_18370,N_18111,N_18166);
and U18371 (N_18371,N_18153,N_18055);
xor U18372 (N_18372,N_18236,N_18130);
or U18373 (N_18373,N_18039,N_18016);
xor U18374 (N_18374,N_18155,N_18232);
or U18375 (N_18375,N_18132,N_18227);
nor U18376 (N_18376,N_18171,N_18002);
xnor U18377 (N_18377,N_18245,N_18146);
xor U18378 (N_18378,N_18092,N_18212);
xnor U18379 (N_18379,N_18038,N_18052);
and U18380 (N_18380,N_18170,N_18174);
or U18381 (N_18381,N_18237,N_18124);
nor U18382 (N_18382,N_18062,N_18229);
nor U18383 (N_18383,N_18158,N_18075);
or U18384 (N_18384,N_18080,N_18093);
xnor U18385 (N_18385,N_18078,N_18124);
and U18386 (N_18386,N_18127,N_18155);
xnor U18387 (N_18387,N_18235,N_18118);
and U18388 (N_18388,N_18224,N_18156);
nand U18389 (N_18389,N_18166,N_18058);
and U18390 (N_18390,N_18171,N_18102);
and U18391 (N_18391,N_18113,N_18016);
xor U18392 (N_18392,N_18000,N_18191);
nor U18393 (N_18393,N_18228,N_18192);
and U18394 (N_18394,N_18059,N_18032);
nand U18395 (N_18395,N_18073,N_18001);
nand U18396 (N_18396,N_18164,N_18146);
xnor U18397 (N_18397,N_18041,N_18073);
nand U18398 (N_18398,N_18098,N_18114);
xnor U18399 (N_18399,N_18094,N_18028);
nand U18400 (N_18400,N_18150,N_18249);
or U18401 (N_18401,N_18204,N_18048);
and U18402 (N_18402,N_18148,N_18222);
and U18403 (N_18403,N_18001,N_18112);
xnor U18404 (N_18404,N_18171,N_18099);
and U18405 (N_18405,N_18020,N_18107);
nand U18406 (N_18406,N_18070,N_18199);
or U18407 (N_18407,N_18241,N_18043);
xnor U18408 (N_18408,N_18128,N_18156);
xor U18409 (N_18409,N_18071,N_18198);
nor U18410 (N_18410,N_18032,N_18188);
or U18411 (N_18411,N_18109,N_18177);
and U18412 (N_18412,N_18092,N_18149);
nand U18413 (N_18413,N_18028,N_18242);
and U18414 (N_18414,N_18009,N_18189);
nor U18415 (N_18415,N_18196,N_18159);
or U18416 (N_18416,N_18067,N_18179);
and U18417 (N_18417,N_18172,N_18155);
xor U18418 (N_18418,N_18180,N_18044);
xnor U18419 (N_18419,N_18149,N_18246);
or U18420 (N_18420,N_18152,N_18006);
xor U18421 (N_18421,N_18010,N_18123);
and U18422 (N_18422,N_18200,N_18205);
or U18423 (N_18423,N_18082,N_18186);
and U18424 (N_18424,N_18101,N_18134);
nor U18425 (N_18425,N_18080,N_18189);
or U18426 (N_18426,N_18043,N_18039);
xor U18427 (N_18427,N_18098,N_18131);
nor U18428 (N_18428,N_18198,N_18010);
nand U18429 (N_18429,N_18121,N_18067);
nand U18430 (N_18430,N_18096,N_18100);
nor U18431 (N_18431,N_18162,N_18200);
nor U18432 (N_18432,N_18027,N_18228);
or U18433 (N_18433,N_18201,N_18215);
and U18434 (N_18434,N_18197,N_18234);
xor U18435 (N_18435,N_18025,N_18022);
nand U18436 (N_18436,N_18069,N_18058);
xnor U18437 (N_18437,N_18162,N_18089);
xnor U18438 (N_18438,N_18189,N_18213);
or U18439 (N_18439,N_18204,N_18027);
and U18440 (N_18440,N_18214,N_18079);
nor U18441 (N_18441,N_18098,N_18036);
or U18442 (N_18442,N_18234,N_18212);
and U18443 (N_18443,N_18154,N_18239);
nand U18444 (N_18444,N_18072,N_18220);
or U18445 (N_18445,N_18012,N_18023);
nor U18446 (N_18446,N_18159,N_18103);
and U18447 (N_18447,N_18216,N_18218);
or U18448 (N_18448,N_18033,N_18118);
nor U18449 (N_18449,N_18002,N_18100);
xnor U18450 (N_18450,N_18134,N_18178);
and U18451 (N_18451,N_18202,N_18039);
and U18452 (N_18452,N_18080,N_18102);
and U18453 (N_18453,N_18113,N_18195);
or U18454 (N_18454,N_18093,N_18003);
or U18455 (N_18455,N_18086,N_18179);
xor U18456 (N_18456,N_18202,N_18147);
nand U18457 (N_18457,N_18242,N_18019);
nor U18458 (N_18458,N_18210,N_18151);
and U18459 (N_18459,N_18152,N_18042);
nor U18460 (N_18460,N_18219,N_18222);
and U18461 (N_18461,N_18220,N_18154);
xor U18462 (N_18462,N_18002,N_18112);
nand U18463 (N_18463,N_18018,N_18179);
nand U18464 (N_18464,N_18046,N_18088);
nand U18465 (N_18465,N_18114,N_18047);
nand U18466 (N_18466,N_18118,N_18029);
nor U18467 (N_18467,N_18174,N_18084);
or U18468 (N_18468,N_18048,N_18091);
nor U18469 (N_18469,N_18167,N_18249);
xnor U18470 (N_18470,N_18018,N_18103);
and U18471 (N_18471,N_18078,N_18189);
or U18472 (N_18472,N_18101,N_18221);
and U18473 (N_18473,N_18092,N_18124);
and U18474 (N_18474,N_18094,N_18027);
nand U18475 (N_18475,N_18013,N_18038);
or U18476 (N_18476,N_18234,N_18188);
xnor U18477 (N_18477,N_18024,N_18099);
or U18478 (N_18478,N_18115,N_18066);
and U18479 (N_18479,N_18237,N_18222);
or U18480 (N_18480,N_18163,N_18009);
or U18481 (N_18481,N_18184,N_18004);
nor U18482 (N_18482,N_18038,N_18032);
and U18483 (N_18483,N_18227,N_18234);
nand U18484 (N_18484,N_18243,N_18166);
nor U18485 (N_18485,N_18184,N_18129);
or U18486 (N_18486,N_18058,N_18047);
nand U18487 (N_18487,N_18084,N_18075);
or U18488 (N_18488,N_18207,N_18149);
nor U18489 (N_18489,N_18039,N_18215);
or U18490 (N_18490,N_18177,N_18215);
or U18491 (N_18491,N_18162,N_18206);
xnor U18492 (N_18492,N_18172,N_18184);
xnor U18493 (N_18493,N_18130,N_18157);
nor U18494 (N_18494,N_18040,N_18074);
nor U18495 (N_18495,N_18021,N_18198);
and U18496 (N_18496,N_18187,N_18232);
or U18497 (N_18497,N_18146,N_18117);
or U18498 (N_18498,N_18227,N_18036);
or U18499 (N_18499,N_18199,N_18026);
nor U18500 (N_18500,N_18465,N_18354);
xnor U18501 (N_18501,N_18380,N_18370);
nand U18502 (N_18502,N_18363,N_18252);
and U18503 (N_18503,N_18272,N_18290);
nand U18504 (N_18504,N_18484,N_18427);
xnor U18505 (N_18505,N_18399,N_18491);
or U18506 (N_18506,N_18324,N_18446);
and U18507 (N_18507,N_18385,N_18358);
nor U18508 (N_18508,N_18326,N_18323);
nand U18509 (N_18509,N_18459,N_18360);
or U18510 (N_18510,N_18490,N_18454);
nor U18511 (N_18511,N_18453,N_18395);
nor U18512 (N_18512,N_18458,N_18288);
and U18513 (N_18513,N_18353,N_18477);
nor U18514 (N_18514,N_18280,N_18338);
nand U18515 (N_18515,N_18268,N_18476);
nor U18516 (N_18516,N_18406,N_18325);
and U18517 (N_18517,N_18388,N_18349);
and U18518 (N_18518,N_18452,N_18373);
nor U18519 (N_18519,N_18261,N_18377);
nand U18520 (N_18520,N_18258,N_18313);
or U18521 (N_18521,N_18265,N_18404);
or U18522 (N_18522,N_18493,N_18462);
nand U18523 (N_18523,N_18294,N_18348);
nand U18524 (N_18524,N_18309,N_18467);
nand U18525 (N_18525,N_18461,N_18424);
or U18526 (N_18526,N_18411,N_18456);
nand U18527 (N_18527,N_18293,N_18291);
or U18528 (N_18528,N_18441,N_18311);
nor U18529 (N_18529,N_18418,N_18438);
and U18530 (N_18530,N_18421,N_18410);
xnor U18531 (N_18531,N_18304,N_18301);
nand U18532 (N_18532,N_18285,N_18351);
and U18533 (N_18533,N_18402,N_18383);
xnor U18534 (N_18534,N_18425,N_18396);
or U18535 (N_18535,N_18480,N_18469);
or U18536 (N_18536,N_18356,N_18431);
or U18537 (N_18537,N_18332,N_18281);
or U18538 (N_18538,N_18361,N_18322);
nor U18539 (N_18539,N_18444,N_18440);
nor U18540 (N_18540,N_18328,N_18299);
or U18541 (N_18541,N_18282,N_18333);
or U18542 (N_18542,N_18352,N_18307);
or U18543 (N_18543,N_18319,N_18375);
xnor U18544 (N_18544,N_18340,N_18344);
nand U18545 (N_18545,N_18442,N_18369);
and U18546 (N_18546,N_18419,N_18310);
nand U18547 (N_18547,N_18479,N_18350);
nand U18548 (N_18548,N_18317,N_18487);
nor U18549 (N_18549,N_18355,N_18306);
or U18550 (N_18550,N_18345,N_18278);
and U18551 (N_18551,N_18368,N_18259);
nand U18552 (N_18552,N_18331,N_18390);
xor U18553 (N_18553,N_18297,N_18433);
xnor U18554 (N_18554,N_18412,N_18494);
xor U18555 (N_18555,N_18336,N_18423);
or U18556 (N_18556,N_18463,N_18339);
xor U18557 (N_18557,N_18498,N_18372);
or U18558 (N_18558,N_18273,N_18365);
and U18559 (N_18559,N_18284,N_18266);
or U18560 (N_18560,N_18475,N_18426);
nor U18561 (N_18561,N_18384,N_18405);
and U18562 (N_18562,N_18382,N_18409);
xor U18563 (N_18563,N_18447,N_18296);
nor U18564 (N_18564,N_18389,N_18393);
or U18565 (N_18565,N_18318,N_18286);
nor U18566 (N_18566,N_18416,N_18376);
nor U18567 (N_18567,N_18379,N_18267);
or U18568 (N_18568,N_18392,N_18422);
nand U18569 (N_18569,N_18414,N_18346);
or U18570 (N_18570,N_18295,N_18337);
and U18571 (N_18571,N_18437,N_18474);
nor U18572 (N_18572,N_18478,N_18359);
xor U18573 (N_18573,N_18366,N_18473);
xnor U18574 (N_18574,N_18492,N_18445);
nor U18575 (N_18575,N_18460,N_18443);
nor U18576 (N_18576,N_18253,N_18362);
xnor U18577 (N_18577,N_18401,N_18300);
nand U18578 (N_18578,N_18420,N_18435);
and U18579 (N_18579,N_18308,N_18457);
and U18580 (N_18580,N_18330,N_18378);
and U18581 (N_18581,N_18312,N_18429);
and U18582 (N_18582,N_18343,N_18298);
xnor U18583 (N_18583,N_18466,N_18496);
nor U18584 (N_18584,N_18450,N_18263);
or U18585 (N_18585,N_18341,N_18251);
nand U18586 (N_18586,N_18279,N_18274);
and U18587 (N_18587,N_18451,N_18449);
xnor U18588 (N_18588,N_18262,N_18386);
nor U18589 (N_18589,N_18314,N_18485);
and U18590 (N_18590,N_18256,N_18287);
nand U18591 (N_18591,N_18320,N_18470);
nor U18592 (N_18592,N_18391,N_18434);
xnor U18593 (N_18593,N_18250,N_18374);
xor U18594 (N_18594,N_18283,N_18483);
and U18595 (N_18595,N_18270,N_18257);
nand U18596 (N_18596,N_18381,N_18455);
nor U18597 (N_18597,N_18387,N_18471);
and U18598 (N_18598,N_18397,N_18400);
xnor U18599 (N_18599,N_18367,N_18347);
xnor U18600 (N_18600,N_18482,N_18486);
or U18601 (N_18601,N_18417,N_18436);
and U18602 (N_18602,N_18305,N_18254);
nand U18603 (N_18603,N_18335,N_18357);
xnor U18604 (N_18604,N_18321,N_18269);
and U18605 (N_18605,N_18275,N_18276);
and U18606 (N_18606,N_18413,N_18302);
nand U18607 (N_18607,N_18448,N_18497);
nor U18608 (N_18608,N_18472,N_18316);
xor U18609 (N_18609,N_18398,N_18481);
or U18610 (N_18610,N_18289,N_18403);
and U18611 (N_18611,N_18432,N_18495);
xor U18612 (N_18612,N_18264,N_18292);
or U18613 (N_18613,N_18439,N_18415);
xnor U18614 (N_18614,N_18303,N_18255);
nor U18615 (N_18615,N_18329,N_18371);
nor U18616 (N_18616,N_18277,N_18260);
or U18617 (N_18617,N_18394,N_18334);
xor U18618 (N_18618,N_18342,N_18364);
nor U18619 (N_18619,N_18499,N_18327);
and U18620 (N_18620,N_18489,N_18271);
nor U18621 (N_18621,N_18468,N_18430);
xor U18622 (N_18622,N_18464,N_18488);
nor U18623 (N_18623,N_18408,N_18407);
or U18624 (N_18624,N_18315,N_18428);
nand U18625 (N_18625,N_18496,N_18467);
nor U18626 (N_18626,N_18476,N_18265);
nand U18627 (N_18627,N_18361,N_18410);
nand U18628 (N_18628,N_18460,N_18476);
or U18629 (N_18629,N_18335,N_18468);
or U18630 (N_18630,N_18347,N_18457);
nand U18631 (N_18631,N_18458,N_18358);
nand U18632 (N_18632,N_18409,N_18492);
xnor U18633 (N_18633,N_18372,N_18445);
xor U18634 (N_18634,N_18281,N_18256);
nor U18635 (N_18635,N_18413,N_18451);
xor U18636 (N_18636,N_18435,N_18350);
nor U18637 (N_18637,N_18393,N_18361);
xor U18638 (N_18638,N_18440,N_18385);
or U18639 (N_18639,N_18269,N_18263);
nor U18640 (N_18640,N_18472,N_18382);
or U18641 (N_18641,N_18296,N_18433);
or U18642 (N_18642,N_18298,N_18456);
xnor U18643 (N_18643,N_18357,N_18415);
xor U18644 (N_18644,N_18265,N_18322);
or U18645 (N_18645,N_18465,N_18440);
or U18646 (N_18646,N_18337,N_18306);
and U18647 (N_18647,N_18361,N_18349);
and U18648 (N_18648,N_18339,N_18346);
nand U18649 (N_18649,N_18321,N_18405);
xor U18650 (N_18650,N_18323,N_18319);
xor U18651 (N_18651,N_18389,N_18309);
nor U18652 (N_18652,N_18418,N_18348);
xnor U18653 (N_18653,N_18304,N_18361);
and U18654 (N_18654,N_18431,N_18483);
or U18655 (N_18655,N_18468,N_18425);
nor U18656 (N_18656,N_18438,N_18393);
nand U18657 (N_18657,N_18283,N_18409);
nand U18658 (N_18658,N_18267,N_18432);
and U18659 (N_18659,N_18335,N_18313);
and U18660 (N_18660,N_18384,N_18440);
or U18661 (N_18661,N_18317,N_18446);
nand U18662 (N_18662,N_18300,N_18284);
xor U18663 (N_18663,N_18494,N_18488);
and U18664 (N_18664,N_18298,N_18328);
or U18665 (N_18665,N_18346,N_18434);
and U18666 (N_18666,N_18436,N_18399);
or U18667 (N_18667,N_18325,N_18252);
and U18668 (N_18668,N_18402,N_18274);
nand U18669 (N_18669,N_18266,N_18278);
or U18670 (N_18670,N_18353,N_18412);
or U18671 (N_18671,N_18284,N_18425);
nand U18672 (N_18672,N_18337,N_18475);
and U18673 (N_18673,N_18284,N_18355);
or U18674 (N_18674,N_18444,N_18347);
xnor U18675 (N_18675,N_18272,N_18274);
nor U18676 (N_18676,N_18441,N_18450);
nand U18677 (N_18677,N_18407,N_18271);
xor U18678 (N_18678,N_18360,N_18486);
nor U18679 (N_18679,N_18484,N_18274);
xnor U18680 (N_18680,N_18359,N_18419);
and U18681 (N_18681,N_18384,N_18267);
and U18682 (N_18682,N_18259,N_18468);
or U18683 (N_18683,N_18490,N_18477);
xnor U18684 (N_18684,N_18279,N_18404);
nand U18685 (N_18685,N_18443,N_18317);
and U18686 (N_18686,N_18379,N_18265);
and U18687 (N_18687,N_18498,N_18389);
xnor U18688 (N_18688,N_18300,N_18387);
nand U18689 (N_18689,N_18410,N_18488);
or U18690 (N_18690,N_18437,N_18357);
nor U18691 (N_18691,N_18367,N_18364);
nand U18692 (N_18692,N_18360,N_18347);
nand U18693 (N_18693,N_18424,N_18273);
nand U18694 (N_18694,N_18372,N_18471);
nand U18695 (N_18695,N_18312,N_18318);
nor U18696 (N_18696,N_18363,N_18438);
xor U18697 (N_18697,N_18429,N_18434);
or U18698 (N_18698,N_18401,N_18296);
and U18699 (N_18699,N_18388,N_18442);
nor U18700 (N_18700,N_18360,N_18431);
nand U18701 (N_18701,N_18254,N_18386);
or U18702 (N_18702,N_18404,N_18393);
xor U18703 (N_18703,N_18299,N_18309);
or U18704 (N_18704,N_18454,N_18412);
xnor U18705 (N_18705,N_18372,N_18415);
nand U18706 (N_18706,N_18346,N_18400);
or U18707 (N_18707,N_18304,N_18455);
nand U18708 (N_18708,N_18493,N_18475);
nor U18709 (N_18709,N_18382,N_18283);
nor U18710 (N_18710,N_18411,N_18262);
nor U18711 (N_18711,N_18411,N_18466);
nor U18712 (N_18712,N_18430,N_18372);
or U18713 (N_18713,N_18412,N_18449);
or U18714 (N_18714,N_18342,N_18440);
or U18715 (N_18715,N_18408,N_18289);
xor U18716 (N_18716,N_18402,N_18278);
nand U18717 (N_18717,N_18371,N_18267);
xor U18718 (N_18718,N_18353,N_18432);
nor U18719 (N_18719,N_18270,N_18365);
nor U18720 (N_18720,N_18407,N_18253);
nand U18721 (N_18721,N_18431,N_18419);
nor U18722 (N_18722,N_18272,N_18307);
nor U18723 (N_18723,N_18323,N_18456);
and U18724 (N_18724,N_18437,N_18356);
and U18725 (N_18725,N_18311,N_18429);
and U18726 (N_18726,N_18254,N_18360);
or U18727 (N_18727,N_18405,N_18388);
nand U18728 (N_18728,N_18400,N_18446);
nand U18729 (N_18729,N_18352,N_18440);
xnor U18730 (N_18730,N_18297,N_18440);
and U18731 (N_18731,N_18309,N_18272);
xor U18732 (N_18732,N_18282,N_18396);
xnor U18733 (N_18733,N_18381,N_18449);
or U18734 (N_18734,N_18303,N_18495);
nor U18735 (N_18735,N_18433,N_18265);
nand U18736 (N_18736,N_18311,N_18360);
nand U18737 (N_18737,N_18314,N_18289);
nor U18738 (N_18738,N_18348,N_18330);
and U18739 (N_18739,N_18447,N_18418);
nor U18740 (N_18740,N_18268,N_18331);
nand U18741 (N_18741,N_18299,N_18406);
and U18742 (N_18742,N_18255,N_18254);
nand U18743 (N_18743,N_18469,N_18251);
nor U18744 (N_18744,N_18346,N_18345);
nand U18745 (N_18745,N_18494,N_18324);
nand U18746 (N_18746,N_18432,N_18480);
nor U18747 (N_18747,N_18418,N_18448);
or U18748 (N_18748,N_18407,N_18313);
and U18749 (N_18749,N_18496,N_18493);
xnor U18750 (N_18750,N_18537,N_18682);
nand U18751 (N_18751,N_18550,N_18523);
and U18752 (N_18752,N_18562,N_18587);
and U18753 (N_18753,N_18681,N_18508);
nor U18754 (N_18754,N_18532,N_18571);
nand U18755 (N_18755,N_18737,N_18505);
or U18756 (N_18756,N_18676,N_18703);
nand U18757 (N_18757,N_18654,N_18736);
and U18758 (N_18758,N_18618,N_18626);
xnor U18759 (N_18759,N_18513,N_18563);
xor U18760 (N_18760,N_18664,N_18597);
nand U18761 (N_18761,N_18610,N_18539);
nand U18762 (N_18762,N_18616,N_18666);
nor U18763 (N_18763,N_18500,N_18567);
or U18764 (N_18764,N_18605,N_18714);
and U18765 (N_18765,N_18619,N_18514);
and U18766 (N_18766,N_18633,N_18582);
xnor U18767 (N_18767,N_18733,N_18645);
nor U18768 (N_18768,N_18623,N_18602);
nand U18769 (N_18769,N_18740,N_18564);
and U18770 (N_18770,N_18728,N_18544);
xor U18771 (N_18771,N_18746,N_18519);
xnor U18772 (N_18772,N_18635,N_18691);
and U18773 (N_18773,N_18661,N_18636);
nor U18774 (N_18774,N_18522,N_18684);
or U18775 (N_18775,N_18578,N_18570);
xnor U18776 (N_18776,N_18632,N_18712);
or U18777 (N_18777,N_18656,N_18518);
nand U18778 (N_18778,N_18698,N_18708);
and U18779 (N_18779,N_18615,N_18695);
nand U18780 (N_18780,N_18579,N_18515);
and U18781 (N_18781,N_18548,N_18672);
or U18782 (N_18782,N_18629,N_18685);
nand U18783 (N_18783,N_18652,N_18647);
nand U18784 (N_18784,N_18592,N_18673);
nand U18785 (N_18785,N_18706,N_18517);
nand U18786 (N_18786,N_18699,N_18668);
nor U18787 (N_18787,N_18547,N_18510);
nor U18788 (N_18788,N_18646,N_18671);
nor U18789 (N_18789,N_18509,N_18575);
nand U18790 (N_18790,N_18683,N_18722);
nor U18791 (N_18791,N_18711,N_18614);
xor U18792 (N_18792,N_18576,N_18612);
nand U18793 (N_18793,N_18607,N_18600);
xnor U18794 (N_18794,N_18589,N_18729);
xnor U18795 (N_18795,N_18639,N_18603);
or U18796 (N_18796,N_18637,N_18526);
and U18797 (N_18797,N_18701,N_18546);
nor U18798 (N_18798,N_18549,N_18586);
nand U18799 (N_18799,N_18719,N_18667);
xor U18800 (N_18800,N_18721,N_18558);
and U18801 (N_18801,N_18697,N_18557);
xor U18802 (N_18802,N_18502,N_18627);
xnor U18803 (N_18803,N_18606,N_18609);
and U18804 (N_18804,N_18732,N_18554);
nor U18805 (N_18805,N_18631,N_18731);
nor U18806 (N_18806,N_18555,N_18588);
nor U18807 (N_18807,N_18566,N_18604);
or U18808 (N_18808,N_18662,N_18574);
and U18809 (N_18809,N_18713,N_18601);
nor U18810 (N_18810,N_18584,N_18524);
xor U18811 (N_18811,N_18747,N_18545);
nor U18812 (N_18812,N_18725,N_18677);
nand U18813 (N_18813,N_18577,N_18591);
nand U18814 (N_18814,N_18687,N_18704);
nor U18815 (N_18815,N_18594,N_18533);
nor U18816 (N_18816,N_18534,N_18540);
or U18817 (N_18817,N_18595,N_18613);
xnor U18818 (N_18818,N_18560,N_18658);
nand U18819 (N_18819,N_18700,N_18527);
and U18820 (N_18820,N_18717,N_18599);
xor U18821 (N_18821,N_18749,N_18739);
xnor U18822 (N_18822,N_18742,N_18565);
nand U18823 (N_18823,N_18622,N_18650);
and U18824 (N_18824,N_18596,N_18688);
nand U18825 (N_18825,N_18504,N_18679);
and U18826 (N_18826,N_18724,N_18608);
nand U18827 (N_18827,N_18503,N_18598);
nor U18828 (N_18828,N_18561,N_18669);
nor U18829 (N_18829,N_18634,N_18709);
xnor U18830 (N_18830,N_18638,N_18680);
or U18831 (N_18831,N_18520,N_18674);
or U18832 (N_18832,N_18621,N_18624);
or U18833 (N_18833,N_18593,N_18556);
xor U18834 (N_18834,N_18580,N_18741);
nor U18835 (N_18835,N_18531,N_18748);
and U18836 (N_18836,N_18628,N_18705);
or U18837 (N_18837,N_18653,N_18727);
xnor U18838 (N_18838,N_18541,N_18660);
and U18839 (N_18839,N_18572,N_18516);
nand U18840 (N_18840,N_18644,N_18686);
nor U18841 (N_18841,N_18694,N_18630);
nand U18842 (N_18842,N_18715,N_18665);
nor U18843 (N_18843,N_18501,N_18506);
nand U18844 (N_18844,N_18583,N_18559);
or U18845 (N_18845,N_18670,N_18640);
nand U18846 (N_18846,N_18569,N_18611);
nor U18847 (N_18847,N_18543,N_18625);
and U18848 (N_18848,N_18692,N_18585);
xor U18849 (N_18849,N_18511,N_18529);
nor U18850 (N_18850,N_18743,N_18528);
xor U18851 (N_18851,N_18690,N_18738);
nand U18852 (N_18852,N_18643,N_18590);
nor U18853 (N_18853,N_18651,N_18675);
xnor U18854 (N_18854,N_18551,N_18659);
nand U18855 (N_18855,N_18512,N_18617);
nand U18856 (N_18856,N_18716,N_18521);
nand U18857 (N_18857,N_18710,N_18723);
xnor U18858 (N_18858,N_18720,N_18568);
xor U18859 (N_18859,N_18735,N_18745);
and U18860 (N_18860,N_18581,N_18507);
nor U18861 (N_18861,N_18707,N_18734);
nor U18862 (N_18862,N_18536,N_18642);
or U18863 (N_18863,N_18538,N_18663);
xor U18864 (N_18864,N_18649,N_18573);
and U18865 (N_18865,N_18552,N_18657);
xnor U18866 (N_18866,N_18535,N_18696);
xor U18867 (N_18867,N_18726,N_18718);
nor U18868 (N_18868,N_18542,N_18648);
nand U18869 (N_18869,N_18689,N_18693);
xor U18870 (N_18870,N_18678,N_18530);
and U18871 (N_18871,N_18744,N_18525);
nand U18872 (N_18872,N_18641,N_18702);
nor U18873 (N_18873,N_18553,N_18620);
xnor U18874 (N_18874,N_18730,N_18655);
nand U18875 (N_18875,N_18500,N_18700);
or U18876 (N_18876,N_18502,N_18716);
or U18877 (N_18877,N_18520,N_18533);
xor U18878 (N_18878,N_18679,N_18604);
nand U18879 (N_18879,N_18507,N_18519);
nand U18880 (N_18880,N_18748,N_18602);
and U18881 (N_18881,N_18604,N_18722);
nand U18882 (N_18882,N_18683,N_18637);
nand U18883 (N_18883,N_18628,N_18684);
or U18884 (N_18884,N_18672,N_18730);
xor U18885 (N_18885,N_18534,N_18593);
nand U18886 (N_18886,N_18547,N_18676);
or U18887 (N_18887,N_18600,N_18740);
xnor U18888 (N_18888,N_18642,N_18558);
xnor U18889 (N_18889,N_18515,N_18746);
or U18890 (N_18890,N_18659,N_18535);
and U18891 (N_18891,N_18716,N_18566);
xnor U18892 (N_18892,N_18618,N_18591);
xnor U18893 (N_18893,N_18720,N_18580);
and U18894 (N_18894,N_18500,N_18598);
nand U18895 (N_18895,N_18689,N_18543);
and U18896 (N_18896,N_18737,N_18553);
nand U18897 (N_18897,N_18650,N_18516);
nor U18898 (N_18898,N_18747,N_18722);
xor U18899 (N_18899,N_18542,N_18626);
nand U18900 (N_18900,N_18607,N_18603);
or U18901 (N_18901,N_18516,N_18648);
or U18902 (N_18902,N_18527,N_18592);
nand U18903 (N_18903,N_18726,N_18609);
nor U18904 (N_18904,N_18627,N_18601);
xnor U18905 (N_18905,N_18623,N_18576);
nor U18906 (N_18906,N_18743,N_18747);
or U18907 (N_18907,N_18542,N_18532);
and U18908 (N_18908,N_18583,N_18742);
or U18909 (N_18909,N_18544,N_18634);
nand U18910 (N_18910,N_18537,N_18564);
and U18911 (N_18911,N_18616,N_18633);
or U18912 (N_18912,N_18541,N_18524);
xor U18913 (N_18913,N_18547,N_18589);
xor U18914 (N_18914,N_18513,N_18691);
and U18915 (N_18915,N_18704,N_18618);
xor U18916 (N_18916,N_18710,N_18634);
xnor U18917 (N_18917,N_18500,N_18580);
nand U18918 (N_18918,N_18729,N_18699);
xnor U18919 (N_18919,N_18518,N_18701);
and U18920 (N_18920,N_18746,N_18683);
nand U18921 (N_18921,N_18677,N_18664);
xor U18922 (N_18922,N_18520,N_18691);
nor U18923 (N_18923,N_18536,N_18596);
xnor U18924 (N_18924,N_18632,N_18574);
and U18925 (N_18925,N_18627,N_18691);
and U18926 (N_18926,N_18582,N_18583);
nor U18927 (N_18927,N_18569,N_18697);
and U18928 (N_18928,N_18550,N_18532);
or U18929 (N_18929,N_18687,N_18551);
xor U18930 (N_18930,N_18656,N_18538);
nand U18931 (N_18931,N_18528,N_18748);
xor U18932 (N_18932,N_18607,N_18588);
nor U18933 (N_18933,N_18614,N_18581);
nand U18934 (N_18934,N_18723,N_18621);
xnor U18935 (N_18935,N_18587,N_18620);
and U18936 (N_18936,N_18608,N_18583);
xnor U18937 (N_18937,N_18514,N_18739);
nand U18938 (N_18938,N_18677,N_18652);
and U18939 (N_18939,N_18737,N_18566);
or U18940 (N_18940,N_18575,N_18500);
xnor U18941 (N_18941,N_18557,N_18549);
or U18942 (N_18942,N_18600,N_18572);
or U18943 (N_18943,N_18608,N_18627);
nor U18944 (N_18944,N_18748,N_18536);
nand U18945 (N_18945,N_18653,N_18655);
nand U18946 (N_18946,N_18598,N_18637);
and U18947 (N_18947,N_18520,N_18555);
nor U18948 (N_18948,N_18560,N_18713);
nand U18949 (N_18949,N_18536,N_18731);
nor U18950 (N_18950,N_18592,N_18665);
nor U18951 (N_18951,N_18621,N_18738);
or U18952 (N_18952,N_18642,N_18532);
and U18953 (N_18953,N_18600,N_18624);
and U18954 (N_18954,N_18546,N_18608);
or U18955 (N_18955,N_18622,N_18732);
xor U18956 (N_18956,N_18743,N_18687);
nand U18957 (N_18957,N_18502,N_18703);
xnor U18958 (N_18958,N_18555,N_18648);
or U18959 (N_18959,N_18669,N_18642);
nand U18960 (N_18960,N_18599,N_18746);
nor U18961 (N_18961,N_18738,N_18528);
and U18962 (N_18962,N_18576,N_18729);
and U18963 (N_18963,N_18530,N_18592);
nor U18964 (N_18964,N_18582,N_18748);
nor U18965 (N_18965,N_18575,N_18528);
nand U18966 (N_18966,N_18711,N_18682);
xnor U18967 (N_18967,N_18663,N_18520);
xnor U18968 (N_18968,N_18719,N_18535);
or U18969 (N_18969,N_18606,N_18578);
xor U18970 (N_18970,N_18712,N_18731);
xor U18971 (N_18971,N_18710,N_18567);
and U18972 (N_18972,N_18599,N_18646);
or U18973 (N_18973,N_18619,N_18501);
or U18974 (N_18974,N_18702,N_18606);
and U18975 (N_18975,N_18735,N_18678);
nor U18976 (N_18976,N_18706,N_18503);
or U18977 (N_18977,N_18663,N_18552);
or U18978 (N_18978,N_18565,N_18523);
and U18979 (N_18979,N_18643,N_18527);
nor U18980 (N_18980,N_18672,N_18644);
or U18981 (N_18981,N_18619,N_18749);
nand U18982 (N_18982,N_18698,N_18733);
and U18983 (N_18983,N_18590,N_18644);
nand U18984 (N_18984,N_18717,N_18679);
nand U18985 (N_18985,N_18532,N_18531);
xnor U18986 (N_18986,N_18697,N_18749);
xor U18987 (N_18987,N_18707,N_18591);
xor U18988 (N_18988,N_18721,N_18584);
nand U18989 (N_18989,N_18686,N_18621);
xor U18990 (N_18990,N_18511,N_18705);
xor U18991 (N_18991,N_18514,N_18748);
xor U18992 (N_18992,N_18531,N_18578);
nand U18993 (N_18993,N_18608,N_18554);
nand U18994 (N_18994,N_18548,N_18730);
xor U18995 (N_18995,N_18628,N_18689);
xor U18996 (N_18996,N_18537,N_18651);
xnor U18997 (N_18997,N_18745,N_18501);
nor U18998 (N_18998,N_18547,N_18524);
nor U18999 (N_18999,N_18615,N_18648);
or U19000 (N_19000,N_18932,N_18838);
nor U19001 (N_19001,N_18832,N_18942);
or U19002 (N_19002,N_18877,N_18906);
nor U19003 (N_19003,N_18813,N_18983);
nor U19004 (N_19004,N_18885,N_18995);
nor U19005 (N_19005,N_18764,N_18848);
and U19006 (N_19006,N_18771,N_18962);
and U19007 (N_19007,N_18947,N_18815);
nor U19008 (N_19008,N_18905,N_18992);
or U19009 (N_19009,N_18913,N_18978);
xnor U19010 (N_19010,N_18860,N_18951);
xor U19011 (N_19011,N_18984,N_18914);
or U19012 (N_19012,N_18895,N_18946);
nand U19013 (N_19013,N_18757,N_18909);
and U19014 (N_19014,N_18840,N_18948);
nor U19015 (N_19015,N_18907,N_18869);
nand U19016 (N_19016,N_18940,N_18896);
xor U19017 (N_19017,N_18780,N_18875);
or U19018 (N_19018,N_18965,N_18761);
or U19019 (N_19019,N_18822,N_18765);
or U19020 (N_19020,N_18827,N_18835);
xnor U19021 (N_19021,N_18849,N_18981);
nor U19022 (N_19022,N_18982,N_18778);
nor U19023 (N_19023,N_18831,N_18891);
xnor U19024 (N_19024,N_18814,N_18911);
xor U19025 (N_19025,N_18949,N_18921);
and U19026 (N_19026,N_18971,N_18816);
or U19027 (N_19027,N_18766,N_18867);
or U19028 (N_19028,N_18807,N_18991);
nor U19029 (N_19029,N_18989,N_18900);
and U19030 (N_19030,N_18936,N_18927);
nand U19031 (N_19031,N_18868,N_18833);
or U19032 (N_19032,N_18985,N_18776);
xor U19033 (N_19033,N_18830,N_18783);
or U19034 (N_19034,N_18812,N_18853);
xnor U19035 (N_19035,N_18821,N_18934);
and U19036 (N_19036,N_18829,N_18800);
nand U19037 (N_19037,N_18987,N_18820);
nor U19038 (N_19038,N_18990,N_18902);
and U19039 (N_19039,N_18903,N_18836);
xor U19040 (N_19040,N_18953,N_18861);
nand U19041 (N_19041,N_18882,N_18808);
and U19042 (N_19042,N_18923,N_18975);
nand U19043 (N_19043,N_18873,N_18912);
and U19044 (N_19044,N_18837,N_18925);
and U19045 (N_19045,N_18939,N_18889);
and U19046 (N_19046,N_18928,N_18762);
or U19047 (N_19047,N_18781,N_18917);
nand U19048 (N_19048,N_18842,N_18870);
nor U19049 (N_19049,N_18892,N_18858);
xor U19050 (N_19050,N_18960,N_18810);
nand U19051 (N_19051,N_18930,N_18834);
and U19052 (N_19052,N_18996,N_18846);
nand U19053 (N_19053,N_18938,N_18943);
xor U19054 (N_19054,N_18802,N_18750);
nor U19055 (N_19055,N_18931,N_18797);
nand U19056 (N_19056,N_18769,N_18796);
or U19057 (N_19057,N_18919,N_18997);
and U19058 (N_19058,N_18878,N_18804);
and U19059 (N_19059,N_18809,N_18844);
nand U19060 (N_19060,N_18920,N_18979);
and U19061 (N_19061,N_18972,N_18763);
and U19062 (N_19062,N_18785,N_18863);
xnor U19063 (N_19063,N_18824,N_18897);
nor U19064 (N_19064,N_18803,N_18888);
xnor U19065 (N_19065,N_18999,N_18904);
and U19066 (N_19066,N_18973,N_18899);
nor U19067 (N_19067,N_18886,N_18841);
nand U19068 (N_19068,N_18890,N_18941);
or U19069 (N_19069,N_18933,N_18944);
or U19070 (N_19070,N_18767,N_18986);
or U19071 (N_19071,N_18789,N_18794);
and U19072 (N_19072,N_18828,N_18759);
nor U19073 (N_19073,N_18924,N_18792);
nor U19074 (N_19074,N_18819,N_18855);
xnor U19075 (N_19075,N_18798,N_18806);
nand U19076 (N_19076,N_18976,N_18922);
nor U19077 (N_19077,N_18864,N_18876);
nor U19078 (N_19078,N_18970,N_18856);
and U19079 (N_19079,N_18774,N_18773);
and U19080 (N_19080,N_18751,N_18926);
nand U19081 (N_19081,N_18883,N_18854);
xnor U19082 (N_19082,N_18880,N_18817);
or U19083 (N_19083,N_18811,N_18957);
or U19084 (N_19084,N_18994,N_18908);
nand U19085 (N_19085,N_18754,N_18801);
xnor U19086 (N_19086,N_18850,N_18799);
nor U19087 (N_19087,N_18969,N_18977);
nand U19088 (N_19088,N_18839,N_18859);
or U19089 (N_19089,N_18788,N_18825);
and U19090 (N_19090,N_18893,N_18756);
or U19091 (N_19091,N_18775,N_18760);
or U19092 (N_19092,N_18918,N_18966);
xnor U19093 (N_19093,N_18935,N_18787);
nor U19094 (N_19094,N_18964,N_18955);
nor U19095 (N_19095,N_18950,N_18866);
xnor U19096 (N_19096,N_18937,N_18768);
nor U19097 (N_19097,N_18872,N_18887);
xor U19098 (N_19098,N_18777,N_18770);
xor U19099 (N_19099,N_18784,N_18793);
and U19100 (N_19100,N_18898,N_18884);
xnor U19101 (N_19101,N_18786,N_18871);
and U19102 (N_19102,N_18755,N_18790);
nand U19103 (N_19103,N_18874,N_18782);
and U19104 (N_19104,N_18963,N_18881);
xor U19105 (N_19105,N_18865,N_18956);
nand U19106 (N_19106,N_18954,N_18980);
xnor U19107 (N_19107,N_18805,N_18952);
nand U19108 (N_19108,N_18993,N_18845);
xor U19109 (N_19109,N_18752,N_18910);
nand U19110 (N_19110,N_18901,N_18958);
nor U19111 (N_19111,N_18974,N_18823);
or U19112 (N_19112,N_18929,N_18772);
or U19113 (N_19113,N_18988,N_18857);
and U19114 (N_19114,N_18852,N_18753);
or U19115 (N_19115,N_18998,N_18894);
and U19116 (N_19116,N_18916,N_18961);
and U19117 (N_19117,N_18915,N_18968);
nor U19118 (N_19118,N_18791,N_18779);
xor U19119 (N_19119,N_18945,N_18851);
nand U19120 (N_19120,N_18959,N_18818);
xor U19121 (N_19121,N_18826,N_18879);
nor U19122 (N_19122,N_18758,N_18967);
and U19123 (N_19123,N_18862,N_18795);
or U19124 (N_19124,N_18843,N_18847);
and U19125 (N_19125,N_18941,N_18753);
or U19126 (N_19126,N_18901,N_18897);
or U19127 (N_19127,N_18872,N_18814);
nor U19128 (N_19128,N_18878,N_18852);
or U19129 (N_19129,N_18786,N_18875);
xnor U19130 (N_19130,N_18945,N_18890);
and U19131 (N_19131,N_18913,N_18937);
and U19132 (N_19132,N_18824,N_18820);
xnor U19133 (N_19133,N_18962,N_18903);
nor U19134 (N_19134,N_18759,N_18938);
nor U19135 (N_19135,N_18821,N_18940);
nor U19136 (N_19136,N_18796,N_18879);
nand U19137 (N_19137,N_18914,N_18983);
and U19138 (N_19138,N_18788,N_18813);
nor U19139 (N_19139,N_18948,N_18893);
xnor U19140 (N_19140,N_18825,N_18900);
xnor U19141 (N_19141,N_18854,N_18944);
and U19142 (N_19142,N_18874,N_18899);
nand U19143 (N_19143,N_18834,N_18860);
nor U19144 (N_19144,N_18848,N_18909);
xor U19145 (N_19145,N_18888,N_18856);
and U19146 (N_19146,N_18980,N_18783);
nor U19147 (N_19147,N_18919,N_18846);
nor U19148 (N_19148,N_18943,N_18908);
nor U19149 (N_19149,N_18755,N_18895);
nor U19150 (N_19150,N_18864,N_18859);
xnor U19151 (N_19151,N_18871,N_18828);
or U19152 (N_19152,N_18867,N_18974);
nand U19153 (N_19153,N_18939,N_18819);
nor U19154 (N_19154,N_18876,N_18987);
nor U19155 (N_19155,N_18791,N_18784);
or U19156 (N_19156,N_18936,N_18838);
and U19157 (N_19157,N_18981,N_18998);
nor U19158 (N_19158,N_18878,N_18932);
nor U19159 (N_19159,N_18859,N_18990);
or U19160 (N_19160,N_18896,N_18764);
nand U19161 (N_19161,N_18997,N_18896);
xor U19162 (N_19162,N_18811,N_18932);
nand U19163 (N_19163,N_18762,N_18809);
or U19164 (N_19164,N_18939,N_18909);
nand U19165 (N_19165,N_18975,N_18889);
xor U19166 (N_19166,N_18803,N_18910);
xor U19167 (N_19167,N_18844,N_18875);
and U19168 (N_19168,N_18975,N_18779);
nand U19169 (N_19169,N_18790,N_18869);
xnor U19170 (N_19170,N_18973,N_18926);
nor U19171 (N_19171,N_18858,N_18808);
or U19172 (N_19172,N_18962,N_18856);
and U19173 (N_19173,N_18906,N_18750);
xor U19174 (N_19174,N_18875,N_18937);
xor U19175 (N_19175,N_18939,N_18915);
nand U19176 (N_19176,N_18889,N_18752);
nand U19177 (N_19177,N_18948,N_18947);
nand U19178 (N_19178,N_18910,N_18905);
nor U19179 (N_19179,N_18866,N_18820);
xor U19180 (N_19180,N_18940,N_18961);
nor U19181 (N_19181,N_18825,N_18840);
nand U19182 (N_19182,N_18797,N_18810);
xor U19183 (N_19183,N_18751,N_18895);
xor U19184 (N_19184,N_18933,N_18891);
or U19185 (N_19185,N_18859,N_18858);
or U19186 (N_19186,N_18861,N_18982);
nor U19187 (N_19187,N_18789,N_18874);
nor U19188 (N_19188,N_18796,N_18840);
nor U19189 (N_19189,N_18948,N_18901);
xor U19190 (N_19190,N_18943,N_18911);
nor U19191 (N_19191,N_18977,N_18840);
or U19192 (N_19192,N_18976,N_18762);
nor U19193 (N_19193,N_18906,N_18834);
or U19194 (N_19194,N_18888,N_18765);
nand U19195 (N_19195,N_18866,N_18994);
and U19196 (N_19196,N_18819,N_18785);
nand U19197 (N_19197,N_18884,N_18918);
nor U19198 (N_19198,N_18751,N_18769);
and U19199 (N_19199,N_18971,N_18860);
or U19200 (N_19200,N_18953,N_18993);
and U19201 (N_19201,N_18962,N_18754);
nor U19202 (N_19202,N_18763,N_18918);
xor U19203 (N_19203,N_18962,N_18848);
and U19204 (N_19204,N_18948,N_18922);
or U19205 (N_19205,N_18996,N_18864);
nor U19206 (N_19206,N_18754,N_18798);
xnor U19207 (N_19207,N_18997,N_18772);
nand U19208 (N_19208,N_18996,N_18792);
or U19209 (N_19209,N_18867,N_18895);
nor U19210 (N_19210,N_18803,N_18935);
nand U19211 (N_19211,N_18950,N_18827);
xnor U19212 (N_19212,N_18883,N_18912);
and U19213 (N_19213,N_18817,N_18847);
nand U19214 (N_19214,N_18889,N_18809);
xor U19215 (N_19215,N_18998,N_18820);
and U19216 (N_19216,N_18814,N_18968);
and U19217 (N_19217,N_18922,N_18970);
and U19218 (N_19218,N_18771,N_18894);
nor U19219 (N_19219,N_18795,N_18857);
nand U19220 (N_19220,N_18882,N_18951);
nor U19221 (N_19221,N_18935,N_18819);
xor U19222 (N_19222,N_18778,N_18899);
and U19223 (N_19223,N_18979,N_18935);
nor U19224 (N_19224,N_18979,N_18981);
and U19225 (N_19225,N_18890,N_18891);
or U19226 (N_19226,N_18861,N_18930);
and U19227 (N_19227,N_18771,N_18847);
or U19228 (N_19228,N_18884,N_18930);
nand U19229 (N_19229,N_18864,N_18916);
and U19230 (N_19230,N_18850,N_18938);
nor U19231 (N_19231,N_18764,N_18926);
xnor U19232 (N_19232,N_18822,N_18848);
xnor U19233 (N_19233,N_18811,N_18980);
nand U19234 (N_19234,N_18791,N_18938);
xor U19235 (N_19235,N_18911,N_18848);
nand U19236 (N_19236,N_18901,N_18973);
xnor U19237 (N_19237,N_18980,N_18958);
nand U19238 (N_19238,N_18954,N_18913);
nand U19239 (N_19239,N_18843,N_18906);
xnor U19240 (N_19240,N_18849,N_18787);
xnor U19241 (N_19241,N_18861,N_18845);
nand U19242 (N_19242,N_18899,N_18806);
nand U19243 (N_19243,N_18940,N_18825);
nand U19244 (N_19244,N_18959,N_18794);
xnor U19245 (N_19245,N_18923,N_18913);
xor U19246 (N_19246,N_18843,N_18763);
or U19247 (N_19247,N_18985,N_18795);
nor U19248 (N_19248,N_18980,N_18946);
and U19249 (N_19249,N_18881,N_18830);
xnor U19250 (N_19250,N_19118,N_19119);
xor U19251 (N_19251,N_19171,N_19202);
or U19252 (N_19252,N_19134,N_19074);
nand U19253 (N_19253,N_19136,N_19093);
nor U19254 (N_19254,N_19002,N_19138);
nor U19255 (N_19255,N_19054,N_19009);
nand U19256 (N_19256,N_19063,N_19004);
or U19257 (N_19257,N_19192,N_19066);
nor U19258 (N_19258,N_19064,N_19200);
xor U19259 (N_19259,N_19082,N_19198);
and U19260 (N_19260,N_19079,N_19100);
nand U19261 (N_19261,N_19097,N_19163);
nor U19262 (N_19262,N_19104,N_19206);
nand U19263 (N_19263,N_19006,N_19039);
nand U19264 (N_19264,N_19193,N_19061);
nand U19265 (N_19265,N_19130,N_19166);
nor U19266 (N_19266,N_19022,N_19249);
or U19267 (N_19267,N_19209,N_19232);
nor U19268 (N_19268,N_19145,N_19129);
or U19269 (N_19269,N_19148,N_19019);
nor U19270 (N_19270,N_19159,N_19011);
nor U19271 (N_19271,N_19229,N_19131);
nor U19272 (N_19272,N_19184,N_19243);
and U19273 (N_19273,N_19091,N_19246);
xor U19274 (N_19274,N_19121,N_19228);
nor U19275 (N_19275,N_19141,N_19245);
nand U19276 (N_19276,N_19216,N_19111);
and U19277 (N_19277,N_19175,N_19040);
or U19278 (N_19278,N_19047,N_19168);
and U19279 (N_19279,N_19089,N_19109);
nand U19280 (N_19280,N_19084,N_19146);
or U19281 (N_19281,N_19036,N_19115);
and U19282 (N_19282,N_19230,N_19113);
xnor U19283 (N_19283,N_19194,N_19218);
xor U19284 (N_19284,N_19075,N_19023);
xnor U19285 (N_19285,N_19030,N_19083);
and U19286 (N_19286,N_19003,N_19045);
xor U19287 (N_19287,N_19162,N_19067);
xnor U19288 (N_19288,N_19122,N_19173);
nand U19289 (N_19289,N_19087,N_19211);
and U19290 (N_19290,N_19053,N_19106);
or U19291 (N_19291,N_19167,N_19048);
xor U19292 (N_19292,N_19239,N_19013);
xor U19293 (N_19293,N_19227,N_19070);
nor U19294 (N_19294,N_19028,N_19116);
nand U19295 (N_19295,N_19186,N_19103);
nand U19296 (N_19296,N_19024,N_19157);
or U19297 (N_19297,N_19078,N_19038);
nand U19298 (N_19298,N_19219,N_19085);
and U19299 (N_19299,N_19077,N_19164);
nand U19300 (N_19300,N_19076,N_19179);
xor U19301 (N_19301,N_19247,N_19195);
and U19302 (N_19302,N_19191,N_19213);
xor U19303 (N_19303,N_19026,N_19010);
xor U19304 (N_19304,N_19094,N_19062);
and U19305 (N_19305,N_19034,N_19222);
xor U19306 (N_19306,N_19199,N_19043);
nand U19307 (N_19307,N_19095,N_19244);
or U19308 (N_19308,N_19234,N_19088);
nor U19309 (N_19309,N_19236,N_19041);
nor U19310 (N_19310,N_19126,N_19016);
nand U19311 (N_19311,N_19226,N_19144);
xor U19312 (N_19312,N_19224,N_19137);
nor U19313 (N_19313,N_19059,N_19102);
nand U19314 (N_19314,N_19117,N_19032);
and U19315 (N_19315,N_19182,N_19021);
nand U19316 (N_19316,N_19001,N_19203);
or U19317 (N_19317,N_19014,N_19073);
nand U19318 (N_19318,N_19237,N_19196);
nor U19319 (N_19319,N_19248,N_19049);
or U19320 (N_19320,N_19133,N_19174);
xnor U19321 (N_19321,N_19052,N_19205);
and U19322 (N_19322,N_19156,N_19068);
nor U19323 (N_19323,N_19210,N_19132);
nand U19324 (N_19324,N_19207,N_19112);
and U19325 (N_19325,N_19212,N_19037);
xor U19326 (N_19326,N_19238,N_19181);
xor U19327 (N_19327,N_19046,N_19050);
or U19328 (N_19328,N_19217,N_19072);
xor U19329 (N_19329,N_19015,N_19044);
xor U19330 (N_19330,N_19105,N_19086);
or U19331 (N_19331,N_19235,N_19185);
or U19332 (N_19332,N_19081,N_19018);
or U19333 (N_19333,N_19177,N_19140);
nor U19334 (N_19334,N_19080,N_19169);
and U19335 (N_19335,N_19127,N_19142);
nor U19336 (N_19336,N_19007,N_19124);
xor U19337 (N_19337,N_19020,N_19178);
xnor U19338 (N_19338,N_19208,N_19005);
nor U19339 (N_19339,N_19151,N_19051);
xnor U19340 (N_19340,N_19033,N_19096);
nor U19341 (N_19341,N_19110,N_19042);
nand U19342 (N_19342,N_19135,N_19204);
xor U19343 (N_19343,N_19108,N_19147);
xor U19344 (N_19344,N_19000,N_19240);
xor U19345 (N_19345,N_19183,N_19180);
nor U19346 (N_19346,N_19154,N_19187);
nor U19347 (N_19347,N_19158,N_19017);
xnor U19348 (N_19348,N_19143,N_19128);
and U19349 (N_19349,N_19223,N_19214);
and U19350 (N_19350,N_19225,N_19092);
nand U19351 (N_19351,N_19139,N_19152);
or U19352 (N_19352,N_19025,N_19165);
xnor U19353 (N_19353,N_19149,N_19057);
nand U19354 (N_19354,N_19233,N_19056);
nand U19355 (N_19355,N_19170,N_19221);
xnor U19356 (N_19356,N_19155,N_19031);
nor U19357 (N_19357,N_19101,N_19190);
nor U19358 (N_19358,N_19058,N_19197);
nand U19359 (N_19359,N_19125,N_19069);
nand U19360 (N_19360,N_19160,N_19241);
nand U19361 (N_19361,N_19153,N_19188);
nand U19362 (N_19362,N_19231,N_19114);
nand U19363 (N_19363,N_19012,N_19242);
nor U19364 (N_19364,N_19107,N_19065);
and U19365 (N_19365,N_19220,N_19090);
or U19366 (N_19366,N_19176,N_19189);
or U19367 (N_19367,N_19161,N_19120);
and U19368 (N_19368,N_19060,N_19215);
nand U19369 (N_19369,N_19008,N_19035);
or U19370 (N_19370,N_19027,N_19029);
nand U19371 (N_19371,N_19055,N_19172);
nand U19372 (N_19372,N_19071,N_19098);
or U19373 (N_19373,N_19123,N_19150);
nor U19374 (N_19374,N_19201,N_19099);
and U19375 (N_19375,N_19215,N_19239);
and U19376 (N_19376,N_19060,N_19051);
or U19377 (N_19377,N_19154,N_19176);
or U19378 (N_19378,N_19018,N_19028);
nand U19379 (N_19379,N_19229,N_19083);
xor U19380 (N_19380,N_19058,N_19209);
or U19381 (N_19381,N_19198,N_19241);
nand U19382 (N_19382,N_19040,N_19009);
xnor U19383 (N_19383,N_19013,N_19104);
or U19384 (N_19384,N_19100,N_19060);
nor U19385 (N_19385,N_19089,N_19063);
xnor U19386 (N_19386,N_19153,N_19114);
and U19387 (N_19387,N_19015,N_19211);
xor U19388 (N_19388,N_19005,N_19209);
xnor U19389 (N_19389,N_19195,N_19212);
xnor U19390 (N_19390,N_19137,N_19065);
nor U19391 (N_19391,N_19116,N_19067);
and U19392 (N_19392,N_19011,N_19172);
and U19393 (N_19393,N_19036,N_19229);
and U19394 (N_19394,N_19002,N_19100);
or U19395 (N_19395,N_19140,N_19192);
and U19396 (N_19396,N_19152,N_19142);
nand U19397 (N_19397,N_19073,N_19211);
and U19398 (N_19398,N_19079,N_19011);
xnor U19399 (N_19399,N_19153,N_19088);
xor U19400 (N_19400,N_19056,N_19068);
and U19401 (N_19401,N_19237,N_19140);
nand U19402 (N_19402,N_19230,N_19194);
xor U19403 (N_19403,N_19138,N_19133);
or U19404 (N_19404,N_19166,N_19109);
nand U19405 (N_19405,N_19162,N_19179);
xnor U19406 (N_19406,N_19148,N_19230);
nor U19407 (N_19407,N_19246,N_19074);
xor U19408 (N_19408,N_19134,N_19034);
or U19409 (N_19409,N_19211,N_19145);
nor U19410 (N_19410,N_19211,N_19146);
xnor U19411 (N_19411,N_19024,N_19079);
nor U19412 (N_19412,N_19020,N_19009);
nor U19413 (N_19413,N_19209,N_19199);
and U19414 (N_19414,N_19008,N_19056);
nand U19415 (N_19415,N_19127,N_19020);
nor U19416 (N_19416,N_19152,N_19001);
nand U19417 (N_19417,N_19221,N_19004);
or U19418 (N_19418,N_19058,N_19082);
xor U19419 (N_19419,N_19102,N_19118);
xor U19420 (N_19420,N_19027,N_19118);
nor U19421 (N_19421,N_19205,N_19110);
and U19422 (N_19422,N_19042,N_19130);
nand U19423 (N_19423,N_19173,N_19142);
xnor U19424 (N_19424,N_19170,N_19141);
and U19425 (N_19425,N_19086,N_19097);
xor U19426 (N_19426,N_19089,N_19102);
and U19427 (N_19427,N_19117,N_19014);
nor U19428 (N_19428,N_19230,N_19102);
or U19429 (N_19429,N_19228,N_19204);
xnor U19430 (N_19430,N_19049,N_19117);
xnor U19431 (N_19431,N_19241,N_19210);
nor U19432 (N_19432,N_19021,N_19248);
nor U19433 (N_19433,N_19002,N_19186);
xnor U19434 (N_19434,N_19135,N_19200);
xor U19435 (N_19435,N_19096,N_19011);
or U19436 (N_19436,N_19085,N_19234);
nand U19437 (N_19437,N_19142,N_19133);
or U19438 (N_19438,N_19024,N_19026);
nand U19439 (N_19439,N_19209,N_19014);
xor U19440 (N_19440,N_19051,N_19054);
nor U19441 (N_19441,N_19135,N_19220);
nand U19442 (N_19442,N_19004,N_19079);
nand U19443 (N_19443,N_19157,N_19242);
and U19444 (N_19444,N_19002,N_19196);
or U19445 (N_19445,N_19097,N_19232);
nor U19446 (N_19446,N_19237,N_19167);
xnor U19447 (N_19447,N_19212,N_19005);
or U19448 (N_19448,N_19207,N_19038);
or U19449 (N_19449,N_19078,N_19022);
and U19450 (N_19450,N_19139,N_19233);
or U19451 (N_19451,N_19223,N_19099);
nor U19452 (N_19452,N_19224,N_19131);
or U19453 (N_19453,N_19182,N_19097);
nand U19454 (N_19454,N_19152,N_19161);
nand U19455 (N_19455,N_19070,N_19087);
and U19456 (N_19456,N_19025,N_19046);
nand U19457 (N_19457,N_19117,N_19170);
or U19458 (N_19458,N_19158,N_19021);
or U19459 (N_19459,N_19233,N_19052);
nor U19460 (N_19460,N_19119,N_19030);
or U19461 (N_19461,N_19018,N_19107);
or U19462 (N_19462,N_19154,N_19134);
nand U19463 (N_19463,N_19090,N_19187);
or U19464 (N_19464,N_19136,N_19106);
nor U19465 (N_19465,N_19005,N_19106);
or U19466 (N_19466,N_19180,N_19194);
nor U19467 (N_19467,N_19091,N_19094);
or U19468 (N_19468,N_19111,N_19170);
nor U19469 (N_19469,N_19096,N_19085);
and U19470 (N_19470,N_19003,N_19182);
xor U19471 (N_19471,N_19194,N_19197);
and U19472 (N_19472,N_19184,N_19002);
and U19473 (N_19473,N_19049,N_19216);
xor U19474 (N_19474,N_19221,N_19243);
xnor U19475 (N_19475,N_19062,N_19030);
nand U19476 (N_19476,N_19006,N_19204);
and U19477 (N_19477,N_19054,N_19053);
nand U19478 (N_19478,N_19148,N_19110);
nand U19479 (N_19479,N_19002,N_19245);
or U19480 (N_19480,N_19103,N_19109);
nor U19481 (N_19481,N_19103,N_19239);
xnor U19482 (N_19482,N_19238,N_19228);
and U19483 (N_19483,N_19233,N_19115);
nor U19484 (N_19484,N_19214,N_19042);
or U19485 (N_19485,N_19180,N_19031);
nand U19486 (N_19486,N_19086,N_19059);
nor U19487 (N_19487,N_19051,N_19108);
or U19488 (N_19488,N_19119,N_19207);
nand U19489 (N_19489,N_19216,N_19071);
and U19490 (N_19490,N_19024,N_19153);
xnor U19491 (N_19491,N_19239,N_19221);
or U19492 (N_19492,N_19141,N_19179);
nor U19493 (N_19493,N_19101,N_19001);
or U19494 (N_19494,N_19102,N_19084);
nand U19495 (N_19495,N_19195,N_19153);
and U19496 (N_19496,N_19101,N_19156);
or U19497 (N_19497,N_19045,N_19147);
and U19498 (N_19498,N_19177,N_19040);
nor U19499 (N_19499,N_19155,N_19113);
nor U19500 (N_19500,N_19492,N_19316);
or U19501 (N_19501,N_19366,N_19350);
nor U19502 (N_19502,N_19395,N_19482);
nand U19503 (N_19503,N_19352,N_19456);
and U19504 (N_19504,N_19369,N_19406);
nand U19505 (N_19505,N_19301,N_19266);
nand U19506 (N_19506,N_19341,N_19373);
and U19507 (N_19507,N_19409,N_19273);
nor U19508 (N_19508,N_19302,N_19453);
and U19509 (N_19509,N_19441,N_19313);
xnor U19510 (N_19510,N_19436,N_19268);
and U19511 (N_19511,N_19413,N_19357);
or U19512 (N_19512,N_19274,N_19472);
and U19513 (N_19513,N_19499,N_19279);
nand U19514 (N_19514,N_19392,N_19495);
xor U19515 (N_19515,N_19332,N_19254);
xnor U19516 (N_19516,N_19337,N_19293);
xor U19517 (N_19517,N_19464,N_19407);
or U19518 (N_19518,N_19402,N_19346);
xor U19519 (N_19519,N_19351,N_19281);
and U19520 (N_19520,N_19416,N_19287);
or U19521 (N_19521,N_19421,N_19449);
xor U19522 (N_19522,N_19305,N_19419);
xor U19523 (N_19523,N_19426,N_19312);
nor U19524 (N_19524,N_19380,N_19272);
nand U19525 (N_19525,N_19418,N_19448);
or U19526 (N_19526,N_19251,N_19289);
nand U19527 (N_19527,N_19378,N_19300);
nand U19528 (N_19528,N_19461,N_19423);
and U19529 (N_19529,N_19259,N_19280);
nor U19530 (N_19530,N_19282,N_19382);
xnor U19531 (N_19531,N_19438,N_19454);
or U19532 (N_19532,N_19435,N_19466);
xnor U19533 (N_19533,N_19473,N_19362);
nor U19534 (N_19534,N_19304,N_19404);
xnor U19535 (N_19535,N_19487,N_19260);
and U19536 (N_19536,N_19445,N_19458);
or U19537 (N_19537,N_19256,N_19481);
nand U19538 (N_19538,N_19286,N_19315);
xor U19539 (N_19539,N_19360,N_19470);
or U19540 (N_19540,N_19322,N_19451);
nor U19541 (N_19541,N_19271,N_19390);
xor U19542 (N_19542,N_19307,N_19348);
or U19543 (N_19543,N_19338,N_19463);
and U19544 (N_19544,N_19469,N_19399);
xnor U19545 (N_19545,N_19371,N_19270);
xnor U19546 (N_19546,N_19319,N_19494);
xnor U19547 (N_19547,N_19465,N_19411);
and U19548 (N_19548,N_19468,N_19292);
or U19549 (N_19549,N_19389,N_19427);
nand U19550 (N_19550,N_19335,N_19276);
xnor U19551 (N_19551,N_19384,N_19347);
nor U19552 (N_19552,N_19367,N_19308);
nor U19553 (N_19553,N_19283,N_19264);
nand U19554 (N_19554,N_19326,N_19471);
nand U19555 (N_19555,N_19364,N_19269);
xor U19556 (N_19556,N_19342,N_19432);
and U19557 (N_19557,N_19320,N_19467);
nor U19558 (N_19558,N_19354,N_19333);
and U19559 (N_19559,N_19314,N_19412);
or U19560 (N_19560,N_19379,N_19370);
or U19561 (N_19561,N_19285,N_19368);
or U19562 (N_19562,N_19299,N_19277);
nor U19563 (N_19563,N_19400,N_19278);
or U19564 (N_19564,N_19457,N_19284);
and U19565 (N_19565,N_19394,N_19345);
and U19566 (N_19566,N_19397,N_19252);
and U19567 (N_19567,N_19443,N_19340);
nand U19568 (N_19568,N_19358,N_19425);
nor U19569 (N_19569,N_19475,N_19306);
xnor U19570 (N_19570,N_19349,N_19330);
nor U19571 (N_19571,N_19258,N_19297);
or U19572 (N_19572,N_19477,N_19429);
nor U19573 (N_19573,N_19359,N_19459);
or U19574 (N_19574,N_19396,N_19462);
nand U19575 (N_19575,N_19493,N_19414);
nand U19576 (N_19576,N_19440,N_19336);
nor U19577 (N_19577,N_19329,N_19321);
nor U19578 (N_19578,N_19262,N_19415);
or U19579 (N_19579,N_19491,N_19444);
and U19580 (N_19580,N_19486,N_19331);
or U19581 (N_19581,N_19478,N_19497);
and U19582 (N_19582,N_19383,N_19265);
and U19583 (N_19583,N_19257,N_19328);
nand U19584 (N_19584,N_19489,N_19485);
nor U19585 (N_19585,N_19311,N_19339);
or U19586 (N_19586,N_19488,N_19317);
nor U19587 (N_19587,N_19401,N_19261);
xnor U19588 (N_19588,N_19430,N_19385);
or U19589 (N_19589,N_19355,N_19388);
nand U19590 (N_19590,N_19496,N_19442);
nand U19591 (N_19591,N_19403,N_19408);
nand U19592 (N_19592,N_19476,N_19250);
and U19593 (N_19593,N_19327,N_19428);
and U19594 (N_19594,N_19291,N_19361);
nor U19595 (N_19595,N_19267,N_19376);
and U19596 (N_19596,N_19363,N_19295);
nand U19597 (N_19597,N_19447,N_19298);
xnor U19598 (N_19598,N_19323,N_19391);
or U19599 (N_19599,N_19431,N_19460);
or U19600 (N_19600,N_19433,N_19424);
and U19601 (N_19601,N_19381,N_19479);
and U19602 (N_19602,N_19325,N_19417);
or U19603 (N_19603,N_19375,N_19455);
nor U19604 (N_19604,N_19318,N_19253);
nand U19605 (N_19605,N_19498,N_19446);
or U19606 (N_19606,N_19365,N_19309);
and U19607 (N_19607,N_19263,N_19303);
nor U19608 (N_19608,N_19290,N_19393);
or U19609 (N_19609,N_19324,N_19386);
xor U19610 (N_19610,N_19377,N_19398);
and U19611 (N_19611,N_19296,N_19353);
xnor U19612 (N_19612,N_19356,N_19422);
nand U19613 (N_19613,N_19334,N_19483);
or U19614 (N_19614,N_19437,N_19344);
nor U19615 (N_19615,N_19374,N_19310);
nand U19616 (N_19616,N_19490,N_19452);
nand U19617 (N_19617,N_19372,N_19405);
and U19618 (N_19618,N_19255,N_19294);
or U19619 (N_19619,N_19387,N_19480);
nand U19620 (N_19620,N_19288,N_19410);
and U19621 (N_19621,N_19450,N_19484);
or U19622 (N_19622,N_19275,N_19434);
or U19623 (N_19623,N_19420,N_19439);
or U19624 (N_19624,N_19474,N_19343);
nand U19625 (N_19625,N_19314,N_19360);
xor U19626 (N_19626,N_19320,N_19270);
nor U19627 (N_19627,N_19410,N_19417);
nand U19628 (N_19628,N_19390,N_19480);
or U19629 (N_19629,N_19280,N_19392);
and U19630 (N_19630,N_19431,N_19480);
or U19631 (N_19631,N_19339,N_19317);
or U19632 (N_19632,N_19316,N_19468);
and U19633 (N_19633,N_19440,N_19301);
and U19634 (N_19634,N_19349,N_19481);
xor U19635 (N_19635,N_19455,N_19418);
and U19636 (N_19636,N_19430,N_19428);
xor U19637 (N_19637,N_19342,N_19294);
nand U19638 (N_19638,N_19363,N_19434);
or U19639 (N_19639,N_19450,N_19332);
or U19640 (N_19640,N_19438,N_19476);
nand U19641 (N_19641,N_19297,N_19406);
xor U19642 (N_19642,N_19307,N_19474);
nor U19643 (N_19643,N_19378,N_19279);
or U19644 (N_19644,N_19468,N_19374);
nor U19645 (N_19645,N_19340,N_19468);
nand U19646 (N_19646,N_19480,N_19324);
or U19647 (N_19647,N_19299,N_19287);
and U19648 (N_19648,N_19306,N_19470);
and U19649 (N_19649,N_19265,N_19400);
and U19650 (N_19650,N_19407,N_19277);
xnor U19651 (N_19651,N_19499,N_19337);
xnor U19652 (N_19652,N_19490,N_19460);
xnor U19653 (N_19653,N_19370,N_19380);
or U19654 (N_19654,N_19497,N_19394);
nand U19655 (N_19655,N_19398,N_19410);
nor U19656 (N_19656,N_19380,N_19494);
xor U19657 (N_19657,N_19375,N_19340);
nand U19658 (N_19658,N_19433,N_19334);
or U19659 (N_19659,N_19442,N_19255);
or U19660 (N_19660,N_19254,N_19275);
or U19661 (N_19661,N_19380,N_19373);
xnor U19662 (N_19662,N_19464,N_19270);
or U19663 (N_19663,N_19326,N_19369);
nand U19664 (N_19664,N_19279,N_19429);
and U19665 (N_19665,N_19406,N_19318);
xnor U19666 (N_19666,N_19401,N_19316);
and U19667 (N_19667,N_19372,N_19313);
or U19668 (N_19668,N_19323,N_19276);
xor U19669 (N_19669,N_19400,N_19396);
xor U19670 (N_19670,N_19269,N_19357);
and U19671 (N_19671,N_19435,N_19300);
or U19672 (N_19672,N_19346,N_19268);
xnor U19673 (N_19673,N_19335,N_19375);
xnor U19674 (N_19674,N_19334,N_19301);
nor U19675 (N_19675,N_19419,N_19319);
nor U19676 (N_19676,N_19320,N_19450);
xnor U19677 (N_19677,N_19477,N_19427);
and U19678 (N_19678,N_19466,N_19487);
or U19679 (N_19679,N_19337,N_19313);
and U19680 (N_19680,N_19276,N_19262);
nor U19681 (N_19681,N_19490,N_19265);
nand U19682 (N_19682,N_19365,N_19431);
xor U19683 (N_19683,N_19412,N_19309);
nand U19684 (N_19684,N_19408,N_19291);
and U19685 (N_19685,N_19492,N_19320);
xor U19686 (N_19686,N_19485,N_19423);
and U19687 (N_19687,N_19390,N_19406);
xor U19688 (N_19688,N_19385,N_19344);
nand U19689 (N_19689,N_19431,N_19283);
xor U19690 (N_19690,N_19367,N_19435);
xnor U19691 (N_19691,N_19266,N_19275);
or U19692 (N_19692,N_19391,N_19260);
xor U19693 (N_19693,N_19489,N_19380);
or U19694 (N_19694,N_19322,N_19296);
nor U19695 (N_19695,N_19252,N_19387);
nand U19696 (N_19696,N_19385,N_19264);
and U19697 (N_19697,N_19491,N_19408);
xor U19698 (N_19698,N_19366,N_19455);
and U19699 (N_19699,N_19437,N_19380);
nor U19700 (N_19700,N_19332,N_19273);
nand U19701 (N_19701,N_19317,N_19281);
or U19702 (N_19702,N_19394,N_19340);
xor U19703 (N_19703,N_19427,N_19333);
or U19704 (N_19704,N_19310,N_19474);
and U19705 (N_19705,N_19394,N_19480);
nor U19706 (N_19706,N_19330,N_19321);
nor U19707 (N_19707,N_19263,N_19471);
nand U19708 (N_19708,N_19414,N_19292);
xnor U19709 (N_19709,N_19269,N_19290);
nand U19710 (N_19710,N_19466,N_19251);
or U19711 (N_19711,N_19322,N_19476);
or U19712 (N_19712,N_19282,N_19496);
nor U19713 (N_19713,N_19373,N_19329);
nand U19714 (N_19714,N_19364,N_19405);
or U19715 (N_19715,N_19453,N_19300);
xor U19716 (N_19716,N_19489,N_19355);
xor U19717 (N_19717,N_19394,N_19265);
nand U19718 (N_19718,N_19384,N_19298);
xnor U19719 (N_19719,N_19306,N_19413);
or U19720 (N_19720,N_19408,N_19323);
nor U19721 (N_19721,N_19444,N_19370);
and U19722 (N_19722,N_19407,N_19380);
xnor U19723 (N_19723,N_19498,N_19380);
and U19724 (N_19724,N_19483,N_19363);
nor U19725 (N_19725,N_19314,N_19338);
nand U19726 (N_19726,N_19297,N_19498);
nor U19727 (N_19727,N_19417,N_19422);
nand U19728 (N_19728,N_19382,N_19492);
or U19729 (N_19729,N_19459,N_19434);
nor U19730 (N_19730,N_19263,N_19466);
nor U19731 (N_19731,N_19450,N_19379);
or U19732 (N_19732,N_19253,N_19450);
or U19733 (N_19733,N_19261,N_19353);
and U19734 (N_19734,N_19432,N_19279);
nand U19735 (N_19735,N_19420,N_19382);
and U19736 (N_19736,N_19455,N_19266);
nand U19737 (N_19737,N_19398,N_19327);
xnor U19738 (N_19738,N_19341,N_19330);
nor U19739 (N_19739,N_19282,N_19250);
and U19740 (N_19740,N_19305,N_19378);
or U19741 (N_19741,N_19297,N_19490);
nor U19742 (N_19742,N_19439,N_19280);
nor U19743 (N_19743,N_19338,N_19402);
nand U19744 (N_19744,N_19369,N_19365);
xor U19745 (N_19745,N_19344,N_19471);
nor U19746 (N_19746,N_19411,N_19405);
or U19747 (N_19747,N_19411,N_19430);
nand U19748 (N_19748,N_19316,N_19311);
or U19749 (N_19749,N_19316,N_19298);
nor U19750 (N_19750,N_19602,N_19500);
nor U19751 (N_19751,N_19621,N_19657);
xor U19752 (N_19752,N_19576,N_19641);
and U19753 (N_19753,N_19510,N_19543);
xor U19754 (N_19754,N_19566,N_19716);
nor U19755 (N_19755,N_19652,N_19741);
nor U19756 (N_19756,N_19549,N_19683);
and U19757 (N_19757,N_19724,N_19646);
or U19758 (N_19758,N_19742,N_19611);
and U19759 (N_19759,N_19540,N_19670);
nor U19760 (N_19760,N_19586,N_19572);
nand U19761 (N_19761,N_19718,N_19582);
or U19762 (N_19762,N_19589,N_19673);
nand U19763 (N_19763,N_19653,N_19517);
xnor U19764 (N_19764,N_19666,N_19710);
nand U19765 (N_19765,N_19520,N_19608);
nand U19766 (N_19766,N_19717,N_19681);
and U19767 (N_19767,N_19544,N_19743);
nor U19768 (N_19768,N_19633,N_19592);
nand U19769 (N_19769,N_19684,N_19746);
or U19770 (N_19770,N_19532,N_19584);
nand U19771 (N_19771,N_19747,N_19596);
or U19772 (N_19772,N_19606,N_19577);
nand U19773 (N_19773,N_19559,N_19732);
xor U19774 (N_19774,N_19739,N_19645);
and U19775 (N_19775,N_19610,N_19548);
nand U19776 (N_19776,N_19578,N_19658);
and U19777 (N_19777,N_19600,N_19601);
or U19778 (N_19778,N_19617,N_19526);
nand U19779 (N_19779,N_19697,N_19671);
nand U19780 (N_19780,N_19706,N_19662);
and U19781 (N_19781,N_19635,N_19689);
and U19782 (N_19782,N_19649,N_19636);
and U19783 (N_19783,N_19714,N_19708);
or U19784 (N_19784,N_19682,N_19539);
nand U19785 (N_19785,N_19723,N_19531);
nand U19786 (N_19786,N_19622,N_19693);
or U19787 (N_19787,N_19555,N_19504);
and U19788 (N_19788,N_19660,N_19628);
nand U19789 (N_19789,N_19607,N_19525);
nor U19790 (N_19790,N_19749,N_19744);
nand U19791 (N_19791,N_19687,N_19748);
xor U19792 (N_19792,N_19736,N_19677);
xor U19793 (N_19793,N_19712,N_19588);
nand U19794 (N_19794,N_19557,N_19629);
nor U19795 (N_19795,N_19725,N_19574);
xor U19796 (N_19796,N_19581,N_19734);
xnor U19797 (N_19797,N_19614,N_19560);
nor U19798 (N_19798,N_19599,N_19516);
nand U19799 (N_19799,N_19533,N_19536);
xor U19800 (N_19800,N_19616,N_19575);
nand U19801 (N_19801,N_19542,N_19508);
and U19802 (N_19802,N_19678,N_19650);
xor U19803 (N_19803,N_19627,N_19685);
nor U19804 (N_19804,N_19514,N_19691);
or U19805 (N_19805,N_19707,N_19654);
and U19806 (N_19806,N_19709,N_19669);
nand U19807 (N_19807,N_19583,N_19623);
and U19808 (N_19808,N_19570,N_19625);
and U19809 (N_19809,N_19643,N_19558);
and U19810 (N_19810,N_19647,N_19580);
nor U19811 (N_19811,N_19603,N_19651);
xor U19812 (N_19812,N_19521,N_19630);
or U19813 (N_19813,N_19637,N_19719);
and U19814 (N_19814,N_19524,N_19711);
and U19815 (N_19815,N_19529,N_19509);
or U19816 (N_19816,N_19728,N_19605);
xnor U19817 (N_19817,N_19585,N_19661);
nor U19818 (N_19818,N_19676,N_19597);
xor U19819 (N_19819,N_19726,N_19665);
nand U19820 (N_19820,N_19615,N_19702);
nand U19821 (N_19821,N_19594,N_19642);
nor U19822 (N_19822,N_19561,N_19668);
nor U19823 (N_19823,N_19730,N_19735);
and U19824 (N_19824,N_19619,N_19530);
nand U19825 (N_19825,N_19639,N_19527);
or U19826 (N_19826,N_19612,N_19618);
nor U19827 (N_19827,N_19656,N_19569);
xnor U19828 (N_19828,N_19688,N_19675);
xnor U19829 (N_19829,N_19648,N_19631);
nor U19830 (N_19830,N_19513,N_19563);
nor U19831 (N_19831,N_19545,N_19564);
and U19832 (N_19832,N_19694,N_19664);
or U19833 (N_19833,N_19733,N_19727);
xor U19834 (N_19834,N_19528,N_19640);
nand U19835 (N_19835,N_19745,N_19565);
and U19836 (N_19836,N_19550,N_19655);
xnor U19837 (N_19837,N_19505,N_19512);
nor U19838 (N_19838,N_19591,N_19595);
or U19839 (N_19839,N_19534,N_19626);
nand U19840 (N_19840,N_19729,N_19511);
nand U19841 (N_19841,N_19695,N_19674);
nand U19842 (N_19842,N_19679,N_19554);
or U19843 (N_19843,N_19552,N_19690);
or U19844 (N_19844,N_19551,N_19553);
or U19845 (N_19845,N_19568,N_19541);
nand U19846 (N_19846,N_19522,N_19535);
nand U19847 (N_19847,N_19537,N_19686);
or U19848 (N_19848,N_19634,N_19713);
or U19849 (N_19849,N_19672,N_19507);
nor U19850 (N_19850,N_19556,N_19562);
and U19851 (N_19851,N_19523,N_19644);
or U19852 (N_19852,N_19579,N_19738);
nand U19853 (N_19853,N_19547,N_19659);
or U19854 (N_19854,N_19519,N_19609);
and U19855 (N_19855,N_19613,N_19604);
nor U19856 (N_19856,N_19692,N_19680);
nor U19857 (N_19857,N_19703,N_19620);
or U19858 (N_19858,N_19667,N_19632);
and U19859 (N_19859,N_19546,N_19701);
and U19860 (N_19860,N_19699,N_19704);
nand U19861 (N_19861,N_19502,N_19700);
xnor U19862 (N_19862,N_19737,N_19705);
xor U19863 (N_19863,N_19721,N_19624);
nand U19864 (N_19864,N_19698,N_19722);
nor U19865 (N_19865,N_19567,N_19503);
or U19866 (N_19866,N_19518,N_19590);
xnor U19867 (N_19867,N_19593,N_19501);
xor U19868 (N_19868,N_19696,N_19598);
nor U19869 (N_19869,N_19506,N_19538);
xnor U19870 (N_19870,N_19731,N_19740);
and U19871 (N_19871,N_19663,N_19720);
nor U19872 (N_19872,N_19573,N_19587);
nand U19873 (N_19873,N_19715,N_19515);
xnor U19874 (N_19874,N_19571,N_19638);
nand U19875 (N_19875,N_19716,N_19541);
and U19876 (N_19876,N_19734,N_19709);
nand U19877 (N_19877,N_19746,N_19590);
nand U19878 (N_19878,N_19741,N_19532);
or U19879 (N_19879,N_19576,N_19606);
nor U19880 (N_19880,N_19506,N_19743);
nor U19881 (N_19881,N_19584,N_19602);
nor U19882 (N_19882,N_19594,N_19661);
and U19883 (N_19883,N_19737,N_19542);
and U19884 (N_19884,N_19655,N_19645);
or U19885 (N_19885,N_19738,N_19706);
xor U19886 (N_19886,N_19721,N_19636);
and U19887 (N_19887,N_19619,N_19521);
nor U19888 (N_19888,N_19595,N_19569);
nor U19889 (N_19889,N_19717,N_19737);
nor U19890 (N_19890,N_19582,N_19528);
nand U19891 (N_19891,N_19659,N_19520);
nand U19892 (N_19892,N_19573,N_19678);
nand U19893 (N_19893,N_19710,N_19662);
and U19894 (N_19894,N_19689,N_19575);
nor U19895 (N_19895,N_19673,N_19713);
xor U19896 (N_19896,N_19527,N_19644);
nor U19897 (N_19897,N_19589,N_19693);
or U19898 (N_19898,N_19721,N_19618);
nand U19899 (N_19899,N_19570,N_19745);
xnor U19900 (N_19900,N_19599,N_19730);
nor U19901 (N_19901,N_19517,N_19625);
nand U19902 (N_19902,N_19613,N_19616);
xor U19903 (N_19903,N_19592,N_19642);
xor U19904 (N_19904,N_19554,N_19577);
and U19905 (N_19905,N_19522,N_19546);
and U19906 (N_19906,N_19536,N_19678);
xor U19907 (N_19907,N_19632,N_19638);
and U19908 (N_19908,N_19621,N_19522);
nand U19909 (N_19909,N_19661,N_19544);
nand U19910 (N_19910,N_19739,N_19747);
or U19911 (N_19911,N_19529,N_19566);
nand U19912 (N_19912,N_19650,N_19664);
and U19913 (N_19913,N_19630,N_19532);
xnor U19914 (N_19914,N_19694,N_19593);
xnor U19915 (N_19915,N_19746,N_19730);
nand U19916 (N_19916,N_19710,N_19530);
or U19917 (N_19917,N_19548,N_19510);
xnor U19918 (N_19918,N_19539,N_19583);
or U19919 (N_19919,N_19674,N_19722);
nand U19920 (N_19920,N_19581,N_19536);
or U19921 (N_19921,N_19738,N_19675);
and U19922 (N_19922,N_19543,N_19735);
nand U19923 (N_19923,N_19634,N_19686);
or U19924 (N_19924,N_19595,N_19662);
xnor U19925 (N_19925,N_19696,N_19596);
xnor U19926 (N_19926,N_19687,N_19511);
or U19927 (N_19927,N_19548,N_19581);
nand U19928 (N_19928,N_19549,N_19559);
nand U19929 (N_19929,N_19686,N_19714);
nand U19930 (N_19930,N_19668,N_19647);
and U19931 (N_19931,N_19570,N_19635);
or U19932 (N_19932,N_19584,N_19670);
nor U19933 (N_19933,N_19595,N_19578);
and U19934 (N_19934,N_19617,N_19632);
xor U19935 (N_19935,N_19506,N_19574);
or U19936 (N_19936,N_19678,N_19521);
nor U19937 (N_19937,N_19733,N_19528);
or U19938 (N_19938,N_19666,N_19558);
nor U19939 (N_19939,N_19592,N_19503);
nand U19940 (N_19940,N_19634,N_19653);
and U19941 (N_19941,N_19730,N_19524);
nor U19942 (N_19942,N_19648,N_19597);
nand U19943 (N_19943,N_19532,N_19556);
xnor U19944 (N_19944,N_19663,N_19512);
nand U19945 (N_19945,N_19629,N_19611);
nand U19946 (N_19946,N_19748,N_19564);
nand U19947 (N_19947,N_19670,N_19664);
nand U19948 (N_19948,N_19742,N_19609);
and U19949 (N_19949,N_19606,N_19637);
and U19950 (N_19950,N_19589,N_19681);
and U19951 (N_19951,N_19589,N_19536);
or U19952 (N_19952,N_19535,N_19576);
or U19953 (N_19953,N_19533,N_19659);
nor U19954 (N_19954,N_19571,N_19597);
nor U19955 (N_19955,N_19543,N_19583);
nand U19956 (N_19956,N_19671,N_19603);
or U19957 (N_19957,N_19582,N_19714);
and U19958 (N_19958,N_19594,N_19588);
or U19959 (N_19959,N_19703,N_19625);
xnor U19960 (N_19960,N_19725,N_19693);
and U19961 (N_19961,N_19588,N_19668);
nand U19962 (N_19962,N_19694,N_19610);
nand U19963 (N_19963,N_19733,N_19556);
nor U19964 (N_19964,N_19679,N_19718);
nand U19965 (N_19965,N_19510,N_19732);
or U19966 (N_19966,N_19716,N_19565);
and U19967 (N_19967,N_19570,N_19528);
nor U19968 (N_19968,N_19696,N_19708);
nand U19969 (N_19969,N_19573,N_19534);
or U19970 (N_19970,N_19629,N_19549);
nor U19971 (N_19971,N_19617,N_19514);
nor U19972 (N_19972,N_19686,N_19549);
and U19973 (N_19973,N_19713,N_19675);
nor U19974 (N_19974,N_19514,N_19650);
and U19975 (N_19975,N_19743,N_19595);
nand U19976 (N_19976,N_19545,N_19727);
xor U19977 (N_19977,N_19724,N_19743);
nand U19978 (N_19978,N_19721,N_19620);
nor U19979 (N_19979,N_19660,N_19676);
nor U19980 (N_19980,N_19715,N_19736);
xnor U19981 (N_19981,N_19704,N_19707);
or U19982 (N_19982,N_19731,N_19595);
or U19983 (N_19983,N_19640,N_19564);
nand U19984 (N_19984,N_19589,N_19714);
nand U19985 (N_19985,N_19645,N_19541);
and U19986 (N_19986,N_19728,N_19714);
and U19987 (N_19987,N_19598,N_19566);
and U19988 (N_19988,N_19678,N_19630);
or U19989 (N_19989,N_19639,N_19685);
nand U19990 (N_19990,N_19647,N_19621);
nor U19991 (N_19991,N_19593,N_19542);
and U19992 (N_19992,N_19694,N_19577);
and U19993 (N_19993,N_19572,N_19722);
nor U19994 (N_19994,N_19597,N_19513);
xnor U19995 (N_19995,N_19625,N_19636);
or U19996 (N_19996,N_19555,N_19598);
nor U19997 (N_19997,N_19645,N_19708);
or U19998 (N_19998,N_19550,N_19623);
nand U19999 (N_19999,N_19663,N_19574);
or UO_0 (O_0,N_19796,N_19820);
nor UO_1 (O_1,N_19899,N_19805);
nor UO_2 (O_2,N_19926,N_19879);
or UO_3 (O_3,N_19932,N_19993);
xnor UO_4 (O_4,N_19983,N_19843);
and UO_5 (O_5,N_19929,N_19982);
nor UO_6 (O_6,N_19827,N_19989);
xor UO_7 (O_7,N_19845,N_19871);
nor UO_8 (O_8,N_19958,N_19876);
or UO_9 (O_9,N_19868,N_19838);
nor UO_10 (O_10,N_19927,N_19831);
xnor UO_11 (O_11,N_19863,N_19857);
or UO_12 (O_12,N_19758,N_19782);
xor UO_13 (O_13,N_19772,N_19974);
nor UO_14 (O_14,N_19877,N_19991);
and UO_15 (O_15,N_19948,N_19840);
nor UO_16 (O_16,N_19860,N_19901);
and UO_17 (O_17,N_19751,N_19808);
nor UO_18 (O_18,N_19769,N_19768);
nor UO_19 (O_19,N_19903,N_19781);
nand UO_20 (O_20,N_19874,N_19855);
nor UO_21 (O_21,N_19846,N_19887);
xor UO_22 (O_22,N_19944,N_19867);
nand UO_23 (O_23,N_19955,N_19767);
nand UO_24 (O_24,N_19854,N_19849);
and UO_25 (O_25,N_19859,N_19888);
and UO_26 (O_26,N_19971,N_19825);
nor UO_27 (O_27,N_19783,N_19806);
and UO_28 (O_28,N_19788,N_19986);
nand UO_29 (O_29,N_19801,N_19980);
nor UO_30 (O_30,N_19947,N_19880);
nor UO_31 (O_31,N_19940,N_19978);
or UO_32 (O_32,N_19878,N_19902);
and UO_33 (O_33,N_19951,N_19814);
and UO_34 (O_34,N_19913,N_19937);
or UO_35 (O_35,N_19786,N_19842);
nor UO_36 (O_36,N_19952,N_19870);
or UO_37 (O_37,N_19897,N_19984);
or UO_38 (O_38,N_19985,N_19754);
or UO_39 (O_39,N_19925,N_19856);
and UO_40 (O_40,N_19914,N_19996);
nand UO_41 (O_41,N_19823,N_19976);
and UO_42 (O_42,N_19818,N_19904);
and UO_43 (O_43,N_19852,N_19968);
nor UO_44 (O_44,N_19793,N_19905);
or UO_45 (O_45,N_19803,N_19775);
and UO_46 (O_46,N_19909,N_19858);
nor UO_47 (O_47,N_19963,N_19804);
and UO_48 (O_48,N_19922,N_19777);
nor UO_49 (O_49,N_19773,N_19875);
and UO_50 (O_50,N_19864,N_19938);
xor UO_51 (O_51,N_19988,N_19764);
and UO_52 (O_52,N_19995,N_19946);
nor UO_53 (O_53,N_19894,N_19873);
nand UO_54 (O_54,N_19953,N_19795);
and UO_55 (O_55,N_19815,N_19882);
and UO_56 (O_56,N_19826,N_19872);
nor UO_57 (O_57,N_19760,N_19979);
or UO_58 (O_58,N_19969,N_19931);
nand UO_59 (O_59,N_19966,N_19930);
and UO_60 (O_60,N_19906,N_19889);
nand UO_61 (O_61,N_19822,N_19778);
xor UO_62 (O_62,N_19753,N_19812);
and UO_63 (O_63,N_19780,N_19981);
nand UO_64 (O_64,N_19841,N_19918);
nor UO_65 (O_65,N_19817,N_19798);
nor UO_66 (O_66,N_19844,N_19766);
nor UO_67 (O_67,N_19911,N_19816);
nor UO_68 (O_68,N_19908,N_19920);
xor UO_69 (O_69,N_19945,N_19848);
and UO_70 (O_70,N_19835,N_19779);
nand UO_71 (O_71,N_19802,N_19910);
xnor UO_72 (O_72,N_19790,N_19886);
nor UO_73 (O_73,N_19994,N_19975);
nor UO_74 (O_74,N_19851,N_19936);
xor UO_75 (O_75,N_19861,N_19896);
or UO_76 (O_76,N_19830,N_19791);
xnor UO_77 (O_77,N_19949,N_19761);
xnor UO_78 (O_78,N_19999,N_19885);
and UO_79 (O_79,N_19939,N_19884);
or UO_80 (O_80,N_19977,N_19765);
xnor UO_81 (O_81,N_19869,N_19784);
nand UO_82 (O_82,N_19912,N_19972);
or UO_83 (O_83,N_19960,N_19832);
and UO_84 (O_84,N_19891,N_19924);
nor UO_85 (O_85,N_19964,N_19759);
xnor UO_86 (O_86,N_19935,N_19789);
xnor UO_87 (O_87,N_19809,N_19755);
nor UO_88 (O_88,N_19900,N_19916);
or UO_89 (O_89,N_19829,N_19792);
xor UO_90 (O_90,N_19828,N_19839);
or UO_91 (O_91,N_19883,N_19810);
xor UO_92 (O_92,N_19813,N_19917);
or UO_93 (O_93,N_19890,N_19762);
xnor UO_94 (O_94,N_19973,N_19824);
nor UO_95 (O_95,N_19752,N_19770);
xnor UO_96 (O_96,N_19965,N_19915);
nand UO_97 (O_97,N_19800,N_19797);
nand UO_98 (O_98,N_19756,N_19954);
and UO_99 (O_99,N_19990,N_19970);
xnor UO_100 (O_100,N_19962,N_19771);
or UO_101 (O_101,N_19811,N_19956);
xor UO_102 (O_102,N_19998,N_19794);
nand UO_103 (O_103,N_19850,N_19893);
xor UO_104 (O_104,N_19837,N_19865);
and UO_105 (O_105,N_19967,N_19834);
nor UO_106 (O_106,N_19959,N_19942);
and UO_107 (O_107,N_19933,N_19774);
or UO_108 (O_108,N_19957,N_19821);
xor UO_109 (O_109,N_19866,N_19750);
or UO_110 (O_110,N_19921,N_19776);
xor UO_111 (O_111,N_19847,N_19943);
xnor UO_112 (O_112,N_19895,N_19941);
or UO_113 (O_113,N_19950,N_19907);
nand UO_114 (O_114,N_19836,N_19853);
nand UO_115 (O_115,N_19928,N_19881);
or UO_116 (O_116,N_19819,N_19987);
nor UO_117 (O_117,N_19757,N_19997);
xnor UO_118 (O_118,N_19898,N_19862);
nor UO_119 (O_119,N_19892,N_19992);
xnor UO_120 (O_120,N_19919,N_19934);
xor UO_121 (O_121,N_19785,N_19833);
xnor UO_122 (O_122,N_19923,N_19961);
xor UO_123 (O_123,N_19807,N_19787);
or UO_124 (O_124,N_19763,N_19799);
or UO_125 (O_125,N_19938,N_19861);
and UO_126 (O_126,N_19830,N_19942);
or UO_127 (O_127,N_19846,N_19860);
or UO_128 (O_128,N_19762,N_19785);
xnor UO_129 (O_129,N_19829,N_19849);
or UO_130 (O_130,N_19933,N_19810);
and UO_131 (O_131,N_19970,N_19946);
xor UO_132 (O_132,N_19941,N_19883);
or UO_133 (O_133,N_19931,N_19983);
xor UO_134 (O_134,N_19927,N_19771);
nor UO_135 (O_135,N_19909,N_19826);
nand UO_136 (O_136,N_19786,N_19799);
or UO_137 (O_137,N_19821,N_19761);
and UO_138 (O_138,N_19993,N_19972);
nand UO_139 (O_139,N_19990,N_19772);
or UO_140 (O_140,N_19994,N_19800);
and UO_141 (O_141,N_19891,N_19970);
and UO_142 (O_142,N_19875,N_19948);
nand UO_143 (O_143,N_19964,N_19893);
or UO_144 (O_144,N_19802,N_19813);
nor UO_145 (O_145,N_19981,N_19893);
nand UO_146 (O_146,N_19899,N_19777);
nor UO_147 (O_147,N_19827,N_19990);
and UO_148 (O_148,N_19968,N_19812);
nor UO_149 (O_149,N_19920,N_19909);
or UO_150 (O_150,N_19991,N_19811);
or UO_151 (O_151,N_19924,N_19983);
or UO_152 (O_152,N_19887,N_19862);
or UO_153 (O_153,N_19932,N_19764);
or UO_154 (O_154,N_19987,N_19975);
nor UO_155 (O_155,N_19935,N_19922);
nand UO_156 (O_156,N_19914,N_19793);
and UO_157 (O_157,N_19766,N_19765);
or UO_158 (O_158,N_19801,N_19963);
and UO_159 (O_159,N_19915,N_19894);
or UO_160 (O_160,N_19815,N_19785);
nor UO_161 (O_161,N_19854,N_19994);
nor UO_162 (O_162,N_19898,N_19793);
or UO_163 (O_163,N_19927,N_19900);
or UO_164 (O_164,N_19807,N_19960);
xor UO_165 (O_165,N_19912,N_19833);
xor UO_166 (O_166,N_19768,N_19807);
and UO_167 (O_167,N_19943,N_19922);
and UO_168 (O_168,N_19995,N_19765);
xnor UO_169 (O_169,N_19860,N_19981);
nand UO_170 (O_170,N_19866,N_19844);
nor UO_171 (O_171,N_19998,N_19966);
and UO_172 (O_172,N_19971,N_19972);
xor UO_173 (O_173,N_19936,N_19937);
or UO_174 (O_174,N_19759,N_19820);
nor UO_175 (O_175,N_19773,N_19938);
nand UO_176 (O_176,N_19936,N_19799);
and UO_177 (O_177,N_19954,N_19818);
xnor UO_178 (O_178,N_19889,N_19935);
nand UO_179 (O_179,N_19795,N_19779);
nand UO_180 (O_180,N_19850,N_19904);
and UO_181 (O_181,N_19969,N_19874);
nand UO_182 (O_182,N_19766,N_19815);
or UO_183 (O_183,N_19973,N_19814);
nor UO_184 (O_184,N_19904,N_19906);
and UO_185 (O_185,N_19802,N_19769);
nor UO_186 (O_186,N_19751,N_19912);
xor UO_187 (O_187,N_19906,N_19834);
or UO_188 (O_188,N_19991,N_19819);
nand UO_189 (O_189,N_19994,N_19776);
nand UO_190 (O_190,N_19866,N_19885);
nand UO_191 (O_191,N_19888,N_19842);
nand UO_192 (O_192,N_19751,N_19815);
nor UO_193 (O_193,N_19866,N_19937);
xor UO_194 (O_194,N_19822,N_19781);
or UO_195 (O_195,N_19866,N_19800);
or UO_196 (O_196,N_19812,N_19998);
and UO_197 (O_197,N_19919,N_19809);
nand UO_198 (O_198,N_19958,N_19989);
xnor UO_199 (O_199,N_19825,N_19897);
xnor UO_200 (O_200,N_19924,N_19908);
and UO_201 (O_201,N_19837,N_19886);
or UO_202 (O_202,N_19996,N_19802);
and UO_203 (O_203,N_19783,N_19993);
and UO_204 (O_204,N_19916,N_19753);
nand UO_205 (O_205,N_19965,N_19993);
and UO_206 (O_206,N_19899,N_19966);
nor UO_207 (O_207,N_19895,N_19814);
nor UO_208 (O_208,N_19756,N_19816);
nand UO_209 (O_209,N_19996,N_19907);
or UO_210 (O_210,N_19823,N_19931);
nand UO_211 (O_211,N_19954,N_19803);
or UO_212 (O_212,N_19811,N_19787);
nor UO_213 (O_213,N_19998,N_19789);
and UO_214 (O_214,N_19807,N_19876);
nor UO_215 (O_215,N_19963,N_19860);
nand UO_216 (O_216,N_19840,N_19933);
nand UO_217 (O_217,N_19866,N_19816);
nand UO_218 (O_218,N_19973,N_19916);
xor UO_219 (O_219,N_19945,N_19924);
or UO_220 (O_220,N_19989,N_19835);
nor UO_221 (O_221,N_19828,N_19788);
nor UO_222 (O_222,N_19886,N_19846);
nand UO_223 (O_223,N_19852,N_19792);
nor UO_224 (O_224,N_19948,N_19900);
xor UO_225 (O_225,N_19793,N_19868);
or UO_226 (O_226,N_19815,N_19966);
nor UO_227 (O_227,N_19984,N_19920);
or UO_228 (O_228,N_19982,N_19809);
and UO_229 (O_229,N_19850,N_19890);
xor UO_230 (O_230,N_19870,N_19822);
xnor UO_231 (O_231,N_19879,N_19822);
xor UO_232 (O_232,N_19953,N_19963);
xor UO_233 (O_233,N_19996,N_19878);
or UO_234 (O_234,N_19950,N_19777);
and UO_235 (O_235,N_19969,N_19850);
nand UO_236 (O_236,N_19763,N_19774);
and UO_237 (O_237,N_19801,N_19976);
or UO_238 (O_238,N_19780,N_19948);
or UO_239 (O_239,N_19837,N_19770);
xnor UO_240 (O_240,N_19987,N_19860);
nand UO_241 (O_241,N_19785,N_19782);
and UO_242 (O_242,N_19780,N_19976);
and UO_243 (O_243,N_19921,N_19822);
nand UO_244 (O_244,N_19928,N_19788);
and UO_245 (O_245,N_19791,N_19954);
or UO_246 (O_246,N_19927,N_19858);
nand UO_247 (O_247,N_19807,N_19990);
nand UO_248 (O_248,N_19954,N_19761);
and UO_249 (O_249,N_19880,N_19928);
nor UO_250 (O_250,N_19955,N_19878);
and UO_251 (O_251,N_19751,N_19983);
xor UO_252 (O_252,N_19936,N_19860);
or UO_253 (O_253,N_19773,N_19910);
and UO_254 (O_254,N_19803,N_19755);
nand UO_255 (O_255,N_19842,N_19913);
or UO_256 (O_256,N_19973,N_19988);
or UO_257 (O_257,N_19833,N_19975);
nand UO_258 (O_258,N_19770,N_19766);
and UO_259 (O_259,N_19930,N_19922);
xor UO_260 (O_260,N_19919,N_19821);
nor UO_261 (O_261,N_19970,N_19849);
and UO_262 (O_262,N_19896,N_19826);
xnor UO_263 (O_263,N_19969,N_19869);
or UO_264 (O_264,N_19954,N_19994);
nor UO_265 (O_265,N_19842,N_19874);
nor UO_266 (O_266,N_19814,N_19829);
nor UO_267 (O_267,N_19845,N_19982);
nand UO_268 (O_268,N_19867,N_19831);
xnor UO_269 (O_269,N_19917,N_19774);
and UO_270 (O_270,N_19905,N_19822);
nand UO_271 (O_271,N_19788,N_19791);
and UO_272 (O_272,N_19872,N_19774);
nand UO_273 (O_273,N_19818,N_19856);
xor UO_274 (O_274,N_19759,N_19919);
xnor UO_275 (O_275,N_19841,N_19995);
nor UO_276 (O_276,N_19751,N_19752);
nand UO_277 (O_277,N_19929,N_19973);
xnor UO_278 (O_278,N_19766,N_19953);
nor UO_279 (O_279,N_19922,N_19884);
or UO_280 (O_280,N_19890,N_19993);
nand UO_281 (O_281,N_19825,N_19837);
nand UO_282 (O_282,N_19987,N_19794);
xor UO_283 (O_283,N_19783,N_19812);
and UO_284 (O_284,N_19837,N_19814);
and UO_285 (O_285,N_19965,N_19891);
nand UO_286 (O_286,N_19872,N_19934);
nand UO_287 (O_287,N_19822,N_19825);
nand UO_288 (O_288,N_19792,N_19907);
nor UO_289 (O_289,N_19990,N_19836);
or UO_290 (O_290,N_19956,N_19826);
and UO_291 (O_291,N_19821,N_19966);
nor UO_292 (O_292,N_19969,N_19752);
nor UO_293 (O_293,N_19925,N_19794);
nand UO_294 (O_294,N_19759,N_19887);
xor UO_295 (O_295,N_19774,N_19980);
nor UO_296 (O_296,N_19956,N_19807);
nor UO_297 (O_297,N_19882,N_19961);
xor UO_298 (O_298,N_19854,N_19817);
and UO_299 (O_299,N_19872,N_19904);
xnor UO_300 (O_300,N_19854,N_19988);
or UO_301 (O_301,N_19820,N_19792);
nand UO_302 (O_302,N_19818,N_19966);
nand UO_303 (O_303,N_19940,N_19840);
or UO_304 (O_304,N_19807,N_19814);
xor UO_305 (O_305,N_19801,N_19894);
nor UO_306 (O_306,N_19988,N_19869);
nand UO_307 (O_307,N_19941,N_19843);
xor UO_308 (O_308,N_19844,N_19862);
and UO_309 (O_309,N_19929,N_19999);
nor UO_310 (O_310,N_19966,N_19921);
nor UO_311 (O_311,N_19873,N_19928);
nor UO_312 (O_312,N_19881,N_19837);
nand UO_313 (O_313,N_19979,N_19808);
nor UO_314 (O_314,N_19946,N_19969);
nand UO_315 (O_315,N_19912,N_19973);
xnor UO_316 (O_316,N_19854,N_19984);
or UO_317 (O_317,N_19793,N_19888);
xnor UO_318 (O_318,N_19897,N_19899);
and UO_319 (O_319,N_19953,N_19764);
nand UO_320 (O_320,N_19864,N_19774);
or UO_321 (O_321,N_19847,N_19879);
xor UO_322 (O_322,N_19828,N_19770);
and UO_323 (O_323,N_19815,N_19863);
or UO_324 (O_324,N_19864,N_19896);
nand UO_325 (O_325,N_19915,N_19762);
or UO_326 (O_326,N_19790,N_19808);
xnor UO_327 (O_327,N_19923,N_19975);
nand UO_328 (O_328,N_19862,N_19840);
and UO_329 (O_329,N_19939,N_19754);
nand UO_330 (O_330,N_19857,N_19938);
or UO_331 (O_331,N_19931,N_19910);
nor UO_332 (O_332,N_19754,N_19821);
nand UO_333 (O_333,N_19756,N_19834);
and UO_334 (O_334,N_19907,N_19963);
nand UO_335 (O_335,N_19976,N_19752);
nand UO_336 (O_336,N_19954,N_19844);
or UO_337 (O_337,N_19866,N_19932);
xnor UO_338 (O_338,N_19920,N_19813);
and UO_339 (O_339,N_19825,N_19934);
or UO_340 (O_340,N_19922,N_19872);
nand UO_341 (O_341,N_19988,N_19996);
and UO_342 (O_342,N_19945,N_19771);
xor UO_343 (O_343,N_19919,N_19927);
and UO_344 (O_344,N_19767,N_19856);
xnor UO_345 (O_345,N_19800,N_19830);
nand UO_346 (O_346,N_19777,N_19857);
or UO_347 (O_347,N_19775,N_19976);
nand UO_348 (O_348,N_19794,N_19922);
and UO_349 (O_349,N_19858,N_19976);
xor UO_350 (O_350,N_19948,N_19776);
xor UO_351 (O_351,N_19899,N_19770);
nand UO_352 (O_352,N_19841,N_19956);
or UO_353 (O_353,N_19786,N_19860);
and UO_354 (O_354,N_19991,N_19962);
or UO_355 (O_355,N_19974,N_19751);
xor UO_356 (O_356,N_19920,N_19874);
or UO_357 (O_357,N_19790,N_19891);
or UO_358 (O_358,N_19873,N_19870);
or UO_359 (O_359,N_19849,N_19813);
nand UO_360 (O_360,N_19758,N_19921);
xor UO_361 (O_361,N_19887,N_19850);
nor UO_362 (O_362,N_19979,N_19918);
or UO_363 (O_363,N_19770,N_19994);
nand UO_364 (O_364,N_19754,N_19970);
and UO_365 (O_365,N_19750,N_19765);
and UO_366 (O_366,N_19997,N_19874);
or UO_367 (O_367,N_19844,N_19926);
xor UO_368 (O_368,N_19797,N_19928);
nor UO_369 (O_369,N_19852,N_19837);
nand UO_370 (O_370,N_19984,N_19825);
xor UO_371 (O_371,N_19982,N_19817);
nor UO_372 (O_372,N_19820,N_19942);
nor UO_373 (O_373,N_19962,N_19826);
nand UO_374 (O_374,N_19831,N_19999);
nor UO_375 (O_375,N_19855,N_19987);
or UO_376 (O_376,N_19773,N_19876);
nor UO_377 (O_377,N_19893,N_19876);
nand UO_378 (O_378,N_19946,N_19832);
nor UO_379 (O_379,N_19773,N_19952);
and UO_380 (O_380,N_19944,N_19813);
nor UO_381 (O_381,N_19932,N_19803);
xnor UO_382 (O_382,N_19816,N_19951);
or UO_383 (O_383,N_19765,N_19787);
xor UO_384 (O_384,N_19800,N_19992);
and UO_385 (O_385,N_19861,N_19928);
nand UO_386 (O_386,N_19951,N_19893);
nand UO_387 (O_387,N_19945,N_19912);
or UO_388 (O_388,N_19823,N_19847);
or UO_389 (O_389,N_19866,N_19998);
or UO_390 (O_390,N_19927,N_19840);
nand UO_391 (O_391,N_19953,N_19865);
xor UO_392 (O_392,N_19828,N_19860);
or UO_393 (O_393,N_19891,N_19894);
and UO_394 (O_394,N_19778,N_19997);
and UO_395 (O_395,N_19977,N_19968);
or UO_396 (O_396,N_19873,N_19869);
nand UO_397 (O_397,N_19810,N_19977);
and UO_398 (O_398,N_19987,N_19828);
nand UO_399 (O_399,N_19828,N_19873);
and UO_400 (O_400,N_19944,N_19807);
or UO_401 (O_401,N_19922,N_19937);
nand UO_402 (O_402,N_19877,N_19861);
and UO_403 (O_403,N_19907,N_19868);
nand UO_404 (O_404,N_19800,N_19773);
or UO_405 (O_405,N_19929,N_19827);
nor UO_406 (O_406,N_19921,N_19963);
and UO_407 (O_407,N_19827,N_19818);
xnor UO_408 (O_408,N_19861,N_19859);
nor UO_409 (O_409,N_19974,N_19860);
nor UO_410 (O_410,N_19977,N_19821);
and UO_411 (O_411,N_19912,N_19819);
or UO_412 (O_412,N_19970,N_19903);
xnor UO_413 (O_413,N_19916,N_19825);
or UO_414 (O_414,N_19906,N_19888);
nor UO_415 (O_415,N_19765,N_19934);
and UO_416 (O_416,N_19770,N_19821);
nor UO_417 (O_417,N_19956,N_19857);
nor UO_418 (O_418,N_19850,N_19811);
and UO_419 (O_419,N_19902,N_19886);
and UO_420 (O_420,N_19861,N_19934);
nand UO_421 (O_421,N_19919,N_19956);
or UO_422 (O_422,N_19983,N_19839);
xor UO_423 (O_423,N_19861,N_19907);
nor UO_424 (O_424,N_19975,N_19790);
nand UO_425 (O_425,N_19826,N_19763);
or UO_426 (O_426,N_19888,N_19980);
xor UO_427 (O_427,N_19864,N_19832);
xor UO_428 (O_428,N_19764,N_19808);
or UO_429 (O_429,N_19920,N_19900);
xor UO_430 (O_430,N_19804,N_19990);
nand UO_431 (O_431,N_19858,N_19788);
and UO_432 (O_432,N_19980,N_19857);
xnor UO_433 (O_433,N_19839,N_19896);
or UO_434 (O_434,N_19836,N_19985);
nor UO_435 (O_435,N_19911,N_19815);
nand UO_436 (O_436,N_19926,N_19817);
and UO_437 (O_437,N_19976,N_19907);
nor UO_438 (O_438,N_19942,N_19780);
and UO_439 (O_439,N_19754,N_19770);
nor UO_440 (O_440,N_19904,N_19984);
xnor UO_441 (O_441,N_19849,N_19783);
nand UO_442 (O_442,N_19918,N_19904);
nand UO_443 (O_443,N_19924,N_19985);
xnor UO_444 (O_444,N_19933,N_19886);
xor UO_445 (O_445,N_19906,N_19978);
xnor UO_446 (O_446,N_19925,N_19979);
nand UO_447 (O_447,N_19794,N_19890);
and UO_448 (O_448,N_19801,N_19978);
nor UO_449 (O_449,N_19948,N_19764);
nand UO_450 (O_450,N_19784,N_19900);
and UO_451 (O_451,N_19998,N_19928);
or UO_452 (O_452,N_19838,N_19870);
and UO_453 (O_453,N_19953,N_19765);
xnor UO_454 (O_454,N_19936,N_19773);
or UO_455 (O_455,N_19962,N_19769);
or UO_456 (O_456,N_19902,N_19787);
nand UO_457 (O_457,N_19846,N_19840);
nand UO_458 (O_458,N_19903,N_19943);
and UO_459 (O_459,N_19923,N_19921);
xor UO_460 (O_460,N_19986,N_19912);
xnor UO_461 (O_461,N_19831,N_19770);
or UO_462 (O_462,N_19967,N_19781);
nand UO_463 (O_463,N_19990,N_19778);
or UO_464 (O_464,N_19884,N_19913);
nor UO_465 (O_465,N_19892,N_19764);
xnor UO_466 (O_466,N_19974,N_19915);
nor UO_467 (O_467,N_19891,N_19940);
and UO_468 (O_468,N_19757,N_19832);
and UO_469 (O_469,N_19812,N_19992);
nor UO_470 (O_470,N_19863,N_19904);
nor UO_471 (O_471,N_19991,N_19781);
nor UO_472 (O_472,N_19816,N_19918);
and UO_473 (O_473,N_19914,N_19837);
xor UO_474 (O_474,N_19816,N_19958);
nand UO_475 (O_475,N_19896,N_19851);
and UO_476 (O_476,N_19789,N_19756);
xor UO_477 (O_477,N_19807,N_19917);
or UO_478 (O_478,N_19904,N_19889);
or UO_479 (O_479,N_19789,N_19816);
nor UO_480 (O_480,N_19979,N_19784);
xnor UO_481 (O_481,N_19976,N_19888);
xor UO_482 (O_482,N_19983,N_19867);
nor UO_483 (O_483,N_19950,N_19762);
xor UO_484 (O_484,N_19950,N_19901);
nand UO_485 (O_485,N_19965,N_19880);
nand UO_486 (O_486,N_19814,N_19887);
and UO_487 (O_487,N_19896,N_19914);
nand UO_488 (O_488,N_19986,N_19899);
nor UO_489 (O_489,N_19890,N_19822);
or UO_490 (O_490,N_19938,N_19846);
nor UO_491 (O_491,N_19860,N_19954);
nand UO_492 (O_492,N_19993,N_19999);
xor UO_493 (O_493,N_19857,N_19992);
nor UO_494 (O_494,N_19903,N_19972);
xor UO_495 (O_495,N_19877,N_19754);
nand UO_496 (O_496,N_19796,N_19770);
nand UO_497 (O_497,N_19908,N_19876);
or UO_498 (O_498,N_19837,N_19797);
and UO_499 (O_499,N_19816,N_19977);
nand UO_500 (O_500,N_19869,N_19900);
or UO_501 (O_501,N_19927,N_19965);
nand UO_502 (O_502,N_19828,N_19951);
nor UO_503 (O_503,N_19988,N_19915);
or UO_504 (O_504,N_19825,N_19788);
or UO_505 (O_505,N_19784,N_19858);
and UO_506 (O_506,N_19967,N_19995);
nor UO_507 (O_507,N_19975,N_19988);
or UO_508 (O_508,N_19796,N_19862);
and UO_509 (O_509,N_19753,N_19804);
and UO_510 (O_510,N_19844,N_19988);
nand UO_511 (O_511,N_19946,N_19794);
nor UO_512 (O_512,N_19845,N_19969);
nand UO_513 (O_513,N_19936,N_19792);
xnor UO_514 (O_514,N_19787,N_19763);
and UO_515 (O_515,N_19763,N_19904);
and UO_516 (O_516,N_19799,N_19769);
nor UO_517 (O_517,N_19951,N_19993);
nor UO_518 (O_518,N_19835,N_19829);
or UO_519 (O_519,N_19947,N_19936);
xnor UO_520 (O_520,N_19830,N_19893);
nor UO_521 (O_521,N_19794,N_19938);
or UO_522 (O_522,N_19797,N_19938);
and UO_523 (O_523,N_19873,N_19830);
nor UO_524 (O_524,N_19925,N_19824);
nand UO_525 (O_525,N_19867,N_19896);
or UO_526 (O_526,N_19944,N_19825);
nor UO_527 (O_527,N_19908,N_19859);
nand UO_528 (O_528,N_19909,N_19798);
nor UO_529 (O_529,N_19890,N_19796);
nor UO_530 (O_530,N_19753,N_19788);
nand UO_531 (O_531,N_19831,N_19905);
and UO_532 (O_532,N_19829,N_19991);
nor UO_533 (O_533,N_19789,N_19918);
nor UO_534 (O_534,N_19954,N_19813);
and UO_535 (O_535,N_19778,N_19875);
nor UO_536 (O_536,N_19976,N_19939);
nand UO_537 (O_537,N_19821,N_19759);
and UO_538 (O_538,N_19759,N_19784);
xor UO_539 (O_539,N_19800,N_19989);
nand UO_540 (O_540,N_19950,N_19944);
nand UO_541 (O_541,N_19926,N_19988);
nor UO_542 (O_542,N_19806,N_19840);
or UO_543 (O_543,N_19775,N_19998);
nand UO_544 (O_544,N_19863,N_19833);
nor UO_545 (O_545,N_19862,N_19888);
nand UO_546 (O_546,N_19788,N_19809);
and UO_547 (O_547,N_19993,N_19780);
and UO_548 (O_548,N_19880,N_19842);
and UO_549 (O_549,N_19971,N_19989);
and UO_550 (O_550,N_19758,N_19966);
and UO_551 (O_551,N_19885,N_19759);
and UO_552 (O_552,N_19942,N_19761);
xnor UO_553 (O_553,N_19995,N_19977);
xor UO_554 (O_554,N_19961,N_19804);
nand UO_555 (O_555,N_19910,N_19864);
xor UO_556 (O_556,N_19821,N_19948);
nor UO_557 (O_557,N_19959,N_19866);
nand UO_558 (O_558,N_19859,N_19959);
or UO_559 (O_559,N_19862,N_19911);
and UO_560 (O_560,N_19849,N_19947);
nand UO_561 (O_561,N_19858,N_19757);
xnor UO_562 (O_562,N_19936,N_19954);
and UO_563 (O_563,N_19884,N_19933);
xnor UO_564 (O_564,N_19769,N_19973);
or UO_565 (O_565,N_19755,N_19896);
xnor UO_566 (O_566,N_19893,N_19987);
xnor UO_567 (O_567,N_19805,N_19866);
nand UO_568 (O_568,N_19762,N_19769);
nand UO_569 (O_569,N_19814,N_19828);
nor UO_570 (O_570,N_19962,N_19915);
or UO_571 (O_571,N_19896,N_19792);
nand UO_572 (O_572,N_19827,N_19938);
nand UO_573 (O_573,N_19825,N_19785);
and UO_574 (O_574,N_19760,N_19942);
nand UO_575 (O_575,N_19939,N_19964);
and UO_576 (O_576,N_19979,N_19751);
xor UO_577 (O_577,N_19985,N_19891);
or UO_578 (O_578,N_19798,N_19803);
and UO_579 (O_579,N_19855,N_19835);
nand UO_580 (O_580,N_19873,N_19851);
and UO_581 (O_581,N_19981,N_19786);
and UO_582 (O_582,N_19809,N_19878);
nor UO_583 (O_583,N_19858,N_19893);
or UO_584 (O_584,N_19912,N_19780);
nor UO_585 (O_585,N_19815,N_19959);
and UO_586 (O_586,N_19986,N_19874);
or UO_587 (O_587,N_19777,N_19945);
and UO_588 (O_588,N_19955,N_19903);
nand UO_589 (O_589,N_19775,N_19782);
nor UO_590 (O_590,N_19879,N_19963);
xor UO_591 (O_591,N_19766,N_19868);
or UO_592 (O_592,N_19994,N_19825);
xor UO_593 (O_593,N_19773,N_19750);
nor UO_594 (O_594,N_19860,N_19857);
nor UO_595 (O_595,N_19972,N_19805);
xor UO_596 (O_596,N_19774,N_19924);
nor UO_597 (O_597,N_19834,N_19860);
and UO_598 (O_598,N_19864,N_19811);
or UO_599 (O_599,N_19814,N_19802);
nand UO_600 (O_600,N_19950,N_19972);
nor UO_601 (O_601,N_19802,N_19963);
and UO_602 (O_602,N_19774,N_19970);
and UO_603 (O_603,N_19842,N_19970);
or UO_604 (O_604,N_19950,N_19808);
and UO_605 (O_605,N_19894,N_19933);
or UO_606 (O_606,N_19832,N_19999);
nor UO_607 (O_607,N_19976,N_19783);
and UO_608 (O_608,N_19982,N_19844);
nand UO_609 (O_609,N_19989,N_19970);
or UO_610 (O_610,N_19783,N_19793);
or UO_611 (O_611,N_19919,N_19828);
and UO_612 (O_612,N_19855,N_19793);
or UO_613 (O_613,N_19945,N_19990);
nand UO_614 (O_614,N_19871,N_19922);
xor UO_615 (O_615,N_19823,N_19846);
xor UO_616 (O_616,N_19956,N_19920);
nor UO_617 (O_617,N_19926,N_19782);
nand UO_618 (O_618,N_19955,N_19766);
xnor UO_619 (O_619,N_19989,N_19775);
nand UO_620 (O_620,N_19896,N_19984);
or UO_621 (O_621,N_19992,N_19843);
and UO_622 (O_622,N_19953,N_19904);
nand UO_623 (O_623,N_19833,N_19927);
nor UO_624 (O_624,N_19818,N_19795);
and UO_625 (O_625,N_19910,N_19942);
xnor UO_626 (O_626,N_19761,N_19802);
or UO_627 (O_627,N_19951,N_19952);
and UO_628 (O_628,N_19859,N_19800);
nor UO_629 (O_629,N_19754,N_19986);
nor UO_630 (O_630,N_19750,N_19923);
and UO_631 (O_631,N_19779,N_19917);
nor UO_632 (O_632,N_19970,N_19911);
or UO_633 (O_633,N_19903,N_19976);
nor UO_634 (O_634,N_19815,N_19874);
or UO_635 (O_635,N_19898,N_19968);
nand UO_636 (O_636,N_19768,N_19880);
or UO_637 (O_637,N_19982,N_19767);
xor UO_638 (O_638,N_19810,N_19781);
or UO_639 (O_639,N_19828,N_19892);
nand UO_640 (O_640,N_19838,N_19975);
xnor UO_641 (O_641,N_19861,N_19770);
and UO_642 (O_642,N_19965,N_19863);
and UO_643 (O_643,N_19945,N_19811);
and UO_644 (O_644,N_19831,N_19806);
and UO_645 (O_645,N_19993,N_19916);
or UO_646 (O_646,N_19761,N_19978);
nor UO_647 (O_647,N_19776,N_19834);
or UO_648 (O_648,N_19900,N_19895);
nand UO_649 (O_649,N_19885,N_19819);
nand UO_650 (O_650,N_19997,N_19790);
xor UO_651 (O_651,N_19959,N_19970);
or UO_652 (O_652,N_19947,N_19952);
or UO_653 (O_653,N_19865,N_19801);
nor UO_654 (O_654,N_19865,N_19768);
nor UO_655 (O_655,N_19897,N_19876);
xnor UO_656 (O_656,N_19852,N_19751);
nand UO_657 (O_657,N_19823,N_19987);
nor UO_658 (O_658,N_19844,N_19980);
and UO_659 (O_659,N_19776,N_19934);
and UO_660 (O_660,N_19934,N_19947);
or UO_661 (O_661,N_19860,N_19972);
nor UO_662 (O_662,N_19756,N_19985);
nor UO_663 (O_663,N_19981,N_19933);
nor UO_664 (O_664,N_19893,N_19910);
xnor UO_665 (O_665,N_19972,N_19845);
nand UO_666 (O_666,N_19829,N_19889);
nand UO_667 (O_667,N_19763,N_19972);
or UO_668 (O_668,N_19867,N_19814);
or UO_669 (O_669,N_19822,N_19937);
nor UO_670 (O_670,N_19781,N_19820);
or UO_671 (O_671,N_19997,N_19981);
nor UO_672 (O_672,N_19820,N_19845);
or UO_673 (O_673,N_19888,N_19794);
nor UO_674 (O_674,N_19969,N_19818);
and UO_675 (O_675,N_19956,N_19989);
or UO_676 (O_676,N_19787,N_19838);
xor UO_677 (O_677,N_19992,N_19776);
and UO_678 (O_678,N_19802,N_19837);
and UO_679 (O_679,N_19905,N_19897);
xor UO_680 (O_680,N_19951,N_19881);
xnor UO_681 (O_681,N_19897,N_19959);
nand UO_682 (O_682,N_19765,N_19792);
xnor UO_683 (O_683,N_19818,N_19764);
xnor UO_684 (O_684,N_19907,N_19763);
nand UO_685 (O_685,N_19981,N_19801);
or UO_686 (O_686,N_19857,N_19917);
and UO_687 (O_687,N_19944,N_19982);
nand UO_688 (O_688,N_19905,N_19912);
or UO_689 (O_689,N_19752,N_19808);
nor UO_690 (O_690,N_19781,N_19998);
nor UO_691 (O_691,N_19883,N_19756);
or UO_692 (O_692,N_19955,N_19992);
nor UO_693 (O_693,N_19767,N_19891);
xor UO_694 (O_694,N_19982,N_19775);
and UO_695 (O_695,N_19890,N_19919);
nand UO_696 (O_696,N_19777,N_19754);
nand UO_697 (O_697,N_19887,N_19902);
xor UO_698 (O_698,N_19820,N_19789);
and UO_699 (O_699,N_19992,N_19982);
xnor UO_700 (O_700,N_19921,N_19810);
and UO_701 (O_701,N_19890,N_19763);
xor UO_702 (O_702,N_19967,N_19916);
and UO_703 (O_703,N_19963,N_19773);
nand UO_704 (O_704,N_19851,N_19771);
or UO_705 (O_705,N_19921,N_19970);
and UO_706 (O_706,N_19856,N_19775);
nor UO_707 (O_707,N_19996,N_19898);
xor UO_708 (O_708,N_19965,N_19908);
or UO_709 (O_709,N_19940,N_19843);
xnor UO_710 (O_710,N_19870,N_19811);
and UO_711 (O_711,N_19808,N_19775);
or UO_712 (O_712,N_19878,N_19904);
and UO_713 (O_713,N_19812,N_19754);
nor UO_714 (O_714,N_19994,N_19781);
or UO_715 (O_715,N_19895,N_19850);
and UO_716 (O_716,N_19955,N_19787);
xnor UO_717 (O_717,N_19958,N_19863);
xnor UO_718 (O_718,N_19968,N_19952);
or UO_719 (O_719,N_19938,N_19793);
or UO_720 (O_720,N_19875,N_19890);
xor UO_721 (O_721,N_19896,N_19937);
or UO_722 (O_722,N_19938,N_19964);
and UO_723 (O_723,N_19810,N_19890);
nor UO_724 (O_724,N_19861,N_19883);
nand UO_725 (O_725,N_19978,N_19896);
nor UO_726 (O_726,N_19809,N_19979);
nand UO_727 (O_727,N_19923,N_19860);
xnor UO_728 (O_728,N_19758,N_19795);
nor UO_729 (O_729,N_19948,N_19761);
xor UO_730 (O_730,N_19804,N_19923);
nand UO_731 (O_731,N_19888,N_19788);
and UO_732 (O_732,N_19766,N_19931);
xor UO_733 (O_733,N_19829,N_19855);
nor UO_734 (O_734,N_19799,N_19985);
or UO_735 (O_735,N_19883,N_19784);
nand UO_736 (O_736,N_19797,N_19863);
nor UO_737 (O_737,N_19802,N_19949);
nand UO_738 (O_738,N_19896,N_19790);
or UO_739 (O_739,N_19986,N_19751);
nand UO_740 (O_740,N_19947,N_19822);
nor UO_741 (O_741,N_19968,N_19903);
xor UO_742 (O_742,N_19918,N_19791);
nand UO_743 (O_743,N_19927,N_19970);
or UO_744 (O_744,N_19820,N_19978);
xnor UO_745 (O_745,N_19916,N_19951);
nand UO_746 (O_746,N_19819,N_19982);
and UO_747 (O_747,N_19910,N_19998);
xor UO_748 (O_748,N_19944,N_19926);
nand UO_749 (O_749,N_19908,N_19934);
and UO_750 (O_750,N_19921,N_19883);
and UO_751 (O_751,N_19765,N_19989);
or UO_752 (O_752,N_19999,N_19887);
xor UO_753 (O_753,N_19811,N_19858);
or UO_754 (O_754,N_19765,N_19768);
xor UO_755 (O_755,N_19772,N_19835);
nor UO_756 (O_756,N_19929,N_19863);
nor UO_757 (O_757,N_19852,N_19834);
or UO_758 (O_758,N_19850,N_19935);
nor UO_759 (O_759,N_19798,N_19939);
xor UO_760 (O_760,N_19834,N_19977);
nor UO_761 (O_761,N_19945,N_19754);
and UO_762 (O_762,N_19755,N_19849);
nand UO_763 (O_763,N_19850,N_19816);
nand UO_764 (O_764,N_19843,N_19759);
xnor UO_765 (O_765,N_19977,N_19903);
xnor UO_766 (O_766,N_19775,N_19842);
and UO_767 (O_767,N_19850,N_19805);
xnor UO_768 (O_768,N_19892,N_19993);
and UO_769 (O_769,N_19824,N_19981);
nand UO_770 (O_770,N_19798,N_19885);
nand UO_771 (O_771,N_19786,N_19804);
nor UO_772 (O_772,N_19768,N_19844);
or UO_773 (O_773,N_19808,N_19936);
xnor UO_774 (O_774,N_19817,N_19891);
and UO_775 (O_775,N_19952,N_19785);
or UO_776 (O_776,N_19884,N_19958);
or UO_777 (O_777,N_19962,N_19829);
xnor UO_778 (O_778,N_19989,N_19766);
nor UO_779 (O_779,N_19781,N_19999);
nor UO_780 (O_780,N_19920,N_19761);
nor UO_781 (O_781,N_19881,N_19981);
or UO_782 (O_782,N_19933,N_19907);
nor UO_783 (O_783,N_19801,N_19879);
nor UO_784 (O_784,N_19972,N_19886);
and UO_785 (O_785,N_19798,N_19783);
or UO_786 (O_786,N_19951,N_19878);
nor UO_787 (O_787,N_19916,N_19881);
and UO_788 (O_788,N_19998,N_19957);
or UO_789 (O_789,N_19884,N_19877);
nor UO_790 (O_790,N_19935,N_19893);
and UO_791 (O_791,N_19858,N_19986);
nand UO_792 (O_792,N_19916,N_19995);
xor UO_793 (O_793,N_19817,N_19846);
or UO_794 (O_794,N_19979,N_19792);
xnor UO_795 (O_795,N_19936,N_19878);
and UO_796 (O_796,N_19919,N_19850);
nand UO_797 (O_797,N_19869,N_19894);
nor UO_798 (O_798,N_19867,N_19856);
or UO_799 (O_799,N_19990,N_19931);
xor UO_800 (O_800,N_19951,N_19841);
nor UO_801 (O_801,N_19995,N_19889);
and UO_802 (O_802,N_19838,N_19914);
or UO_803 (O_803,N_19946,N_19941);
or UO_804 (O_804,N_19966,N_19842);
and UO_805 (O_805,N_19824,N_19793);
nand UO_806 (O_806,N_19927,N_19995);
or UO_807 (O_807,N_19769,N_19756);
nor UO_808 (O_808,N_19899,N_19785);
xor UO_809 (O_809,N_19980,N_19803);
nand UO_810 (O_810,N_19881,N_19958);
nor UO_811 (O_811,N_19965,N_19807);
nor UO_812 (O_812,N_19957,N_19891);
and UO_813 (O_813,N_19977,N_19875);
nor UO_814 (O_814,N_19926,N_19810);
nand UO_815 (O_815,N_19797,N_19954);
or UO_816 (O_816,N_19935,N_19788);
or UO_817 (O_817,N_19777,N_19784);
xor UO_818 (O_818,N_19784,N_19948);
xor UO_819 (O_819,N_19940,N_19882);
or UO_820 (O_820,N_19966,N_19947);
and UO_821 (O_821,N_19908,N_19800);
nor UO_822 (O_822,N_19763,N_19913);
xor UO_823 (O_823,N_19815,N_19987);
and UO_824 (O_824,N_19817,N_19918);
nor UO_825 (O_825,N_19987,N_19927);
nor UO_826 (O_826,N_19947,N_19788);
nand UO_827 (O_827,N_19931,N_19920);
nor UO_828 (O_828,N_19765,N_19955);
and UO_829 (O_829,N_19800,N_19889);
or UO_830 (O_830,N_19766,N_19850);
xor UO_831 (O_831,N_19925,N_19834);
nor UO_832 (O_832,N_19903,N_19917);
and UO_833 (O_833,N_19944,N_19961);
nor UO_834 (O_834,N_19912,N_19906);
nor UO_835 (O_835,N_19868,N_19801);
and UO_836 (O_836,N_19838,N_19921);
nor UO_837 (O_837,N_19770,N_19963);
and UO_838 (O_838,N_19778,N_19803);
nand UO_839 (O_839,N_19947,N_19789);
xor UO_840 (O_840,N_19876,N_19976);
nand UO_841 (O_841,N_19783,N_19932);
nor UO_842 (O_842,N_19914,N_19870);
nand UO_843 (O_843,N_19783,N_19764);
nor UO_844 (O_844,N_19875,N_19994);
nand UO_845 (O_845,N_19936,N_19871);
nor UO_846 (O_846,N_19934,N_19953);
and UO_847 (O_847,N_19896,N_19900);
xor UO_848 (O_848,N_19956,N_19767);
nor UO_849 (O_849,N_19778,N_19932);
xor UO_850 (O_850,N_19878,N_19930);
and UO_851 (O_851,N_19958,N_19990);
xor UO_852 (O_852,N_19774,N_19923);
nand UO_853 (O_853,N_19969,N_19812);
xor UO_854 (O_854,N_19996,N_19796);
nand UO_855 (O_855,N_19999,N_19860);
nor UO_856 (O_856,N_19974,N_19838);
and UO_857 (O_857,N_19780,N_19934);
nand UO_858 (O_858,N_19810,N_19906);
or UO_859 (O_859,N_19781,N_19789);
nand UO_860 (O_860,N_19923,N_19928);
and UO_861 (O_861,N_19827,N_19829);
and UO_862 (O_862,N_19901,N_19989);
xor UO_863 (O_863,N_19900,N_19982);
nand UO_864 (O_864,N_19853,N_19971);
xor UO_865 (O_865,N_19940,N_19957);
or UO_866 (O_866,N_19951,N_19829);
nor UO_867 (O_867,N_19876,N_19917);
or UO_868 (O_868,N_19944,N_19841);
and UO_869 (O_869,N_19840,N_19995);
and UO_870 (O_870,N_19976,N_19943);
and UO_871 (O_871,N_19901,N_19790);
nor UO_872 (O_872,N_19811,N_19753);
nand UO_873 (O_873,N_19833,N_19949);
and UO_874 (O_874,N_19872,N_19882);
nor UO_875 (O_875,N_19882,N_19995);
and UO_876 (O_876,N_19953,N_19838);
nor UO_877 (O_877,N_19995,N_19893);
and UO_878 (O_878,N_19832,N_19943);
and UO_879 (O_879,N_19798,N_19996);
nor UO_880 (O_880,N_19914,N_19790);
nand UO_881 (O_881,N_19968,N_19870);
nor UO_882 (O_882,N_19773,N_19921);
xnor UO_883 (O_883,N_19980,N_19898);
and UO_884 (O_884,N_19946,N_19773);
or UO_885 (O_885,N_19753,N_19966);
nor UO_886 (O_886,N_19907,N_19779);
or UO_887 (O_887,N_19898,N_19846);
nand UO_888 (O_888,N_19898,N_19915);
nand UO_889 (O_889,N_19821,N_19835);
and UO_890 (O_890,N_19761,N_19764);
nand UO_891 (O_891,N_19825,N_19863);
or UO_892 (O_892,N_19817,N_19949);
or UO_893 (O_893,N_19906,N_19877);
and UO_894 (O_894,N_19800,N_19878);
and UO_895 (O_895,N_19845,N_19868);
nand UO_896 (O_896,N_19995,N_19871);
and UO_897 (O_897,N_19865,N_19845);
and UO_898 (O_898,N_19850,N_19790);
nor UO_899 (O_899,N_19766,N_19980);
and UO_900 (O_900,N_19788,N_19820);
nor UO_901 (O_901,N_19974,N_19793);
xor UO_902 (O_902,N_19803,N_19759);
nand UO_903 (O_903,N_19856,N_19940);
nor UO_904 (O_904,N_19904,N_19804);
nand UO_905 (O_905,N_19859,N_19876);
or UO_906 (O_906,N_19895,N_19773);
nor UO_907 (O_907,N_19828,N_19811);
and UO_908 (O_908,N_19830,N_19985);
or UO_909 (O_909,N_19890,N_19834);
or UO_910 (O_910,N_19998,N_19818);
and UO_911 (O_911,N_19966,N_19819);
or UO_912 (O_912,N_19820,N_19910);
nor UO_913 (O_913,N_19866,N_19792);
xnor UO_914 (O_914,N_19936,N_19815);
and UO_915 (O_915,N_19827,N_19882);
nand UO_916 (O_916,N_19987,N_19825);
and UO_917 (O_917,N_19927,N_19989);
xnor UO_918 (O_918,N_19971,N_19965);
or UO_919 (O_919,N_19815,N_19763);
nand UO_920 (O_920,N_19823,N_19993);
and UO_921 (O_921,N_19856,N_19999);
or UO_922 (O_922,N_19850,N_19791);
or UO_923 (O_923,N_19810,N_19974);
nand UO_924 (O_924,N_19964,N_19800);
nand UO_925 (O_925,N_19994,N_19844);
xor UO_926 (O_926,N_19773,N_19853);
nor UO_927 (O_927,N_19982,N_19885);
nor UO_928 (O_928,N_19866,N_19758);
nor UO_929 (O_929,N_19822,N_19975);
xor UO_930 (O_930,N_19887,N_19924);
xor UO_931 (O_931,N_19833,N_19970);
nor UO_932 (O_932,N_19987,N_19799);
xnor UO_933 (O_933,N_19839,N_19825);
nor UO_934 (O_934,N_19765,N_19873);
or UO_935 (O_935,N_19759,N_19808);
nor UO_936 (O_936,N_19826,N_19824);
or UO_937 (O_937,N_19761,N_19969);
nor UO_938 (O_938,N_19845,N_19775);
nand UO_939 (O_939,N_19980,N_19875);
xor UO_940 (O_940,N_19762,N_19897);
nand UO_941 (O_941,N_19764,N_19881);
xnor UO_942 (O_942,N_19817,N_19834);
nand UO_943 (O_943,N_19885,N_19781);
and UO_944 (O_944,N_19822,N_19889);
and UO_945 (O_945,N_19894,N_19802);
nand UO_946 (O_946,N_19902,N_19867);
nor UO_947 (O_947,N_19768,N_19881);
and UO_948 (O_948,N_19801,N_19952);
nand UO_949 (O_949,N_19787,N_19839);
nand UO_950 (O_950,N_19898,N_19985);
and UO_951 (O_951,N_19996,N_19761);
nor UO_952 (O_952,N_19900,N_19953);
nor UO_953 (O_953,N_19924,N_19930);
nor UO_954 (O_954,N_19801,N_19856);
nor UO_955 (O_955,N_19861,N_19813);
or UO_956 (O_956,N_19980,N_19994);
xnor UO_957 (O_957,N_19768,N_19926);
nor UO_958 (O_958,N_19855,N_19904);
and UO_959 (O_959,N_19995,N_19787);
nor UO_960 (O_960,N_19869,N_19984);
nor UO_961 (O_961,N_19774,N_19902);
or UO_962 (O_962,N_19751,N_19930);
and UO_963 (O_963,N_19879,N_19835);
or UO_964 (O_964,N_19958,N_19838);
nor UO_965 (O_965,N_19969,N_19796);
xor UO_966 (O_966,N_19790,N_19948);
and UO_967 (O_967,N_19923,N_19907);
or UO_968 (O_968,N_19832,N_19947);
or UO_969 (O_969,N_19848,N_19762);
nand UO_970 (O_970,N_19978,N_19958);
nor UO_971 (O_971,N_19752,N_19887);
or UO_972 (O_972,N_19958,N_19973);
or UO_973 (O_973,N_19831,N_19823);
nor UO_974 (O_974,N_19890,N_19975);
xor UO_975 (O_975,N_19913,N_19788);
nand UO_976 (O_976,N_19952,N_19904);
xnor UO_977 (O_977,N_19872,N_19976);
and UO_978 (O_978,N_19793,N_19760);
or UO_979 (O_979,N_19904,N_19777);
nand UO_980 (O_980,N_19982,N_19774);
xnor UO_981 (O_981,N_19875,N_19811);
or UO_982 (O_982,N_19754,N_19837);
xor UO_983 (O_983,N_19883,N_19898);
xor UO_984 (O_984,N_19878,N_19963);
nand UO_985 (O_985,N_19801,N_19924);
and UO_986 (O_986,N_19930,N_19829);
xnor UO_987 (O_987,N_19785,N_19998);
or UO_988 (O_988,N_19780,N_19783);
and UO_989 (O_989,N_19878,N_19758);
or UO_990 (O_990,N_19926,N_19847);
xnor UO_991 (O_991,N_19978,N_19947);
and UO_992 (O_992,N_19935,N_19811);
or UO_993 (O_993,N_19808,N_19825);
nand UO_994 (O_994,N_19812,N_19768);
or UO_995 (O_995,N_19896,N_19815);
or UO_996 (O_996,N_19970,N_19938);
and UO_997 (O_997,N_19963,N_19952);
and UO_998 (O_998,N_19898,N_19835);
or UO_999 (O_999,N_19838,N_19971);
xnor UO_1000 (O_1000,N_19853,N_19763);
nand UO_1001 (O_1001,N_19791,N_19943);
nand UO_1002 (O_1002,N_19895,N_19916);
or UO_1003 (O_1003,N_19997,N_19978);
or UO_1004 (O_1004,N_19902,N_19942);
or UO_1005 (O_1005,N_19883,N_19832);
nor UO_1006 (O_1006,N_19868,N_19839);
or UO_1007 (O_1007,N_19780,N_19974);
or UO_1008 (O_1008,N_19970,N_19857);
and UO_1009 (O_1009,N_19857,N_19755);
nand UO_1010 (O_1010,N_19895,N_19831);
and UO_1011 (O_1011,N_19885,N_19768);
or UO_1012 (O_1012,N_19922,N_19869);
and UO_1013 (O_1013,N_19897,N_19783);
or UO_1014 (O_1014,N_19847,N_19893);
or UO_1015 (O_1015,N_19922,N_19885);
nand UO_1016 (O_1016,N_19784,N_19809);
nand UO_1017 (O_1017,N_19778,N_19998);
xor UO_1018 (O_1018,N_19774,N_19956);
nand UO_1019 (O_1019,N_19859,N_19924);
xnor UO_1020 (O_1020,N_19833,N_19849);
xnor UO_1021 (O_1021,N_19938,N_19933);
or UO_1022 (O_1022,N_19767,N_19812);
and UO_1023 (O_1023,N_19897,N_19968);
or UO_1024 (O_1024,N_19799,N_19816);
nor UO_1025 (O_1025,N_19816,N_19778);
nand UO_1026 (O_1026,N_19811,N_19841);
nand UO_1027 (O_1027,N_19787,N_19897);
xor UO_1028 (O_1028,N_19772,N_19923);
xor UO_1029 (O_1029,N_19763,N_19791);
and UO_1030 (O_1030,N_19771,N_19776);
nand UO_1031 (O_1031,N_19754,N_19853);
xor UO_1032 (O_1032,N_19877,N_19992);
nor UO_1033 (O_1033,N_19904,N_19857);
nand UO_1034 (O_1034,N_19756,N_19785);
nor UO_1035 (O_1035,N_19973,N_19911);
nand UO_1036 (O_1036,N_19974,N_19923);
nor UO_1037 (O_1037,N_19856,N_19855);
or UO_1038 (O_1038,N_19821,N_19897);
nor UO_1039 (O_1039,N_19913,N_19975);
xnor UO_1040 (O_1040,N_19911,N_19813);
xnor UO_1041 (O_1041,N_19870,N_19913);
or UO_1042 (O_1042,N_19887,N_19802);
nor UO_1043 (O_1043,N_19834,N_19785);
or UO_1044 (O_1044,N_19831,N_19845);
and UO_1045 (O_1045,N_19934,N_19972);
xnor UO_1046 (O_1046,N_19968,N_19752);
nand UO_1047 (O_1047,N_19868,N_19798);
or UO_1048 (O_1048,N_19986,N_19950);
nor UO_1049 (O_1049,N_19904,N_19960);
xnor UO_1050 (O_1050,N_19975,N_19933);
nand UO_1051 (O_1051,N_19991,N_19871);
nand UO_1052 (O_1052,N_19799,N_19919);
nor UO_1053 (O_1053,N_19827,N_19937);
nor UO_1054 (O_1054,N_19771,N_19869);
or UO_1055 (O_1055,N_19833,N_19817);
nor UO_1056 (O_1056,N_19955,N_19953);
nand UO_1057 (O_1057,N_19894,N_19784);
xnor UO_1058 (O_1058,N_19919,N_19887);
nand UO_1059 (O_1059,N_19955,N_19822);
or UO_1060 (O_1060,N_19925,N_19917);
and UO_1061 (O_1061,N_19758,N_19774);
nand UO_1062 (O_1062,N_19830,N_19961);
or UO_1063 (O_1063,N_19899,N_19850);
or UO_1064 (O_1064,N_19810,N_19821);
nand UO_1065 (O_1065,N_19812,N_19882);
or UO_1066 (O_1066,N_19822,N_19899);
nand UO_1067 (O_1067,N_19956,N_19931);
nand UO_1068 (O_1068,N_19960,N_19955);
and UO_1069 (O_1069,N_19830,N_19856);
nand UO_1070 (O_1070,N_19941,N_19824);
and UO_1071 (O_1071,N_19969,N_19995);
or UO_1072 (O_1072,N_19987,N_19938);
nor UO_1073 (O_1073,N_19953,N_19822);
nand UO_1074 (O_1074,N_19797,N_19986);
or UO_1075 (O_1075,N_19822,N_19866);
or UO_1076 (O_1076,N_19786,N_19757);
or UO_1077 (O_1077,N_19992,N_19964);
and UO_1078 (O_1078,N_19934,N_19839);
xor UO_1079 (O_1079,N_19859,N_19862);
or UO_1080 (O_1080,N_19880,N_19980);
or UO_1081 (O_1081,N_19969,N_19799);
xor UO_1082 (O_1082,N_19998,N_19982);
and UO_1083 (O_1083,N_19782,N_19937);
and UO_1084 (O_1084,N_19772,N_19967);
and UO_1085 (O_1085,N_19913,N_19894);
and UO_1086 (O_1086,N_19912,N_19804);
xnor UO_1087 (O_1087,N_19843,N_19877);
xnor UO_1088 (O_1088,N_19770,N_19751);
or UO_1089 (O_1089,N_19834,N_19779);
nand UO_1090 (O_1090,N_19978,N_19832);
xor UO_1091 (O_1091,N_19868,N_19926);
nor UO_1092 (O_1092,N_19956,N_19823);
nor UO_1093 (O_1093,N_19955,N_19838);
nor UO_1094 (O_1094,N_19858,N_19874);
xor UO_1095 (O_1095,N_19953,N_19754);
and UO_1096 (O_1096,N_19786,N_19920);
xnor UO_1097 (O_1097,N_19897,N_19764);
xor UO_1098 (O_1098,N_19987,N_19818);
or UO_1099 (O_1099,N_19815,N_19822);
and UO_1100 (O_1100,N_19969,N_19952);
nand UO_1101 (O_1101,N_19964,N_19812);
xor UO_1102 (O_1102,N_19987,N_19832);
nor UO_1103 (O_1103,N_19874,N_19825);
and UO_1104 (O_1104,N_19900,N_19928);
nand UO_1105 (O_1105,N_19948,N_19998);
and UO_1106 (O_1106,N_19906,N_19848);
nor UO_1107 (O_1107,N_19790,N_19785);
xnor UO_1108 (O_1108,N_19797,N_19942);
or UO_1109 (O_1109,N_19759,N_19773);
nand UO_1110 (O_1110,N_19899,N_19780);
nor UO_1111 (O_1111,N_19938,N_19844);
nor UO_1112 (O_1112,N_19821,N_19800);
xnor UO_1113 (O_1113,N_19752,N_19840);
nor UO_1114 (O_1114,N_19863,N_19907);
nand UO_1115 (O_1115,N_19833,N_19889);
or UO_1116 (O_1116,N_19980,N_19835);
or UO_1117 (O_1117,N_19881,N_19827);
nand UO_1118 (O_1118,N_19941,N_19782);
or UO_1119 (O_1119,N_19955,N_19834);
nor UO_1120 (O_1120,N_19907,N_19973);
or UO_1121 (O_1121,N_19882,N_19814);
xor UO_1122 (O_1122,N_19852,N_19955);
and UO_1123 (O_1123,N_19991,N_19870);
and UO_1124 (O_1124,N_19757,N_19862);
xor UO_1125 (O_1125,N_19797,N_19816);
nand UO_1126 (O_1126,N_19909,N_19808);
nor UO_1127 (O_1127,N_19881,N_19765);
and UO_1128 (O_1128,N_19918,N_19812);
xnor UO_1129 (O_1129,N_19857,N_19803);
nor UO_1130 (O_1130,N_19847,N_19843);
and UO_1131 (O_1131,N_19962,N_19935);
nand UO_1132 (O_1132,N_19978,N_19894);
xor UO_1133 (O_1133,N_19953,N_19936);
nand UO_1134 (O_1134,N_19870,N_19854);
xnor UO_1135 (O_1135,N_19999,N_19847);
and UO_1136 (O_1136,N_19882,N_19825);
or UO_1137 (O_1137,N_19898,N_19830);
and UO_1138 (O_1138,N_19808,N_19957);
xor UO_1139 (O_1139,N_19974,N_19910);
and UO_1140 (O_1140,N_19874,N_19890);
nor UO_1141 (O_1141,N_19875,N_19981);
nor UO_1142 (O_1142,N_19895,N_19901);
or UO_1143 (O_1143,N_19871,N_19759);
nor UO_1144 (O_1144,N_19780,N_19898);
nand UO_1145 (O_1145,N_19832,N_19772);
nand UO_1146 (O_1146,N_19865,N_19776);
xnor UO_1147 (O_1147,N_19881,N_19908);
or UO_1148 (O_1148,N_19923,N_19915);
and UO_1149 (O_1149,N_19753,N_19825);
nor UO_1150 (O_1150,N_19889,N_19977);
xnor UO_1151 (O_1151,N_19801,N_19754);
nor UO_1152 (O_1152,N_19805,N_19864);
nand UO_1153 (O_1153,N_19855,N_19753);
or UO_1154 (O_1154,N_19994,N_19972);
nand UO_1155 (O_1155,N_19885,N_19928);
and UO_1156 (O_1156,N_19875,N_19782);
or UO_1157 (O_1157,N_19916,N_19856);
nor UO_1158 (O_1158,N_19903,N_19883);
nor UO_1159 (O_1159,N_19905,N_19844);
or UO_1160 (O_1160,N_19875,N_19835);
xnor UO_1161 (O_1161,N_19899,N_19842);
nor UO_1162 (O_1162,N_19750,N_19989);
nand UO_1163 (O_1163,N_19946,N_19838);
nand UO_1164 (O_1164,N_19790,N_19783);
nand UO_1165 (O_1165,N_19860,N_19973);
or UO_1166 (O_1166,N_19968,N_19892);
or UO_1167 (O_1167,N_19795,N_19899);
xnor UO_1168 (O_1168,N_19777,N_19897);
xor UO_1169 (O_1169,N_19863,N_19754);
or UO_1170 (O_1170,N_19941,N_19842);
or UO_1171 (O_1171,N_19812,N_19824);
nor UO_1172 (O_1172,N_19842,N_19798);
and UO_1173 (O_1173,N_19808,N_19908);
nand UO_1174 (O_1174,N_19963,N_19849);
or UO_1175 (O_1175,N_19937,N_19877);
or UO_1176 (O_1176,N_19826,N_19934);
xor UO_1177 (O_1177,N_19753,N_19813);
xnor UO_1178 (O_1178,N_19760,N_19978);
xor UO_1179 (O_1179,N_19812,N_19841);
xnor UO_1180 (O_1180,N_19960,N_19775);
xor UO_1181 (O_1181,N_19912,N_19948);
and UO_1182 (O_1182,N_19903,N_19979);
and UO_1183 (O_1183,N_19881,N_19983);
xnor UO_1184 (O_1184,N_19814,N_19811);
nand UO_1185 (O_1185,N_19771,N_19765);
nor UO_1186 (O_1186,N_19776,N_19852);
or UO_1187 (O_1187,N_19918,N_19974);
xnor UO_1188 (O_1188,N_19854,N_19802);
or UO_1189 (O_1189,N_19896,N_19803);
nor UO_1190 (O_1190,N_19799,N_19788);
and UO_1191 (O_1191,N_19807,N_19830);
and UO_1192 (O_1192,N_19902,N_19776);
xor UO_1193 (O_1193,N_19963,N_19777);
and UO_1194 (O_1194,N_19904,N_19798);
nor UO_1195 (O_1195,N_19986,N_19841);
nor UO_1196 (O_1196,N_19755,N_19970);
nor UO_1197 (O_1197,N_19845,N_19787);
or UO_1198 (O_1198,N_19949,N_19900);
xor UO_1199 (O_1199,N_19946,N_19974);
nor UO_1200 (O_1200,N_19777,N_19933);
nor UO_1201 (O_1201,N_19759,N_19923);
and UO_1202 (O_1202,N_19985,N_19752);
nand UO_1203 (O_1203,N_19881,N_19863);
and UO_1204 (O_1204,N_19951,N_19875);
nor UO_1205 (O_1205,N_19948,N_19886);
or UO_1206 (O_1206,N_19996,N_19984);
or UO_1207 (O_1207,N_19973,N_19994);
nor UO_1208 (O_1208,N_19954,N_19842);
or UO_1209 (O_1209,N_19911,N_19894);
xnor UO_1210 (O_1210,N_19995,N_19868);
or UO_1211 (O_1211,N_19981,N_19986);
and UO_1212 (O_1212,N_19792,N_19787);
nand UO_1213 (O_1213,N_19800,N_19901);
xnor UO_1214 (O_1214,N_19852,N_19847);
or UO_1215 (O_1215,N_19836,N_19869);
xor UO_1216 (O_1216,N_19752,N_19978);
xnor UO_1217 (O_1217,N_19759,N_19859);
nand UO_1218 (O_1218,N_19904,N_19790);
or UO_1219 (O_1219,N_19755,N_19978);
xnor UO_1220 (O_1220,N_19797,N_19783);
or UO_1221 (O_1221,N_19755,N_19926);
xnor UO_1222 (O_1222,N_19881,N_19848);
and UO_1223 (O_1223,N_19856,N_19910);
and UO_1224 (O_1224,N_19797,N_19867);
xor UO_1225 (O_1225,N_19975,N_19978);
nor UO_1226 (O_1226,N_19883,N_19817);
nand UO_1227 (O_1227,N_19756,N_19775);
or UO_1228 (O_1228,N_19858,N_19942);
xor UO_1229 (O_1229,N_19868,N_19908);
nor UO_1230 (O_1230,N_19991,N_19922);
or UO_1231 (O_1231,N_19944,N_19828);
nand UO_1232 (O_1232,N_19853,N_19920);
nand UO_1233 (O_1233,N_19994,N_19759);
xor UO_1234 (O_1234,N_19946,N_19763);
and UO_1235 (O_1235,N_19963,N_19750);
and UO_1236 (O_1236,N_19862,N_19873);
and UO_1237 (O_1237,N_19783,N_19942);
nand UO_1238 (O_1238,N_19969,N_19891);
nand UO_1239 (O_1239,N_19805,N_19839);
or UO_1240 (O_1240,N_19806,N_19834);
nor UO_1241 (O_1241,N_19782,N_19979);
nor UO_1242 (O_1242,N_19828,N_19880);
and UO_1243 (O_1243,N_19762,N_19833);
nor UO_1244 (O_1244,N_19910,N_19757);
xnor UO_1245 (O_1245,N_19920,N_19812);
nand UO_1246 (O_1246,N_19888,N_19856);
xnor UO_1247 (O_1247,N_19930,N_19981);
nor UO_1248 (O_1248,N_19983,N_19884);
xor UO_1249 (O_1249,N_19967,N_19821);
nor UO_1250 (O_1250,N_19824,N_19854);
or UO_1251 (O_1251,N_19987,N_19801);
or UO_1252 (O_1252,N_19944,N_19943);
or UO_1253 (O_1253,N_19927,N_19875);
xnor UO_1254 (O_1254,N_19794,N_19874);
nand UO_1255 (O_1255,N_19917,N_19930);
nor UO_1256 (O_1256,N_19921,N_19798);
nand UO_1257 (O_1257,N_19937,N_19950);
and UO_1258 (O_1258,N_19764,N_19775);
nor UO_1259 (O_1259,N_19937,N_19752);
or UO_1260 (O_1260,N_19906,N_19890);
xnor UO_1261 (O_1261,N_19848,N_19903);
and UO_1262 (O_1262,N_19890,N_19923);
or UO_1263 (O_1263,N_19864,N_19768);
and UO_1264 (O_1264,N_19790,N_19835);
or UO_1265 (O_1265,N_19985,N_19893);
nor UO_1266 (O_1266,N_19777,N_19838);
and UO_1267 (O_1267,N_19976,N_19890);
xnor UO_1268 (O_1268,N_19960,N_19806);
nor UO_1269 (O_1269,N_19786,N_19771);
xor UO_1270 (O_1270,N_19986,N_19808);
and UO_1271 (O_1271,N_19835,N_19891);
nand UO_1272 (O_1272,N_19821,N_19851);
or UO_1273 (O_1273,N_19807,N_19782);
xor UO_1274 (O_1274,N_19868,N_19762);
and UO_1275 (O_1275,N_19916,N_19974);
or UO_1276 (O_1276,N_19769,N_19944);
or UO_1277 (O_1277,N_19977,N_19859);
or UO_1278 (O_1278,N_19800,N_19925);
nand UO_1279 (O_1279,N_19852,N_19770);
xnor UO_1280 (O_1280,N_19854,N_19888);
nor UO_1281 (O_1281,N_19862,N_19872);
xor UO_1282 (O_1282,N_19819,N_19889);
nor UO_1283 (O_1283,N_19929,N_19951);
and UO_1284 (O_1284,N_19784,N_19818);
nand UO_1285 (O_1285,N_19895,N_19902);
xnor UO_1286 (O_1286,N_19903,N_19755);
xor UO_1287 (O_1287,N_19816,N_19780);
and UO_1288 (O_1288,N_19978,N_19982);
nand UO_1289 (O_1289,N_19760,N_19922);
or UO_1290 (O_1290,N_19902,N_19912);
xor UO_1291 (O_1291,N_19794,N_19876);
and UO_1292 (O_1292,N_19985,N_19994);
or UO_1293 (O_1293,N_19848,N_19812);
and UO_1294 (O_1294,N_19935,N_19853);
nor UO_1295 (O_1295,N_19853,N_19918);
or UO_1296 (O_1296,N_19927,N_19787);
and UO_1297 (O_1297,N_19802,N_19750);
xnor UO_1298 (O_1298,N_19847,N_19792);
xnor UO_1299 (O_1299,N_19959,N_19775);
and UO_1300 (O_1300,N_19907,N_19853);
and UO_1301 (O_1301,N_19972,N_19853);
nor UO_1302 (O_1302,N_19828,N_19847);
nor UO_1303 (O_1303,N_19934,N_19932);
or UO_1304 (O_1304,N_19791,N_19820);
nand UO_1305 (O_1305,N_19864,N_19874);
nor UO_1306 (O_1306,N_19922,N_19993);
nand UO_1307 (O_1307,N_19821,N_19928);
nor UO_1308 (O_1308,N_19770,N_19789);
nor UO_1309 (O_1309,N_19850,N_19981);
or UO_1310 (O_1310,N_19893,N_19785);
nor UO_1311 (O_1311,N_19789,N_19957);
or UO_1312 (O_1312,N_19953,N_19899);
xor UO_1313 (O_1313,N_19887,N_19750);
nor UO_1314 (O_1314,N_19831,N_19779);
xor UO_1315 (O_1315,N_19981,N_19926);
nor UO_1316 (O_1316,N_19965,N_19796);
xor UO_1317 (O_1317,N_19809,N_19945);
nor UO_1318 (O_1318,N_19823,N_19760);
nand UO_1319 (O_1319,N_19997,N_19884);
and UO_1320 (O_1320,N_19857,N_19760);
and UO_1321 (O_1321,N_19752,N_19874);
or UO_1322 (O_1322,N_19950,N_19842);
and UO_1323 (O_1323,N_19820,N_19786);
xor UO_1324 (O_1324,N_19773,N_19908);
or UO_1325 (O_1325,N_19821,N_19990);
nand UO_1326 (O_1326,N_19844,N_19922);
nand UO_1327 (O_1327,N_19976,N_19812);
nand UO_1328 (O_1328,N_19791,N_19885);
nand UO_1329 (O_1329,N_19789,N_19949);
or UO_1330 (O_1330,N_19750,N_19775);
or UO_1331 (O_1331,N_19796,N_19913);
or UO_1332 (O_1332,N_19794,N_19796);
xor UO_1333 (O_1333,N_19978,N_19969);
or UO_1334 (O_1334,N_19903,N_19851);
nor UO_1335 (O_1335,N_19779,N_19935);
nor UO_1336 (O_1336,N_19966,N_19843);
nand UO_1337 (O_1337,N_19870,N_19868);
nor UO_1338 (O_1338,N_19903,N_19798);
and UO_1339 (O_1339,N_19893,N_19819);
nand UO_1340 (O_1340,N_19832,N_19995);
xor UO_1341 (O_1341,N_19909,N_19908);
nor UO_1342 (O_1342,N_19777,N_19797);
xnor UO_1343 (O_1343,N_19868,N_19788);
nand UO_1344 (O_1344,N_19949,N_19884);
nand UO_1345 (O_1345,N_19906,N_19818);
nor UO_1346 (O_1346,N_19811,N_19955);
nor UO_1347 (O_1347,N_19946,N_19928);
and UO_1348 (O_1348,N_19897,N_19851);
nor UO_1349 (O_1349,N_19984,N_19817);
xnor UO_1350 (O_1350,N_19940,N_19950);
nand UO_1351 (O_1351,N_19769,N_19788);
nor UO_1352 (O_1352,N_19776,N_19913);
nand UO_1353 (O_1353,N_19808,N_19877);
nor UO_1354 (O_1354,N_19753,N_19961);
nor UO_1355 (O_1355,N_19953,N_19901);
and UO_1356 (O_1356,N_19826,N_19999);
and UO_1357 (O_1357,N_19775,N_19802);
nor UO_1358 (O_1358,N_19785,N_19994);
nand UO_1359 (O_1359,N_19753,N_19948);
or UO_1360 (O_1360,N_19993,N_19929);
xor UO_1361 (O_1361,N_19914,N_19823);
nor UO_1362 (O_1362,N_19879,N_19782);
and UO_1363 (O_1363,N_19855,N_19967);
nor UO_1364 (O_1364,N_19824,N_19788);
or UO_1365 (O_1365,N_19876,N_19819);
or UO_1366 (O_1366,N_19928,N_19774);
and UO_1367 (O_1367,N_19777,N_19853);
xor UO_1368 (O_1368,N_19985,N_19835);
nor UO_1369 (O_1369,N_19999,N_19851);
and UO_1370 (O_1370,N_19782,N_19878);
and UO_1371 (O_1371,N_19966,N_19846);
or UO_1372 (O_1372,N_19788,N_19957);
nor UO_1373 (O_1373,N_19762,N_19984);
xor UO_1374 (O_1374,N_19763,N_19995);
or UO_1375 (O_1375,N_19807,N_19783);
nand UO_1376 (O_1376,N_19898,N_19945);
nor UO_1377 (O_1377,N_19880,N_19995);
nand UO_1378 (O_1378,N_19841,N_19984);
and UO_1379 (O_1379,N_19975,N_19762);
or UO_1380 (O_1380,N_19869,N_19829);
and UO_1381 (O_1381,N_19823,N_19766);
xnor UO_1382 (O_1382,N_19866,N_19864);
nor UO_1383 (O_1383,N_19911,N_19941);
xor UO_1384 (O_1384,N_19980,N_19832);
or UO_1385 (O_1385,N_19790,N_19935);
and UO_1386 (O_1386,N_19950,N_19839);
nand UO_1387 (O_1387,N_19798,N_19913);
xnor UO_1388 (O_1388,N_19876,N_19762);
nand UO_1389 (O_1389,N_19975,N_19779);
nand UO_1390 (O_1390,N_19966,N_19781);
or UO_1391 (O_1391,N_19931,N_19852);
or UO_1392 (O_1392,N_19808,N_19822);
xnor UO_1393 (O_1393,N_19807,N_19905);
nand UO_1394 (O_1394,N_19754,N_19912);
nand UO_1395 (O_1395,N_19820,N_19896);
or UO_1396 (O_1396,N_19768,N_19985);
nor UO_1397 (O_1397,N_19811,N_19990);
nor UO_1398 (O_1398,N_19955,N_19859);
or UO_1399 (O_1399,N_19793,N_19844);
nand UO_1400 (O_1400,N_19800,N_19987);
nand UO_1401 (O_1401,N_19816,N_19855);
xnor UO_1402 (O_1402,N_19764,N_19941);
nor UO_1403 (O_1403,N_19954,N_19940);
and UO_1404 (O_1404,N_19984,N_19943);
xor UO_1405 (O_1405,N_19887,N_19858);
or UO_1406 (O_1406,N_19819,N_19976);
xor UO_1407 (O_1407,N_19905,N_19983);
xnor UO_1408 (O_1408,N_19931,N_19829);
nor UO_1409 (O_1409,N_19915,N_19895);
nor UO_1410 (O_1410,N_19878,N_19920);
nor UO_1411 (O_1411,N_19848,N_19939);
xnor UO_1412 (O_1412,N_19926,N_19921);
nor UO_1413 (O_1413,N_19789,N_19852);
and UO_1414 (O_1414,N_19940,N_19945);
nor UO_1415 (O_1415,N_19867,N_19937);
or UO_1416 (O_1416,N_19938,N_19865);
nor UO_1417 (O_1417,N_19902,N_19934);
and UO_1418 (O_1418,N_19925,N_19968);
nor UO_1419 (O_1419,N_19883,N_19889);
nor UO_1420 (O_1420,N_19853,N_19881);
nor UO_1421 (O_1421,N_19872,N_19795);
nand UO_1422 (O_1422,N_19865,N_19880);
nor UO_1423 (O_1423,N_19763,N_19869);
and UO_1424 (O_1424,N_19790,N_19976);
nor UO_1425 (O_1425,N_19836,N_19997);
nor UO_1426 (O_1426,N_19855,N_19795);
nor UO_1427 (O_1427,N_19813,N_19949);
or UO_1428 (O_1428,N_19855,N_19811);
or UO_1429 (O_1429,N_19844,N_19876);
xnor UO_1430 (O_1430,N_19837,N_19752);
and UO_1431 (O_1431,N_19958,N_19799);
nand UO_1432 (O_1432,N_19844,N_19823);
and UO_1433 (O_1433,N_19999,N_19877);
or UO_1434 (O_1434,N_19960,N_19883);
and UO_1435 (O_1435,N_19948,N_19770);
or UO_1436 (O_1436,N_19923,N_19851);
nor UO_1437 (O_1437,N_19756,N_19942);
or UO_1438 (O_1438,N_19979,N_19915);
or UO_1439 (O_1439,N_19804,N_19864);
nand UO_1440 (O_1440,N_19940,N_19924);
and UO_1441 (O_1441,N_19762,N_19964);
or UO_1442 (O_1442,N_19750,N_19954);
or UO_1443 (O_1443,N_19860,N_19908);
or UO_1444 (O_1444,N_19812,N_19917);
or UO_1445 (O_1445,N_19840,N_19765);
nor UO_1446 (O_1446,N_19982,N_19762);
xor UO_1447 (O_1447,N_19881,N_19987);
and UO_1448 (O_1448,N_19768,N_19831);
nor UO_1449 (O_1449,N_19964,N_19854);
nand UO_1450 (O_1450,N_19911,N_19784);
or UO_1451 (O_1451,N_19883,N_19963);
nor UO_1452 (O_1452,N_19958,N_19976);
nor UO_1453 (O_1453,N_19832,N_19825);
or UO_1454 (O_1454,N_19784,N_19802);
nor UO_1455 (O_1455,N_19833,N_19911);
nand UO_1456 (O_1456,N_19766,N_19756);
or UO_1457 (O_1457,N_19815,N_19962);
nor UO_1458 (O_1458,N_19985,N_19849);
nand UO_1459 (O_1459,N_19846,N_19993);
and UO_1460 (O_1460,N_19760,N_19997);
xor UO_1461 (O_1461,N_19807,N_19967);
nand UO_1462 (O_1462,N_19896,N_19843);
or UO_1463 (O_1463,N_19934,N_19983);
and UO_1464 (O_1464,N_19813,N_19768);
nand UO_1465 (O_1465,N_19931,N_19775);
nand UO_1466 (O_1466,N_19978,N_19817);
xnor UO_1467 (O_1467,N_19991,N_19986);
xnor UO_1468 (O_1468,N_19999,N_19757);
xnor UO_1469 (O_1469,N_19758,N_19893);
xor UO_1470 (O_1470,N_19966,N_19890);
and UO_1471 (O_1471,N_19845,N_19900);
and UO_1472 (O_1472,N_19961,N_19837);
or UO_1473 (O_1473,N_19924,N_19820);
and UO_1474 (O_1474,N_19987,N_19803);
and UO_1475 (O_1475,N_19752,N_19835);
nand UO_1476 (O_1476,N_19888,N_19870);
nand UO_1477 (O_1477,N_19895,N_19784);
and UO_1478 (O_1478,N_19801,N_19896);
or UO_1479 (O_1479,N_19905,N_19750);
xor UO_1480 (O_1480,N_19910,N_19939);
nand UO_1481 (O_1481,N_19803,N_19892);
and UO_1482 (O_1482,N_19901,N_19853);
and UO_1483 (O_1483,N_19879,N_19933);
and UO_1484 (O_1484,N_19836,N_19808);
or UO_1485 (O_1485,N_19900,N_19967);
or UO_1486 (O_1486,N_19999,N_19871);
and UO_1487 (O_1487,N_19812,N_19899);
or UO_1488 (O_1488,N_19910,N_19763);
and UO_1489 (O_1489,N_19921,N_19885);
xor UO_1490 (O_1490,N_19887,N_19835);
nand UO_1491 (O_1491,N_19803,N_19990);
or UO_1492 (O_1492,N_19763,N_19993);
nand UO_1493 (O_1493,N_19794,N_19833);
or UO_1494 (O_1494,N_19886,N_19957);
nand UO_1495 (O_1495,N_19759,N_19967);
or UO_1496 (O_1496,N_19826,N_19866);
or UO_1497 (O_1497,N_19968,N_19987);
or UO_1498 (O_1498,N_19767,N_19972);
and UO_1499 (O_1499,N_19935,N_19839);
or UO_1500 (O_1500,N_19855,N_19991);
nor UO_1501 (O_1501,N_19756,N_19777);
nand UO_1502 (O_1502,N_19899,N_19957);
nand UO_1503 (O_1503,N_19774,N_19983);
and UO_1504 (O_1504,N_19877,N_19971);
and UO_1505 (O_1505,N_19969,N_19879);
nor UO_1506 (O_1506,N_19782,N_19810);
xor UO_1507 (O_1507,N_19768,N_19896);
or UO_1508 (O_1508,N_19789,N_19848);
xor UO_1509 (O_1509,N_19794,N_19893);
nand UO_1510 (O_1510,N_19971,N_19866);
and UO_1511 (O_1511,N_19980,N_19870);
xor UO_1512 (O_1512,N_19815,N_19784);
or UO_1513 (O_1513,N_19839,N_19789);
nor UO_1514 (O_1514,N_19868,N_19802);
or UO_1515 (O_1515,N_19858,N_19838);
and UO_1516 (O_1516,N_19837,N_19795);
and UO_1517 (O_1517,N_19969,N_19821);
nor UO_1518 (O_1518,N_19781,N_19855);
nand UO_1519 (O_1519,N_19968,N_19845);
nor UO_1520 (O_1520,N_19782,N_19928);
xnor UO_1521 (O_1521,N_19965,N_19872);
or UO_1522 (O_1522,N_19953,N_19987);
xor UO_1523 (O_1523,N_19989,N_19907);
nor UO_1524 (O_1524,N_19829,N_19857);
or UO_1525 (O_1525,N_19997,N_19942);
nor UO_1526 (O_1526,N_19974,N_19814);
and UO_1527 (O_1527,N_19853,N_19949);
nand UO_1528 (O_1528,N_19847,N_19802);
or UO_1529 (O_1529,N_19981,N_19751);
and UO_1530 (O_1530,N_19888,N_19879);
nor UO_1531 (O_1531,N_19953,N_19950);
or UO_1532 (O_1532,N_19994,N_19997);
or UO_1533 (O_1533,N_19925,N_19816);
or UO_1534 (O_1534,N_19852,N_19794);
nand UO_1535 (O_1535,N_19899,N_19835);
xnor UO_1536 (O_1536,N_19838,N_19833);
nor UO_1537 (O_1537,N_19806,N_19987);
nor UO_1538 (O_1538,N_19806,N_19993);
and UO_1539 (O_1539,N_19925,N_19948);
or UO_1540 (O_1540,N_19869,N_19982);
xnor UO_1541 (O_1541,N_19778,N_19838);
xor UO_1542 (O_1542,N_19933,N_19962);
and UO_1543 (O_1543,N_19985,N_19769);
and UO_1544 (O_1544,N_19994,N_19818);
xor UO_1545 (O_1545,N_19812,N_19982);
nand UO_1546 (O_1546,N_19837,N_19844);
or UO_1547 (O_1547,N_19806,N_19884);
nand UO_1548 (O_1548,N_19770,N_19833);
and UO_1549 (O_1549,N_19904,N_19834);
or UO_1550 (O_1550,N_19912,N_19818);
nor UO_1551 (O_1551,N_19800,N_19971);
and UO_1552 (O_1552,N_19838,N_19934);
nand UO_1553 (O_1553,N_19903,N_19776);
nand UO_1554 (O_1554,N_19916,N_19872);
xnor UO_1555 (O_1555,N_19939,N_19889);
nand UO_1556 (O_1556,N_19804,N_19947);
nor UO_1557 (O_1557,N_19924,N_19805);
or UO_1558 (O_1558,N_19885,N_19880);
nand UO_1559 (O_1559,N_19804,N_19850);
nand UO_1560 (O_1560,N_19963,N_19872);
xnor UO_1561 (O_1561,N_19755,N_19832);
nor UO_1562 (O_1562,N_19832,N_19919);
or UO_1563 (O_1563,N_19861,N_19868);
xnor UO_1564 (O_1564,N_19784,N_19923);
nand UO_1565 (O_1565,N_19805,N_19917);
nand UO_1566 (O_1566,N_19807,N_19983);
xor UO_1567 (O_1567,N_19984,N_19862);
or UO_1568 (O_1568,N_19832,N_19790);
nor UO_1569 (O_1569,N_19818,N_19768);
and UO_1570 (O_1570,N_19894,N_19785);
nor UO_1571 (O_1571,N_19940,N_19956);
nand UO_1572 (O_1572,N_19980,N_19904);
nand UO_1573 (O_1573,N_19921,N_19917);
or UO_1574 (O_1574,N_19895,N_19811);
xor UO_1575 (O_1575,N_19909,N_19754);
or UO_1576 (O_1576,N_19864,N_19945);
xnor UO_1577 (O_1577,N_19850,N_19906);
or UO_1578 (O_1578,N_19891,N_19779);
nand UO_1579 (O_1579,N_19964,N_19985);
or UO_1580 (O_1580,N_19901,N_19944);
or UO_1581 (O_1581,N_19977,N_19928);
xor UO_1582 (O_1582,N_19947,N_19835);
nand UO_1583 (O_1583,N_19806,N_19869);
nor UO_1584 (O_1584,N_19774,N_19798);
xnor UO_1585 (O_1585,N_19878,N_19751);
or UO_1586 (O_1586,N_19819,N_19868);
nor UO_1587 (O_1587,N_19995,N_19964);
or UO_1588 (O_1588,N_19906,N_19842);
nor UO_1589 (O_1589,N_19881,N_19872);
nor UO_1590 (O_1590,N_19879,N_19808);
and UO_1591 (O_1591,N_19978,N_19897);
xnor UO_1592 (O_1592,N_19832,N_19935);
nor UO_1593 (O_1593,N_19929,N_19764);
nand UO_1594 (O_1594,N_19972,N_19778);
xnor UO_1595 (O_1595,N_19853,N_19893);
and UO_1596 (O_1596,N_19792,N_19835);
nor UO_1597 (O_1597,N_19983,N_19963);
nor UO_1598 (O_1598,N_19772,N_19904);
or UO_1599 (O_1599,N_19829,N_19870);
or UO_1600 (O_1600,N_19791,N_19919);
nor UO_1601 (O_1601,N_19999,N_19966);
nor UO_1602 (O_1602,N_19819,N_19953);
nor UO_1603 (O_1603,N_19944,N_19815);
nand UO_1604 (O_1604,N_19924,N_19868);
xnor UO_1605 (O_1605,N_19820,N_19936);
nor UO_1606 (O_1606,N_19914,N_19768);
and UO_1607 (O_1607,N_19807,N_19940);
xnor UO_1608 (O_1608,N_19792,N_19877);
or UO_1609 (O_1609,N_19976,N_19841);
nand UO_1610 (O_1610,N_19893,N_19811);
nand UO_1611 (O_1611,N_19762,N_19941);
xor UO_1612 (O_1612,N_19973,N_19990);
xnor UO_1613 (O_1613,N_19769,N_19906);
and UO_1614 (O_1614,N_19836,N_19928);
and UO_1615 (O_1615,N_19947,N_19770);
and UO_1616 (O_1616,N_19986,N_19819);
or UO_1617 (O_1617,N_19872,N_19936);
nor UO_1618 (O_1618,N_19919,N_19926);
and UO_1619 (O_1619,N_19901,N_19913);
xor UO_1620 (O_1620,N_19900,N_19829);
and UO_1621 (O_1621,N_19990,N_19768);
nor UO_1622 (O_1622,N_19940,N_19892);
nand UO_1623 (O_1623,N_19759,N_19839);
or UO_1624 (O_1624,N_19953,N_19998);
and UO_1625 (O_1625,N_19918,N_19864);
nand UO_1626 (O_1626,N_19998,N_19787);
and UO_1627 (O_1627,N_19871,N_19805);
nand UO_1628 (O_1628,N_19943,N_19949);
and UO_1629 (O_1629,N_19997,N_19915);
or UO_1630 (O_1630,N_19966,N_19886);
and UO_1631 (O_1631,N_19876,N_19793);
xor UO_1632 (O_1632,N_19803,N_19859);
nand UO_1633 (O_1633,N_19939,N_19911);
nand UO_1634 (O_1634,N_19830,N_19914);
and UO_1635 (O_1635,N_19799,N_19920);
xor UO_1636 (O_1636,N_19885,N_19894);
nor UO_1637 (O_1637,N_19934,N_19927);
and UO_1638 (O_1638,N_19833,N_19790);
xor UO_1639 (O_1639,N_19898,N_19998);
nand UO_1640 (O_1640,N_19956,N_19794);
nor UO_1641 (O_1641,N_19905,N_19967);
and UO_1642 (O_1642,N_19821,N_19866);
or UO_1643 (O_1643,N_19931,N_19944);
and UO_1644 (O_1644,N_19826,N_19802);
nand UO_1645 (O_1645,N_19781,N_19861);
and UO_1646 (O_1646,N_19860,N_19827);
and UO_1647 (O_1647,N_19887,N_19827);
nor UO_1648 (O_1648,N_19899,N_19855);
xnor UO_1649 (O_1649,N_19968,N_19907);
or UO_1650 (O_1650,N_19792,N_19951);
xnor UO_1651 (O_1651,N_19930,N_19882);
or UO_1652 (O_1652,N_19935,N_19785);
nand UO_1653 (O_1653,N_19933,N_19958);
or UO_1654 (O_1654,N_19763,N_19822);
xor UO_1655 (O_1655,N_19845,N_19846);
or UO_1656 (O_1656,N_19849,N_19908);
xor UO_1657 (O_1657,N_19758,N_19947);
nor UO_1658 (O_1658,N_19797,N_19996);
nand UO_1659 (O_1659,N_19937,N_19962);
xor UO_1660 (O_1660,N_19762,N_19927);
and UO_1661 (O_1661,N_19939,N_19864);
nor UO_1662 (O_1662,N_19815,N_19861);
nand UO_1663 (O_1663,N_19780,N_19784);
or UO_1664 (O_1664,N_19824,N_19827);
nand UO_1665 (O_1665,N_19907,N_19759);
or UO_1666 (O_1666,N_19888,N_19874);
and UO_1667 (O_1667,N_19770,N_19971);
nand UO_1668 (O_1668,N_19988,N_19759);
and UO_1669 (O_1669,N_19866,N_19994);
or UO_1670 (O_1670,N_19994,N_19856);
nand UO_1671 (O_1671,N_19875,N_19775);
or UO_1672 (O_1672,N_19821,N_19834);
xnor UO_1673 (O_1673,N_19831,N_19865);
nor UO_1674 (O_1674,N_19953,N_19863);
xnor UO_1675 (O_1675,N_19784,N_19841);
nor UO_1676 (O_1676,N_19768,N_19945);
and UO_1677 (O_1677,N_19821,N_19868);
and UO_1678 (O_1678,N_19934,N_19876);
nor UO_1679 (O_1679,N_19953,N_19787);
nor UO_1680 (O_1680,N_19911,N_19926);
xor UO_1681 (O_1681,N_19873,N_19772);
nand UO_1682 (O_1682,N_19939,N_19903);
nand UO_1683 (O_1683,N_19756,N_19780);
xor UO_1684 (O_1684,N_19830,N_19997);
xnor UO_1685 (O_1685,N_19771,N_19928);
nor UO_1686 (O_1686,N_19861,N_19929);
and UO_1687 (O_1687,N_19843,N_19830);
xnor UO_1688 (O_1688,N_19892,N_19854);
xor UO_1689 (O_1689,N_19964,N_19900);
nand UO_1690 (O_1690,N_19835,N_19851);
nand UO_1691 (O_1691,N_19914,N_19942);
xor UO_1692 (O_1692,N_19758,N_19890);
nand UO_1693 (O_1693,N_19978,N_19877);
or UO_1694 (O_1694,N_19919,N_19833);
nand UO_1695 (O_1695,N_19960,N_19858);
nor UO_1696 (O_1696,N_19893,N_19776);
or UO_1697 (O_1697,N_19925,N_19867);
or UO_1698 (O_1698,N_19947,N_19941);
or UO_1699 (O_1699,N_19760,N_19963);
nand UO_1700 (O_1700,N_19874,N_19929);
or UO_1701 (O_1701,N_19951,N_19995);
xor UO_1702 (O_1702,N_19979,N_19904);
xnor UO_1703 (O_1703,N_19781,N_19895);
and UO_1704 (O_1704,N_19881,N_19796);
nor UO_1705 (O_1705,N_19951,N_19865);
nand UO_1706 (O_1706,N_19824,N_19760);
nand UO_1707 (O_1707,N_19885,N_19780);
nand UO_1708 (O_1708,N_19826,N_19761);
nor UO_1709 (O_1709,N_19760,N_19836);
and UO_1710 (O_1710,N_19930,N_19768);
nor UO_1711 (O_1711,N_19905,N_19951);
xnor UO_1712 (O_1712,N_19967,N_19878);
xor UO_1713 (O_1713,N_19997,N_19801);
or UO_1714 (O_1714,N_19766,N_19840);
xor UO_1715 (O_1715,N_19964,N_19777);
nand UO_1716 (O_1716,N_19830,N_19770);
nor UO_1717 (O_1717,N_19864,N_19958);
xor UO_1718 (O_1718,N_19810,N_19759);
nor UO_1719 (O_1719,N_19823,N_19977);
nand UO_1720 (O_1720,N_19861,N_19872);
xnor UO_1721 (O_1721,N_19800,N_19907);
or UO_1722 (O_1722,N_19923,N_19872);
or UO_1723 (O_1723,N_19984,N_19767);
and UO_1724 (O_1724,N_19959,N_19760);
nor UO_1725 (O_1725,N_19968,N_19885);
or UO_1726 (O_1726,N_19810,N_19798);
nand UO_1727 (O_1727,N_19858,N_19855);
nand UO_1728 (O_1728,N_19818,N_19929);
nand UO_1729 (O_1729,N_19750,N_19824);
xor UO_1730 (O_1730,N_19888,N_19785);
nand UO_1731 (O_1731,N_19975,N_19787);
nor UO_1732 (O_1732,N_19949,N_19808);
or UO_1733 (O_1733,N_19773,N_19944);
nand UO_1734 (O_1734,N_19755,N_19770);
xnor UO_1735 (O_1735,N_19916,N_19914);
and UO_1736 (O_1736,N_19856,N_19785);
nor UO_1737 (O_1737,N_19974,N_19928);
or UO_1738 (O_1738,N_19934,N_19887);
xor UO_1739 (O_1739,N_19774,N_19903);
and UO_1740 (O_1740,N_19769,N_19861);
xnor UO_1741 (O_1741,N_19899,N_19809);
and UO_1742 (O_1742,N_19879,N_19908);
xor UO_1743 (O_1743,N_19908,N_19799);
nor UO_1744 (O_1744,N_19869,N_19979);
nand UO_1745 (O_1745,N_19879,N_19774);
nor UO_1746 (O_1746,N_19830,N_19841);
nor UO_1747 (O_1747,N_19981,N_19790);
nor UO_1748 (O_1748,N_19775,N_19780);
xor UO_1749 (O_1749,N_19757,N_19803);
and UO_1750 (O_1750,N_19814,N_19816);
xnor UO_1751 (O_1751,N_19768,N_19773);
or UO_1752 (O_1752,N_19764,N_19853);
and UO_1753 (O_1753,N_19760,N_19803);
nand UO_1754 (O_1754,N_19794,N_19750);
and UO_1755 (O_1755,N_19787,N_19759);
nand UO_1756 (O_1756,N_19754,N_19818);
or UO_1757 (O_1757,N_19773,N_19795);
nand UO_1758 (O_1758,N_19969,N_19807);
nand UO_1759 (O_1759,N_19788,N_19896);
or UO_1760 (O_1760,N_19945,N_19817);
nand UO_1761 (O_1761,N_19847,N_19861);
xnor UO_1762 (O_1762,N_19878,N_19884);
and UO_1763 (O_1763,N_19912,N_19753);
nand UO_1764 (O_1764,N_19954,N_19929);
and UO_1765 (O_1765,N_19857,N_19824);
and UO_1766 (O_1766,N_19778,N_19882);
nand UO_1767 (O_1767,N_19840,N_19839);
and UO_1768 (O_1768,N_19757,N_19873);
and UO_1769 (O_1769,N_19992,N_19884);
and UO_1770 (O_1770,N_19987,N_19847);
xnor UO_1771 (O_1771,N_19889,N_19894);
and UO_1772 (O_1772,N_19991,N_19889);
and UO_1773 (O_1773,N_19862,N_19992);
nand UO_1774 (O_1774,N_19852,N_19821);
nor UO_1775 (O_1775,N_19867,N_19985);
xnor UO_1776 (O_1776,N_19771,N_19770);
or UO_1777 (O_1777,N_19765,N_19956);
nand UO_1778 (O_1778,N_19995,N_19895);
or UO_1779 (O_1779,N_19796,N_19944);
nand UO_1780 (O_1780,N_19998,N_19761);
or UO_1781 (O_1781,N_19946,N_19968);
nand UO_1782 (O_1782,N_19983,N_19866);
xor UO_1783 (O_1783,N_19909,N_19780);
nor UO_1784 (O_1784,N_19978,N_19753);
nand UO_1785 (O_1785,N_19779,N_19943);
or UO_1786 (O_1786,N_19784,N_19844);
nor UO_1787 (O_1787,N_19767,N_19755);
or UO_1788 (O_1788,N_19898,N_19791);
nor UO_1789 (O_1789,N_19793,N_19825);
nor UO_1790 (O_1790,N_19983,N_19838);
or UO_1791 (O_1791,N_19826,N_19923);
or UO_1792 (O_1792,N_19943,N_19971);
nor UO_1793 (O_1793,N_19826,N_19782);
or UO_1794 (O_1794,N_19872,N_19887);
nand UO_1795 (O_1795,N_19904,N_19911);
or UO_1796 (O_1796,N_19914,N_19806);
nor UO_1797 (O_1797,N_19955,N_19872);
nand UO_1798 (O_1798,N_19957,N_19778);
xnor UO_1799 (O_1799,N_19785,N_19855);
or UO_1800 (O_1800,N_19946,N_19989);
nor UO_1801 (O_1801,N_19830,N_19767);
nand UO_1802 (O_1802,N_19794,N_19840);
and UO_1803 (O_1803,N_19876,N_19953);
nand UO_1804 (O_1804,N_19958,N_19991);
or UO_1805 (O_1805,N_19866,N_19870);
nand UO_1806 (O_1806,N_19970,N_19976);
and UO_1807 (O_1807,N_19752,N_19932);
and UO_1808 (O_1808,N_19845,N_19937);
or UO_1809 (O_1809,N_19873,N_19888);
and UO_1810 (O_1810,N_19827,N_19812);
nor UO_1811 (O_1811,N_19798,N_19862);
nand UO_1812 (O_1812,N_19914,N_19986);
nor UO_1813 (O_1813,N_19891,N_19968);
and UO_1814 (O_1814,N_19807,N_19767);
or UO_1815 (O_1815,N_19833,N_19967);
nor UO_1816 (O_1816,N_19780,N_19911);
xor UO_1817 (O_1817,N_19861,N_19836);
nand UO_1818 (O_1818,N_19859,N_19900);
and UO_1819 (O_1819,N_19764,N_19995);
nand UO_1820 (O_1820,N_19948,N_19891);
xnor UO_1821 (O_1821,N_19853,N_19817);
xor UO_1822 (O_1822,N_19936,N_19823);
and UO_1823 (O_1823,N_19850,N_19936);
or UO_1824 (O_1824,N_19803,N_19947);
xor UO_1825 (O_1825,N_19787,N_19794);
and UO_1826 (O_1826,N_19803,N_19810);
nand UO_1827 (O_1827,N_19892,N_19781);
or UO_1828 (O_1828,N_19928,N_19813);
nand UO_1829 (O_1829,N_19877,N_19996);
and UO_1830 (O_1830,N_19980,N_19778);
and UO_1831 (O_1831,N_19837,N_19913);
nor UO_1832 (O_1832,N_19799,N_19851);
nor UO_1833 (O_1833,N_19850,N_19761);
nand UO_1834 (O_1834,N_19867,N_19900);
and UO_1835 (O_1835,N_19901,N_19755);
and UO_1836 (O_1836,N_19768,N_19950);
and UO_1837 (O_1837,N_19930,N_19845);
nor UO_1838 (O_1838,N_19758,N_19853);
nor UO_1839 (O_1839,N_19919,N_19894);
nor UO_1840 (O_1840,N_19994,N_19794);
or UO_1841 (O_1841,N_19938,N_19807);
and UO_1842 (O_1842,N_19975,N_19886);
and UO_1843 (O_1843,N_19753,N_19887);
xor UO_1844 (O_1844,N_19849,N_19972);
xor UO_1845 (O_1845,N_19818,N_19992);
or UO_1846 (O_1846,N_19861,N_19793);
and UO_1847 (O_1847,N_19972,N_19929);
nor UO_1848 (O_1848,N_19956,N_19819);
or UO_1849 (O_1849,N_19785,N_19827);
and UO_1850 (O_1850,N_19972,N_19862);
or UO_1851 (O_1851,N_19960,N_19875);
nor UO_1852 (O_1852,N_19929,N_19792);
or UO_1853 (O_1853,N_19774,N_19955);
or UO_1854 (O_1854,N_19985,N_19890);
and UO_1855 (O_1855,N_19998,N_19823);
or UO_1856 (O_1856,N_19761,N_19794);
nor UO_1857 (O_1857,N_19877,N_19807);
or UO_1858 (O_1858,N_19867,N_19829);
xor UO_1859 (O_1859,N_19904,N_19902);
or UO_1860 (O_1860,N_19876,N_19966);
nand UO_1861 (O_1861,N_19755,N_19971);
nand UO_1862 (O_1862,N_19939,N_19818);
nand UO_1863 (O_1863,N_19950,N_19836);
xnor UO_1864 (O_1864,N_19996,N_19932);
and UO_1865 (O_1865,N_19832,N_19920);
or UO_1866 (O_1866,N_19949,N_19913);
or UO_1867 (O_1867,N_19856,N_19900);
nand UO_1868 (O_1868,N_19953,N_19914);
nor UO_1869 (O_1869,N_19860,N_19967);
xnor UO_1870 (O_1870,N_19895,N_19987);
or UO_1871 (O_1871,N_19977,N_19798);
nand UO_1872 (O_1872,N_19975,N_19849);
xnor UO_1873 (O_1873,N_19800,N_19886);
and UO_1874 (O_1874,N_19898,N_19970);
or UO_1875 (O_1875,N_19955,N_19889);
xnor UO_1876 (O_1876,N_19961,N_19769);
and UO_1877 (O_1877,N_19994,N_19883);
and UO_1878 (O_1878,N_19836,N_19975);
nor UO_1879 (O_1879,N_19826,N_19961);
nand UO_1880 (O_1880,N_19906,N_19990);
xor UO_1881 (O_1881,N_19810,N_19751);
and UO_1882 (O_1882,N_19926,N_19922);
or UO_1883 (O_1883,N_19946,N_19853);
nand UO_1884 (O_1884,N_19984,N_19935);
nor UO_1885 (O_1885,N_19892,N_19931);
or UO_1886 (O_1886,N_19756,N_19909);
xor UO_1887 (O_1887,N_19791,N_19917);
nor UO_1888 (O_1888,N_19886,N_19888);
nand UO_1889 (O_1889,N_19874,N_19808);
or UO_1890 (O_1890,N_19802,N_19942);
or UO_1891 (O_1891,N_19778,N_19787);
nor UO_1892 (O_1892,N_19864,N_19776);
and UO_1893 (O_1893,N_19779,N_19977);
and UO_1894 (O_1894,N_19835,N_19987);
nor UO_1895 (O_1895,N_19806,N_19876);
nor UO_1896 (O_1896,N_19957,N_19868);
xor UO_1897 (O_1897,N_19967,N_19760);
nor UO_1898 (O_1898,N_19794,N_19860);
and UO_1899 (O_1899,N_19966,N_19870);
and UO_1900 (O_1900,N_19918,N_19754);
nand UO_1901 (O_1901,N_19995,N_19773);
or UO_1902 (O_1902,N_19943,N_19881);
xnor UO_1903 (O_1903,N_19801,N_19965);
and UO_1904 (O_1904,N_19846,N_19872);
or UO_1905 (O_1905,N_19899,N_19993);
nor UO_1906 (O_1906,N_19895,N_19789);
or UO_1907 (O_1907,N_19982,N_19916);
nand UO_1908 (O_1908,N_19792,N_19931);
nor UO_1909 (O_1909,N_19768,N_19992);
and UO_1910 (O_1910,N_19928,N_19952);
nor UO_1911 (O_1911,N_19860,N_19962);
and UO_1912 (O_1912,N_19755,N_19776);
xnor UO_1913 (O_1913,N_19933,N_19863);
or UO_1914 (O_1914,N_19926,N_19901);
nor UO_1915 (O_1915,N_19771,N_19787);
or UO_1916 (O_1916,N_19847,N_19871);
nand UO_1917 (O_1917,N_19778,N_19831);
nand UO_1918 (O_1918,N_19791,N_19896);
and UO_1919 (O_1919,N_19802,N_19879);
and UO_1920 (O_1920,N_19849,N_19823);
nand UO_1921 (O_1921,N_19772,N_19985);
and UO_1922 (O_1922,N_19895,N_19860);
and UO_1923 (O_1923,N_19929,N_19943);
xor UO_1924 (O_1924,N_19977,N_19947);
nand UO_1925 (O_1925,N_19810,N_19830);
and UO_1926 (O_1926,N_19917,N_19920);
nor UO_1927 (O_1927,N_19817,N_19794);
and UO_1928 (O_1928,N_19905,N_19786);
or UO_1929 (O_1929,N_19792,N_19860);
or UO_1930 (O_1930,N_19880,N_19884);
and UO_1931 (O_1931,N_19755,N_19852);
and UO_1932 (O_1932,N_19822,N_19944);
nor UO_1933 (O_1933,N_19978,N_19936);
nor UO_1934 (O_1934,N_19940,N_19996);
or UO_1935 (O_1935,N_19809,N_19763);
nand UO_1936 (O_1936,N_19961,N_19839);
nand UO_1937 (O_1937,N_19852,N_19953);
xor UO_1938 (O_1938,N_19939,N_19855);
xor UO_1939 (O_1939,N_19969,N_19935);
and UO_1940 (O_1940,N_19794,N_19806);
xnor UO_1941 (O_1941,N_19789,N_19758);
nand UO_1942 (O_1942,N_19928,N_19907);
xor UO_1943 (O_1943,N_19915,N_19953);
or UO_1944 (O_1944,N_19970,N_19956);
nand UO_1945 (O_1945,N_19923,N_19904);
nand UO_1946 (O_1946,N_19944,N_19775);
or UO_1947 (O_1947,N_19752,N_19907);
nand UO_1948 (O_1948,N_19797,N_19905);
nor UO_1949 (O_1949,N_19816,N_19815);
xor UO_1950 (O_1950,N_19801,N_19858);
xnor UO_1951 (O_1951,N_19796,N_19946);
nand UO_1952 (O_1952,N_19961,N_19930);
nand UO_1953 (O_1953,N_19882,N_19847);
nor UO_1954 (O_1954,N_19958,N_19802);
and UO_1955 (O_1955,N_19907,N_19790);
or UO_1956 (O_1956,N_19823,N_19984);
nor UO_1957 (O_1957,N_19881,N_19763);
xnor UO_1958 (O_1958,N_19924,N_19756);
and UO_1959 (O_1959,N_19756,N_19917);
nor UO_1960 (O_1960,N_19818,N_19792);
nor UO_1961 (O_1961,N_19978,N_19994);
and UO_1962 (O_1962,N_19816,N_19880);
and UO_1963 (O_1963,N_19765,N_19791);
nand UO_1964 (O_1964,N_19811,N_19944);
nand UO_1965 (O_1965,N_19751,N_19937);
nor UO_1966 (O_1966,N_19848,N_19761);
xnor UO_1967 (O_1967,N_19961,N_19850);
or UO_1968 (O_1968,N_19887,N_19826);
nor UO_1969 (O_1969,N_19873,N_19755);
nor UO_1970 (O_1970,N_19935,N_19995);
or UO_1971 (O_1971,N_19771,N_19942);
and UO_1972 (O_1972,N_19954,N_19801);
and UO_1973 (O_1973,N_19787,N_19921);
nor UO_1974 (O_1974,N_19853,N_19838);
xnor UO_1975 (O_1975,N_19876,N_19877);
nand UO_1976 (O_1976,N_19848,N_19980);
nand UO_1977 (O_1977,N_19930,N_19770);
and UO_1978 (O_1978,N_19969,N_19940);
nand UO_1979 (O_1979,N_19908,N_19979);
or UO_1980 (O_1980,N_19802,N_19849);
nand UO_1981 (O_1981,N_19832,N_19879);
or UO_1982 (O_1982,N_19928,N_19801);
and UO_1983 (O_1983,N_19963,N_19827);
xor UO_1984 (O_1984,N_19906,N_19775);
nor UO_1985 (O_1985,N_19939,N_19807);
or UO_1986 (O_1986,N_19832,N_19814);
and UO_1987 (O_1987,N_19956,N_19808);
xnor UO_1988 (O_1988,N_19940,N_19921);
xor UO_1989 (O_1989,N_19819,N_19777);
and UO_1990 (O_1990,N_19972,N_19874);
nor UO_1991 (O_1991,N_19968,N_19970);
or UO_1992 (O_1992,N_19924,N_19993);
xor UO_1993 (O_1993,N_19881,N_19915);
and UO_1994 (O_1994,N_19932,N_19782);
nor UO_1995 (O_1995,N_19952,N_19809);
nand UO_1996 (O_1996,N_19963,N_19943);
or UO_1997 (O_1997,N_19787,N_19956);
and UO_1998 (O_1998,N_19821,N_19914);
nand UO_1999 (O_1999,N_19956,N_19918);
xor UO_2000 (O_2000,N_19761,N_19921);
or UO_2001 (O_2001,N_19756,N_19971);
or UO_2002 (O_2002,N_19791,N_19996);
or UO_2003 (O_2003,N_19886,N_19782);
xnor UO_2004 (O_2004,N_19969,N_19898);
nor UO_2005 (O_2005,N_19808,N_19954);
nand UO_2006 (O_2006,N_19770,N_19795);
and UO_2007 (O_2007,N_19996,N_19848);
or UO_2008 (O_2008,N_19925,N_19955);
or UO_2009 (O_2009,N_19905,N_19919);
xor UO_2010 (O_2010,N_19888,N_19887);
xnor UO_2011 (O_2011,N_19851,N_19900);
xnor UO_2012 (O_2012,N_19899,N_19751);
and UO_2013 (O_2013,N_19941,N_19769);
nand UO_2014 (O_2014,N_19782,N_19754);
and UO_2015 (O_2015,N_19987,N_19992);
nor UO_2016 (O_2016,N_19921,N_19842);
or UO_2017 (O_2017,N_19973,N_19975);
nor UO_2018 (O_2018,N_19981,N_19859);
nor UO_2019 (O_2019,N_19843,N_19969);
or UO_2020 (O_2020,N_19931,N_19928);
nand UO_2021 (O_2021,N_19924,N_19858);
or UO_2022 (O_2022,N_19968,N_19790);
nand UO_2023 (O_2023,N_19994,N_19879);
or UO_2024 (O_2024,N_19848,N_19818);
or UO_2025 (O_2025,N_19999,N_19782);
nand UO_2026 (O_2026,N_19768,N_19923);
nor UO_2027 (O_2027,N_19959,N_19806);
nand UO_2028 (O_2028,N_19809,N_19856);
nand UO_2029 (O_2029,N_19958,N_19967);
nor UO_2030 (O_2030,N_19758,N_19762);
or UO_2031 (O_2031,N_19788,N_19750);
nor UO_2032 (O_2032,N_19757,N_19868);
or UO_2033 (O_2033,N_19926,N_19918);
nor UO_2034 (O_2034,N_19817,N_19841);
nand UO_2035 (O_2035,N_19961,N_19802);
and UO_2036 (O_2036,N_19771,N_19780);
nor UO_2037 (O_2037,N_19949,N_19963);
or UO_2038 (O_2038,N_19941,N_19916);
nand UO_2039 (O_2039,N_19811,N_19777);
and UO_2040 (O_2040,N_19751,N_19779);
nor UO_2041 (O_2041,N_19832,N_19982);
or UO_2042 (O_2042,N_19798,N_19797);
nor UO_2043 (O_2043,N_19917,N_19983);
nor UO_2044 (O_2044,N_19842,N_19764);
xnor UO_2045 (O_2045,N_19958,N_19888);
nand UO_2046 (O_2046,N_19860,N_19797);
xor UO_2047 (O_2047,N_19925,N_19928);
or UO_2048 (O_2048,N_19788,N_19934);
nor UO_2049 (O_2049,N_19873,N_19866);
nand UO_2050 (O_2050,N_19758,N_19874);
or UO_2051 (O_2051,N_19844,N_19916);
or UO_2052 (O_2052,N_19839,N_19807);
and UO_2053 (O_2053,N_19829,N_19975);
nor UO_2054 (O_2054,N_19924,N_19871);
and UO_2055 (O_2055,N_19846,N_19989);
or UO_2056 (O_2056,N_19970,N_19937);
xor UO_2057 (O_2057,N_19948,N_19936);
nor UO_2058 (O_2058,N_19881,N_19871);
nor UO_2059 (O_2059,N_19887,N_19795);
xor UO_2060 (O_2060,N_19850,N_19996);
xor UO_2061 (O_2061,N_19854,N_19774);
xnor UO_2062 (O_2062,N_19892,N_19945);
or UO_2063 (O_2063,N_19976,N_19879);
nand UO_2064 (O_2064,N_19869,N_19967);
nor UO_2065 (O_2065,N_19983,N_19823);
xor UO_2066 (O_2066,N_19931,N_19847);
xnor UO_2067 (O_2067,N_19762,N_19823);
and UO_2068 (O_2068,N_19901,N_19999);
or UO_2069 (O_2069,N_19753,N_19768);
or UO_2070 (O_2070,N_19798,N_19768);
or UO_2071 (O_2071,N_19751,N_19830);
and UO_2072 (O_2072,N_19820,N_19785);
and UO_2073 (O_2073,N_19779,N_19948);
xor UO_2074 (O_2074,N_19958,N_19856);
nand UO_2075 (O_2075,N_19964,N_19856);
or UO_2076 (O_2076,N_19858,N_19871);
nand UO_2077 (O_2077,N_19858,N_19915);
nor UO_2078 (O_2078,N_19856,N_19828);
or UO_2079 (O_2079,N_19917,N_19928);
nor UO_2080 (O_2080,N_19922,N_19976);
or UO_2081 (O_2081,N_19779,N_19858);
and UO_2082 (O_2082,N_19909,N_19841);
or UO_2083 (O_2083,N_19969,N_19903);
nand UO_2084 (O_2084,N_19870,N_19878);
nor UO_2085 (O_2085,N_19775,N_19752);
and UO_2086 (O_2086,N_19970,N_19885);
or UO_2087 (O_2087,N_19853,N_19977);
xor UO_2088 (O_2088,N_19992,N_19970);
xnor UO_2089 (O_2089,N_19830,N_19988);
xnor UO_2090 (O_2090,N_19832,N_19811);
xor UO_2091 (O_2091,N_19955,N_19808);
nand UO_2092 (O_2092,N_19900,N_19778);
and UO_2093 (O_2093,N_19756,N_19842);
xnor UO_2094 (O_2094,N_19873,N_19917);
xor UO_2095 (O_2095,N_19879,N_19991);
or UO_2096 (O_2096,N_19807,N_19991);
nor UO_2097 (O_2097,N_19912,N_19968);
xor UO_2098 (O_2098,N_19937,N_19906);
xor UO_2099 (O_2099,N_19796,N_19925);
nor UO_2100 (O_2100,N_19785,N_19965);
or UO_2101 (O_2101,N_19921,N_19954);
nor UO_2102 (O_2102,N_19864,N_19785);
or UO_2103 (O_2103,N_19907,N_19793);
and UO_2104 (O_2104,N_19954,N_19869);
or UO_2105 (O_2105,N_19959,N_19915);
nand UO_2106 (O_2106,N_19863,N_19842);
or UO_2107 (O_2107,N_19929,N_19867);
and UO_2108 (O_2108,N_19932,N_19964);
nand UO_2109 (O_2109,N_19821,N_19854);
or UO_2110 (O_2110,N_19996,N_19936);
and UO_2111 (O_2111,N_19848,N_19786);
xnor UO_2112 (O_2112,N_19830,N_19783);
nand UO_2113 (O_2113,N_19794,N_19855);
and UO_2114 (O_2114,N_19972,N_19813);
and UO_2115 (O_2115,N_19987,N_19753);
or UO_2116 (O_2116,N_19941,N_19781);
or UO_2117 (O_2117,N_19954,N_19977);
nor UO_2118 (O_2118,N_19886,N_19958);
or UO_2119 (O_2119,N_19849,N_19992);
nand UO_2120 (O_2120,N_19939,N_19833);
nor UO_2121 (O_2121,N_19881,N_19751);
nor UO_2122 (O_2122,N_19882,N_19906);
and UO_2123 (O_2123,N_19758,N_19981);
nand UO_2124 (O_2124,N_19908,N_19875);
or UO_2125 (O_2125,N_19892,N_19950);
nor UO_2126 (O_2126,N_19974,N_19781);
xor UO_2127 (O_2127,N_19820,N_19996);
nand UO_2128 (O_2128,N_19787,N_19904);
nor UO_2129 (O_2129,N_19845,N_19936);
or UO_2130 (O_2130,N_19962,N_19981);
or UO_2131 (O_2131,N_19901,N_19931);
or UO_2132 (O_2132,N_19781,N_19896);
nand UO_2133 (O_2133,N_19936,N_19995);
and UO_2134 (O_2134,N_19988,N_19949);
xnor UO_2135 (O_2135,N_19949,N_19896);
nor UO_2136 (O_2136,N_19996,N_19935);
nor UO_2137 (O_2137,N_19873,N_19950);
or UO_2138 (O_2138,N_19800,N_19942);
xor UO_2139 (O_2139,N_19752,N_19784);
nor UO_2140 (O_2140,N_19782,N_19874);
nor UO_2141 (O_2141,N_19997,N_19983);
nor UO_2142 (O_2142,N_19827,N_19855);
and UO_2143 (O_2143,N_19897,N_19966);
nand UO_2144 (O_2144,N_19843,N_19788);
nand UO_2145 (O_2145,N_19760,N_19977);
nand UO_2146 (O_2146,N_19823,N_19955);
nand UO_2147 (O_2147,N_19881,N_19961);
nand UO_2148 (O_2148,N_19887,N_19837);
xor UO_2149 (O_2149,N_19879,N_19873);
nor UO_2150 (O_2150,N_19887,N_19910);
nand UO_2151 (O_2151,N_19986,N_19856);
and UO_2152 (O_2152,N_19820,N_19919);
or UO_2153 (O_2153,N_19881,N_19820);
or UO_2154 (O_2154,N_19787,N_19914);
and UO_2155 (O_2155,N_19784,N_19950);
or UO_2156 (O_2156,N_19756,N_19869);
xnor UO_2157 (O_2157,N_19765,N_19991);
or UO_2158 (O_2158,N_19769,N_19965);
or UO_2159 (O_2159,N_19975,N_19877);
xnor UO_2160 (O_2160,N_19850,N_19977);
and UO_2161 (O_2161,N_19967,N_19773);
xor UO_2162 (O_2162,N_19964,N_19822);
and UO_2163 (O_2163,N_19998,N_19983);
xnor UO_2164 (O_2164,N_19865,N_19848);
and UO_2165 (O_2165,N_19976,N_19955);
nor UO_2166 (O_2166,N_19825,N_19835);
and UO_2167 (O_2167,N_19811,N_19860);
xnor UO_2168 (O_2168,N_19756,N_19929);
or UO_2169 (O_2169,N_19828,N_19913);
and UO_2170 (O_2170,N_19754,N_19778);
or UO_2171 (O_2171,N_19963,N_19769);
or UO_2172 (O_2172,N_19776,N_19847);
xor UO_2173 (O_2173,N_19768,N_19983);
and UO_2174 (O_2174,N_19947,N_19905);
nor UO_2175 (O_2175,N_19833,N_19888);
or UO_2176 (O_2176,N_19968,N_19947);
or UO_2177 (O_2177,N_19976,N_19897);
and UO_2178 (O_2178,N_19847,N_19788);
or UO_2179 (O_2179,N_19917,N_19954);
nor UO_2180 (O_2180,N_19862,N_19938);
and UO_2181 (O_2181,N_19961,N_19833);
nor UO_2182 (O_2182,N_19833,N_19750);
xor UO_2183 (O_2183,N_19849,N_19860);
nor UO_2184 (O_2184,N_19957,N_19950);
nor UO_2185 (O_2185,N_19861,N_19760);
nand UO_2186 (O_2186,N_19801,N_19892);
or UO_2187 (O_2187,N_19783,N_19782);
xor UO_2188 (O_2188,N_19896,N_19977);
and UO_2189 (O_2189,N_19956,N_19946);
or UO_2190 (O_2190,N_19861,N_19871);
and UO_2191 (O_2191,N_19996,N_19909);
and UO_2192 (O_2192,N_19949,N_19793);
or UO_2193 (O_2193,N_19779,N_19842);
nor UO_2194 (O_2194,N_19898,N_19781);
or UO_2195 (O_2195,N_19849,N_19751);
xnor UO_2196 (O_2196,N_19828,N_19976);
nand UO_2197 (O_2197,N_19935,N_19966);
xnor UO_2198 (O_2198,N_19893,N_19919);
xnor UO_2199 (O_2199,N_19911,N_19771);
or UO_2200 (O_2200,N_19879,N_19920);
nor UO_2201 (O_2201,N_19880,N_19961);
and UO_2202 (O_2202,N_19883,N_19794);
and UO_2203 (O_2203,N_19930,N_19844);
nor UO_2204 (O_2204,N_19999,N_19761);
and UO_2205 (O_2205,N_19881,N_19960);
or UO_2206 (O_2206,N_19860,N_19957);
xor UO_2207 (O_2207,N_19934,N_19858);
xnor UO_2208 (O_2208,N_19925,N_19965);
and UO_2209 (O_2209,N_19806,N_19853);
nor UO_2210 (O_2210,N_19772,N_19891);
xor UO_2211 (O_2211,N_19862,N_19971);
nor UO_2212 (O_2212,N_19992,N_19858);
and UO_2213 (O_2213,N_19987,N_19925);
and UO_2214 (O_2214,N_19828,N_19774);
and UO_2215 (O_2215,N_19970,N_19806);
or UO_2216 (O_2216,N_19892,N_19955);
or UO_2217 (O_2217,N_19831,N_19807);
or UO_2218 (O_2218,N_19925,N_19976);
and UO_2219 (O_2219,N_19762,N_19934);
and UO_2220 (O_2220,N_19752,N_19908);
nand UO_2221 (O_2221,N_19880,N_19805);
nor UO_2222 (O_2222,N_19860,N_19870);
or UO_2223 (O_2223,N_19774,N_19755);
nor UO_2224 (O_2224,N_19974,N_19765);
or UO_2225 (O_2225,N_19775,N_19774);
xnor UO_2226 (O_2226,N_19755,N_19949);
and UO_2227 (O_2227,N_19794,N_19773);
nand UO_2228 (O_2228,N_19818,N_19989);
nor UO_2229 (O_2229,N_19980,N_19989);
or UO_2230 (O_2230,N_19949,N_19918);
xor UO_2231 (O_2231,N_19986,N_19911);
nor UO_2232 (O_2232,N_19912,N_19876);
nand UO_2233 (O_2233,N_19879,N_19794);
nor UO_2234 (O_2234,N_19858,N_19985);
xnor UO_2235 (O_2235,N_19928,N_19826);
and UO_2236 (O_2236,N_19842,N_19902);
nor UO_2237 (O_2237,N_19867,N_19765);
or UO_2238 (O_2238,N_19797,N_19945);
and UO_2239 (O_2239,N_19871,N_19768);
nand UO_2240 (O_2240,N_19774,N_19916);
nor UO_2241 (O_2241,N_19914,N_19800);
or UO_2242 (O_2242,N_19978,N_19843);
xnor UO_2243 (O_2243,N_19799,N_19842);
nor UO_2244 (O_2244,N_19883,N_19816);
or UO_2245 (O_2245,N_19862,N_19802);
xnor UO_2246 (O_2246,N_19957,N_19829);
nor UO_2247 (O_2247,N_19850,N_19889);
nand UO_2248 (O_2248,N_19926,N_19870);
or UO_2249 (O_2249,N_19751,N_19750);
and UO_2250 (O_2250,N_19779,N_19966);
xnor UO_2251 (O_2251,N_19888,N_19905);
nor UO_2252 (O_2252,N_19972,N_19871);
and UO_2253 (O_2253,N_19877,N_19848);
xor UO_2254 (O_2254,N_19815,N_19757);
nor UO_2255 (O_2255,N_19962,N_19807);
nand UO_2256 (O_2256,N_19827,N_19965);
or UO_2257 (O_2257,N_19938,N_19916);
xnor UO_2258 (O_2258,N_19808,N_19885);
nand UO_2259 (O_2259,N_19961,N_19796);
or UO_2260 (O_2260,N_19792,N_19758);
xor UO_2261 (O_2261,N_19757,N_19765);
and UO_2262 (O_2262,N_19816,N_19862);
or UO_2263 (O_2263,N_19759,N_19996);
or UO_2264 (O_2264,N_19966,N_19956);
and UO_2265 (O_2265,N_19848,N_19788);
nor UO_2266 (O_2266,N_19842,N_19795);
nor UO_2267 (O_2267,N_19899,N_19970);
or UO_2268 (O_2268,N_19864,N_19781);
nand UO_2269 (O_2269,N_19780,N_19772);
or UO_2270 (O_2270,N_19867,N_19954);
nand UO_2271 (O_2271,N_19959,N_19763);
xor UO_2272 (O_2272,N_19907,N_19937);
nor UO_2273 (O_2273,N_19783,N_19967);
and UO_2274 (O_2274,N_19963,N_19763);
or UO_2275 (O_2275,N_19799,N_19941);
xor UO_2276 (O_2276,N_19853,N_19811);
xnor UO_2277 (O_2277,N_19844,N_19843);
xnor UO_2278 (O_2278,N_19900,N_19936);
or UO_2279 (O_2279,N_19813,N_19906);
nand UO_2280 (O_2280,N_19974,N_19874);
or UO_2281 (O_2281,N_19795,N_19998);
or UO_2282 (O_2282,N_19817,N_19769);
or UO_2283 (O_2283,N_19852,N_19984);
xor UO_2284 (O_2284,N_19936,N_19934);
nand UO_2285 (O_2285,N_19751,N_19803);
nor UO_2286 (O_2286,N_19903,N_19779);
nor UO_2287 (O_2287,N_19881,N_19938);
or UO_2288 (O_2288,N_19894,N_19750);
or UO_2289 (O_2289,N_19821,N_19865);
nor UO_2290 (O_2290,N_19969,N_19776);
and UO_2291 (O_2291,N_19973,N_19964);
nor UO_2292 (O_2292,N_19793,N_19966);
or UO_2293 (O_2293,N_19973,N_19800);
or UO_2294 (O_2294,N_19785,N_19954);
xnor UO_2295 (O_2295,N_19900,N_19970);
or UO_2296 (O_2296,N_19786,N_19991);
and UO_2297 (O_2297,N_19868,N_19756);
nand UO_2298 (O_2298,N_19852,N_19831);
nand UO_2299 (O_2299,N_19912,N_19879);
or UO_2300 (O_2300,N_19854,N_19879);
and UO_2301 (O_2301,N_19781,N_19851);
and UO_2302 (O_2302,N_19895,N_19801);
and UO_2303 (O_2303,N_19911,N_19776);
nand UO_2304 (O_2304,N_19773,N_19991);
xnor UO_2305 (O_2305,N_19818,N_19830);
and UO_2306 (O_2306,N_19971,N_19834);
and UO_2307 (O_2307,N_19902,N_19769);
nor UO_2308 (O_2308,N_19973,N_19896);
nand UO_2309 (O_2309,N_19868,N_19993);
or UO_2310 (O_2310,N_19801,N_19867);
nand UO_2311 (O_2311,N_19799,N_19991);
nor UO_2312 (O_2312,N_19772,N_19890);
nor UO_2313 (O_2313,N_19851,N_19854);
or UO_2314 (O_2314,N_19935,N_19856);
nand UO_2315 (O_2315,N_19960,N_19805);
xor UO_2316 (O_2316,N_19865,N_19926);
or UO_2317 (O_2317,N_19963,N_19828);
xor UO_2318 (O_2318,N_19985,N_19853);
xnor UO_2319 (O_2319,N_19876,N_19786);
xnor UO_2320 (O_2320,N_19931,N_19752);
and UO_2321 (O_2321,N_19963,N_19961);
nand UO_2322 (O_2322,N_19997,N_19787);
nor UO_2323 (O_2323,N_19771,N_19887);
xnor UO_2324 (O_2324,N_19856,N_19995);
nor UO_2325 (O_2325,N_19994,N_19937);
and UO_2326 (O_2326,N_19806,N_19942);
and UO_2327 (O_2327,N_19936,N_19932);
and UO_2328 (O_2328,N_19846,N_19991);
or UO_2329 (O_2329,N_19884,N_19753);
and UO_2330 (O_2330,N_19915,N_19865);
and UO_2331 (O_2331,N_19760,N_19838);
and UO_2332 (O_2332,N_19845,N_19916);
nand UO_2333 (O_2333,N_19980,N_19913);
nor UO_2334 (O_2334,N_19768,N_19754);
or UO_2335 (O_2335,N_19895,N_19949);
and UO_2336 (O_2336,N_19877,N_19927);
xnor UO_2337 (O_2337,N_19791,N_19929);
nor UO_2338 (O_2338,N_19919,N_19876);
xor UO_2339 (O_2339,N_19939,N_19872);
nor UO_2340 (O_2340,N_19846,N_19779);
nand UO_2341 (O_2341,N_19923,N_19839);
and UO_2342 (O_2342,N_19924,N_19906);
nand UO_2343 (O_2343,N_19835,N_19785);
xor UO_2344 (O_2344,N_19972,N_19987);
or UO_2345 (O_2345,N_19910,N_19875);
xnor UO_2346 (O_2346,N_19812,N_19972);
nand UO_2347 (O_2347,N_19955,N_19959);
and UO_2348 (O_2348,N_19921,N_19859);
nand UO_2349 (O_2349,N_19887,N_19878);
or UO_2350 (O_2350,N_19944,N_19758);
xor UO_2351 (O_2351,N_19986,N_19777);
and UO_2352 (O_2352,N_19858,N_19990);
and UO_2353 (O_2353,N_19979,N_19921);
or UO_2354 (O_2354,N_19773,N_19916);
xnor UO_2355 (O_2355,N_19959,N_19757);
nor UO_2356 (O_2356,N_19759,N_19804);
or UO_2357 (O_2357,N_19963,N_19817);
or UO_2358 (O_2358,N_19808,N_19891);
or UO_2359 (O_2359,N_19958,N_19997);
or UO_2360 (O_2360,N_19879,N_19781);
and UO_2361 (O_2361,N_19971,N_19782);
nor UO_2362 (O_2362,N_19966,N_19949);
nor UO_2363 (O_2363,N_19855,N_19932);
xnor UO_2364 (O_2364,N_19911,N_19958);
or UO_2365 (O_2365,N_19979,N_19885);
and UO_2366 (O_2366,N_19897,N_19835);
nand UO_2367 (O_2367,N_19943,N_19786);
and UO_2368 (O_2368,N_19779,N_19772);
nand UO_2369 (O_2369,N_19903,N_19791);
nand UO_2370 (O_2370,N_19774,N_19888);
and UO_2371 (O_2371,N_19804,N_19752);
nand UO_2372 (O_2372,N_19945,N_19948);
nor UO_2373 (O_2373,N_19975,N_19874);
nor UO_2374 (O_2374,N_19785,N_19976);
nor UO_2375 (O_2375,N_19862,N_19822);
nand UO_2376 (O_2376,N_19870,N_19887);
nor UO_2377 (O_2377,N_19836,N_19991);
nor UO_2378 (O_2378,N_19856,N_19781);
xor UO_2379 (O_2379,N_19951,N_19773);
nor UO_2380 (O_2380,N_19864,N_19822);
nor UO_2381 (O_2381,N_19988,N_19840);
or UO_2382 (O_2382,N_19807,N_19835);
nand UO_2383 (O_2383,N_19909,N_19883);
xor UO_2384 (O_2384,N_19920,N_19824);
nand UO_2385 (O_2385,N_19903,N_19850);
nand UO_2386 (O_2386,N_19991,N_19921);
xor UO_2387 (O_2387,N_19870,N_19786);
nor UO_2388 (O_2388,N_19907,N_19814);
xor UO_2389 (O_2389,N_19814,N_19943);
or UO_2390 (O_2390,N_19808,N_19866);
xor UO_2391 (O_2391,N_19810,N_19939);
nor UO_2392 (O_2392,N_19991,N_19875);
xnor UO_2393 (O_2393,N_19799,N_19801);
nor UO_2394 (O_2394,N_19968,N_19901);
xor UO_2395 (O_2395,N_19806,N_19821);
or UO_2396 (O_2396,N_19874,N_19978);
nand UO_2397 (O_2397,N_19822,N_19997);
or UO_2398 (O_2398,N_19807,N_19812);
and UO_2399 (O_2399,N_19930,N_19756);
and UO_2400 (O_2400,N_19753,N_19883);
nor UO_2401 (O_2401,N_19814,N_19845);
nand UO_2402 (O_2402,N_19791,N_19863);
nand UO_2403 (O_2403,N_19832,N_19826);
xnor UO_2404 (O_2404,N_19769,N_19890);
nand UO_2405 (O_2405,N_19962,N_19819);
or UO_2406 (O_2406,N_19843,N_19888);
or UO_2407 (O_2407,N_19779,N_19797);
nand UO_2408 (O_2408,N_19950,N_19884);
nor UO_2409 (O_2409,N_19979,N_19825);
nor UO_2410 (O_2410,N_19921,N_19827);
nand UO_2411 (O_2411,N_19800,N_19843);
or UO_2412 (O_2412,N_19840,N_19764);
xor UO_2413 (O_2413,N_19806,N_19941);
and UO_2414 (O_2414,N_19870,N_19848);
xnor UO_2415 (O_2415,N_19828,N_19946);
and UO_2416 (O_2416,N_19801,N_19914);
nand UO_2417 (O_2417,N_19778,N_19881);
xor UO_2418 (O_2418,N_19752,N_19862);
nor UO_2419 (O_2419,N_19856,N_19754);
nor UO_2420 (O_2420,N_19974,N_19809);
and UO_2421 (O_2421,N_19752,N_19950);
xor UO_2422 (O_2422,N_19983,N_19827);
and UO_2423 (O_2423,N_19895,N_19943);
or UO_2424 (O_2424,N_19878,N_19804);
nand UO_2425 (O_2425,N_19948,N_19968);
or UO_2426 (O_2426,N_19826,N_19831);
xor UO_2427 (O_2427,N_19760,N_19802);
and UO_2428 (O_2428,N_19825,N_19790);
nand UO_2429 (O_2429,N_19774,N_19920);
or UO_2430 (O_2430,N_19900,N_19774);
xnor UO_2431 (O_2431,N_19919,N_19864);
nand UO_2432 (O_2432,N_19858,N_19847);
nand UO_2433 (O_2433,N_19859,N_19874);
xor UO_2434 (O_2434,N_19890,N_19930);
xnor UO_2435 (O_2435,N_19781,N_19762);
xor UO_2436 (O_2436,N_19958,N_19861);
nor UO_2437 (O_2437,N_19794,N_19779);
and UO_2438 (O_2438,N_19979,N_19986);
and UO_2439 (O_2439,N_19753,N_19842);
nand UO_2440 (O_2440,N_19752,N_19882);
xnor UO_2441 (O_2441,N_19852,N_19919);
nand UO_2442 (O_2442,N_19965,N_19938);
or UO_2443 (O_2443,N_19920,N_19835);
xor UO_2444 (O_2444,N_19849,N_19814);
nor UO_2445 (O_2445,N_19969,N_19779);
xor UO_2446 (O_2446,N_19878,N_19805);
and UO_2447 (O_2447,N_19945,N_19982);
nor UO_2448 (O_2448,N_19868,N_19830);
xor UO_2449 (O_2449,N_19972,N_19920);
and UO_2450 (O_2450,N_19833,N_19881);
nand UO_2451 (O_2451,N_19815,N_19834);
xnor UO_2452 (O_2452,N_19821,N_19939);
or UO_2453 (O_2453,N_19835,N_19818);
nand UO_2454 (O_2454,N_19789,N_19872);
nand UO_2455 (O_2455,N_19933,N_19757);
nor UO_2456 (O_2456,N_19790,N_19930);
or UO_2457 (O_2457,N_19797,N_19970);
xor UO_2458 (O_2458,N_19923,N_19973);
xnor UO_2459 (O_2459,N_19934,N_19852);
nor UO_2460 (O_2460,N_19759,N_19979);
xnor UO_2461 (O_2461,N_19948,N_19807);
or UO_2462 (O_2462,N_19800,N_19845);
nor UO_2463 (O_2463,N_19840,N_19870);
nand UO_2464 (O_2464,N_19868,N_19754);
xor UO_2465 (O_2465,N_19754,N_19987);
and UO_2466 (O_2466,N_19798,N_19844);
xnor UO_2467 (O_2467,N_19959,N_19909);
nand UO_2468 (O_2468,N_19959,N_19861);
nor UO_2469 (O_2469,N_19779,N_19874);
xor UO_2470 (O_2470,N_19991,N_19979);
and UO_2471 (O_2471,N_19804,N_19761);
xor UO_2472 (O_2472,N_19902,N_19782);
nand UO_2473 (O_2473,N_19918,N_19948);
nand UO_2474 (O_2474,N_19954,N_19996);
or UO_2475 (O_2475,N_19922,N_19987);
or UO_2476 (O_2476,N_19843,N_19833);
or UO_2477 (O_2477,N_19787,N_19793);
and UO_2478 (O_2478,N_19878,N_19888);
and UO_2479 (O_2479,N_19780,N_19969);
nor UO_2480 (O_2480,N_19980,N_19897);
nor UO_2481 (O_2481,N_19766,N_19990);
or UO_2482 (O_2482,N_19986,N_19803);
xnor UO_2483 (O_2483,N_19908,N_19968);
or UO_2484 (O_2484,N_19751,N_19948);
nand UO_2485 (O_2485,N_19823,N_19870);
or UO_2486 (O_2486,N_19874,N_19995);
and UO_2487 (O_2487,N_19758,N_19937);
nor UO_2488 (O_2488,N_19873,N_19962);
xor UO_2489 (O_2489,N_19966,N_19927);
or UO_2490 (O_2490,N_19930,N_19772);
nor UO_2491 (O_2491,N_19938,N_19863);
nor UO_2492 (O_2492,N_19783,N_19873);
nand UO_2493 (O_2493,N_19777,N_19859);
xor UO_2494 (O_2494,N_19824,N_19923);
and UO_2495 (O_2495,N_19907,N_19903);
nand UO_2496 (O_2496,N_19889,N_19812);
nand UO_2497 (O_2497,N_19937,N_19980);
nor UO_2498 (O_2498,N_19831,N_19900);
nand UO_2499 (O_2499,N_19820,N_19821);
endmodule